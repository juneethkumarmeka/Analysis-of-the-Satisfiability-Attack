module basic_2000_20000_2500_4_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1030,In_1878);
and U1 (N_1,In_1120,In_917);
nor U2 (N_2,In_831,In_1440);
xor U3 (N_3,In_1840,In_1885);
and U4 (N_4,In_1527,In_372);
nor U5 (N_5,In_1017,In_252);
and U6 (N_6,In_745,In_1753);
nand U7 (N_7,In_1538,In_120);
nor U8 (N_8,In_1430,In_1323);
or U9 (N_9,In_1646,In_1478);
or U10 (N_10,In_223,In_1250);
xor U11 (N_11,In_933,In_1916);
or U12 (N_12,In_1855,In_313);
nand U13 (N_13,In_692,In_610);
nand U14 (N_14,In_337,In_1812);
nor U15 (N_15,In_1044,In_44);
or U16 (N_16,In_1881,In_536);
nor U17 (N_17,In_825,In_57);
or U18 (N_18,In_1827,In_1273);
xor U19 (N_19,In_909,In_1787);
nor U20 (N_20,In_843,In_998);
nor U21 (N_21,In_1870,In_1903);
or U22 (N_22,In_226,In_432);
and U23 (N_23,In_1856,In_1589);
xor U24 (N_24,In_817,In_152);
nor U25 (N_25,In_1052,In_1462);
nand U26 (N_26,In_781,In_1637);
and U27 (N_27,In_1691,In_1800);
nand U28 (N_28,In_1936,In_377);
and U29 (N_29,In_1111,In_819);
or U30 (N_30,In_486,In_161);
xnor U31 (N_31,In_117,In_1858);
and U32 (N_32,In_670,In_1002);
xnor U33 (N_33,In_30,In_204);
nor U34 (N_34,In_724,In_450);
nand U35 (N_35,In_1288,In_1399);
and U36 (N_36,In_1846,In_904);
or U37 (N_37,In_119,In_701);
nor U38 (N_38,In_466,In_62);
or U39 (N_39,In_139,In_1785);
and U40 (N_40,In_560,In_227);
or U41 (N_41,In_1365,In_1619);
nand U42 (N_42,In_45,In_1295);
nor U43 (N_43,In_425,In_416);
nand U44 (N_44,In_13,In_894);
xor U45 (N_45,In_1270,In_690);
nand U46 (N_46,In_926,In_1229);
nor U47 (N_47,In_1919,In_1978);
nand U48 (N_48,In_1027,In_1436);
or U49 (N_49,In_1915,In_1359);
xor U50 (N_50,In_1743,In_746);
and U51 (N_51,In_1501,In_233);
nand U52 (N_52,In_1824,In_704);
or U53 (N_53,In_1245,In_1214);
and U54 (N_54,In_1434,In_193);
nand U55 (N_55,In_1191,In_1341);
nand U56 (N_56,In_51,In_581);
nor U57 (N_57,In_1121,In_648);
or U58 (N_58,In_140,In_1364);
and U59 (N_59,In_167,In_236);
xor U60 (N_60,In_50,In_1426);
and U61 (N_61,In_1072,In_842);
xor U62 (N_62,In_1581,In_1660);
and U63 (N_63,In_1570,In_409);
xnor U64 (N_64,In_754,In_1068);
and U65 (N_65,In_1090,In_628);
nor U66 (N_66,In_731,In_687);
or U67 (N_67,In_1710,In_1933);
nand U68 (N_68,In_1777,In_575);
and U69 (N_69,In_829,In_703);
nor U70 (N_70,In_1427,In_1627);
or U71 (N_71,In_467,In_1975);
and U72 (N_72,In_989,In_525);
xor U73 (N_73,In_640,In_939);
xor U74 (N_74,In_945,In_1586);
xor U75 (N_75,In_1709,In_65);
and U76 (N_76,In_1651,In_1571);
nand U77 (N_77,In_1465,In_1456);
or U78 (N_78,In_1639,In_1860);
xnor U79 (N_79,In_66,In_215);
and U80 (N_80,In_1481,In_228);
nor U81 (N_81,In_306,In_895);
nand U82 (N_82,In_615,In_578);
nor U83 (N_83,In_1285,In_698);
and U84 (N_84,In_796,In_711);
nand U85 (N_85,In_153,In_21);
and U86 (N_86,In_1305,In_159);
nor U87 (N_87,In_484,In_906);
nand U88 (N_88,In_782,In_1882);
xnor U89 (N_89,In_191,In_1720);
xnor U90 (N_90,In_369,In_811);
nand U91 (N_91,In_1009,In_763);
xor U92 (N_92,In_492,In_693);
and U93 (N_93,In_1150,In_1007);
nand U94 (N_94,In_1474,In_1839);
xor U95 (N_95,In_559,In_868);
or U96 (N_96,In_1037,In_554);
xnor U97 (N_97,In_538,In_1874);
nor U98 (N_98,In_1061,In_410);
or U99 (N_99,In_296,In_299);
nor U100 (N_100,In_1036,In_1767);
and U101 (N_101,In_497,In_1739);
nand U102 (N_102,In_254,In_86);
nor U103 (N_103,In_977,In_102);
nor U104 (N_104,In_613,In_1751);
and U105 (N_105,In_113,In_637);
xor U106 (N_106,In_1263,In_1721);
xnor U107 (N_107,In_1868,In_882);
nor U108 (N_108,In_553,In_1417);
xnor U109 (N_109,In_1649,In_736);
or U110 (N_110,In_1587,In_1039);
xor U111 (N_111,In_442,In_803);
xor U112 (N_112,In_951,In_1485);
nor U113 (N_113,In_722,In_1325);
nand U114 (N_114,In_878,In_1560);
nand U115 (N_115,In_319,In_1504);
nor U116 (N_116,In_1237,In_1507);
nand U117 (N_117,In_433,In_728);
nand U118 (N_118,In_92,In_1692);
nor U119 (N_119,In_1284,In_1954);
and U120 (N_120,In_587,In_279);
nor U121 (N_121,In_1940,In_1979);
or U122 (N_122,In_762,In_1930);
nor U123 (N_123,In_590,In_1154);
xor U124 (N_124,In_1892,In_1566);
or U125 (N_125,In_1744,In_510);
nor U126 (N_126,In_269,In_747);
or U127 (N_127,In_1883,In_1439);
and U128 (N_128,In_922,In_18);
nor U129 (N_129,In_1287,In_1764);
xor U130 (N_130,In_1451,In_14);
or U131 (N_131,In_1588,In_935);
nand U132 (N_132,In_1190,In_1424);
xnor U133 (N_133,In_1182,In_1849);
and U134 (N_134,In_149,In_528);
xnor U135 (N_135,In_1642,In_1084);
nor U136 (N_136,In_1144,In_676);
nor U137 (N_137,In_99,In_1816);
and U138 (N_138,In_181,In_847);
and U139 (N_139,In_137,In_323);
nand U140 (N_140,In_1558,In_1733);
nand U141 (N_141,In_1471,In_28);
xor U142 (N_142,In_7,In_1663);
nor U143 (N_143,In_1708,In_1648);
nor U144 (N_144,In_596,In_1333);
and U145 (N_145,In_1138,In_1717);
or U146 (N_146,In_1185,In_1040);
and U147 (N_147,In_642,In_329);
or U148 (N_148,In_1384,In_1131);
or U149 (N_149,In_1549,In_1752);
or U150 (N_150,In_790,In_1477);
and U151 (N_151,In_923,In_143);
nor U152 (N_152,In_761,In_622);
and U153 (N_153,In_1048,In_1838);
nand U154 (N_154,In_1161,In_365);
xor U155 (N_155,In_958,In_74);
and U156 (N_156,In_320,In_1873);
nand U157 (N_157,In_476,In_1115);
xnor U158 (N_158,In_645,In_1126);
nor U159 (N_159,In_265,In_1593);
xor U160 (N_160,In_439,In_680);
xnor U161 (N_161,In_619,In_292);
xor U162 (N_162,In_534,In_871);
nor U163 (N_163,In_608,In_1445);
or U164 (N_164,In_1932,In_577);
or U165 (N_165,In_1572,In_422);
nor U166 (N_166,In_624,In_1791);
xor U167 (N_167,In_1595,In_83);
and U168 (N_168,In_1276,In_1974);
nand U169 (N_169,In_947,In_87);
nor U170 (N_170,In_562,In_1740);
and U171 (N_171,In_408,In_1047);
nand U172 (N_172,In_591,In_1666);
or U173 (N_173,In_1266,In_469);
and U174 (N_174,In_991,In_478);
nor U175 (N_175,In_1100,In_1086);
nor U176 (N_176,In_866,In_79);
nor U177 (N_177,In_1844,In_163);
and U178 (N_178,In_1802,In_1832);
xor U179 (N_179,In_1407,In_737);
and U180 (N_180,In_1329,In_1255);
or U181 (N_181,In_605,In_780);
nor U182 (N_182,In_1971,In_740);
nor U183 (N_183,In_1685,In_700);
nor U184 (N_184,In_1600,In_1447);
xor U185 (N_185,In_996,In_348);
nor U186 (N_186,In_558,In_828);
nor U187 (N_187,In_1205,In_527);
and U188 (N_188,In_1830,In_1807);
nor U189 (N_189,In_1810,In_15);
nor U190 (N_190,In_795,In_530);
nand U191 (N_191,In_1521,In_1309);
nand U192 (N_192,In_1992,In_1050);
or U193 (N_193,In_705,In_571);
xnor U194 (N_194,In_373,In_207);
xnor U195 (N_195,In_238,In_1184);
nor U196 (N_196,In_599,In_1177);
nor U197 (N_197,In_1041,In_1563);
nand U198 (N_198,In_1062,In_101);
nor U199 (N_199,In_1917,In_1962);
xor U200 (N_200,In_234,In_1112);
nand U201 (N_201,In_186,In_165);
or U202 (N_202,In_979,In_573);
or U203 (N_203,In_1057,In_1582);
nor U204 (N_204,In_1677,In_1348);
xor U205 (N_205,In_1897,In_589);
xor U206 (N_206,In_1332,In_1748);
and U207 (N_207,In_1562,In_1557);
and U208 (N_208,In_124,In_282);
and U209 (N_209,In_1955,In_1901);
nor U210 (N_210,In_1028,In_235);
and U211 (N_211,In_1053,In_1905);
xor U212 (N_212,In_1152,In_1706);
or U213 (N_213,In_849,In_1322);
or U214 (N_214,In_808,In_1271);
or U215 (N_215,In_658,In_1388);
xor U216 (N_216,In_976,In_97);
or U217 (N_217,In_148,In_1226);
xor U218 (N_218,In_1713,In_1995);
nand U219 (N_219,In_1404,In_824);
nor U220 (N_220,In_1159,In_1934);
xor U221 (N_221,In_1898,In_1984);
nor U222 (N_222,In_390,In_529);
nor U223 (N_223,In_157,In_49);
or U224 (N_224,In_1151,In_1551);
or U225 (N_225,In_760,In_1833);
nand U226 (N_226,In_860,In_1893);
and U227 (N_227,In_259,In_770);
and U228 (N_228,In_1645,In_170);
and U229 (N_229,In_1109,In_230);
or U230 (N_230,In_283,In_1188);
and U231 (N_231,In_1054,In_503);
nor U232 (N_232,In_1715,In_980);
or U233 (N_233,In_696,In_607);
nor U234 (N_234,In_1524,In_1358);
and U235 (N_235,In_863,In_482);
and U236 (N_236,In_1512,In_429);
nand U237 (N_237,In_1944,In_331);
and U238 (N_238,In_496,In_556);
nor U239 (N_239,In_1400,In_1380);
and U240 (N_240,In_726,In_924);
nor U241 (N_241,In_26,In_1272);
nand U242 (N_242,In_602,In_792);
or U243 (N_243,In_545,In_988);
and U244 (N_244,In_60,In_1568);
nor U245 (N_245,In_1443,In_1775);
and U246 (N_246,In_1218,In_603);
and U247 (N_247,In_861,In_121);
nand U248 (N_248,In_403,In_244);
or U249 (N_249,In_752,In_973);
or U250 (N_250,In_555,In_1886);
nand U251 (N_251,In_1500,In_75);
or U252 (N_252,In_84,In_1441);
and U253 (N_253,In_1489,In_1761);
nand U254 (N_254,In_1069,In_1700);
xor U255 (N_255,In_526,In_315);
or U256 (N_256,In_1470,In_750);
xor U257 (N_257,In_444,In_1852);
nand U258 (N_258,In_1246,In_1371);
nor U259 (N_259,In_69,In_1135);
or U260 (N_260,In_1731,In_185);
nor U261 (N_261,In_253,In_1820);
nor U262 (N_262,In_196,In_1476);
or U263 (N_263,In_1981,In_470);
and U264 (N_264,In_764,In_174);
and U265 (N_265,In_1727,In_798);
nand U266 (N_266,In_1909,In_1372);
xor U267 (N_267,In_1884,In_1804);
nand U268 (N_268,In_506,In_73);
and U269 (N_269,In_1450,In_543);
xnor U270 (N_270,In_383,In_473);
nand U271 (N_271,In_354,In_1075);
xnor U272 (N_272,In_29,In_1950);
or U273 (N_273,In_1612,In_1834);
xor U274 (N_274,In_1343,In_1051);
nor U275 (N_275,In_115,In_1356);
nor U276 (N_276,In_1398,In_147);
or U277 (N_277,In_956,In_1031);
or U278 (N_278,In_1005,In_1292);
xor U279 (N_279,In_1654,In_943);
nand U280 (N_280,In_1679,In_31);
nand U281 (N_281,In_1165,In_1610);
and U282 (N_282,In_400,In_967);
nand U283 (N_283,In_1758,In_1);
and U284 (N_284,In_633,In_109);
nand U285 (N_285,In_1196,In_430);
xor U286 (N_286,In_1669,In_928);
and U287 (N_287,In_453,In_1723);
nor U288 (N_288,In_1861,In_686);
or U289 (N_289,In_656,In_17);
xor U290 (N_290,In_356,In_1118);
or U291 (N_291,In_626,In_1703);
nor U292 (N_292,In_1147,In_158);
xor U293 (N_293,In_994,In_59);
nor U294 (N_294,In_366,In_1197);
and U295 (N_295,In_1446,In_667);
or U296 (N_296,In_990,In_1049);
or U297 (N_297,In_440,In_1798);
or U298 (N_298,In_195,In_511);
nand U299 (N_299,In_838,In_182);
nor U300 (N_300,In_96,In_1542);
nor U301 (N_301,In_130,In_823);
nand U302 (N_302,In_561,In_1224);
or U303 (N_303,In_310,In_614);
nor U304 (N_304,In_907,In_583);
nor U305 (N_305,In_229,In_198);
and U306 (N_306,In_890,In_1594);
nand U307 (N_307,In_710,In_948);
or U308 (N_308,In_1484,In_1926);
xnor U309 (N_309,In_567,In_1863);
or U310 (N_310,In_565,In_1302);
xor U311 (N_311,In_39,In_291);
or U312 (N_312,In_1296,In_474);
or U313 (N_313,In_783,In_1393);
or U314 (N_314,In_1657,In_415);
xnor U315 (N_315,In_1584,In_1503);
nor U316 (N_316,In_166,In_123);
nor U317 (N_317,In_1004,In_20);
or U318 (N_318,In_1490,In_1724);
xor U319 (N_319,In_1643,In_1737);
nor U320 (N_320,In_216,In_1518);
xnor U321 (N_321,In_1479,In_885);
nand U322 (N_322,In_1534,In_104);
and U323 (N_323,In_1961,In_112);
xor U324 (N_324,In_779,In_1070);
or U325 (N_325,In_1986,In_222);
or U326 (N_326,In_1106,In_1415);
xor U327 (N_327,In_1107,In_1281);
nand U328 (N_328,In_171,In_1460);
or U329 (N_329,In_508,In_649);
xnor U330 (N_330,In_1577,In_1795);
and U331 (N_331,In_1728,In_1083);
or U332 (N_332,In_1334,In_1851);
xnor U333 (N_333,In_954,In_892);
nand U334 (N_334,In_955,In_490);
nand U335 (N_335,In_392,In_1122);
and U336 (N_336,In_1312,In_1038);
nor U337 (N_337,In_1776,In_1349);
and U338 (N_338,In_1972,In_1841);
and U339 (N_339,In_1499,In_1468);
nor U340 (N_340,In_643,In_1908);
nand U341 (N_341,In_952,In_220);
and U342 (N_342,In_616,In_862);
nor U343 (N_343,In_1513,In_1300);
or U344 (N_344,In_379,In_1402);
or U345 (N_345,In_368,In_769);
nor U346 (N_346,In_271,In_897);
and U347 (N_347,In_1401,In_1444);
nor U348 (N_348,In_1442,In_515);
nand U349 (N_349,In_593,In_475);
nand U350 (N_350,In_91,In_802);
xnor U351 (N_351,In_1410,In_1265);
nor U352 (N_352,In_682,In_815);
nor U353 (N_353,In_1353,In_1192);
nand U354 (N_354,In_217,In_814);
or U355 (N_355,In_1960,In_625);
or U356 (N_356,In_1429,In_1228);
nand U357 (N_357,In_777,In_33);
or U358 (N_358,In_566,In_1307);
and U359 (N_359,In_1578,In_1517);
xor U360 (N_360,In_1003,In_1136);
nand U361 (N_361,In_720,In_513);
or U362 (N_362,In_1668,In_839);
nand U363 (N_363,In_1078,In_1769);
nor U364 (N_364,In_1127,In_1902);
and U365 (N_365,In_959,In_1298);
nor U366 (N_366,In_1203,In_1613);
and U367 (N_367,In_930,In_1806);
nor U368 (N_368,In_1071,In_1799);
nor U369 (N_369,In_162,In_324);
nand U370 (N_370,In_1472,In_1698);
and U371 (N_371,In_301,In_774);
nand U372 (N_372,In_1094,In_723);
nor U373 (N_373,In_1956,In_1826);
nor U374 (N_374,In_1686,In_332);
nand U375 (N_375,In_1350,In_404);
nand U376 (N_376,In_1313,In_141);
nor U377 (N_377,In_1406,In_1162);
or U378 (N_378,In_267,In_1983);
nand U379 (N_379,In_509,In_1869);
nand U380 (N_380,In_1336,In_1605);
or U381 (N_381,In_1483,In_1779);
and U382 (N_382,In_1045,In_6);
nor U383 (N_383,In_10,In_1297);
or U384 (N_384,In_1019,In_1314);
xnor U385 (N_385,In_540,In_328);
nand U386 (N_386,In_970,In_1516);
nand U387 (N_387,In_70,In_1428);
nand U388 (N_388,In_445,In_455);
nand U389 (N_389,In_968,In_1601);
nor U390 (N_390,In_1008,In_1033);
xnor U391 (N_391,In_679,In_1615);
nand U392 (N_392,In_201,In_789);
nand U393 (N_393,In_118,In_1209);
xnor U394 (N_394,In_342,In_303);
nand U395 (N_395,In_1792,In_1701);
nand U396 (N_396,In_1347,In_477);
nand U397 (N_397,In_683,In_1875);
or U398 (N_398,In_1023,In_576);
nand U399 (N_399,In_172,In_1545);
nand U400 (N_400,In_813,In_1058);
or U401 (N_401,In_192,In_1414);
or U402 (N_402,In_168,In_135);
or U403 (N_403,In_1585,In_133);
xor U404 (N_404,In_1469,In_1103);
nand U405 (N_405,In_899,In_689);
nor U406 (N_406,In_749,In_499);
or U407 (N_407,In_1000,In_821);
xnor U408 (N_408,In_1634,In_1219);
xnor U409 (N_409,In_612,In_1101);
nand U410 (N_410,In_800,In_845);
xor U411 (N_411,In_1644,In_756);
and U412 (N_412,In_1815,In_1609);
xor U413 (N_413,In_1772,In_716);
or U414 (N_414,In_1020,In_1495);
nand U415 (N_415,In_1969,In_169);
and U416 (N_416,In_953,In_184);
and U417 (N_417,In_1042,In_1553);
or U418 (N_418,In_1620,In_1064);
or U419 (N_419,In_1319,In_1174);
nand U420 (N_420,In_114,In_1531);
nor U421 (N_421,In_804,In_684);
and U422 (N_422,In_1964,In_569);
nand U423 (N_423,In_500,In_1360);
xnor U424 (N_424,In_1320,In_155);
or U425 (N_425,In_67,In_1965);
and U426 (N_426,In_1729,In_1169);
or U427 (N_427,In_1425,In_1963);
and U428 (N_428,In_1695,In_1662);
and U429 (N_429,In_1317,In_1110);
or U430 (N_430,In_1920,In_1528);
or U431 (N_431,In_582,In_491);
nor U432 (N_432,In_631,In_435);
xor U433 (N_433,In_739,In_721);
and U434 (N_434,In_786,In_1506);
or U435 (N_435,In_350,In_827);
and U436 (N_436,In_1105,In_1195);
nor U437 (N_437,In_1164,In_258);
nand U438 (N_438,In_1034,In_212);
or U439 (N_439,In_743,In_714);
and U440 (N_440,In_911,In_1330);
and U441 (N_441,In_1511,In_1149);
and U442 (N_442,In_1432,In_1491);
nor U443 (N_443,In_888,In_1665);
and U444 (N_444,In_335,In_936);
and U445 (N_445,In_434,In_1200);
nor U446 (N_446,In_1555,In_1722);
or U447 (N_447,In_1959,In_966);
and U448 (N_448,In_1535,In_1683);
xor U449 (N_449,In_106,In_652);
xor U450 (N_450,In_934,In_1013);
nand U451 (N_451,In_1821,In_294);
xor U452 (N_452,In_1732,In_116);
nand U453 (N_453,In_384,In_1148);
and U454 (N_454,In_801,In_77);
xor U455 (N_455,In_1976,In_1712);
nand U456 (N_456,In_982,In_176);
nand U457 (N_457,In_1381,In_1694);
and U458 (N_458,In_1552,In_1327);
and U459 (N_459,In_1240,In_441);
and U460 (N_460,In_601,In_1340);
xor U461 (N_461,In_903,In_1793);
or U462 (N_462,In_1173,In_1597);
or U463 (N_463,In_183,In_1900);
or U464 (N_464,In_43,In_702);
and U465 (N_465,In_856,In_518);
and U466 (N_466,In_787,In_531);
nor U467 (N_467,In_1696,In_1487);
or U468 (N_468,In_347,In_250);
xor U469 (N_469,In_832,In_1918);
nor U470 (N_470,In_1213,In_333);
xnor U471 (N_471,In_910,In_879);
nor U472 (N_472,In_1906,In_443);
nand U473 (N_473,In_918,In_80);
nand U474 (N_474,In_549,In_1966);
nand U475 (N_475,In_398,In_1208);
or U476 (N_476,In_1947,In_210);
nand U477 (N_477,In_358,In_32);
or U478 (N_478,In_64,In_108);
or U479 (N_479,In_399,In_993);
or U480 (N_480,In_1508,In_1590);
and U481 (N_481,In_418,In_664);
nand U482 (N_482,In_893,In_1622);
nand U483 (N_483,In_8,In_1843);
nor U484 (N_484,In_1635,In_1750);
nor U485 (N_485,In_391,In_1006);
or U486 (N_486,In_338,In_431);
and U487 (N_487,In_846,In_604);
nor U488 (N_488,In_1699,In_1248);
xor U489 (N_489,In_1606,In_858);
or U490 (N_490,In_805,In_437);
nor U491 (N_491,In_452,In_1746);
nand U492 (N_492,In_1670,In_1523);
xor U493 (N_493,In_1129,In_411);
or U494 (N_494,In_732,In_665);
and U495 (N_495,In_1390,In_785);
nand U496 (N_496,In_1194,In_364);
nand U497 (N_497,In_1095,In_464);
and U498 (N_498,In_1957,In_797);
nor U499 (N_499,In_997,In_1848);
nor U500 (N_500,In_1080,In_1636);
and U501 (N_501,In_48,In_9);
nand U502 (N_502,In_1186,In_929);
nor U503 (N_503,In_675,In_992);
or U504 (N_504,In_659,In_1502);
xnor U505 (N_505,In_1257,In_532);
or U506 (N_506,In_1099,In_1486);
and U507 (N_507,In_1970,In_1537);
nand U508 (N_508,In_1990,In_1289);
nand U509 (N_509,In_1201,In_1012);
and U510 (N_510,In_1338,In_630);
or U511 (N_511,In_1817,In_1653);
xnor U512 (N_512,In_231,In_1056);
nand U513 (N_513,In_1206,In_1621);
nand U514 (N_514,In_393,In_1459);
nand U515 (N_515,In_902,In_396);
xor U516 (N_516,In_1242,In_751);
and U517 (N_517,In_1383,In_1423);
or U518 (N_518,In_278,In_56);
xor U519 (N_519,In_1128,In_1805);
and U520 (N_520,In_533,In_131);
nor U521 (N_521,In_1158,In_1525);
xnor U522 (N_522,In_784,In_1464);
xor U523 (N_523,In_1141,In_1420);
and U524 (N_524,In_1367,In_502);
and U525 (N_525,In_1324,In_465);
nor U526 (N_526,In_1994,In_1980);
xor U527 (N_527,In_1286,In_1658);
nor U528 (N_528,In_867,In_1556);
or U529 (N_529,In_454,In_937);
or U530 (N_530,In_519,In_188);
or U531 (N_531,In_251,In_1714);
and U532 (N_532,In_1923,In_1738);
and U533 (N_533,In_1014,In_621);
nand U534 (N_534,In_405,In_639);
or U535 (N_535,In_620,In_1193);
nand U536 (N_536,In_913,In_1633);
xnor U537 (N_537,In_1303,In_1304);
xor U538 (N_538,In_428,In_1467);
and U539 (N_539,In_1046,In_1766);
and U540 (N_540,In_394,In_1029);
and U541 (N_541,In_809,In_1611);
xor U542 (N_542,In_807,In_276);
nor U543 (N_543,In_793,In_835);
nand U544 (N_544,In_757,In_1362);
or U545 (N_545,In_771,In_205);
nand U546 (N_546,In_485,In_1244);
nor U547 (N_547,In_1187,In_1475);
xnor U548 (N_548,In_1408,In_1280);
xnor U549 (N_549,In_1641,In_1896);
xnor U550 (N_550,In_964,In_16);
xor U551 (N_551,In_1290,In_1889);
or U552 (N_552,In_908,In_501);
and U553 (N_553,In_419,In_1262);
nor U554 (N_554,In_1656,In_915);
xor U555 (N_555,In_592,In_1842);
nand U556 (N_556,In_1098,In_458);
nor U557 (N_557,In_1711,In_685);
nor U558 (N_558,In_1825,In_280);
xnor U559 (N_559,In_427,In_1386);
nor U560 (N_560,In_830,In_810);
nand U561 (N_561,In_1941,In_1409);
nand U562 (N_562,In_678,In_1283);
nor U563 (N_563,In_1172,In_1774);
xnor U564 (N_564,In_834,In_218);
or U565 (N_565,In_734,In_180);
or U566 (N_566,In_1171,In_1331);
xnor U567 (N_567,In_1124,In_107);
nor U568 (N_568,In_1096,In_961);
or U569 (N_569,In_742,In_456);
nand U570 (N_570,In_361,In_1249);
or U571 (N_571,In_42,In_1973);
nand U572 (N_572,In_853,In_1747);
nor U573 (N_573,In_901,In_483);
and U574 (N_574,In_55,In_983);
or U575 (N_575,In_874,In_588);
or U576 (N_576,In_1759,In_1243);
nand U577 (N_577,In_95,In_1803);
xnor U578 (N_578,In_190,In_1421);
nor U579 (N_579,In_1321,In_288);
xnor U580 (N_580,In_242,In_1076);
or U581 (N_581,In_11,In_1554);
nor U582 (N_582,In_1215,In_1310);
or U583 (N_583,In_145,In_875);
xor U584 (N_584,In_551,In_1631);
and U585 (N_585,In_1559,In_1749);
nor U586 (N_586,In_1828,In_1888);
nor U587 (N_587,In_1702,In_1431);
or U588 (N_588,In_641,In_1181);
or U589 (N_589,In_644,In_5);
nor U590 (N_590,In_851,In_1134);
or U591 (N_591,In_1596,In_1435);
nor U592 (N_592,In_1942,In_128);
nor U593 (N_593,In_1707,In_1232);
or U594 (N_594,In_1130,In_877);
nor U595 (N_595,In_1236,In_256);
xnor U596 (N_596,In_1032,In_1894);
and U597 (N_597,In_88,In_663);
or U598 (N_598,In_1220,In_295);
xnor U599 (N_599,In_636,In_606);
xor U600 (N_600,In_1230,In_1306);
xor U601 (N_601,In_1629,In_111);
nor U602 (N_602,In_1392,In_1617);
nor U603 (N_603,In_1801,In_326);
xor U604 (N_604,In_493,In_960);
and U605 (N_605,In_799,In_896);
nand U606 (N_606,In_850,In_1077);
nor U607 (N_607,In_505,In_262);
nor U608 (N_608,In_841,In_1375);
xnor U609 (N_609,In_1233,In_611);
or U610 (N_610,In_46,In_206);
or U611 (N_611,In_1880,In_1790);
and U612 (N_612,In_246,In_962);
nand U613 (N_613,In_708,In_1123);
nor U614 (N_614,In_187,In_54);
and U615 (N_615,In_1235,In_1675);
nand U616 (N_616,In_240,In_887);
nor U617 (N_617,In_426,In_243);
xnor U618 (N_618,In_327,In_1411);
nand U619 (N_619,In_632,In_1952);
nand U620 (N_620,In_1291,In_1279);
or U621 (N_621,In_1395,In_1261);
xor U622 (N_622,In_1339,In_225);
xor U623 (N_623,In_311,In_1985);
and U624 (N_624,In_1389,In_468);
nor U625 (N_625,In_200,In_1010);
or U626 (N_626,In_1575,In_1533);
or U627 (N_627,In_766,In_1678);
nor U628 (N_628,In_1796,In_820);
nor U629 (N_629,In_312,In_1452);
or U630 (N_630,In_260,In_1837);
xnor U631 (N_631,In_1368,In_1659);
nand U632 (N_632,In_1867,In_446);
and U633 (N_633,In_1278,In_448);
nand U634 (N_634,In_677,In_768);
nand U635 (N_635,In_1035,In_1982);
nor U636 (N_636,In_1866,In_395);
or U637 (N_637,In_1337,In_655);
and U638 (N_638,In_461,In_681);
nor U639 (N_639,In_1768,In_305);
or U640 (N_640,In_376,In_1797);
nor U641 (N_641,In_24,In_1529);
and U642 (N_642,In_1342,In_919);
nand U643 (N_643,In_209,In_1931);
xnor U644 (N_644,In_522,In_1693);
and U645 (N_645,In_600,In_1377);
and U646 (N_646,In_699,In_4);
nor U647 (N_647,In_266,In_1418);
nor U648 (N_648,In_1180,In_791);
nor U649 (N_649,In_1786,In_816);
xor U650 (N_650,In_938,In_488);
and U651 (N_651,In_1911,In_759);
nand U652 (N_652,In_707,In_367);
or U653 (N_653,In_1773,In_1308);
nand U654 (N_654,In_564,In_334);
nand U655 (N_655,In_822,In_353);
nand U656 (N_656,In_512,In_1346);
nor U657 (N_657,In_634,In_1092);
nand U658 (N_658,In_869,In_1505);
xor U659 (N_659,In_208,In_330);
and U660 (N_660,In_572,In_1741);
xnor U661 (N_661,In_773,In_753);
or U662 (N_662,In_1872,In_37);
xnor U663 (N_663,In_25,In_214);
xor U664 (N_664,In_1216,In_1183);
nand U665 (N_665,In_1879,In_1770);
or U666 (N_666,In_1604,In_58);
nand U667 (N_667,In_1116,In_173);
nor U668 (N_668,In_308,In_660);
nand U669 (N_669,In_1156,In_688);
nor U670 (N_670,In_1780,In_178);
or U671 (N_671,In_1602,In_1864);
nor U672 (N_672,In_1808,In_1988);
nand U673 (N_673,In_1063,In_1207);
and U674 (N_674,In_1082,In_142);
and U675 (N_675,In_1223,In_916);
and U676 (N_676,In_1550,In_1087);
nor U677 (N_677,In_1592,In_436);
xnor U678 (N_678,In_160,In_523);
or U679 (N_679,In_1253,In_406);
and U680 (N_680,In_1433,In_950);
or U681 (N_681,In_268,In_695);
nand U682 (N_682,In_1788,In_972);
xnor U683 (N_683,In_963,In_719);
nand U684 (N_684,In_1599,In_1146);
xor U685 (N_685,In_1277,In_1403);
or U686 (N_686,In_1394,In_694);
and U687 (N_687,In_981,In_1416);
or U688 (N_688,In_1113,In_1845);
nand U689 (N_689,In_247,In_568);
nand U690 (N_690,In_609,In_748);
xor U691 (N_691,In_413,In_146);
nand U692 (N_692,In_1929,In_281);
nor U693 (N_693,In_1176,In_889);
nor U694 (N_694,In_203,In_136);
nand U695 (N_695,In_1163,In_715);
nand U696 (N_696,In_1379,In_1945);
nand U697 (N_697,In_1114,In_219);
xnor U698 (N_698,In_1132,In_623);
or U699 (N_699,In_352,In_1924);
or U700 (N_700,In_417,In_548);
nor U701 (N_701,In_1254,In_1093);
and U702 (N_702,In_122,In_884);
xnor U703 (N_703,In_547,In_100);
xor U704 (N_704,In_127,In_579);
nor U705 (N_705,In_1373,In_1536);
xnor U706 (N_706,In_669,In_386);
or U707 (N_707,In_1921,In_98);
xor U708 (N_708,In_635,In_1457);
and U709 (N_709,In_1251,In_1419);
xor U710 (N_710,In_586,In_1822);
nand U711 (N_711,In_1638,In_1519);
nor U712 (N_712,In_1652,In_978);
and U713 (N_713,In_1412,In_1655);
nand U714 (N_714,In_345,In_661);
nor U715 (N_715,In_629,In_472);
nand U716 (N_716,In_876,In_82);
nor U717 (N_717,In_110,In_1282);
xor U718 (N_718,In_1376,In_1104);
and U719 (N_719,In_504,In_1260);
or U720 (N_720,In_460,In_375);
or U721 (N_721,In_1546,In_1097);
and U722 (N_722,In_286,In_1315);
xor U723 (N_723,In_103,In_1569);
nand U724 (N_724,In_1024,In_22);
nand U725 (N_725,In_264,In_1765);
xnor U726 (N_726,In_563,In_126);
nand U727 (N_727,In_189,In_1967);
xnor U728 (N_728,In_1354,In_1374);
nand U729 (N_729,In_1690,In_1664);
nand U730 (N_730,In_302,In_125);
nor U731 (N_731,In_672,In_293);
nor U732 (N_732,In_872,In_718);
or U733 (N_733,In_1937,In_585);
and U734 (N_734,In_1989,In_1540);
nand U735 (N_735,In_1073,In_541);
or U736 (N_736,In_339,In_1730);
nand U737 (N_737,In_1762,In_1264);
nand U738 (N_738,In_346,In_535);
nor U739 (N_739,In_1927,In_199);
or U740 (N_740,In_985,In_1405);
xnor U741 (N_741,In_852,In_537);
nor U742 (N_742,In_1968,In_341);
nand U743 (N_743,In_1997,In_1238);
nor U744 (N_744,In_273,In_357);
or U745 (N_745,In_755,In_975);
xor U746 (N_746,In_668,In_552);
xor U747 (N_747,In_725,In_974);
nand U748 (N_748,In_304,In_68);
or U749 (N_749,In_480,In_1922);
nand U750 (N_750,In_1274,In_156);
or U751 (N_751,In_1928,In_1060);
or U752 (N_752,In_481,In_1591);
nand U753 (N_753,In_300,In_421);
xor U754 (N_754,In_1632,In_942);
xnor U755 (N_755,In_1344,In_758);
or U756 (N_756,In_1267,In_1225);
or U757 (N_757,In_1522,In_941);
nand U758 (N_758,In_1782,In_580);
or U759 (N_759,In_1951,In_1091);
nor U760 (N_760,In_1227,In_1139);
nand U761 (N_761,In_520,In_2);
xor U762 (N_762,In_969,In_1085);
or U763 (N_763,In_1539,In_646);
or U764 (N_764,In_1170,In_1854);
or U765 (N_765,In_1914,In_1168);
and U766 (N_766,In_1526,In_387);
and U767 (N_767,In_27,In_1026);
nand U768 (N_768,In_1771,In_1199);
xnor U769 (N_769,In_420,In_1157);
xor U770 (N_770,In_733,In_1021);
nor U771 (N_771,In_1899,In_775);
nand U772 (N_772,In_776,In_1067);
or U773 (N_773,In_1378,In_1482);
or U774 (N_774,In_397,In_881);
xnor U775 (N_775,In_883,In_1887);
nor U776 (N_776,In_709,In_340);
xnor U777 (N_777,In_1811,In_594);
and U778 (N_778,In_1573,In_129);
nor U779 (N_779,In_638,In_462);
and U780 (N_780,In_1498,In_1202);
nor U781 (N_781,In_94,In_274);
nand U782 (N_782,In_778,In_1705);
nor U783 (N_783,In_1370,In_925);
nor U784 (N_784,In_653,In_463);
nand U785 (N_785,In_1515,In_1736);
nor U786 (N_786,In_495,In_971);
and U787 (N_787,In_284,In_498);
or U788 (N_788,In_1831,In_351);
nor U789 (N_789,In_957,In_1530);
nor U790 (N_790,In_880,In_1102);
nand U791 (N_791,In_1231,In_314);
xor U792 (N_792,In_298,In_53);
nand U793 (N_793,In_1603,In_19);
xnor U794 (N_794,In_1361,In_898);
nand U795 (N_795,In_237,In_940);
or U796 (N_796,In_1681,In_741);
nand U797 (N_797,In_542,In_287);
nand U798 (N_798,In_1544,In_794);
or U799 (N_799,In_744,In_1625);
nor U800 (N_800,In_1256,In_912);
or U801 (N_801,In_263,In_697);
nor U802 (N_802,In_1081,In_1859);
or U803 (N_803,In_1809,In_1853);
and U804 (N_804,In_1904,In_921);
and U805 (N_805,In_1241,In_539);
and U806 (N_806,In_211,In_1907);
xor U807 (N_807,In_1671,In_1189);
or U808 (N_808,In_864,In_999);
nor U809 (N_809,In_1366,In_627);
or U810 (N_810,In_257,In_1865);
or U811 (N_811,In_1458,In_550);
xnor U812 (N_812,In_1509,In_1835);
or U813 (N_813,In_1142,In_344);
and U814 (N_814,In_213,In_514);
or U815 (N_815,In_1119,In_1734);
xor U816 (N_816,In_570,In_1948);
nor U817 (N_817,In_1543,In_34);
xnor U818 (N_818,In_459,In_1680);
xnor U819 (N_819,In_859,In_309);
nor U820 (N_820,In_873,In_1318);
nand U821 (N_821,In_1125,In_1876);
nand U822 (N_822,In_81,In_61);
nand U823 (N_823,In_1640,In_447);
nor U824 (N_824,In_1754,In_1673);
nor U825 (N_825,In_1813,In_245);
nand U826 (N_826,In_41,In_1268);
and U827 (N_827,In_965,In_402);
xnor U828 (N_828,In_837,In_202);
or U829 (N_829,In_389,In_1725);
xor U830 (N_830,In_1437,In_255);
xor U831 (N_831,In_1357,In_1871);
xnor U832 (N_832,In_854,In_618);
nor U833 (N_833,In_322,In_855);
nor U834 (N_834,In_1756,In_574);
nor U835 (N_835,In_151,In_1143);
and U836 (N_836,In_1155,In_1001);
and U837 (N_837,In_175,In_1204);
nand U838 (N_838,In_1438,In_355);
xnor U839 (N_839,In_0,In_1211);
or U840 (N_840,In_647,In_72);
nand U841 (N_841,In_1065,In_150);
nor U842 (N_842,In_371,In_836);
and U843 (N_843,In_239,In_598);
or U844 (N_844,In_1133,In_584);
nand U845 (N_845,In_1857,In_944);
and U846 (N_846,In_1345,In_71);
or U847 (N_847,In_90,In_489);
or U848 (N_848,In_1221,In_1814);
or U849 (N_849,In_1547,In_449);
xor U850 (N_850,In_1454,In_507);
nand U851 (N_851,In_1492,In_1647);
nor U852 (N_852,In_1862,In_1946);
nor U853 (N_853,In_325,In_1448);
or U854 (N_854,In_1466,In_772);
nand U855 (N_855,In_1269,In_1449);
nor U856 (N_856,In_674,In_844);
xnor U857 (N_857,In_438,In_706);
xor U858 (N_858,In_1667,In_1140);
xor U859 (N_859,In_224,In_1488);
and U860 (N_860,In_1166,In_1385);
or U861 (N_861,In_765,In_1212);
and U862 (N_862,In_1561,In_412);
and U863 (N_863,In_154,In_457);
or U864 (N_864,In_1328,In_1623);
and U865 (N_865,In_63,In_1794);
nand U866 (N_866,In_521,In_1850);
or U867 (N_867,In_1745,In_1217);
or U868 (N_868,In_1778,In_729);
and U869 (N_869,In_1674,In_1925);
xnor U870 (N_870,In_946,In_1074);
and U871 (N_871,In_1949,In_1565);
nor U872 (N_872,In_1935,In_1299);
nand U873 (N_873,In_407,In_401);
nand U874 (N_874,In_1614,In_47);
and U875 (N_875,In_1576,In_1497);
and U876 (N_876,In_317,In_657);
xnor U877 (N_877,In_833,In_524);
nand U878 (N_878,In_857,In_134);
or U879 (N_879,In_516,In_471);
xnor U880 (N_880,In_1137,In_378);
nor U881 (N_881,In_380,In_1079);
or U882 (N_882,In_336,In_318);
and U883 (N_883,In_451,In_1781);
nand U884 (N_884,In_1496,In_1616);
nand U885 (N_885,In_289,In_1958);
xnor U886 (N_886,In_1089,In_1608);
nor U887 (N_887,In_597,In_717);
and U888 (N_888,In_1719,In_1676);
and U889 (N_889,In_35,In_1301);
nor U890 (N_890,In_1829,In_1055);
nand U891 (N_891,In_241,In_1258);
or U892 (N_892,In_1016,In_712);
xor U893 (N_893,In_1913,In_363);
nor U894 (N_894,In_360,In_132);
xnor U895 (N_895,In_3,In_23);
xnor U896 (N_896,In_1953,In_1718);
nor U897 (N_897,In_1532,In_1661);
or U898 (N_898,In_1234,In_1755);
nor U899 (N_899,In_1823,In_1088);
nand U900 (N_900,In_1351,In_52);
nand U901 (N_901,In_920,In_1891);
nor U902 (N_902,In_650,In_1987);
or U903 (N_903,In_927,In_494);
nand U904 (N_904,In_249,In_1996);
or U905 (N_905,In_1630,In_1998);
or U906 (N_906,In_1991,In_1473);
xnor U907 (N_907,In_1252,In_423);
and U908 (N_908,In_691,In_1735);
nor U909 (N_909,In_1912,In_1397);
or U910 (N_910,In_362,In_986);
xnor U911 (N_911,In_995,In_1618);
or U912 (N_912,In_85,In_713);
nor U913 (N_913,In_374,In_1783);
or U914 (N_914,In_78,In_1650);
nor U915 (N_915,In_1520,In_1567);
and U916 (N_916,In_730,In_93);
nor U917 (N_917,In_1938,In_1939);
nor U918 (N_918,In_1117,In_277);
xnor U919 (N_919,In_826,In_1910);
and U920 (N_920,In_12,In_1895);
nor U921 (N_921,In_932,In_285);
or U922 (N_922,In_1598,In_1355);
nand U923 (N_923,In_1382,In_1059);
and U924 (N_924,In_76,In_316);
or U925 (N_925,In_1836,In_248);
nor U926 (N_926,In_1977,In_487);
nor U927 (N_927,In_1387,In_1043);
xnor U928 (N_928,In_984,In_221);
nand U929 (N_929,In_424,In_840);
xnor U930 (N_930,In_382,In_1422);
or U931 (N_931,In_1461,In_1687);
nand U932 (N_932,In_1025,In_1784);
and U933 (N_933,In_1259,In_1396);
and U934 (N_934,In_1145,In_1688);
and U935 (N_935,In_1222,In_1018);
nand U936 (N_936,In_1993,In_343);
or U937 (N_937,In_38,In_36);
xnor U938 (N_938,In_1890,In_1179);
nand U939 (N_939,In_1763,In_1326);
nand U940 (N_940,In_1716,In_738);
xnor U941 (N_941,In_179,In_1022);
nand U942 (N_942,In_479,In_194);
nor U943 (N_943,In_767,In_517);
xor U944 (N_944,In_388,In_1153);
nor U945 (N_945,In_1198,In_164);
xnor U946 (N_946,In_1167,In_1818);
or U947 (N_947,In_1335,In_1541);
or U948 (N_948,In_914,In_1015);
and U949 (N_949,In_806,In_1626);
and U950 (N_950,In_1789,In_546);
nor U951 (N_951,In_1999,In_949);
xnor U952 (N_952,In_1704,In_321);
and U953 (N_953,In_727,In_1108);
nor U954 (N_954,In_89,In_349);
nand U955 (N_955,In_1877,In_370);
or U956 (N_956,In_1684,In_557);
or U957 (N_957,In_307,In_870);
nand U958 (N_958,In_1697,In_1275);
nor U959 (N_959,In_1175,In_1178);
nand U960 (N_960,In_197,In_931);
nor U961 (N_961,In_595,In_1494);
nor U962 (N_962,In_270,In_1316);
or U963 (N_963,In_1689,In_900);
nor U964 (N_964,In_1480,In_905);
and U965 (N_965,In_1624,In_617);
nor U966 (N_966,In_1672,In_1574);
nor U967 (N_967,In_891,In_1607);
or U968 (N_968,In_1363,In_138);
nor U969 (N_969,In_1311,In_261);
and U970 (N_970,In_290,In_788);
or U971 (N_971,In_1579,In_1352);
nand U972 (N_972,In_812,In_144);
and U973 (N_973,In_1391,In_381);
nor U974 (N_974,In_1294,In_1453);
and U975 (N_975,In_1413,In_1548);
xnor U976 (N_976,In_272,In_1760);
nor U977 (N_977,In_1682,In_1757);
nor U978 (N_978,In_232,In_105);
nand U979 (N_979,In_1011,In_673);
xnor U980 (N_980,In_654,In_1247);
nand U981 (N_981,In_987,In_1066);
nand U982 (N_982,In_666,In_1742);
xnor U983 (N_983,In_177,In_651);
nand U984 (N_984,In_1455,In_297);
xor U985 (N_985,In_544,In_1847);
nor U986 (N_986,In_359,In_848);
or U987 (N_987,In_275,In_735);
and U988 (N_988,In_818,In_865);
nor U989 (N_989,In_1514,In_1726);
xor U990 (N_990,In_671,In_1463);
and U991 (N_991,In_414,In_1239);
nor U992 (N_992,In_1580,In_1819);
nand U993 (N_993,In_1510,In_886);
nand U994 (N_994,In_1564,In_1160);
xnor U995 (N_995,In_1493,In_1943);
and U996 (N_996,In_1369,In_1293);
or U997 (N_997,In_1628,In_1210);
xor U998 (N_998,In_40,In_385);
or U999 (N_999,In_662,In_1583);
nand U1000 (N_1000,In_1302,In_1012);
nor U1001 (N_1001,In_610,In_396);
or U1002 (N_1002,In_1904,In_662);
nor U1003 (N_1003,In_404,In_7);
nor U1004 (N_1004,In_1999,In_1897);
or U1005 (N_1005,In_1532,In_1695);
xnor U1006 (N_1006,In_1072,In_137);
nand U1007 (N_1007,In_442,In_1858);
and U1008 (N_1008,In_382,In_629);
and U1009 (N_1009,In_1620,In_988);
xnor U1010 (N_1010,In_1267,In_1246);
nor U1011 (N_1011,In_470,In_932);
and U1012 (N_1012,In_1864,In_495);
and U1013 (N_1013,In_529,In_736);
nand U1014 (N_1014,In_1297,In_355);
or U1015 (N_1015,In_1054,In_246);
nand U1016 (N_1016,In_1684,In_781);
or U1017 (N_1017,In_1811,In_142);
or U1018 (N_1018,In_1384,In_1751);
or U1019 (N_1019,In_1603,In_1398);
nand U1020 (N_1020,In_1925,In_712);
and U1021 (N_1021,In_171,In_87);
nor U1022 (N_1022,In_1785,In_1558);
and U1023 (N_1023,In_589,In_663);
and U1024 (N_1024,In_665,In_1430);
and U1025 (N_1025,In_1251,In_262);
and U1026 (N_1026,In_715,In_956);
nand U1027 (N_1027,In_994,In_1265);
nor U1028 (N_1028,In_361,In_1559);
nor U1029 (N_1029,In_636,In_1179);
nand U1030 (N_1030,In_755,In_1100);
and U1031 (N_1031,In_768,In_738);
or U1032 (N_1032,In_1090,In_771);
nor U1033 (N_1033,In_1323,In_438);
and U1034 (N_1034,In_1681,In_1820);
and U1035 (N_1035,In_1466,In_1436);
nand U1036 (N_1036,In_1165,In_1745);
and U1037 (N_1037,In_366,In_1905);
xor U1038 (N_1038,In_604,In_177);
nor U1039 (N_1039,In_844,In_186);
or U1040 (N_1040,In_1663,In_1460);
nor U1041 (N_1041,In_134,In_1570);
xnor U1042 (N_1042,In_1091,In_1394);
xor U1043 (N_1043,In_1929,In_1088);
nand U1044 (N_1044,In_789,In_1055);
xnor U1045 (N_1045,In_1986,In_1715);
nand U1046 (N_1046,In_1459,In_345);
nand U1047 (N_1047,In_264,In_221);
xnor U1048 (N_1048,In_1210,In_1437);
or U1049 (N_1049,In_633,In_530);
xnor U1050 (N_1050,In_1530,In_1521);
and U1051 (N_1051,In_1436,In_1989);
and U1052 (N_1052,In_14,In_234);
nand U1053 (N_1053,In_662,In_1864);
or U1054 (N_1054,In_699,In_967);
nor U1055 (N_1055,In_694,In_763);
nand U1056 (N_1056,In_1975,In_1041);
or U1057 (N_1057,In_612,In_1919);
xnor U1058 (N_1058,In_1864,In_576);
nor U1059 (N_1059,In_1525,In_632);
nor U1060 (N_1060,In_1145,In_598);
xnor U1061 (N_1061,In_173,In_190);
nor U1062 (N_1062,In_1314,In_403);
and U1063 (N_1063,In_1073,In_534);
and U1064 (N_1064,In_1348,In_224);
and U1065 (N_1065,In_1967,In_791);
nand U1066 (N_1066,In_692,In_190);
nand U1067 (N_1067,In_782,In_548);
nand U1068 (N_1068,In_214,In_1869);
xor U1069 (N_1069,In_1032,In_1744);
xnor U1070 (N_1070,In_1301,In_1800);
or U1071 (N_1071,In_682,In_754);
or U1072 (N_1072,In_1454,In_1115);
nand U1073 (N_1073,In_1246,In_1075);
and U1074 (N_1074,In_841,In_670);
nand U1075 (N_1075,In_140,In_868);
and U1076 (N_1076,In_219,In_141);
or U1077 (N_1077,In_345,In_1161);
and U1078 (N_1078,In_1517,In_856);
and U1079 (N_1079,In_866,In_1205);
or U1080 (N_1080,In_1924,In_836);
and U1081 (N_1081,In_122,In_11);
and U1082 (N_1082,In_949,In_1818);
or U1083 (N_1083,In_270,In_1833);
or U1084 (N_1084,In_1751,In_923);
nor U1085 (N_1085,In_365,In_1313);
nor U1086 (N_1086,In_818,In_1868);
nand U1087 (N_1087,In_130,In_1404);
or U1088 (N_1088,In_1309,In_349);
xor U1089 (N_1089,In_131,In_1546);
nor U1090 (N_1090,In_150,In_247);
or U1091 (N_1091,In_541,In_1236);
or U1092 (N_1092,In_694,In_747);
nand U1093 (N_1093,In_207,In_609);
and U1094 (N_1094,In_1407,In_678);
and U1095 (N_1095,In_268,In_1616);
xnor U1096 (N_1096,In_1586,In_1238);
xor U1097 (N_1097,In_676,In_1448);
nand U1098 (N_1098,In_377,In_480);
and U1099 (N_1099,In_1207,In_1034);
xor U1100 (N_1100,In_1583,In_1095);
or U1101 (N_1101,In_669,In_1551);
or U1102 (N_1102,In_867,In_735);
and U1103 (N_1103,In_1661,In_1167);
nor U1104 (N_1104,In_648,In_170);
and U1105 (N_1105,In_1543,In_1039);
nand U1106 (N_1106,In_1695,In_1813);
nor U1107 (N_1107,In_985,In_390);
nor U1108 (N_1108,In_1176,In_1331);
or U1109 (N_1109,In_1985,In_116);
xnor U1110 (N_1110,In_1138,In_1110);
nand U1111 (N_1111,In_1497,In_1338);
xnor U1112 (N_1112,In_702,In_530);
and U1113 (N_1113,In_1981,In_1331);
nand U1114 (N_1114,In_1851,In_1854);
and U1115 (N_1115,In_10,In_914);
and U1116 (N_1116,In_877,In_898);
or U1117 (N_1117,In_1783,In_1629);
nor U1118 (N_1118,In_817,In_1661);
xnor U1119 (N_1119,In_80,In_1750);
or U1120 (N_1120,In_1286,In_1903);
or U1121 (N_1121,In_1244,In_513);
xnor U1122 (N_1122,In_756,In_1993);
or U1123 (N_1123,In_555,In_899);
nand U1124 (N_1124,In_282,In_228);
and U1125 (N_1125,In_136,In_121);
xnor U1126 (N_1126,In_1051,In_906);
nand U1127 (N_1127,In_1465,In_769);
nor U1128 (N_1128,In_821,In_178);
nor U1129 (N_1129,In_689,In_1843);
nand U1130 (N_1130,In_320,In_106);
nor U1131 (N_1131,In_1496,In_72);
nand U1132 (N_1132,In_918,In_35);
or U1133 (N_1133,In_1310,In_427);
and U1134 (N_1134,In_783,In_531);
xnor U1135 (N_1135,In_1697,In_560);
nor U1136 (N_1136,In_120,In_699);
nor U1137 (N_1137,In_1514,In_155);
xnor U1138 (N_1138,In_1575,In_1065);
or U1139 (N_1139,In_1203,In_1168);
nand U1140 (N_1140,In_1789,In_100);
and U1141 (N_1141,In_719,In_1299);
and U1142 (N_1142,In_1645,In_949);
nand U1143 (N_1143,In_686,In_662);
xor U1144 (N_1144,In_189,In_1644);
nand U1145 (N_1145,In_266,In_454);
and U1146 (N_1146,In_1538,In_812);
or U1147 (N_1147,In_504,In_1371);
nor U1148 (N_1148,In_772,In_1494);
nand U1149 (N_1149,In_1357,In_1717);
and U1150 (N_1150,In_894,In_1987);
xor U1151 (N_1151,In_232,In_1383);
xor U1152 (N_1152,In_1187,In_821);
nand U1153 (N_1153,In_1897,In_928);
or U1154 (N_1154,In_1468,In_294);
nand U1155 (N_1155,In_1925,In_1157);
nor U1156 (N_1156,In_124,In_1130);
and U1157 (N_1157,In_1105,In_1024);
nand U1158 (N_1158,In_1257,In_895);
nor U1159 (N_1159,In_775,In_1139);
nand U1160 (N_1160,In_383,In_1195);
and U1161 (N_1161,In_585,In_1946);
xor U1162 (N_1162,In_1957,In_214);
xor U1163 (N_1163,In_867,In_334);
nor U1164 (N_1164,In_43,In_145);
xnor U1165 (N_1165,In_116,In_1734);
nand U1166 (N_1166,In_964,In_321);
and U1167 (N_1167,In_787,In_1589);
xnor U1168 (N_1168,In_1729,In_1464);
or U1169 (N_1169,In_363,In_1239);
and U1170 (N_1170,In_372,In_592);
and U1171 (N_1171,In_1362,In_1815);
nor U1172 (N_1172,In_1900,In_1826);
xor U1173 (N_1173,In_11,In_1671);
or U1174 (N_1174,In_252,In_1569);
or U1175 (N_1175,In_264,In_1885);
or U1176 (N_1176,In_1603,In_1595);
nand U1177 (N_1177,In_861,In_1025);
and U1178 (N_1178,In_332,In_1253);
and U1179 (N_1179,In_985,In_1670);
xor U1180 (N_1180,In_845,In_33);
xnor U1181 (N_1181,In_923,In_1990);
xnor U1182 (N_1182,In_902,In_697);
and U1183 (N_1183,In_977,In_791);
nand U1184 (N_1184,In_309,In_99);
nand U1185 (N_1185,In_1139,In_1328);
nand U1186 (N_1186,In_1049,In_202);
nand U1187 (N_1187,In_200,In_425);
or U1188 (N_1188,In_1622,In_1068);
xor U1189 (N_1189,In_918,In_249);
or U1190 (N_1190,In_1569,In_33);
nor U1191 (N_1191,In_1099,In_101);
xnor U1192 (N_1192,In_552,In_518);
or U1193 (N_1193,In_339,In_1097);
nand U1194 (N_1194,In_1856,In_1724);
nand U1195 (N_1195,In_664,In_456);
xor U1196 (N_1196,In_1326,In_743);
xor U1197 (N_1197,In_1250,In_551);
or U1198 (N_1198,In_1322,In_1369);
nor U1199 (N_1199,In_441,In_324);
nor U1200 (N_1200,In_889,In_978);
nor U1201 (N_1201,In_639,In_1720);
xnor U1202 (N_1202,In_496,In_1022);
xnor U1203 (N_1203,In_1542,In_341);
nand U1204 (N_1204,In_251,In_1845);
or U1205 (N_1205,In_1448,In_550);
and U1206 (N_1206,In_1199,In_1439);
xor U1207 (N_1207,In_119,In_1806);
and U1208 (N_1208,In_1165,In_426);
xnor U1209 (N_1209,In_124,In_1399);
xnor U1210 (N_1210,In_61,In_218);
xor U1211 (N_1211,In_864,In_530);
nor U1212 (N_1212,In_1877,In_1661);
nor U1213 (N_1213,In_363,In_620);
or U1214 (N_1214,In_147,In_942);
and U1215 (N_1215,In_543,In_0);
xor U1216 (N_1216,In_1697,In_1150);
or U1217 (N_1217,In_195,In_1222);
and U1218 (N_1218,In_1257,In_629);
nor U1219 (N_1219,In_1158,In_1990);
nor U1220 (N_1220,In_1945,In_903);
nand U1221 (N_1221,In_620,In_1800);
nor U1222 (N_1222,In_438,In_184);
and U1223 (N_1223,In_743,In_808);
or U1224 (N_1224,In_281,In_1126);
xor U1225 (N_1225,In_863,In_31);
xor U1226 (N_1226,In_759,In_1355);
and U1227 (N_1227,In_1315,In_1678);
or U1228 (N_1228,In_783,In_1318);
xnor U1229 (N_1229,In_1974,In_1858);
nand U1230 (N_1230,In_1518,In_1150);
nor U1231 (N_1231,In_1912,In_285);
nand U1232 (N_1232,In_1066,In_1344);
nor U1233 (N_1233,In_1766,In_1023);
and U1234 (N_1234,In_1664,In_839);
nand U1235 (N_1235,In_953,In_1145);
and U1236 (N_1236,In_1287,In_288);
or U1237 (N_1237,In_486,In_425);
nand U1238 (N_1238,In_332,In_1297);
xnor U1239 (N_1239,In_549,In_180);
xor U1240 (N_1240,In_1795,In_1264);
xor U1241 (N_1241,In_744,In_418);
or U1242 (N_1242,In_1270,In_1954);
and U1243 (N_1243,In_1326,In_1754);
or U1244 (N_1244,In_1144,In_1401);
xnor U1245 (N_1245,In_1282,In_1117);
xor U1246 (N_1246,In_1851,In_1202);
nand U1247 (N_1247,In_1883,In_639);
and U1248 (N_1248,In_873,In_1010);
nand U1249 (N_1249,In_1394,In_630);
and U1250 (N_1250,In_587,In_1650);
nand U1251 (N_1251,In_358,In_1012);
or U1252 (N_1252,In_704,In_483);
or U1253 (N_1253,In_877,In_470);
and U1254 (N_1254,In_1742,In_1582);
and U1255 (N_1255,In_1274,In_354);
xnor U1256 (N_1256,In_1246,In_272);
xnor U1257 (N_1257,In_1693,In_155);
nor U1258 (N_1258,In_266,In_1006);
or U1259 (N_1259,In_290,In_864);
nor U1260 (N_1260,In_733,In_517);
and U1261 (N_1261,In_309,In_1432);
nand U1262 (N_1262,In_1943,In_520);
nor U1263 (N_1263,In_548,In_563);
or U1264 (N_1264,In_1111,In_730);
xor U1265 (N_1265,In_1942,In_1936);
nand U1266 (N_1266,In_913,In_1220);
and U1267 (N_1267,In_1121,In_1360);
nor U1268 (N_1268,In_97,In_836);
nor U1269 (N_1269,In_308,In_1333);
nor U1270 (N_1270,In_382,In_83);
nand U1271 (N_1271,In_19,In_1797);
or U1272 (N_1272,In_932,In_1545);
nor U1273 (N_1273,In_803,In_552);
and U1274 (N_1274,In_643,In_1116);
nand U1275 (N_1275,In_1752,In_804);
nand U1276 (N_1276,In_1160,In_1104);
nor U1277 (N_1277,In_142,In_1106);
xor U1278 (N_1278,In_1642,In_578);
nor U1279 (N_1279,In_1328,In_1227);
nand U1280 (N_1280,In_130,In_1356);
and U1281 (N_1281,In_1097,In_1880);
xnor U1282 (N_1282,In_161,In_120);
xor U1283 (N_1283,In_1201,In_172);
or U1284 (N_1284,In_501,In_1875);
or U1285 (N_1285,In_1278,In_1470);
xor U1286 (N_1286,In_298,In_1005);
xor U1287 (N_1287,In_405,In_565);
nor U1288 (N_1288,In_940,In_1627);
or U1289 (N_1289,In_1914,In_639);
xor U1290 (N_1290,In_1763,In_1280);
and U1291 (N_1291,In_1858,In_1477);
xnor U1292 (N_1292,In_1689,In_1039);
nor U1293 (N_1293,In_159,In_489);
nand U1294 (N_1294,In_604,In_587);
or U1295 (N_1295,In_946,In_635);
xnor U1296 (N_1296,In_63,In_1965);
or U1297 (N_1297,In_906,In_1412);
nand U1298 (N_1298,In_858,In_35);
or U1299 (N_1299,In_551,In_1518);
xor U1300 (N_1300,In_1131,In_1205);
nand U1301 (N_1301,In_1074,In_1648);
nand U1302 (N_1302,In_1995,In_1171);
or U1303 (N_1303,In_1579,In_937);
and U1304 (N_1304,In_627,In_1435);
and U1305 (N_1305,In_1845,In_972);
xnor U1306 (N_1306,In_143,In_113);
and U1307 (N_1307,In_599,In_494);
and U1308 (N_1308,In_1056,In_1081);
xor U1309 (N_1309,In_1300,In_411);
nor U1310 (N_1310,In_416,In_269);
and U1311 (N_1311,In_1070,In_1102);
nor U1312 (N_1312,In_1114,In_25);
or U1313 (N_1313,In_648,In_1517);
nand U1314 (N_1314,In_1986,In_1014);
nand U1315 (N_1315,In_1147,In_194);
nor U1316 (N_1316,In_665,In_1362);
nand U1317 (N_1317,In_316,In_43);
xnor U1318 (N_1318,In_864,In_332);
and U1319 (N_1319,In_1634,In_1130);
and U1320 (N_1320,In_331,In_1112);
nor U1321 (N_1321,In_7,In_1391);
nand U1322 (N_1322,In_758,In_368);
or U1323 (N_1323,In_705,In_75);
and U1324 (N_1324,In_1889,In_345);
and U1325 (N_1325,In_1918,In_327);
or U1326 (N_1326,In_1947,In_232);
nand U1327 (N_1327,In_1901,In_1688);
nand U1328 (N_1328,In_1589,In_1278);
nor U1329 (N_1329,In_1061,In_1167);
nor U1330 (N_1330,In_1170,In_1369);
nor U1331 (N_1331,In_1224,In_1226);
xor U1332 (N_1332,In_1614,In_1984);
and U1333 (N_1333,In_378,In_1357);
or U1334 (N_1334,In_74,In_221);
xnor U1335 (N_1335,In_293,In_544);
nor U1336 (N_1336,In_1025,In_392);
nor U1337 (N_1337,In_63,In_1824);
nand U1338 (N_1338,In_1974,In_1833);
or U1339 (N_1339,In_724,In_1200);
or U1340 (N_1340,In_417,In_1481);
xnor U1341 (N_1341,In_1974,In_731);
and U1342 (N_1342,In_1110,In_1606);
and U1343 (N_1343,In_1674,In_736);
xor U1344 (N_1344,In_160,In_936);
and U1345 (N_1345,In_1724,In_632);
and U1346 (N_1346,In_1331,In_257);
xnor U1347 (N_1347,In_454,In_978);
or U1348 (N_1348,In_264,In_801);
nor U1349 (N_1349,In_1603,In_1288);
nor U1350 (N_1350,In_1792,In_1589);
or U1351 (N_1351,In_1372,In_1276);
nand U1352 (N_1352,In_187,In_810);
nor U1353 (N_1353,In_1657,In_1399);
nand U1354 (N_1354,In_1597,In_1371);
and U1355 (N_1355,In_21,In_437);
xnor U1356 (N_1356,In_119,In_649);
and U1357 (N_1357,In_100,In_1899);
xnor U1358 (N_1358,In_334,In_974);
nor U1359 (N_1359,In_1868,In_1988);
xnor U1360 (N_1360,In_1584,In_228);
and U1361 (N_1361,In_109,In_1537);
xor U1362 (N_1362,In_168,In_960);
and U1363 (N_1363,In_1606,In_151);
and U1364 (N_1364,In_1102,In_170);
nand U1365 (N_1365,In_1980,In_39);
nand U1366 (N_1366,In_1351,In_530);
and U1367 (N_1367,In_1698,In_1467);
nand U1368 (N_1368,In_1949,In_1233);
xnor U1369 (N_1369,In_1699,In_344);
nand U1370 (N_1370,In_1134,In_249);
or U1371 (N_1371,In_993,In_743);
and U1372 (N_1372,In_631,In_1569);
xor U1373 (N_1373,In_1087,In_632);
xnor U1374 (N_1374,In_1369,In_1848);
nor U1375 (N_1375,In_786,In_1574);
or U1376 (N_1376,In_912,In_1977);
xor U1377 (N_1377,In_1954,In_1227);
xor U1378 (N_1378,In_1518,In_1491);
nand U1379 (N_1379,In_1495,In_990);
and U1380 (N_1380,In_325,In_1993);
nor U1381 (N_1381,In_507,In_429);
nor U1382 (N_1382,In_834,In_577);
or U1383 (N_1383,In_800,In_344);
nor U1384 (N_1384,In_1912,In_54);
or U1385 (N_1385,In_711,In_1551);
nor U1386 (N_1386,In_638,In_1157);
or U1387 (N_1387,In_720,In_254);
and U1388 (N_1388,In_892,In_641);
or U1389 (N_1389,In_1759,In_1733);
xor U1390 (N_1390,In_1325,In_1329);
xnor U1391 (N_1391,In_704,In_1925);
and U1392 (N_1392,In_1454,In_513);
xnor U1393 (N_1393,In_823,In_1367);
xor U1394 (N_1394,In_31,In_6);
or U1395 (N_1395,In_961,In_1571);
or U1396 (N_1396,In_933,In_428);
xnor U1397 (N_1397,In_924,In_736);
and U1398 (N_1398,In_525,In_1015);
xnor U1399 (N_1399,In_723,In_320);
and U1400 (N_1400,In_1204,In_1810);
xnor U1401 (N_1401,In_801,In_1598);
nand U1402 (N_1402,In_848,In_487);
xnor U1403 (N_1403,In_522,In_1790);
nand U1404 (N_1404,In_1318,In_1205);
or U1405 (N_1405,In_1215,In_968);
nor U1406 (N_1406,In_677,In_277);
and U1407 (N_1407,In_1055,In_1703);
nand U1408 (N_1408,In_1202,In_1516);
xnor U1409 (N_1409,In_1573,In_1973);
nor U1410 (N_1410,In_1501,In_866);
nand U1411 (N_1411,In_421,In_191);
nor U1412 (N_1412,In_775,In_447);
nand U1413 (N_1413,In_1044,In_826);
and U1414 (N_1414,In_358,In_975);
nand U1415 (N_1415,In_1050,In_1486);
and U1416 (N_1416,In_920,In_606);
and U1417 (N_1417,In_1760,In_812);
and U1418 (N_1418,In_1655,In_1303);
nor U1419 (N_1419,In_878,In_664);
xnor U1420 (N_1420,In_310,In_434);
and U1421 (N_1421,In_457,In_117);
xor U1422 (N_1422,In_1632,In_836);
or U1423 (N_1423,In_1734,In_1480);
and U1424 (N_1424,In_1614,In_1608);
nand U1425 (N_1425,In_1347,In_1709);
and U1426 (N_1426,In_1290,In_1813);
nand U1427 (N_1427,In_812,In_1381);
xor U1428 (N_1428,In_955,In_22);
or U1429 (N_1429,In_1130,In_1466);
or U1430 (N_1430,In_775,In_1789);
nand U1431 (N_1431,In_693,In_992);
nand U1432 (N_1432,In_1461,In_900);
xnor U1433 (N_1433,In_987,In_1287);
nor U1434 (N_1434,In_1084,In_1100);
nand U1435 (N_1435,In_550,In_522);
nor U1436 (N_1436,In_409,In_1312);
or U1437 (N_1437,In_1523,In_262);
xnor U1438 (N_1438,In_163,In_982);
nand U1439 (N_1439,In_1903,In_1239);
or U1440 (N_1440,In_962,In_601);
and U1441 (N_1441,In_1676,In_198);
nand U1442 (N_1442,In_940,In_1369);
or U1443 (N_1443,In_1985,In_322);
nand U1444 (N_1444,In_1081,In_509);
and U1445 (N_1445,In_1407,In_42);
nor U1446 (N_1446,In_38,In_15);
nor U1447 (N_1447,In_120,In_1112);
or U1448 (N_1448,In_260,In_1116);
and U1449 (N_1449,In_1271,In_189);
nand U1450 (N_1450,In_971,In_139);
and U1451 (N_1451,In_10,In_498);
or U1452 (N_1452,In_403,In_340);
nand U1453 (N_1453,In_1743,In_534);
nor U1454 (N_1454,In_755,In_850);
nand U1455 (N_1455,In_32,In_1076);
xnor U1456 (N_1456,In_1309,In_1331);
nor U1457 (N_1457,In_1779,In_1553);
nand U1458 (N_1458,In_1488,In_1396);
nand U1459 (N_1459,In_976,In_709);
or U1460 (N_1460,In_1063,In_1349);
and U1461 (N_1461,In_1552,In_1234);
and U1462 (N_1462,In_770,In_877);
nor U1463 (N_1463,In_440,In_108);
xnor U1464 (N_1464,In_437,In_1343);
nand U1465 (N_1465,In_1882,In_914);
or U1466 (N_1466,In_815,In_1917);
xnor U1467 (N_1467,In_1500,In_189);
or U1468 (N_1468,In_923,In_1783);
nand U1469 (N_1469,In_783,In_1458);
nand U1470 (N_1470,In_1151,In_50);
or U1471 (N_1471,In_1122,In_736);
xor U1472 (N_1472,In_272,In_569);
and U1473 (N_1473,In_778,In_358);
or U1474 (N_1474,In_72,In_228);
and U1475 (N_1475,In_560,In_1544);
nor U1476 (N_1476,In_595,In_242);
xnor U1477 (N_1477,In_224,In_1408);
or U1478 (N_1478,In_1451,In_1241);
or U1479 (N_1479,In_340,In_561);
xnor U1480 (N_1480,In_1706,In_1866);
or U1481 (N_1481,In_1398,In_386);
nor U1482 (N_1482,In_796,In_855);
and U1483 (N_1483,In_1639,In_126);
or U1484 (N_1484,In_1117,In_1491);
or U1485 (N_1485,In_881,In_507);
and U1486 (N_1486,In_775,In_10);
or U1487 (N_1487,In_985,In_1624);
nor U1488 (N_1488,In_1862,In_235);
and U1489 (N_1489,In_1087,In_1616);
and U1490 (N_1490,In_1287,In_912);
and U1491 (N_1491,In_784,In_714);
xor U1492 (N_1492,In_1905,In_1760);
or U1493 (N_1493,In_1032,In_1800);
xnor U1494 (N_1494,In_1591,In_521);
nand U1495 (N_1495,In_412,In_1508);
or U1496 (N_1496,In_339,In_1992);
xnor U1497 (N_1497,In_1761,In_1335);
nand U1498 (N_1498,In_581,In_833);
and U1499 (N_1499,In_596,In_200);
nor U1500 (N_1500,In_170,In_1709);
or U1501 (N_1501,In_1831,In_245);
nand U1502 (N_1502,In_1104,In_682);
xor U1503 (N_1503,In_800,In_1121);
xor U1504 (N_1504,In_567,In_653);
nand U1505 (N_1505,In_249,In_1656);
and U1506 (N_1506,In_1244,In_1139);
xor U1507 (N_1507,In_1585,In_1974);
nor U1508 (N_1508,In_1795,In_1996);
xor U1509 (N_1509,In_1737,In_1298);
nor U1510 (N_1510,In_1417,In_525);
xnor U1511 (N_1511,In_1986,In_286);
nand U1512 (N_1512,In_1415,In_424);
and U1513 (N_1513,In_520,In_1068);
xor U1514 (N_1514,In_1218,In_1426);
xor U1515 (N_1515,In_1665,In_186);
and U1516 (N_1516,In_1444,In_756);
xnor U1517 (N_1517,In_772,In_1241);
nand U1518 (N_1518,In_1181,In_790);
xnor U1519 (N_1519,In_1626,In_910);
nor U1520 (N_1520,In_1989,In_848);
xor U1521 (N_1521,In_812,In_116);
and U1522 (N_1522,In_1015,In_1375);
or U1523 (N_1523,In_1520,In_266);
or U1524 (N_1524,In_558,In_1644);
and U1525 (N_1525,In_354,In_697);
nand U1526 (N_1526,In_502,In_936);
or U1527 (N_1527,In_898,In_1271);
nor U1528 (N_1528,In_28,In_435);
or U1529 (N_1529,In_1087,In_1689);
xnor U1530 (N_1530,In_1795,In_584);
and U1531 (N_1531,In_907,In_913);
and U1532 (N_1532,In_1071,In_960);
nor U1533 (N_1533,In_1232,In_1467);
and U1534 (N_1534,In_450,In_467);
and U1535 (N_1535,In_699,In_620);
or U1536 (N_1536,In_656,In_1380);
nand U1537 (N_1537,In_993,In_398);
xnor U1538 (N_1538,In_1499,In_717);
nand U1539 (N_1539,In_1655,In_1099);
and U1540 (N_1540,In_1771,In_1459);
nand U1541 (N_1541,In_284,In_301);
nand U1542 (N_1542,In_1099,In_641);
xnor U1543 (N_1543,In_399,In_1182);
or U1544 (N_1544,In_321,In_1524);
xor U1545 (N_1545,In_859,In_1907);
nor U1546 (N_1546,In_1378,In_888);
and U1547 (N_1547,In_1149,In_853);
and U1548 (N_1548,In_178,In_1754);
xnor U1549 (N_1549,In_1735,In_1924);
and U1550 (N_1550,In_1864,In_1419);
nor U1551 (N_1551,In_1668,In_506);
nand U1552 (N_1552,In_1840,In_202);
nor U1553 (N_1553,In_1813,In_1186);
xor U1554 (N_1554,In_973,In_540);
and U1555 (N_1555,In_667,In_1023);
xor U1556 (N_1556,In_1776,In_1514);
nor U1557 (N_1557,In_485,In_1631);
or U1558 (N_1558,In_1928,In_701);
xnor U1559 (N_1559,In_1360,In_1701);
nor U1560 (N_1560,In_1584,In_1094);
xor U1561 (N_1561,In_215,In_894);
nor U1562 (N_1562,In_339,In_765);
nor U1563 (N_1563,In_497,In_1110);
xnor U1564 (N_1564,In_1500,In_392);
and U1565 (N_1565,In_925,In_1818);
nor U1566 (N_1566,In_242,In_1395);
nor U1567 (N_1567,In_1511,In_20);
and U1568 (N_1568,In_727,In_1691);
nor U1569 (N_1569,In_201,In_1693);
or U1570 (N_1570,In_1427,In_1937);
or U1571 (N_1571,In_1304,In_879);
nand U1572 (N_1572,In_1342,In_1799);
nand U1573 (N_1573,In_208,In_512);
and U1574 (N_1574,In_228,In_531);
nor U1575 (N_1575,In_1580,In_1257);
xor U1576 (N_1576,In_1695,In_940);
nor U1577 (N_1577,In_799,In_1586);
nand U1578 (N_1578,In_1567,In_331);
nor U1579 (N_1579,In_559,In_1540);
xor U1580 (N_1580,In_70,In_1968);
xor U1581 (N_1581,In_1908,In_1757);
xor U1582 (N_1582,In_1408,In_1744);
xor U1583 (N_1583,In_1292,In_330);
nand U1584 (N_1584,In_1558,In_545);
and U1585 (N_1585,In_475,In_1430);
or U1586 (N_1586,In_1719,In_1940);
nand U1587 (N_1587,In_966,In_1838);
nand U1588 (N_1588,In_229,In_1103);
and U1589 (N_1589,In_152,In_1276);
and U1590 (N_1590,In_1802,In_930);
or U1591 (N_1591,In_1394,In_820);
or U1592 (N_1592,In_749,In_971);
nor U1593 (N_1593,In_567,In_627);
xnor U1594 (N_1594,In_552,In_195);
and U1595 (N_1595,In_207,In_497);
xnor U1596 (N_1596,In_1200,In_1758);
xnor U1597 (N_1597,In_1630,In_1538);
nor U1598 (N_1598,In_549,In_1133);
and U1599 (N_1599,In_1833,In_948);
or U1600 (N_1600,In_883,In_50);
or U1601 (N_1601,In_1103,In_342);
nor U1602 (N_1602,In_1927,In_1412);
xnor U1603 (N_1603,In_913,In_691);
and U1604 (N_1604,In_1080,In_142);
and U1605 (N_1605,In_1984,In_1565);
and U1606 (N_1606,In_762,In_976);
or U1607 (N_1607,In_647,In_1333);
nand U1608 (N_1608,In_1053,In_578);
and U1609 (N_1609,In_337,In_1976);
xor U1610 (N_1610,In_298,In_1679);
xnor U1611 (N_1611,In_1266,In_1306);
nand U1612 (N_1612,In_1753,In_1227);
nor U1613 (N_1613,In_1873,In_973);
or U1614 (N_1614,In_58,In_1396);
nand U1615 (N_1615,In_1875,In_1393);
nand U1616 (N_1616,In_1715,In_744);
nor U1617 (N_1617,In_1137,In_359);
nor U1618 (N_1618,In_1275,In_1450);
nand U1619 (N_1619,In_363,In_718);
and U1620 (N_1620,In_60,In_853);
nor U1621 (N_1621,In_717,In_1296);
or U1622 (N_1622,In_85,In_1119);
and U1623 (N_1623,In_634,In_1024);
nor U1624 (N_1624,In_1362,In_1562);
nor U1625 (N_1625,In_899,In_201);
and U1626 (N_1626,In_791,In_86);
nor U1627 (N_1627,In_1059,In_1380);
or U1628 (N_1628,In_1508,In_713);
xnor U1629 (N_1629,In_368,In_1530);
nand U1630 (N_1630,In_866,In_1282);
nand U1631 (N_1631,In_1323,In_1092);
or U1632 (N_1632,In_109,In_735);
or U1633 (N_1633,In_1593,In_856);
nand U1634 (N_1634,In_105,In_999);
nor U1635 (N_1635,In_1238,In_1013);
xnor U1636 (N_1636,In_1492,In_1341);
nand U1637 (N_1637,In_749,In_1243);
or U1638 (N_1638,In_1346,In_1727);
nand U1639 (N_1639,In_1855,In_898);
nor U1640 (N_1640,In_908,In_1971);
nand U1641 (N_1641,In_1941,In_383);
or U1642 (N_1642,In_1088,In_593);
nor U1643 (N_1643,In_1468,In_1226);
xnor U1644 (N_1644,In_1868,In_731);
nand U1645 (N_1645,In_551,In_634);
and U1646 (N_1646,In_296,In_1413);
nand U1647 (N_1647,In_1522,In_1137);
nor U1648 (N_1648,In_1409,In_1796);
nand U1649 (N_1649,In_1435,In_1576);
and U1650 (N_1650,In_1338,In_830);
and U1651 (N_1651,In_1722,In_739);
xor U1652 (N_1652,In_521,In_1645);
nand U1653 (N_1653,In_1755,In_577);
nor U1654 (N_1654,In_1032,In_224);
or U1655 (N_1655,In_1688,In_516);
xor U1656 (N_1656,In_244,In_437);
and U1657 (N_1657,In_815,In_330);
or U1658 (N_1658,In_1669,In_675);
and U1659 (N_1659,In_1783,In_1661);
nor U1660 (N_1660,In_1122,In_363);
nor U1661 (N_1661,In_1451,In_1642);
and U1662 (N_1662,In_840,In_210);
nand U1663 (N_1663,In_802,In_1938);
xnor U1664 (N_1664,In_1625,In_1669);
or U1665 (N_1665,In_1297,In_1504);
xor U1666 (N_1666,In_1572,In_1930);
or U1667 (N_1667,In_1779,In_1997);
nor U1668 (N_1668,In_1251,In_16);
nand U1669 (N_1669,In_1136,In_631);
nor U1670 (N_1670,In_400,In_1341);
xor U1671 (N_1671,In_1921,In_815);
nand U1672 (N_1672,In_1361,In_1236);
and U1673 (N_1673,In_1556,In_1101);
nand U1674 (N_1674,In_646,In_94);
and U1675 (N_1675,In_1954,In_362);
or U1676 (N_1676,In_1448,In_331);
nor U1677 (N_1677,In_1846,In_1690);
or U1678 (N_1678,In_1637,In_935);
nor U1679 (N_1679,In_470,In_309);
and U1680 (N_1680,In_352,In_596);
or U1681 (N_1681,In_1313,In_1133);
nand U1682 (N_1682,In_1204,In_1469);
and U1683 (N_1683,In_338,In_239);
nand U1684 (N_1684,In_1671,In_1627);
and U1685 (N_1685,In_324,In_100);
nand U1686 (N_1686,In_256,In_192);
nor U1687 (N_1687,In_1582,In_724);
nor U1688 (N_1688,In_955,In_1680);
and U1689 (N_1689,In_220,In_195);
nand U1690 (N_1690,In_1751,In_198);
xor U1691 (N_1691,In_1913,In_1972);
nand U1692 (N_1692,In_1932,In_1810);
and U1693 (N_1693,In_676,In_1274);
or U1694 (N_1694,In_1963,In_1875);
nor U1695 (N_1695,In_1380,In_1784);
nor U1696 (N_1696,In_1824,In_1115);
xnor U1697 (N_1697,In_129,In_120);
xnor U1698 (N_1698,In_34,In_232);
and U1699 (N_1699,In_1414,In_453);
nand U1700 (N_1700,In_878,In_905);
nand U1701 (N_1701,In_749,In_336);
or U1702 (N_1702,In_727,In_1927);
nor U1703 (N_1703,In_459,In_1970);
xor U1704 (N_1704,In_1755,In_1448);
nand U1705 (N_1705,In_1441,In_1921);
or U1706 (N_1706,In_425,In_253);
and U1707 (N_1707,In_1960,In_1649);
nand U1708 (N_1708,In_1011,In_1565);
xnor U1709 (N_1709,In_1112,In_1764);
nand U1710 (N_1710,In_1345,In_1911);
nand U1711 (N_1711,In_114,In_432);
nand U1712 (N_1712,In_1177,In_904);
or U1713 (N_1713,In_1388,In_919);
or U1714 (N_1714,In_1988,In_1239);
xor U1715 (N_1715,In_1117,In_1190);
nand U1716 (N_1716,In_1839,In_476);
nand U1717 (N_1717,In_1948,In_1048);
xor U1718 (N_1718,In_280,In_354);
nand U1719 (N_1719,In_703,In_1298);
xnor U1720 (N_1720,In_892,In_1128);
nand U1721 (N_1721,In_1574,In_1807);
and U1722 (N_1722,In_11,In_31);
xor U1723 (N_1723,In_282,In_146);
nand U1724 (N_1724,In_596,In_718);
nand U1725 (N_1725,In_828,In_1206);
or U1726 (N_1726,In_49,In_1910);
xor U1727 (N_1727,In_973,In_506);
and U1728 (N_1728,In_29,In_947);
nor U1729 (N_1729,In_1814,In_219);
xor U1730 (N_1730,In_1087,In_965);
and U1731 (N_1731,In_1700,In_848);
nor U1732 (N_1732,In_1207,In_1845);
or U1733 (N_1733,In_271,In_274);
and U1734 (N_1734,In_1463,In_506);
nand U1735 (N_1735,In_1606,In_1838);
nand U1736 (N_1736,In_319,In_171);
or U1737 (N_1737,In_1664,In_1339);
or U1738 (N_1738,In_494,In_1100);
nand U1739 (N_1739,In_201,In_1870);
nand U1740 (N_1740,In_1363,In_1288);
and U1741 (N_1741,In_1708,In_292);
xnor U1742 (N_1742,In_1268,In_122);
and U1743 (N_1743,In_460,In_608);
xnor U1744 (N_1744,In_82,In_1873);
xor U1745 (N_1745,In_1385,In_1321);
nand U1746 (N_1746,In_735,In_1118);
or U1747 (N_1747,In_1387,In_829);
nand U1748 (N_1748,In_584,In_347);
nor U1749 (N_1749,In_1416,In_536);
nor U1750 (N_1750,In_1037,In_1956);
nand U1751 (N_1751,In_393,In_1763);
xor U1752 (N_1752,In_1530,In_68);
and U1753 (N_1753,In_1701,In_452);
and U1754 (N_1754,In_1648,In_1508);
xor U1755 (N_1755,In_1453,In_1649);
and U1756 (N_1756,In_1264,In_1136);
nor U1757 (N_1757,In_282,In_759);
and U1758 (N_1758,In_1724,In_1126);
xnor U1759 (N_1759,In_41,In_697);
xnor U1760 (N_1760,In_624,In_677);
or U1761 (N_1761,In_1561,In_1124);
nor U1762 (N_1762,In_1919,In_833);
nand U1763 (N_1763,In_418,In_1372);
nor U1764 (N_1764,In_242,In_1249);
xor U1765 (N_1765,In_1786,In_1711);
nand U1766 (N_1766,In_816,In_1315);
and U1767 (N_1767,In_173,In_138);
xor U1768 (N_1768,In_753,In_906);
nor U1769 (N_1769,In_1623,In_1352);
xnor U1770 (N_1770,In_1374,In_368);
nor U1771 (N_1771,In_905,In_115);
or U1772 (N_1772,In_317,In_1167);
xor U1773 (N_1773,In_792,In_1112);
nand U1774 (N_1774,In_1875,In_7);
xor U1775 (N_1775,In_545,In_234);
and U1776 (N_1776,In_920,In_1463);
xor U1777 (N_1777,In_755,In_1358);
xor U1778 (N_1778,In_282,In_1773);
nor U1779 (N_1779,In_966,In_640);
or U1780 (N_1780,In_1174,In_113);
and U1781 (N_1781,In_741,In_1542);
and U1782 (N_1782,In_67,In_700);
or U1783 (N_1783,In_333,In_1614);
or U1784 (N_1784,In_1044,In_726);
and U1785 (N_1785,In_1072,In_856);
and U1786 (N_1786,In_551,In_4);
xor U1787 (N_1787,In_1024,In_1008);
and U1788 (N_1788,In_942,In_270);
and U1789 (N_1789,In_1550,In_1159);
nor U1790 (N_1790,In_179,In_1702);
xor U1791 (N_1791,In_954,In_1958);
xor U1792 (N_1792,In_1532,In_165);
and U1793 (N_1793,In_1123,In_608);
nor U1794 (N_1794,In_1820,In_97);
and U1795 (N_1795,In_1292,In_970);
nand U1796 (N_1796,In_625,In_1817);
nor U1797 (N_1797,In_1687,In_1318);
xor U1798 (N_1798,In_1167,In_21);
nor U1799 (N_1799,In_794,In_1643);
and U1800 (N_1800,In_1428,In_1731);
and U1801 (N_1801,In_358,In_654);
nor U1802 (N_1802,In_1964,In_1250);
and U1803 (N_1803,In_1096,In_1604);
and U1804 (N_1804,In_1364,In_894);
xnor U1805 (N_1805,In_1471,In_142);
or U1806 (N_1806,In_899,In_1955);
or U1807 (N_1807,In_113,In_1035);
and U1808 (N_1808,In_915,In_1256);
nor U1809 (N_1809,In_851,In_246);
nor U1810 (N_1810,In_12,In_1669);
nor U1811 (N_1811,In_821,In_1276);
nand U1812 (N_1812,In_705,In_678);
xor U1813 (N_1813,In_1844,In_230);
nand U1814 (N_1814,In_1312,In_1894);
xnor U1815 (N_1815,In_1529,In_1772);
and U1816 (N_1816,In_1110,In_1723);
nand U1817 (N_1817,In_557,In_1632);
nor U1818 (N_1818,In_61,In_1518);
and U1819 (N_1819,In_1698,In_415);
nor U1820 (N_1820,In_1354,In_1840);
nand U1821 (N_1821,In_156,In_1563);
nor U1822 (N_1822,In_1825,In_1687);
nand U1823 (N_1823,In_536,In_798);
xor U1824 (N_1824,In_908,In_1746);
nand U1825 (N_1825,In_1339,In_1323);
nor U1826 (N_1826,In_1871,In_1447);
nor U1827 (N_1827,In_141,In_1724);
or U1828 (N_1828,In_488,In_158);
xor U1829 (N_1829,In_915,In_286);
nand U1830 (N_1830,In_1795,In_1767);
nor U1831 (N_1831,In_1742,In_404);
or U1832 (N_1832,In_724,In_1689);
nor U1833 (N_1833,In_68,In_897);
or U1834 (N_1834,In_1778,In_178);
nor U1835 (N_1835,In_336,In_286);
nand U1836 (N_1836,In_607,In_937);
and U1837 (N_1837,In_257,In_425);
xnor U1838 (N_1838,In_1950,In_1105);
or U1839 (N_1839,In_1817,In_1920);
nor U1840 (N_1840,In_1089,In_414);
xor U1841 (N_1841,In_993,In_666);
xor U1842 (N_1842,In_1109,In_494);
nor U1843 (N_1843,In_1965,In_1502);
xnor U1844 (N_1844,In_1847,In_1292);
xnor U1845 (N_1845,In_1109,In_164);
xnor U1846 (N_1846,In_229,In_1623);
xor U1847 (N_1847,In_1004,In_1324);
nor U1848 (N_1848,In_1016,In_350);
nor U1849 (N_1849,In_701,In_470);
and U1850 (N_1850,In_712,In_1408);
and U1851 (N_1851,In_1993,In_992);
nand U1852 (N_1852,In_1692,In_1788);
and U1853 (N_1853,In_1086,In_1653);
nor U1854 (N_1854,In_1117,In_779);
xnor U1855 (N_1855,In_1983,In_605);
nand U1856 (N_1856,In_963,In_69);
and U1857 (N_1857,In_1389,In_471);
nand U1858 (N_1858,In_814,In_254);
or U1859 (N_1859,In_1089,In_1960);
or U1860 (N_1860,In_1663,In_1037);
nand U1861 (N_1861,In_1538,In_1955);
nand U1862 (N_1862,In_140,In_1751);
and U1863 (N_1863,In_399,In_417);
nor U1864 (N_1864,In_522,In_1600);
nand U1865 (N_1865,In_801,In_618);
nor U1866 (N_1866,In_1953,In_104);
nand U1867 (N_1867,In_514,In_347);
xor U1868 (N_1868,In_1389,In_1045);
or U1869 (N_1869,In_157,In_1901);
nor U1870 (N_1870,In_1553,In_387);
nor U1871 (N_1871,In_727,In_1452);
nand U1872 (N_1872,In_786,In_740);
and U1873 (N_1873,In_702,In_1878);
or U1874 (N_1874,In_18,In_1593);
nand U1875 (N_1875,In_352,In_975);
or U1876 (N_1876,In_1599,In_1958);
and U1877 (N_1877,In_425,In_1987);
xor U1878 (N_1878,In_30,In_1131);
and U1879 (N_1879,In_475,In_1136);
nor U1880 (N_1880,In_827,In_1825);
or U1881 (N_1881,In_739,In_1943);
xnor U1882 (N_1882,In_1238,In_1195);
and U1883 (N_1883,In_1149,In_1682);
nand U1884 (N_1884,In_1590,In_996);
nand U1885 (N_1885,In_115,In_705);
or U1886 (N_1886,In_474,In_1195);
xor U1887 (N_1887,In_191,In_1882);
xor U1888 (N_1888,In_195,In_1351);
xnor U1889 (N_1889,In_1475,In_1529);
xor U1890 (N_1890,In_65,In_1429);
nor U1891 (N_1891,In_1616,In_110);
nor U1892 (N_1892,In_1981,In_1034);
nand U1893 (N_1893,In_490,In_891);
nor U1894 (N_1894,In_629,In_428);
nand U1895 (N_1895,In_425,In_1681);
and U1896 (N_1896,In_1222,In_61);
or U1897 (N_1897,In_110,In_1128);
xnor U1898 (N_1898,In_768,In_1751);
nor U1899 (N_1899,In_649,In_1543);
nor U1900 (N_1900,In_225,In_816);
nand U1901 (N_1901,In_1574,In_387);
or U1902 (N_1902,In_336,In_1486);
or U1903 (N_1903,In_873,In_1559);
xor U1904 (N_1904,In_247,In_278);
nor U1905 (N_1905,In_38,In_903);
nor U1906 (N_1906,In_224,In_1239);
and U1907 (N_1907,In_1488,In_1570);
and U1908 (N_1908,In_681,In_1925);
or U1909 (N_1909,In_927,In_1452);
nand U1910 (N_1910,In_1174,In_1841);
or U1911 (N_1911,In_384,In_396);
and U1912 (N_1912,In_1420,In_337);
xor U1913 (N_1913,In_247,In_708);
xor U1914 (N_1914,In_235,In_437);
nand U1915 (N_1915,In_1789,In_1008);
nor U1916 (N_1916,In_1385,In_587);
nand U1917 (N_1917,In_1722,In_165);
nor U1918 (N_1918,In_826,In_401);
nand U1919 (N_1919,In_480,In_932);
xnor U1920 (N_1920,In_1485,In_715);
nand U1921 (N_1921,In_1105,In_1330);
nor U1922 (N_1922,In_1347,In_1235);
or U1923 (N_1923,In_1616,In_916);
or U1924 (N_1924,In_1601,In_177);
and U1925 (N_1925,In_821,In_119);
nand U1926 (N_1926,In_1638,In_730);
xor U1927 (N_1927,In_737,In_1277);
nor U1928 (N_1928,In_760,In_356);
and U1929 (N_1929,In_140,In_1471);
nand U1930 (N_1930,In_1519,In_667);
xnor U1931 (N_1931,In_1920,In_1540);
nor U1932 (N_1932,In_1181,In_858);
xor U1933 (N_1933,In_118,In_1736);
xor U1934 (N_1934,In_1015,In_343);
or U1935 (N_1935,In_1466,In_1390);
nand U1936 (N_1936,In_398,In_809);
nor U1937 (N_1937,In_310,In_57);
xor U1938 (N_1938,In_850,In_60);
nand U1939 (N_1939,In_147,In_41);
xnor U1940 (N_1940,In_1538,In_895);
nand U1941 (N_1941,In_1538,In_923);
and U1942 (N_1942,In_1078,In_1371);
nand U1943 (N_1943,In_1502,In_729);
and U1944 (N_1944,In_17,In_47);
or U1945 (N_1945,In_365,In_966);
nor U1946 (N_1946,In_414,In_419);
nand U1947 (N_1947,In_756,In_466);
and U1948 (N_1948,In_794,In_740);
xor U1949 (N_1949,In_87,In_437);
nand U1950 (N_1950,In_1983,In_724);
and U1951 (N_1951,In_254,In_1294);
xnor U1952 (N_1952,In_553,In_999);
nor U1953 (N_1953,In_1898,In_1759);
or U1954 (N_1954,In_181,In_1087);
xnor U1955 (N_1955,In_553,In_136);
nand U1956 (N_1956,In_1001,In_1432);
or U1957 (N_1957,In_1801,In_551);
nor U1958 (N_1958,In_704,In_1572);
nor U1959 (N_1959,In_184,In_289);
xnor U1960 (N_1960,In_1827,In_920);
or U1961 (N_1961,In_1138,In_67);
nor U1962 (N_1962,In_743,In_784);
and U1963 (N_1963,In_1343,In_145);
xor U1964 (N_1964,In_1401,In_963);
or U1965 (N_1965,In_1667,In_1922);
nand U1966 (N_1966,In_1751,In_741);
xnor U1967 (N_1967,In_1967,In_312);
nor U1968 (N_1968,In_873,In_1794);
or U1969 (N_1969,In_1471,In_175);
and U1970 (N_1970,In_791,In_1215);
nor U1971 (N_1971,In_1143,In_487);
nand U1972 (N_1972,In_1130,In_676);
nand U1973 (N_1973,In_1265,In_1301);
nand U1974 (N_1974,In_182,In_399);
and U1975 (N_1975,In_1327,In_1867);
and U1976 (N_1976,In_1511,In_1387);
nor U1977 (N_1977,In_976,In_1661);
nand U1978 (N_1978,In_34,In_834);
xnor U1979 (N_1979,In_1892,In_1930);
nor U1980 (N_1980,In_998,In_1034);
or U1981 (N_1981,In_1342,In_810);
or U1982 (N_1982,In_744,In_20);
nand U1983 (N_1983,In_976,In_1812);
nor U1984 (N_1984,In_752,In_1071);
nor U1985 (N_1985,In_1070,In_591);
and U1986 (N_1986,In_1107,In_11);
xor U1987 (N_1987,In_1603,In_870);
xor U1988 (N_1988,In_1960,In_1877);
xor U1989 (N_1989,In_151,In_721);
nand U1990 (N_1990,In_963,In_1782);
nor U1991 (N_1991,In_205,In_1944);
xnor U1992 (N_1992,In_1251,In_448);
nor U1993 (N_1993,In_1212,In_1415);
xnor U1994 (N_1994,In_1020,In_351);
xnor U1995 (N_1995,In_1496,In_1177);
nand U1996 (N_1996,In_1299,In_1654);
xor U1997 (N_1997,In_14,In_1074);
xnor U1998 (N_1998,In_1198,In_1904);
xnor U1999 (N_1999,In_448,In_1230);
nand U2000 (N_2000,In_1432,In_1681);
nor U2001 (N_2001,In_1657,In_1523);
xnor U2002 (N_2002,In_514,In_990);
or U2003 (N_2003,In_564,In_638);
or U2004 (N_2004,In_386,In_1436);
xor U2005 (N_2005,In_925,In_946);
or U2006 (N_2006,In_1155,In_1172);
or U2007 (N_2007,In_89,In_903);
and U2008 (N_2008,In_967,In_554);
or U2009 (N_2009,In_1108,In_1710);
nand U2010 (N_2010,In_1876,In_683);
nand U2011 (N_2011,In_607,In_1792);
nand U2012 (N_2012,In_1546,In_32);
nand U2013 (N_2013,In_1524,In_1075);
and U2014 (N_2014,In_1853,In_1891);
or U2015 (N_2015,In_1958,In_1635);
and U2016 (N_2016,In_1206,In_264);
xnor U2017 (N_2017,In_32,In_1583);
nor U2018 (N_2018,In_1535,In_1695);
nor U2019 (N_2019,In_17,In_746);
and U2020 (N_2020,In_897,In_694);
xor U2021 (N_2021,In_1933,In_745);
xor U2022 (N_2022,In_1075,In_1230);
nor U2023 (N_2023,In_1679,In_1592);
nand U2024 (N_2024,In_137,In_363);
and U2025 (N_2025,In_1433,In_626);
or U2026 (N_2026,In_1990,In_1908);
nor U2027 (N_2027,In_1940,In_753);
or U2028 (N_2028,In_1186,In_1108);
nor U2029 (N_2029,In_360,In_268);
xor U2030 (N_2030,In_1545,In_46);
or U2031 (N_2031,In_199,In_1984);
and U2032 (N_2032,In_1569,In_189);
and U2033 (N_2033,In_1322,In_1061);
xor U2034 (N_2034,In_943,In_1494);
nor U2035 (N_2035,In_74,In_683);
nand U2036 (N_2036,In_1062,In_1127);
xnor U2037 (N_2037,In_393,In_988);
and U2038 (N_2038,In_64,In_1231);
and U2039 (N_2039,In_107,In_355);
xor U2040 (N_2040,In_1255,In_1766);
and U2041 (N_2041,In_226,In_1232);
or U2042 (N_2042,In_697,In_873);
or U2043 (N_2043,In_253,In_940);
nand U2044 (N_2044,In_608,In_1593);
and U2045 (N_2045,In_845,In_1507);
nor U2046 (N_2046,In_1974,In_1566);
nor U2047 (N_2047,In_747,In_1686);
and U2048 (N_2048,In_1887,In_857);
xor U2049 (N_2049,In_1019,In_877);
xor U2050 (N_2050,In_999,In_131);
or U2051 (N_2051,In_118,In_1370);
nand U2052 (N_2052,In_602,In_1093);
nor U2053 (N_2053,In_791,In_1362);
or U2054 (N_2054,In_1028,In_457);
or U2055 (N_2055,In_1749,In_1098);
xnor U2056 (N_2056,In_1998,In_1245);
nor U2057 (N_2057,In_1299,In_1451);
nor U2058 (N_2058,In_1773,In_5);
nand U2059 (N_2059,In_1853,In_1031);
nand U2060 (N_2060,In_542,In_1509);
nand U2061 (N_2061,In_1048,In_1288);
and U2062 (N_2062,In_669,In_1658);
nand U2063 (N_2063,In_175,In_1374);
nand U2064 (N_2064,In_680,In_1138);
nand U2065 (N_2065,In_1549,In_1816);
or U2066 (N_2066,In_995,In_294);
nand U2067 (N_2067,In_879,In_1941);
nor U2068 (N_2068,In_691,In_1611);
nand U2069 (N_2069,In_1840,In_96);
xor U2070 (N_2070,In_342,In_1695);
nor U2071 (N_2071,In_1279,In_1233);
and U2072 (N_2072,In_1961,In_894);
and U2073 (N_2073,In_1704,In_565);
nor U2074 (N_2074,In_691,In_1026);
nor U2075 (N_2075,In_1778,In_838);
nor U2076 (N_2076,In_480,In_469);
nand U2077 (N_2077,In_1008,In_1779);
nor U2078 (N_2078,In_219,In_271);
and U2079 (N_2079,In_9,In_1710);
xor U2080 (N_2080,In_245,In_1013);
and U2081 (N_2081,In_470,In_344);
xnor U2082 (N_2082,In_1805,In_1244);
and U2083 (N_2083,In_279,In_351);
nor U2084 (N_2084,In_423,In_1910);
nor U2085 (N_2085,In_733,In_246);
and U2086 (N_2086,In_1094,In_1295);
nor U2087 (N_2087,In_83,In_430);
and U2088 (N_2088,In_1951,In_1387);
nand U2089 (N_2089,In_76,In_207);
xor U2090 (N_2090,In_1463,In_959);
nor U2091 (N_2091,In_912,In_53);
nand U2092 (N_2092,In_1748,In_954);
and U2093 (N_2093,In_1569,In_1856);
and U2094 (N_2094,In_1504,In_279);
or U2095 (N_2095,In_1314,In_1380);
nand U2096 (N_2096,In_402,In_134);
or U2097 (N_2097,In_224,In_1190);
or U2098 (N_2098,In_339,In_52);
and U2099 (N_2099,In_1158,In_1194);
nor U2100 (N_2100,In_1983,In_92);
or U2101 (N_2101,In_482,In_1014);
or U2102 (N_2102,In_920,In_1013);
or U2103 (N_2103,In_307,In_258);
and U2104 (N_2104,In_1698,In_1832);
and U2105 (N_2105,In_658,In_1733);
and U2106 (N_2106,In_688,In_242);
nand U2107 (N_2107,In_1124,In_1671);
nor U2108 (N_2108,In_1892,In_1933);
and U2109 (N_2109,In_1999,In_597);
or U2110 (N_2110,In_1131,In_343);
or U2111 (N_2111,In_1515,In_1714);
or U2112 (N_2112,In_654,In_121);
xnor U2113 (N_2113,In_652,In_1943);
xnor U2114 (N_2114,In_586,In_550);
nand U2115 (N_2115,In_1464,In_240);
or U2116 (N_2116,In_762,In_1187);
xor U2117 (N_2117,In_324,In_1053);
or U2118 (N_2118,In_828,In_1427);
and U2119 (N_2119,In_1387,In_1360);
or U2120 (N_2120,In_508,In_615);
and U2121 (N_2121,In_628,In_1502);
nand U2122 (N_2122,In_436,In_631);
or U2123 (N_2123,In_1741,In_1693);
nor U2124 (N_2124,In_1150,In_285);
and U2125 (N_2125,In_1182,In_754);
and U2126 (N_2126,In_1767,In_678);
or U2127 (N_2127,In_1946,In_1192);
xor U2128 (N_2128,In_704,In_47);
and U2129 (N_2129,In_188,In_654);
nand U2130 (N_2130,In_1617,In_115);
nor U2131 (N_2131,In_185,In_940);
and U2132 (N_2132,In_750,In_1497);
nand U2133 (N_2133,In_571,In_563);
nand U2134 (N_2134,In_314,In_1015);
nand U2135 (N_2135,In_494,In_1074);
and U2136 (N_2136,In_1274,In_253);
nand U2137 (N_2137,In_1161,In_1883);
and U2138 (N_2138,In_1172,In_294);
nand U2139 (N_2139,In_86,In_829);
nand U2140 (N_2140,In_486,In_743);
and U2141 (N_2141,In_1938,In_207);
or U2142 (N_2142,In_803,In_1089);
nand U2143 (N_2143,In_607,In_340);
and U2144 (N_2144,In_1815,In_144);
xor U2145 (N_2145,In_609,In_355);
nand U2146 (N_2146,In_171,In_1265);
nor U2147 (N_2147,In_525,In_176);
xnor U2148 (N_2148,In_1581,In_735);
and U2149 (N_2149,In_649,In_927);
nand U2150 (N_2150,In_1671,In_202);
or U2151 (N_2151,In_731,In_338);
nand U2152 (N_2152,In_1168,In_197);
and U2153 (N_2153,In_196,In_77);
or U2154 (N_2154,In_1681,In_1072);
nor U2155 (N_2155,In_406,In_591);
or U2156 (N_2156,In_1277,In_1638);
nand U2157 (N_2157,In_1694,In_1897);
or U2158 (N_2158,In_24,In_1931);
and U2159 (N_2159,In_1637,In_103);
xnor U2160 (N_2160,In_505,In_371);
nor U2161 (N_2161,In_1401,In_1438);
xnor U2162 (N_2162,In_630,In_115);
xnor U2163 (N_2163,In_1092,In_523);
nor U2164 (N_2164,In_1470,In_1764);
nor U2165 (N_2165,In_904,In_1869);
nor U2166 (N_2166,In_96,In_1359);
nor U2167 (N_2167,In_1653,In_1919);
nand U2168 (N_2168,In_1650,In_1194);
nor U2169 (N_2169,In_378,In_1957);
or U2170 (N_2170,In_1314,In_1924);
or U2171 (N_2171,In_770,In_464);
nand U2172 (N_2172,In_1373,In_1646);
xor U2173 (N_2173,In_1016,In_1462);
nand U2174 (N_2174,In_502,In_1333);
nor U2175 (N_2175,In_253,In_1062);
xor U2176 (N_2176,In_843,In_1508);
nor U2177 (N_2177,In_1542,In_1013);
xnor U2178 (N_2178,In_1321,In_1017);
and U2179 (N_2179,In_927,In_1783);
nor U2180 (N_2180,In_1568,In_211);
nor U2181 (N_2181,In_103,In_1369);
and U2182 (N_2182,In_862,In_674);
and U2183 (N_2183,In_1141,In_249);
nand U2184 (N_2184,In_1419,In_930);
or U2185 (N_2185,In_673,In_1817);
and U2186 (N_2186,In_586,In_539);
nor U2187 (N_2187,In_1512,In_1824);
nor U2188 (N_2188,In_429,In_1768);
xor U2189 (N_2189,In_1629,In_1965);
and U2190 (N_2190,In_797,In_1922);
or U2191 (N_2191,In_1598,In_444);
xnor U2192 (N_2192,In_1161,In_900);
or U2193 (N_2193,In_1899,In_593);
and U2194 (N_2194,In_1208,In_731);
xor U2195 (N_2195,In_507,In_874);
or U2196 (N_2196,In_1911,In_941);
xnor U2197 (N_2197,In_535,In_828);
xnor U2198 (N_2198,In_450,In_834);
nor U2199 (N_2199,In_1620,In_638);
nand U2200 (N_2200,In_677,In_945);
xnor U2201 (N_2201,In_647,In_1664);
nor U2202 (N_2202,In_582,In_975);
nand U2203 (N_2203,In_497,In_961);
nand U2204 (N_2204,In_278,In_1825);
xnor U2205 (N_2205,In_368,In_362);
or U2206 (N_2206,In_1665,In_587);
xnor U2207 (N_2207,In_549,In_1281);
nand U2208 (N_2208,In_936,In_388);
or U2209 (N_2209,In_156,In_1550);
and U2210 (N_2210,In_1577,In_1457);
nor U2211 (N_2211,In_126,In_403);
and U2212 (N_2212,In_1972,In_1140);
or U2213 (N_2213,In_105,In_1600);
nor U2214 (N_2214,In_71,In_655);
xnor U2215 (N_2215,In_1114,In_1593);
nor U2216 (N_2216,In_241,In_303);
and U2217 (N_2217,In_1032,In_352);
nand U2218 (N_2218,In_440,In_1165);
nand U2219 (N_2219,In_951,In_677);
and U2220 (N_2220,In_170,In_1779);
and U2221 (N_2221,In_138,In_877);
and U2222 (N_2222,In_1518,In_1678);
nand U2223 (N_2223,In_992,In_1049);
nand U2224 (N_2224,In_1827,In_992);
or U2225 (N_2225,In_1328,In_1059);
xnor U2226 (N_2226,In_166,In_1721);
or U2227 (N_2227,In_1589,In_1638);
nand U2228 (N_2228,In_70,In_744);
xnor U2229 (N_2229,In_550,In_1053);
or U2230 (N_2230,In_946,In_908);
or U2231 (N_2231,In_1572,In_687);
xor U2232 (N_2232,In_1418,In_1124);
nor U2233 (N_2233,In_1192,In_794);
nand U2234 (N_2234,In_1055,In_213);
nand U2235 (N_2235,In_140,In_1538);
and U2236 (N_2236,In_1286,In_1197);
nand U2237 (N_2237,In_1071,In_1182);
or U2238 (N_2238,In_1653,In_1364);
and U2239 (N_2239,In_1417,In_629);
or U2240 (N_2240,In_585,In_91);
nand U2241 (N_2241,In_1371,In_1099);
xnor U2242 (N_2242,In_763,In_53);
nor U2243 (N_2243,In_489,In_1363);
nand U2244 (N_2244,In_1961,In_1451);
and U2245 (N_2245,In_496,In_243);
nor U2246 (N_2246,In_1912,In_606);
nor U2247 (N_2247,In_56,In_1814);
xor U2248 (N_2248,In_939,In_1086);
and U2249 (N_2249,In_160,In_1799);
or U2250 (N_2250,In_1538,In_808);
xor U2251 (N_2251,In_882,In_1269);
nor U2252 (N_2252,In_107,In_11);
and U2253 (N_2253,In_605,In_1414);
nor U2254 (N_2254,In_1554,In_550);
and U2255 (N_2255,In_1579,In_1766);
xnor U2256 (N_2256,In_1682,In_1138);
nor U2257 (N_2257,In_173,In_1113);
xor U2258 (N_2258,In_1852,In_537);
xor U2259 (N_2259,In_1563,In_1271);
nand U2260 (N_2260,In_258,In_662);
nor U2261 (N_2261,In_618,In_1960);
nor U2262 (N_2262,In_1384,In_1828);
nor U2263 (N_2263,In_1120,In_1798);
nor U2264 (N_2264,In_1335,In_1077);
and U2265 (N_2265,In_608,In_1956);
nor U2266 (N_2266,In_98,In_1506);
nand U2267 (N_2267,In_1602,In_1200);
or U2268 (N_2268,In_1317,In_345);
nor U2269 (N_2269,In_1814,In_144);
nor U2270 (N_2270,In_1737,In_69);
nor U2271 (N_2271,In_239,In_1191);
or U2272 (N_2272,In_1185,In_448);
or U2273 (N_2273,In_1307,In_155);
or U2274 (N_2274,In_1535,In_769);
xnor U2275 (N_2275,In_1298,In_417);
nor U2276 (N_2276,In_1840,In_1887);
nand U2277 (N_2277,In_1930,In_1514);
and U2278 (N_2278,In_1534,In_1781);
nand U2279 (N_2279,In_564,In_1398);
and U2280 (N_2280,In_1668,In_585);
xnor U2281 (N_2281,In_1581,In_348);
or U2282 (N_2282,In_852,In_834);
nor U2283 (N_2283,In_1879,In_1636);
xor U2284 (N_2284,In_1618,In_895);
xor U2285 (N_2285,In_1442,In_242);
xor U2286 (N_2286,In_820,In_936);
nand U2287 (N_2287,In_1596,In_732);
xor U2288 (N_2288,In_1721,In_769);
xnor U2289 (N_2289,In_1903,In_946);
xnor U2290 (N_2290,In_651,In_1765);
nand U2291 (N_2291,In_614,In_1663);
xnor U2292 (N_2292,In_1755,In_844);
and U2293 (N_2293,In_69,In_648);
or U2294 (N_2294,In_1277,In_1881);
or U2295 (N_2295,In_1119,In_509);
xnor U2296 (N_2296,In_343,In_426);
and U2297 (N_2297,In_824,In_1725);
and U2298 (N_2298,In_856,In_1107);
nand U2299 (N_2299,In_302,In_621);
or U2300 (N_2300,In_1603,In_860);
nor U2301 (N_2301,In_1554,In_1111);
xnor U2302 (N_2302,In_664,In_952);
or U2303 (N_2303,In_759,In_1865);
xor U2304 (N_2304,In_460,In_32);
or U2305 (N_2305,In_1509,In_1614);
or U2306 (N_2306,In_196,In_752);
or U2307 (N_2307,In_1339,In_94);
and U2308 (N_2308,In_1681,In_614);
nand U2309 (N_2309,In_1270,In_751);
nand U2310 (N_2310,In_139,In_1269);
nor U2311 (N_2311,In_500,In_255);
nand U2312 (N_2312,In_266,In_1756);
nor U2313 (N_2313,In_1849,In_141);
nand U2314 (N_2314,In_800,In_769);
and U2315 (N_2315,In_1185,In_662);
nor U2316 (N_2316,In_1405,In_429);
xnor U2317 (N_2317,In_1202,In_1941);
or U2318 (N_2318,In_887,In_781);
nand U2319 (N_2319,In_1646,In_1049);
nor U2320 (N_2320,In_385,In_1685);
nor U2321 (N_2321,In_1424,In_708);
nor U2322 (N_2322,In_1913,In_1529);
nand U2323 (N_2323,In_580,In_147);
nor U2324 (N_2324,In_663,In_337);
nand U2325 (N_2325,In_1470,In_1587);
and U2326 (N_2326,In_1571,In_386);
xor U2327 (N_2327,In_1869,In_1378);
and U2328 (N_2328,In_158,In_1990);
or U2329 (N_2329,In_734,In_1984);
nor U2330 (N_2330,In_606,In_755);
xnor U2331 (N_2331,In_728,In_484);
nand U2332 (N_2332,In_1160,In_1352);
and U2333 (N_2333,In_730,In_735);
and U2334 (N_2334,In_455,In_711);
nor U2335 (N_2335,In_1062,In_1084);
and U2336 (N_2336,In_1750,In_1794);
and U2337 (N_2337,In_1392,In_314);
and U2338 (N_2338,In_85,In_1794);
xor U2339 (N_2339,In_250,In_75);
nor U2340 (N_2340,In_353,In_1358);
and U2341 (N_2341,In_1661,In_1113);
or U2342 (N_2342,In_930,In_1057);
xnor U2343 (N_2343,In_1542,In_1830);
nor U2344 (N_2344,In_691,In_654);
nor U2345 (N_2345,In_1987,In_1409);
nand U2346 (N_2346,In_1138,In_502);
and U2347 (N_2347,In_1300,In_577);
nand U2348 (N_2348,In_63,In_1889);
nor U2349 (N_2349,In_1266,In_1643);
nand U2350 (N_2350,In_290,In_84);
nor U2351 (N_2351,In_1330,In_716);
or U2352 (N_2352,In_1753,In_766);
xnor U2353 (N_2353,In_797,In_949);
nor U2354 (N_2354,In_1701,In_1835);
nor U2355 (N_2355,In_1676,In_149);
xor U2356 (N_2356,In_126,In_737);
nor U2357 (N_2357,In_1245,In_1148);
nor U2358 (N_2358,In_1033,In_703);
xor U2359 (N_2359,In_829,In_837);
nand U2360 (N_2360,In_1648,In_1847);
xor U2361 (N_2361,In_1504,In_269);
nand U2362 (N_2362,In_1295,In_1620);
nor U2363 (N_2363,In_1801,In_906);
xor U2364 (N_2364,In_1136,In_418);
and U2365 (N_2365,In_1902,In_863);
nor U2366 (N_2366,In_74,In_492);
nand U2367 (N_2367,In_365,In_1671);
or U2368 (N_2368,In_9,In_1120);
xnor U2369 (N_2369,In_1597,In_356);
nand U2370 (N_2370,In_165,In_889);
and U2371 (N_2371,In_72,In_846);
nand U2372 (N_2372,In_1948,In_781);
xor U2373 (N_2373,In_67,In_647);
nand U2374 (N_2374,In_1920,In_1367);
xnor U2375 (N_2375,In_737,In_305);
or U2376 (N_2376,In_145,In_225);
nor U2377 (N_2377,In_287,In_805);
nor U2378 (N_2378,In_668,In_813);
and U2379 (N_2379,In_613,In_1586);
and U2380 (N_2380,In_833,In_1263);
nand U2381 (N_2381,In_1717,In_690);
xnor U2382 (N_2382,In_1452,In_543);
or U2383 (N_2383,In_1031,In_1164);
or U2384 (N_2384,In_587,In_429);
nand U2385 (N_2385,In_1144,In_1725);
xnor U2386 (N_2386,In_845,In_87);
nor U2387 (N_2387,In_1925,In_1760);
xnor U2388 (N_2388,In_1915,In_1864);
nor U2389 (N_2389,In_1945,In_1902);
or U2390 (N_2390,In_408,In_795);
nor U2391 (N_2391,In_1600,In_690);
or U2392 (N_2392,In_402,In_559);
nor U2393 (N_2393,In_58,In_260);
xnor U2394 (N_2394,In_1532,In_1264);
nor U2395 (N_2395,In_1253,In_1833);
and U2396 (N_2396,In_82,In_1019);
nor U2397 (N_2397,In_525,In_527);
or U2398 (N_2398,In_1700,In_1849);
or U2399 (N_2399,In_113,In_1863);
xnor U2400 (N_2400,In_698,In_1680);
xnor U2401 (N_2401,In_350,In_1447);
nor U2402 (N_2402,In_1831,In_542);
nor U2403 (N_2403,In_1172,In_1676);
or U2404 (N_2404,In_1440,In_428);
or U2405 (N_2405,In_491,In_1296);
and U2406 (N_2406,In_1692,In_290);
and U2407 (N_2407,In_780,In_1101);
nor U2408 (N_2408,In_416,In_1218);
and U2409 (N_2409,In_1530,In_1734);
nor U2410 (N_2410,In_160,In_1467);
and U2411 (N_2411,In_151,In_646);
or U2412 (N_2412,In_1873,In_293);
or U2413 (N_2413,In_1365,In_236);
nor U2414 (N_2414,In_1259,In_555);
and U2415 (N_2415,In_1365,In_1140);
nor U2416 (N_2416,In_872,In_1778);
nor U2417 (N_2417,In_1765,In_984);
nand U2418 (N_2418,In_1690,In_1483);
xnor U2419 (N_2419,In_1352,In_823);
xor U2420 (N_2420,In_222,In_1112);
nand U2421 (N_2421,In_555,In_921);
nand U2422 (N_2422,In_403,In_947);
or U2423 (N_2423,In_1739,In_1425);
nor U2424 (N_2424,In_442,In_696);
or U2425 (N_2425,In_125,In_517);
or U2426 (N_2426,In_1478,In_560);
xnor U2427 (N_2427,In_231,In_1904);
nand U2428 (N_2428,In_1232,In_1911);
nor U2429 (N_2429,In_289,In_603);
and U2430 (N_2430,In_1519,In_1293);
xor U2431 (N_2431,In_1330,In_1779);
and U2432 (N_2432,In_1851,In_1783);
nor U2433 (N_2433,In_1135,In_1853);
or U2434 (N_2434,In_1918,In_236);
nand U2435 (N_2435,In_543,In_1148);
xnor U2436 (N_2436,In_1841,In_420);
nand U2437 (N_2437,In_1230,In_921);
xnor U2438 (N_2438,In_1170,In_320);
nor U2439 (N_2439,In_468,In_1747);
or U2440 (N_2440,In_1708,In_1456);
xor U2441 (N_2441,In_164,In_1939);
or U2442 (N_2442,In_884,In_1347);
nand U2443 (N_2443,In_85,In_587);
and U2444 (N_2444,In_1102,In_628);
nand U2445 (N_2445,In_445,In_377);
or U2446 (N_2446,In_120,In_522);
and U2447 (N_2447,In_1798,In_982);
or U2448 (N_2448,In_943,In_1591);
nor U2449 (N_2449,In_1682,In_1739);
nand U2450 (N_2450,In_1994,In_1785);
nor U2451 (N_2451,In_1154,In_1893);
nor U2452 (N_2452,In_369,In_1200);
nand U2453 (N_2453,In_1128,In_1982);
nor U2454 (N_2454,In_687,In_1402);
or U2455 (N_2455,In_826,In_1595);
or U2456 (N_2456,In_932,In_278);
or U2457 (N_2457,In_1321,In_138);
nor U2458 (N_2458,In_899,In_627);
xnor U2459 (N_2459,In_1642,In_1967);
xnor U2460 (N_2460,In_885,In_490);
and U2461 (N_2461,In_330,In_871);
nand U2462 (N_2462,In_871,In_307);
nand U2463 (N_2463,In_152,In_1552);
or U2464 (N_2464,In_230,In_376);
and U2465 (N_2465,In_1069,In_642);
or U2466 (N_2466,In_1260,In_627);
nand U2467 (N_2467,In_1488,In_36);
nand U2468 (N_2468,In_1643,In_1816);
nor U2469 (N_2469,In_1300,In_1428);
xor U2470 (N_2470,In_881,In_1038);
and U2471 (N_2471,In_602,In_603);
or U2472 (N_2472,In_833,In_1855);
and U2473 (N_2473,In_1833,In_1226);
or U2474 (N_2474,In_1546,In_64);
nor U2475 (N_2475,In_1514,In_1752);
xor U2476 (N_2476,In_1935,In_821);
nand U2477 (N_2477,In_1134,In_1443);
nand U2478 (N_2478,In_853,In_571);
nor U2479 (N_2479,In_378,In_1190);
nor U2480 (N_2480,In_103,In_262);
xnor U2481 (N_2481,In_469,In_355);
xnor U2482 (N_2482,In_1092,In_1017);
nor U2483 (N_2483,In_1697,In_680);
nor U2484 (N_2484,In_1249,In_1823);
nand U2485 (N_2485,In_1823,In_1427);
or U2486 (N_2486,In_295,In_1485);
xnor U2487 (N_2487,In_1098,In_1291);
or U2488 (N_2488,In_244,In_33);
xnor U2489 (N_2489,In_1717,In_813);
xnor U2490 (N_2490,In_709,In_901);
or U2491 (N_2491,In_145,In_685);
and U2492 (N_2492,In_1291,In_920);
and U2493 (N_2493,In_1683,In_382);
and U2494 (N_2494,In_980,In_1905);
xnor U2495 (N_2495,In_1106,In_1649);
or U2496 (N_2496,In_362,In_168);
nor U2497 (N_2497,In_166,In_962);
xor U2498 (N_2498,In_215,In_1084);
nor U2499 (N_2499,In_1067,In_1949);
and U2500 (N_2500,In_788,In_1196);
nand U2501 (N_2501,In_1059,In_534);
or U2502 (N_2502,In_643,In_1890);
or U2503 (N_2503,In_504,In_1332);
nor U2504 (N_2504,In_1198,In_1283);
nand U2505 (N_2505,In_1168,In_1600);
and U2506 (N_2506,In_523,In_433);
xnor U2507 (N_2507,In_944,In_1816);
and U2508 (N_2508,In_1489,In_1047);
and U2509 (N_2509,In_378,In_1609);
xor U2510 (N_2510,In_909,In_187);
xor U2511 (N_2511,In_457,In_1227);
nand U2512 (N_2512,In_1602,In_356);
nand U2513 (N_2513,In_1251,In_1186);
xor U2514 (N_2514,In_879,In_1072);
nand U2515 (N_2515,In_552,In_1407);
or U2516 (N_2516,In_1273,In_1747);
xnor U2517 (N_2517,In_295,In_1889);
xor U2518 (N_2518,In_1515,In_14);
and U2519 (N_2519,In_805,In_466);
and U2520 (N_2520,In_176,In_1959);
nand U2521 (N_2521,In_1228,In_1159);
or U2522 (N_2522,In_263,In_503);
or U2523 (N_2523,In_1407,In_564);
and U2524 (N_2524,In_417,In_1221);
nand U2525 (N_2525,In_1774,In_1298);
xnor U2526 (N_2526,In_588,In_1050);
xor U2527 (N_2527,In_887,In_1620);
xnor U2528 (N_2528,In_1441,In_700);
nor U2529 (N_2529,In_406,In_350);
or U2530 (N_2530,In_1152,In_1473);
xor U2531 (N_2531,In_1699,In_1549);
nor U2532 (N_2532,In_1220,In_487);
nor U2533 (N_2533,In_451,In_846);
nor U2534 (N_2534,In_722,In_1071);
and U2535 (N_2535,In_963,In_710);
nor U2536 (N_2536,In_55,In_768);
nand U2537 (N_2537,In_454,In_352);
or U2538 (N_2538,In_191,In_1619);
xnor U2539 (N_2539,In_596,In_798);
nand U2540 (N_2540,In_165,In_1254);
xnor U2541 (N_2541,In_1888,In_1158);
nand U2542 (N_2542,In_1071,In_973);
nor U2543 (N_2543,In_1365,In_98);
xnor U2544 (N_2544,In_147,In_432);
nand U2545 (N_2545,In_1463,In_1319);
nor U2546 (N_2546,In_1248,In_427);
nor U2547 (N_2547,In_1552,In_1679);
or U2548 (N_2548,In_1965,In_757);
nor U2549 (N_2549,In_695,In_1599);
or U2550 (N_2550,In_423,In_1486);
or U2551 (N_2551,In_563,In_1827);
nor U2552 (N_2552,In_1022,In_1482);
or U2553 (N_2553,In_1693,In_609);
or U2554 (N_2554,In_1413,In_1477);
nor U2555 (N_2555,In_271,In_365);
xnor U2556 (N_2556,In_177,In_1571);
nor U2557 (N_2557,In_1716,In_1879);
xor U2558 (N_2558,In_50,In_43);
or U2559 (N_2559,In_1286,In_1458);
nor U2560 (N_2560,In_1072,In_1844);
nand U2561 (N_2561,In_1267,In_973);
nand U2562 (N_2562,In_782,In_709);
nand U2563 (N_2563,In_75,In_381);
nor U2564 (N_2564,In_1219,In_1163);
xor U2565 (N_2565,In_791,In_294);
nor U2566 (N_2566,In_163,In_1636);
and U2567 (N_2567,In_566,In_748);
xor U2568 (N_2568,In_1142,In_1179);
and U2569 (N_2569,In_851,In_1065);
or U2570 (N_2570,In_1191,In_1059);
and U2571 (N_2571,In_491,In_1277);
or U2572 (N_2572,In_976,In_714);
nand U2573 (N_2573,In_130,In_1748);
and U2574 (N_2574,In_1542,In_1026);
and U2575 (N_2575,In_1696,In_197);
or U2576 (N_2576,In_1325,In_279);
nor U2577 (N_2577,In_801,In_1158);
nand U2578 (N_2578,In_50,In_1389);
nand U2579 (N_2579,In_377,In_1060);
and U2580 (N_2580,In_973,In_1505);
xor U2581 (N_2581,In_1583,In_249);
and U2582 (N_2582,In_1820,In_1326);
or U2583 (N_2583,In_231,In_328);
nand U2584 (N_2584,In_1713,In_247);
nor U2585 (N_2585,In_1179,In_584);
xnor U2586 (N_2586,In_236,In_998);
nor U2587 (N_2587,In_1744,In_196);
or U2588 (N_2588,In_1019,In_76);
or U2589 (N_2589,In_1974,In_774);
nor U2590 (N_2590,In_376,In_1995);
or U2591 (N_2591,In_729,In_1836);
and U2592 (N_2592,In_486,In_76);
or U2593 (N_2593,In_1512,In_452);
or U2594 (N_2594,In_1326,In_1480);
nand U2595 (N_2595,In_1430,In_1677);
or U2596 (N_2596,In_1603,In_685);
or U2597 (N_2597,In_1306,In_728);
or U2598 (N_2598,In_1156,In_1166);
xor U2599 (N_2599,In_926,In_888);
nor U2600 (N_2600,In_1031,In_557);
nand U2601 (N_2601,In_67,In_1595);
or U2602 (N_2602,In_1783,In_1633);
and U2603 (N_2603,In_152,In_492);
and U2604 (N_2604,In_1998,In_504);
nor U2605 (N_2605,In_1528,In_569);
and U2606 (N_2606,In_1070,In_1662);
nand U2607 (N_2607,In_1790,In_1140);
or U2608 (N_2608,In_1312,In_52);
nand U2609 (N_2609,In_1536,In_1596);
and U2610 (N_2610,In_1535,In_341);
nand U2611 (N_2611,In_1058,In_1038);
nor U2612 (N_2612,In_711,In_1732);
or U2613 (N_2613,In_1255,In_504);
or U2614 (N_2614,In_1976,In_1248);
xor U2615 (N_2615,In_1953,In_1165);
and U2616 (N_2616,In_1779,In_202);
and U2617 (N_2617,In_1706,In_1106);
xor U2618 (N_2618,In_1940,In_265);
nand U2619 (N_2619,In_1676,In_26);
xor U2620 (N_2620,In_1358,In_87);
nand U2621 (N_2621,In_1181,In_1279);
xnor U2622 (N_2622,In_1739,In_434);
or U2623 (N_2623,In_1672,In_331);
or U2624 (N_2624,In_1646,In_1103);
nand U2625 (N_2625,In_1173,In_1607);
and U2626 (N_2626,In_160,In_1267);
and U2627 (N_2627,In_1611,In_416);
nand U2628 (N_2628,In_1013,In_371);
nor U2629 (N_2629,In_1758,In_1502);
or U2630 (N_2630,In_1764,In_805);
nor U2631 (N_2631,In_1416,In_1823);
nand U2632 (N_2632,In_1391,In_505);
and U2633 (N_2633,In_1518,In_881);
and U2634 (N_2634,In_213,In_1288);
xor U2635 (N_2635,In_892,In_616);
nor U2636 (N_2636,In_1099,In_80);
and U2637 (N_2637,In_131,In_1900);
xnor U2638 (N_2638,In_1137,In_1080);
and U2639 (N_2639,In_307,In_1746);
nor U2640 (N_2640,In_713,In_1325);
and U2641 (N_2641,In_773,In_585);
or U2642 (N_2642,In_1490,In_1901);
nand U2643 (N_2643,In_669,In_226);
and U2644 (N_2644,In_140,In_922);
nand U2645 (N_2645,In_1598,In_1178);
or U2646 (N_2646,In_1718,In_497);
nor U2647 (N_2647,In_421,In_1437);
xor U2648 (N_2648,In_926,In_913);
xnor U2649 (N_2649,In_1831,In_332);
xnor U2650 (N_2650,In_836,In_279);
or U2651 (N_2651,In_1029,In_1152);
xor U2652 (N_2652,In_64,In_1129);
nand U2653 (N_2653,In_747,In_31);
nor U2654 (N_2654,In_980,In_1411);
nand U2655 (N_2655,In_1320,In_277);
or U2656 (N_2656,In_874,In_404);
nand U2657 (N_2657,In_927,In_249);
or U2658 (N_2658,In_868,In_949);
or U2659 (N_2659,In_993,In_1562);
nand U2660 (N_2660,In_1648,In_1345);
xor U2661 (N_2661,In_817,In_821);
and U2662 (N_2662,In_588,In_401);
and U2663 (N_2663,In_1446,In_720);
nand U2664 (N_2664,In_1215,In_541);
nand U2665 (N_2665,In_730,In_447);
and U2666 (N_2666,In_1701,In_708);
and U2667 (N_2667,In_1922,In_165);
and U2668 (N_2668,In_1059,In_1594);
nor U2669 (N_2669,In_1971,In_942);
or U2670 (N_2670,In_931,In_420);
and U2671 (N_2671,In_970,In_1063);
or U2672 (N_2672,In_92,In_1437);
or U2673 (N_2673,In_592,In_1165);
nor U2674 (N_2674,In_448,In_264);
xnor U2675 (N_2675,In_1435,In_1716);
xnor U2676 (N_2676,In_1026,In_711);
or U2677 (N_2677,In_1221,In_1021);
or U2678 (N_2678,In_407,In_1727);
or U2679 (N_2679,In_1842,In_1152);
nor U2680 (N_2680,In_1213,In_1115);
or U2681 (N_2681,In_425,In_1355);
or U2682 (N_2682,In_867,In_601);
nand U2683 (N_2683,In_27,In_517);
or U2684 (N_2684,In_788,In_914);
xor U2685 (N_2685,In_564,In_226);
or U2686 (N_2686,In_1866,In_1943);
or U2687 (N_2687,In_360,In_1054);
xor U2688 (N_2688,In_1958,In_1241);
xnor U2689 (N_2689,In_101,In_155);
nand U2690 (N_2690,In_1160,In_982);
xor U2691 (N_2691,In_1613,In_558);
nand U2692 (N_2692,In_863,In_1678);
xor U2693 (N_2693,In_600,In_277);
and U2694 (N_2694,In_1160,In_853);
nor U2695 (N_2695,In_557,In_1405);
nand U2696 (N_2696,In_1165,In_1860);
or U2697 (N_2697,In_1496,In_1898);
xnor U2698 (N_2698,In_1603,In_283);
or U2699 (N_2699,In_1256,In_890);
nor U2700 (N_2700,In_216,In_1566);
and U2701 (N_2701,In_314,In_1910);
xor U2702 (N_2702,In_1695,In_252);
nand U2703 (N_2703,In_751,In_1479);
nand U2704 (N_2704,In_222,In_218);
xnor U2705 (N_2705,In_177,In_134);
or U2706 (N_2706,In_1032,In_1296);
nand U2707 (N_2707,In_610,In_1162);
nand U2708 (N_2708,In_638,In_712);
nor U2709 (N_2709,In_1195,In_384);
nand U2710 (N_2710,In_366,In_1519);
or U2711 (N_2711,In_1675,In_1525);
xor U2712 (N_2712,In_1476,In_469);
nand U2713 (N_2713,In_121,In_1908);
or U2714 (N_2714,In_990,In_517);
and U2715 (N_2715,In_1413,In_1165);
and U2716 (N_2716,In_1605,In_1279);
nor U2717 (N_2717,In_1583,In_1372);
and U2718 (N_2718,In_1041,In_1341);
or U2719 (N_2719,In_1693,In_1384);
or U2720 (N_2720,In_662,In_1917);
and U2721 (N_2721,In_302,In_525);
nand U2722 (N_2722,In_1654,In_1305);
and U2723 (N_2723,In_984,In_699);
or U2724 (N_2724,In_980,In_693);
and U2725 (N_2725,In_743,In_1363);
or U2726 (N_2726,In_1604,In_1668);
xnor U2727 (N_2727,In_1181,In_1192);
nor U2728 (N_2728,In_502,In_1778);
xnor U2729 (N_2729,In_1657,In_547);
xnor U2730 (N_2730,In_283,In_1762);
or U2731 (N_2731,In_1627,In_363);
nor U2732 (N_2732,In_469,In_539);
or U2733 (N_2733,In_1991,In_902);
or U2734 (N_2734,In_1094,In_884);
nor U2735 (N_2735,In_988,In_1271);
or U2736 (N_2736,In_283,In_1360);
and U2737 (N_2737,In_1015,In_1211);
xnor U2738 (N_2738,In_271,In_1022);
or U2739 (N_2739,In_471,In_1988);
or U2740 (N_2740,In_1869,In_1890);
nand U2741 (N_2741,In_1539,In_564);
nand U2742 (N_2742,In_16,In_1041);
or U2743 (N_2743,In_865,In_738);
and U2744 (N_2744,In_199,In_1122);
nor U2745 (N_2745,In_31,In_245);
nand U2746 (N_2746,In_1819,In_1630);
nand U2747 (N_2747,In_1889,In_347);
or U2748 (N_2748,In_815,In_1712);
or U2749 (N_2749,In_1903,In_1450);
and U2750 (N_2750,In_1726,In_1396);
and U2751 (N_2751,In_1423,In_1530);
and U2752 (N_2752,In_818,In_1088);
nand U2753 (N_2753,In_1619,In_50);
xor U2754 (N_2754,In_1998,In_909);
xor U2755 (N_2755,In_814,In_1814);
nand U2756 (N_2756,In_137,In_709);
and U2757 (N_2757,In_1961,In_1708);
nor U2758 (N_2758,In_1390,In_1456);
nand U2759 (N_2759,In_1804,In_302);
xnor U2760 (N_2760,In_1692,In_1732);
nor U2761 (N_2761,In_1312,In_1471);
and U2762 (N_2762,In_153,In_1289);
or U2763 (N_2763,In_1116,In_1589);
and U2764 (N_2764,In_388,In_1916);
or U2765 (N_2765,In_900,In_1166);
or U2766 (N_2766,In_1050,In_1398);
or U2767 (N_2767,In_50,In_1196);
or U2768 (N_2768,In_456,In_1477);
nand U2769 (N_2769,In_121,In_683);
or U2770 (N_2770,In_679,In_1208);
nor U2771 (N_2771,In_1054,In_1834);
or U2772 (N_2772,In_857,In_724);
xor U2773 (N_2773,In_944,In_539);
nand U2774 (N_2774,In_261,In_1038);
and U2775 (N_2775,In_1568,In_243);
or U2776 (N_2776,In_770,In_401);
and U2777 (N_2777,In_1749,In_949);
or U2778 (N_2778,In_21,In_549);
nor U2779 (N_2779,In_1931,In_762);
nand U2780 (N_2780,In_374,In_269);
and U2781 (N_2781,In_898,In_1585);
nand U2782 (N_2782,In_1192,In_1452);
and U2783 (N_2783,In_929,In_177);
or U2784 (N_2784,In_1261,In_754);
and U2785 (N_2785,In_487,In_465);
and U2786 (N_2786,In_1463,In_1899);
xor U2787 (N_2787,In_678,In_895);
nand U2788 (N_2788,In_1582,In_1796);
and U2789 (N_2789,In_628,In_785);
nor U2790 (N_2790,In_48,In_457);
or U2791 (N_2791,In_258,In_1835);
xnor U2792 (N_2792,In_1242,In_518);
nand U2793 (N_2793,In_1669,In_1624);
or U2794 (N_2794,In_594,In_1825);
and U2795 (N_2795,In_732,In_170);
xor U2796 (N_2796,In_1383,In_944);
nor U2797 (N_2797,In_1405,In_278);
or U2798 (N_2798,In_1413,In_468);
and U2799 (N_2799,In_1357,In_1964);
xnor U2800 (N_2800,In_1002,In_1022);
nand U2801 (N_2801,In_1066,In_1050);
and U2802 (N_2802,In_856,In_1611);
xor U2803 (N_2803,In_802,In_1197);
nand U2804 (N_2804,In_650,In_1650);
or U2805 (N_2805,In_1849,In_151);
nand U2806 (N_2806,In_1527,In_877);
xnor U2807 (N_2807,In_586,In_1021);
nor U2808 (N_2808,In_1535,In_1419);
and U2809 (N_2809,In_238,In_318);
nand U2810 (N_2810,In_492,In_872);
xor U2811 (N_2811,In_831,In_1);
and U2812 (N_2812,In_1594,In_1238);
nand U2813 (N_2813,In_1203,In_1540);
nand U2814 (N_2814,In_677,In_248);
or U2815 (N_2815,In_64,In_762);
nand U2816 (N_2816,In_1495,In_209);
or U2817 (N_2817,In_985,In_1727);
xnor U2818 (N_2818,In_363,In_1968);
xor U2819 (N_2819,In_313,In_1411);
nand U2820 (N_2820,In_1005,In_88);
and U2821 (N_2821,In_1056,In_1962);
nand U2822 (N_2822,In_1090,In_895);
nand U2823 (N_2823,In_735,In_483);
nor U2824 (N_2824,In_1857,In_726);
nor U2825 (N_2825,In_352,In_293);
or U2826 (N_2826,In_386,In_792);
nor U2827 (N_2827,In_18,In_1314);
or U2828 (N_2828,In_340,In_1654);
nor U2829 (N_2829,In_1840,In_27);
xor U2830 (N_2830,In_482,In_1275);
and U2831 (N_2831,In_1408,In_706);
nand U2832 (N_2832,In_770,In_311);
nand U2833 (N_2833,In_1427,In_1369);
nor U2834 (N_2834,In_293,In_910);
xnor U2835 (N_2835,In_729,In_713);
and U2836 (N_2836,In_628,In_267);
xnor U2837 (N_2837,In_1011,In_459);
and U2838 (N_2838,In_834,In_1629);
and U2839 (N_2839,In_257,In_1636);
and U2840 (N_2840,In_1801,In_970);
nand U2841 (N_2841,In_1194,In_1464);
or U2842 (N_2842,In_1350,In_1787);
and U2843 (N_2843,In_668,In_1239);
and U2844 (N_2844,In_1894,In_1824);
nand U2845 (N_2845,In_59,In_360);
or U2846 (N_2846,In_1824,In_150);
or U2847 (N_2847,In_62,In_578);
nor U2848 (N_2848,In_1084,In_1995);
nand U2849 (N_2849,In_644,In_1648);
xor U2850 (N_2850,In_1737,In_473);
nand U2851 (N_2851,In_1034,In_811);
nand U2852 (N_2852,In_1144,In_1918);
and U2853 (N_2853,In_1170,In_391);
or U2854 (N_2854,In_1366,In_1655);
xor U2855 (N_2855,In_1326,In_745);
and U2856 (N_2856,In_1594,In_623);
and U2857 (N_2857,In_1941,In_1126);
xor U2858 (N_2858,In_949,In_1834);
nor U2859 (N_2859,In_1336,In_1148);
and U2860 (N_2860,In_394,In_1212);
and U2861 (N_2861,In_555,In_1382);
nor U2862 (N_2862,In_1097,In_254);
xor U2863 (N_2863,In_847,In_677);
nand U2864 (N_2864,In_937,In_1947);
nor U2865 (N_2865,In_699,In_1286);
xor U2866 (N_2866,In_1708,In_49);
nor U2867 (N_2867,In_837,In_106);
nor U2868 (N_2868,In_754,In_427);
and U2869 (N_2869,In_975,In_1418);
xnor U2870 (N_2870,In_648,In_476);
or U2871 (N_2871,In_168,In_1237);
nand U2872 (N_2872,In_174,In_1805);
and U2873 (N_2873,In_738,In_40);
nand U2874 (N_2874,In_1634,In_1034);
xnor U2875 (N_2875,In_257,In_74);
and U2876 (N_2876,In_44,In_611);
or U2877 (N_2877,In_1280,In_1550);
or U2878 (N_2878,In_1871,In_1501);
xnor U2879 (N_2879,In_1760,In_1424);
nand U2880 (N_2880,In_98,In_280);
or U2881 (N_2881,In_1591,In_1205);
nor U2882 (N_2882,In_1573,In_723);
nand U2883 (N_2883,In_1110,In_681);
xor U2884 (N_2884,In_918,In_1553);
nor U2885 (N_2885,In_914,In_1271);
xnor U2886 (N_2886,In_654,In_1186);
nor U2887 (N_2887,In_1627,In_195);
nor U2888 (N_2888,In_1065,In_381);
xor U2889 (N_2889,In_1916,In_1120);
xor U2890 (N_2890,In_925,In_1470);
nand U2891 (N_2891,In_1661,In_840);
and U2892 (N_2892,In_46,In_274);
or U2893 (N_2893,In_1455,In_8);
xnor U2894 (N_2894,In_1183,In_1167);
or U2895 (N_2895,In_434,In_709);
xor U2896 (N_2896,In_1712,In_1031);
or U2897 (N_2897,In_1721,In_931);
nand U2898 (N_2898,In_1460,In_1139);
xnor U2899 (N_2899,In_1322,In_768);
xnor U2900 (N_2900,In_248,In_406);
and U2901 (N_2901,In_747,In_1118);
xor U2902 (N_2902,In_461,In_1264);
and U2903 (N_2903,In_1154,In_1614);
xor U2904 (N_2904,In_1864,In_1867);
nand U2905 (N_2905,In_729,In_918);
xnor U2906 (N_2906,In_1303,In_806);
or U2907 (N_2907,In_1586,In_597);
or U2908 (N_2908,In_475,In_185);
or U2909 (N_2909,In_409,In_910);
xnor U2910 (N_2910,In_231,In_1258);
or U2911 (N_2911,In_1719,In_963);
xnor U2912 (N_2912,In_662,In_87);
and U2913 (N_2913,In_1530,In_1858);
xor U2914 (N_2914,In_818,In_1590);
nor U2915 (N_2915,In_1632,In_1151);
or U2916 (N_2916,In_1904,In_677);
or U2917 (N_2917,In_1975,In_1017);
and U2918 (N_2918,In_292,In_293);
and U2919 (N_2919,In_646,In_751);
or U2920 (N_2920,In_1064,In_5);
nor U2921 (N_2921,In_1266,In_1320);
nor U2922 (N_2922,In_168,In_1235);
nor U2923 (N_2923,In_1346,In_381);
and U2924 (N_2924,In_253,In_1980);
xnor U2925 (N_2925,In_233,In_901);
nor U2926 (N_2926,In_1020,In_1745);
and U2927 (N_2927,In_714,In_1078);
nand U2928 (N_2928,In_889,In_1332);
or U2929 (N_2929,In_1026,In_618);
xor U2930 (N_2930,In_1009,In_120);
nor U2931 (N_2931,In_1072,In_1791);
nor U2932 (N_2932,In_1630,In_484);
or U2933 (N_2933,In_416,In_1093);
or U2934 (N_2934,In_1768,In_801);
nor U2935 (N_2935,In_709,In_842);
or U2936 (N_2936,In_347,In_357);
nor U2937 (N_2937,In_1389,In_1558);
and U2938 (N_2938,In_1677,In_1201);
xnor U2939 (N_2939,In_1924,In_1202);
or U2940 (N_2940,In_1085,In_1612);
nand U2941 (N_2941,In_474,In_1606);
xnor U2942 (N_2942,In_1952,In_770);
nor U2943 (N_2943,In_95,In_496);
or U2944 (N_2944,In_315,In_19);
and U2945 (N_2945,In_1933,In_1483);
or U2946 (N_2946,In_162,In_82);
nor U2947 (N_2947,In_532,In_1889);
nand U2948 (N_2948,In_1433,In_139);
nor U2949 (N_2949,In_1451,In_663);
nand U2950 (N_2950,In_1281,In_1495);
nand U2951 (N_2951,In_347,In_1901);
or U2952 (N_2952,In_716,In_114);
xnor U2953 (N_2953,In_1130,In_1355);
or U2954 (N_2954,In_897,In_1721);
or U2955 (N_2955,In_1636,In_1307);
nand U2956 (N_2956,In_1245,In_402);
or U2957 (N_2957,In_1286,In_1727);
nor U2958 (N_2958,In_863,In_1730);
xnor U2959 (N_2959,In_68,In_1501);
nand U2960 (N_2960,In_878,In_651);
nor U2961 (N_2961,In_989,In_1843);
and U2962 (N_2962,In_1750,In_1128);
and U2963 (N_2963,In_991,In_499);
xor U2964 (N_2964,In_1223,In_918);
nand U2965 (N_2965,In_1749,In_1998);
xnor U2966 (N_2966,In_497,In_570);
nor U2967 (N_2967,In_1316,In_811);
or U2968 (N_2968,In_1416,In_1425);
nor U2969 (N_2969,In_1799,In_1930);
nor U2970 (N_2970,In_158,In_1631);
xor U2971 (N_2971,In_393,In_1116);
and U2972 (N_2972,In_19,In_816);
nand U2973 (N_2973,In_317,In_226);
nand U2974 (N_2974,In_1323,In_155);
nor U2975 (N_2975,In_1641,In_1583);
xor U2976 (N_2976,In_133,In_1009);
xnor U2977 (N_2977,In_1295,In_1506);
nand U2978 (N_2978,In_1411,In_1432);
xor U2979 (N_2979,In_620,In_1738);
nor U2980 (N_2980,In_118,In_1154);
and U2981 (N_2981,In_1275,In_3);
nor U2982 (N_2982,In_906,In_969);
nor U2983 (N_2983,In_1279,In_1032);
and U2984 (N_2984,In_1611,In_789);
or U2985 (N_2985,In_709,In_1946);
nand U2986 (N_2986,In_641,In_1503);
xnor U2987 (N_2987,In_476,In_1011);
nor U2988 (N_2988,In_1710,In_825);
nand U2989 (N_2989,In_495,In_1546);
and U2990 (N_2990,In_1943,In_1650);
or U2991 (N_2991,In_279,In_292);
and U2992 (N_2992,In_350,In_793);
nor U2993 (N_2993,In_482,In_1545);
nand U2994 (N_2994,In_1543,In_594);
xnor U2995 (N_2995,In_1143,In_891);
or U2996 (N_2996,In_640,In_1138);
nand U2997 (N_2997,In_407,In_732);
and U2998 (N_2998,In_1971,In_648);
and U2999 (N_2999,In_1313,In_935);
nand U3000 (N_3000,In_573,In_36);
and U3001 (N_3001,In_1699,In_1010);
nor U3002 (N_3002,In_1084,In_1263);
nor U3003 (N_3003,In_327,In_1666);
nor U3004 (N_3004,In_1271,In_515);
and U3005 (N_3005,In_403,In_1949);
or U3006 (N_3006,In_431,In_1038);
xnor U3007 (N_3007,In_635,In_1978);
or U3008 (N_3008,In_319,In_136);
nand U3009 (N_3009,In_171,In_899);
and U3010 (N_3010,In_1860,In_1582);
and U3011 (N_3011,In_236,In_1284);
xor U3012 (N_3012,In_1641,In_1180);
and U3013 (N_3013,In_830,In_1591);
or U3014 (N_3014,In_1695,In_1573);
xor U3015 (N_3015,In_1847,In_1751);
nor U3016 (N_3016,In_1983,In_1303);
xnor U3017 (N_3017,In_1936,In_197);
nor U3018 (N_3018,In_405,In_1503);
and U3019 (N_3019,In_1097,In_779);
or U3020 (N_3020,In_1853,In_1181);
or U3021 (N_3021,In_1014,In_381);
and U3022 (N_3022,In_715,In_1497);
nor U3023 (N_3023,In_1368,In_1545);
xnor U3024 (N_3024,In_386,In_1919);
nor U3025 (N_3025,In_1299,In_114);
and U3026 (N_3026,In_585,In_1020);
xnor U3027 (N_3027,In_89,In_1663);
and U3028 (N_3028,In_1755,In_1936);
nand U3029 (N_3029,In_492,In_311);
or U3030 (N_3030,In_343,In_521);
nand U3031 (N_3031,In_97,In_652);
nand U3032 (N_3032,In_1589,In_44);
and U3033 (N_3033,In_449,In_590);
nand U3034 (N_3034,In_704,In_1372);
and U3035 (N_3035,In_868,In_666);
or U3036 (N_3036,In_1600,In_529);
or U3037 (N_3037,In_1464,In_936);
nor U3038 (N_3038,In_457,In_476);
or U3039 (N_3039,In_508,In_413);
or U3040 (N_3040,In_444,In_288);
nor U3041 (N_3041,In_932,In_405);
or U3042 (N_3042,In_1876,In_1830);
or U3043 (N_3043,In_581,In_225);
xnor U3044 (N_3044,In_789,In_1472);
xor U3045 (N_3045,In_1001,In_1194);
nor U3046 (N_3046,In_1789,In_1483);
or U3047 (N_3047,In_1483,In_1541);
nor U3048 (N_3048,In_1731,In_47);
and U3049 (N_3049,In_318,In_1826);
and U3050 (N_3050,In_737,In_568);
xnor U3051 (N_3051,In_1216,In_133);
nand U3052 (N_3052,In_929,In_1340);
nand U3053 (N_3053,In_1565,In_1909);
xor U3054 (N_3054,In_995,In_1352);
and U3055 (N_3055,In_160,In_26);
and U3056 (N_3056,In_585,In_1032);
or U3057 (N_3057,In_1307,In_774);
and U3058 (N_3058,In_832,In_1274);
or U3059 (N_3059,In_1918,In_1582);
xor U3060 (N_3060,In_71,In_1272);
or U3061 (N_3061,In_290,In_1490);
and U3062 (N_3062,In_1353,In_1842);
nor U3063 (N_3063,In_1245,In_912);
and U3064 (N_3064,In_393,In_257);
nor U3065 (N_3065,In_1115,In_814);
nor U3066 (N_3066,In_1160,In_1360);
and U3067 (N_3067,In_1435,In_1268);
or U3068 (N_3068,In_1479,In_1369);
nor U3069 (N_3069,In_949,In_1030);
and U3070 (N_3070,In_1052,In_1378);
xnor U3071 (N_3071,In_760,In_1141);
and U3072 (N_3072,In_1800,In_1378);
nor U3073 (N_3073,In_1754,In_1382);
and U3074 (N_3074,In_1792,In_817);
nor U3075 (N_3075,In_1720,In_1977);
xor U3076 (N_3076,In_282,In_135);
and U3077 (N_3077,In_168,In_1600);
nand U3078 (N_3078,In_1096,In_163);
nor U3079 (N_3079,In_1822,In_756);
nor U3080 (N_3080,In_1247,In_91);
and U3081 (N_3081,In_1801,In_1752);
xnor U3082 (N_3082,In_1362,In_126);
nand U3083 (N_3083,In_1708,In_1022);
or U3084 (N_3084,In_1392,In_1918);
xnor U3085 (N_3085,In_1720,In_508);
nor U3086 (N_3086,In_1722,In_387);
or U3087 (N_3087,In_1021,In_1261);
nand U3088 (N_3088,In_80,In_353);
and U3089 (N_3089,In_1277,In_1255);
xor U3090 (N_3090,In_1017,In_1263);
or U3091 (N_3091,In_229,In_65);
xor U3092 (N_3092,In_1815,In_1984);
nand U3093 (N_3093,In_1243,In_1280);
and U3094 (N_3094,In_3,In_395);
and U3095 (N_3095,In_564,In_1309);
or U3096 (N_3096,In_341,In_513);
xnor U3097 (N_3097,In_89,In_706);
and U3098 (N_3098,In_1634,In_1990);
xnor U3099 (N_3099,In_455,In_11);
or U3100 (N_3100,In_1654,In_94);
nor U3101 (N_3101,In_1953,In_218);
nand U3102 (N_3102,In_710,In_416);
or U3103 (N_3103,In_1958,In_528);
nand U3104 (N_3104,In_361,In_840);
nand U3105 (N_3105,In_933,In_1079);
xor U3106 (N_3106,In_122,In_1669);
nor U3107 (N_3107,In_357,In_1539);
or U3108 (N_3108,In_1082,In_2);
xnor U3109 (N_3109,In_1043,In_164);
nor U3110 (N_3110,In_357,In_9);
nand U3111 (N_3111,In_1822,In_825);
nand U3112 (N_3112,In_1874,In_1901);
nand U3113 (N_3113,In_1611,In_296);
nand U3114 (N_3114,In_934,In_818);
or U3115 (N_3115,In_526,In_1425);
nor U3116 (N_3116,In_1671,In_1466);
xor U3117 (N_3117,In_723,In_1620);
and U3118 (N_3118,In_1955,In_1768);
xnor U3119 (N_3119,In_904,In_1859);
nand U3120 (N_3120,In_310,In_1013);
nor U3121 (N_3121,In_1825,In_1008);
nor U3122 (N_3122,In_1273,In_1485);
nand U3123 (N_3123,In_1801,In_680);
xnor U3124 (N_3124,In_179,In_716);
and U3125 (N_3125,In_9,In_916);
nand U3126 (N_3126,In_1488,In_1231);
nand U3127 (N_3127,In_1048,In_726);
nand U3128 (N_3128,In_658,In_1652);
or U3129 (N_3129,In_732,In_1442);
nor U3130 (N_3130,In_156,In_716);
and U3131 (N_3131,In_238,In_467);
nor U3132 (N_3132,In_1966,In_1373);
xnor U3133 (N_3133,In_265,In_446);
xnor U3134 (N_3134,In_1301,In_1766);
and U3135 (N_3135,In_1998,In_1269);
nor U3136 (N_3136,In_483,In_248);
nand U3137 (N_3137,In_1871,In_1280);
nor U3138 (N_3138,In_1599,In_435);
and U3139 (N_3139,In_748,In_1824);
nor U3140 (N_3140,In_424,In_1859);
nor U3141 (N_3141,In_984,In_1542);
nand U3142 (N_3142,In_1509,In_1058);
nor U3143 (N_3143,In_473,In_989);
or U3144 (N_3144,In_387,In_1504);
or U3145 (N_3145,In_1527,In_1487);
nor U3146 (N_3146,In_1010,In_1266);
xor U3147 (N_3147,In_15,In_1460);
xor U3148 (N_3148,In_1510,In_588);
xor U3149 (N_3149,In_720,In_1891);
nand U3150 (N_3150,In_343,In_1214);
nand U3151 (N_3151,In_1339,In_569);
nor U3152 (N_3152,In_130,In_1880);
and U3153 (N_3153,In_61,In_1495);
or U3154 (N_3154,In_1058,In_1220);
and U3155 (N_3155,In_376,In_597);
and U3156 (N_3156,In_493,In_976);
xor U3157 (N_3157,In_484,In_875);
xor U3158 (N_3158,In_1782,In_292);
and U3159 (N_3159,In_590,In_1084);
nand U3160 (N_3160,In_1020,In_1385);
xor U3161 (N_3161,In_259,In_660);
nor U3162 (N_3162,In_886,In_1690);
nand U3163 (N_3163,In_298,In_473);
nand U3164 (N_3164,In_752,In_461);
nand U3165 (N_3165,In_781,In_346);
nor U3166 (N_3166,In_571,In_1825);
nand U3167 (N_3167,In_1726,In_1134);
xnor U3168 (N_3168,In_1492,In_1403);
or U3169 (N_3169,In_576,In_1675);
nor U3170 (N_3170,In_437,In_573);
nand U3171 (N_3171,In_609,In_1499);
or U3172 (N_3172,In_693,In_1127);
nor U3173 (N_3173,In_1393,In_1707);
nand U3174 (N_3174,In_798,In_90);
or U3175 (N_3175,In_828,In_1334);
xor U3176 (N_3176,In_1516,In_581);
and U3177 (N_3177,In_1638,In_1458);
or U3178 (N_3178,In_956,In_713);
nand U3179 (N_3179,In_1676,In_963);
nor U3180 (N_3180,In_1902,In_1723);
xnor U3181 (N_3181,In_1568,In_1138);
nor U3182 (N_3182,In_1406,In_5);
nor U3183 (N_3183,In_385,In_1773);
and U3184 (N_3184,In_1787,In_657);
xor U3185 (N_3185,In_1231,In_1906);
nor U3186 (N_3186,In_896,In_857);
or U3187 (N_3187,In_1075,In_1617);
nor U3188 (N_3188,In_253,In_855);
nor U3189 (N_3189,In_1773,In_1653);
nand U3190 (N_3190,In_701,In_1989);
and U3191 (N_3191,In_609,In_1287);
and U3192 (N_3192,In_1233,In_1666);
or U3193 (N_3193,In_1621,In_556);
and U3194 (N_3194,In_580,In_1500);
nor U3195 (N_3195,In_1965,In_1089);
nand U3196 (N_3196,In_1352,In_1817);
nand U3197 (N_3197,In_389,In_709);
or U3198 (N_3198,In_324,In_196);
and U3199 (N_3199,In_1573,In_557);
nand U3200 (N_3200,In_1902,In_1437);
nor U3201 (N_3201,In_1598,In_73);
xor U3202 (N_3202,In_440,In_802);
nor U3203 (N_3203,In_1837,In_624);
xor U3204 (N_3204,In_1735,In_525);
nor U3205 (N_3205,In_192,In_1419);
nor U3206 (N_3206,In_944,In_1483);
and U3207 (N_3207,In_683,In_43);
nand U3208 (N_3208,In_1844,In_68);
or U3209 (N_3209,In_417,In_1552);
or U3210 (N_3210,In_627,In_573);
xor U3211 (N_3211,In_1907,In_1481);
nor U3212 (N_3212,In_1956,In_1369);
or U3213 (N_3213,In_1964,In_1264);
xnor U3214 (N_3214,In_905,In_1687);
xor U3215 (N_3215,In_441,In_1573);
nor U3216 (N_3216,In_66,In_1673);
and U3217 (N_3217,In_254,In_574);
nand U3218 (N_3218,In_1752,In_1847);
or U3219 (N_3219,In_1369,In_1029);
and U3220 (N_3220,In_1019,In_1616);
and U3221 (N_3221,In_1286,In_369);
nand U3222 (N_3222,In_275,In_658);
or U3223 (N_3223,In_1967,In_25);
or U3224 (N_3224,In_233,In_678);
nand U3225 (N_3225,In_607,In_398);
or U3226 (N_3226,In_858,In_1276);
xor U3227 (N_3227,In_1376,In_1927);
and U3228 (N_3228,In_200,In_535);
and U3229 (N_3229,In_1626,In_1159);
and U3230 (N_3230,In_1465,In_1761);
nand U3231 (N_3231,In_940,In_1689);
xnor U3232 (N_3232,In_1848,In_176);
nand U3233 (N_3233,In_1478,In_1631);
and U3234 (N_3234,In_1551,In_1627);
nor U3235 (N_3235,In_530,In_409);
or U3236 (N_3236,In_344,In_1917);
xnor U3237 (N_3237,In_777,In_827);
xor U3238 (N_3238,In_1482,In_660);
and U3239 (N_3239,In_560,In_1037);
or U3240 (N_3240,In_884,In_1365);
and U3241 (N_3241,In_1440,In_979);
xnor U3242 (N_3242,In_655,In_1552);
nor U3243 (N_3243,In_423,In_471);
xor U3244 (N_3244,In_5,In_861);
xnor U3245 (N_3245,In_800,In_1972);
and U3246 (N_3246,In_986,In_1106);
nand U3247 (N_3247,In_1249,In_940);
and U3248 (N_3248,In_1734,In_24);
xor U3249 (N_3249,In_486,In_296);
and U3250 (N_3250,In_1339,In_852);
and U3251 (N_3251,In_183,In_565);
or U3252 (N_3252,In_535,In_906);
nor U3253 (N_3253,In_899,In_324);
or U3254 (N_3254,In_548,In_1771);
or U3255 (N_3255,In_1868,In_1335);
or U3256 (N_3256,In_509,In_755);
nor U3257 (N_3257,In_1537,In_1334);
nand U3258 (N_3258,In_733,In_1790);
nand U3259 (N_3259,In_1155,In_1765);
or U3260 (N_3260,In_1958,In_265);
or U3261 (N_3261,In_113,In_562);
nor U3262 (N_3262,In_171,In_1288);
nor U3263 (N_3263,In_124,In_669);
xor U3264 (N_3264,In_1230,In_1542);
xnor U3265 (N_3265,In_1040,In_961);
xnor U3266 (N_3266,In_759,In_339);
and U3267 (N_3267,In_980,In_930);
nor U3268 (N_3268,In_60,In_1534);
xnor U3269 (N_3269,In_902,In_439);
or U3270 (N_3270,In_672,In_499);
and U3271 (N_3271,In_162,In_939);
and U3272 (N_3272,In_51,In_1978);
nand U3273 (N_3273,In_1061,In_829);
xor U3274 (N_3274,In_1018,In_214);
and U3275 (N_3275,In_1552,In_1881);
and U3276 (N_3276,In_1588,In_1125);
or U3277 (N_3277,In_1698,In_29);
nand U3278 (N_3278,In_362,In_945);
nor U3279 (N_3279,In_610,In_298);
or U3280 (N_3280,In_321,In_1972);
and U3281 (N_3281,In_739,In_1161);
nand U3282 (N_3282,In_362,In_638);
xor U3283 (N_3283,In_1253,In_1487);
or U3284 (N_3284,In_1401,In_1750);
nor U3285 (N_3285,In_1628,In_333);
xor U3286 (N_3286,In_453,In_661);
nor U3287 (N_3287,In_721,In_1727);
nand U3288 (N_3288,In_82,In_62);
and U3289 (N_3289,In_1575,In_1942);
and U3290 (N_3290,In_1820,In_691);
or U3291 (N_3291,In_1868,In_261);
and U3292 (N_3292,In_1370,In_438);
and U3293 (N_3293,In_1059,In_1840);
nand U3294 (N_3294,In_1168,In_48);
nand U3295 (N_3295,In_880,In_393);
or U3296 (N_3296,In_1017,In_1882);
and U3297 (N_3297,In_423,In_124);
xnor U3298 (N_3298,In_1277,In_1531);
or U3299 (N_3299,In_403,In_916);
nor U3300 (N_3300,In_1005,In_1316);
nand U3301 (N_3301,In_1311,In_1473);
xor U3302 (N_3302,In_649,In_239);
xnor U3303 (N_3303,In_532,In_916);
nor U3304 (N_3304,In_1885,In_995);
nor U3305 (N_3305,In_1214,In_1190);
xor U3306 (N_3306,In_1097,In_1766);
xor U3307 (N_3307,In_1503,In_1779);
or U3308 (N_3308,In_104,In_1084);
or U3309 (N_3309,In_418,In_699);
nand U3310 (N_3310,In_367,In_1352);
and U3311 (N_3311,In_899,In_1455);
nand U3312 (N_3312,In_1134,In_598);
and U3313 (N_3313,In_599,In_1762);
and U3314 (N_3314,In_332,In_1415);
xor U3315 (N_3315,In_1860,In_725);
or U3316 (N_3316,In_811,In_1300);
nor U3317 (N_3317,In_1933,In_1029);
nand U3318 (N_3318,In_1144,In_291);
or U3319 (N_3319,In_1596,In_1694);
nand U3320 (N_3320,In_1736,In_634);
nor U3321 (N_3321,In_1459,In_337);
and U3322 (N_3322,In_367,In_1380);
and U3323 (N_3323,In_1132,In_86);
nand U3324 (N_3324,In_1064,In_1602);
and U3325 (N_3325,In_1632,In_1768);
and U3326 (N_3326,In_1370,In_1377);
xnor U3327 (N_3327,In_1403,In_1125);
xor U3328 (N_3328,In_997,In_1009);
xor U3329 (N_3329,In_684,In_870);
or U3330 (N_3330,In_1646,In_788);
nor U3331 (N_3331,In_1120,In_1601);
or U3332 (N_3332,In_1168,In_837);
and U3333 (N_3333,In_468,In_52);
xor U3334 (N_3334,In_739,In_1326);
nand U3335 (N_3335,In_1963,In_436);
nor U3336 (N_3336,In_791,In_1267);
or U3337 (N_3337,In_371,In_1374);
xor U3338 (N_3338,In_1564,In_546);
nor U3339 (N_3339,In_1877,In_1751);
nor U3340 (N_3340,In_1776,In_1906);
nand U3341 (N_3341,In_918,In_995);
or U3342 (N_3342,In_1136,In_1433);
or U3343 (N_3343,In_985,In_131);
or U3344 (N_3344,In_1027,In_854);
or U3345 (N_3345,In_1595,In_737);
xor U3346 (N_3346,In_41,In_353);
or U3347 (N_3347,In_375,In_1933);
nor U3348 (N_3348,In_74,In_286);
nor U3349 (N_3349,In_1784,In_1101);
xnor U3350 (N_3350,In_1382,In_965);
or U3351 (N_3351,In_513,In_210);
or U3352 (N_3352,In_973,In_697);
or U3353 (N_3353,In_467,In_471);
or U3354 (N_3354,In_1523,In_608);
xnor U3355 (N_3355,In_1837,In_816);
nor U3356 (N_3356,In_728,In_396);
xnor U3357 (N_3357,In_1462,In_1530);
and U3358 (N_3358,In_1365,In_522);
nor U3359 (N_3359,In_1705,In_339);
or U3360 (N_3360,In_649,In_337);
or U3361 (N_3361,In_1053,In_1886);
nand U3362 (N_3362,In_371,In_1490);
or U3363 (N_3363,In_1992,In_1751);
or U3364 (N_3364,In_1962,In_1726);
and U3365 (N_3365,In_748,In_1729);
nor U3366 (N_3366,In_195,In_800);
nor U3367 (N_3367,In_1677,In_1406);
nand U3368 (N_3368,In_139,In_1008);
nor U3369 (N_3369,In_70,In_1579);
or U3370 (N_3370,In_630,In_1509);
or U3371 (N_3371,In_34,In_1038);
or U3372 (N_3372,In_95,In_1752);
and U3373 (N_3373,In_123,In_844);
or U3374 (N_3374,In_931,In_817);
nor U3375 (N_3375,In_1398,In_209);
nor U3376 (N_3376,In_434,In_739);
nor U3377 (N_3377,In_462,In_312);
and U3378 (N_3378,In_1874,In_1017);
or U3379 (N_3379,In_1094,In_534);
nor U3380 (N_3380,In_1494,In_255);
and U3381 (N_3381,In_309,In_1233);
nand U3382 (N_3382,In_1377,In_1872);
or U3383 (N_3383,In_566,In_973);
xnor U3384 (N_3384,In_671,In_1249);
or U3385 (N_3385,In_1340,In_362);
or U3386 (N_3386,In_907,In_565);
or U3387 (N_3387,In_34,In_971);
nor U3388 (N_3388,In_1758,In_1336);
and U3389 (N_3389,In_1084,In_1148);
nor U3390 (N_3390,In_1202,In_270);
nand U3391 (N_3391,In_376,In_72);
xnor U3392 (N_3392,In_1950,In_562);
and U3393 (N_3393,In_1763,In_1328);
and U3394 (N_3394,In_75,In_1732);
nand U3395 (N_3395,In_1705,In_1454);
and U3396 (N_3396,In_532,In_1894);
or U3397 (N_3397,In_739,In_1760);
or U3398 (N_3398,In_1472,In_1110);
nor U3399 (N_3399,In_793,In_868);
and U3400 (N_3400,In_973,In_1054);
xor U3401 (N_3401,In_1949,In_986);
or U3402 (N_3402,In_40,In_427);
xnor U3403 (N_3403,In_982,In_1476);
or U3404 (N_3404,In_1956,In_1465);
nor U3405 (N_3405,In_1437,In_649);
and U3406 (N_3406,In_1091,In_221);
nor U3407 (N_3407,In_1279,In_345);
xor U3408 (N_3408,In_1259,In_749);
or U3409 (N_3409,In_615,In_1477);
nand U3410 (N_3410,In_219,In_1492);
xor U3411 (N_3411,In_886,In_193);
nand U3412 (N_3412,In_1876,In_1092);
nor U3413 (N_3413,In_686,In_1117);
and U3414 (N_3414,In_1221,In_541);
or U3415 (N_3415,In_804,In_1530);
and U3416 (N_3416,In_1762,In_1528);
and U3417 (N_3417,In_1163,In_1079);
or U3418 (N_3418,In_244,In_125);
nor U3419 (N_3419,In_1926,In_56);
nor U3420 (N_3420,In_1345,In_486);
or U3421 (N_3421,In_1475,In_70);
nor U3422 (N_3422,In_1074,In_963);
and U3423 (N_3423,In_95,In_1347);
nand U3424 (N_3424,In_408,In_1252);
nor U3425 (N_3425,In_1539,In_1069);
nand U3426 (N_3426,In_362,In_335);
xor U3427 (N_3427,In_637,In_844);
or U3428 (N_3428,In_1805,In_129);
xor U3429 (N_3429,In_1008,In_595);
or U3430 (N_3430,In_414,In_425);
xor U3431 (N_3431,In_951,In_1222);
or U3432 (N_3432,In_671,In_1586);
nand U3433 (N_3433,In_682,In_1618);
and U3434 (N_3434,In_1433,In_1905);
and U3435 (N_3435,In_855,In_497);
xor U3436 (N_3436,In_1355,In_407);
nand U3437 (N_3437,In_1231,In_1447);
nor U3438 (N_3438,In_561,In_1294);
and U3439 (N_3439,In_1501,In_1843);
or U3440 (N_3440,In_555,In_1579);
xnor U3441 (N_3441,In_1708,In_434);
xnor U3442 (N_3442,In_1703,In_1388);
nand U3443 (N_3443,In_1115,In_725);
xor U3444 (N_3444,In_1977,In_1804);
xor U3445 (N_3445,In_266,In_422);
xnor U3446 (N_3446,In_361,In_937);
and U3447 (N_3447,In_386,In_1884);
or U3448 (N_3448,In_1531,In_296);
xor U3449 (N_3449,In_785,In_1354);
xnor U3450 (N_3450,In_274,In_1363);
nor U3451 (N_3451,In_386,In_1800);
xor U3452 (N_3452,In_1315,In_1138);
nor U3453 (N_3453,In_965,In_1183);
nor U3454 (N_3454,In_761,In_462);
xor U3455 (N_3455,In_1239,In_1925);
nor U3456 (N_3456,In_802,In_169);
xnor U3457 (N_3457,In_411,In_297);
nand U3458 (N_3458,In_1971,In_1856);
nand U3459 (N_3459,In_1716,In_1948);
nand U3460 (N_3460,In_287,In_1129);
and U3461 (N_3461,In_1487,In_461);
and U3462 (N_3462,In_1323,In_1707);
nand U3463 (N_3463,In_1111,In_934);
nand U3464 (N_3464,In_1169,In_1028);
or U3465 (N_3465,In_26,In_1441);
nor U3466 (N_3466,In_807,In_257);
nand U3467 (N_3467,In_1706,In_1266);
xor U3468 (N_3468,In_817,In_1282);
nor U3469 (N_3469,In_1483,In_977);
nand U3470 (N_3470,In_1435,In_409);
nor U3471 (N_3471,In_595,In_763);
xor U3472 (N_3472,In_1465,In_708);
nor U3473 (N_3473,In_1652,In_937);
or U3474 (N_3474,In_25,In_997);
nor U3475 (N_3475,In_1284,In_1438);
and U3476 (N_3476,In_1830,In_1226);
xnor U3477 (N_3477,In_633,In_913);
xor U3478 (N_3478,In_1784,In_385);
nor U3479 (N_3479,In_332,In_408);
nor U3480 (N_3480,In_1826,In_1845);
nand U3481 (N_3481,In_679,In_1045);
or U3482 (N_3482,In_558,In_1614);
and U3483 (N_3483,In_989,In_790);
or U3484 (N_3484,In_1111,In_1804);
xnor U3485 (N_3485,In_426,In_836);
xnor U3486 (N_3486,In_1320,In_1717);
nor U3487 (N_3487,In_12,In_1727);
nor U3488 (N_3488,In_421,In_207);
or U3489 (N_3489,In_436,In_1663);
nor U3490 (N_3490,In_1379,In_1212);
nor U3491 (N_3491,In_1883,In_852);
or U3492 (N_3492,In_102,In_415);
nor U3493 (N_3493,In_1653,In_122);
xnor U3494 (N_3494,In_516,In_896);
nor U3495 (N_3495,In_1160,In_467);
or U3496 (N_3496,In_42,In_1402);
or U3497 (N_3497,In_1659,In_1084);
or U3498 (N_3498,In_1697,In_148);
nor U3499 (N_3499,In_1557,In_573);
or U3500 (N_3500,In_1746,In_62);
or U3501 (N_3501,In_1624,In_59);
and U3502 (N_3502,In_1054,In_1571);
nand U3503 (N_3503,In_426,In_838);
xnor U3504 (N_3504,In_832,In_1971);
nand U3505 (N_3505,In_834,In_639);
and U3506 (N_3506,In_990,In_406);
and U3507 (N_3507,In_345,In_1039);
or U3508 (N_3508,In_1660,In_1027);
xor U3509 (N_3509,In_1170,In_1067);
nand U3510 (N_3510,In_1962,In_1897);
nand U3511 (N_3511,In_1377,In_1830);
nand U3512 (N_3512,In_1620,In_970);
xor U3513 (N_3513,In_1840,In_476);
nor U3514 (N_3514,In_1833,In_646);
or U3515 (N_3515,In_1513,In_1743);
and U3516 (N_3516,In_344,In_1648);
and U3517 (N_3517,In_1155,In_1295);
xnor U3518 (N_3518,In_1686,In_1346);
and U3519 (N_3519,In_1446,In_635);
or U3520 (N_3520,In_1318,In_546);
and U3521 (N_3521,In_1211,In_1430);
and U3522 (N_3522,In_456,In_1235);
xnor U3523 (N_3523,In_944,In_1864);
or U3524 (N_3524,In_724,In_877);
nor U3525 (N_3525,In_1497,In_774);
and U3526 (N_3526,In_1339,In_67);
xor U3527 (N_3527,In_708,In_1244);
nand U3528 (N_3528,In_1573,In_449);
xor U3529 (N_3529,In_1693,In_1195);
nor U3530 (N_3530,In_1866,In_636);
nor U3531 (N_3531,In_1516,In_1151);
nand U3532 (N_3532,In_602,In_270);
xor U3533 (N_3533,In_569,In_722);
and U3534 (N_3534,In_1145,In_927);
and U3535 (N_3535,In_1759,In_868);
or U3536 (N_3536,In_963,In_1174);
xnor U3537 (N_3537,In_1765,In_1208);
xnor U3538 (N_3538,In_1566,In_1956);
xnor U3539 (N_3539,In_494,In_1172);
or U3540 (N_3540,In_1042,In_749);
xor U3541 (N_3541,In_1454,In_1219);
nor U3542 (N_3542,In_729,In_959);
nand U3543 (N_3543,In_720,In_194);
or U3544 (N_3544,In_162,In_990);
or U3545 (N_3545,In_1968,In_1217);
or U3546 (N_3546,In_1063,In_1229);
nand U3547 (N_3547,In_1797,In_195);
nor U3548 (N_3548,In_349,In_782);
nor U3549 (N_3549,In_86,In_1730);
and U3550 (N_3550,In_953,In_1286);
or U3551 (N_3551,In_1008,In_1102);
or U3552 (N_3552,In_1894,In_1900);
nor U3553 (N_3553,In_1980,In_184);
or U3554 (N_3554,In_245,In_1503);
nor U3555 (N_3555,In_1198,In_1979);
nand U3556 (N_3556,In_839,In_403);
xor U3557 (N_3557,In_1699,In_917);
nand U3558 (N_3558,In_1999,In_1706);
xor U3559 (N_3559,In_926,In_929);
nor U3560 (N_3560,In_1102,In_1840);
nand U3561 (N_3561,In_1011,In_653);
xor U3562 (N_3562,In_1248,In_1679);
xor U3563 (N_3563,In_448,In_1553);
nor U3564 (N_3564,In_1994,In_562);
xnor U3565 (N_3565,In_134,In_180);
or U3566 (N_3566,In_996,In_636);
xor U3567 (N_3567,In_757,In_787);
nand U3568 (N_3568,In_1681,In_1336);
nor U3569 (N_3569,In_1312,In_952);
and U3570 (N_3570,In_315,In_71);
nand U3571 (N_3571,In_1318,In_1187);
xnor U3572 (N_3572,In_1461,In_1274);
and U3573 (N_3573,In_43,In_517);
nor U3574 (N_3574,In_788,In_956);
xor U3575 (N_3575,In_286,In_898);
xnor U3576 (N_3576,In_415,In_1556);
and U3577 (N_3577,In_640,In_1591);
nand U3578 (N_3578,In_1984,In_1887);
xnor U3579 (N_3579,In_1251,In_1048);
or U3580 (N_3580,In_1913,In_551);
xnor U3581 (N_3581,In_873,In_1531);
nand U3582 (N_3582,In_1640,In_44);
xor U3583 (N_3583,In_182,In_1717);
and U3584 (N_3584,In_612,In_103);
nor U3585 (N_3585,In_61,In_1149);
or U3586 (N_3586,In_851,In_946);
nor U3587 (N_3587,In_637,In_756);
xor U3588 (N_3588,In_984,In_351);
or U3589 (N_3589,In_1896,In_582);
or U3590 (N_3590,In_1815,In_1501);
nand U3591 (N_3591,In_868,In_41);
or U3592 (N_3592,In_1440,In_978);
and U3593 (N_3593,In_1774,In_1579);
and U3594 (N_3594,In_1188,In_390);
nor U3595 (N_3595,In_760,In_1178);
nand U3596 (N_3596,In_1086,In_1768);
and U3597 (N_3597,In_776,In_1112);
nand U3598 (N_3598,In_340,In_300);
nand U3599 (N_3599,In_352,In_619);
nand U3600 (N_3600,In_468,In_1622);
xor U3601 (N_3601,In_1146,In_61);
xnor U3602 (N_3602,In_1375,In_1268);
xor U3603 (N_3603,In_1473,In_1231);
nand U3604 (N_3604,In_1272,In_31);
nand U3605 (N_3605,In_1191,In_1452);
and U3606 (N_3606,In_979,In_58);
nand U3607 (N_3607,In_475,In_828);
nor U3608 (N_3608,In_1884,In_1556);
nor U3609 (N_3609,In_86,In_1563);
xnor U3610 (N_3610,In_386,In_897);
nand U3611 (N_3611,In_104,In_1649);
or U3612 (N_3612,In_689,In_90);
nor U3613 (N_3613,In_1379,In_1207);
nor U3614 (N_3614,In_351,In_1565);
nand U3615 (N_3615,In_1426,In_683);
and U3616 (N_3616,In_1163,In_1273);
nand U3617 (N_3617,In_1001,In_1058);
nor U3618 (N_3618,In_1107,In_1145);
nor U3619 (N_3619,In_1480,In_958);
or U3620 (N_3620,In_589,In_1748);
and U3621 (N_3621,In_668,In_1038);
nor U3622 (N_3622,In_74,In_1986);
and U3623 (N_3623,In_1969,In_399);
and U3624 (N_3624,In_624,In_1800);
nand U3625 (N_3625,In_1896,In_557);
xor U3626 (N_3626,In_1109,In_117);
and U3627 (N_3627,In_1661,In_663);
or U3628 (N_3628,In_334,In_148);
nor U3629 (N_3629,In_1992,In_1792);
nand U3630 (N_3630,In_965,In_1141);
xor U3631 (N_3631,In_1179,In_1613);
xnor U3632 (N_3632,In_9,In_1548);
or U3633 (N_3633,In_964,In_1740);
nor U3634 (N_3634,In_1790,In_1398);
xnor U3635 (N_3635,In_128,In_294);
nor U3636 (N_3636,In_762,In_1665);
and U3637 (N_3637,In_527,In_1423);
or U3638 (N_3638,In_1431,In_116);
and U3639 (N_3639,In_1181,In_838);
and U3640 (N_3640,In_281,In_1260);
nor U3641 (N_3641,In_797,In_81);
nand U3642 (N_3642,In_602,In_1152);
or U3643 (N_3643,In_201,In_651);
xnor U3644 (N_3644,In_792,In_151);
or U3645 (N_3645,In_833,In_261);
nand U3646 (N_3646,In_708,In_210);
or U3647 (N_3647,In_1713,In_1141);
or U3648 (N_3648,In_994,In_270);
xnor U3649 (N_3649,In_745,In_1560);
xor U3650 (N_3650,In_1805,In_557);
nor U3651 (N_3651,In_587,In_909);
xnor U3652 (N_3652,In_1789,In_305);
nor U3653 (N_3653,In_1102,In_1220);
nor U3654 (N_3654,In_1375,In_51);
nand U3655 (N_3655,In_198,In_2);
xor U3656 (N_3656,In_1859,In_1324);
nor U3657 (N_3657,In_1243,In_1206);
nor U3658 (N_3658,In_1023,In_1758);
nor U3659 (N_3659,In_980,In_658);
or U3660 (N_3660,In_98,In_1811);
nor U3661 (N_3661,In_1684,In_1936);
xor U3662 (N_3662,In_1841,In_1267);
nand U3663 (N_3663,In_1831,In_1972);
nor U3664 (N_3664,In_1054,In_1243);
nor U3665 (N_3665,In_1252,In_1611);
nor U3666 (N_3666,In_1083,In_693);
nor U3667 (N_3667,In_1873,In_754);
and U3668 (N_3668,In_1773,In_719);
or U3669 (N_3669,In_452,In_1148);
nor U3670 (N_3670,In_794,In_1962);
xnor U3671 (N_3671,In_1959,In_1822);
or U3672 (N_3672,In_1820,In_796);
nor U3673 (N_3673,In_605,In_815);
and U3674 (N_3674,In_1394,In_1263);
xor U3675 (N_3675,In_572,In_1497);
nand U3676 (N_3676,In_1758,In_992);
xnor U3677 (N_3677,In_1862,In_1645);
nand U3678 (N_3678,In_806,In_944);
or U3679 (N_3679,In_423,In_956);
and U3680 (N_3680,In_1767,In_1690);
nand U3681 (N_3681,In_1664,In_392);
xnor U3682 (N_3682,In_162,In_860);
nor U3683 (N_3683,In_1508,In_735);
nor U3684 (N_3684,In_1800,In_1868);
nor U3685 (N_3685,In_1682,In_547);
xnor U3686 (N_3686,In_1841,In_776);
xnor U3687 (N_3687,In_1943,In_1047);
xnor U3688 (N_3688,In_1154,In_587);
nand U3689 (N_3689,In_1632,In_301);
xnor U3690 (N_3690,In_1927,In_1511);
nand U3691 (N_3691,In_1241,In_1458);
and U3692 (N_3692,In_1164,In_488);
nand U3693 (N_3693,In_1054,In_550);
and U3694 (N_3694,In_1171,In_343);
nand U3695 (N_3695,In_969,In_684);
nand U3696 (N_3696,In_1170,In_1562);
or U3697 (N_3697,In_1205,In_1243);
and U3698 (N_3698,In_476,In_321);
or U3699 (N_3699,In_1461,In_336);
nor U3700 (N_3700,In_965,In_279);
and U3701 (N_3701,In_861,In_237);
nand U3702 (N_3702,In_1005,In_1998);
and U3703 (N_3703,In_260,In_895);
xnor U3704 (N_3704,In_1327,In_1844);
and U3705 (N_3705,In_867,In_1350);
nor U3706 (N_3706,In_736,In_1249);
nand U3707 (N_3707,In_684,In_1413);
xor U3708 (N_3708,In_1501,In_1934);
xnor U3709 (N_3709,In_752,In_1224);
or U3710 (N_3710,In_1422,In_1178);
or U3711 (N_3711,In_891,In_264);
nand U3712 (N_3712,In_1991,In_1241);
or U3713 (N_3713,In_1721,In_414);
nor U3714 (N_3714,In_677,In_1428);
xnor U3715 (N_3715,In_1393,In_1213);
nor U3716 (N_3716,In_438,In_134);
nor U3717 (N_3717,In_806,In_794);
xor U3718 (N_3718,In_1769,In_676);
nand U3719 (N_3719,In_1754,In_733);
xnor U3720 (N_3720,In_1818,In_1784);
nand U3721 (N_3721,In_1491,In_774);
or U3722 (N_3722,In_1961,In_81);
nor U3723 (N_3723,In_1191,In_565);
xor U3724 (N_3724,In_108,In_298);
nand U3725 (N_3725,In_329,In_1966);
and U3726 (N_3726,In_486,In_1221);
and U3727 (N_3727,In_131,In_271);
xnor U3728 (N_3728,In_551,In_172);
nand U3729 (N_3729,In_162,In_822);
nor U3730 (N_3730,In_1259,In_882);
nand U3731 (N_3731,In_315,In_1573);
nand U3732 (N_3732,In_522,In_105);
and U3733 (N_3733,In_14,In_1763);
nand U3734 (N_3734,In_864,In_752);
nand U3735 (N_3735,In_245,In_419);
and U3736 (N_3736,In_1837,In_1318);
nor U3737 (N_3737,In_931,In_1621);
nor U3738 (N_3738,In_1670,In_39);
nand U3739 (N_3739,In_1589,In_1837);
xor U3740 (N_3740,In_813,In_357);
nor U3741 (N_3741,In_0,In_387);
nor U3742 (N_3742,In_1838,In_755);
nor U3743 (N_3743,In_824,In_1471);
xnor U3744 (N_3744,In_632,In_861);
xnor U3745 (N_3745,In_1105,In_474);
nand U3746 (N_3746,In_1547,In_679);
nand U3747 (N_3747,In_1058,In_330);
nand U3748 (N_3748,In_959,In_1446);
nor U3749 (N_3749,In_1797,In_632);
nor U3750 (N_3750,In_754,In_1348);
nand U3751 (N_3751,In_1875,In_314);
or U3752 (N_3752,In_837,In_88);
and U3753 (N_3753,In_629,In_773);
or U3754 (N_3754,In_1170,In_410);
or U3755 (N_3755,In_163,In_1566);
xnor U3756 (N_3756,In_1029,In_644);
nor U3757 (N_3757,In_652,In_833);
or U3758 (N_3758,In_1471,In_875);
xor U3759 (N_3759,In_676,In_817);
and U3760 (N_3760,In_1870,In_1780);
or U3761 (N_3761,In_1382,In_1874);
nand U3762 (N_3762,In_1679,In_351);
xnor U3763 (N_3763,In_1747,In_596);
nand U3764 (N_3764,In_1646,In_771);
and U3765 (N_3765,In_1711,In_1788);
or U3766 (N_3766,In_1382,In_399);
and U3767 (N_3767,In_1496,In_1907);
and U3768 (N_3768,In_378,In_1486);
nand U3769 (N_3769,In_1389,In_1173);
nor U3770 (N_3770,In_1738,In_1082);
xor U3771 (N_3771,In_1814,In_2);
nor U3772 (N_3772,In_306,In_1756);
xor U3773 (N_3773,In_1591,In_265);
nor U3774 (N_3774,In_988,In_1677);
and U3775 (N_3775,In_1019,In_1624);
nor U3776 (N_3776,In_1440,In_518);
xnor U3777 (N_3777,In_347,In_1764);
nor U3778 (N_3778,In_1308,In_866);
xor U3779 (N_3779,In_1304,In_612);
and U3780 (N_3780,In_1698,In_101);
and U3781 (N_3781,In_1131,In_1724);
xor U3782 (N_3782,In_75,In_574);
nor U3783 (N_3783,In_1535,In_267);
or U3784 (N_3784,In_7,In_1353);
nor U3785 (N_3785,In_515,In_1064);
nand U3786 (N_3786,In_1811,In_161);
xnor U3787 (N_3787,In_915,In_660);
xor U3788 (N_3788,In_887,In_158);
or U3789 (N_3789,In_665,In_289);
nand U3790 (N_3790,In_592,In_344);
nor U3791 (N_3791,In_1015,In_1764);
nor U3792 (N_3792,In_1444,In_14);
nand U3793 (N_3793,In_1893,In_74);
and U3794 (N_3794,In_1510,In_1401);
or U3795 (N_3795,In_986,In_1506);
xor U3796 (N_3796,In_1022,In_1481);
or U3797 (N_3797,In_906,In_1473);
nand U3798 (N_3798,In_1603,In_1196);
and U3799 (N_3799,In_1094,In_86);
nand U3800 (N_3800,In_920,In_527);
nor U3801 (N_3801,In_226,In_1663);
or U3802 (N_3802,In_1064,In_764);
or U3803 (N_3803,In_639,In_1731);
nand U3804 (N_3804,In_1070,In_876);
nand U3805 (N_3805,In_1076,In_365);
xnor U3806 (N_3806,In_835,In_44);
or U3807 (N_3807,In_741,In_1553);
or U3808 (N_3808,In_1367,In_812);
xnor U3809 (N_3809,In_928,In_1793);
nor U3810 (N_3810,In_1606,In_1502);
or U3811 (N_3811,In_105,In_575);
xor U3812 (N_3812,In_1460,In_1754);
nand U3813 (N_3813,In_746,In_1702);
nor U3814 (N_3814,In_833,In_872);
xnor U3815 (N_3815,In_647,In_95);
xnor U3816 (N_3816,In_371,In_1079);
or U3817 (N_3817,In_1615,In_530);
or U3818 (N_3818,In_319,In_337);
xnor U3819 (N_3819,In_1181,In_1351);
or U3820 (N_3820,In_1586,In_1013);
or U3821 (N_3821,In_487,In_57);
and U3822 (N_3822,In_1451,In_58);
nor U3823 (N_3823,In_122,In_438);
xnor U3824 (N_3824,In_863,In_1248);
nand U3825 (N_3825,In_1060,In_656);
xnor U3826 (N_3826,In_165,In_76);
nand U3827 (N_3827,In_1418,In_361);
nand U3828 (N_3828,In_275,In_1995);
nor U3829 (N_3829,In_799,In_1456);
nor U3830 (N_3830,In_1847,In_458);
and U3831 (N_3831,In_1917,In_1739);
and U3832 (N_3832,In_658,In_1456);
or U3833 (N_3833,In_1777,In_658);
nand U3834 (N_3834,In_908,In_818);
xnor U3835 (N_3835,In_659,In_1364);
nor U3836 (N_3836,In_1737,In_575);
and U3837 (N_3837,In_1224,In_125);
xor U3838 (N_3838,In_1467,In_1710);
nor U3839 (N_3839,In_454,In_1990);
nor U3840 (N_3840,In_249,In_1899);
or U3841 (N_3841,In_1953,In_1649);
nand U3842 (N_3842,In_484,In_65);
and U3843 (N_3843,In_1595,In_946);
xor U3844 (N_3844,In_955,In_1178);
nor U3845 (N_3845,In_1199,In_1176);
xnor U3846 (N_3846,In_1499,In_1018);
nand U3847 (N_3847,In_497,In_1152);
nor U3848 (N_3848,In_1443,In_902);
nand U3849 (N_3849,In_1321,In_246);
nand U3850 (N_3850,In_1487,In_1662);
nand U3851 (N_3851,In_1959,In_181);
nor U3852 (N_3852,In_976,In_1421);
nand U3853 (N_3853,In_303,In_495);
and U3854 (N_3854,In_1448,In_1540);
and U3855 (N_3855,In_1480,In_1977);
nand U3856 (N_3856,In_1400,In_1646);
xor U3857 (N_3857,In_61,In_1165);
or U3858 (N_3858,In_1468,In_1200);
nor U3859 (N_3859,In_1182,In_924);
nand U3860 (N_3860,In_1849,In_1063);
nand U3861 (N_3861,In_336,In_1577);
or U3862 (N_3862,In_581,In_448);
and U3863 (N_3863,In_1613,In_1928);
xor U3864 (N_3864,In_494,In_1755);
nand U3865 (N_3865,In_624,In_1213);
or U3866 (N_3866,In_1000,In_1360);
or U3867 (N_3867,In_1123,In_725);
nor U3868 (N_3868,In_717,In_704);
xnor U3869 (N_3869,In_103,In_351);
or U3870 (N_3870,In_1915,In_1335);
or U3871 (N_3871,In_444,In_1255);
nand U3872 (N_3872,In_653,In_1470);
nand U3873 (N_3873,In_154,In_1957);
nor U3874 (N_3874,In_1931,In_899);
and U3875 (N_3875,In_245,In_1005);
nor U3876 (N_3876,In_1340,In_372);
and U3877 (N_3877,In_1647,In_760);
nand U3878 (N_3878,In_963,In_229);
and U3879 (N_3879,In_991,In_1370);
nand U3880 (N_3880,In_349,In_964);
xnor U3881 (N_3881,In_1073,In_483);
or U3882 (N_3882,In_1232,In_354);
nor U3883 (N_3883,In_1011,In_944);
or U3884 (N_3884,In_489,In_334);
nand U3885 (N_3885,In_1919,In_918);
and U3886 (N_3886,In_1228,In_1933);
xnor U3887 (N_3887,In_292,In_183);
or U3888 (N_3888,In_198,In_216);
and U3889 (N_3889,In_564,In_792);
nor U3890 (N_3890,In_569,In_641);
xor U3891 (N_3891,In_1809,In_1399);
or U3892 (N_3892,In_621,In_340);
nor U3893 (N_3893,In_872,In_1111);
nand U3894 (N_3894,In_990,In_811);
or U3895 (N_3895,In_683,In_106);
nor U3896 (N_3896,In_67,In_1706);
or U3897 (N_3897,In_532,In_164);
or U3898 (N_3898,In_84,In_1735);
xnor U3899 (N_3899,In_1130,In_1192);
and U3900 (N_3900,In_928,In_143);
xnor U3901 (N_3901,In_1062,In_1083);
and U3902 (N_3902,In_1761,In_612);
and U3903 (N_3903,In_417,In_1162);
and U3904 (N_3904,In_1763,In_181);
and U3905 (N_3905,In_1845,In_392);
or U3906 (N_3906,In_1572,In_1334);
xnor U3907 (N_3907,In_1432,In_1145);
xnor U3908 (N_3908,In_1799,In_710);
nor U3909 (N_3909,In_62,In_1834);
nor U3910 (N_3910,In_178,In_1879);
nor U3911 (N_3911,In_1133,In_593);
nor U3912 (N_3912,In_408,In_1812);
or U3913 (N_3913,In_16,In_78);
and U3914 (N_3914,In_928,In_1612);
nand U3915 (N_3915,In_784,In_1861);
nor U3916 (N_3916,In_346,In_1273);
xor U3917 (N_3917,In_1280,In_1686);
nand U3918 (N_3918,In_1502,In_639);
or U3919 (N_3919,In_1892,In_1381);
nand U3920 (N_3920,In_1120,In_1476);
and U3921 (N_3921,In_82,In_1981);
nor U3922 (N_3922,In_1721,In_248);
or U3923 (N_3923,In_1952,In_1638);
nor U3924 (N_3924,In_1100,In_1580);
nor U3925 (N_3925,In_1676,In_1521);
and U3926 (N_3926,In_1584,In_415);
nor U3927 (N_3927,In_1012,In_1308);
nor U3928 (N_3928,In_1542,In_485);
nand U3929 (N_3929,In_507,In_652);
or U3930 (N_3930,In_958,In_162);
or U3931 (N_3931,In_401,In_232);
xor U3932 (N_3932,In_1084,In_1012);
or U3933 (N_3933,In_1318,In_254);
or U3934 (N_3934,In_1693,In_1902);
nand U3935 (N_3935,In_1843,In_1694);
xor U3936 (N_3936,In_1271,In_667);
or U3937 (N_3937,In_17,In_986);
xor U3938 (N_3938,In_315,In_1449);
or U3939 (N_3939,In_409,In_1194);
xnor U3940 (N_3940,In_627,In_1031);
nand U3941 (N_3941,In_1669,In_182);
or U3942 (N_3942,In_943,In_1796);
or U3943 (N_3943,In_1465,In_926);
nand U3944 (N_3944,In_541,In_1682);
xor U3945 (N_3945,In_1628,In_962);
xor U3946 (N_3946,In_315,In_1471);
nor U3947 (N_3947,In_1446,In_1337);
nand U3948 (N_3948,In_581,In_1159);
or U3949 (N_3949,In_766,In_1766);
and U3950 (N_3950,In_672,In_1836);
nand U3951 (N_3951,In_1078,In_934);
xor U3952 (N_3952,In_1725,In_402);
nand U3953 (N_3953,In_174,In_1265);
and U3954 (N_3954,In_479,In_281);
nor U3955 (N_3955,In_161,In_1136);
xor U3956 (N_3956,In_1635,In_505);
or U3957 (N_3957,In_86,In_22);
or U3958 (N_3958,In_1542,In_1333);
xnor U3959 (N_3959,In_989,In_324);
xnor U3960 (N_3960,In_39,In_1135);
nor U3961 (N_3961,In_1043,In_609);
or U3962 (N_3962,In_651,In_1434);
xor U3963 (N_3963,In_740,In_1123);
nor U3964 (N_3964,In_997,In_805);
nand U3965 (N_3965,In_1994,In_724);
nand U3966 (N_3966,In_1308,In_640);
xor U3967 (N_3967,In_837,In_527);
nand U3968 (N_3968,In_481,In_978);
and U3969 (N_3969,In_906,In_1392);
xnor U3970 (N_3970,In_1699,In_1771);
nor U3971 (N_3971,In_202,In_1150);
xnor U3972 (N_3972,In_1725,In_959);
or U3973 (N_3973,In_1292,In_529);
nand U3974 (N_3974,In_732,In_168);
or U3975 (N_3975,In_1407,In_181);
or U3976 (N_3976,In_1198,In_319);
nor U3977 (N_3977,In_679,In_1316);
and U3978 (N_3978,In_16,In_90);
or U3979 (N_3979,In_786,In_473);
or U3980 (N_3980,In_1253,In_922);
and U3981 (N_3981,In_265,In_1721);
nor U3982 (N_3982,In_1769,In_1986);
xnor U3983 (N_3983,In_701,In_1495);
and U3984 (N_3984,In_1847,In_548);
xnor U3985 (N_3985,In_1613,In_839);
nor U3986 (N_3986,In_1287,In_525);
xor U3987 (N_3987,In_1570,In_589);
nand U3988 (N_3988,In_1626,In_1911);
and U3989 (N_3989,In_1821,In_1733);
xnor U3990 (N_3990,In_1430,In_1402);
nor U3991 (N_3991,In_1882,In_235);
nand U3992 (N_3992,In_354,In_110);
or U3993 (N_3993,In_1342,In_507);
or U3994 (N_3994,In_1089,In_1700);
nor U3995 (N_3995,In_1911,In_1005);
nor U3996 (N_3996,In_907,In_1744);
xor U3997 (N_3997,In_832,In_953);
nand U3998 (N_3998,In_1198,In_277);
xnor U3999 (N_3999,In_1799,In_570);
nand U4000 (N_4000,In_859,In_1504);
xor U4001 (N_4001,In_1317,In_1127);
nor U4002 (N_4002,In_1711,In_682);
nor U4003 (N_4003,In_826,In_753);
xnor U4004 (N_4004,In_787,In_1902);
and U4005 (N_4005,In_1364,In_1600);
nor U4006 (N_4006,In_1528,In_515);
nand U4007 (N_4007,In_1795,In_5);
xor U4008 (N_4008,In_1688,In_338);
nor U4009 (N_4009,In_471,In_809);
nand U4010 (N_4010,In_1144,In_697);
or U4011 (N_4011,In_396,In_189);
or U4012 (N_4012,In_375,In_1969);
nor U4013 (N_4013,In_786,In_1036);
nor U4014 (N_4014,In_1818,In_28);
xor U4015 (N_4015,In_1160,In_131);
and U4016 (N_4016,In_1905,In_157);
and U4017 (N_4017,In_1904,In_1578);
nand U4018 (N_4018,In_475,In_1848);
nand U4019 (N_4019,In_1423,In_1667);
and U4020 (N_4020,In_825,In_1941);
xor U4021 (N_4021,In_842,In_1009);
nor U4022 (N_4022,In_1664,In_1765);
nor U4023 (N_4023,In_423,In_1559);
or U4024 (N_4024,In_397,In_1843);
and U4025 (N_4025,In_689,In_803);
or U4026 (N_4026,In_755,In_1113);
or U4027 (N_4027,In_294,In_1485);
nor U4028 (N_4028,In_1127,In_545);
nand U4029 (N_4029,In_1576,In_652);
and U4030 (N_4030,In_419,In_1658);
or U4031 (N_4031,In_523,In_397);
nor U4032 (N_4032,In_278,In_1995);
and U4033 (N_4033,In_1471,In_840);
xnor U4034 (N_4034,In_1152,In_1784);
nor U4035 (N_4035,In_107,In_349);
nand U4036 (N_4036,In_847,In_1239);
xor U4037 (N_4037,In_1660,In_206);
or U4038 (N_4038,In_1977,In_969);
nand U4039 (N_4039,In_1827,In_1338);
nor U4040 (N_4040,In_740,In_1663);
xor U4041 (N_4041,In_1478,In_1718);
and U4042 (N_4042,In_280,In_647);
nor U4043 (N_4043,In_1627,In_1236);
xnor U4044 (N_4044,In_155,In_1315);
nor U4045 (N_4045,In_615,In_1031);
nand U4046 (N_4046,In_1029,In_365);
and U4047 (N_4047,In_373,In_1317);
or U4048 (N_4048,In_578,In_790);
and U4049 (N_4049,In_1684,In_759);
and U4050 (N_4050,In_401,In_109);
nand U4051 (N_4051,In_72,In_1767);
nor U4052 (N_4052,In_391,In_972);
or U4053 (N_4053,In_1102,In_361);
nor U4054 (N_4054,In_1682,In_963);
xnor U4055 (N_4055,In_1159,In_1144);
and U4056 (N_4056,In_41,In_708);
xnor U4057 (N_4057,In_306,In_575);
or U4058 (N_4058,In_32,In_1901);
nor U4059 (N_4059,In_314,In_1691);
nor U4060 (N_4060,In_106,In_905);
xor U4061 (N_4061,In_86,In_886);
nor U4062 (N_4062,In_618,In_1524);
or U4063 (N_4063,In_1011,In_116);
nand U4064 (N_4064,In_1839,In_773);
xnor U4065 (N_4065,In_1488,In_538);
or U4066 (N_4066,In_598,In_1572);
nor U4067 (N_4067,In_882,In_1459);
or U4068 (N_4068,In_1747,In_712);
nor U4069 (N_4069,In_1178,In_168);
xor U4070 (N_4070,In_310,In_1037);
and U4071 (N_4071,In_536,In_1525);
nor U4072 (N_4072,In_1113,In_182);
nand U4073 (N_4073,In_1715,In_1895);
nand U4074 (N_4074,In_1914,In_1193);
or U4075 (N_4075,In_448,In_1457);
nand U4076 (N_4076,In_268,In_1391);
nor U4077 (N_4077,In_1986,In_1473);
or U4078 (N_4078,In_1678,In_373);
nor U4079 (N_4079,In_582,In_702);
or U4080 (N_4080,In_473,In_1824);
xor U4081 (N_4081,In_1878,In_1562);
nor U4082 (N_4082,In_820,In_1309);
or U4083 (N_4083,In_1520,In_202);
xnor U4084 (N_4084,In_853,In_1275);
nand U4085 (N_4085,In_1672,In_1098);
nand U4086 (N_4086,In_743,In_1918);
and U4087 (N_4087,In_1903,In_648);
nand U4088 (N_4088,In_1272,In_1983);
nand U4089 (N_4089,In_1705,In_43);
or U4090 (N_4090,In_799,In_1096);
and U4091 (N_4091,In_1080,In_353);
nand U4092 (N_4092,In_1421,In_1699);
or U4093 (N_4093,In_1215,In_1851);
or U4094 (N_4094,In_1033,In_1601);
and U4095 (N_4095,In_928,In_1177);
nand U4096 (N_4096,In_1590,In_1258);
xnor U4097 (N_4097,In_1005,In_1562);
nor U4098 (N_4098,In_1049,In_426);
xor U4099 (N_4099,In_1310,In_1014);
nand U4100 (N_4100,In_1452,In_615);
and U4101 (N_4101,In_1704,In_536);
or U4102 (N_4102,In_1196,In_1523);
nor U4103 (N_4103,In_169,In_1201);
nand U4104 (N_4104,In_689,In_1435);
nand U4105 (N_4105,In_900,In_405);
and U4106 (N_4106,In_1101,In_308);
and U4107 (N_4107,In_514,In_1009);
xnor U4108 (N_4108,In_1476,In_1392);
xnor U4109 (N_4109,In_633,In_1603);
or U4110 (N_4110,In_881,In_1903);
nand U4111 (N_4111,In_391,In_969);
xor U4112 (N_4112,In_467,In_727);
nor U4113 (N_4113,In_1960,In_387);
or U4114 (N_4114,In_1664,In_1977);
or U4115 (N_4115,In_1346,In_233);
xnor U4116 (N_4116,In_544,In_685);
xor U4117 (N_4117,In_1840,In_239);
and U4118 (N_4118,In_982,In_1615);
nor U4119 (N_4119,In_575,In_442);
or U4120 (N_4120,In_1308,In_1669);
nor U4121 (N_4121,In_1572,In_1055);
nand U4122 (N_4122,In_134,In_936);
nand U4123 (N_4123,In_27,In_572);
xor U4124 (N_4124,In_2,In_1302);
xor U4125 (N_4125,In_113,In_1545);
xnor U4126 (N_4126,In_481,In_477);
nand U4127 (N_4127,In_995,In_903);
nand U4128 (N_4128,In_1373,In_1090);
nand U4129 (N_4129,In_1439,In_862);
xor U4130 (N_4130,In_825,In_561);
nor U4131 (N_4131,In_808,In_1091);
or U4132 (N_4132,In_1622,In_1825);
and U4133 (N_4133,In_775,In_477);
nand U4134 (N_4134,In_1854,In_1582);
xnor U4135 (N_4135,In_1739,In_1240);
nand U4136 (N_4136,In_1722,In_906);
or U4137 (N_4137,In_1608,In_319);
and U4138 (N_4138,In_684,In_931);
xor U4139 (N_4139,In_611,In_1313);
nand U4140 (N_4140,In_1301,In_117);
nor U4141 (N_4141,In_782,In_424);
or U4142 (N_4142,In_848,In_1269);
nand U4143 (N_4143,In_1846,In_1588);
xor U4144 (N_4144,In_1206,In_1950);
or U4145 (N_4145,In_1518,In_676);
or U4146 (N_4146,In_837,In_1410);
or U4147 (N_4147,In_457,In_836);
nand U4148 (N_4148,In_361,In_635);
and U4149 (N_4149,In_861,In_710);
nand U4150 (N_4150,In_594,In_454);
xor U4151 (N_4151,In_1604,In_372);
xor U4152 (N_4152,In_339,In_321);
xor U4153 (N_4153,In_1434,In_105);
nor U4154 (N_4154,In_1258,In_1002);
or U4155 (N_4155,In_1527,In_1047);
nand U4156 (N_4156,In_625,In_1446);
and U4157 (N_4157,In_810,In_1239);
nand U4158 (N_4158,In_1039,In_1866);
nor U4159 (N_4159,In_965,In_1594);
nor U4160 (N_4160,In_902,In_102);
xor U4161 (N_4161,In_1454,In_1257);
or U4162 (N_4162,In_970,In_351);
nand U4163 (N_4163,In_88,In_794);
or U4164 (N_4164,In_634,In_794);
nand U4165 (N_4165,In_1956,In_1098);
and U4166 (N_4166,In_1668,In_349);
nand U4167 (N_4167,In_448,In_1335);
nand U4168 (N_4168,In_210,In_918);
or U4169 (N_4169,In_1152,In_1165);
nand U4170 (N_4170,In_1950,In_1230);
or U4171 (N_4171,In_1980,In_1624);
and U4172 (N_4172,In_1442,In_1910);
nand U4173 (N_4173,In_620,In_1168);
nor U4174 (N_4174,In_1663,In_633);
nor U4175 (N_4175,In_1349,In_1384);
and U4176 (N_4176,In_658,In_979);
nand U4177 (N_4177,In_98,In_759);
xnor U4178 (N_4178,In_1656,In_12);
or U4179 (N_4179,In_1902,In_1396);
nor U4180 (N_4180,In_532,In_1065);
and U4181 (N_4181,In_1838,In_1074);
nor U4182 (N_4182,In_1511,In_603);
or U4183 (N_4183,In_1078,In_531);
xor U4184 (N_4184,In_502,In_4);
nand U4185 (N_4185,In_962,In_1616);
xor U4186 (N_4186,In_1866,In_1100);
and U4187 (N_4187,In_40,In_1342);
xnor U4188 (N_4188,In_584,In_1802);
nand U4189 (N_4189,In_1228,In_706);
and U4190 (N_4190,In_861,In_706);
xnor U4191 (N_4191,In_1719,In_868);
and U4192 (N_4192,In_1577,In_986);
or U4193 (N_4193,In_1204,In_1815);
nor U4194 (N_4194,In_578,In_713);
nand U4195 (N_4195,In_1659,In_1458);
xor U4196 (N_4196,In_674,In_336);
and U4197 (N_4197,In_434,In_1056);
nand U4198 (N_4198,In_1040,In_274);
or U4199 (N_4199,In_250,In_822);
xnor U4200 (N_4200,In_50,In_574);
nand U4201 (N_4201,In_1229,In_442);
nand U4202 (N_4202,In_395,In_879);
nor U4203 (N_4203,In_809,In_940);
nand U4204 (N_4204,In_1491,In_143);
and U4205 (N_4205,In_1723,In_925);
or U4206 (N_4206,In_1567,In_596);
nor U4207 (N_4207,In_723,In_1297);
xnor U4208 (N_4208,In_1109,In_776);
nand U4209 (N_4209,In_1267,In_1269);
or U4210 (N_4210,In_1573,In_809);
nor U4211 (N_4211,In_290,In_1988);
or U4212 (N_4212,In_1457,In_1475);
nand U4213 (N_4213,In_977,In_1092);
and U4214 (N_4214,In_1849,In_1379);
nor U4215 (N_4215,In_550,In_683);
xnor U4216 (N_4216,In_159,In_438);
xor U4217 (N_4217,In_43,In_1079);
and U4218 (N_4218,In_702,In_427);
nor U4219 (N_4219,In_299,In_1674);
nand U4220 (N_4220,In_1752,In_1431);
or U4221 (N_4221,In_228,In_760);
xnor U4222 (N_4222,In_1919,In_164);
xor U4223 (N_4223,In_836,In_1199);
nor U4224 (N_4224,In_828,In_1645);
nor U4225 (N_4225,In_625,In_1503);
nand U4226 (N_4226,In_1629,In_1472);
nor U4227 (N_4227,In_1871,In_1818);
or U4228 (N_4228,In_1380,In_537);
or U4229 (N_4229,In_1014,In_1701);
nor U4230 (N_4230,In_1428,In_1302);
and U4231 (N_4231,In_630,In_1796);
nor U4232 (N_4232,In_75,In_890);
xor U4233 (N_4233,In_1216,In_1289);
or U4234 (N_4234,In_892,In_1937);
xor U4235 (N_4235,In_72,In_210);
and U4236 (N_4236,In_499,In_1766);
and U4237 (N_4237,In_114,In_1174);
or U4238 (N_4238,In_564,In_472);
xor U4239 (N_4239,In_436,In_1676);
xnor U4240 (N_4240,In_1898,In_981);
xor U4241 (N_4241,In_1522,In_1136);
or U4242 (N_4242,In_1241,In_343);
nor U4243 (N_4243,In_194,In_612);
or U4244 (N_4244,In_868,In_1738);
nand U4245 (N_4245,In_259,In_197);
and U4246 (N_4246,In_878,In_860);
and U4247 (N_4247,In_635,In_791);
and U4248 (N_4248,In_1729,In_675);
nor U4249 (N_4249,In_1457,In_768);
or U4250 (N_4250,In_515,In_1943);
and U4251 (N_4251,In_1385,In_414);
or U4252 (N_4252,In_486,In_676);
or U4253 (N_4253,In_583,In_13);
and U4254 (N_4254,In_131,In_972);
nor U4255 (N_4255,In_1548,In_1979);
or U4256 (N_4256,In_556,In_56);
xnor U4257 (N_4257,In_606,In_1546);
nor U4258 (N_4258,In_186,In_907);
xor U4259 (N_4259,In_222,In_147);
nand U4260 (N_4260,In_442,In_1942);
and U4261 (N_4261,In_442,In_769);
or U4262 (N_4262,In_1609,In_782);
or U4263 (N_4263,In_1654,In_209);
xnor U4264 (N_4264,In_641,In_943);
xnor U4265 (N_4265,In_1525,In_669);
nor U4266 (N_4266,In_1390,In_53);
or U4267 (N_4267,In_1279,In_1502);
nand U4268 (N_4268,In_1224,In_1326);
xor U4269 (N_4269,In_984,In_823);
nand U4270 (N_4270,In_166,In_1148);
nand U4271 (N_4271,In_1333,In_1669);
and U4272 (N_4272,In_993,In_421);
xor U4273 (N_4273,In_1783,In_721);
and U4274 (N_4274,In_1111,In_1434);
nor U4275 (N_4275,In_159,In_496);
and U4276 (N_4276,In_1552,In_577);
xor U4277 (N_4277,In_1124,In_140);
nand U4278 (N_4278,In_867,In_1035);
xnor U4279 (N_4279,In_1514,In_1818);
nand U4280 (N_4280,In_1916,In_1018);
or U4281 (N_4281,In_1313,In_1647);
and U4282 (N_4282,In_190,In_1839);
and U4283 (N_4283,In_415,In_984);
nand U4284 (N_4284,In_1771,In_1811);
xnor U4285 (N_4285,In_988,In_1739);
nand U4286 (N_4286,In_1347,In_472);
or U4287 (N_4287,In_1689,In_349);
nand U4288 (N_4288,In_1053,In_1283);
or U4289 (N_4289,In_259,In_1192);
xnor U4290 (N_4290,In_1462,In_40);
nand U4291 (N_4291,In_827,In_127);
xnor U4292 (N_4292,In_1571,In_1642);
or U4293 (N_4293,In_1578,In_1078);
and U4294 (N_4294,In_606,In_1498);
xnor U4295 (N_4295,In_1953,In_1272);
xor U4296 (N_4296,In_552,In_1200);
nand U4297 (N_4297,In_207,In_1477);
xor U4298 (N_4298,In_1144,In_273);
and U4299 (N_4299,In_699,In_1927);
nor U4300 (N_4300,In_1154,In_371);
xnor U4301 (N_4301,In_91,In_1644);
or U4302 (N_4302,In_754,In_4);
nand U4303 (N_4303,In_1349,In_1318);
nand U4304 (N_4304,In_1509,In_846);
nor U4305 (N_4305,In_747,In_175);
xnor U4306 (N_4306,In_1333,In_912);
xor U4307 (N_4307,In_1269,In_1961);
xor U4308 (N_4308,In_1521,In_1787);
or U4309 (N_4309,In_1505,In_1921);
nor U4310 (N_4310,In_1005,In_842);
and U4311 (N_4311,In_1057,In_1421);
and U4312 (N_4312,In_687,In_1893);
nand U4313 (N_4313,In_581,In_545);
nand U4314 (N_4314,In_1392,In_1000);
nand U4315 (N_4315,In_1046,In_1012);
and U4316 (N_4316,In_473,In_1672);
and U4317 (N_4317,In_502,In_531);
and U4318 (N_4318,In_680,In_1719);
nor U4319 (N_4319,In_371,In_746);
or U4320 (N_4320,In_1591,In_904);
or U4321 (N_4321,In_1529,In_1033);
xnor U4322 (N_4322,In_905,In_1567);
and U4323 (N_4323,In_751,In_1721);
nor U4324 (N_4324,In_941,In_1504);
nor U4325 (N_4325,In_426,In_1391);
xor U4326 (N_4326,In_1357,In_1463);
or U4327 (N_4327,In_1884,In_528);
or U4328 (N_4328,In_628,In_1385);
or U4329 (N_4329,In_1510,In_382);
nor U4330 (N_4330,In_1447,In_271);
nand U4331 (N_4331,In_109,In_115);
xnor U4332 (N_4332,In_1615,In_653);
nand U4333 (N_4333,In_603,In_1758);
nor U4334 (N_4334,In_1261,In_1498);
or U4335 (N_4335,In_1960,In_478);
nor U4336 (N_4336,In_1418,In_1476);
nor U4337 (N_4337,In_838,In_703);
or U4338 (N_4338,In_1921,In_521);
nand U4339 (N_4339,In_320,In_1716);
or U4340 (N_4340,In_917,In_1493);
xnor U4341 (N_4341,In_1209,In_214);
nor U4342 (N_4342,In_85,In_910);
xor U4343 (N_4343,In_1506,In_343);
or U4344 (N_4344,In_1777,In_812);
and U4345 (N_4345,In_753,In_442);
xnor U4346 (N_4346,In_1833,In_374);
xor U4347 (N_4347,In_1455,In_583);
nor U4348 (N_4348,In_1879,In_311);
and U4349 (N_4349,In_1118,In_1732);
nor U4350 (N_4350,In_1463,In_1845);
xnor U4351 (N_4351,In_1314,In_1144);
or U4352 (N_4352,In_1116,In_1613);
nor U4353 (N_4353,In_311,In_1070);
nor U4354 (N_4354,In_37,In_423);
nor U4355 (N_4355,In_101,In_608);
or U4356 (N_4356,In_1190,In_485);
xor U4357 (N_4357,In_1706,In_1777);
or U4358 (N_4358,In_865,In_727);
and U4359 (N_4359,In_1221,In_1053);
xor U4360 (N_4360,In_1179,In_1261);
xnor U4361 (N_4361,In_839,In_935);
nor U4362 (N_4362,In_1042,In_618);
and U4363 (N_4363,In_11,In_611);
xnor U4364 (N_4364,In_877,In_1650);
and U4365 (N_4365,In_390,In_729);
nor U4366 (N_4366,In_1535,In_1510);
and U4367 (N_4367,In_949,In_1678);
nor U4368 (N_4368,In_1116,In_1288);
nand U4369 (N_4369,In_504,In_635);
nor U4370 (N_4370,In_62,In_1662);
xnor U4371 (N_4371,In_1076,In_929);
nor U4372 (N_4372,In_284,In_783);
nand U4373 (N_4373,In_1613,In_918);
or U4374 (N_4374,In_1976,In_972);
nand U4375 (N_4375,In_1495,In_1710);
nand U4376 (N_4376,In_1169,In_1416);
nor U4377 (N_4377,In_1386,In_1100);
nand U4378 (N_4378,In_510,In_730);
and U4379 (N_4379,In_133,In_455);
nand U4380 (N_4380,In_1623,In_828);
xnor U4381 (N_4381,In_1941,In_1111);
nor U4382 (N_4382,In_618,In_1358);
or U4383 (N_4383,In_1462,In_78);
or U4384 (N_4384,In_1180,In_1077);
nor U4385 (N_4385,In_1917,In_218);
nand U4386 (N_4386,In_562,In_1399);
nor U4387 (N_4387,In_1744,In_860);
or U4388 (N_4388,In_400,In_1070);
xor U4389 (N_4389,In_617,In_151);
nor U4390 (N_4390,In_155,In_1664);
nand U4391 (N_4391,In_1242,In_875);
or U4392 (N_4392,In_355,In_465);
nor U4393 (N_4393,In_1005,In_1399);
nand U4394 (N_4394,In_602,In_728);
and U4395 (N_4395,In_1385,In_1729);
nor U4396 (N_4396,In_1712,In_719);
nand U4397 (N_4397,In_1820,In_493);
and U4398 (N_4398,In_731,In_1923);
nor U4399 (N_4399,In_560,In_995);
xnor U4400 (N_4400,In_397,In_1226);
nor U4401 (N_4401,In_1868,In_1773);
and U4402 (N_4402,In_218,In_711);
nand U4403 (N_4403,In_208,In_375);
nand U4404 (N_4404,In_997,In_1579);
or U4405 (N_4405,In_1068,In_568);
nor U4406 (N_4406,In_718,In_1355);
or U4407 (N_4407,In_1083,In_856);
xnor U4408 (N_4408,In_306,In_1790);
or U4409 (N_4409,In_1510,In_966);
or U4410 (N_4410,In_808,In_1387);
or U4411 (N_4411,In_1962,In_523);
and U4412 (N_4412,In_103,In_509);
and U4413 (N_4413,In_286,In_1650);
nand U4414 (N_4414,In_1637,In_1024);
nor U4415 (N_4415,In_1900,In_214);
or U4416 (N_4416,In_737,In_1072);
or U4417 (N_4417,In_1479,In_1493);
xnor U4418 (N_4418,In_1334,In_522);
nor U4419 (N_4419,In_914,In_1684);
xor U4420 (N_4420,In_23,In_1058);
nand U4421 (N_4421,In_565,In_1544);
nand U4422 (N_4422,In_1221,In_1450);
and U4423 (N_4423,In_1311,In_1945);
nor U4424 (N_4424,In_348,In_1754);
nor U4425 (N_4425,In_111,In_1835);
nor U4426 (N_4426,In_1736,In_878);
or U4427 (N_4427,In_59,In_782);
nor U4428 (N_4428,In_984,In_1405);
or U4429 (N_4429,In_976,In_112);
or U4430 (N_4430,In_1444,In_1569);
or U4431 (N_4431,In_1386,In_649);
nand U4432 (N_4432,In_1327,In_554);
nor U4433 (N_4433,In_1592,In_565);
or U4434 (N_4434,In_1254,In_1883);
nand U4435 (N_4435,In_1176,In_1475);
or U4436 (N_4436,In_392,In_1266);
and U4437 (N_4437,In_542,In_1093);
nand U4438 (N_4438,In_634,In_1699);
nor U4439 (N_4439,In_1482,In_1016);
nor U4440 (N_4440,In_1446,In_1058);
nor U4441 (N_4441,In_982,In_30);
nand U4442 (N_4442,In_71,In_1093);
nand U4443 (N_4443,In_121,In_1659);
or U4444 (N_4444,In_1634,In_774);
and U4445 (N_4445,In_1713,In_372);
and U4446 (N_4446,In_386,In_437);
nor U4447 (N_4447,In_1961,In_1435);
nand U4448 (N_4448,In_365,In_464);
nand U4449 (N_4449,In_687,In_1501);
nand U4450 (N_4450,In_985,In_1065);
and U4451 (N_4451,In_380,In_712);
and U4452 (N_4452,In_1918,In_614);
or U4453 (N_4453,In_408,In_765);
and U4454 (N_4454,In_767,In_527);
nor U4455 (N_4455,In_631,In_598);
nor U4456 (N_4456,In_1167,In_1332);
xor U4457 (N_4457,In_989,In_706);
and U4458 (N_4458,In_1758,In_829);
or U4459 (N_4459,In_194,In_1164);
or U4460 (N_4460,In_1017,In_1227);
xnor U4461 (N_4461,In_1719,In_1204);
nand U4462 (N_4462,In_996,In_1651);
and U4463 (N_4463,In_936,In_1168);
or U4464 (N_4464,In_932,In_756);
nand U4465 (N_4465,In_923,In_2);
and U4466 (N_4466,In_785,In_1988);
xor U4467 (N_4467,In_1393,In_126);
nand U4468 (N_4468,In_1811,In_1801);
nand U4469 (N_4469,In_743,In_1511);
nor U4470 (N_4470,In_1472,In_267);
nand U4471 (N_4471,In_1173,In_870);
or U4472 (N_4472,In_695,In_978);
nand U4473 (N_4473,In_1918,In_1957);
nor U4474 (N_4474,In_1595,In_857);
nand U4475 (N_4475,In_926,In_1596);
xnor U4476 (N_4476,In_933,In_1332);
xnor U4477 (N_4477,In_1076,In_1398);
xnor U4478 (N_4478,In_957,In_869);
nor U4479 (N_4479,In_1432,In_1003);
nand U4480 (N_4480,In_1340,In_193);
or U4481 (N_4481,In_270,In_277);
xnor U4482 (N_4482,In_1286,In_139);
xor U4483 (N_4483,In_49,In_1273);
xor U4484 (N_4484,In_658,In_796);
nor U4485 (N_4485,In_1867,In_452);
and U4486 (N_4486,In_135,In_1344);
xnor U4487 (N_4487,In_1463,In_822);
or U4488 (N_4488,In_1582,In_1373);
or U4489 (N_4489,In_377,In_1180);
or U4490 (N_4490,In_1713,In_792);
and U4491 (N_4491,In_742,In_564);
and U4492 (N_4492,In_161,In_1875);
and U4493 (N_4493,In_811,In_38);
and U4494 (N_4494,In_1709,In_628);
nand U4495 (N_4495,In_1827,In_1013);
nand U4496 (N_4496,In_1873,In_1827);
or U4497 (N_4497,In_1523,In_1584);
xor U4498 (N_4498,In_50,In_3);
xnor U4499 (N_4499,In_1399,In_1879);
nor U4500 (N_4500,In_253,In_137);
nand U4501 (N_4501,In_993,In_1946);
xnor U4502 (N_4502,In_1018,In_26);
nor U4503 (N_4503,In_706,In_584);
nand U4504 (N_4504,In_906,In_308);
nor U4505 (N_4505,In_608,In_833);
and U4506 (N_4506,In_1941,In_1538);
nor U4507 (N_4507,In_45,In_1467);
and U4508 (N_4508,In_17,In_1803);
nand U4509 (N_4509,In_1858,In_1454);
nand U4510 (N_4510,In_1373,In_326);
or U4511 (N_4511,In_617,In_298);
nand U4512 (N_4512,In_1705,In_1025);
xor U4513 (N_4513,In_299,In_1293);
or U4514 (N_4514,In_1557,In_455);
nand U4515 (N_4515,In_1914,In_1474);
or U4516 (N_4516,In_1074,In_179);
and U4517 (N_4517,In_1472,In_88);
or U4518 (N_4518,In_1761,In_1285);
or U4519 (N_4519,In_903,In_1967);
and U4520 (N_4520,In_1686,In_1259);
nand U4521 (N_4521,In_20,In_1572);
xor U4522 (N_4522,In_851,In_485);
xor U4523 (N_4523,In_247,In_1840);
nand U4524 (N_4524,In_843,In_1181);
or U4525 (N_4525,In_998,In_433);
nor U4526 (N_4526,In_7,In_1903);
nand U4527 (N_4527,In_73,In_1742);
or U4528 (N_4528,In_1940,In_1265);
nor U4529 (N_4529,In_1693,In_962);
and U4530 (N_4530,In_143,In_1931);
or U4531 (N_4531,In_1754,In_871);
and U4532 (N_4532,In_1727,In_1692);
nand U4533 (N_4533,In_398,In_177);
and U4534 (N_4534,In_432,In_659);
nor U4535 (N_4535,In_1035,In_515);
xor U4536 (N_4536,In_1658,In_1445);
and U4537 (N_4537,In_1523,In_824);
nand U4538 (N_4538,In_182,In_1568);
nor U4539 (N_4539,In_309,In_1140);
xnor U4540 (N_4540,In_1030,In_1384);
or U4541 (N_4541,In_789,In_198);
xor U4542 (N_4542,In_1559,In_235);
or U4543 (N_4543,In_816,In_1921);
nand U4544 (N_4544,In_15,In_1095);
or U4545 (N_4545,In_1986,In_952);
xor U4546 (N_4546,In_1099,In_158);
and U4547 (N_4547,In_719,In_118);
nand U4548 (N_4548,In_1007,In_518);
or U4549 (N_4549,In_1263,In_818);
and U4550 (N_4550,In_1855,In_977);
and U4551 (N_4551,In_52,In_692);
or U4552 (N_4552,In_1034,In_539);
xor U4553 (N_4553,In_402,In_359);
and U4554 (N_4554,In_1419,In_1247);
and U4555 (N_4555,In_1853,In_570);
and U4556 (N_4556,In_655,In_965);
and U4557 (N_4557,In_302,In_346);
or U4558 (N_4558,In_1578,In_1267);
and U4559 (N_4559,In_396,In_1292);
or U4560 (N_4560,In_427,In_893);
nand U4561 (N_4561,In_729,In_1654);
nand U4562 (N_4562,In_642,In_72);
nand U4563 (N_4563,In_1210,In_1908);
and U4564 (N_4564,In_330,In_126);
xor U4565 (N_4565,In_1019,In_120);
or U4566 (N_4566,In_1901,In_1784);
nand U4567 (N_4567,In_927,In_10);
xnor U4568 (N_4568,In_736,In_190);
nor U4569 (N_4569,In_1436,In_422);
or U4570 (N_4570,In_1836,In_1051);
nand U4571 (N_4571,In_1198,In_1931);
xnor U4572 (N_4572,In_122,In_212);
xnor U4573 (N_4573,In_1375,In_1433);
nand U4574 (N_4574,In_1210,In_1474);
nor U4575 (N_4575,In_1579,In_465);
nor U4576 (N_4576,In_1633,In_1041);
xor U4577 (N_4577,In_1673,In_501);
xor U4578 (N_4578,In_1423,In_934);
nand U4579 (N_4579,In_151,In_791);
xnor U4580 (N_4580,In_1166,In_1958);
or U4581 (N_4581,In_962,In_1810);
nand U4582 (N_4582,In_396,In_703);
and U4583 (N_4583,In_1674,In_1444);
xnor U4584 (N_4584,In_49,In_1230);
xnor U4585 (N_4585,In_159,In_1244);
nor U4586 (N_4586,In_824,In_1453);
nand U4587 (N_4587,In_1169,In_1891);
nand U4588 (N_4588,In_362,In_502);
xor U4589 (N_4589,In_539,In_1400);
or U4590 (N_4590,In_1318,In_284);
or U4591 (N_4591,In_123,In_1909);
xor U4592 (N_4592,In_130,In_1697);
xor U4593 (N_4593,In_1577,In_976);
nor U4594 (N_4594,In_1635,In_591);
or U4595 (N_4595,In_1094,In_1460);
nand U4596 (N_4596,In_1368,In_242);
nor U4597 (N_4597,In_1910,In_514);
or U4598 (N_4598,In_119,In_141);
nand U4599 (N_4599,In_1117,In_949);
nor U4600 (N_4600,In_1557,In_1926);
and U4601 (N_4601,In_1215,In_1895);
nor U4602 (N_4602,In_819,In_66);
or U4603 (N_4603,In_1205,In_1954);
xor U4604 (N_4604,In_446,In_587);
and U4605 (N_4605,In_1634,In_1783);
or U4606 (N_4606,In_1298,In_1303);
and U4607 (N_4607,In_712,In_1096);
nor U4608 (N_4608,In_1105,In_1074);
xnor U4609 (N_4609,In_56,In_749);
nor U4610 (N_4610,In_1307,In_392);
or U4611 (N_4611,In_455,In_166);
and U4612 (N_4612,In_1917,In_597);
and U4613 (N_4613,In_340,In_1452);
or U4614 (N_4614,In_1347,In_923);
and U4615 (N_4615,In_1415,In_1570);
and U4616 (N_4616,In_817,In_255);
and U4617 (N_4617,In_61,In_1527);
nand U4618 (N_4618,In_237,In_1704);
or U4619 (N_4619,In_1692,In_1749);
nand U4620 (N_4620,In_17,In_742);
nor U4621 (N_4621,In_1585,In_1242);
or U4622 (N_4622,In_276,In_168);
or U4623 (N_4623,In_1727,In_1256);
xnor U4624 (N_4624,In_638,In_115);
xor U4625 (N_4625,In_1818,In_1918);
or U4626 (N_4626,In_1492,In_393);
and U4627 (N_4627,In_1503,In_1398);
nand U4628 (N_4628,In_1958,In_380);
and U4629 (N_4629,In_1850,In_761);
or U4630 (N_4630,In_1125,In_1271);
nand U4631 (N_4631,In_1072,In_1043);
and U4632 (N_4632,In_894,In_1098);
or U4633 (N_4633,In_869,In_1587);
xnor U4634 (N_4634,In_1982,In_1416);
nor U4635 (N_4635,In_285,In_1635);
xor U4636 (N_4636,In_57,In_1284);
or U4637 (N_4637,In_134,In_1317);
and U4638 (N_4638,In_624,In_1619);
or U4639 (N_4639,In_1231,In_334);
nor U4640 (N_4640,In_1054,In_1573);
xnor U4641 (N_4641,In_1674,In_974);
or U4642 (N_4642,In_891,In_1113);
and U4643 (N_4643,In_1301,In_1211);
nor U4644 (N_4644,In_404,In_983);
nand U4645 (N_4645,In_28,In_1718);
or U4646 (N_4646,In_992,In_484);
nor U4647 (N_4647,In_272,In_1427);
nand U4648 (N_4648,In_1785,In_103);
xor U4649 (N_4649,In_1343,In_1598);
or U4650 (N_4650,In_288,In_81);
xor U4651 (N_4651,In_1339,In_453);
nor U4652 (N_4652,In_892,In_1529);
nor U4653 (N_4653,In_1951,In_1243);
nand U4654 (N_4654,In_1688,In_1130);
nand U4655 (N_4655,In_1424,In_349);
and U4656 (N_4656,In_601,In_159);
and U4657 (N_4657,In_1229,In_415);
nand U4658 (N_4658,In_112,In_1631);
and U4659 (N_4659,In_361,In_1168);
xnor U4660 (N_4660,In_959,In_1917);
and U4661 (N_4661,In_614,In_1374);
and U4662 (N_4662,In_56,In_870);
and U4663 (N_4663,In_1542,In_1540);
xor U4664 (N_4664,In_783,In_228);
and U4665 (N_4665,In_1415,In_1805);
nand U4666 (N_4666,In_1750,In_1406);
and U4667 (N_4667,In_1826,In_1924);
nor U4668 (N_4668,In_1033,In_440);
xnor U4669 (N_4669,In_1846,In_1446);
xor U4670 (N_4670,In_11,In_180);
and U4671 (N_4671,In_1783,In_691);
nor U4672 (N_4672,In_1658,In_1346);
and U4673 (N_4673,In_1765,In_1841);
nor U4674 (N_4674,In_885,In_736);
or U4675 (N_4675,In_849,In_296);
nand U4676 (N_4676,In_1630,In_46);
xor U4677 (N_4677,In_1758,In_1897);
nor U4678 (N_4678,In_1064,In_791);
or U4679 (N_4679,In_916,In_930);
nand U4680 (N_4680,In_52,In_950);
nand U4681 (N_4681,In_409,In_1360);
xor U4682 (N_4682,In_297,In_1122);
or U4683 (N_4683,In_1005,In_1206);
nor U4684 (N_4684,In_1775,In_1521);
or U4685 (N_4685,In_193,In_1481);
or U4686 (N_4686,In_1889,In_800);
xor U4687 (N_4687,In_1583,In_1681);
xor U4688 (N_4688,In_1128,In_1781);
and U4689 (N_4689,In_1965,In_699);
and U4690 (N_4690,In_1748,In_897);
xnor U4691 (N_4691,In_60,In_972);
nor U4692 (N_4692,In_1587,In_192);
xor U4693 (N_4693,In_210,In_1593);
or U4694 (N_4694,In_334,In_89);
nor U4695 (N_4695,In_934,In_1664);
nor U4696 (N_4696,In_1904,In_1305);
or U4697 (N_4697,In_1332,In_1550);
nand U4698 (N_4698,In_1475,In_1979);
or U4699 (N_4699,In_1930,In_1216);
nor U4700 (N_4700,In_1855,In_1482);
or U4701 (N_4701,In_684,In_603);
nand U4702 (N_4702,In_1897,In_1652);
xor U4703 (N_4703,In_367,In_1111);
nand U4704 (N_4704,In_1434,In_1763);
nor U4705 (N_4705,In_1845,In_1510);
or U4706 (N_4706,In_1402,In_952);
nand U4707 (N_4707,In_54,In_1240);
or U4708 (N_4708,In_1158,In_866);
and U4709 (N_4709,In_1774,In_1893);
xnor U4710 (N_4710,In_1597,In_1655);
nand U4711 (N_4711,In_81,In_1311);
or U4712 (N_4712,In_1838,In_1655);
nor U4713 (N_4713,In_342,In_1952);
xnor U4714 (N_4714,In_966,In_1542);
nand U4715 (N_4715,In_238,In_572);
or U4716 (N_4716,In_1179,In_958);
or U4717 (N_4717,In_1192,In_321);
or U4718 (N_4718,In_131,In_1395);
nor U4719 (N_4719,In_285,In_1458);
nor U4720 (N_4720,In_173,In_14);
nand U4721 (N_4721,In_1502,In_1528);
xnor U4722 (N_4722,In_1154,In_541);
or U4723 (N_4723,In_383,In_1820);
xnor U4724 (N_4724,In_965,In_11);
or U4725 (N_4725,In_1562,In_1409);
and U4726 (N_4726,In_1167,In_1578);
nor U4727 (N_4727,In_228,In_773);
and U4728 (N_4728,In_206,In_1614);
xnor U4729 (N_4729,In_1023,In_254);
or U4730 (N_4730,In_1543,In_1628);
and U4731 (N_4731,In_504,In_1764);
nor U4732 (N_4732,In_1996,In_142);
nor U4733 (N_4733,In_451,In_1702);
nand U4734 (N_4734,In_1333,In_259);
nand U4735 (N_4735,In_1472,In_1535);
nor U4736 (N_4736,In_98,In_640);
xnor U4737 (N_4737,In_292,In_1308);
and U4738 (N_4738,In_1169,In_1121);
or U4739 (N_4739,In_1062,In_925);
xor U4740 (N_4740,In_1705,In_429);
nand U4741 (N_4741,In_1543,In_545);
and U4742 (N_4742,In_1817,In_1855);
xnor U4743 (N_4743,In_1720,In_1729);
or U4744 (N_4744,In_1935,In_474);
xnor U4745 (N_4745,In_1566,In_541);
or U4746 (N_4746,In_1279,In_865);
or U4747 (N_4747,In_482,In_449);
xor U4748 (N_4748,In_1723,In_1240);
or U4749 (N_4749,In_1643,In_760);
nand U4750 (N_4750,In_910,In_1984);
xor U4751 (N_4751,In_1046,In_441);
nand U4752 (N_4752,In_1021,In_1497);
or U4753 (N_4753,In_1748,In_1839);
and U4754 (N_4754,In_861,In_1761);
nor U4755 (N_4755,In_1626,In_74);
xnor U4756 (N_4756,In_123,In_1983);
nand U4757 (N_4757,In_431,In_1172);
and U4758 (N_4758,In_1174,In_334);
nand U4759 (N_4759,In_1178,In_1203);
nor U4760 (N_4760,In_146,In_1969);
and U4761 (N_4761,In_1855,In_643);
or U4762 (N_4762,In_1146,In_42);
xnor U4763 (N_4763,In_1257,In_127);
or U4764 (N_4764,In_1125,In_1896);
xor U4765 (N_4765,In_190,In_693);
nand U4766 (N_4766,In_1341,In_1988);
xor U4767 (N_4767,In_472,In_532);
xor U4768 (N_4768,In_473,In_743);
nor U4769 (N_4769,In_1163,In_910);
nand U4770 (N_4770,In_424,In_345);
or U4771 (N_4771,In_771,In_1774);
xnor U4772 (N_4772,In_612,In_1343);
nand U4773 (N_4773,In_1414,In_1568);
or U4774 (N_4774,In_441,In_1291);
xnor U4775 (N_4775,In_1939,In_1748);
or U4776 (N_4776,In_1437,In_555);
xnor U4777 (N_4777,In_949,In_1884);
or U4778 (N_4778,In_1947,In_1925);
or U4779 (N_4779,In_1524,In_405);
nand U4780 (N_4780,In_1867,In_1028);
nand U4781 (N_4781,In_1023,In_1324);
nor U4782 (N_4782,In_1995,In_778);
or U4783 (N_4783,In_141,In_1956);
nor U4784 (N_4784,In_395,In_1832);
nand U4785 (N_4785,In_1105,In_1325);
or U4786 (N_4786,In_401,In_677);
nand U4787 (N_4787,In_1422,In_1789);
and U4788 (N_4788,In_670,In_1493);
xnor U4789 (N_4789,In_567,In_227);
nor U4790 (N_4790,In_1814,In_1396);
nand U4791 (N_4791,In_525,In_649);
and U4792 (N_4792,In_875,In_242);
and U4793 (N_4793,In_1362,In_999);
xor U4794 (N_4794,In_1739,In_742);
nor U4795 (N_4795,In_1223,In_1912);
xnor U4796 (N_4796,In_230,In_1200);
nand U4797 (N_4797,In_1957,In_570);
nor U4798 (N_4798,In_282,In_145);
xor U4799 (N_4799,In_1178,In_590);
and U4800 (N_4800,In_1716,In_340);
nand U4801 (N_4801,In_1862,In_463);
xor U4802 (N_4802,In_714,In_760);
and U4803 (N_4803,In_1281,In_968);
and U4804 (N_4804,In_1451,In_1490);
or U4805 (N_4805,In_1066,In_5);
and U4806 (N_4806,In_1974,In_1545);
nor U4807 (N_4807,In_1263,In_783);
and U4808 (N_4808,In_1817,In_1901);
xnor U4809 (N_4809,In_1130,In_1309);
xor U4810 (N_4810,In_40,In_162);
xor U4811 (N_4811,In_1954,In_646);
and U4812 (N_4812,In_17,In_1523);
nor U4813 (N_4813,In_72,In_1166);
xnor U4814 (N_4814,In_1169,In_1717);
nor U4815 (N_4815,In_1529,In_658);
and U4816 (N_4816,In_10,In_1352);
or U4817 (N_4817,In_567,In_1084);
and U4818 (N_4818,In_1761,In_1802);
nor U4819 (N_4819,In_763,In_808);
or U4820 (N_4820,In_309,In_466);
or U4821 (N_4821,In_1935,In_1794);
nand U4822 (N_4822,In_661,In_1491);
and U4823 (N_4823,In_1607,In_932);
and U4824 (N_4824,In_749,In_1218);
xor U4825 (N_4825,In_1564,In_1321);
and U4826 (N_4826,In_1677,In_1786);
and U4827 (N_4827,In_1,In_195);
nor U4828 (N_4828,In_1672,In_75);
nor U4829 (N_4829,In_991,In_1079);
nand U4830 (N_4830,In_1133,In_1709);
nor U4831 (N_4831,In_90,In_471);
xnor U4832 (N_4832,In_797,In_862);
or U4833 (N_4833,In_1322,In_73);
nor U4834 (N_4834,In_47,In_1499);
xor U4835 (N_4835,In_1040,In_745);
nor U4836 (N_4836,In_487,In_325);
or U4837 (N_4837,In_406,In_1057);
and U4838 (N_4838,In_1364,In_755);
nand U4839 (N_4839,In_1623,In_947);
xor U4840 (N_4840,In_1540,In_1256);
and U4841 (N_4841,In_1822,In_1437);
nor U4842 (N_4842,In_176,In_908);
nand U4843 (N_4843,In_1365,In_1383);
and U4844 (N_4844,In_1302,In_1250);
or U4845 (N_4845,In_747,In_1107);
and U4846 (N_4846,In_551,In_1863);
xnor U4847 (N_4847,In_1149,In_587);
and U4848 (N_4848,In_1163,In_549);
nand U4849 (N_4849,In_481,In_853);
and U4850 (N_4850,In_1938,In_1044);
nand U4851 (N_4851,In_541,In_53);
or U4852 (N_4852,In_1021,In_506);
or U4853 (N_4853,In_802,In_223);
and U4854 (N_4854,In_933,In_841);
nor U4855 (N_4855,In_97,In_132);
and U4856 (N_4856,In_769,In_1770);
nand U4857 (N_4857,In_1439,In_842);
nor U4858 (N_4858,In_246,In_370);
nand U4859 (N_4859,In_748,In_1753);
nor U4860 (N_4860,In_841,In_1292);
nand U4861 (N_4861,In_541,In_1440);
or U4862 (N_4862,In_447,In_1407);
xnor U4863 (N_4863,In_1024,In_1154);
nand U4864 (N_4864,In_320,In_1538);
nand U4865 (N_4865,In_595,In_999);
nor U4866 (N_4866,In_245,In_1488);
and U4867 (N_4867,In_1426,In_818);
or U4868 (N_4868,In_1253,In_1313);
xor U4869 (N_4869,In_101,In_118);
or U4870 (N_4870,In_948,In_873);
and U4871 (N_4871,In_1126,In_1691);
and U4872 (N_4872,In_1879,In_296);
and U4873 (N_4873,In_65,In_66);
nand U4874 (N_4874,In_1462,In_851);
nand U4875 (N_4875,In_883,In_1843);
xnor U4876 (N_4876,In_598,In_830);
nand U4877 (N_4877,In_126,In_1327);
and U4878 (N_4878,In_1497,In_989);
xnor U4879 (N_4879,In_698,In_1923);
nand U4880 (N_4880,In_1822,In_224);
nor U4881 (N_4881,In_1753,In_1234);
nor U4882 (N_4882,In_1519,In_1532);
or U4883 (N_4883,In_1749,In_695);
nand U4884 (N_4884,In_1062,In_1093);
nand U4885 (N_4885,In_917,In_262);
or U4886 (N_4886,In_1910,In_718);
xnor U4887 (N_4887,In_1847,In_989);
and U4888 (N_4888,In_1638,In_1863);
nor U4889 (N_4889,In_156,In_425);
nand U4890 (N_4890,In_150,In_15);
nand U4891 (N_4891,In_503,In_857);
or U4892 (N_4892,In_40,In_1158);
or U4893 (N_4893,In_469,In_922);
and U4894 (N_4894,In_277,In_822);
and U4895 (N_4895,In_766,In_430);
nand U4896 (N_4896,In_520,In_872);
nor U4897 (N_4897,In_319,In_1522);
and U4898 (N_4898,In_1174,In_1955);
nor U4899 (N_4899,In_660,In_1100);
and U4900 (N_4900,In_1152,In_336);
nor U4901 (N_4901,In_110,In_928);
and U4902 (N_4902,In_665,In_1286);
nor U4903 (N_4903,In_1343,In_1081);
or U4904 (N_4904,In_974,In_641);
or U4905 (N_4905,In_1204,In_1604);
xnor U4906 (N_4906,In_1478,In_1620);
or U4907 (N_4907,In_1750,In_234);
xor U4908 (N_4908,In_45,In_904);
xnor U4909 (N_4909,In_1115,In_467);
and U4910 (N_4910,In_527,In_1326);
xnor U4911 (N_4911,In_1532,In_606);
nand U4912 (N_4912,In_1178,In_1821);
xor U4913 (N_4913,In_1648,In_1791);
and U4914 (N_4914,In_756,In_1345);
nand U4915 (N_4915,In_192,In_391);
nor U4916 (N_4916,In_974,In_833);
nor U4917 (N_4917,In_674,In_1704);
nor U4918 (N_4918,In_273,In_812);
nor U4919 (N_4919,In_542,In_966);
xnor U4920 (N_4920,In_1264,In_591);
xor U4921 (N_4921,In_195,In_503);
nand U4922 (N_4922,In_1712,In_432);
nand U4923 (N_4923,In_267,In_823);
and U4924 (N_4924,In_1764,In_951);
xor U4925 (N_4925,In_562,In_958);
xnor U4926 (N_4926,In_1199,In_78);
and U4927 (N_4927,In_1545,In_975);
or U4928 (N_4928,In_133,In_1294);
xor U4929 (N_4929,In_872,In_698);
or U4930 (N_4930,In_1971,In_655);
nand U4931 (N_4931,In_143,In_426);
nand U4932 (N_4932,In_873,In_1480);
nor U4933 (N_4933,In_1772,In_700);
xnor U4934 (N_4934,In_1654,In_1503);
xor U4935 (N_4935,In_1574,In_1077);
and U4936 (N_4936,In_114,In_1495);
nand U4937 (N_4937,In_1312,In_1672);
and U4938 (N_4938,In_305,In_804);
nor U4939 (N_4939,In_1947,In_205);
or U4940 (N_4940,In_1066,In_1118);
nor U4941 (N_4941,In_94,In_1332);
nor U4942 (N_4942,In_1791,In_59);
xnor U4943 (N_4943,In_396,In_459);
nor U4944 (N_4944,In_285,In_650);
xor U4945 (N_4945,In_134,In_504);
nor U4946 (N_4946,In_1000,In_620);
or U4947 (N_4947,In_936,In_996);
and U4948 (N_4948,In_1592,In_1889);
xor U4949 (N_4949,In_1699,In_1664);
xor U4950 (N_4950,In_1442,In_456);
or U4951 (N_4951,In_338,In_698);
and U4952 (N_4952,In_1537,In_235);
nor U4953 (N_4953,In_909,In_44);
and U4954 (N_4954,In_1791,In_1953);
nand U4955 (N_4955,In_237,In_698);
nand U4956 (N_4956,In_463,In_1460);
or U4957 (N_4957,In_232,In_1920);
and U4958 (N_4958,In_640,In_1995);
nand U4959 (N_4959,In_135,In_1109);
xnor U4960 (N_4960,In_1245,In_523);
nand U4961 (N_4961,In_1055,In_1222);
nor U4962 (N_4962,In_665,In_254);
nor U4963 (N_4963,In_1409,In_1823);
and U4964 (N_4964,In_1474,In_288);
xor U4965 (N_4965,In_1886,In_184);
or U4966 (N_4966,In_1581,In_1495);
and U4967 (N_4967,In_1021,In_1266);
nand U4968 (N_4968,In_557,In_716);
or U4969 (N_4969,In_1885,In_1722);
nor U4970 (N_4970,In_618,In_1050);
or U4971 (N_4971,In_604,In_1738);
nand U4972 (N_4972,In_576,In_1627);
or U4973 (N_4973,In_344,In_619);
nand U4974 (N_4974,In_544,In_31);
and U4975 (N_4975,In_881,In_1834);
nand U4976 (N_4976,In_1902,In_1345);
xor U4977 (N_4977,In_304,In_639);
and U4978 (N_4978,In_1318,In_635);
or U4979 (N_4979,In_26,In_312);
or U4980 (N_4980,In_426,In_1644);
nand U4981 (N_4981,In_1245,In_481);
and U4982 (N_4982,In_295,In_503);
or U4983 (N_4983,In_394,In_757);
or U4984 (N_4984,In_1837,In_755);
nand U4985 (N_4985,In_64,In_1666);
nor U4986 (N_4986,In_1335,In_1571);
nand U4987 (N_4987,In_476,In_860);
and U4988 (N_4988,In_1432,In_1719);
nand U4989 (N_4989,In_909,In_120);
and U4990 (N_4990,In_1706,In_1573);
and U4991 (N_4991,In_382,In_1509);
xnor U4992 (N_4992,In_1052,In_634);
and U4993 (N_4993,In_239,In_1715);
xor U4994 (N_4994,In_88,In_463);
or U4995 (N_4995,In_699,In_612);
nand U4996 (N_4996,In_370,In_1287);
or U4997 (N_4997,In_189,In_1908);
and U4998 (N_4998,In_524,In_1782);
nand U4999 (N_4999,In_1576,In_840);
nand U5000 (N_5000,N_4815,N_2989);
nand U5001 (N_5001,N_1518,N_3535);
nor U5002 (N_5002,N_821,N_3121);
and U5003 (N_5003,N_343,N_1047);
and U5004 (N_5004,N_3413,N_3617);
nand U5005 (N_5005,N_3651,N_1863);
and U5006 (N_5006,N_812,N_3742);
xor U5007 (N_5007,N_3782,N_505);
nor U5008 (N_5008,N_1666,N_242);
and U5009 (N_5009,N_3602,N_92);
nand U5010 (N_5010,N_576,N_1897);
xor U5011 (N_5011,N_1430,N_3129);
and U5012 (N_5012,N_2225,N_4655);
nand U5013 (N_5013,N_3548,N_654);
nand U5014 (N_5014,N_4706,N_4249);
nor U5015 (N_5015,N_602,N_4278);
or U5016 (N_5016,N_3492,N_2789);
nor U5017 (N_5017,N_4760,N_3331);
xnor U5018 (N_5018,N_4596,N_985);
nor U5019 (N_5019,N_2947,N_3905);
nor U5020 (N_5020,N_1218,N_1439);
and U5021 (N_5021,N_2640,N_3877);
xnor U5022 (N_5022,N_4821,N_2160);
or U5023 (N_5023,N_2595,N_856);
or U5024 (N_5024,N_52,N_3159);
and U5025 (N_5025,N_884,N_4835);
xnor U5026 (N_5026,N_969,N_4687);
and U5027 (N_5027,N_4506,N_4568);
or U5028 (N_5028,N_3537,N_2249);
nand U5029 (N_5029,N_855,N_2173);
or U5030 (N_5030,N_4657,N_2761);
or U5031 (N_5031,N_287,N_1542);
or U5032 (N_5032,N_4554,N_3780);
nor U5033 (N_5033,N_104,N_125);
nor U5034 (N_5034,N_732,N_3449);
or U5035 (N_5035,N_1348,N_2265);
and U5036 (N_5036,N_1488,N_3618);
or U5037 (N_5037,N_1973,N_2938);
or U5038 (N_5038,N_562,N_1743);
xor U5039 (N_5039,N_2479,N_1510);
xor U5040 (N_5040,N_3670,N_4961);
xor U5041 (N_5041,N_351,N_4284);
nor U5042 (N_5042,N_1061,N_3634);
or U5043 (N_5043,N_2154,N_4861);
nand U5044 (N_5044,N_500,N_3363);
xor U5045 (N_5045,N_3063,N_3244);
and U5046 (N_5046,N_21,N_862);
and U5047 (N_5047,N_4226,N_502);
and U5048 (N_5048,N_4865,N_453);
xor U5049 (N_5049,N_3606,N_249);
or U5050 (N_5050,N_582,N_2836);
nand U5051 (N_5051,N_2923,N_618);
nand U5052 (N_5052,N_1583,N_2770);
or U5053 (N_5053,N_4668,N_4597);
xor U5054 (N_5054,N_1018,N_2200);
and U5055 (N_5055,N_2385,N_2894);
nor U5056 (N_5056,N_1643,N_1117);
and U5057 (N_5057,N_544,N_3157);
xnor U5058 (N_5058,N_492,N_726);
nand U5059 (N_5059,N_1454,N_1005);
xnor U5060 (N_5060,N_1686,N_3570);
and U5061 (N_5061,N_3937,N_3946);
or U5062 (N_5062,N_3864,N_4494);
xor U5063 (N_5063,N_3242,N_366);
and U5064 (N_5064,N_2283,N_4920);
or U5065 (N_5065,N_695,N_439);
xor U5066 (N_5066,N_3303,N_2591);
xor U5067 (N_5067,N_2170,N_1924);
nand U5068 (N_5068,N_4031,N_4064);
nor U5069 (N_5069,N_1720,N_606);
or U5070 (N_5070,N_4935,N_1023);
nand U5071 (N_5071,N_956,N_1232);
nand U5072 (N_5072,N_123,N_4072);
xor U5073 (N_5073,N_4167,N_2963);
nor U5074 (N_5074,N_4156,N_3639);
nor U5075 (N_5075,N_3724,N_2686);
and U5076 (N_5076,N_3783,N_1532);
or U5077 (N_5077,N_1537,N_3404);
nand U5078 (N_5078,N_286,N_2497);
xor U5079 (N_5079,N_3172,N_4244);
nor U5080 (N_5080,N_3220,N_3723);
and U5081 (N_5081,N_3731,N_2831);
nand U5082 (N_5082,N_165,N_1648);
nor U5083 (N_5083,N_109,N_4137);
xor U5084 (N_5084,N_4140,N_3869);
nor U5085 (N_5085,N_3356,N_3156);
nand U5086 (N_5086,N_3900,N_1129);
and U5087 (N_5087,N_1441,N_2703);
nor U5088 (N_5088,N_3423,N_4091);
xor U5089 (N_5089,N_3348,N_2885);
nand U5090 (N_5090,N_1652,N_1257);
xnor U5091 (N_5091,N_4689,N_1093);
xor U5092 (N_5092,N_4897,N_4627);
or U5093 (N_5093,N_1144,N_4148);
and U5094 (N_5094,N_1298,N_570);
nor U5095 (N_5095,N_2784,N_4598);
nand U5096 (N_5096,N_1295,N_3978);
nor U5097 (N_5097,N_3674,N_2237);
or U5098 (N_5098,N_644,N_3643);
xor U5099 (N_5099,N_1269,N_1500);
xnor U5100 (N_5100,N_4536,N_1830);
and U5101 (N_5101,N_2313,N_4008);
and U5102 (N_5102,N_3901,N_2721);
xor U5103 (N_5103,N_635,N_811);
xor U5104 (N_5104,N_3005,N_1695);
nand U5105 (N_5105,N_694,N_4878);
nor U5106 (N_5106,N_3292,N_4459);
xnor U5107 (N_5107,N_4857,N_4968);
xnor U5108 (N_5108,N_4937,N_4652);
or U5109 (N_5109,N_4138,N_2544);
nand U5110 (N_5110,N_4853,N_4400);
or U5111 (N_5111,N_2169,N_4283);
nor U5112 (N_5112,N_1568,N_3216);
or U5113 (N_5113,N_871,N_1185);
xnor U5114 (N_5114,N_4600,N_4621);
or U5115 (N_5115,N_912,N_796);
xor U5116 (N_5116,N_2267,N_2391);
and U5117 (N_5117,N_3099,N_4851);
or U5118 (N_5118,N_1880,N_4161);
xnor U5119 (N_5119,N_404,N_3104);
or U5120 (N_5120,N_1688,N_3462);
or U5121 (N_5121,N_1696,N_247);
xnor U5122 (N_5122,N_2910,N_4427);
xnor U5123 (N_5123,N_2733,N_10);
nor U5124 (N_5124,N_1127,N_1501);
nor U5125 (N_5125,N_195,N_3071);
nand U5126 (N_5126,N_3977,N_406);
and U5127 (N_5127,N_4000,N_2229);
or U5128 (N_5128,N_739,N_1584);
xnor U5129 (N_5129,N_2131,N_3081);
or U5130 (N_5130,N_3231,N_2731);
nand U5131 (N_5131,N_954,N_1546);
nor U5132 (N_5132,N_1881,N_3466);
nor U5133 (N_5133,N_4368,N_1980);
or U5134 (N_5134,N_1827,N_1140);
nor U5135 (N_5135,N_4364,N_2757);
nand U5136 (N_5136,N_2227,N_2375);
xnor U5137 (N_5137,N_1256,N_895);
nor U5138 (N_5138,N_2402,N_1646);
and U5139 (N_5139,N_2769,N_3726);
xor U5140 (N_5140,N_1572,N_2900);
xnor U5141 (N_5141,N_1226,N_4240);
nor U5142 (N_5142,N_3197,N_520);
and U5143 (N_5143,N_4874,N_4288);
xor U5144 (N_5144,N_1115,N_4006);
xor U5145 (N_5145,N_3831,N_4817);
xnor U5146 (N_5146,N_1110,N_2880);
or U5147 (N_5147,N_3779,N_70);
or U5148 (N_5148,N_3525,N_20);
and U5149 (N_5149,N_4358,N_4341);
or U5150 (N_5150,N_2748,N_620);
xnor U5151 (N_5151,N_1280,N_2041);
and U5152 (N_5152,N_2157,N_672);
nor U5153 (N_5153,N_629,N_3968);
nand U5154 (N_5154,N_1623,N_1244);
or U5155 (N_5155,N_3673,N_3122);
nand U5156 (N_5156,N_4952,N_4232);
nand U5157 (N_5157,N_3253,N_133);
nor U5158 (N_5158,N_3246,N_634);
or U5159 (N_5159,N_1995,N_2744);
or U5160 (N_5160,N_710,N_4108);
or U5161 (N_5161,N_917,N_2351);
nor U5162 (N_5162,N_2483,N_4455);
nor U5163 (N_5163,N_3085,N_1889);
nand U5164 (N_5164,N_4017,N_1736);
or U5165 (N_5165,N_3571,N_4214);
nand U5166 (N_5166,N_1319,N_3507);
nor U5167 (N_5167,N_198,N_1098);
nor U5168 (N_5168,N_3550,N_2407);
nand U5169 (N_5169,N_4545,N_359);
and U5170 (N_5170,N_2725,N_3872);
nor U5171 (N_5171,N_3545,N_3421);
xor U5172 (N_5172,N_1692,N_1859);
or U5173 (N_5173,N_2631,N_3647);
or U5174 (N_5174,N_1741,N_4460);
xor U5175 (N_5175,N_4109,N_4026);
and U5176 (N_5176,N_965,N_1581);
nand U5177 (N_5177,N_1610,N_2981);
nor U5178 (N_5178,N_2023,N_34);
nor U5179 (N_5179,N_3811,N_3041);
nor U5180 (N_5180,N_1912,N_3436);
nand U5181 (N_5181,N_2768,N_2025);
or U5182 (N_5182,N_1408,N_1262);
or U5183 (N_5183,N_4508,N_4542);
and U5184 (N_5184,N_3415,N_141);
xnor U5185 (N_5185,N_2302,N_3728);
and U5186 (N_5186,N_489,N_1871);
xnor U5187 (N_5187,N_4149,N_4521);
nand U5188 (N_5188,N_2785,N_4188);
or U5189 (N_5189,N_3696,N_170);
xor U5190 (N_5190,N_2967,N_3008);
nand U5191 (N_5191,N_2969,N_1901);
nor U5192 (N_5192,N_3610,N_1003);
nand U5193 (N_5193,N_988,N_4365);
xnor U5194 (N_5194,N_1103,N_2408);
xnor U5195 (N_5195,N_3187,N_1763);
xnor U5196 (N_5196,N_1204,N_2103);
xor U5197 (N_5197,N_4942,N_4361);
xnor U5198 (N_5198,N_2798,N_932);
nor U5199 (N_5199,N_2608,N_4704);
and U5200 (N_5200,N_3391,N_2362);
or U5201 (N_5201,N_4967,N_622);
and U5202 (N_5202,N_2257,N_4089);
and U5203 (N_5203,N_4466,N_2822);
or U5204 (N_5204,N_2182,N_3684);
nand U5205 (N_5205,N_3270,N_4969);
nor U5206 (N_5206,N_2845,N_961);
and U5207 (N_5207,N_138,N_866);
xor U5208 (N_5208,N_1544,N_1953);
nand U5209 (N_5209,N_3894,N_4312);
and U5210 (N_5210,N_1687,N_3036);
nand U5211 (N_5211,N_2274,N_299);
and U5212 (N_5212,N_1788,N_2504);
nor U5213 (N_5213,N_3793,N_4281);
xnor U5214 (N_5214,N_874,N_4943);
nor U5215 (N_5215,N_2600,N_4746);
or U5216 (N_5216,N_4322,N_3441);
xor U5217 (N_5217,N_1999,N_1470);
xor U5218 (N_5218,N_3196,N_4224);
and U5219 (N_5219,N_1007,N_1528);
xnor U5220 (N_5220,N_2100,N_3543);
xnor U5221 (N_5221,N_1054,N_3629);
nand U5222 (N_5222,N_1443,N_4454);
nand U5223 (N_5223,N_2141,N_679);
nor U5224 (N_5224,N_2395,N_3454);
or U5225 (N_5225,N_3215,N_3383);
xnor U5226 (N_5226,N_590,N_4928);
or U5227 (N_5227,N_3965,N_444);
nand U5228 (N_5228,N_4362,N_2951);
or U5229 (N_5229,N_2932,N_3353);
nor U5230 (N_5230,N_3173,N_370);
nand U5231 (N_5231,N_1576,N_545);
nand U5232 (N_5232,N_1458,N_1312);
nand U5233 (N_5233,N_3201,N_4966);
nor U5234 (N_5234,N_4437,N_877);
and U5235 (N_5235,N_842,N_3710);
xor U5236 (N_5236,N_1377,N_3145);
nand U5237 (N_5237,N_3013,N_12);
xor U5238 (N_5238,N_2851,N_3457);
xor U5239 (N_5239,N_4192,N_4329);
nand U5240 (N_5240,N_805,N_4318);
or U5241 (N_5241,N_4163,N_223);
nor U5242 (N_5242,N_4005,N_3269);
nand U5243 (N_5243,N_3885,N_3746);
nor U5244 (N_5244,N_714,N_1189);
or U5245 (N_5245,N_1234,N_220);
or U5246 (N_5246,N_183,N_2069);
xnor U5247 (N_5247,N_1989,N_2081);
nand U5248 (N_5248,N_181,N_771);
nor U5249 (N_5249,N_4090,N_1251);
nor U5250 (N_5250,N_2833,N_616);
or U5251 (N_5251,N_1702,N_3918);
nand U5252 (N_5252,N_2444,N_281);
or U5253 (N_5253,N_3974,N_1163);
and U5254 (N_5254,N_897,N_3790);
nor U5255 (N_5255,N_1772,N_1245);
nor U5256 (N_5256,N_1268,N_6);
and U5257 (N_5257,N_107,N_4080);
nand U5258 (N_5258,N_3660,N_607);
nor U5259 (N_5259,N_1073,N_4674);
nand U5260 (N_5260,N_4294,N_3433);
nand U5261 (N_5261,N_4480,N_2763);
nand U5262 (N_5262,N_15,N_1357);
xnor U5263 (N_5263,N_795,N_1856);
nor U5264 (N_5264,N_128,N_3890);
and U5265 (N_5265,N_137,N_2862);
xnor U5266 (N_5266,N_848,N_1857);
xor U5267 (N_5267,N_899,N_4884);
xnor U5268 (N_5268,N_2427,N_4269);
xnor U5269 (N_5269,N_1690,N_4628);
nor U5270 (N_5270,N_2239,N_609);
nand U5271 (N_5271,N_3337,N_3450);
or U5272 (N_5272,N_1492,N_3867);
and U5273 (N_5273,N_2516,N_3359);
xor U5274 (N_5274,N_2468,N_94);
nor U5275 (N_5275,N_569,N_1013);
and U5276 (N_5276,N_1105,N_3169);
nor U5277 (N_5277,N_498,N_1814);
nor U5278 (N_5278,N_2745,N_510);
nor U5279 (N_5279,N_2209,N_1595);
nor U5280 (N_5280,N_4242,N_3054);
and U5281 (N_5281,N_2448,N_3330);
nand U5282 (N_5282,N_4429,N_2);
nor U5283 (N_5283,N_2406,N_1944);
nand U5284 (N_5284,N_39,N_2156);
nand U5285 (N_5285,N_883,N_3300);
nor U5286 (N_5286,N_3347,N_2288);
and U5287 (N_5287,N_4397,N_1959);
or U5288 (N_5288,N_927,N_797);
and U5289 (N_5289,N_1230,N_4836);
or U5290 (N_5290,N_31,N_390);
nor U5291 (N_5291,N_3791,N_3962);
nor U5292 (N_5292,N_416,N_4287);
nor U5293 (N_5293,N_3214,N_4112);
or U5294 (N_5294,N_4450,N_2827);
nor U5295 (N_5295,N_4958,N_2093);
nor U5296 (N_5296,N_4843,N_2475);
xor U5297 (N_5297,N_275,N_578);
xor U5298 (N_5298,N_911,N_4561);
nand U5299 (N_5299,N_791,N_2062);
or U5300 (N_5300,N_2092,N_1640);
nor U5301 (N_5301,N_1008,N_3392);
and U5302 (N_5302,N_3338,N_3473);
or U5303 (N_5303,N_1842,N_4557);
and U5304 (N_5304,N_506,N_4859);
and U5305 (N_5305,N_4613,N_1057);
nor U5306 (N_5306,N_1020,N_3440);
or U5307 (N_5307,N_3568,N_459);
and U5308 (N_5308,N_2122,N_2289);
or U5309 (N_5309,N_2487,N_3828);
or U5310 (N_5310,N_1472,N_3097);
and U5311 (N_5311,N_3838,N_205);
nand U5312 (N_5312,N_2113,N_1920);
xnor U5313 (N_5313,N_2604,N_3304);
nor U5314 (N_5314,N_3717,N_2645);
xor U5315 (N_5315,N_4753,N_987);
or U5316 (N_5316,N_4713,N_1258);
nor U5317 (N_5317,N_3534,N_2802);
nand U5318 (N_5318,N_2044,N_823);
or U5319 (N_5319,N_75,N_2364);
nor U5320 (N_5320,N_2664,N_1487);
and U5321 (N_5321,N_4899,N_2212);
xnor U5322 (N_5322,N_4349,N_2942);
or U5323 (N_5323,N_2056,N_2334);
nor U5324 (N_5324,N_4514,N_769);
xor U5325 (N_5325,N_1012,N_3422);
nor U5326 (N_5326,N_4441,N_4464);
and U5327 (N_5327,N_4754,N_2118);
and U5328 (N_5328,N_423,N_4303);
or U5329 (N_5329,N_331,N_3664);
nand U5330 (N_5330,N_4317,N_4366);
or U5331 (N_5331,N_588,N_2639);
nand U5332 (N_5332,N_1081,N_2979);
and U5333 (N_5333,N_4528,N_1084);
or U5334 (N_5334,N_4009,N_3829);
nand U5335 (N_5335,N_124,N_4814);
or U5336 (N_5336,N_3313,N_1207);
nor U5337 (N_5337,N_2722,N_3718);
xor U5338 (N_5338,N_231,N_1341);
or U5339 (N_5339,N_3753,N_3418);
and U5340 (N_5340,N_1867,N_446);
nor U5341 (N_5341,N_1865,N_1101);
xnor U5342 (N_5342,N_3352,N_3018);
or U5343 (N_5343,N_4592,N_3034);
or U5344 (N_5344,N_4462,N_160);
nand U5345 (N_5345,N_1118,N_554);
or U5346 (N_5346,N_2693,N_2772);
xor U5347 (N_5347,N_4707,N_1451);
nor U5348 (N_5348,N_2767,N_3556);
nor U5349 (N_5349,N_976,N_1992);
or U5350 (N_5350,N_3042,N_1352);
or U5351 (N_5351,N_2097,N_2457);
and U5352 (N_5352,N_2959,N_495);
and U5353 (N_5353,N_2756,N_1113);
and U5354 (N_5354,N_2801,N_4905);
and U5355 (N_5355,N_3306,N_2127);
or U5356 (N_5356,N_25,N_2204);
nand U5357 (N_5357,N_4549,N_835);
xor U5358 (N_5358,N_4953,N_4203);
or U5359 (N_5359,N_1321,N_2853);
nor U5360 (N_5360,N_2913,N_4539);
and U5361 (N_5361,N_2117,N_3682);
nand U5362 (N_5362,N_380,N_3049);
nor U5363 (N_5363,N_3911,N_553);
or U5364 (N_5364,N_3262,N_3594);
and U5365 (N_5365,N_2751,N_3512);
or U5366 (N_5366,N_4710,N_312);
xnor U5367 (N_5367,N_3103,N_1386);
nand U5368 (N_5368,N_3892,N_3478);
xnor U5369 (N_5369,N_4417,N_852);
and U5370 (N_5370,N_3060,N_3032);
and U5371 (N_5371,N_4096,N_1423);
and U5372 (N_5372,N_3904,N_4712);
and U5373 (N_5373,N_164,N_4914);
and U5374 (N_5374,N_4946,N_1668);
xor U5375 (N_5375,N_4190,N_2795);
and U5376 (N_5376,N_185,N_1770);
or U5377 (N_5377,N_4761,N_2336);
xnor U5378 (N_5378,N_555,N_3120);
nor U5379 (N_5379,N_2707,N_773);
or U5380 (N_5380,N_4608,N_3561);
xor U5381 (N_5381,N_4693,N_3374);
or U5382 (N_5382,N_2379,N_4559);
nand U5383 (N_5383,N_989,N_1751);
nor U5384 (N_5384,N_265,N_766);
xnor U5385 (N_5385,N_1063,N_4808);
nand U5386 (N_5386,N_3027,N_2863);
nand U5387 (N_5387,N_3860,N_2397);
and U5388 (N_5388,N_3598,N_4660);
and U5389 (N_5389,N_29,N_3690);
nor U5390 (N_5390,N_3888,N_2493);
or U5391 (N_5391,N_1965,N_2382);
nand U5392 (N_5392,N_1169,N_2984);
nand U5393 (N_5393,N_2138,N_2464);
or U5394 (N_5394,N_276,N_691);
or U5395 (N_5395,N_4635,N_960);
and U5396 (N_5396,N_4324,N_754);
nor U5397 (N_5397,N_4998,N_4744);
and U5398 (N_5398,N_3957,N_2149);
nand U5399 (N_5399,N_2201,N_2776);
nand U5400 (N_5400,N_2294,N_783);
and U5401 (N_5401,N_4419,N_4513);
and U5402 (N_5402,N_365,N_2553);
xnor U5403 (N_5403,N_4881,N_1925);
and U5404 (N_5404,N_3309,N_2803);
or U5405 (N_5405,N_2490,N_3212);
and U5406 (N_5406,N_2451,N_2857);
nor U5407 (N_5407,N_121,N_1402);
and U5408 (N_5408,N_660,N_733);
or U5409 (N_5409,N_3916,N_4565);
xor U5410 (N_5410,N_4556,N_3850);
nand U5411 (N_5411,N_674,N_3523);
or U5412 (N_5412,N_1250,N_1119);
nand U5413 (N_5413,N_3031,N_4496);
xnor U5414 (N_5414,N_2440,N_610);
nand U5415 (N_5415,N_2386,N_3991);
and U5416 (N_5416,N_707,N_838);
xor U5417 (N_5417,N_3721,N_234);
nand U5418 (N_5418,N_2996,N_1571);
nor U5419 (N_5419,N_4113,N_4023);
and U5420 (N_5420,N_2718,N_2578);
nand U5421 (N_5421,N_2569,N_631);
nor U5422 (N_5422,N_4171,N_2366);
nand U5423 (N_5423,N_2280,N_3110);
or U5424 (N_5424,N_4453,N_4423);
xnor U5425 (N_5425,N_105,N_3951);
xnor U5426 (N_5426,N_2861,N_3371);
xnor U5427 (N_5427,N_1930,N_1050);
and U5428 (N_5428,N_1214,N_2501);
xnor U5429 (N_5429,N_740,N_4728);
and U5430 (N_5430,N_3672,N_1070);
nor U5431 (N_5431,N_3952,N_2650);
or U5432 (N_5432,N_1318,N_146);
nor U5433 (N_5433,N_4833,N_3083);
nand U5434 (N_5434,N_3135,N_1582);
xor U5435 (N_5435,N_1287,N_1415);
or U5436 (N_5436,N_2758,N_4959);
nand U5437 (N_5437,N_937,N_2710);
xnor U5438 (N_5438,N_532,N_3393);
nor U5439 (N_5439,N_1124,N_549);
nand U5440 (N_5440,N_2356,N_3896);
nand U5441 (N_5441,N_1642,N_786);
and U5442 (N_5442,N_4220,N_2814);
xnor U5443 (N_5443,N_1817,N_2287);
and U5444 (N_5444,N_1588,N_2076);
or U5445 (N_5445,N_4921,N_889);
or U5446 (N_5446,N_3064,N_1832);
nand U5447 (N_5447,N_2164,N_4619);
and U5448 (N_5448,N_3140,N_3686);
xor U5449 (N_5449,N_3816,N_2343);
nor U5450 (N_5450,N_1424,N_344);
or U5451 (N_5451,N_1854,N_3198);
nor U5452 (N_5452,N_3070,N_640);
or U5453 (N_5453,N_1718,N_4566);
nand U5454 (N_5454,N_3613,N_3748);
xnor U5455 (N_5455,N_112,N_3472);
nor U5456 (N_5456,N_3572,N_967);
nand U5457 (N_5457,N_4371,N_1428);
or U5458 (N_5458,N_1270,N_3050);
or U5459 (N_5459,N_1340,N_4540);
nand U5460 (N_5460,N_4511,N_854);
or U5461 (N_5461,N_2291,N_3924);
nor U5462 (N_5462,N_1802,N_1190);
and U5463 (N_5463,N_2898,N_4088);
or U5464 (N_5464,N_1154,N_3075);
nor U5465 (N_5465,N_132,N_361);
xnor U5466 (N_5466,N_4623,N_4123);
and U5467 (N_5467,N_1206,N_1815);
nor U5468 (N_5468,N_2125,N_604);
and U5469 (N_5469,N_54,N_2316);
nor U5470 (N_5470,N_1264,N_4791);
nor U5471 (N_5471,N_4810,N_397);
nand U5472 (N_5472,N_3772,N_2482);
and U5473 (N_5473,N_3310,N_2521);
nand U5474 (N_5474,N_1028,N_2114);
and U5475 (N_5475,N_3994,N_2206);
xnor U5476 (N_5476,N_1917,N_1596);
and U5477 (N_5477,N_1067,N_4426);
nand U5478 (N_5478,N_2676,N_3597);
xor U5479 (N_5479,N_3514,N_4049);
nand U5480 (N_5480,N_3380,N_1171);
nand U5481 (N_5481,N_1782,N_1673);
nor U5482 (N_5482,N_4991,N_4263);
or U5483 (N_5483,N_3935,N_4601);
nand U5484 (N_5484,N_718,N_2263);
nand U5485 (N_5485,N_4142,N_980);
or U5486 (N_5486,N_4230,N_816);
xor U5487 (N_5487,N_2774,N_3278);
xnor U5488 (N_5488,N_197,N_3117);
and U5489 (N_5489,N_3221,N_3927);
or U5490 (N_5490,N_2931,N_3076);
xnor U5491 (N_5491,N_2186,N_3652);
nor U5492 (N_5492,N_1161,N_4236);
xor U5493 (N_5493,N_4306,N_3265);
nand U5494 (N_5494,N_1387,N_418);
and U5495 (N_5495,N_3627,N_2371);
and U5496 (N_5496,N_415,N_719);
nor U5497 (N_5497,N_4986,N_4742);
nand U5498 (N_5498,N_1622,N_3107);
nor U5499 (N_5499,N_1861,N_3861);
or U5500 (N_5500,N_136,N_4825);
xor U5501 (N_5501,N_3863,N_2140);
and U5502 (N_5502,N_2966,N_336);
and U5503 (N_5503,N_2542,N_3882);
and U5504 (N_5504,N_1591,N_3555);
and U5505 (N_5505,N_1240,N_3871);
nor U5506 (N_5506,N_1463,N_1448);
or U5507 (N_5507,N_4421,N_3465);
nand U5508 (N_5508,N_3825,N_561);
or U5509 (N_5509,N_3516,N_257);
nor U5510 (N_5510,N_2161,N_4954);
xor U5511 (N_5511,N_743,N_4243);
nor U5512 (N_5512,N_4779,N_4880);
or U5513 (N_5513,N_4768,N_4097);
nor U5514 (N_5514,N_1767,N_4356);
xor U5515 (N_5515,N_2270,N_1891);
or U5516 (N_5516,N_1427,N_1496);
nor U5517 (N_5517,N_2077,N_4277);
nand U5518 (N_5518,N_1805,N_232);
nor U5519 (N_5519,N_2370,N_2278);
nand U5520 (N_5520,N_1665,N_1828);
nand U5521 (N_5521,N_237,N_1075);
nand U5522 (N_5522,N_1397,N_4174);
nand U5523 (N_5523,N_781,N_2341);
nand U5524 (N_5524,N_4893,N_713);
or U5525 (N_5525,N_2309,N_3805);
nand U5526 (N_5526,N_4359,N_2559);
nand U5527 (N_5527,N_4941,N_1356);
nand U5528 (N_5528,N_3377,N_3653);
xor U5529 (N_5529,N_3903,N_3067);
xor U5530 (N_5530,N_1036,N_1894);
nand U5531 (N_5531,N_649,N_1136);
xor U5532 (N_5532,N_166,N_3840);
or U5533 (N_5533,N_4485,N_4898);
and U5534 (N_5534,N_1417,N_1438);
xnor U5535 (N_5535,N_3323,N_278);
nor U5536 (N_5536,N_228,N_3592);
nor U5537 (N_5537,N_2180,N_161);
nand U5538 (N_5538,N_2215,N_3764);
nand U5539 (N_5539,N_537,N_4103);
nand U5540 (N_5540,N_3604,N_1526);
nand U5541 (N_5541,N_4039,N_4068);
and U5542 (N_5542,N_2766,N_1996);
or U5543 (N_5543,N_4143,N_202);
xor U5544 (N_5544,N_4879,N_4705);
xor U5545 (N_5545,N_4342,N_4343);
xnor U5546 (N_5546,N_1593,N_4307);
nor U5547 (N_5547,N_1533,N_4569);
or U5548 (N_5548,N_1506,N_309);
nor U5549 (N_5549,N_2933,N_2068);
xnor U5550 (N_5550,N_1564,N_1305);
nand U5551 (N_5551,N_784,N_2380);
xnor U5552 (N_5552,N_4896,N_3565);
nand U5553 (N_5553,N_2988,N_3154);
xnor U5554 (N_5554,N_2050,N_2054);
or U5555 (N_5555,N_3607,N_2474);
nor U5556 (N_5556,N_2807,N_2162);
nand U5557 (N_5557,N_667,N_1964);
or U5558 (N_5558,N_3553,N_1354);
or U5559 (N_5559,N_3274,N_1714);
nand U5560 (N_5560,N_2296,N_4326);
nor U5561 (N_5561,N_2485,N_2531);
xnor U5562 (N_5562,N_1128,N_3224);
xnor U5563 (N_5563,N_472,N_2476);
nor U5564 (N_5564,N_564,N_819);
or U5565 (N_5565,N_1486,N_2060);
or U5566 (N_5566,N_2134,N_1637);
and U5567 (N_5567,N_2449,N_4215);
xnor U5568 (N_5568,N_3130,N_953);
xnor U5569 (N_5569,N_3938,N_4960);
nand U5570 (N_5570,N_1179,N_4792);
and U5571 (N_5571,N_772,N_4204);
xor U5572 (N_5572,N_4221,N_1835);
and U5573 (N_5573,N_3954,N_3539);
nand U5574 (N_5574,N_1655,N_260);
nand U5575 (N_5575,N_268,N_1299);
nand U5576 (N_5576,N_2588,N_2403);
or U5577 (N_5577,N_3038,N_3209);
or U5578 (N_5578,N_4045,N_4647);
xnor U5579 (N_5579,N_2008,N_4196);
and U5580 (N_5580,N_2152,N_992);
xnor U5581 (N_5581,N_2236,N_3759);
nand U5582 (N_5582,N_4157,N_2390);
and U5583 (N_5583,N_3430,N_4337);
xnor U5584 (N_5584,N_1951,N_3487);
and U5585 (N_5585,N_1645,N_1168);
nand U5586 (N_5586,N_4260,N_662);
or U5587 (N_5587,N_1811,N_1219);
xnor U5588 (N_5588,N_57,N_3118);
or U5589 (N_5589,N_4116,N_681);
or U5590 (N_5590,N_4618,N_3980);
nor U5591 (N_5591,N_2579,N_174);
and U5592 (N_5592,N_4011,N_2532);
or U5593 (N_5593,N_4066,N_567);
nor U5594 (N_5594,N_3162,N_2153);
nor U5595 (N_5595,N_2228,N_2443);
nor U5596 (N_5596,N_175,N_4139);
and U5597 (N_5597,N_4331,N_4594);
or U5598 (N_5598,N_3865,N_4439);
and U5599 (N_5599,N_284,N_194);
xor U5600 (N_5600,N_2357,N_1764);
nor U5601 (N_5601,N_88,N_1547);
xnor U5602 (N_5602,N_1442,N_3662);
and U5603 (N_5603,N_1139,N_2037);
or U5604 (N_5604,N_4560,N_1091);
nor U5605 (N_5605,N_2621,N_1351);
and U5606 (N_5606,N_1505,N_959);
or U5607 (N_5607,N_4769,N_2788);
and U5608 (N_5608,N_319,N_2874);
nor U5609 (N_5609,N_263,N_1909);
nor U5610 (N_5610,N_4637,N_1845);
and U5611 (N_5611,N_1866,N_4588);
nand U5612 (N_5612,N_1700,N_190);
or U5613 (N_5613,N_145,N_1303);
nand U5614 (N_5614,N_4062,N_4338);
and U5615 (N_5615,N_466,N_763);
and U5616 (N_5616,N_2572,N_1934);
or U5617 (N_5617,N_3025,N_2387);
nor U5618 (N_5618,N_3026,N_4305);
nor U5619 (N_5619,N_4778,N_4716);
nor U5620 (N_5620,N_81,N_4053);
and U5621 (N_5621,N_2251,N_3447);
nand U5622 (N_5622,N_1723,N_3112);
xor U5623 (N_5623,N_64,N_915);
nand U5624 (N_5624,N_3969,N_3248);
nand U5625 (N_5625,N_2430,N_4648);
xnor U5626 (N_5626,N_1907,N_4087);
or U5627 (N_5627,N_1478,N_2659);
nor U5628 (N_5628,N_1540,N_4512);
or U5629 (N_5629,N_2095,N_2971);
nand U5630 (N_5630,N_840,N_977);
xnor U5631 (N_5631,N_3887,N_4134);
nor U5632 (N_5632,N_2714,N_1991);
and U5633 (N_5633,N_108,N_4370);
nand U5634 (N_5634,N_3972,N_774);
nor U5635 (N_5635,N_2668,N_1431);
or U5636 (N_5636,N_4438,N_4870);
and U5637 (N_5637,N_470,N_2708);
xnor U5638 (N_5638,N_2825,N_3518);
xor U5639 (N_5639,N_2871,N_2004);
xnor U5640 (N_5640,N_1449,N_4178);
nand U5641 (N_5641,N_3149,N_4258);
nand U5642 (N_5642,N_4503,N_1624);
and U5643 (N_5643,N_3229,N_3459);
or U5644 (N_5644,N_2024,N_3416);
nor U5645 (N_5645,N_1294,N_863);
and U5646 (N_5646,N_1719,N_958);
or U5647 (N_5647,N_3301,N_1928);
nand U5648 (N_5648,N_3495,N_4405);
or U5649 (N_5649,N_3844,N_1514);
and U5650 (N_5650,N_3982,N_900);
nand U5651 (N_5651,N_2079,N_2571);
nor U5652 (N_5652,N_1585,N_4990);
or U5653 (N_5653,N_1892,N_503);
xnor U5654 (N_5654,N_3087,N_3252);
or U5655 (N_5655,N_4626,N_2794);
and U5656 (N_5656,N_2472,N_3372);
or U5657 (N_5657,N_3999,N_4872);
xnor U5658 (N_5658,N_2096,N_3228);
nor U5659 (N_5659,N_1482,N_4686);
nor U5660 (N_5660,N_3327,N_2216);
nand U5661 (N_5661,N_1188,N_3502);
nand U5662 (N_5662,N_4564,N_4854);
nor U5663 (N_5663,N_3908,N_2848);
nor U5664 (N_5664,N_4862,N_1198);
or U5665 (N_5665,N_4730,N_919);
or U5666 (N_5666,N_2507,N_2899);
or U5667 (N_5667,N_1521,N_2878);
nand U5668 (N_5668,N_2298,N_4978);
nor U5669 (N_5669,N_4177,N_2867);
xnor U5670 (N_5670,N_1167,N_1812);
xor U5671 (N_5671,N_114,N_4677);
nand U5672 (N_5672,N_1783,N_4683);
and U5673 (N_5673,N_4353,N_3661);
and U5674 (N_5674,N_2613,N_3414);
or U5675 (N_5675,N_1053,N_1634);
or U5676 (N_5676,N_357,N_3128);
or U5677 (N_5677,N_241,N_4070);
xnor U5678 (N_5678,N_851,N_4018);
and U5679 (N_5679,N_1799,N_1286);
and U5680 (N_5680,N_4997,N_424);
nor U5681 (N_5681,N_3544,N_3515);
xor U5682 (N_5682,N_2450,N_1704);
or U5683 (N_5683,N_1987,N_490);
xor U5684 (N_5684,N_4906,N_3057);
nand U5685 (N_5685,N_1418,N_2462);
xnor U5686 (N_5686,N_4128,N_1210);
xnor U5687 (N_5687,N_2253,N_4518);
xnor U5688 (N_5688,N_1051,N_3261);
nor U5689 (N_5689,N_2873,N_2723);
and U5690 (N_5690,N_509,N_296);
nor U5691 (N_5691,N_711,N_3584);
nor U5692 (N_5692,N_2210,N_4581);
xor U5693 (N_5693,N_3803,N_215);
nand U5694 (N_5694,N_2155,N_4543);
or U5695 (N_5695,N_4916,N_4535);
xor U5696 (N_5696,N_2121,N_3773);
xor U5697 (N_5697,N_1313,N_27);
nand U5698 (N_5698,N_3663,N_2124);
and U5699 (N_5699,N_48,N_1381);
and U5700 (N_5700,N_2311,N_3461);
nor U5701 (N_5701,N_1950,N_1037);
nand U5702 (N_5702,N_3250,N_2073);
and U5703 (N_5703,N_4829,N_837);
nor U5704 (N_5704,N_1236,N_3479);
and U5705 (N_5705,N_4737,N_1765);
nor U5706 (N_5706,N_1752,N_2685);
nor U5707 (N_5707,N_1888,N_2046);
nand U5708 (N_5708,N_4904,N_1263);
and U5709 (N_5709,N_1104,N_1931);
nand U5710 (N_5710,N_4154,N_3388);
xor U5711 (N_5711,N_113,N_645);
and U5712 (N_5712,N_2922,N_1422);
nor U5713 (N_5713,N_475,N_3986);
nor U5714 (N_5714,N_225,N_2840);
and U5715 (N_5715,N_270,N_474);
xor U5716 (N_5716,N_1165,N_2610);
xor U5717 (N_5717,N_3835,N_4684);
nand U5718 (N_5718,N_4490,N_2304);
and U5719 (N_5719,N_4929,N_1983);
xor U5720 (N_5720,N_2299,N_2051);
or U5721 (N_5721,N_375,N_3233);
or U5722 (N_5722,N_3621,N_1731);
or U5723 (N_5723,N_3438,N_2328);
or U5724 (N_5724,N_300,N_2226);
and U5725 (N_5725,N_463,N_1790);
nand U5726 (N_5726,N_2945,N_4416);
and U5727 (N_5727,N_1086,N_2702);
and U5728 (N_5728,N_2649,N_2350);
or U5729 (N_5729,N_2528,N_4685);
nand U5730 (N_5730,N_2339,N_4191);
and U5731 (N_5731,N_4505,N_2983);
nor U5732 (N_5732,N_402,N_1726);
nand U5733 (N_5733,N_3603,N_896);
nor U5734 (N_5734,N_1460,N_2243);
and U5735 (N_5735,N_4268,N_1644);
nand U5736 (N_5736,N_4672,N_2480);
xnor U5737 (N_5737,N_3101,N_4931);
nand U5738 (N_5738,N_2584,N_646);
nor U5739 (N_5739,N_2465,N_3993);
and U5740 (N_5740,N_3503,N_4748);
or U5741 (N_5741,N_179,N_785);
xnor U5742 (N_5742,N_4606,N_1071);
or U5743 (N_5743,N_1495,N_628);
xnor U5744 (N_5744,N_1279,N_4722);
and U5745 (N_5745,N_4575,N_2711);
or U5746 (N_5746,N_1242,N_3912);
xor U5747 (N_5747,N_778,N_3435);
nand U5748 (N_5748,N_2234,N_941);
xnor U5749 (N_5749,N_3362,N_4849);
nand U5750 (N_5750,N_1626,N_3317);
and U5751 (N_5751,N_2509,N_1461);
or U5752 (N_5752,N_4121,N_2432);
xor U5753 (N_5753,N_1705,N_4335);
nand U5754 (N_5754,N_1523,N_4298);
nor U5755 (N_5755,N_3366,N_888);
and U5756 (N_5756,N_3147,N_4227);
nand U5757 (N_5757,N_273,N_1121);
nand U5758 (N_5758,N_2400,N_2272);
nor U5759 (N_5759,N_3668,N_3815);
and U5760 (N_5760,N_3691,N_1615);
nand U5761 (N_5761,N_4315,N_1159);
and U5762 (N_5762,N_2843,N_2638);
xor U5763 (N_5763,N_787,N_3056);
xor U5764 (N_5764,N_2057,N_952);
nand U5765 (N_5765,N_435,N_3804);
xnor U5766 (N_5766,N_550,N_2344);
or U5767 (N_5767,N_2308,N_4484);
xor U5768 (N_5768,N_4377,N_4264);
or U5769 (N_5769,N_2523,N_3917);
nand U5770 (N_5770,N_149,N_3314);
or U5771 (N_5771,N_4700,N_3186);
xor U5772 (N_5772,N_4584,N_2536);
and U5773 (N_5773,N_4919,N_1918);
nor U5774 (N_5774,N_3302,N_1511);
nand U5775 (N_5775,N_4497,N_2961);
nor U5776 (N_5776,N_2810,N_501);
and U5777 (N_5777,N_2090,N_3800);
nor U5778 (N_5778,N_656,N_1905);
and U5779 (N_5779,N_4352,N_1371);
nand U5780 (N_5780,N_2184,N_2478);
nand U5781 (N_5781,N_245,N_1217);
or U5782 (N_5782,N_3961,N_3612);
xnor U5783 (N_5783,N_3463,N_1120);
nand U5784 (N_5784,N_4392,N_3909);
or U5785 (N_5785,N_2455,N_1657);
nor U5786 (N_5786,N_1137,N_4458);
and U5787 (N_5787,N_4697,N_3702);
and U5788 (N_5788,N_3964,N_1942);
xnor U5789 (N_5789,N_4917,N_3094);
xor U5790 (N_5790,N_873,N_1078);
and U5791 (N_5791,N_4310,N_4933);
and U5792 (N_5792,N_3305,N_2735);
or U5793 (N_5793,N_4404,N_203);
or U5794 (N_5794,N_1941,N_246);
xnor U5795 (N_5795,N_3715,N_3326);
nand U5796 (N_5796,N_1952,N_2190);
or U5797 (N_5797,N_4446,N_2625);
nand U5798 (N_5798,N_3755,N_2290);
or U5799 (N_5799,N_737,N_3852);
and U5800 (N_5800,N_1724,N_2671);
or U5801 (N_5801,N_1010,N_892);
xor U5802 (N_5802,N_4079,N_1580);
and U5803 (N_5803,N_4770,N_1399);
xnor U5804 (N_5804,N_3931,N_3849);
and U5805 (N_5805,N_868,N_750);
nand U5806 (N_5806,N_782,N_1017);
or U5807 (N_5807,N_4297,N_3021);
nor U5808 (N_5808,N_1574,N_338);
and U5809 (N_5809,N_3382,N_2013);
and U5810 (N_5810,N_1869,N_2997);
nor U5811 (N_5811,N_3369,N_393);
nand U5812 (N_5812,N_4963,N_3223);
and U5813 (N_5813,N_4482,N_2098);
nand U5814 (N_5814,N_1160,N_3203);
xnor U5815 (N_5815,N_1803,N_1046);
nor U5816 (N_5816,N_2256,N_2286);
nand U5817 (N_5817,N_3219,N_1011);
or U5818 (N_5818,N_720,N_1874);
or U5819 (N_5819,N_2953,N_269);
and U5820 (N_5820,N_2423,N_4544);
nor U5821 (N_5821,N_4027,N_597);
nor U5822 (N_5822,N_1984,N_3679);
nand U5823 (N_5823,N_3802,N_3497);
nand U5824 (N_5824,N_4250,N_2929);
and U5825 (N_5825,N_2901,N_4075);
nand U5826 (N_5826,N_668,N_2826);
or U5827 (N_5827,N_3817,N_3408);
or U5828 (N_5828,N_1481,N_4993);
nor U5829 (N_5829,N_2145,N_4617);
and U5830 (N_5830,N_986,N_4382);
and U5831 (N_5831,N_2615,N_1216);
or U5832 (N_5832,N_2819,N_3019);
or U5833 (N_5833,N_4325,N_708);
and U5834 (N_5834,N_2797,N_3072);
and U5835 (N_5835,N_2709,N_2805);
and U5836 (N_5836,N_3020,N_162);
nand U5837 (N_5837,N_2860,N_4688);
nand U5838 (N_5838,N_1573,N_4624);
nand U5839 (N_5839,N_824,N_1722);
or U5840 (N_5840,N_1365,N_4300);
nand U5841 (N_5841,N_3033,N_4602);
or U5842 (N_5842,N_4444,N_951);
and U5843 (N_5843,N_1579,N_2321);
nor U5844 (N_5844,N_4772,N_2537);
nor U5845 (N_5845,N_4152,N_1949);
or U5846 (N_5846,N_2208,N_2641);
or U5847 (N_5847,N_519,N_79);
and U5848 (N_5848,N_955,N_721);
nand U5849 (N_5849,N_421,N_931);
nor U5850 (N_5850,N_384,N_2948);
nand U5851 (N_5851,N_2679,N_2594);
and U5852 (N_5852,N_3650,N_2275);
nor U5853 (N_5853,N_2368,N_3177);
and U5854 (N_5854,N_3458,N_3426);
and U5855 (N_5855,N_2884,N_2746);
nor U5856 (N_5856,N_2540,N_2318);
or U5857 (N_5857,N_4168,N_4210);
and U5858 (N_5858,N_4891,N_86);
nand U5859 (N_5859,N_3958,N_2248);
nor U5860 (N_5860,N_926,N_2259);
nand U5861 (N_5861,N_999,N_3754);
and U5862 (N_5862,N_3123,N_3146);
or U5863 (N_5863,N_2762,N_3786);
or U5864 (N_5864,N_3513,N_4115);
nand U5865 (N_5865,N_4531,N_4431);
nor U5866 (N_5866,N_3165,N_458);
and U5867 (N_5867,N_1721,N_3411);
xor U5868 (N_5868,N_828,N_2779);
nor U5869 (N_5869,N_4029,N_3355);
nand U5870 (N_5870,N_4727,N_3493);
nor U5871 (N_5871,N_1376,N_1469);
and U5872 (N_5872,N_971,N_3929);
nand U5873 (N_5873,N_3700,N_3895);
xnor U5874 (N_5874,N_1215,N_3329);
xnor U5875 (N_5875,N_579,N_4902);
xor U5876 (N_5876,N_3339,N_2626);
nand U5877 (N_5877,N_326,N_1477);
and U5878 (N_5878,N_3541,N_1519);
and U5879 (N_5879,N_2101,N_4119);
nand U5880 (N_5880,N_3361,N_729);
and U5881 (N_5881,N_2914,N_214);
nand U5882 (N_5882,N_341,N_460);
nor U5883 (N_5883,N_1040,N_1969);
and U5884 (N_5884,N_3601,N_3659);
nand U5885 (N_5885,N_535,N_2085);
and U5886 (N_5886,N_3569,N_2696);
and U5887 (N_5887,N_2441,N_1956);
nor U5888 (N_5888,N_3599,N_3637);
or U5889 (N_5889,N_3088,N_3258);
or U5890 (N_5890,N_552,N_2783);
xnor U5891 (N_5891,N_3859,N_156);
and U5892 (N_5892,N_2273,N_1777);
nand U5893 (N_5893,N_4802,N_752);
and U5894 (N_5894,N_3168,N_4641);
nor U5895 (N_5895,N_3716,N_4720);
xnor U5896 (N_5896,N_4146,N_585);
nor U5897 (N_5897,N_2782,N_3126);
nor U5898 (N_5898,N_4481,N_4478);
and U5899 (N_5899,N_4603,N_830);
xnor U5900 (N_5900,N_2713,N_1948);
nand U5901 (N_5901,N_2066,N_437);
nand U5902 (N_5902,N_3712,N_267);
xor U5903 (N_5903,N_1679,N_2868);
nand U5904 (N_5904,N_3125,N_1249);
nor U5905 (N_5905,N_2527,N_1551);
xor U5906 (N_5906,N_457,N_3004);
nor U5907 (N_5907,N_1068,N_23);
or U5908 (N_5908,N_2887,N_876);
or U5909 (N_5909,N_1612,N_3729);
and U5910 (N_5910,N_2720,N_1380);
or U5911 (N_5911,N_764,N_2958);
or U5912 (N_5912,N_1758,N_3722);
nor U5913 (N_5913,N_1978,N_264);
or U5914 (N_5914,N_2870,N_2549);
xor U5915 (N_5915,N_4229,N_445);
xor U5916 (N_5916,N_3394,N_4582);
nor U5917 (N_5917,N_3906,N_4837);
or U5918 (N_5918,N_3047,N_1557);
xor U5919 (N_5919,N_4471,N_1122);
xor U5920 (N_5920,N_2486,N_2585);
and U5921 (N_5921,N_2358,N_3002);
nand U5922 (N_5922,N_738,N_3528);
nand U5923 (N_5923,N_4043,N_2295);
or U5924 (N_5924,N_1293,N_1932);
nand U5925 (N_5925,N_557,N_625);
nand U5926 (N_5926,N_1683,N_41);
nand U5927 (N_5927,N_3644,N_2574);
nand U5928 (N_5928,N_3296,N_3480);
or U5929 (N_5929,N_2048,N_1133);
or U5930 (N_5930,N_2904,N_2755);
and U5931 (N_5931,N_1599,N_663);
xnor U5932 (N_5932,N_4407,N_1288);
nor U5933 (N_5933,N_497,N_89);
xnor U5934 (N_5934,N_4735,N_3564);
nor U5935 (N_5935,N_1604,N_940);
nor U5936 (N_5936,N_2310,N_546);
nor U5937 (N_5937,N_705,N_3558);
and U5938 (N_5938,N_3766,N_4645);
nor U5939 (N_5939,N_3704,N_46);
nor U5940 (N_5940,N_4669,N_4165);
xnor U5941 (N_5941,N_3971,N_339);
nor U5942 (N_5942,N_1329,N_3151);
and U5943 (N_5943,N_689,N_3240);
xor U5944 (N_5944,N_3566,N_2198);
xnor U5945 (N_5945,N_860,N_1697);
nand U5946 (N_5946,N_4934,N_4270);
nor U5947 (N_5947,N_4595,N_2908);
xnor U5948 (N_5948,N_4054,N_568);
or U5949 (N_5949,N_4830,N_1824);
or U5950 (N_5950,N_864,N_831);
nor U5951 (N_5951,N_3910,N_950);
xnor U5952 (N_5952,N_2583,N_1749);
xnor U5953 (N_5953,N_3148,N_1346);
xor U5954 (N_5954,N_2349,N_394);
xor U5955 (N_5955,N_1290,N_2189);
xor U5956 (N_5956,N_4869,N_2728);
nor U5957 (N_5957,N_4388,N_1497);
and U5958 (N_5958,N_184,N_2799);
nor U5959 (N_5959,N_683,N_1389);
and U5960 (N_5960,N_1884,N_2674);
or U5961 (N_5961,N_3655,N_2545);
xnor U5962 (N_5962,N_4985,N_559);
xor U5963 (N_5963,N_3397,N_178);
and U5964 (N_5964,N_4845,N_4633);
nand U5965 (N_5965,N_1271,N_4415);
nor U5966 (N_5966,N_666,N_208);
nand U5967 (N_5967,N_1044,N_157);
or U5968 (N_5968,N_2130,N_4763);
or U5969 (N_5969,N_2750,N_2628);
nand U5970 (N_5970,N_3876,N_2192);
xnor U5971 (N_5971,N_4915,N_55);
nor U5972 (N_5972,N_651,N_3845);
or U5973 (N_5973,N_4756,N_4913);
nor U5974 (N_5974,N_3284,N_815);
nand U5975 (N_5975,N_4670,N_1808);
nor U5976 (N_5976,N_2519,N_1416);
or U5977 (N_5977,N_1260,N_2598);
nand U5978 (N_5978,N_4940,N_5);
nand U5979 (N_5979,N_1398,N_2242);
and U5980 (N_5980,N_3848,N_4650);
xnor U5981 (N_5981,N_2602,N_3322);
and U5982 (N_5982,N_3445,N_3471);
or U5983 (N_5983,N_706,N_4345);
nand U5984 (N_5984,N_1677,N_751);
xor U5985 (N_5985,N_289,N_258);
nand U5986 (N_5986,N_1971,N_4767);
xor U5987 (N_5987,N_2247,N_3656);
xnor U5988 (N_5988,N_3751,N_2563);
nand U5989 (N_5989,N_3434,N_4701);
nor U5990 (N_5990,N_4254,N_3182);
or U5991 (N_5991,N_3343,N_151);
xnor U5992 (N_5992,N_2960,N_637);
or U5993 (N_5993,N_993,N_2151);
nand U5994 (N_5994,N_1033,N_1338);
nor U5995 (N_5995,N_4396,N_2644);
xor U5996 (N_5996,N_2596,N_4562);
or U5997 (N_5997,N_1238,N_3689);
nand U5998 (N_5998,N_1493,N_1388);
and U5999 (N_5999,N_2181,N_844);
nand U6000 (N_6000,N_4553,N_563);
and U6001 (N_6001,N_1850,N_256);
nand U6002 (N_6002,N_294,N_389);
xor U6003 (N_6003,N_42,N_2398);
nand U6004 (N_6004,N_2891,N_909);
nand U6005 (N_6005,N_4949,N_4493);
xor U6006 (N_6006,N_1779,N_1911);
nor U6007 (N_6007,N_2781,N_4483);
or U6008 (N_6008,N_3379,N_4936);
and U6009 (N_6009,N_4001,N_1654);
or U6010 (N_6010,N_4106,N_3373);
nor U6011 (N_6011,N_1886,N_3809);
nand U6012 (N_6012,N_3501,N_3051);
and U6013 (N_6013,N_3636,N_2724);
xor U6014 (N_6014,N_4025,N_3960);
nor U6015 (N_6015,N_2442,N_3035);
xnor U6016 (N_6016,N_3346,N_2775);
or U6017 (N_6017,N_1394,N_3580);
xnor U6018 (N_6018,N_1801,N_3499);
and U6019 (N_6019,N_4127,N_4739);
and U6020 (N_6020,N_2305,N_140);
xnor U6021 (N_6021,N_1676,N_2075);
nor U6022 (N_6022,N_701,N_4820);
nand U6023 (N_6023,N_2458,N_4181);
nor U6024 (N_6024,N_40,N_2244);
and U6025 (N_6025,N_914,N_1029);
nand U6026 (N_6026,N_4194,N_3963);
and U6027 (N_6027,N_827,N_187);
and U6028 (N_6028,N_1785,N_236);
and U6029 (N_6029,N_3155,N_1939);
xnor U6030 (N_6030,N_4743,N_3360);
or U6031 (N_6031,N_3137,N_580);
xnor U6032 (N_6032,N_4013,N_3866);
or U6033 (N_6033,N_1818,N_19);
nand U6034 (N_6034,N_371,N_1097);
and U6035 (N_6035,N_2132,N_4172);
xor U6036 (N_6036,N_4856,N_3195);
or U6037 (N_6037,N_3873,N_1675);
and U6038 (N_6038,N_2590,N_990);
nand U6039 (N_6039,N_310,N_4774);
and U6040 (N_6040,N_3736,N_159);
and U6041 (N_6041,N_1125,N_3092);
xor U6042 (N_6042,N_4980,N_4410);
or U6043 (N_6043,N_2194,N_2467);
xor U6044 (N_6044,N_3915,N_2034);
or U6045 (N_6045,N_4863,N_1411);
nor U6046 (N_6046,N_1328,N_2832);
or U6047 (N_6047,N_3160,N_826);
nand U6048 (N_6048,N_33,N_1343);
or U6049 (N_6049,N_2178,N_4046);
or U6050 (N_6050,N_3190,N_4486);
nor U6051 (N_6051,N_3666,N_2137);
and U6052 (N_6052,N_4614,N_1450);
nand U6053 (N_6053,N_1323,N_1164);
and U6054 (N_6054,N_1034,N_4745);
nor U6055 (N_6055,N_4957,N_692);
xnor U6056 (N_6056,N_4979,N_3632);
nand U6057 (N_6057,N_53,N_2315);
and U6058 (N_6058,N_4866,N_4680);
nand U6059 (N_6059,N_1962,N_4925);
and U6060 (N_6060,N_1266,N_669);
nand U6061 (N_6061,N_2176,N_207);
or U6062 (N_6062,N_2133,N_788);
nand U6063 (N_6063,N_3345,N_511);
and U6064 (N_6064,N_4775,N_1089);
nor U6065 (N_6065,N_3475,N_272);
xor U6066 (N_6066,N_1531,N_2207);
nor U6067 (N_6067,N_2734,N_1278);
or U6068 (N_6068,N_139,N_2974);
or U6069 (N_6069,N_2306,N_2993);
nor U6070 (N_6070,N_638,N_1858);
xnor U6071 (N_6071,N_2855,N_3288);
and U6072 (N_6072,N_3941,N_2330);
nor U6073 (N_6073,N_2844,N_731);
nand U6074 (N_6074,N_4724,N_4984);
nand U6075 (N_6075,N_982,N_893);
or U6076 (N_6076,N_168,N_334);
nor U6077 (N_6077,N_3683,N_4828);
xor U6078 (N_6078,N_2300,N_4509);
nor U6079 (N_6079,N_2030,N_1339);
or U6080 (N_6080,N_1,N_963);
or U6081 (N_6081,N_3546,N_879);
nand U6082 (N_6082,N_1041,N_4373);
nor U6083 (N_6083,N_1494,N_163);
and U6084 (N_6084,N_2561,N_1178);
or U6085 (N_6085,N_2067,N_1395);
nor U6086 (N_6086,N_3281,N_1231);
nor U6087 (N_6087,N_4956,N_3039);
and U6088 (N_6088,N_3595,N_427);
xor U6089 (N_6089,N_2558,N_4363);
nor U6090 (N_6090,N_757,N_901);
nor U6091 (N_6091,N_2541,N_2575);
and U6092 (N_6092,N_493,N_1875);
or U6093 (N_6093,N_867,N_2061);
xor U6094 (N_6094,N_3210,N_2567);
nand U6095 (N_6095,N_3705,N_1774);
xor U6096 (N_6096,N_2882,N_1064);
and U6097 (N_6097,N_2429,N_4731);
nand U6098 (N_6098,N_1038,N_2515);
nand U6099 (N_6099,N_747,N_4132);
nor U6100 (N_6100,N_2503,N_3667);
and U6101 (N_6101,N_1701,N_2888);
nor U6102 (N_6102,N_4434,N_1499);
and U6103 (N_6103,N_3098,N_3506);
or U6104 (N_6104,N_945,N_4567);
or U6105 (N_6105,N_1804,N_1906);
and U6106 (N_6106,N_2935,N_4534);
or U6107 (N_6107,N_853,N_1106);
and U6108 (N_6108,N_1550,N_321);
and U6109 (N_6109,N_1565,N_2624);
xor U6110 (N_6110,N_3940,N_3297);
xor U6111 (N_6111,N_994,N_3062);
xnor U6112 (N_6112,N_4262,N_4579);
or U6113 (N_6113,N_3855,N_3);
nor U6114 (N_6114,N_3235,N_4818);
nor U6115 (N_6115,N_1425,N_2438);
xnor U6116 (N_6116,N_1543,N_4890);
and U6117 (N_6117,N_4267,N_1590);
nor U6118 (N_6118,N_1876,N_2965);
nand U6119 (N_6119,N_1847,N_4333);
nor U6120 (N_6120,N_1362,N_4708);
nor U6121 (N_6121,N_1069,N_923);
nand U6122 (N_6122,N_1823,N_2972);
nor U6123 (N_6123,N_4032,N_4261);
or U6124 (N_6124,N_1200,N_4472);
nand U6125 (N_6125,N_3818,N_3234);
nor U6126 (N_6126,N_66,N_4638);
xor U6127 (N_6127,N_1291,N_1586);
and U6128 (N_6128,N_407,N_624);
xnor U6129 (N_6129,N_1693,N_4099);
nand U6130 (N_6130,N_3163,N_3378);
nand U6131 (N_6131,N_1739,N_1829);
and U6132 (N_6132,N_2740,N_409);
xor U6133 (N_6133,N_4440,N_1684);
xnor U6134 (N_6134,N_3158,N_2017);
nand U6135 (N_6135,N_342,N_3029);
nand U6136 (N_6136,N_2691,N_3184);
and U6137 (N_6137,N_1186,N_1311);
nand U6138 (N_6138,N_2992,N_2980);
or U6139 (N_6139,N_4823,N_4801);
nor U6140 (N_6140,N_3066,N_4246);
and U6141 (N_6141,N_1509,N_3671);
nand U6142 (N_6142,N_517,N_1780);
or U6143 (N_6143,N_1879,N_2006);
nand U6144 (N_6144,N_368,N_4275);
xor U6145 (N_6145,N_405,N_3669);
xor U6146 (N_6146,N_3821,N_4199);
nor U6147 (N_6147,N_1613,N_4133);
and U6148 (N_6148,N_3620,N_306);
xor U6149 (N_6149,N_3048,N_2678);
xor U6150 (N_6150,N_4574,N_3843);
xor U6151 (N_6151,N_2001,N_3600);
xnor U6152 (N_6152,N_4951,N_3989);
nand U6153 (N_6153,N_1307,N_3778);
xor U6154 (N_6154,N_4981,N_3257);
or U6155 (N_6155,N_2193,N_4432);
xnor U6156 (N_6156,N_4982,N_4219);
nor U6157 (N_6157,N_3325,N_4758);
or U6158 (N_6158,N_2284,N_1146);
xnor U6159 (N_6159,N_1647,N_4408);
nor U6160 (N_6160,N_2562,N_1900);
and U6161 (N_6161,N_699,N_859);
xor U6162 (N_6162,N_2957,N_4135);
nand U6163 (N_6163,N_4649,N_3109);
and U6164 (N_6164,N_2698,N_556);
nand U6165 (N_6165,N_839,N_167);
xnor U6166 (N_6166,N_2548,N_3987);
and U6167 (N_6167,N_2264,N_4401);
or U6168 (N_6168,N_3044,N_907);
and U6169 (N_6169,N_239,N_4159);
xnor U6170 (N_6170,N_2576,N_3588);
nor U6171 (N_6171,N_2820,N_277);
nor U6172 (N_6172,N_117,N_4111);
or U6173 (N_6173,N_3768,N_240);
and U6174 (N_6174,N_846,N_3794);
nor U6175 (N_6175,N_3365,N_933);
xor U6176 (N_6176,N_3396,N_4537);
or U6177 (N_6177,N_658,N_2682);
and U6178 (N_6178,N_4831,N_2399);
nor U6179 (N_6179,N_127,N_3024);
and U6180 (N_6180,N_3277,N_1088);
nand U6181 (N_6181,N_1938,N_2347);
xor U6182 (N_6182,N_1966,N_1473);
nor U6183 (N_6183,N_1076,N_2492);
nor U6184 (N_6184,N_1558,N_4022);
and U6185 (N_6185,N_1370,N_4380);
nand U6186 (N_6186,N_4622,N_1484);
nor U6187 (N_6187,N_916,N_3847);
or U6188 (N_6188,N_2329,N_1625);
and U6189 (N_6189,N_2704,N_800);
nand U6190 (N_6190,N_1904,N_1221);
nor U6191 (N_6191,N_4796,N_487);
xor U6192 (N_6192,N_2197,N_3164);
and U6193 (N_6193,N_4418,N_3206);
nand U6194 (N_6194,N_4360,N_4036);
xnor U6195 (N_6195,N_4213,N_2730);
or U6196 (N_6196,N_221,N_2241);
nand U6197 (N_6197,N_0,N_3268);
nand U6198 (N_6198,N_1885,N_3340);
or U6199 (N_6199,N_4065,N_1746);
or U6200 (N_6200,N_4976,N_504);
and U6201 (N_6201,N_2159,N_3760);
nand U6202 (N_6202,N_274,N_2599);
xor U6203 (N_6203,N_4894,N_1085);
and U6204 (N_6204,N_523,N_1030);
or U6205 (N_6205,N_2424,N_2335);
or U6206 (N_6206,N_1862,N_4336);
and U6207 (N_6207,N_3527,N_1059);
or U6208 (N_6208,N_1243,N_792);
nor U6209 (N_6209,N_1627,N_2606);
and U6210 (N_6210,N_2238,N_688);
xor U6211 (N_6211,N_3881,N_2854);
xnor U6212 (N_6212,N_4301,N_1756);
xnor U6213 (N_6213,N_3053,N_1220);
or U6214 (N_6214,N_288,N_1403);
or U6215 (N_6215,N_2811,N_465);
and U6216 (N_6216,N_3878,N_4806);
and U6217 (N_6217,N_2042,N_2890);
nand U6218 (N_6218,N_584,N_2654);
xor U6219 (N_6219,N_1090,N_1650);
nor U6220 (N_6220,N_2511,N_2471);
nor U6221 (N_6221,N_2035,N_1667);
nand U6222 (N_6222,N_3583,N_2279);
nor U6223 (N_6223,N_2003,N_4020);
or U6224 (N_6224,N_3777,N_3256);
or U6225 (N_6225,N_63,N_1833);
nor U6226 (N_6226,N_2393,N_2392);
or U6227 (N_6227,N_3319,N_252);
and U6228 (N_6228,N_2297,N_2892);
or U6229 (N_6229,N_4813,N_4679);
nor U6230 (N_6230,N_3926,N_2374);
and U6231 (N_6231,N_1755,N_403);
nor U6232 (N_6232,N_1349,N_587);
nor U6233 (N_6233,N_9,N_3387);
and U6234 (N_6234,N_4038,N_3150);
or U6235 (N_6235,N_4141,N_3677);
nor U6236 (N_6236,N_4607,N_934);
nand U6237 (N_6237,N_725,N_703);
or U6238 (N_6238,N_2342,N_97);
nand U6239 (N_6239,N_2520,N_1561);
or U6240 (N_6240,N_1893,N_1589);
or U6241 (N_6241,N_1466,N_1024);
nand U6242 (N_6242,N_2246,N_3489);
nor U6243 (N_6243,N_1350,N_4805);
and U6244 (N_6244,N_3174,N_1988);
nand U6245 (N_6245,N_574,N_1325);
xnor U6246 (N_6246,N_3006,N_2188);
nand U6247 (N_6247,N_98,N_4489);
nand U6248 (N_6248,N_4449,N_4765);
and U6249 (N_6249,N_3007,N_1761);
or U6250 (N_6250,N_3254,N_4021);
and U6251 (N_6251,N_3227,N_2669);
nor U6252 (N_6252,N_4819,N_279);
xnor U6253 (N_6253,N_2934,N_4576);
xor U6254 (N_6254,N_4319,N_4738);
nand U6255 (N_6255,N_4507,N_4164);
and U6256 (N_6256,N_2635,N_3001);
or U6257 (N_6257,N_186,N_1285);
nor U6258 (N_6258,N_3500,N_1201);
and U6259 (N_6259,N_372,N_2185);
and U6260 (N_6260,N_2586,N_2086);
or U6261 (N_6261,N_118,N_765);
xor U6262 (N_6262,N_2240,N_4042);
nor U6263 (N_6263,N_4572,N_4339);
nor U6264 (N_6264,N_755,N_3059);
nand U6265 (N_6265,N_4500,N_4987);
or U6266 (N_6266,N_3131,N_4274);
xor U6267 (N_6267,N_3452,N_3412);
xnor U6268 (N_6268,N_74,N_379);
or U6269 (N_6269,N_1816,N_2716);
xnor U6270 (N_6270,N_4907,N_2043);
and U6271 (N_6271,N_2705,N_1748);
nand U6272 (N_6272,N_4965,N_3827);
and U6273 (N_6273,N_1412,N_3642);
nand U6274 (N_6274,N_476,N_4402);
nor U6275 (N_6275,N_4945,N_1691);
xnor U6276 (N_6276,N_4256,N_4741);
xor U6277 (N_6277,N_2552,N_1156);
xor U6278 (N_6278,N_3161,N_2865);
nor U6279 (N_6279,N_4253,N_2700);
or U6280 (N_6280,N_3769,N_619);
xnor U6281 (N_6281,N_3260,N_1407);
or U6282 (N_6282,N_2684,N_1621);
or U6283 (N_6283,N_4266,N_3533);
and U6284 (N_6284,N_4803,N_1308);
or U6285 (N_6285,N_2902,N_398);
or U6286 (N_6286,N_4200,N_4811);
xor U6287 (N_6287,N_4547,N_1364);
nand U6288 (N_6288,N_182,N_4546);
nor U6289 (N_6289,N_76,N_1296);
nor U6290 (N_6290,N_3799,N_4425);
or U6291 (N_6291,N_1130,N_3037);
xor U6292 (N_6292,N_142,N_325);
nand U6293 (N_6293,N_2605,N_2538);
xor U6294 (N_6294,N_4285,N_119);
and U6295 (N_6295,N_2614,N_1414);
nor U6296 (N_6296,N_841,N_3708);
nand U6297 (N_6297,N_857,N_2271);
nor U6298 (N_6298,N_3898,N_2109);
xnor U6299 (N_6299,N_24,N_3468);
and U6300 (N_6300,N_1095,N_3180);
nor U6301 (N_6301,N_2616,N_4413);
or U6302 (N_6302,N_3756,N_3282);
nand U6303 (N_6303,N_3208,N_1837);
or U6304 (N_6304,N_4272,N_2088);
xor U6305 (N_6305,N_3318,N_1316);
nor U6306 (N_6306,N_2701,N_894);
xor U6307 (N_6307,N_650,N_4892);
or U6308 (N_6308,N_3046,N_4883);
nor U6309 (N_6309,N_2036,N_1594);
xnor U6310 (N_6310,N_1347,N_3255);
nand U6311 (N_6311,N_3285,N_144);
nand U6312 (N_6312,N_1562,N_1649);
nand U6313 (N_6313,N_3747,N_56);
nor U6314 (N_6314,N_1947,N_2022);
and U6315 (N_6315,N_2506,N_1459);
or U6316 (N_6316,N_35,N_250);
nor U6317 (N_6317,N_51,N_4292);
xor U6318 (N_6318,N_3945,N_2546);
xnor U6319 (N_6319,N_2007,N_4975);
nor U6320 (N_6320,N_1246,N_2706);
or U6321 (N_6321,N_2964,N_2428);
or U6322 (N_6322,N_4822,N_524);
or U6323 (N_6323,N_2555,N_2396);
or U6324 (N_6324,N_1709,N_2697);
or U6325 (N_6325,N_36,N_4384);
and U6326 (N_6326,N_322,N_2879);
and U6327 (N_6327,N_2849,N_4422);
nand U6328 (N_6328,N_4475,N_4886);
and U6329 (N_6329,N_1554,N_4867);
and U6330 (N_6330,N_1277,N_3925);
and U6331 (N_6331,N_4747,N_4777);
nor U6332 (N_6332,N_2747,N_891);
nor U6333 (N_6333,N_4457,N_947);
nand U6334 (N_6334,N_1180,N_3272);
nand U6335 (N_6335,N_2677,N_759);
and U6336 (N_6336,N_2817,N_1324);
nor U6337 (N_6337,N_3432,N_298);
and U6338 (N_6338,N_2982,N_4992);
nand U6339 (N_6339,N_1916,N_3111);
or U6340 (N_6340,N_1849,N_2361);
or U6341 (N_6341,N_3467,N_1383);
xor U6342 (N_6342,N_4715,N_3334);
and U6343 (N_6343,N_4625,N_3891);
and U6344 (N_6344,N_452,N_4876);
xor U6345 (N_6345,N_1940,N_3697);
or U6346 (N_6346,N_3949,N_4100);
or U6347 (N_6347,N_430,N_676);
and U6348 (N_6348,N_4850,N_3733);
nand U6349 (N_6349,N_1049,N_18);
nor U6350 (N_6350,N_1192,N_1838);
nand U6351 (N_6351,N_1681,N_3185);
and U6352 (N_6352,N_1112,N_1843);
and U6353 (N_6353,N_3074,N_949);
nand U6354 (N_6354,N_1203,N_468);
nor U6355 (N_6355,N_1452,N_2754);
or U6356 (N_6356,N_3832,N_4291);
xnor U6357 (N_6357,N_1176,N_400);
or U6358 (N_6358,N_1252,N_206);
and U6359 (N_6359,N_2417,N_979);
or U6360 (N_6360,N_4092,N_50);
nand U6361 (N_6361,N_488,N_3633);
nor U6362 (N_6362,N_1698,N_87);
nand U6363 (N_6363,N_870,N_1114);
or U6364 (N_6364,N_1502,N_4681);
nand U6365 (N_6365,N_1680,N_3474);
nor U6366 (N_6366,N_3797,N_1967);
xnor U6367 (N_6367,N_1658,N_1363);
nor U6368 (N_6368,N_2314,N_1986);
nor U6369 (N_6369,N_834,N_4709);
and U6370 (N_6370,N_1809,N_3619);
nor U6371 (N_6371,N_1405,N_3735);
or U6372 (N_6372,N_4145,N_3171);
or U6373 (N_6373,N_2673,N_486);
and U6374 (N_6374,N_1255,N_2529);
nor U6375 (N_6375,N_2262,N_3170);
and U6376 (N_6376,N_4832,N_558);
and U6377 (N_6377,N_3959,N_4782);
xnor U6378 (N_6378,N_2944,N_2551);
or U6379 (N_6379,N_3402,N_2609);
or U6380 (N_6380,N_2276,N_1304);
or U6381 (N_6381,N_3966,N_3734);
nand U6382 (N_6382,N_803,N_2809);
or U6383 (N_6383,N_3267,N_4578);
and U6384 (N_6384,N_216,N_3455);
and U6385 (N_6385,N_1345,N_1052);
and U6386 (N_6386,N_103,N_3554);
or U6387 (N_6387,N_3692,N_780);
or U6388 (N_6388,N_2568,N_591);
nor U6389 (N_6389,N_1195,N_885);
and U6390 (N_6390,N_3249,N_4428);
nand U6391 (N_6391,N_2658,N_4580);
nand U6392 (N_6392,N_3785,N_630);
nand U6393 (N_6393,N_434,N_3504);
xor U6394 (N_6394,N_4599,N_148);
nand U6395 (N_6395,N_1015,N_1001);
nor U6396 (N_6396,N_3922,N_1685);
nor U6397 (N_6397,N_2823,N_4323);
and U6398 (N_6398,N_2842,N_2841);
and U6399 (N_6399,N_2687,N_2232);
nand U6400 (N_6400,N_3645,N_3680);
nand U6401 (N_6401,N_1762,N_3727);
nand U6402 (N_6402,N_869,N_429);
or U6403 (N_6403,N_3113,N_1919);
or U6404 (N_6404,N_939,N_608);
nor U6405 (N_6405,N_1401,N_2514);
nand U6406 (N_6406,N_150,N_391);
nor U6407 (N_6407,N_448,N_3524);
or U6408 (N_6408,N_2383,N_4824);
nor U6409 (N_6409,N_4007,N_1072);
and U6410 (N_6410,N_4465,N_3028);
nor U6411 (N_6411,N_3990,N_3017);
and U6412 (N_6412,N_2683,N_1993);
and U6413 (N_6413,N_1337,N_1464);
nor U6414 (N_6414,N_2573,N_4279);
nor U6415 (N_6415,N_1820,N_1914);
nand U6416 (N_6416,N_3011,N_1836);
or U6417 (N_6417,N_2675,N_991);
nand U6418 (N_6418,N_4776,N_4094);
nor U6419 (N_6419,N_3520,N_62);
nand U6420 (N_6420,N_4551,N_1222);
xnor U6421 (N_6421,N_4903,N_4643);
and U6422 (N_6422,N_4461,N_507);
and U6423 (N_6423,N_2388,N_4646);
xor U6424 (N_6424,N_1759,N_648);
and U6425 (N_6425,N_1248,N_2352);
xnor U6426 (N_6426,N_1522,N_285);
and U6427 (N_6427,N_2525,N_1689);
nand U6428 (N_6428,N_702,N_513);
and U6429 (N_6429,N_1570,N_3437);
nand U6430 (N_6430,N_4736,N_3065);
and U6431 (N_6431,N_4378,N_1406);
and U6432 (N_6432,N_3443,N_3701);
and U6433 (N_6433,N_364,N_612);
or U6434 (N_6434,N_722,N_3862);
nor U6435 (N_6435,N_847,N_906);
xor U6436 (N_6436,N_3530,N_4393);
nand U6437 (N_6437,N_376,N_4211);
nor U6438 (N_6438,N_903,N_3496);
xor U6439 (N_6439,N_974,N_2688);
nand U6440 (N_6440,N_3806,N_603);
xor U6441 (N_6441,N_4223,N_3970);
nor U6442 (N_6442,N_4469,N_2828);
nand U6443 (N_6443,N_4375,N_1327);
nor U6444 (N_6444,N_8,N_793);
xor U6445 (N_6445,N_4809,N_80);
and U6446 (N_6446,N_4271,N_4840);
xnor U6447 (N_6447,N_3739,N_4124);
xnor U6448 (N_6448,N_2260,N_209);
xor U6449 (N_6449,N_2925,N_1378);
xor U6450 (N_6450,N_1744,N_3836);
xnor U6451 (N_6451,N_2171,N_2955);
nand U6452 (N_6452,N_779,N_2906);
nand U6453 (N_6453,N_1841,N_2166);
nor U6454 (N_6454,N_4644,N_3178);
or U6455 (N_6455,N_1961,N_3139);
nand U6456 (N_6456,N_318,N_1527);
xor U6457 (N_6457,N_2886,N_1182);
nor U6458 (N_6458,N_4147,N_2040);
or U6459 (N_6459,N_111,N_526);
nand U6460 (N_6460,N_1760,N_724);
and U6461 (N_6461,N_2058,N_1517);
or U6462 (N_6462,N_4947,N_3442);
xnor U6463 (N_6463,N_2943,N_3243);
nor U6464 (N_6464,N_3976,N_3143);
xor U6465 (N_6465,N_4864,N_1157);
or U6466 (N_6466,N_2147,N_3611);
and U6467 (N_6467,N_335,N_2791);
and U6468 (N_6468,N_1148,N_704);
xor U6469 (N_6469,N_1840,N_807);
and U6470 (N_6470,N_3476,N_881);
and U6471 (N_6471,N_2656,N_4044);
nor U6472 (N_6472,N_753,N_685);
xnor U6473 (N_6473,N_1334,N_1922);
nor U6474 (N_6474,N_60,N_3095);
and U6475 (N_6475,N_4520,N_533);
and U6476 (N_6476,N_2872,N_2726);
nand U6477 (N_6477,N_2582,N_1392);
nor U6478 (N_6478,N_295,N_1087);
and U6479 (N_6479,N_3375,N_1834);
nor U6480 (N_6480,N_2418,N_4541);
or U6481 (N_6481,N_3942,N_1491);
xor U6482 (N_6482,N_790,N_4900);
nor U6483 (N_6483,N_1444,N_2915);
nor U6484 (N_6484,N_1766,N_813);
or U6485 (N_6485,N_2016,N_3551);
or U6486 (N_6486,N_2883,N_4390);
nor U6487 (N_6487,N_2866,N_2087);
or U6488 (N_6488,N_3984,N_3336);
and U6489 (N_6489,N_2859,N_1000);
nand U6490 (N_6490,N_1710,N_4104);
or U6491 (N_6491,N_4827,N_3289);
and U6492 (N_6492,N_3114,N_716);
or U6493 (N_6493,N_1503,N_4733);
nor U6494 (N_6494,N_4812,N_2293);
nand U6495 (N_6495,N_3483,N_2510);
nand U6496 (N_6496,N_4651,N_512);
nor U6497 (N_6497,N_1745,N_3531);
nor U6498 (N_6498,N_2470,N_456);
and U6499 (N_6499,N_2790,N_4609);
xor U6500 (N_6500,N_4630,N_2404);
or U6501 (N_6501,N_843,N_3283);
nand U6502 (N_6502,N_1747,N_4293);
and U6503 (N_6503,N_110,N_4340);
and U6504 (N_6504,N_2401,N_1661);
and U6505 (N_6505,N_1490,N_3511);
nand U6506 (N_6506,N_1413,N_516);
nor U6507 (N_6507,N_538,N_1170);
nand U6508 (N_6508,N_4615,N_3589);
or U6509 (N_6509,N_1143,N_3750);
and U6510 (N_6510,N_2084,N_3830);
xor U6511 (N_6511,N_2301,N_4385);
xor U6512 (N_6512,N_1228,N_422);
and U6513 (N_6513,N_3385,N_211);
or U6514 (N_6514,N_1775,N_4344);
nand U6515 (N_6515,N_2320,N_1882);
and U6516 (N_6516,N_158,N_4409);
xor U6517 (N_6517,N_1123,N_1555);
xor U6518 (N_6518,N_575,N_1292);
and U6519 (N_6519,N_283,N_943);
or U6520 (N_6520,N_3631,N_4877);
and U6521 (N_6521,N_355,N_4653);
xnor U6522 (N_6522,N_1066,N_1923);
nand U6523 (N_6523,N_173,N_3324);
nand U6524 (N_6524,N_2717,N_4048);
or U6525 (N_6525,N_1158,N_1162);
or U6526 (N_6526,N_4855,N_2778);
or U6527 (N_6527,N_1651,N_1768);
nor U6528 (N_6528,N_728,N_2796);
xor U6529 (N_6529,N_1541,N_3526);
and U6530 (N_6530,N_970,N_508);
and U6531 (N_6531,N_1669,N_3646);
or U6532 (N_6532,N_2144,N_1778);
nor U6533 (N_6533,N_4445,N_641);
nand U6534 (N_6534,N_4328,N_77);
or U6535 (N_6535,N_1022,N_1199);
or U6536 (N_6536,N_2323,N_4729);
and U6537 (N_6537,N_2199,N_328);
nor U6538 (N_6538,N_4930,N_3144);
nand U6539 (N_6539,N_3819,N_2564);
xor U6540 (N_6540,N_2459,N_3699);
nand U6541 (N_6541,N_4604,N_1355);
nand U6542 (N_6542,N_2987,N_4895);
xnor U6543 (N_6543,N_4252,N_600);
or U6544 (N_6544,N_627,N_3226);
nand U6545 (N_6545,N_4448,N_746);
or U6546 (N_6546,N_583,N_2905);
and U6547 (N_6547,N_3429,N_1132);
nor U6548 (N_6548,N_101,N_798);
nor U6549 (N_6549,N_3693,N_3955);
or U6550 (N_6550,N_3628,N_433);
or U6551 (N_6551,N_4816,N_2412);
nor U6552 (N_6552,N_3176,N_1077);
or U6553 (N_6553,N_4430,N_382);
nand U6554 (N_6554,N_2128,N_11);
and U6555 (N_6555,N_1620,N_1535);
nor U6556 (N_6556,N_68,N_2053);
nor U6557 (N_6557,N_3720,N_2167);
nor U6558 (N_6558,N_4308,N_2919);
or U6559 (N_6559,N_3953,N_4755);
xnor U6560 (N_6560,N_1474,N_3241);
xnor U6561 (N_6561,N_1225,N_2252);
and U6562 (N_6562,N_303,N_4189);
nor U6563 (N_6563,N_308,N_4955);
nand U6564 (N_6564,N_2771,N_2858);
and U6565 (N_6565,N_820,N_172);
nand U6566 (N_6566,N_594,N_1520);
nor U6567 (N_6567,N_4218,N_1102);
and U6568 (N_6568,N_3767,N_1929);
or U6569 (N_6569,N_1516,N_4316);
nand U6570 (N_6570,N_4182,N_2522);
xor U6571 (N_6571,N_4037,N_2765);
or U6572 (N_6572,N_2285,N_1890);
nor U6573 (N_6573,N_4752,N_3133);
or U6574 (N_6574,N_1142,N_2838);
nor U6575 (N_6575,N_443,N_2331);
xor U6576 (N_6576,N_2219,N_687);
nor U6577 (N_6577,N_1014,N_3522);
xnor U6578 (N_6578,N_1539,N_3132);
xnor U6579 (N_6579,N_395,N_2895);
nand U6580 (N_6580,N_2646,N_224);
or U6581 (N_6581,N_981,N_1259);
nand U6582 (N_6582,N_2102,N_1126);
or U6583 (N_6583,N_4082,N_3737);
nand U6584 (N_6584,N_1335,N_3576);
xnor U6585 (N_6585,N_921,N_259);
xor U6586 (N_6586,N_675,N_4019);
xnor U6587 (N_6587,N_3557,N_2049);
nor U6588 (N_6588,N_4632,N_4093);
nand U6589 (N_6589,N_3307,N_1042);
nor U6590 (N_6590,N_4492,N_2494);
or U6591 (N_6591,N_2530,N_4634);
nand U6592 (N_6592,N_930,N_4988);
xnor U6593 (N_6593,N_2324,N_3678);
and U6594 (N_6594,N_2365,N_1895);
xor U6595 (N_6595,N_3419,N_4473);
or U6596 (N_6596,N_2094,N_1360);
and U6597 (N_6597,N_2968,N_4295);
nor U6598 (N_6598,N_2603,N_3350);
nor U6599 (N_6599,N_3936,N_204);
nor U6600 (N_6600,N_314,N_1465);
xnor U6601 (N_6601,N_1921,N_1559);
nand U6602 (N_6602,N_2292,N_2752);
xor U6603 (N_6603,N_4950,N_2410);
nand U6604 (N_6604,N_3519,N_4495);
and U6605 (N_6605,N_1712,N_1913);
xor U6606 (N_6606,N_4550,N_347);
nor U6607 (N_6607,N_399,N_2699);
xor U6608 (N_6608,N_534,N_67);
nor U6609 (N_6609,N_2793,N_4357);
nand U6610 (N_6610,N_126,N_4184);
and U6611 (N_6611,N_2517,N_745);
or U6612 (N_6612,N_4412,N_420);
xnor U6613 (N_6613,N_315,N_4858);
nand U6614 (N_6614,N_1846,N_4783);
nand U6615 (N_6615,N_3273,N_4391);
or U6616 (N_6616,N_2749,N_1784);
xor U6617 (N_6617,N_3108,N_2736);
or U6618 (N_6618,N_2695,N_547);
or U6619 (N_6619,N_2777,N_3798);
or U6620 (N_6620,N_3295,N_2986);
nand U6621 (N_6621,N_1935,N_4110);
or U6622 (N_6622,N_4524,N_4793);
xnor U6623 (N_6623,N_4926,N_4794);
nor U6624 (N_6624,N_3105,N_131);
and U6625 (N_6625,N_3068,N_2533);
xnor U6626 (N_6626,N_1301,N_3837);
xnor U6627 (N_6627,N_2985,N_966);
or U6628 (N_6628,N_134,N_1636);
or U6629 (N_6629,N_4452,N_2657);
nor U6630 (N_6630,N_712,N_2738);
or U6631 (N_6631,N_2367,N_1616);
nor U6632 (N_6632,N_388,N_3808);
and U6633 (N_6633,N_693,N_4666);
or U6634 (N_6634,N_887,N_3287);
nand U6635 (N_6635,N_4015,N_2804);
and U6636 (N_6636,N_1936,N_2737);
xor U6637 (N_6637,N_3609,N_1344);
and U6638 (N_6638,N_71,N_3774);
and U6639 (N_6639,N_47,N_543);
or U6640 (N_6640,N_4085,N_2513);
nand U6641 (N_6641,N_799,N_2453);
nand U6642 (N_6642,N_2489,N_1663);
or U6643 (N_6643,N_2389,N_3752);
nor U6644 (N_6644,N_392,N_4186);
xnor U6645 (N_6645,N_2896,N_307);
nand U6646 (N_6646,N_4101,N_432);
or U6647 (N_6647,N_4789,N_1330);
xnor U6648 (N_6648,N_2622,N_4255);
nand U6649 (N_6649,N_266,N_964);
or U6650 (N_6650,N_367,N_845);
nand U6651 (N_6651,N_327,N_2218);
and U6652 (N_6652,N_2881,N_4552);
xor U6653 (N_6653,N_4447,N_4424);
nor U6654 (N_6654,N_3706,N_316);
nor U6655 (N_6655,N_73,N_2431);
xor U6656 (N_6656,N_2729,N_4587);
nor U6657 (N_6657,N_3486,N_4517);
nand U6658 (N_6658,N_480,N_4369);
or U6659 (N_6659,N_3833,N_3425);
nor U6660 (N_6660,N_3834,N_1504);
nand U6661 (N_6661,N_925,N_684);
and U6662 (N_6662,N_3796,N_2135);
xnor U6663 (N_6663,N_1632,N_3641);
xnor U6664 (N_6664,N_3077,N_1670);
nand U6665 (N_6665,N_1447,N_3787);
or U6666 (N_6666,N_4795,N_4376);
and U6667 (N_6667,N_670,N_2643);
or U6668 (N_6668,N_3933,N_354);
xnor U6669 (N_6669,N_3694,N_4346);
xor U6670 (N_6670,N_3630,N_4034);
nand U6671 (N_6671,N_1813,N_3605);
or U6672 (N_6672,N_4558,N_4012);
or U6673 (N_6673,N_349,N_4386);
nand U6674 (N_6674,N_2787,N_4028);
nor U6675 (N_6675,N_2539,N_1960);
nor U6676 (N_6676,N_849,N_4846);
nand U6677 (N_6677,N_345,N_2893);
or U6678 (N_6678,N_1946,N_918);
xnor U6679 (N_6679,N_2250,N_875);
or U6680 (N_6680,N_528,N_2764);
xor U6681 (N_6681,N_3115,N_4962);
and U6682 (N_6682,N_2063,N_2384);
nand U6683 (N_6683,N_995,N_4309);
xor U6684 (N_6684,N_1587,N_898);
or U6685 (N_6685,N_332,N_1455);
nand U6686 (N_6686,N_1628,N_1852);
and U6687 (N_6687,N_4302,N_1601);
nor U6688 (N_6688,N_957,N_1605);
nand U6689 (N_6689,N_1205,N_4206);
nand U6690 (N_6690,N_58,N_4695);
nor U6691 (N_6691,N_4347,N_4003);
nor U6692 (N_6692,N_3236,N_2317);
or U6693 (N_6693,N_601,N_385);
and U6694 (N_6694,N_1974,N_1099);
nand U6695 (N_6695,N_3529,N_1577);
xor U6696 (N_6696,N_1915,N_2995);
and U6697 (N_6697,N_2082,N_4725);
and U6698 (N_6698,N_3807,N_3749);
and U6699 (N_6699,N_3299,N_2498);
and U6700 (N_6700,N_3795,N_1674);
xor U6701 (N_6701,N_3826,N_3134);
xnor U6702 (N_6702,N_243,N_4245);
and U6703 (N_6703,N_572,N_4664);
or U6704 (N_6704,N_329,N_3820);
nor U6705 (N_6705,N_1873,N_4151);
nand U6706 (N_6706,N_1409,N_1725);
nor U6707 (N_6707,N_1437,N_4235);
nand U6708 (N_6708,N_1297,N_2220);
or U6709 (N_6709,N_1241,N_3237);
and U6710 (N_6710,N_3370,N_3741);
nand U6711 (N_6711,N_1600,N_1284);
xor U6712 (N_6712,N_2150,N_3096);
xor U6713 (N_6713,N_1453,N_922);
nand U6714 (N_6714,N_1306,N_2435);
and U6715 (N_6715,N_1135,N_4433);
nand U6716 (N_6716,N_1197,N_2211);
nand U6717 (N_6717,N_1831,N_2116);
and U6718 (N_6718,N_177,N_1471);
xnor U6719 (N_6719,N_3192,N_2612);
xnor U6720 (N_6720,N_1943,N_78);
and U6721 (N_6721,N_3484,N_2994);
or U6722 (N_6722,N_44,N_3189);
xnor U6723 (N_6723,N_4063,N_810);
nor U6724 (N_6724,N_2560,N_1963);
nor U6725 (N_6725,N_2083,N_2743);
xnor U6726 (N_6726,N_972,N_30);
and U6727 (N_6727,N_4882,N_4398);
and U6728 (N_6728,N_2333,N_4130);
or U6729 (N_6729,N_4995,N_3932);
nand U6730 (N_6730,N_2488,N_2372);
or U6731 (N_6731,N_462,N_3858);
nand U6732 (N_6732,N_3743,N_2719);
and U6733 (N_6733,N_2876,N_4002);
or U6734 (N_6734,N_3264,N_219);
and U6735 (N_6735,N_2183,N_2694);
nand U6736 (N_6736,N_2889,N_4120);
nand U6737 (N_6737,N_682,N_4529);
nand U6738 (N_6738,N_589,N_3084);
nand U6739 (N_6739,N_3012,N_438);
xnor U6740 (N_6740,N_1810,N_2630);
nand U6741 (N_6741,N_192,N_3508);
and U6742 (N_6742,N_4671,N_1202);
and U6743 (N_6743,N_1728,N_440);
or U6744 (N_6744,N_655,N_3822);
nor U6745 (N_6745,N_2617,N_4667);
and U6746 (N_6746,N_4611,N_337);
nor U6747 (N_6747,N_3332,N_291);
nand U6748 (N_6748,N_734,N_386);
or U6749 (N_6749,N_904,N_3213);
xor U6750 (N_6750,N_878,N_4086);
nor U6751 (N_6751,N_1694,N_3810);
xnor U6752 (N_6752,N_4321,N_1972);
nor U6753 (N_6753,N_3368,N_413);
or U6754 (N_6754,N_2928,N_4162);
and U6755 (N_6755,N_4395,N_4055);
nand U6756 (N_6756,N_832,N_1433);
or U6757 (N_6757,N_4067,N_3191);
or U6758 (N_6758,N_3078,N_3781);
nand U6759 (N_6759,N_2195,N_1619);
nand U6760 (N_6760,N_615,N_1432);
nand U6761 (N_6761,N_14,N_212);
xnor U6762 (N_6762,N_1426,N_3981);
nor U6763 (N_6763,N_4839,N_3685);
or U6764 (N_6764,N_1631,N_2954);
and U6765 (N_6765,N_542,N_3973);
or U6766 (N_6766,N_2535,N_1498);
nor U6767 (N_6767,N_479,N_4024);
and U6768 (N_6768,N_4265,N_4798);
and U6769 (N_6769,N_2104,N_715);
or U6770 (N_6770,N_230,N_1213);
and U6771 (N_6771,N_3517,N_3175);
xor U6772 (N_6772,N_2026,N_213);
nand U6773 (N_6773,N_3886,N_3540);
xnor U6774 (N_6774,N_3294,N_902);
and U6775 (N_6775,N_2415,N_4762);
or U6776 (N_6776,N_3944,N_566);
xor U6777 (N_6777,N_3245,N_2254);
nand U6778 (N_6778,N_2524,N_4563);
xnor U6779 (N_6779,N_4173,N_1549);
or U6780 (N_6780,N_2812,N_1083);
or U6781 (N_6781,N_4470,N_176);
and U6782 (N_6782,N_22,N_3758);
and U6783 (N_6783,N_1475,N_2690);
xor U6784 (N_6784,N_2998,N_348);
xnor U6785 (N_6785,N_2281,N_1534);
xnor U6786 (N_6786,N_2111,N_1235);
or U6787 (N_6787,N_4289,N_4676);
nor U6788 (N_6788,N_1757,N_2924);
xnor U6789 (N_6789,N_1092,N_4479);
and U6790 (N_6790,N_2363,N_311);
nor U6791 (N_6791,N_3100,N_3841);
nand U6792 (N_6792,N_317,N_3625);
or U6793 (N_6793,N_736,N_436);
and U6794 (N_6794,N_661,N_4530);
nor U6795 (N_6795,N_2172,N_1957);
and U6796 (N_6796,N_3709,N_16);
xor U6797 (N_6797,N_3762,N_4692);
xor U6798 (N_6798,N_1797,N_4661);
or U6799 (N_6799,N_2593,N_4871);
nand U6800 (N_6800,N_560,N_836);
and U6801 (N_6801,N_3488,N_3376);
nand U6802 (N_6802,N_4977,N_2126);
or U6803 (N_6803,N_735,N_346);
xor U6804 (N_6804,N_115,N_4420);
nor U6805 (N_6805,N_2165,N_636);
or U6806 (N_6806,N_1563,N_2481);
and U6807 (N_6807,N_1134,N_2661);
xor U6808 (N_6808,N_924,N_962);
or U6809 (N_6809,N_908,N_2607);
xnor U6810 (N_6810,N_3902,N_4212);
xor U6811 (N_6811,N_2652,N_521);
and U6812 (N_6812,N_2877,N_1738);
and U6813 (N_6813,N_467,N_882);
and U6814 (N_6814,N_4527,N_408);
xnor U6815 (N_6815,N_1456,N_1678);
and U6816 (N_6816,N_1597,N_26);
nand U6817 (N_6817,N_1633,N_1883);
nor U6818 (N_6818,N_4711,N_2064);
xnor U6819 (N_6819,N_3536,N_2917);
nand U6820 (N_6820,N_2970,N_4593);
and U6821 (N_6821,N_1062,N_3563);
and U6822 (N_6822,N_614,N_2727);
xnor U6823 (N_6823,N_1229,N_872);
and U6824 (N_6824,N_1026,N_2818);
or U6825 (N_6825,N_3884,N_3552);
nor U6826 (N_6826,N_3579,N_196);
xnor U6827 (N_6827,N_2224,N_3482);
nor U6828 (N_6828,N_1552,N_814);
nor U6829 (N_6829,N_3868,N_1436);
nand U6830 (N_6830,N_1223,N_2454);
nand U6831 (N_6831,N_2419,N_2976);
and U6832 (N_6832,N_3357,N_116);
nand U6833 (N_6833,N_4868,N_3276);
nor U6834 (N_6834,N_2303,N_153);
nand U6835 (N_6835,N_2005,N_2837);
or U6836 (N_6836,N_4403,N_913);
nor U6837 (N_6837,N_1706,N_1641);
xor U6838 (N_6838,N_861,N_4734);
nand U6839 (N_6839,N_2505,N_4826);
and U6840 (N_6840,N_4784,N_2821);
and U6841 (N_6841,N_514,N_762);
or U6842 (N_6842,N_3985,N_2019);
xnor U6843 (N_6843,N_4239,N_1368);
or U6844 (N_6844,N_2580,N_984);
and U6845 (N_6845,N_4780,N_3205);
and U6846 (N_6846,N_304,N_2377);
nand U6847 (N_6847,N_2508,N_700);
or U6848 (N_6848,N_377,N_632);
or U6849 (N_6849,N_3395,N_1480);
or U6850 (N_6850,N_2484,N_4225);
and U6851 (N_6851,N_1209,N_4372);
xor U6852 (N_6852,N_2031,N_621);
or U6853 (N_6853,N_313,N_4944);
nor U6854 (N_6854,N_3030,N_3939);
or U6855 (N_6855,N_65,N_496);
nor U6856 (N_6856,N_2123,N_4698);
xnor U6857 (N_6857,N_4299,N_829);
and U6858 (N_6858,N_1193,N_3023);
nand U6859 (N_6859,N_4548,N_1792);
nand U6860 (N_6860,N_3333,N_1187);
or U6861 (N_6861,N_1715,N_244);
and U6862 (N_6862,N_3559,N_3914);
and U6863 (N_6863,N_4004,N_2021);
or U6864 (N_6864,N_4488,N_3218);
or U6865 (N_6865,N_2163,N_4908);
and U6866 (N_6866,N_3045,N_461);
nand U6867 (N_6867,N_3073,N_767);
and U6868 (N_6868,N_4468,N_3119);
nor U6869 (N_6869,N_3675,N_419);
xnor U6870 (N_6870,N_3451,N_1908);
and U6871 (N_6871,N_2009,N_302);
xor U6872 (N_6872,N_261,N_3022);
nor U6873 (N_6873,N_363,N_3188);
nor U6874 (N_6874,N_37,N_4750);
and U6875 (N_6875,N_1798,N_227);
nand U6876 (N_6876,N_1819,N_217);
nor U6877 (N_6877,N_369,N_717);
nand U6878 (N_6878,N_4797,N_293);
and U6879 (N_6879,N_1796,N_4314);
xnor U6880 (N_6880,N_3321,N_3398);
and U6881 (N_6881,N_1794,N_758);
or U6882 (N_6882,N_2577,N_102);
nand U6883 (N_6883,N_4187,N_374);
nand U6884 (N_6884,N_2990,N_1058);
and U6885 (N_6885,N_301,N_1429);
nor U6886 (N_6886,N_1769,N_1578);
xor U6887 (N_6887,N_2629,N_2800);
nor U6888 (N_6888,N_2773,N_742);
and U6889 (N_6889,N_4999,N_1390);
and U6890 (N_6890,N_4041,N_3874);
nand U6891 (N_6891,N_3857,N_1603);
or U6892 (N_6892,N_2712,N_4901);
xnor U6893 (N_6893,N_1374,N_613);
xor U6894 (N_6894,N_4740,N_1740);
xor U6895 (N_6895,N_2187,N_378);
nand U6896 (N_6896,N_3069,N_3745);
nand U6897 (N_6897,N_3788,N_4989);
nor U6898 (N_6898,N_3279,N_3344);
or U6899 (N_6899,N_3998,N_2907);
nand U6900 (N_6900,N_1789,N_975);
xor U6901 (N_6901,N_777,N_4059);
nor U6902 (N_6902,N_2070,N_2020);
nand U6903 (N_6903,N_626,N_1045);
or U6904 (N_6904,N_2434,N_946);
xnor U6905 (N_6905,N_4205,N_3676);
nor U6906 (N_6906,N_2815,N_414);
nand U6907 (N_6907,N_3923,N_551);
nor U6908 (N_6908,N_482,N_1734);
xor U6909 (N_6909,N_4327,N_2813);
nor U6910 (N_6910,N_3090,N_3384);
nand U6911 (N_6911,N_32,N_3052);
and U6912 (N_6912,N_2177,N_2634);
or U6913 (N_6913,N_3608,N_450);
nor U6914 (N_6914,N_2340,N_3770);
nor U6915 (N_6915,N_2000,N_2875);
and U6916 (N_6916,N_3950,N_2059);
nand U6917 (N_6917,N_2011,N_130);
and U6918 (N_6918,N_2550,N_3919);
nor U6919 (N_6919,N_973,N_3444);
nand U6920 (N_6920,N_1183,N_1434);
or U6921 (N_6921,N_3956,N_3654);
or U6922 (N_6922,N_396,N_1855);
and U6923 (N_6923,N_3930,N_1282);
or U6924 (N_6924,N_491,N_4350);
nand U6925 (N_6925,N_3342,N_3707);
and U6926 (N_6926,N_3889,N_1598);
nor U6927 (N_6927,N_2949,N_744);
xnor U6928 (N_6928,N_3623,N_290);
xnor U6929 (N_6929,N_2230,N_1233);
and U6930 (N_6930,N_653,N_1369);
or U6931 (N_6931,N_85,N_4040);
nor U6932 (N_6932,N_1682,N_4273);
nand U6933 (N_6933,N_4538,N_2032);
xnor U6934 (N_6934,N_1111,N_45);
and U6935 (N_6935,N_4076,N_2518);
xnor U6936 (N_6936,N_1887,N_3658);
nor U6937 (N_6937,N_3247,N_1602);
and U6938 (N_6938,N_4927,N_4047);
or U6939 (N_6939,N_2446,N_2202);
nor U6940 (N_6940,N_2477,N_4948);
and U6941 (N_6941,N_2107,N_3542);
and U6942 (N_6942,N_1382,N_387);
and U6943 (N_6943,N_808,N_1420);
or U6944 (N_6944,N_4533,N_3573);
xor U6945 (N_6945,N_531,N_1699);
or U6946 (N_6946,N_2680,N_441);
nand U6947 (N_6947,N_2648,N_3509);
and U6948 (N_6948,N_428,N_1750);
and U6949 (N_6949,N_201,N_499);
nor U6950 (N_6950,N_4932,N_3424);
and U6951 (N_6951,N_2543,N_2378);
and U6952 (N_6952,N_2233,N_3477);
nand U6953 (N_6953,N_3199,N_1507);
nand U6954 (N_6954,N_478,N_4033);
nand U6955 (N_6955,N_2213,N_2829);
or U6956 (N_6956,N_639,N_770);
xor U6957 (N_6957,N_3271,N_1009);
xnor U6958 (N_6958,N_3061,N_1776);
or U6959 (N_6959,N_2864,N_2936);
nor U6960 (N_6960,N_3792,N_4399);
nand U6961 (N_6961,N_4202,N_2620);
and U6962 (N_6962,N_1317,N_978);
xnor U6963 (N_6963,N_4675,N_4180);
and U6964 (N_6964,N_3813,N_850);
nand U6965 (N_6965,N_1274,N_1853);
and U6966 (N_6966,N_3298,N_1435);
nand U6967 (N_6967,N_518,N_3824);
or U6968 (N_6968,N_3638,N_4785);
and U6969 (N_6969,N_3167,N_193);
or U6970 (N_6970,N_4074,N_1795);
xnor U6971 (N_6971,N_4155,N_1309);
and U6972 (N_6972,N_2601,N_4394);
xnor U6973 (N_6973,N_352,N_1019);
nor U6974 (N_6974,N_3854,N_4726);
nor U6975 (N_6975,N_730,N_3947);
nand U6976 (N_6976,N_1566,N_3814);
xor U6977 (N_6977,N_2592,N_3230);
and U6978 (N_6978,N_3400,N_2856);
or U6979 (N_6979,N_4442,N_152);
nand U6980 (N_6980,N_3616,N_2338);
nand U6981 (N_6981,N_280,N_4166);
and U6982 (N_6982,N_2015,N_4702);
nor U6983 (N_6983,N_3538,N_3761);
nand U6984 (N_6984,N_2473,N_690);
or U6985 (N_6985,N_1975,N_3626);
xor U6986 (N_6986,N_1016,N_4406);
nand U6987 (N_6987,N_282,N_1896);
nor U6988 (N_6988,N_218,N_2381);
or U6989 (N_6989,N_4348,N_4663);
or U6990 (N_6990,N_1877,N_2322);
or U6991 (N_6991,N_1247,N_1332);
nand U6992 (N_6992,N_4771,N_3386);
or U6993 (N_6993,N_2091,N_61);
nor U6994 (N_6994,N_417,N_3238);
or U6995 (N_6995,N_4259,N_1131);
xnor U6996 (N_6996,N_4443,N_4071);
xor U6997 (N_6997,N_4248,N_2912);
or U6998 (N_6998,N_1806,N_4056);
and U6999 (N_6999,N_4570,N_3194);
or U7000 (N_7000,N_2952,N_3582);
or U7001 (N_7001,N_2466,N_1848);
nor U7002 (N_7002,N_948,N_3846);
nor U7003 (N_7003,N_271,N_2570);
nor U7004 (N_7004,N_3635,N_1476);
nand U7005 (N_7005,N_2692,N_3481);
nand U7006 (N_7006,N_2071,N_4620);
nor U7007 (N_7007,N_3259,N_1361);
nor U7008 (N_7008,N_1265,N_3967);
nor U7009 (N_7009,N_997,N_1954);
nor U7010 (N_7010,N_3549,N_2456);
xor U7011 (N_7011,N_2089,N_4983);
nor U7012 (N_7012,N_3079,N_2534);
nand U7013 (N_7013,N_1393,N_2816);
or U7014 (N_7014,N_154,N_2214);
or U7015 (N_7015,N_2760,N_4233);
or U7016 (N_7016,N_3364,N_4160);
or U7017 (N_7017,N_2047,N_1462);
or U7018 (N_7018,N_2637,N_49);
nand U7019 (N_7019,N_2655,N_2911);
or U7020 (N_7020,N_2581,N_571);
or U7021 (N_7021,N_1639,N_3490);
or U7022 (N_7022,N_2353,N_2359);
or U7023 (N_7023,N_697,N_1844);
and U7024 (N_7024,N_1826,N_2937);
xor U7025 (N_7025,N_4585,N_2780);
nor U7026 (N_7026,N_4477,N_3996);
xnor U7027 (N_7027,N_983,N_1283);
and U7028 (N_7028,N_1138,N_238);
xnor U7029 (N_7029,N_1275,N_2447);
and U7030 (N_7030,N_3290,N_2647);
nor U7031 (N_7031,N_4010,N_1707);
xor U7032 (N_7032,N_3615,N_3732);
nor U7033 (N_7033,N_1080,N_3470);
and U7034 (N_7034,N_3420,N_3593);
xor U7035 (N_7035,N_540,N_3934);
nor U7036 (N_7036,N_3293,N_936);
nor U7037 (N_7037,N_4238,N_3124);
or U7038 (N_7038,N_1659,N_330);
or U7039 (N_7039,N_3744,N_412);
and U7040 (N_7040,N_3771,N_4586);
nor U7041 (N_7041,N_2460,N_2143);
nor U7042 (N_7042,N_652,N_2411);
or U7043 (N_7043,N_4885,N_657);
nor U7044 (N_7044,N_3491,N_4605);
or U7045 (N_7045,N_1672,N_4525);
and U7046 (N_7046,N_4721,N_1404);
xor U7047 (N_7047,N_2436,N_1141);
nand U7048 (N_7048,N_2179,N_4665);
and U7049 (N_7049,N_4788,N_4237);
or U7050 (N_7050,N_1006,N_4759);
xor U7051 (N_7051,N_1851,N_2421);
xor U7052 (N_7052,N_1446,N_4122);
or U7053 (N_7053,N_3320,N_3217);
and U7054 (N_7054,N_1239,N_1976);
and U7055 (N_7055,N_2651,N_3581);
or U7056 (N_7056,N_4050,N_4061);
xnor U7057 (N_7057,N_2627,N_425);
nand U7058 (N_7058,N_1716,N_727);
or U7059 (N_7059,N_3315,N_665);
nand U7060 (N_7060,N_4282,N_4516);
xnor U7061 (N_7061,N_4383,N_2205);
and U7062 (N_7062,N_129,N_617);
or U7063 (N_7063,N_1968,N_741);
nor U7064 (N_7064,N_4502,N_2916);
nor U7065 (N_7065,N_3913,N_297);
and U7066 (N_7066,N_4515,N_2978);
nand U7067 (N_7067,N_2619,N_548);
xnor U7068 (N_7068,N_4860,N_4467);
or U7069 (N_7069,N_4964,N_449);
xnor U7070 (N_7070,N_1990,N_4751);
xnor U7071 (N_7071,N_1367,N_3698);
xnor U7072 (N_7072,N_4841,N_1713);
nor U7073 (N_7073,N_2642,N_4217);
xnor U7074 (N_7074,N_1079,N_4176);
or U7075 (N_7075,N_1184,N_2566);
nand U7076 (N_7076,N_4057,N_4573);
xnor U7077 (N_7077,N_1868,N_4654);
nor U7078 (N_7078,N_3328,N_4911);
xnor U7079 (N_7079,N_2175,N_1773);
xor U7080 (N_7080,N_4807,N_4640);
nor U7081 (N_7081,N_2715,N_254);
nor U7082 (N_7082,N_2547,N_1864);
nor U7083 (N_7083,N_2420,N_3899);
or U7084 (N_7084,N_226,N_4095);
and U7085 (N_7085,N_4351,N_4058);
nor U7086 (N_7086,N_2999,N_1771);
nand U7087 (N_7087,N_1366,N_2346);
and U7088 (N_7088,N_84,N_2741);
nor U7089 (N_7089,N_599,N_1981);
or U7090 (N_7090,N_1737,N_3089);
xnor U7091 (N_7091,N_647,N_381);
nand U7092 (N_7092,N_4354,N_3417);
nand U7093 (N_7093,N_2033,N_4522);
and U7094 (N_7094,N_2439,N_4125);
xor U7095 (N_7095,N_1630,N_4499);
nand U7096 (N_7096,N_1787,N_3875);
nand U7097 (N_7097,N_4153,N_3080);
or U7098 (N_7098,N_3407,N_2139);
nor U7099 (N_7099,N_2416,N_3928);
and U7100 (N_7100,N_2759,N_928);
and U7101 (N_7101,N_1400,N_4228);
nand U7102 (N_7102,N_1742,N_3138);
nor U7103 (N_7103,N_593,N_494);
nor U7104 (N_7104,N_3763,N_2222);
xor U7105 (N_7105,N_4656,N_3312);
and U7106 (N_7106,N_356,N_1181);
and U7107 (N_7107,N_4216,N_642);
xnor U7108 (N_7108,N_2921,N_565);
xor U7109 (N_7109,N_191,N_3251);
nand U7110 (N_7110,N_1096,N_1660);
and U7111 (N_7111,N_2266,N_3116);
nor U7112 (N_7112,N_3058,N_4060);
nor U7113 (N_7113,N_106,N_4247);
xnor U7114 (N_7114,N_199,N_189);
or U7115 (N_7115,N_3494,N_3562);
xnor U7116 (N_7116,N_3547,N_233);
nor U7117 (N_7117,N_4170,N_4924);
nand U7118 (N_7118,N_1512,N_4590);
nand U7119 (N_7119,N_2120,N_1421);
nand U7120 (N_7120,N_4555,N_822);
nor U7121 (N_7121,N_2469,N_1109);
or U7122 (N_7122,N_1039,N_1569);
nor U7123 (N_7123,N_4616,N_1191);
xnor U7124 (N_7124,N_3725,N_4231);
or U7125 (N_7125,N_2491,N_83);
or U7126 (N_7126,N_28,N_1004);
nor U7127 (N_7127,N_2611,N_59);
nand U7128 (N_7128,N_4175,N_171);
or U7129 (N_7129,N_426,N_3222);
nand U7130 (N_7130,N_4678,N_709);
and U7131 (N_7131,N_3141,N_1151);
nand U7132 (N_7132,N_3703,N_4591);
and U7133 (N_7133,N_2045,N_3640);
nor U7134 (N_7134,N_3997,N_1653);
or U7135 (N_7135,N_1358,N_4118);
nor U7136 (N_7136,N_471,N_677);
xor U7137 (N_7137,N_2739,N_1955);
and U7138 (N_7138,N_2835,N_2277);
xor U7139 (N_7139,N_100,N_4504);
nor U7140 (N_7140,N_4150,N_4703);
xnor U7141 (N_7141,N_2950,N_1082);
or U7142 (N_7142,N_2394,N_4717);
nand U7143 (N_7143,N_1211,N_13);
nand U7144 (N_7144,N_4757,N_686);
xor U7145 (N_7145,N_3577,N_3308);
nand U7146 (N_7146,N_3921,N_2115);
xnor U7147 (N_7147,N_2554,N_4912);
nand U7148 (N_7148,N_4852,N_3688);
or U7149 (N_7149,N_210,N_1530);
and U7150 (N_7150,N_4208,N_4179);
xnor U7151 (N_7151,N_411,N_3082);
nor U7152 (N_7152,N_3485,N_2512);
xor U7153 (N_7153,N_4367,N_2926);
xnor U7154 (N_7154,N_2146,N_2667);
nor U7155 (N_7155,N_3801,N_4673);
nand U7156 (N_7156,N_2080,N_3010);
or U7157 (N_7157,N_3687,N_2110);
nor U7158 (N_7158,N_929,N_998);
or U7159 (N_7159,N_2846,N_340);
nor U7160 (N_7160,N_4847,N_1781);
xnor U7161 (N_7161,N_4257,N_135);
nand U7162 (N_7162,N_1065,N_2445);
nor U7163 (N_7163,N_3016,N_4909);
nand U7164 (N_7164,N_522,N_3142);
xnor U7165 (N_7165,N_3204,N_825);
and U7166 (N_7166,N_1730,N_1638);
nand U7167 (N_7167,N_605,N_2072);
xor U7168 (N_7168,N_1048,N_333);
nor U7169 (N_7169,N_2463,N_1899);
and U7170 (N_7170,N_1147,N_1379);
xor U7171 (N_7171,N_323,N_1302);
nor U7172 (N_7172,N_1671,N_596);
xnor U7173 (N_7173,N_3975,N_1276);
nor U7174 (N_7174,N_1419,N_91);
nand U7175 (N_7175,N_2941,N_833);
nor U7176 (N_7176,N_235,N_2897);
or U7177 (N_7177,N_2742,N_1727);
xor U7178 (N_7178,N_1384,N_3367);
xnor U7179 (N_7179,N_4,N_4612);
nor U7180 (N_7180,N_4790,N_4718);
or U7181 (N_7181,N_4332,N_1479);
and U7182 (N_7182,N_4994,N_1145);
xnor U7183 (N_7183,N_749,N_4487);
xnor U7184 (N_7184,N_4723,N_944);
nor U7185 (N_7185,N_529,N_3596);
or U7186 (N_7186,N_2258,N_2405);
nand U7187 (N_7187,N_2332,N_477);
nor U7188 (N_7188,N_2345,N_2589);
or U7189 (N_7189,N_2681,N_2038);
and U7190 (N_7190,N_1903,N_2597);
or U7191 (N_7191,N_671,N_2158);
nand U7192 (N_7192,N_4510,N_4636);
nand U7193 (N_7193,N_2852,N_3870);
nor U7194 (N_7194,N_4498,N_1489);
nand U7195 (N_7195,N_2196,N_760);
nand U7196 (N_7196,N_3586,N_4631);
and U7197 (N_7197,N_1315,N_3469);
or U7198 (N_7198,N_968,N_4330);
and U7199 (N_7199,N_890,N_2495);
or U7200 (N_7200,N_1933,N_2903);
or U7201 (N_7201,N_3427,N_4970);
nand U7202 (N_7202,N_1525,N_4234);
nand U7203 (N_7203,N_680,N_4526);
nor U7204 (N_7204,N_82,N_383);
nand U7205 (N_7205,N_809,N_4732);
nand U7206 (N_7206,N_4875,N_1331);
or U7207 (N_7207,N_2930,N_1998);
nor U7208 (N_7208,N_3853,N_696);
nand U7209 (N_7209,N_1208,N_93);
and U7210 (N_7210,N_1703,N_4696);
xor U7211 (N_7211,N_4474,N_723);
nand U7212 (N_7212,N_539,N_3275);
nand U7213 (N_7213,N_817,N_595);
and U7214 (N_7214,N_4185,N_4131);
nor U7215 (N_7215,N_1553,N_1056);
and U7216 (N_7216,N_4209,N_3948);
and U7217 (N_7217,N_2065,N_801);
and U7218 (N_7218,N_4280,N_169);
nand U7219 (N_7219,N_2268,N_4873);
xnor U7220 (N_7220,N_2587,N_4117);
nand U7221 (N_7221,N_1385,N_3839);
and U7222 (N_7222,N_4659,N_442);
nor U7223 (N_7223,N_2106,N_4699);
nand U7224 (N_7224,N_4077,N_3883);
xnor U7225 (N_7225,N_2940,N_4764);
nand U7226 (N_7226,N_1606,N_4073);
nand U7227 (N_7227,N_4887,N_1043);
or U7228 (N_7228,N_1822,N_473);
or U7229 (N_7229,N_1212,N_4532);
or U7230 (N_7230,N_678,N_3127);
nor U7231 (N_7231,N_2502,N_1002);
and U7232 (N_7232,N_4799,N_3263);
nand U7233 (N_7233,N_1027,N_2839);
nor U7234 (N_7234,N_4787,N_2413);
nor U7235 (N_7235,N_1107,N_2354);
or U7236 (N_7236,N_2235,N_4577);
nand U7237 (N_7237,N_4014,N_1173);
and U7238 (N_7238,N_2312,N_527);
xor U7239 (N_7239,N_2927,N_1729);
and U7240 (N_7240,N_802,N_4691);
or U7241 (N_7241,N_4523,N_592);
or U7242 (N_7242,N_7,N_2327);
or U7243 (N_7243,N_350,N_4682);
or U7244 (N_7244,N_4105,N_515);
xnor U7245 (N_7245,N_3200,N_2099);
nand U7246 (N_7246,N_2850,N_4129);
or U7247 (N_7247,N_3460,N_1536);
or U7248 (N_7248,N_4923,N_90);
nand U7249 (N_7249,N_1166,N_3464);
nor U7250 (N_7250,N_4197,N_410);
nand U7251 (N_7251,N_2663,N_2806);
and U7252 (N_7252,N_2119,N_4193);
xor U7253 (N_7253,N_1410,N_886);
nor U7254 (N_7254,N_1254,N_1440);
xor U7255 (N_7255,N_3590,N_3498);
nor U7256 (N_7256,N_292,N_4773);
xor U7257 (N_7257,N_248,N_4848);
xnor U7258 (N_7258,N_942,N_2824);
nor U7259 (N_7259,N_2231,N_3335);
nand U7260 (N_7260,N_3401,N_2425);
nor U7261 (N_7261,N_4251,N_2623);
nor U7262 (N_7262,N_1898,N_320);
nand U7263 (N_7263,N_72,N_2847);
nor U7264 (N_7264,N_4436,N_3575);
and U7265 (N_7265,N_4198,N_1359);
and U7266 (N_7266,N_3453,N_469);
nand U7267 (N_7267,N_38,N_1194);
or U7268 (N_7268,N_1196,N_3152);
nor U7269 (N_7269,N_3995,N_1754);
xor U7270 (N_7270,N_1614,N_4973);
xor U7271 (N_7271,N_2029,N_3907);
nand U7272 (N_7272,N_794,N_255);
xnor U7273 (N_7273,N_1994,N_1608);
and U7274 (N_7274,N_3765,N_3730);
xor U7275 (N_7275,N_3681,N_4766);
nand U7276 (N_7276,N_3587,N_3789);
nor U7277 (N_7277,N_2808,N_1025);
or U7278 (N_7278,N_2732,N_4241);
or U7279 (N_7279,N_4387,N_1149);
or U7280 (N_7280,N_804,N_4974);
or U7281 (N_7281,N_2834,N_4084);
or U7282 (N_7282,N_4276,N_2319);
and U7283 (N_7283,N_1153,N_4838);
xnor U7284 (N_7284,N_3439,N_1662);
or U7285 (N_7285,N_4629,N_3043);
and U7286 (N_7286,N_2526,N_1237);
nor U7287 (N_7287,N_454,N_4069);
and U7288 (N_7288,N_180,N_1396);
nor U7289 (N_7289,N_4888,N_4476);
xnor U7290 (N_7290,N_3311,N_485);
xnor U7291 (N_7291,N_484,N_1753);
xnor U7292 (N_7292,N_2129,N_2662);
nor U7293 (N_7293,N_1372,N_1839);
or U7294 (N_7294,N_1791,N_2422);
nor U7295 (N_7295,N_1567,N_2909);
xnor U7296 (N_7296,N_1538,N_1735);
nand U7297 (N_7297,N_756,N_95);
or U7298 (N_7298,N_4451,N_4389);
nand U7299 (N_7299,N_2203,N_3291);
and U7300 (N_7300,N_3740,N_1108);
or U7301 (N_7301,N_4078,N_1997);
nor U7302 (N_7302,N_3351,N_4786);
or U7303 (N_7303,N_1800,N_2255);
nor U7304 (N_7304,N_4114,N_2461);
xnor U7305 (N_7305,N_69,N_3510);
nor U7306 (N_7306,N_865,N_4311);
xnor U7307 (N_7307,N_1656,N_905);
nand U7308 (N_7308,N_1342,N_2221);
xnor U7309 (N_7309,N_1609,N_643);
nand U7310 (N_7310,N_2753,N_1100);
nor U7311 (N_7311,N_2282,N_2148);
nand U7312 (N_7312,N_4491,N_996);
and U7313 (N_7313,N_1664,N_2174);
or U7314 (N_7314,N_1958,N_2557);
nor U7315 (N_7315,N_455,N_3179);
nor U7316 (N_7316,N_3624,N_200);
nor U7317 (N_7317,N_2556,N_431);
xor U7318 (N_7318,N_1926,N_4642);
or U7319 (N_7319,N_3280,N_3521);
nor U7320 (N_7320,N_4571,N_536);
and U7321 (N_7321,N_1175,N_4938);
nand U7322 (N_7322,N_4749,N_3015);
nor U7323 (N_7323,N_262,N_1060);
or U7324 (N_7324,N_3286,N_3014);
nor U7325 (N_7325,N_3354,N_451);
nand U7326 (N_7326,N_2962,N_3695);
nor U7327 (N_7327,N_1267,N_2991);
and U7328 (N_7328,N_4030,N_1375);
nand U7329 (N_7329,N_3823,N_1977);
or U7330 (N_7330,N_3316,N_3776);
or U7331 (N_7331,N_4158,N_3410);
or U7332 (N_7332,N_3102,N_2039);
and U7333 (N_7333,N_1945,N_4918);
xnor U7334 (N_7334,N_251,N_188);
xnor U7335 (N_7335,N_2373,N_4136);
and U7336 (N_7336,N_1937,N_3988);
nand U7337 (N_7337,N_143,N_1910);
and U7338 (N_7338,N_2946,N_2052);
nor U7339 (N_7339,N_4583,N_3614);
or U7340 (N_7340,N_1529,N_3239);
or U7341 (N_7341,N_1617,N_3943);
nand U7342 (N_7342,N_673,N_2792);
nor U7343 (N_7343,N_1281,N_2168);
nand U7344 (N_7344,N_2028,N_1253);
nand U7345 (N_7345,N_1055,N_789);
nand U7346 (N_7346,N_4844,N_1618);
xnor U7347 (N_7347,N_2414,N_3622);
nor U7348 (N_7348,N_360,N_4922);
and U7349 (N_7349,N_3713,N_577);
and U7350 (N_7350,N_4381,N_4519);
and U7351 (N_7351,N_4834,N_4144);
and U7352 (N_7352,N_1878,N_1508);
nand U7353 (N_7353,N_1515,N_2672);
or U7354 (N_7354,N_3880,N_4098);
or U7355 (N_7355,N_2105,N_1807);
or U7356 (N_7356,N_481,N_2010);
and U7357 (N_7357,N_4781,N_1860);
xnor U7358 (N_7358,N_1116,N_3979);
or U7359 (N_7359,N_3166,N_1733);
or U7360 (N_7360,N_761,N_2977);
xnor U7361 (N_7361,N_3775,N_3183);
and U7362 (N_7362,N_1902,N_229);
xor U7363 (N_7363,N_4694,N_1870);
nor U7364 (N_7364,N_775,N_2452);
or U7365 (N_7365,N_4971,N_3560);
and U7366 (N_7366,N_3405,N_3648);
nand U7367 (N_7367,N_1732,N_1391);
and U7368 (N_7368,N_2078,N_1979);
and U7369 (N_7369,N_3381,N_3009);
nor U7370 (N_7370,N_664,N_17);
or U7371 (N_7371,N_1320,N_3585);
or U7372 (N_7372,N_1272,N_222);
and U7373 (N_7373,N_2437,N_4290);
and U7374 (N_7374,N_4126,N_3784);
or U7375 (N_7375,N_748,N_525);
and U7376 (N_7376,N_1556,N_633);
nor U7377 (N_7377,N_2307,N_2660);
or U7378 (N_7378,N_1457,N_3665);
nor U7379 (N_7379,N_3358,N_3055);
xnor U7380 (N_7380,N_1150,N_1326);
xor U7381 (N_7381,N_530,N_2920);
nand U7382 (N_7382,N_806,N_1592);
nor U7383 (N_7383,N_1021,N_2653);
or U7384 (N_7384,N_3893,N_4910);
nor U7385 (N_7385,N_4035,N_598);
xnor U7386 (N_7386,N_3211,N_2360);
xor U7387 (N_7387,N_401,N_3456);
nor U7388 (N_7388,N_611,N_2376);
and U7389 (N_7389,N_4052,N_1467);
and U7390 (N_7390,N_2409,N_2012);
xor U7391 (N_7391,N_4207,N_1289);
xnor U7392 (N_7392,N_2665,N_2433);
nand U7393 (N_7393,N_3181,N_96);
nor U7394 (N_7394,N_1353,N_3431);
and U7395 (N_7395,N_2326,N_43);
or U7396 (N_7396,N_1717,N_2369);
nand U7397 (N_7397,N_3403,N_1485);
xnor U7398 (N_7398,N_4639,N_2142);
or U7399 (N_7399,N_1793,N_4889);
or U7400 (N_7400,N_3225,N_2939);
nor U7401 (N_7401,N_4320,N_1310);
nand U7402 (N_7402,N_3399,N_3649);
nand U7403 (N_7403,N_2245,N_4939);
and U7404 (N_7404,N_1483,N_4195);
xor U7405 (N_7405,N_3406,N_1575);
or U7406 (N_7406,N_4379,N_3897);
nor U7407 (N_7407,N_147,N_4183);
or U7408 (N_7408,N_4463,N_3591);
xnor U7409 (N_7409,N_768,N_2918);
or U7410 (N_7410,N_2786,N_2108);
nand U7411 (N_7411,N_4610,N_4714);
xnor U7412 (N_7412,N_464,N_698);
nand U7413 (N_7413,N_2018,N_3578);
nor U7414 (N_7414,N_4051,N_4355);
and U7415 (N_7415,N_3879,N_3842);
or U7416 (N_7416,N_1031,N_4662);
and U7417 (N_7417,N_4411,N_4107);
nand U7418 (N_7418,N_1155,N_920);
and U7419 (N_7419,N_3714,N_447);
and U7420 (N_7420,N_2055,N_2670);
nand U7421 (N_7421,N_3389,N_4414);
nand U7422 (N_7422,N_1560,N_4304);
or U7423 (N_7423,N_659,N_1314);
nand U7424 (N_7424,N_3856,N_3409);
nor U7425 (N_7425,N_3505,N_4501);
nor U7426 (N_7426,N_4083,N_2499);
xnor U7427 (N_7427,N_1985,N_1172);
nor U7428 (N_7428,N_1074,N_1611);
xnor U7429 (N_7429,N_2636,N_3532);
nand U7430 (N_7430,N_2074,N_3086);
nand U7431 (N_7431,N_2325,N_1174);
xnor U7432 (N_7432,N_4658,N_1035);
and U7433 (N_7433,N_1872,N_358);
or U7434 (N_7434,N_2666,N_3193);
nor U7435 (N_7435,N_586,N_1524);
and U7436 (N_7436,N_938,N_4201);
xnor U7437 (N_7437,N_1224,N_3738);
nand U7438 (N_7438,N_4690,N_2869);
xor U7439 (N_7439,N_3207,N_4996);
and U7440 (N_7440,N_1821,N_2337);
nand U7441 (N_7441,N_2261,N_2269);
nor U7442 (N_7442,N_573,N_2618);
and U7443 (N_7443,N_4222,N_3446);
and U7444 (N_7444,N_1629,N_3341);
or U7445 (N_7445,N_4334,N_1548);
xor U7446 (N_7446,N_3983,N_3349);
or U7447 (N_7447,N_1373,N_3657);
nor U7448 (N_7448,N_4296,N_3812);
or U7449 (N_7449,N_4456,N_1545);
or U7450 (N_7450,N_3093,N_1635);
nor U7451 (N_7451,N_373,N_3390);
xor U7452 (N_7452,N_1333,N_2348);
nor U7453 (N_7453,N_2633,N_4800);
or U7454 (N_7454,N_2830,N_910);
xnor U7455 (N_7455,N_1336,N_3106);
or U7456 (N_7456,N_3202,N_1970);
and U7457 (N_7457,N_3574,N_4102);
or U7458 (N_7458,N_155,N_4313);
and U7459 (N_7459,N_1786,N_3719);
or U7460 (N_7460,N_4016,N_2355);
nand U7461 (N_7461,N_1322,N_1825);
nor U7462 (N_7462,N_2956,N_2689);
xnor U7463 (N_7463,N_4374,N_3040);
or U7464 (N_7464,N_4589,N_818);
and U7465 (N_7465,N_1711,N_1177);
and U7466 (N_7466,N_1261,N_1513);
and U7467 (N_7467,N_2565,N_2973);
or U7468 (N_7468,N_4286,N_2632);
xnor U7469 (N_7469,N_1927,N_2014);
or U7470 (N_7470,N_581,N_120);
nand U7471 (N_7471,N_483,N_4804);
nor U7472 (N_7472,N_4842,N_4972);
nand U7473 (N_7473,N_324,N_1708);
or U7474 (N_7474,N_253,N_3153);
nand U7475 (N_7475,N_1445,N_3428);
nand U7476 (N_7476,N_2112,N_353);
xnor U7477 (N_7477,N_1094,N_776);
or U7478 (N_7478,N_3851,N_1227);
nand U7479 (N_7479,N_3266,N_1468);
or U7480 (N_7480,N_99,N_880);
and U7481 (N_7481,N_305,N_1607);
nand U7482 (N_7482,N_4435,N_122);
nand U7483 (N_7483,N_2975,N_3232);
nand U7484 (N_7484,N_362,N_2223);
nor U7485 (N_7485,N_1982,N_541);
and U7486 (N_7486,N_2136,N_3992);
and U7487 (N_7487,N_2217,N_2496);
xnor U7488 (N_7488,N_935,N_858);
and U7489 (N_7489,N_623,N_1273);
and U7490 (N_7490,N_3000,N_3003);
or U7491 (N_7491,N_4081,N_3711);
nor U7492 (N_7492,N_4719,N_2027);
or U7493 (N_7493,N_2002,N_2500);
and U7494 (N_7494,N_3757,N_1152);
nand U7495 (N_7495,N_3920,N_3091);
or U7496 (N_7496,N_2426,N_1032);
nor U7497 (N_7497,N_4169,N_3136);
and U7498 (N_7498,N_1300,N_3567);
nand U7499 (N_7499,N_2191,N_3448);
nand U7500 (N_7500,N_1604,N_1526);
and U7501 (N_7501,N_1347,N_4077);
and U7502 (N_7502,N_3812,N_770);
xnor U7503 (N_7503,N_664,N_929);
nor U7504 (N_7504,N_2021,N_3376);
nor U7505 (N_7505,N_4740,N_1110);
nor U7506 (N_7506,N_2247,N_3667);
nor U7507 (N_7507,N_568,N_3104);
xor U7508 (N_7508,N_1138,N_4401);
nand U7509 (N_7509,N_354,N_4365);
nand U7510 (N_7510,N_1277,N_1663);
nand U7511 (N_7511,N_1312,N_271);
nand U7512 (N_7512,N_3096,N_4683);
or U7513 (N_7513,N_3781,N_2788);
or U7514 (N_7514,N_57,N_1755);
nor U7515 (N_7515,N_741,N_3688);
or U7516 (N_7516,N_1625,N_2355);
nand U7517 (N_7517,N_4920,N_3243);
and U7518 (N_7518,N_3782,N_3457);
or U7519 (N_7519,N_4436,N_3531);
nor U7520 (N_7520,N_4322,N_1906);
nand U7521 (N_7521,N_770,N_3809);
nand U7522 (N_7522,N_125,N_2243);
xnor U7523 (N_7523,N_593,N_401);
nor U7524 (N_7524,N_3875,N_3973);
or U7525 (N_7525,N_653,N_1391);
xor U7526 (N_7526,N_4839,N_1002);
or U7527 (N_7527,N_2680,N_2325);
and U7528 (N_7528,N_872,N_167);
xnor U7529 (N_7529,N_2174,N_2768);
nor U7530 (N_7530,N_1946,N_1201);
and U7531 (N_7531,N_2671,N_2898);
nor U7532 (N_7532,N_4141,N_3710);
nor U7533 (N_7533,N_562,N_912);
xor U7534 (N_7534,N_2732,N_2075);
or U7535 (N_7535,N_3151,N_4136);
nand U7536 (N_7536,N_313,N_4927);
and U7537 (N_7537,N_2232,N_4576);
nand U7538 (N_7538,N_666,N_538);
and U7539 (N_7539,N_4260,N_1995);
and U7540 (N_7540,N_2183,N_4334);
or U7541 (N_7541,N_1814,N_2291);
nor U7542 (N_7542,N_88,N_4053);
and U7543 (N_7543,N_4636,N_1388);
nand U7544 (N_7544,N_4461,N_4540);
and U7545 (N_7545,N_3711,N_515);
and U7546 (N_7546,N_1243,N_3959);
or U7547 (N_7547,N_4949,N_3015);
and U7548 (N_7548,N_344,N_1968);
nor U7549 (N_7549,N_3298,N_3464);
or U7550 (N_7550,N_697,N_4667);
nor U7551 (N_7551,N_4844,N_2947);
xnor U7552 (N_7552,N_1124,N_3698);
or U7553 (N_7553,N_1569,N_3222);
nor U7554 (N_7554,N_4608,N_1337);
or U7555 (N_7555,N_3765,N_189);
or U7556 (N_7556,N_2729,N_3072);
xor U7557 (N_7557,N_3843,N_4464);
xnor U7558 (N_7558,N_1104,N_2004);
nand U7559 (N_7559,N_4211,N_1460);
or U7560 (N_7560,N_3964,N_3787);
xnor U7561 (N_7561,N_3101,N_1141);
and U7562 (N_7562,N_1610,N_1140);
xnor U7563 (N_7563,N_3443,N_2971);
nor U7564 (N_7564,N_947,N_2937);
xor U7565 (N_7565,N_1697,N_3382);
nor U7566 (N_7566,N_4796,N_256);
and U7567 (N_7567,N_4189,N_296);
xnor U7568 (N_7568,N_2077,N_1855);
xor U7569 (N_7569,N_2635,N_3704);
and U7570 (N_7570,N_1883,N_2268);
and U7571 (N_7571,N_2884,N_888);
and U7572 (N_7572,N_2882,N_1805);
nor U7573 (N_7573,N_2,N_4017);
and U7574 (N_7574,N_4747,N_183);
or U7575 (N_7575,N_1998,N_1245);
nor U7576 (N_7576,N_3392,N_2571);
nand U7577 (N_7577,N_3358,N_609);
or U7578 (N_7578,N_3019,N_2242);
nand U7579 (N_7579,N_1802,N_2359);
and U7580 (N_7580,N_2050,N_4970);
xnor U7581 (N_7581,N_2273,N_505);
and U7582 (N_7582,N_2386,N_4621);
xnor U7583 (N_7583,N_1140,N_3158);
nand U7584 (N_7584,N_2898,N_4640);
xnor U7585 (N_7585,N_588,N_657);
or U7586 (N_7586,N_4375,N_3330);
nand U7587 (N_7587,N_181,N_3288);
nor U7588 (N_7588,N_4574,N_3612);
or U7589 (N_7589,N_4540,N_3029);
nor U7590 (N_7590,N_51,N_897);
nand U7591 (N_7591,N_1736,N_2724);
or U7592 (N_7592,N_4332,N_4180);
or U7593 (N_7593,N_4538,N_4871);
nor U7594 (N_7594,N_1446,N_2857);
or U7595 (N_7595,N_3076,N_2197);
and U7596 (N_7596,N_1150,N_1691);
and U7597 (N_7597,N_3710,N_417);
or U7598 (N_7598,N_3584,N_4301);
nand U7599 (N_7599,N_4445,N_2206);
xor U7600 (N_7600,N_645,N_4530);
xnor U7601 (N_7601,N_448,N_2765);
nand U7602 (N_7602,N_4480,N_1425);
or U7603 (N_7603,N_3470,N_4788);
xor U7604 (N_7604,N_2779,N_246);
nor U7605 (N_7605,N_1399,N_1859);
or U7606 (N_7606,N_2624,N_4921);
nor U7607 (N_7607,N_3401,N_2624);
nand U7608 (N_7608,N_1999,N_648);
xnor U7609 (N_7609,N_2170,N_774);
xor U7610 (N_7610,N_1017,N_153);
nand U7611 (N_7611,N_3865,N_3113);
and U7612 (N_7612,N_4992,N_3675);
nand U7613 (N_7613,N_2686,N_4686);
xor U7614 (N_7614,N_4779,N_310);
xor U7615 (N_7615,N_2052,N_3708);
nand U7616 (N_7616,N_219,N_4877);
xor U7617 (N_7617,N_3314,N_2025);
and U7618 (N_7618,N_2013,N_4402);
xnor U7619 (N_7619,N_4574,N_3000);
nor U7620 (N_7620,N_4837,N_228);
nor U7621 (N_7621,N_436,N_4993);
nand U7622 (N_7622,N_2311,N_2959);
nand U7623 (N_7623,N_2281,N_2693);
xnor U7624 (N_7624,N_3143,N_1592);
or U7625 (N_7625,N_2711,N_1382);
nor U7626 (N_7626,N_811,N_1858);
nor U7627 (N_7627,N_137,N_556);
and U7628 (N_7628,N_3405,N_2615);
xor U7629 (N_7629,N_2930,N_2330);
or U7630 (N_7630,N_3859,N_777);
nand U7631 (N_7631,N_2012,N_644);
xnor U7632 (N_7632,N_777,N_354);
or U7633 (N_7633,N_3346,N_180);
nand U7634 (N_7634,N_1102,N_2468);
or U7635 (N_7635,N_1945,N_2443);
nand U7636 (N_7636,N_3219,N_2039);
nor U7637 (N_7637,N_3302,N_1286);
nor U7638 (N_7638,N_1155,N_4015);
nand U7639 (N_7639,N_1233,N_4060);
or U7640 (N_7640,N_362,N_3253);
and U7641 (N_7641,N_2340,N_2116);
nor U7642 (N_7642,N_2321,N_3930);
nand U7643 (N_7643,N_1848,N_3174);
or U7644 (N_7644,N_4209,N_3035);
xnor U7645 (N_7645,N_3129,N_4449);
and U7646 (N_7646,N_2593,N_3084);
and U7647 (N_7647,N_1412,N_243);
nand U7648 (N_7648,N_527,N_1179);
or U7649 (N_7649,N_3894,N_924);
nand U7650 (N_7650,N_288,N_3531);
or U7651 (N_7651,N_2857,N_824);
and U7652 (N_7652,N_1173,N_217);
and U7653 (N_7653,N_3273,N_2903);
or U7654 (N_7654,N_3245,N_1559);
nor U7655 (N_7655,N_8,N_4675);
or U7656 (N_7656,N_2675,N_2456);
or U7657 (N_7657,N_358,N_132);
nand U7658 (N_7658,N_1113,N_3120);
xor U7659 (N_7659,N_60,N_332);
nand U7660 (N_7660,N_1717,N_4505);
or U7661 (N_7661,N_3539,N_2595);
or U7662 (N_7662,N_2545,N_3187);
or U7663 (N_7663,N_1671,N_4795);
and U7664 (N_7664,N_3536,N_2249);
xnor U7665 (N_7665,N_1959,N_4784);
or U7666 (N_7666,N_166,N_4647);
xor U7667 (N_7667,N_2187,N_4327);
xnor U7668 (N_7668,N_2022,N_3028);
nand U7669 (N_7669,N_4934,N_2249);
and U7670 (N_7670,N_4080,N_3899);
nand U7671 (N_7671,N_3696,N_4503);
nor U7672 (N_7672,N_335,N_2594);
nand U7673 (N_7673,N_4636,N_628);
or U7674 (N_7674,N_4614,N_1796);
nor U7675 (N_7675,N_928,N_2446);
and U7676 (N_7676,N_814,N_4493);
nand U7677 (N_7677,N_1960,N_3453);
xor U7678 (N_7678,N_3705,N_1971);
xor U7679 (N_7679,N_19,N_2597);
xnor U7680 (N_7680,N_320,N_1671);
nor U7681 (N_7681,N_3897,N_4851);
xnor U7682 (N_7682,N_4258,N_2607);
xnor U7683 (N_7683,N_220,N_1560);
xnor U7684 (N_7684,N_746,N_781);
and U7685 (N_7685,N_2156,N_4575);
nand U7686 (N_7686,N_836,N_3746);
or U7687 (N_7687,N_479,N_620);
and U7688 (N_7688,N_4413,N_1226);
nor U7689 (N_7689,N_1882,N_775);
and U7690 (N_7690,N_310,N_3350);
and U7691 (N_7691,N_752,N_4754);
xor U7692 (N_7692,N_1353,N_4177);
and U7693 (N_7693,N_2148,N_4718);
and U7694 (N_7694,N_2881,N_3206);
nand U7695 (N_7695,N_2629,N_2113);
xnor U7696 (N_7696,N_1892,N_3556);
xor U7697 (N_7697,N_4316,N_2107);
nand U7698 (N_7698,N_3157,N_1512);
and U7699 (N_7699,N_4896,N_519);
nor U7700 (N_7700,N_2162,N_3765);
xor U7701 (N_7701,N_825,N_0);
or U7702 (N_7702,N_924,N_3226);
nor U7703 (N_7703,N_854,N_216);
nand U7704 (N_7704,N_643,N_1399);
or U7705 (N_7705,N_3712,N_2925);
xnor U7706 (N_7706,N_1125,N_3423);
and U7707 (N_7707,N_4644,N_2060);
xor U7708 (N_7708,N_3321,N_33);
and U7709 (N_7709,N_2511,N_286);
nand U7710 (N_7710,N_1244,N_169);
or U7711 (N_7711,N_1280,N_2029);
nand U7712 (N_7712,N_3371,N_3994);
xnor U7713 (N_7713,N_873,N_760);
or U7714 (N_7714,N_2681,N_131);
and U7715 (N_7715,N_3517,N_4422);
or U7716 (N_7716,N_4538,N_326);
nand U7717 (N_7717,N_1565,N_905);
and U7718 (N_7718,N_2858,N_141);
and U7719 (N_7719,N_2955,N_1033);
nand U7720 (N_7720,N_3608,N_2991);
nand U7721 (N_7721,N_4413,N_1795);
and U7722 (N_7722,N_2042,N_2429);
xnor U7723 (N_7723,N_2575,N_355);
nand U7724 (N_7724,N_3156,N_66);
or U7725 (N_7725,N_125,N_1543);
nand U7726 (N_7726,N_3362,N_405);
xor U7727 (N_7727,N_2285,N_1370);
and U7728 (N_7728,N_2210,N_3111);
and U7729 (N_7729,N_1375,N_868);
xnor U7730 (N_7730,N_183,N_3898);
and U7731 (N_7731,N_3500,N_905);
and U7732 (N_7732,N_3833,N_238);
xor U7733 (N_7733,N_855,N_4480);
or U7734 (N_7734,N_2588,N_557);
nor U7735 (N_7735,N_4407,N_1375);
or U7736 (N_7736,N_320,N_1172);
nand U7737 (N_7737,N_1502,N_1796);
nand U7738 (N_7738,N_2468,N_2026);
nor U7739 (N_7739,N_4383,N_4115);
or U7740 (N_7740,N_2428,N_2086);
and U7741 (N_7741,N_3703,N_4586);
nor U7742 (N_7742,N_2304,N_865);
or U7743 (N_7743,N_961,N_3681);
nand U7744 (N_7744,N_2243,N_1409);
or U7745 (N_7745,N_1512,N_573);
and U7746 (N_7746,N_2576,N_144);
or U7747 (N_7747,N_4779,N_1713);
xor U7748 (N_7748,N_502,N_1201);
nand U7749 (N_7749,N_1207,N_48);
or U7750 (N_7750,N_697,N_1813);
nor U7751 (N_7751,N_2401,N_752);
nor U7752 (N_7752,N_3933,N_153);
xor U7753 (N_7753,N_1513,N_620);
nor U7754 (N_7754,N_535,N_4796);
xnor U7755 (N_7755,N_3380,N_2780);
nand U7756 (N_7756,N_4307,N_1487);
xnor U7757 (N_7757,N_3430,N_4738);
nor U7758 (N_7758,N_1268,N_714);
or U7759 (N_7759,N_3078,N_4359);
and U7760 (N_7760,N_1625,N_2437);
nor U7761 (N_7761,N_3312,N_1838);
nand U7762 (N_7762,N_326,N_4987);
and U7763 (N_7763,N_4526,N_3837);
xor U7764 (N_7764,N_4038,N_1059);
nand U7765 (N_7765,N_890,N_963);
or U7766 (N_7766,N_2339,N_3502);
nand U7767 (N_7767,N_4851,N_4013);
nand U7768 (N_7768,N_188,N_1695);
or U7769 (N_7769,N_1168,N_2902);
or U7770 (N_7770,N_256,N_2925);
xor U7771 (N_7771,N_4215,N_3533);
and U7772 (N_7772,N_2084,N_4597);
nor U7773 (N_7773,N_1823,N_37);
nor U7774 (N_7774,N_2836,N_449);
xor U7775 (N_7775,N_4062,N_3112);
or U7776 (N_7776,N_1372,N_3879);
and U7777 (N_7777,N_2954,N_1498);
nor U7778 (N_7778,N_4905,N_2933);
or U7779 (N_7779,N_108,N_2863);
and U7780 (N_7780,N_3555,N_2312);
nor U7781 (N_7781,N_3831,N_3895);
and U7782 (N_7782,N_3577,N_4977);
xnor U7783 (N_7783,N_128,N_2507);
nand U7784 (N_7784,N_304,N_844);
nor U7785 (N_7785,N_716,N_2988);
nor U7786 (N_7786,N_3941,N_3950);
nor U7787 (N_7787,N_1158,N_2774);
nor U7788 (N_7788,N_1382,N_811);
and U7789 (N_7789,N_3146,N_3888);
nand U7790 (N_7790,N_3269,N_1346);
nor U7791 (N_7791,N_1914,N_712);
and U7792 (N_7792,N_3782,N_757);
and U7793 (N_7793,N_204,N_1860);
xor U7794 (N_7794,N_3632,N_2065);
nor U7795 (N_7795,N_138,N_1693);
nor U7796 (N_7796,N_2879,N_1304);
nor U7797 (N_7797,N_3794,N_310);
nand U7798 (N_7798,N_4252,N_3345);
and U7799 (N_7799,N_531,N_3691);
nor U7800 (N_7800,N_2682,N_1888);
xor U7801 (N_7801,N_109,N_3478);
nand U7802 (N_7802,N_447,N_2028);
or U7803 (N_7803,N_3712,N_687);
xor U7804 (N_7804,N_1806,N_3849);
or U7805 (N_7805,N_2667,N_1857);
nor U7806 (N_7806,N_4362,N_2196);
nor U7807 (N_7807,N_1953,N_776);
nor U7808 (N_7808,N_4522,N_4111);
xor U7809 (N_7809,N_4169,N_1281);
and U7810 (N_7810,N_1357,N_3890);
nor U7811 (N_7811,N_3365,N_35);
nand U7812 (N_7812,N_3295,N_2382);
nand U7813 (N_7813,N_2052,N_2977);
nand U7814 (N_7814,N_382,N_546);
nor U7815 (N_7815,N_3703,N_847);
nand U7816 (N_7816,N_4070,N_3339);
nor U7817 (N_7817,N_1688,N_4587);
nand U7818 (N_7818,N_2784,N_1531);
nor U7819 (N_7819,N_2397,N_4668);
nor U7820 (N_7820,N_2547,N_2587);
nor U7821 (N_7821,N_414,N_1785);
nor U7822 (N_7822,N_460,N_3338);
xor U7823 (N_7823,N_3298,N_4720);
nand U7824 (N_7824,N_4730,N_3673);
and U7825 (N_7825,N_1232,N_3122);
xor U7826 (N_7826,N_2877,N_3554);
nor U7827 (N_7827,N_2707,N_4682);
or U7828 (N_7828,N_3253,N_930);
or U7829 (N_7829,N_682,N_4678);
and U7830 (N_7830,N_3956,N_1148);
or U7831 (N_7831,N_4615,N_3497);
and U7832 (N_7832,N_4696,N_2118);
nor U7833 (N_7833,N_248,N_290);
nand U7834 (N_7834,N_4735,N_4806);
or U7835 (N_7835,N_4561,N_4062);
nand U7836 (N_7836,N_1330,N_1752);
xnor U7837 (N_7837,N_3277,N_2236);
xnor U7838 (N_7838,N_1214,N_205);
and U7839 (N_7839,N_3346,N_1621);
nand U7840 (N_7840,N_238,N_1136);
and U7841 (N_7841,N_2009,N_2617);
nor U7842 (N_7842,N_1513,N_3346);
or U7843 (N_7843,N_3430,N_1962);
nand U7844 (N_7844,N_1149,N_4603);
or U7845 (N_7845,N_379,N_3196);
nand U7846 (N_7846,N_1662,N_3631);
nand U7847 (N_7847,N_1050,N_3288);
and U7848 (N_7848,N_703,N_2715);
nor U7849 (N_7849,N_3320,N_626);
xnor U7850 (N_7850,N_4992,N_4051);
or U7851 (N_7851,N_1739,N_1432);
or U7852 (N_7852,N_4726,N_1612);
or U7853 (N_7853,N_782,N_440);
nor U7854 (N_7854,N_3082,N_183);
nand U7855 (N_7855,N_822,N_248);
or U7856 (N_7856,N_4920,N_1195);
or U7857 (N_7857,N_3713,N_1350);
nor U7858 (N_7858,N_3478,N_3849);
nand U7859 (N_7859,N_775,N_3402);
or U7860 (N_7860,N_1572,N_4842);
or U7861 (N_7861,N_2298,N_2675);
nor U7862 (N_7862,N_588,N_2794);
nand U7863 (N_7863,N_2719,N_164);
nand U7864 (N_7864,N_1765,N_2792);
and U7865 (N_7865,N_3301,N_1245);
xnor U7866 (N_7866,N_3466,N_2417);
or U7867 (N_7867,N_208,N_1608);
nor U7868 (N_7868,N_1278,N_497);
nor U7869 (N_7869,N_126,N_992);
and U7870 (N_7870,N_495,N_2311);
nor U7871 (N_7871,N_383,N_2550);
nor U7872 (N_7872,N_1983,N_1768);
nor U7873 (N_7873,N_4625,N_2841);
and U7874 (N_7874,N_4447,N_2792);
or U7875 (N_7875,N_4156,N_1882);
and U7876 (N_7876,N_4286,N_174);
nand U7877 (N_7877,N_624,N_1274);
nand U7878 (N_7878,N_3173,N_4527);
or U7879 (N_7879,N_712,N_1548);
or U7880 (N_7880,N_4176,N_2402);
and U7881 (N_7881,N_806,N_4274);
or U7882 (N_7882,N_2805,N_1246);
nor U7883 (N_7883,N_3072,N_85);
nor U7884 (N_7884,N_2598,N_2628);
or U7885 (N_7885,N_3835,N_4983);
or U7886 (N_7886,N_3277,N_1827);
nand U7887 (N_7887,N_3131,N_3563);
nor U7888 (N_7888,N_2472,N_1851);
nand U7889 (N_7889,N_1442,N_3819);
xnor U7890 (N_7890,N_1586,N_2131);
and U7891 (N_7891,N_176,N_1876);
nand U7892 (N_7892,N_979,N_1824);
xor U7893 (N_7893,N_4875,N_3982);
or U7894 (N_7894,N_3956,N_4183);
or U7895 (N_7895,N_4042,N_1557);
nor U7896 (N_7896,N_4691,N_3551);
or U7897 (N_7897,N_4990,N_3062);
nand U7898 (N_7898,N_1102,N_1073);
nor U7899 (N_7899,N_2099,N_3041);
xnor U7900 (N_7900,N_640,N_4175);
xor U7901 (N_7901,N_4379,N_2347);
nand U7902 (N_7902,N_194,N_1221);
nand U7903 (N_7903,N_4381,N_3024);
or U7904 (N_7904,N_3728,N_835);
and U7905 (N_7905,N_3268,N_2188);
xor U7906 (N_7906,N_2891,N_3834);
or U7907 (N_7907,N_2475,N_3520);
nor U7908 (N_7908,N_1573,N_1688);
or U7909 (N_7909,N_4446,N_196);
and U7910 (N_7910,N_2625,N_1021);
xor U7911 (N_7911,N_595,N_2427);
nor U7912 (N_7912,N_1619,N_2108);
nand U7913 (N_7913,N_4650,N_1022);
xnor U7914 (N_7914,N_2994,N_91);
and U7915 (N_7915,N_255,N_4783);
nand U7916 (N_7916,N_3300,N_4015);
and U7917 (N_7917,N_2741,N_1907);
and U7918 (N_7918,N_3290,N_2516);
or U7919 (N_7919,N_66,N_2896);
xor U7920 (N_7920,N_309,N_3868);
and U7921 (N_7921,N_2077,N_2032);
or U7922 (N_7922,N_3125,N_1452);
xnor U7923 (N_7923,N_2800,N_4635);
and U7924 (N_7924,N_919,N_1079);
xnor U7925 (N_7925,N_2700,N_2729);
or U7926 (N_7926,N_1537,N_235);
nand U7927 (N_7927,N_3444,N_4843);
xor U7928 (N_7928,N_3350,N_4163);
nand U7929 (N_7929,N_4802,N_1211);
xnor U7930 (N_7930,N_3354,N_3654);
nand U7931 (N_7931,N_3959,N_2818);
and U7932 (N_7932,N_3723,N_4117);
nand U7933 (N_7933,N_3696,N_4946);
and U7934 (N_7934,N_3782,N_1387);
nand U7935 (N_7935,N_2250,N_3172);
nand U7936 (N_7936,N_2463,N_2270);
or U7937 (N_7937,N_230,N_1439);
nor U7938 (N_7938,N_2394,N_4799);
nand U7939 (N_7939,N_3789,N_4702);
nand U7940 (N_7940,N_951,N_1147);
nor U7941 (N_7941,N_4065,N_1953);
or U7942 (N_7942,N_3370,N_3712);
and U7943 (N_7943,N_3661,N_1731);
nor U7944 (N_7944,N_680,N_3557);
and U7945 (N_7945,N_2695,N_304);
nor U7946 (N_7946,N_163,N_3193);
nor U7947 (N_7947,N_91,N_1421);
nor U7948 (N_7948,N_1328,N_3627);
xor U7949 (N_7949,N_1205,N_277);
nor U7950 (N_7950,N_3562,N_3132);
nand U7951 (N_7951,N_1663,N_4942);
nor U7952 (N_7952,N_4051,N_2117);
and U7953 (N_7953,N_2918,N_3909);
xor U7954 (N_7954,N_2617,N_2883);
nor U7955 (N_7955,N_2033,N_2832);
xor U7956 (N_7956,N_3009,N_1121);
nor U7957 (N_7957,N_3901,N_339);
nor U7958 (N_7958,N_2739,N_369);
nor U7959 (N_7959,N_1994,N_1002);
nand U7960 (N_7960,N_4861,N_1246);
or U7961 (N_7961,N_4755,N_3572);
nor U7962 (N_7962,N_940,N_3323);
nand U7963 (N_7963,N_4943,N_2246);
nor U7964 (N_7964,N_4997,N_1170);
xor U7965 (N_7965,N_3440,N_4517);
or U7966 (N_7966,N_4625,N_2182);
nand U7967 (N_7967,N_2905,N_149);
or U7968 (N_7968,N_285,N_2923);
and U7969 (N_7969,N_3552,N_3904);
nor U7970 (N_7970,N_2837,N_4926);
nor U7971 (N_7971,N_4823,N_1024);
and U7972 (N_7972,N_3569,N_644);
or U7973 (N_7973,N_1776,N_4643);
and U7974 (N_7974,N_4941,N_452);
and U7975 (N_7975,N_194,N_4276);
nor U7976 (N_7976,N_3736,N_4458);
nor U7977 (N_7977,N_266,N_4363);
nor U7978 (N_7978,N_227,N_1992);
and U7979 (N_7979,N_3378,N_2671);
xnor U7980 (N_7980,N_3524,N_65);
and U7981 (N_7981,N_2893,N_4009);
and U7982 (N_7982,N_3724,N_393);
xor U7983 (N_7983,N_2926,N_3499);
and U7984 (N_7984,N_259,N_2483);
nand U7985 (N_7985,N_4217,N_460);
nand U7986 (N_7986,N_3540,N_1415);
nand U7987 (N_7987,N_3821,N_3184);
xor U7988 (N_7988,N_4761,N_4377);
and U7989 (N_7989,N_1977,N_3943);
xor U7990 (N_7990,N_201,N_2002);
nand U7991 (N_7991,N_624,N_2390);
nand U7992 (N_7992,N_3201,N_4066);
nor U7993 (N_7993,N_4557,N_491);
nor U7994 (N_7994,N_4612,N_3091);
xor U7995 (N_7995,N_1830,N_1941);
and U7996 (N_7996,N_2535,N_2958);
nor U7997 (N_7997,N_4687,N_4341);
nor U7998 (N_7998,N_1697,N_3731);
nor U7999 (N_7999,N_3446,N_2317);
and U8000 (N_8000,N_1684,N_3053);
nand U8001 (N_8001,N_4572,N_3254);
nand U8002 (N_8002,N_1137,N_3873);
nor U8003 (N_8003,N_4351,N_2976);
xor U8004 (N_8004,N_3344,N_256);
nor U8005 (N_8005,N_4348,N_806);
and U8006 (N_8006,N_1255,N_3951);
xor U8007 (N_8007,N_2585,N_307);
nor U8008 (N_8008,N_2075,N_767);
xor U8009 (N_8009,N_4206,N_619);
and U8010 (N_8010,N_4641,N_3051);
xnor U8011 (N_8011,N_3267,N_4378);
nor U8012 (N_8012,N_3428,N_2405);
xor U8013 (N_8013,N_3506,N_3020);
xnor U8014 (N_8014,N_687,N_2222);
nor U8015 (N_8015,N_3029,N_1300);
nor U8016 (N_8016,N_3798,N_2077);
nor U8017 (N_8017,N_3063,N_3752);
or U8018 (N_8018,N_4793,N_1052);
nor U8019 (N_8019,N_990,N_1411);
nor U8020 (N_8020,N_2934,N_1896);
and U8021 (N_8021,N_3303,N_3971);
nand U8022 (N_8022,N_413,N_2692);
and U8023 (N_8023,N_937,N_1969);
xor U8024 (N_8024,N_4048,N_48);
nand U8025 (N_8025,N_3361,N_3380);
and U8026 (N_8026,N_4904,N_4567);
or U8027 (N_8027,N_3051,N_1141);
and U8028 (N_8028,N_1529,N_2829);
nand U8029 (N_8029,N_1275,N_4120);
xor U8030 (N_8030,N_3119,N_4391);
or U8031 (N_8031,N_4205,N_2124);
xnor U8032 (N_8032,N_3847,N_4937);
and U8033 (N_8033,N_1804,N_3458);
xor U8034 (N_8034,N_546,N_1546);
nand U8035 (N_8035,N_3126,N_4186);
nor U8036 (N_8036,N_436,N_3047);
or U8037 (N_8037,N_4073,N_3391);
nand U8038 (N_8038,N_1080,N_1801);
nor U8039 (N_8039,N_2838,N_4076);
and U8040 (N_8040,N_1681,N_1401);
and U8041 (N_8041,N_1723,N_1313);
or U8042 (N_8042,N_3574,N_2020);
nand U8043 (N_8043,N_2316,N_4393);
xor U8044 (N_8044,N_566,N_1541);
nor U8045 (N_8045,N_706,N_2461);
nand U8046 (N_8046,N_4140,N_3061);
nand U8047 (N_8047,N_2969,N_1713);
and U8048 (N_8048,N_4091,N_2850);
nor U8049 (N_8049,N_1890,N_4953);
xnor U8050 (N_8050,N_3027,N_4750);
nor U8051 (N_8051,N_444,N_1480);
xor U8052 (N_8052,N_3923,N_2808);
nor U8053 (N_8053,N_3965,N_1606);
and U8054 (N_8054,N_4905,N_291);
and U8055 (N_8055,N_99,N_4397);
or U8056 (N_8056,N_4291,N_1021);
nand U8057 (N_8057,N_2725,N_2076);
xnor U8058 (N_8058,N_2855,N_2376);
xnor U8059 (N_8059,N_2074,N_3398);
or U8060 (N_8060,N_783,N_705);
nand U8061 (N_8061,N_673,N_3788);
nand U8062 (N_8062,N_3993,N_1671);
and U8063 (N_8063,N_621,N_312);
or U8064 (N_8064,N_2891,N_1112);
or U8065 (N_8065,N_4988,N_4076);
nand U8066 (N_8066,N_1939,N_3177);
nand U8067 (N_8067,N_2953,N_1490);
xnor U8068 (N_8068,N_1023,N_1679);
and U8069 (N_8069,N_3798,N_1364);
nor U8070 (N_8070,N_774,N_2773);
xnor U8071 (N_8071,N_2397,N_4873);
xor U8072 (N_8072,N_4692,N_3962);
and U8073 (N_8073,N_3182,N_1538);
xor U8074 (N_8074,N_4244,N_1997);
nand U8075 (N_8075,N_3195,N_224);
or U8076 (N_8076,N_132,N_1388);
xnor U8077 (N_8077,N_3399,N_2413);
xor U8078 (N_8078,N_1163,N_3585);
or U8079 (N_8079,N_1263,N_1264);
nand U8080 (N_8080,N_248,N_2440);
nor U8081 (N_8081,N_40,N_4594);
xnor U8082 (N_8082,N_577,N_4126);
nor U8083 (N_8083,N_1223,N_217);
nor U8084 (N_8084,N_1717,N_2498);
nand U8085 (N_8085,N_1555,N_4778);
or U8086 (N_8086,N_3087,N_4136);
or U8087 (N_8087,N_3895,N_4959);
nor U8088 (N_8088,N_3327,N_2462);
xnor U8089 (N_8089,N_2224,N_3060);
xnor U8090 (N_8090,N_1634,N_4925);
xor U8091 (N_8091,N_261,N_4273);
and U8092 (N_8092,N_2783,N_3562);
and U8093 (N_8093,N_4246,N_4421);
and U8094 (N_8094,N_4193,N_4327);
nand U8095 (N_8095,N_608,N_2937);
nand U8096 (N_8096,N_4821,N_4665);
and U8097 (N_8097,N_1924,N_3020);
or U8098 (N_8098,N_2488,N_2215);
nand U8099 (N_8099,N_4666,N_3290);
nor U8100 (N_8100,N_2514,N_3408);
and U8101 (N_8101,N_3869,N_2289);
and U8102 (N_8102,N_3840,N_2386);
nor U8103 (N_8103,N_4572,N_4167);
nand U8104 (N_8104,N_3714,N_3769);
nor U8105 (N_8105,N_1124,N_1);
xnor U8106 (N_8106,N_4739,N_71);
xor U8107 (N_8107,N_4664,N_1945);
xnor U8108 (N_8108,N_3535,N_2677);
or U8109 (N_8109,N_3595,N_663);
or U8110 (N_8110,N_1380,N_2839);
nand U8111 (N_8111,N_4564,N_2);
xnor U8112 (N_8112,N_279,N_4637);
xor U8113 (N_8113,N_1767,N_1661);
or U8114 (N_8114,N_4031,N_753);
or U8115 (N_8115,N_4551,N_771);
or U8116 (N_8116,N_2659,N_2656);
and U8117 (N_8117,N_254,N_1198);
and U8118 (N_8118,N_4299,N_2017);
nand U8119 (N_8119,N_3842,N_402);
nand U8120 (N_8120,N_38,N_4177);
and U8121 (N_8121,N_2167,N_4342);
xor U8122 (N_8122,N_154,N_3014);
nand U8123 (N_8123,N_1188,N_4985);
nor U8124 (N_8124,N_2996,N_2193);
and U8125 (N_8125,N_633,N_2509);
or U8126 (N_8126,N_2844,N_2424);
or U8127 (N_8127,N_2657,N_3202);
nand U8128 (N_8128,N_2829,N_1717);
nand U8129 (N_8129,N_4114,N_3953);
xor U8130 (N_8130,N_3398,N_4767);
or U8131 (N_8131,N_3952,N_3181);
nand U8132 (N_8132,N_4431,N_591);
and U8133 (N_8133,N_2713,N_3956);
xnor U8134 (N_8134,N_3022,N_3782);
or U8135 (N_8135,N_4454,N_3139);
or U8136 (N_8136,N_4166,N_2313);
and U8137 (N_8137,N_3321,N_1844);
nor U8138 (N_8138,N_4852,N_2746);
xnor U8139 (N_8139,N_2900,N_2640);
nor U8140 (N_8140,N_3182,N_483);
nor U8141 (N_8141,N_74,N_691);
xnor U8142 (N_8142,N_1751,N_2815);
xor U8143 (N_8143,N_3991,N_2282);
or U8144 (N_8144,N_160,N_2435);
or U8145 (N_8145,N_859,N_2187);
or U8146 (N_8146,N_3946,N_3111);
nor U8147 (N_8147,N_2971,N_1476);
or U8148 (N_8148,N_1899,N_3685);
nor U8149 (N_8149,N_507,N_541);
nor U8150 (N_8150,N_1238,N_3736);
and U8151 (N_8151,N_2359,N_2409);
and U8152 (N_8152,N_2107,N_2868);
nor U8153 (N_8153,N_171,N_3549);
nor U8154 (N_8154,N_2537,N_4646);
nand U8155 (N_8155,N_14,N_2683);
or U8156 (N_8156,N_3882,N_3523);
nand U8157 (N_8157,N_4018,N_1035);
and U8158 (N_8158,N_589,N_1653);
nand U8159 (N_8159,N_3684,N_4905);
nand U8160 (N_8160,N_3524,N_4126);
nand U8161 (N_8161,N_4519,N_3718);
or U8162 (N_8162,N_4103,N_4660);
nand U8163 (N_8163,N_275,N_903);
xnor U8164 (N_8164,N_1142,N_859);
xnor U8165 (N_8165,N_1754,N_1922);
nand U8166 (N_8166,N_145,N_3739);
nand U8167 (N_8167,N_846,N_110);
and U8168 (N_8168,N_3368,N_2357);
nand U8169 (N_8169,N_4527,N_1637);
xnor U8170 (N_8170,N_4087,N_4534);
or U8171 (N_8171,N_49,N_1846);
and U8172 (N_8172,N_3495,N_2469);
nor U8173 (N_8173,N_3701,N_1019);
nand U8174 (N_8174,N_4459,N_4307);
or U8175 (N_8175,N_1005,N_3642);
nand U8176 (N_8176,N_1010,N_451);
and U8177 (N_8177,N_142,N_363);
nor U8178 (N_8178,N_3810,N_4973);
or U8179 (N_8179,N_522,N_1517);
nand U8180 (N_8180,N_1095,N_2259);
nor U8181 (N_8181,N_1827,N_4161);
nand U8182 (N_8182,N_1607,N_4716);
and U8183 (N_8183,N_137,N_3895);
nand U8184 (N_8184,N_2825,N_3897);
xnor U8185 (N_8185,N_4576,N_2560);
xnor U8186 (N_8186,N_1982,N_1263);
nand U8187 (N_8187,N_4104,N_2269);
and U8188 (N_8188,N_401,N_2901);
nand U8189 (N_8189,N_2336,N_43);
xnor U8190 (N_8190,N_2029,N_3605);
and U8191 (N_8191,N_3111,N_3413);
or U8192 (N_8192,N_3104,N_2829);
or U8193 (N_8193,N_857,N_1685);
nor U8194 (N_8194,N_2134,N_2748);
and U8195 (N_8195,N_4957,N_2174);
nor U8196 (N_8196,N_587,N_23);
xnor U8197 (N_8197,N_4520,N_1826);
and U8198 (N_8198,N_171,N_3946);
nor U8199 (N_8199,N_3352,N_3209);
nand U8200 (N_8200,N_1350,N_2867);
nor U8201 (N_8201,N_3766,N_3262);
nor U8202 (N_8202,N_1099,N_3228);
xnor U8203 (N_8203,N_1719,N_397);
nand U8204 (N_8204,N_1494,N_22);
and U8205 (N_8205,N_4943,N_278);
nor U8206 (N_8206,N_3536,N_506);
nand U8207 (N_8207,N_3368,N_2639);
and U8208 (N_8208,N_2775,N_1222);
and U8209 (N_8209,N_250,N_2830);
xor U8210 (N_8210,N_3170,N_3306);
and U8211 (N_8211,N_3873,N_2617);
xnor U8212 (N_8212,N_3893,N_3218);
and U8213 (N_8213,N_1762,N_2075);
and U8214 (N_8214,N_68,N_4575);
xor U8215 (N_8215,N_1863,N_2183);
nand U8216 (N_8216,N_3185,N_310);
or U8217 (N_8217,N_3544,N_695);
and U8218 (N_8218,N_900,N_133);
or U8219 (N_8219,N_3426,N_2066);
xnor U8220 (N_8220,N_1646,N_4672);
nor U8221 (N_8221,N_2114,N_884);
and U8222 (N_8222,N_2669,N_4310);
or U8223 (N_8223,N_2190,N_485);
nor U8224 (N_8224,N_2153,N_3759);
nand U8225 (N_8225,N_951,N_926);
nor U8226 (N_8226,N_4893,N_1027);
and U8227 (N_8227,N_3211,N_209);
nand U8228 (N_8228,N_4769,N_3636);
or U8229 (N_8229,N_2924,N_4615);
xnor U8230 (N_8230,N_2206,N_228);
or U8231 (N_8231,N_1880,N_4561);
nor U8232 (N_8232,N_3072,N_3826);
and U8233 (N_8233,N_285,N_3054);
nand U8234 (N_8234,N_3744,N_1084);
xor U8235 (N_8235,N_4968,N_3861);
nand U8236 (N_8236,N_2439,N_3162);
nor U8237 (N_8237,N_4148,N_4225);
or U8238 (N_8238,N_2101,N_4238);
nor U8239 (N_8239,N_4645,N_1725);
xor U8240 (N_8240,N_1288,N_2706);
or U8241 (N_8241,N_1275,N_4652);
and U8242 (N_8242,N_1071,N_607);
nor U8243 (N_8243,N_4539,N_484);
or U8244 (N_8244,N_4949,N_3229);
and U8245 (N_8245,N_1060,N_2508);
or U8246 (N_8246,N_2707,N_4303);
nor U8247 (N_8247,N_370,N_4929);
or U8248 (N_8248,N_2746,N_2917);
nor U8249 (N_8249,N_1381,N_3904);
xor U8250 (N_8250,N_3587,N_2061);
nor U8251 (N_8251,N_4362,N_1414);
nand U8252 (N_8252,N_4391,N_1548);
nor U8253 (N_8253,N_3004,N_823);
or U8254 (N_8254,N_120,N_1379);
or U8255 (N_8255,N_3339,N_1049);
or U8256 (N_8256,N_4467,N_2641);
xor U8257 (N_8257,N_1017,N_1297);
nand U8258 (N_8258,N_1115,N_1703);
xnor U8259 (N_8259,N_1904,N_299);
and U8260 (N_8260,N_1231,N_4483);
xor U8261 (N_8261,N_3956,N_705);
nor U8262 (N_8262,N_2666,N_1348);
nor U8263 (N_8263,N_1986,N_377);
nor U8264 (N_8264,N_2568,N_3911);
nand U8265 (N_8265,N_3964,N_1623);
or U8266 (N_8266,N_3876,N_1684);
and U8267 (N_8267,N_3963,N_1585);
and U8268 (N_8268,N_2055,N_1454);
nand U8269 (N_8269,N_1733,N_2109);
or U8270 (N_8270,N_391,N_2670);
xnor U8271 (N_8271,N_1708,N_3456);
xnor U8272 (N_8272,N_736,N_2656);
nor U8273 (N_8273,N_3092,N_3332);
and U8274 (N_8274,N_518,N_1423);
nand U8275 (N_8275,N_4568,N_2469);
or U8276 (N_8276,N_2552,N_1602);
xor U8277 (N_8277,N_3258,N_4165);
nand U8278 (N_8278,N_3705,N_2676);
nor U8279 (N_8279,N_210,N_4998);
nand U8280 (N_8280,N_1692,N_1600);
and U8281 (N_8281,N_4118,N_3386);
xnor U8282 (N_8282,N_3886,N_3399);
xnor U8283 (N_8283,N_1585,N_2250);
nand U8284 (N_8284,N_4077,N_617);
xnor U8285 (N_8285,N_2371,N_2937);
nand U8286 (N_8286,N_2678,N_4275);
or U8287 (N_8287,N_2322,N_4094);
nand U8288 (N_8288,N_83,N_4061);
nor U8289 (N_8289,N_4669,N_2039);
and U8290 (N_8290,N_2447,N_2476);
nand U8291 (N_8291,N_3315,N_2448);
nor U8292 (N_8292,N_3074,N_35);
nand U8293 (N_8293,N_2601,N_2439);
nor U8294 (N_8294,N_3345,N_2340);
and U8295 (N_8295,N_2105,N_3855);
nor U8296 (N_8296,N_1227,N_3574);
and U8297 (N_8297,N_2109,N_1434);
nor U8298 (N_8298,N_1696,N_1463);
or U8299 (N_8299,N_2004,N_1263);
and U8300 (N_8300,N_2426,N_2066);
and U8301 (N_8301,N_2659,N_955);
nor U8302 (N_8302,N_4846,N_2992);
or U8303 (N_8303,N_3213,N_2941);
or U8304 (N_8304,N_612,N_1403);
nor U8305 (N_8305,N_4766,N_2521);
xor U8306 (N_8306,N_3360,N_2791);
xnor U8307 (N_8307,N_599,N_1839);
nor U8308 (N_8308,N_4980,N_3464);
nor U8309 (N_8309,N_3406,N_2980);
nor U8310 (N_8310,N_2401,N_2996);
xnor U8311 (N_8311,N_2907,N_3120);
xnor U8312 (N_8312,N_3213,N_3149);
nor U8313 (N_8313,N_34,N_1078);
and U8314 (N_8314,N_3352,N_409);
and U8315 (N_8315,N_1648,N_4512);
xor U8316 (N_8316,N_66,N_1133);
nand U8317 (N_8317,N_4570,N_203);
and U8318 (N_8318,N_1503,N_2203);
nor U8319 (N_8319,N_878,N_3333);
xor U8320 (N_8320,N_3316,N_3082);
nor U8321 (N_8321,N_3142,N_869);
xnor U8322 (N_8322,N_3896,N_3771);
xnor U8323 (N_8323,N_3638,N_3014);
xnor U8324 (N_8324,N_4461,N_640);
nand U8325 (N_8325,N_691,N_3702);
nor U8326 (N_8326,N_2599,N_618);
xnor U8327 (N_8327,N_1048,N_4999);
nor U8328 (N_8328,N_647,N_3246);
and U8329 (N_8329,N_3258,N_4306);
xor U8330 (N_8330,N_1830,N_3058);
nor U8331 (N_8331,N_941,N_2202);
nor U8332 (N_8332,N_1439,N_1954);
nor U8333 (N_8333,N_3953,N_3409);
nand U8334 (N_8334,N_3297,N_1801);
xor U8335 (N_8335,N_1468,N_4697);
or U8336 (N_8336,N_836,N_2099);
and U8337 (N_8337,N_1906,N_3019);
or U8338 (N_8338,N_2679,N_2296);
and U8339 (N_8339,N_4010,N_750);
xor U8340 (N_8340,N_3684,N_3190);
or U8341 (N_8341,N_2067,N_698);
xnor U8342 (N_8342,N_218,N_4530);
or U8343 (N_8343,N_3955,N_961);
nand U8344 (N_8344,N_2724,N_3656);
or U8345 (N_8345,N_1171,N_1897);
and U8346 (N_8346,N_2920,N_2896);
xor U8347 (N_8347,N_2074,N_4212);
nand U8348 (N_8348,N_2236,N_2966);
nand U8349 (N_8349,N_495,N_2644);
nor U8350 (N_8350,N_2858,N_2507);
xor U8351 (N_8351,N_2517,N_4719);
and U8352 (N_8352,N_4824,N_2795);
and U8353 (N_8353,N_4665,N_4123);
xor U8354 (N_8354,N_2374,N_2863);
xnor U8355 (N_8355,N_3923,N_1044);
or U8356 (N_8356,N_3964,N_4640);
nand U8357 (N_8357,N_2435,N_75);
nand U8358 (N_8358,N_3087,N_2626);
nor U8359 (N_8359,N_405,N_3526);
or U8360 (N_8360,N_3397,N_329);
nor U8361 (N_8361,N_1937,N_2621);
nor U8362 (N_8362,N_1142,N_3258);
nor U8363 (N_8363,N_3063,N_1402);
or U8364 (N_8364,N_2108,N_1466);
or U8365 (N_8365,N_4885,N_4497);
and U8366 (N_8366,N_2846,N_4421);
or U8367 (N_8367,N_1956,N_1296);
and U8368 (N_8368,N_651,N_3252);
xor U8369 (N_8369,N_4954,N_1711);
xor U8370 (N_8370,N_3168,N_3846);
nand U8371 (N_8371,N_1162,N_852);
nor U8372 (N_8372,N_1907,N_4248);
xor U8373 (N_8373,N_1997,N_3905);
nor U8374 (N_8374,N_4063,N_115);
and U8375 (N_8375,N_4881,N_2359);
nand U8376 (N_8376,N_3512,N_2220);
and U8377 (N_8377,N_3977,N_1630);
nand U8378 (N_8378,N_4225,N_905);
or U8379 (N_8379,N_3190,N_2659);
xnor U8380 (N_8380,N_374,N_4827);
or U8381 (N_8381,N_2162,N_4617);
nand U8382 (N_8382,N_128,N_764);
nor U8383 (N_8383,N_1765,N_3866);
xnor U8384 (N_8384,N_25,N_3317);
or U8385 (N_8385,N_682,N_1499);
nor U8386 (N_8386,N_3748,N_781);
xnor U8387 (N_8387,N_953,N_983);
nand U8388 (N_8388,N_67,N_2561);
nand U8389 (N_8389,N_4612,N_4891);
nor U8390 (N_8390,N_4407,N_2112);
nand U8391 (N_8391,N_1225,N_4465);
xor U8392 (N_8392,N_2809,N_2683);
nor U8393 (N_8393,N_4002,N_3261);
or U8394 (N_8394,N_1007,N_1617);
or U8395 (N_8395,N_3159,N_2989);
nand U8396 (N_8396,N_2101,N_58);
and U8397 (N_8397,N_2569,N_4580);
or U8398 (N_8398,N_2588,N_1324);
or U8399 (N_8399,N_4831,N_81);
nand U8400 (N_8400,N_2118,N_4333);
and U8401 (N_8401,N_1433,N_4998);
nand U8402 (N_8402,N_1461,N_2994);
xor U8403 (N_8403,N_498,N_2284);
nand U8404 (N_8404,N_3681,N_995);
or U8405 (N_8405,N_3103,N_3817);
and U8406 (N_8406,N_1965,N_2232);
xnor U8407 (N_8407,N_4981,N_3876);
nor U8408 (N_8408,N_1743,N_1695);
or U8409 (N_8409,N_1265,N_985);
nor U8410 (N_8410,N_1780,N_3741);
or U8411 (N_8411,N_444,N_453);
xor U8412 (N_8412,N_795,N_4187);
nor U8413 (N_8413,N_3566,N_3016);
xnor U8414 (N_8414,N_4641,N_3177);
xnor U8415 (N_8415,N_2748,N_2654);
or U8416 (N_8416,N_3560,N_449);
or U8417 (N_8417,N_1446,N_3505);
and U8418 (N_8418,N_2149,N_2607);
or U8419 (N_8419,N_1457,N_1530);
nand U8420 (N_8420,N_3624,N_1845);
nand U8421 (N_8421,N_2517,N_2600);
and U8422 (N_8422,N_443,N_4525);
xor U8423 (N_8423,N_2736,N_3005);
xnor U8424 (N_8424,N_509,N_1528);
xor U8425 (N_8425,N_4791,N_3162);
or U8426 (N_8426,N_225,N_3849);
or U8427 (N_8427,N_1614,N_4878);
or U8428 (N_8428,N_1201,N_3506);
or U8429 (N_8429,N_3684,N_1875);
or U8430 (N_8430,N_4887,N_878);
xnor U8431 (N_8431,N_2877,N_553);
xnor U8432 (N_8432,N_4436,N_461);
xor U8433 (N_8433,N_3919,N_3124);
xnor U8434 (N_8434,N_1582,N_3372);
and U8435 (N_8435,N_3568,N_2220);
or U8436 (N_8436,N_622,N_4167);
nand U8437 (N_8437,N_4957,N_1766);
nor U8438 (N_8438,N_2289,N_2411);
xnor U8439 (N_8439,N_3027,N_2463);
and U8440 (N_8440,N_4193,N_3370);
and U8441 (N_8441,N_2941,N_291);
or U8442 (N_8442,N_1712,N_4464);
nor U8443 (N_8443,N_3687,N_2863);
nand U8444 (N_8444,N_132,N_1514);
and U8445 (N_8445,N_595,N_3264);
nand U8446 (N_8446,N_4079,N_4963);
xor U8447 (N_8447,N_1504,N_900);
xnor U8448 (N_8448,N_2476,N_685);
xnor U8449 (N_8449,N_3740,N_877);
nor U8450 (N_8450,N_2526,N_2976);
nand U8451 (N_8451,N_3303,N_1617);
or U8452 (N_8452,N_3736,N_703);
xnor U8453 (N_8453,N_3715,N_3265);
or U8454 (N_8454,N_941,N_2174);
xor U8455 (N_8455,N_689,N_4805);
xor U8456 (N_8456,N_81,N_4165);
and U8457 (N_8457,N_1471,N_3450);
xor U8458 (N_8458,N_4084,N_2443);
xnor U8459 (N_8459,N_4574,N_2688);
and U8460 (N_8460,N_66,N_3973);
nor U8461 (N_8461,N_706,N_2853);
xnor U8462 (N_8462,N_3248,N_4885);
nand U8463 (N_8463,N_3520,N_717);
and U8464 (N_8464,N_1973,N_3174);
nand U8465 (N_8465,N_463,N_3735);
or U8466 (N_8466,N_3711,N_2369);
xor U8467 (N_8467,N_4273,N_4715);
nor U8468 (N_8468,N_1478,N_3609);
and U8469 (N_8469,N_1561,N_3971);
or U8470 (N_8470,N_1175,N_3369);
nand U8471 (N_8471,N_635,N_3309);
or U8472 (N_8472,N_2727,N_4328);
or U8473 (N_8473,N_2165,N_2236);
and U8474 (N_8474,N_671,N_708);
xor U8475 (N_8475,N_2283,N_4297);
nand U8476 (N_8476,N_2002,N_2374);
nand U8477 (N_8477,N_603,N_3265);
xor U8478 (N_8478,N_3903,N_3383);
and U8479 (N_8479,N_3979,N_810);
nor U8480 (N_8480,N_41,N_87);
or U8481 (N_8481,N_2783,N_4207);
xnor U8482 (N_8482,N_2737,N_3559);
xor U8483 (N_8483,N_535,N_3908);
nand U8484 (N_8484,N_4394,N_342);
xnor U8485 (N_8485,N_834,N_3549);
nor U8486 (N_8486,N_3028,N_2265);
xor U8487 (N_8487,N_3198,N_4506);
nor U8488 (N_8488,N_157,N_1349);
xnor U8489 (N_8489,N_1366,N_2737);
xnor U8490 (N_8490,N_2410,N_1606);
or U8491 (N_8491,N_3192,N_1361);
and U8492 (N_8492,N_532,N_266);
nand U8493 (N_8493,N_356,N_2647);
nor U8494 (N_8494,N_2024,N_4150);
nor U8495 (N_8495,N_520,N_2465);
or U8496 (N_8496,N_1604,N_1454);
and U8497 (N_8497,N_4350,N_1104);
nand U8498 (N_8498,N_2161,N_4651);
and U8499 (N_8499,N_88,N_792);
nor U8500 (N_8500,N_4111,N_174);
nand U8501 (N_8501,N_3921,N_4027);
xor U8502 (N_8502,N_2690,N_1816);
or U8503 (N_8503,N_1770,N_192);
and U8504 (N_8504,N_2690,N_2972);
nand U8505 (N_8505,N_2942,N_1564);
nor U8506 (N_8506,N_3464,N_3556);
or U8507 (N_8507,N_522,N_4561);
nand U8508 (N_8508,N_867,N_3522);
nand U8509 (N_8509,N_2972,N_3787);
or U8510 (N_8510,N_1919,N_4004);
or U8511 (N_8511,N_3836,N_284);
and U8512 (N_8512,N_106,N_3275);
xnor U8513 (N_8513,N_631,N_4011);
and U8514 (N_8514,N_4785,N_2171);
or U8515 (N_8515,N_3208,N_4633);
nand U8516 (N_8516,N_3697,N_2672);
nand U8517 (N_8517,N_3847,N_2353);
xnor U8518 (N_8518,N_2504,N_699);
and U8519 (N_8519,N_4666,N_3037);
or U8520 (N_8520,N_1264,N_2461);
nor U8521 (N_8521,N_1491,N_3081);
or U8522 (N_8522,N_2579,N_1080);
nand U8523 (N_8523,N_3643,N_1234);
or U8524 (N_8524,N_1763,N_1299);
xor U8525 (N_8525,N_1323,N_1166);
nor U8526 (N_8526,N_1406,N_3408);
nor U8527 (N_8527,N_4900,N_3842);
nand U8528 (N_8528,N_4955,N_3195);
or U8529 (N_8529,N_55,N_35);
nor U8530 (N_8530,N_4086,N_1854);
nor U8531 (N_8531,N_1402,N_1273);
xor U8532 (N_8532,N_2507,N_394);
xor U8533 (N_8533,N_1075,N_2749);
or U8534 (N_8534,N_3627,N_980);
nor U8535 (N_8535,N_2222,N_1098);
xor U8536 (N_8536,N_3866,N_3318);
xor U8537 (N_8537,N_3761,N_2927);
xnor U8538 (N_8538,N_3974,N_3114);
and U8539 (N_8539,N_3863,N_1358);
xnor U8540 (N_8540,N_98,N_1888);
nor U8541 (N_8541,N_1074,N_3577);
and U8542 (N_8542,N_4815,N_723);
and U8543 (N_8543,N_213,N_3555);
xnor U8544 (N_8544,N_2955,N_3498);
or U8545 (N_8545,N_1685,N_4603);
xor U8546 (N_8546,N_4554,N_1992);
and U8547 (N_8547,N_3329,N_4665);
and U8548 (N_8548,N_4256,N_3173);
nor U8549 (N_8549,N_654,N_4961);
nand U8550 (N_8550,N_2527,N_2405);
or U8551 (N_8551,N_1694,N_3064);
and U8552 (N_8552,N_4992,N_20);
nand U8553 (N_8553,N_2005,N_3957);
xor U8554 (N_8554,N_3359,N_1558);
and U8555 (N_8555,N_3388,N_4178);
or U8556 (N_8556,N_393,N_4850);
xnor U8557 (N_8557,N_2461,N_3299);
nor U8558 (N_8558,N_3259,N_1854);
nor U8559 (N_8559,N_3573,N_3763);
and U8560 (N_8560,N_3141,N_4646);
nand U8561 (N_8561,N_4793,N_1222);
nand U8562 (N_8562,N_4535,N_806);
and U8563 (N_8563,N_618,N_1353);
and U8564 (N_8564,N_4224,N_487);
and U8565 (N_8565,N_2554,N_4018);
nand U8566 (N_8566,N_4446,N_4144);
nor U8567 (N_8567,N_2234,N_3024);
or U8568 (N_8568,N_325,N_1115);
xnor U8569 (N_8569,N_3334,N_3204);
xor U8570 (N_8570,N_4642,N_4511);
nor U8571 (N_8571,N_3865,N_3275);
nand U8572 (N_8572,N_371,N_1459);
or U8573 (N_8573,N_1977,N_2499);
nor U8574 (N_8574,N_1484,N_2247);
nand U8575 (N_8575,N_4429,N_1869);
xnor U8576 (N_8576,N_3214,N_200);
xor U8577 (N_8577,N_503,N_1458);
or U8578 (N_8578,N_2690,N_770);
nand U8579 (N_8579,N_4622,N_1900);
nand U8580 (N_8580,N_1374,N_2322);
or U8581 (N_8581,N_3948,N_1561);
xnor U8582 (N_8582,N_2963,N_3469);
and U8583 (N_8583,N_2848,N_2758);
xor U8584 (N_8584,N_4548,N_3014);
nand U8585 (N_8585,N_1232,N_239);
and U8586 (N_8586,N_2034,N_2640);
nand U8587 (N_8587,N_615,N_405);
xor U8588 (N_8588,N_315,N_4283);
or U8589 (N_8589,N_2422,N_1207);
nor U8590 (N_8590,N_1987,N_4044);
nand U8591 (N_8591,N_1468,N_1293);
nor U8592 (N_8592,N_2632,N_3288);
nand U8593 (N_8593,N_4595,N_4643);
and U8594 (N_8594,N_1808,N_3784);
nand U8595 (N_8595,N_172,N_2790);
and U8596 (N_8596,N_4211,N_4240);
nand U8597 (N_8597,N_509,N_2480);
and U8598 (N_8598,N_475,N_4723);
and U8599 (N_8599,N_4098,N_3508);
xnor U8600 (N_8600,N_1695,N_2231);
nor U8601 (N_8601,N_2820,N_1305);
nor U8602 (N_8602,N_4461,N_59);
xnor U8603 (N_8603,N_2825,N_4587);
nor U8604 (N_8604,N_217,N_3289);
xor U8605 (N_8605,N_1006,N_2415);
or U8606 (N_8606,N_2448,N_1364);
nor U8607 (N_8607,N_2785,N_969);
nand U8608 (N_8608,N_2793,N_4938);
or U8609 (N_8609,N_3954,N_1154);
or U8610 (N_8610,N_1826,N_1761);
nand U8611 (N_8611,N_769,N_2758);
nand U8612 (N_8612,N_3305,N_3392);
or U8613 (N_8613,N_4498,N_3594);
nand U8614 (N_8614,N_589,N_3998);
nand U8615 (N_8615,N_2869,N_4643);
xnor U8616 (N_8616,N_2216,N_710);
or U8617 (N_8617,N_787,N_2049);
nor U8618 (N_8618,N_2596,N_2209);
and U8619 (N_8619,N_4348,N_32);
nand U8620 (N_8620,N_4672,N_1912);
nand U8621 (N_8621,N_850,N_3917);
or U8622 (N_8622,N_3103,N_2456);
xor U8623 (N_8623,N_3060,N_4464);
or U8624 (N_8624,N_2654,N_975);
nor U8625 (N_8625,N_21,N_4029);
nand U8626 (N_8626,N_4474,N_1080);
nand U8627 (N_8627,N_3425,N_2445);
or U8628 (N_8628,N_4789,N_2671);
or U8629 (N_8629,N_4104,N_2954);
nand U8630 (N_8630,N_678,N_795);
nand U8631 (N_8631,N_4449,N_255);
nor U8632 (N_8632,N_4886,N_3283);
nor U8633 (N_8633,N_609,N_4983);
or U8634 (N_8634,N_3862,N_2681);
and U8635 (N_8635,N_1974,N_1197);
and U8636 (N_8636,N_1179,N_2054);
xor U8637 (N_8637,N_359,N_4058);
nor U8638 (N_8638,N_4555,N_2730);
and U8639 (N_8639,N_4789,N_2342);
xnor U8640 (N_8640,N_1355,N_3187);
and U8641 (N_8641,N_3335,N_136);
and U8642 (N_8642,N_1318,N_2169);
and U8643 (N_8643,N_2668,N_178);
nor U8644 (N_8644,N_45,N_1488);
nand U8645 (N_8645,N_108,N_4259);
and U8646 (N_8646,N_1994,N_4117);
and U8647 (N_8647,N_1306,N_910);
and U8648 (N_8648,N_4572,N_3527);
nor U8649 (N_8649,N_4063,N_2816);
or U8650 (N_8650,N_1011,N_503);
nand U8651 (N_8651,N_4167,N_913);
or U8652 (N_8652,N_1278,N_377);
nand U8653 (N_8653,N_2817,N_2954);
and U8654 (N_8654,N_3335,N_4392);
nor U8655 (N_8655,N_3499,N_3877);
xor U8656 (N_8656,N_323,N_292);
nor U8657 (N_8657,N_21,N_3162);
nor U8658 (N_8658,N_2850,N_2713);
and U8659 (N_8659,N_815,N_1198);
and U8660 (N_8660,N_165,N_1631);
and U8661 (N_8661,N_4328,N_1907);
xnor U8662 (N_8662,N_2536,N_762);
or U8663 (N_8663,N_2217,N_4433);
nor U8664 (N_8664,N_1359,N_1022);
nor U8665 (N_8665,N_586,N_2504);
nand U8666 (N_8666,N_1778,N_1559);
and U8667 (N_8667,N_2005,N_1376);
nor U8668 (N_8668,N_966,N_861);
xnor U8669 (N_8669,N_899,N_270);
nand U8670 (N_8670,N_4722,N_2958);
or U8671 (N_8671,N_522,N_4598);
xor U8672 (N_8672,N_2298,N_408);
nor U8673 (N_8673,N_1369,N_2530);
xnor U8674 (N_8674,N_402,N_2721);
xor U8675 (N_8675,N_3334,N_4239);
nand U8676 (N_8676,N_4422,N_86);
and U8677 (N_8677,N_1168,N_4590);
nor U8678 (N_8678,N_1145,N_4094);
nor U8679 (N_8679,N_65,N_1502);
nand U8680 (N_8680,N_3884,N_4573);
nand U8681 (N_8681,N_263,N_2691);
or U8682 (N_8682,N_1753,N_2260);
xnor U8683 (N_8683,N_3951,N_483);
nor U8684 (N_8684,N_41,N_692);
or U8685 (N_8685,N_4696,N_2562);
nor U8686 (N_8686,N_1434,N_3883);
xnor U8687 (N_8687,N_4787,N_4496);
nand U8688 (N_8688,N_4089,N_4273);
nand U8689 (N_8689,N_2711,N_3425);
and U8690 (N_8690,N_4700,N_3897);
or U8691 (N_8691,N_2455,N_1931);
nand U8692 (N_8692,N_2760,N_1791);
xnor U8693 (N_8693,N_3214,N_1890);
nor U8694 (N_8694,N_559,N_2788);
xor U8695 (N_8695,N_175,N_1858);
nand U8696 (N_8696,N_1583,N_4128);
nand U8697 (N_8697,N_117,N_463);
xnor U8698 (N_8698,N_428,N_1440);
nor U8699 (N_8699,N_1432,N_2631);
and U8700 (N_8700,N_1251,N_386);
and U8701 (N_8701,N_3245,N_3071);
or U8702 (N_8702,N_1250,N_1808);
xor U8703 (N_8703,N_120,N_4864);
xor U8704 (N_8704,N_2011,N_2135);
xnor U8705 (N_8705,N_4802,N_3500);
and U8706 (N_8706,N_1415,N_472);
or U8707 (N_8707,N_4174,N_808);
nor U8708 (N_8708,N_2244,N_1292);
nor U8709 (N_8709,N_2706,N_4525);
nand U8710 (N_8710,N_4613,N_4205);
xnor U8711 (N_8711,N_595,N_760);
and U8712 (N_8712,N_445,N_3381);
and U8713 (N_8713,N_2578,N_4801);
nand U8714 (N_8714,N_2141,N_1231);
and U8715 (N_8715,N_1311,N_2614);
nand U8716 (N_8716,N_726,N_604);
xnor U8717 (N_8717,N_572,N_4227);
nand U8718 (N_8718,N_4839,N_2468);
or U8719 (N_8719,N_4896,N_165);
and U8720 (N_8720,N_3841,N_2155);
or U8721 (N_8721,N_3189,N_25);
or U8722 (N_8722,N_247,N_671);
xor U8723 (N_8723,N_3174,N_2911);
and U8724 (N_8724,N_258,N_2958);
and U8725 (N_8725,N_3032,N_1359);
nor U8726 (N_8726,N_157,N_1330);
nand U8727 (N_8727,N_1040,N_625);
and U8728 (N_8728,N_2515,N_2443);
or U8729 (N_8729,N_4606,N_1932);
nor U8730 (N_8730,N_3553,N_2130);
nor U8731 (N_8731,N_919,N_1432);
xnor U8732 (N_8732,N_396,N_983);
nor U8733 (N_8733,N_3663,N_4938);
nor U8734 (N_8734,N_4455,N_3601);
nor U8735 (N_8735,N_1257,N_3161);
or U8736 (N_8736,N_1942,N_1555);
xor U8737 (N_8737,N_1052,N_2832);
or U8738 (N_8738,N_1055,N_4004);
or U8739 (N_8739,N_4566,N_260);
xnor U8740 (N_8740,N_2755,N_4396);
nand U8741 (N_8741,N_180,N_4729);
nor U8742 (N_8742,N_1190,N_3264);
nor U8743 (N_8743,N_3637,N_2532);
nand U8744 (N_8744,N_2387,N_2521);
or U8745 (N_8745,N_979,N_2541);
or U8746 (N_8746,N_3965,N_4718);
or U8747 (N_8747,N_1014,N_4299);
or U8748 (N_8748,N_1421,N_3744);
and U8749 (N_8749,N_2446,N_1411);
nor U8750 (N_8750,N_2611,N_1410);
nand U8751 (N_8751,N_2784,N_4136);
xor U8752 (N_8752,N_1379,N_4510);
nand U8753 (N_8753,N_4487,N_2149);
xnor U8754 (N_8754,N_3249,N_3218);
nor U8755 (N_8755,N_1459,N_2492);
and U8756 (N_8756,N_3093,N_4665);
and U8757 (N_8757,N_4992,N_1347);
or U8758 (N_8758,N_220,N_1028);
nor U8759 (N_8759,N_20,N_4141);
xor U8760 (N_8760,N_34,N_1966);
or U8761 (N_8761,N_2241,N_4576);
nor U8762 (N_8762,N_1947,N_3548);
or U8763 (N_8763,N_1984,N_3074);
and U8764 (N_8764,N_3467,N_4482);
nor U8765 (N_8765,N_1707,N_4880);
nor U8766 (N_8766,N_3536,N_3191);
xor U8767 (N_8767,N_687,N_503);
and U8768 (N_8768,N_1403,N_451);
nor U8769 (N_8769,N_3896,N_453);
nor U8770 (N_8770,N_778,N_3102);
xnor U8771 (N_8771,N_1117,N_1242);
or U8772 (N_8772,N_3660,N_4217);
or U8773 (N_8773,N_2394,N_758);
xnor U8774 (N_8774,N_2328,N_4918);
nor U8775 (N_8775,N_4489,N_1178);
nor U8776 (N_8776,N_4954,N_770);
nor U8777 (N_8777,N_1408,N_4005);
nor U8778 (N_8778,N_4075,N_681);
or U8779 (N_8779,N_4202,N_4688);
xor U8780 (N_8780,N_2968,N_33);
nor U8781 (N_8781,N_628,N_1637);
xnor U8782 (N_8782,N_1342,N_2736);
nor U8783 (N_8783,N_55,N_2663);
or U8784 (N_8784,N_2635,N_2922);
or U8785 (N_8785,N_4539,N_3521);
nand U8786 (N_8786,N_2853,N_289);
and U8787 (N_8787,N_3782,N_3697);
xnor U8788 (N_8788,N_349,N_4582);
xnor U8789 (N_8789,N_1527,N_4723);
xor U8790 (N_8790,N_3963,N_1850);
or U8791 (N_8791,N_2937,N_2934);
nand U8792 (N_8792,N_4045,N_218);
nor U8793 (N_8793,N_3421,N_3346);
xnor U8794 (N_8794,N_767,N_1709);
xor U8795 (N_8795,N_2501,N_2623);
xor U8796 (N_8796,N_2752,N_2641);
xor U8797 (N_8797,N_4380,N_125);
xor U8798 (N_8798,N_418,N_162);
nand U8799 (N_8799,N_3853,N_1161);
and U8800 (N_8800,N_489,N_3916);
and U8801 (N_8801,N_3391,N_3751);
and U8802 (N_8802,N_4565,N_4781);
or U8803 (N_8803,N_1170,N_3269);
and U8804 (N_8804,N_1727,N_2371);
nand U8805 (N_8805,N_4943,N_3972);
and U8806 (N_8806,N_2091,N_344);
and U8807 (N_8807,N_954,N_4447);
and U8808 (N_8808,N_2635,N_4303);
or U8809 (N_8809,N_4136,N_2919);
nor U8810 (N_8810,N_3883,N_4898);
or U8811 (N_8811,N_4265,N_796);
nor U8812 (N_8812,N_1113,N_695);
xnor U8813 (N_8813,N_4826,N_4378);
nand U8814 (N_8814,N_4075,N_3422);
nand U8815 (N_8815,N_2081,N_3776);
and U8816 (N_8816,N_4664,N_2743);
nand U8817 (N_8817,N_3075,N_4940);
nor U8818 (N_8818,N_404,N_4054);
xor U8819 (N_8819,N_3617,N_2296);
xor U8820 (N_8820,N_2474,N_3059);
nor U8821 (N_8821,N_1027,N_2519);
nand U8822 (N_8822,N_3055,N_532);
xnor U8823 (N_8823,N_2453,N_2285);
nand U8824 (N_8824,N_3547,N_1550);
and U8825 (N_8825,N_668,N_2952);
xor U8826 (N_8826,N_4688,N_4531);
nand U8827 (N_8827,N_4734,N_4118);
nor U8828 (N_8828,N_1316,N_2745);
nand U8829 (N_8829,N_3897,N_2072);
and U8830 (N_8830,N_2636,N_4720);
or U8831 (N_8831,N_543,N_1611);
and U8832 (N_8832,N_4906,N_2583);
xnor U8833 (N_8833,N_1883,N_2576);
nand U8834 (N_8834,N_1484,N_2541);
and U8835 (N_8835,N_634,N_55);
or U8836 (N_8836,N_3070,N_2079);
or U8837 (N_8837,N_4533,N_4419);
xor U8838 (N_8838,N_3595,N_851);
nor U8839 (N_8839,N_852,N_3373);
nor U8840 (N_8840,N_526,N_3705);
and U8841 (N_8841,N_1786,N_2234);
nor U8842 (N_8842,N_2990,N_1188);
nor U8843 (N_8843,N_3000,N_1795);
nand U8844 (N_8844,N_3969,N_4548);
and U8845 (N_8845,N_1717,N_1802);
nor U8846 (N_8846,N_2160,N_3995);
or U8847 (N_8847,N_3896,N_3527);
nor U8848 (N_8848,N_4997,N_4795);
nand U8849 (N_8849,N_1119,N_2393);
xnor U8850 (N_8850,N_3488,N_2946);
nand U8851 (N_8851,N_2012,N_771);
nor U8852 (N_8852,N_2849,N_2459);
or U8853 (N_8853,N_801,N_4964);
nor U8854 (N_8854,N_2497,N_2630);
xnor U8855 (N_8855,N_360,N_792);
nor U8856 (N_8856,N_2686,N_359);
nand U8857 (N_8857,N_97,N_2631);
nand U8858 (N_8858,N_3536,N_3200);
xor U8859 (N_8859,N_3350,N_1108);
nand U8860 (N_8860,N_3868,N_833);
or U8861 (N_8861,N_1512,N_1008);
xnor U8862 (N_8862,N_2580,N_600);
nand U8863 (N_8863,N_29,N_2665);
nor U8864 (N_8864,N_1072,N_857);
and U8865 (N_8865,N_3100,N_1436);
or U8866 (N_8866,N_683,N_3735);
nor U8867 (N_8867,N_2702,N_3076);
or U8868 (N_8868,N_4656,N_1620);
nand U8869 (N_8869,N_4716,N_3945);
and U8870 (N_8870,N_2450,N_3488);
xnor U8871 (N_8871,N_1056,N_2012);
or U8872 (N_8872,N_4639,N_2256);
and U8873 (N_8873,N_2986,N_1691);
nor U8874 (N_8874,N_595,N_541);
and U8875 (N_8875,N_4402,N_3362);
xnor U8876 (N_8876,N_685,N_1494);
or U8877 (N_8877,N_4666,N_2541);
nand U8878 (N_8878,N_4292,N_1111);
xor U8879 (N_8879,N_492,N_390);
or U8880 (N_8880,N_2698,N_4592);
or U8881 (N_8881,N_3104,N_279);
nor U8882 (N_8882,N_2950,N_4127);
xnor U8883 (N_8883,N_1582,N_1889);
nand U8884 (N_8884,N_456,N_2143);
xnor U8885 (N_8885,N_4333,N_4201);
or U8886 (N_8886,N_1096,N_1632);
or U8887 (N_8887,N_1991,N_3543);
and U8888 (N_8888,N_4748,N_694);
nor U8889 (N_8889,N_1286,N_1721);
nor U8890 (N_8890,N_4124,N_2967);
xor U8891 (N_8891,N_4477,N_3915);
nor U8892 (N_8892,N_3457,N_1501);
xor U8893 (N_8893,N_792,N_1744);
nand U8894 (N_8894,N_1977,N_3328);
nor U8895 (N_8895,N_2862,N_4082);
xor U8896 (N_8896,N_2169,N_3622);
nor U8897 (N_8897,N_3891,N_165);
and U8898 (N_8898,N_2859,N_178);
nor U8899 (N_8899,N_3574,N_721);
nor U8900 (N_8900,N_4810,N_4250);
or U8901 (N_8901,N_3143,N_2891);
nand U8902 (N_8902,N_3577,N_3295);
or U8903 (N_8903,N_1794,N_510);
xor U8904 (N_8904,N_2501,N_3740);
or U8905 (N_8905,N_385,N_3647);
nand U8906 (N_8906,N_1608,N_1776);
xnor U8907 (N_8907,N_2588,N_3078);
nor U8908 (N_8908,N_204,N_63);
nor U8909 (N_8909,N_3288,N_1908);
or U8910 (N_8910,N_2537,N_307);
nand U8911 (N_8911,N_2603,N_1084);
nand U8912 (N_8912,N_680,N_1379);
xnor U8913 (N_8913,N_2062,N_4623);
nand U8914 (N_8914,N_2608,N_1273);
or U8915 (N_8915,N_4344,N_4445);
nand U8916 (N_8916,N_1931,N_4347);
or U8917 (N_8917,N_3428,N_1398);
and U8918 (N_8918,N_4627,N_3243);
xor U8919 (N_8919,N_4864,N_4540);
or U8920 (N_8920,N_2088,N_3037);
nand U8921 (N_8921,N_1289,N_2960);
or U8922 (N_8922,N_2539,N_2083);
nor U8923 (N_8923,N_2615,N_439);
nand U8924 (N_8924,N_4717,N_3399);
nand U8925 (N_8925,N_1646,N_3517);
and U8926 (N_8926,N_3156,N_923);
or U8927 (N_8927,N_4190,N_4789);
and U8928 (N_8928,N_3374,N_2064);
or U8929 (N_8929,N_2764,N_4790);
and U8930 (N_8930,N_341,N_311);
and U8931 (N_8931,N_4419,N_4330);
nand U8932 (N_8932,N_1841,N_3878);
nor U8933 (N_8933,N_3263,N_3934);
and U8934 (N_8934,N_2214,N_234);
nand U8935 (N_8935,N_4001,N_3634);
xnor U8936 (N_8936,N_668,N_3779);
nand U8937 (N_8937,N_1495,N_469);
and U8938 (N_8938,N_559,N_2537);
xor U8939 (N_8939,N_170,N_421);
nand U8940 (N_8940,N_203,N_4094);
nand U8941 (N_8941,N_3181,N_1659);
nand U8942 (N_8942,N_1022,N_106);
and U8943 (N_8943,N_3682,N_344);
or U8944 (N_8944,N_3421,N_2527);
or U8945 (N_8945,N_847,N_3240);
xor U8946 (N_8946,N_3571,N_559);
or U8947 (N_8947,N_2218,N_3252);
and U8948 (N_8948,N_4124,N_2617);
xnor U8949 (N_8949,N_3728,N_4210);
and U8950 (N_8950,N_2232,N_3638);
nor U8951 (N_8951,N_4011,N_4061);
nor U8952 (N_8952,N_1169,N_1973);
xor U8953 (N_8953,N_273,N_650);
nor U8954 (N_8954,N_3297,N_4067);
nor U8955 (N_8955,N_3833,N_4684);
nor U8956 (N_8956,N_181,N_2077);
nor U8957 (N_8957,N_2646,N_4166);
nor U8958 (N_8958,N_3355,N_3021);
or U8959 (N_8959,N_470,N_3769);
or U8960 (N_8960,N_3997,N_1621);
nor U8961 (N_8961,N_2306,N_2714);
nor U8962 (N_8962,N_3598,N_3747);
nor U8963 (N_8963,N_3698,N_1802);
nor U8964 (N_8964,N_2037,N_467);
or U8965 (N_8965,N_4111,N_2075);
or U8966 (N_8966,N_3265,N_4190);
nand U8967 (N_8967,N_3660,N_1234);
and U8968 (N_8968,N_1644,N_1339);
or U8969 (N_8969,N_111,N_3192);
xor U8970 (N_8970,N_1195,N_4552);
nand U8971 (N_8971,N_3586,N_2797);
nand U8972 (N_8972,N_3837,N_2092);
xor U8973 (N_8973,N_4731,N_509);
or U8974 (N_8974,N_764,N_1916);
xor U8975 (N_8975,N_590,N_4903);
and U8976 (N_8976,N_4079,N_2894);
and U8977 (N_8977,N_2251,N_865);
nand U8978 (N_8978,N_2336,N_155);
nand U8979 (N_8979,N_3461,N_4645);
or U8980 (N_8980,N_1146,N_2519);
nor U8981 (N_8981,N_3358,N_3196);
nor U8982 (N_8982,N_200,N_386);
nand U8983 (N_8983,N_2155,N_3507);
nor U8984 (N_8984,N_1366,N_2720);
xnor U8985 (N_8985,N_4015,N_4689);
or U8986 (N_8986,N_614,N_3248);
or U8987 (N_8987,N_156,N_2609);
or U8988 (N_8988,N_277,N_1731);
or U8989 (N_8989,N_2779,N_4062);
or U8990 (N_8990,N_1127,N_3781);
or U8991 (N_8991,N_953,N_2148);
and U8992 (N_8992,N_900,N_2197);
nor U8993 (N_8993,N_2508,N_4083);
and U8994 (N_8994,N_1995,N_3297);
nand U8995 (N_8995,N_2058,N_509);
and U8996 (N_8996,N_182,N_3655);
nand U8997 (N_8997,N_4464,N_1825);
or U8998 (N_8998,N_1601,N_1886);
or U8999 (N_8999,N_1772,N_2148);
and U9000 (N_9000,N_916,N_939);
and U9001 (N_9001,N_4823,N_4416);
or U9002 (N_9002,N_4723,N_1777);
xor U9003 (N_9003,N_4625,N_2430);
or U9004 (N_9004,N_3151,N_1417);
nor U9005 (N_9005,N_4060,N_2143);
xnor U9006 (N_9006,N_3975,N_1753);
nand U9007 (N_9007,N_431,N_332);
or U9008 (N_9008,N_4893,N_303);
and U9009 (N_9009,N_1399,N_2674);
nand U9010 (N_9010,N_4845,N_1714);
nor U9011 (N_9011,N_1095,N_4669);
xor U9012 (N_9012,N_4357,N_706);
nand U9013 (N_9013,N_163,N_4807);
and U9014 (N_9014,N_4721,N_976);
nor U9015 (N_9015,N_976,N_4171);
or U9016 (N_9016,N_4206,N_4298);
nand U9017 (N_9017,N_907,N_4724);
or U9018 (N_9018,N_626,N_1965);
or U9019 (N_9019,N_4729,N_1665);
nor U9020 (N_9020,N_4253,N_2244);
xor U9021 (N_9021,N_688,N_1828);
xor U9022 (N_9022,N_1732,N_2688);
xnor U9023 (N_9023,N_2820,N_3089);
and U9024 (N_9024,N_289,N_4129);
nor U9025 (N_9025,N_1337,N_1229);
and U9026 (N_9026,N_4403,N_4441);
nand U9027 (N_9027,N_4032,N_4845);
nor U9028 (N_9028,N_3643,N_4310);
or U9029 (N_9029,N_4691,N_55);
or U9030 (N_9030,N_775,N_912);
or U9031 (N_9031,N_200,N_3847);
and U9032 (N_9032,N_2720,N_3151);
nor U9033 (N_9033,N_3737,N_1134);
and U9034 (N_9034,N_2310,N_1411);
xnor U9035 (N_9035,N_104,N_3882);
nor U9036 (N_9036,N_274,N_1033);
or U9037 (N_9037,N_1480,N_2898);
or U9038 (N_9038,N_4490,N_4091);
xnor U9039 (N_9039,N_2362,N_1478);
nor U9040 (N_9040,N_3983,N_2668);
nor U9041 (N_9041,N_3427,N_1483);
nor U9042 (N_9042,N_4509,N_1677);
and U9043 (N_9043,N_1971,N_4267);
nand U9044 (N_9044,N_2034,N_1746);
nor U9045 (N_9045,N_4643,N_2735);
or U9046 (N_9046,N_3531,N_2848);
nand U9047 (N_9047,N_4441,N_3867);
nand U9048 (N_9048,N_75,N_1516);
nor U9049 (N_9049,N_2859,N_4611);
nor U9050 (N_9050,N_1369,N_2415);
nand U9051 (N_9051,N_3111,N_3270);
nor U9052 (N_9052,N_2631,N_153);
and U9053 (N_9053,N_977,N_790);
xnor U9054 (N_9054,N_4360,N_4391);
and U9055 (N_9055,N_2369,N_4077);
nand U9056 (N_9056,N_786,N_1949);
nand U9057 (N_9057,N_4761,N_1775);
nor U9058 (N_9058,N_4814,N_1122);
nand U9059 (N_9059,N_3438,N_1115);
and U9060 (N_9060,N_4421,N_671);
and U9061 (N_9061,N_854,N_4228);
nor U9062 (N_9062,N_671,N_1605);
nor U9063 (N_9063,N_4489,N_3316);
or U9064 (N_9064,N_2082,N_2517);
nand U9065 (N_9065,N_1782,N_4744);
nor U9066 (N_9066,N_2553,N_1745);
and U9067 (N_9067,N_2917,N_4639);
nor U9068 (N_9068,N_3871,N_4701);
nand U9069 (N_9069,N_1422,N_900);
and U9070 (N_9070,N_4762,N_779);
or U9071 (N_9071,N_3335,N_1443);
nand U9072 (N_9072,N_3027,N_692);
nand U9073 (N_9073,N_708,N_4280);
nor U9074 (N_9074,N_209,N_1779);
and U9075 (N_9075,N_4668,N_3916);
or U9076 (N_9076,N_1241,N_4066);
nor U9077 (N_9077,N_4073,N_4203);
xor U9078 (N_9078,N_1543,N_4085);
and U9079 (N_9079,N_1371,N_537);
nand U9080 (N_9080,N_2155,N_3291);
nor U9081 (N_9081,N_3521,N_2982);
xnor U9082 (N_9082,N_4944,N_4254);
nor U9083 (N_9083,N_3802,N_109);
nand U9084 (N_9084,N_1640,N_4603);
xor U9085 (N_9085,N_4384,N_3116);
nor U9086 (N_9086,N_2150,N_2848);
or U9087 (N_9087,N_2737,N_3251);
nand U9088 (N_9088,N_423,N_2765);
nand U9089 (N_9089,N_1986,N_2243);
xnor U9090 (N_9090,N_4961,N_981);
nand U9091 (N_9091,N_4692,N_2072);
xor U9092 (N_9092,N_3679,N_2748);
and U9093 (N_9093,N_2472,N_1661);
nor U9094 (N_9094,N_3756,N_935);
xor U9095 (N_9095,N_3971,N_1407);
nor U9096 (N_9096,N_575,N_3989);
xor U9097 (N_9097,N_4395,N_2953);
and U9098 (N_9098,N_3306,N_3327);
and U9099 (N_9099,N_1374,N_2193);
nand U9100 (N_9100,N_4280,N_2316);
nor U9101 (N_9101,N_4180,N_4461);
nor U9102 (N_9102,N_2175,N_2355);
and U9103 (N_9103,N_3007,N_811);
nor U9104 (N_9104,N_4262,N_883);
or U9105 (N_9105,N_4419,N_2267);
nand U9106 (N_9106,N_1977,N_628);
or U9107 (N_9107,N_2238,N_2652);
and U9108 (N_9108,N_4848,N_3753);
nand U9109 (N_9109,N_3257,N_3462);
or U9110 (N_9110,N_1564,N_1296);
xor U9111 (N_9111,N_244,N_4030);
xnor U9112 (N_9112,N_1315,N_1482);
nor U9113 (N_9113,N_4659,N_4140);
xnor U9114 (N_9114,N_2102,N_2254);
xnor U9115 (N_9115,N_1169,N_1245);
xor U9116 (N_9116,N_4507,N_3820);
xnor U9117 (N_9117,N_2971,N_5);
and U9118 (N_9118,N_615,N_3693);
nor U9119 (N_9119,N_3895,N_772);
or U9120 (N_9120,N_2308,N_4101);
and U9121 (N_9121,N_767,N_4064);
nor U9122 (N_9122,N_108,N_2110);
xnor U9123 (N_9123,N_3006,N_1535);
and U9124 (N_9124,N_3423,N_2528);
and U9125 (N_9125,N_1475,N_362);
and U9126 (N_9126,N_4488,N_147);
xor U9127 (N_9127,N_4692,N_3518);
or U9128 (N_9128,N_585,N_1817);
and U9129 (N_9129,N_3971,N_4954);
nand U9130 (N_9130,N_410,N_1625);
xor U9131 (N_9131,N_2481,N_2233);
nor U9132 (N_9132,N_3846,N_2934);
or U9133 (N_9133,N_452,N_1499);
or U9134 (N_9134,N_735,N_1321);
xor U9135 (N_9135,N_3100,N_315);
nand U9136 (N_9136,N_2359,N_2967);
and U9137 (N_9137,N_3516,N_2564);
and U9138 (N_9138,N_2826,N_1074);
nor U9139 (N_9139,N_534,N_1768);
nand U9140 (N_9140,N_2280,N_2983);
and U9141 (N_9141,N_1276,N_2301);
or U9142 (N_9142,N_3763,N_2914);
xor U9143 (N_9143,N_4903,N_657);
xnor U9144 (N_9144,N_1370,N_3192);
xnor U9145 (N_9145,N_3412,N_1713);
or U9146 (N_9146,N_3493,N_3212);
xor U9147 (N_9147,N_466,N_1236);
nand U9148 (N_9148,N_2005,N_1907);
or U9149 (N_9149,N_1245,N_4798);
xor U9150 (N_9150,N_402,N_186);
nor U9151 (N_9151,N_911,N_834);
nand U9152 (N_9152,N_3845,N_3510);
xor U9153 (N_9153,N_380,N_1573);
xor U9154 (N_9154,N_2593,N_2729);
and U9155 (N_9155,N_2101,N_2454);
nor U9156 (N_9156,N_2786,N_4371);
xnor U9157 (N_9157,N_4312,N_49);
or U9158 (N_9158,N_2641,N_2979);
nand U9159 (N_9159,N_2922,N_4782);
xnor U9160 (N_9160,N_4434,N_759);
xor U9161 (N_9161,N_4441,N_4102);
xor U9162 (N_9162,N_3276,N_3237);
xor U9163 (N_9163,N_4091,N_4786);
nor U9164 (N_9164,N_590,N_1621);
nor U9165 (N_9165,N_204,N_2684);
and U9166 (N_9166,N_4494,N_3896);
nor U9167 (N_9167,N_1748,N_1088);
nand U9168 (N_9168,N_3502,N_136);
or U9169 (N_9169,N_3882,N_3496);
nand U9170 (N_9170,N_2013,N_1960);
or U9171 (N_9171,N_3051,N_1327);
or U9172 (N_9172,N_4498,N_4061);
xnor U9173 (N_9173,N_1896,N_3693);
nand U9174 (N_9174,N_3615,N_3);
nand U9175 (N_9175,N_1544,N_3776);
and U9176 (N_9176,N_4693,N_164);
nor U9177 (N_9177,N_2307,N_1863);
nand U9178 (N_9178,N_860,N_3292);
nor U9179 (N_9179,N_1417,N_423);
nand U9180 (N_9180,N_2959,N_4839);
nor U9181 (N_9181,N_1005,N_2155);
and U9182 (N_9182,N_3196,N_2461);
nand U9183 (N_9183,N_360,N_4502);
or U9184 (N_9184,N_2021,N_2607);
and U9185 (N_9185,N_2,N_264);
xnor U9186 (N_9186,N_3568,N_4101);
xor U9187 (N_9187,N_1973,N_4731);
xnor U9188 (N_9188,N_2181,N_1434);
xor U9189 (N_9189,N_3194,N_1479);
or U9190 (N_9190,N_4570,N_637);
or U9191 (N_9191,N_1966,N_1162);
xor U9192 (N_9192,N_832,N_3316);
xor U9193 (N_9193,N_4021,N_3277);
or U9194 (N_9194,N_1119,N_957);
xor U9195 (N_9195,N_4920,N_249);
or U9196 (N_9196,N_928,N_3649);
and U9197 (N_9197,N_3726,N_3184);
nand U9198 (N_9198,N_731,N_3361);
or U9199 (N_9199,N_3763,N_1908);
nor U9200 (N_9200,N_3361,N_2432);
xor U9201 (N_9201,N_3592,N_2036);
and U9202 (N_9202,N_2576,N_4371);
nand U9203 (N_9203,N_3160,N_2116);
or U9204 (N_9204,N_2135,N_4318);
xnor U9205 (N_9205,N_2158,N_1932);
nand U9206 (N_9206,N_1041,N_144);
and U9207 (N_9207,N_1670,N_4737);
xnor U9208 (N_9208,N_1058,N_2675);
and U9209 (N_9209,N_3456,N_2601);
or U9210 (N_9210,N_4501,N_20);
or U9211 (N_9211,N_8,N_1919);
or U9212 (N_9212,N_2713,N_168);
or U9213 (N_9213,N_3021,N_2935);
nand U9214 (N_9214,N_3688,N_1095);
or U9215 (N_9215,N_2239,N_4319);
nor U9216 (N_9216,N_2670,N_2079);
nor U9217 (N_9217,N_1773,N_3333);
or U9218 (N_9218,N_2740,N_3695);
or U9219 (N_9219,N_4644,N_1614);
and U9220 (N_9220,N_46,N_4766);
and U9221 (N_9221,N_2308,N_4758);
nor U9222 (N_9222,N_2052,N_3259);
nand U9223 (N_9223,N_1676,N_3171);
nor U9224 (N_9224,N_1167,N_3031);
nand U9225 (N_9225,N_2856,N_1128);
xor U9226 (N_9226,N_4646,N_1669);
or U9227 (N_9227,N_3193,N_1123);
nand U9228 (N_9228,N_4780,N_2855);
xnor U9229 (N_9229,N_4147,N_4391);
xor U9230 (N_9230,N_4100,N_2096);
xnor U9231 (N_9231,N_970,N_2633);
or U9232 (N_9232,N_2332,N_3430);
nand U9233 (N_9233,N_3152,N_4866);
or U9234 (N_9234,N_1129,N_3552);
or U9235 (N_9235,N_2673,N_3625);
xnor U9236 (N_9236,N_1812,N_4336);
and U9237 (N_9237,N_2467,N_3262);
xnor U9238 (N_9238,N_691,N_70);
nor U9239 (N_9239,N_4423,N_2271);
nand U9240 (N_9240,N_1548,N_4913);
and U9241 (N_9241,N_1817,N_1968);
or U9242 (N_9242,N_1334,N_4152);
xor U9243 (N_9243,N_884,N_4232);
xnor U9244 (N_9244,N_3341,N_4180);
and U9245 (N_9245,N_2336,N_4294);
and U9246 (N_9246,N_4481,N_810);
xor U9247 (N_9247,N_1222,N_650);
xor U9248 (N_9248,N_3792,N_3265);
and U9249 (N_9249,N_1399,N_4697);
xor U9250 (N_9250,N_2887,N_3033);
xor U9251 (N_9251,N_1646,N_4215);
or U9252 (N_9252,N_3380,N_2968);
and U9253 (N_9253,N_3121,N_4157);
nor U9254 (N_9254,N_173,N_1885);
and U9255 (N_9255,N_1101,N_1055);
or U9256 (N_9256,N_232,N_3380);
or U9257 (N_9257,N_600,N_1831);
nor U9258 (N_9258,N_4473,N_3493);
and U9259 (N_9259,N_2904,N_3364);
nor U9260 (N_9260,N_1029,N_835);
or U9261 (N_9261,N_3334,N_3435);
nand U9262 (N_9262,N_3770,N_1846);
nor U9263 (N_9263,N_1050,N_2757);
nor U9264 (N_9264,N_1439,N_1668);
xor U9265 (N_9265,N_1700,N_3441);
nand U9266 (N_9266,N_1661,N_1448);
or U9267 (N_9267,N_4600,N_1820);
and U9268 (N_9268,N_1082,N_2244);
and U9269 (N_9269,N_4898,N_1129);
nand U9270 (N_9270,N_4848,N_4649);
xor U9271 (N_9271,N_1425,N_1555);
or U9272 (N_9272,N_1068,N_1679);
nand U9273 (N_9273,N_3071,N_1216);
xor U9274 (N_9274,N_207,N_247);
and U9275 (N_9275,N_1710,N_4349);
or U9276 (N_9276,N_116,N_879);
nor U9277 (N_9277,N_1122,N_2333);
or U9278 (N_9278,N_3361,N_3365);
nand U9279 (N_9279,N_4498,N_3738);
xnor U9280 (N_9280,N_2842,N_2575);
nand U9281 (N_9281,N_967,N_1834);
and U9282 (N_9282,N_3984,N_2528);
nor U9283 (N_9283,N_3789,N_1523);
nor U9284 (N_9284,N_4600,N_2735);
nor U9285 (N_9285,N_1743,N_2894);
nand U9286 (N_9286,N_3805,N_2813);
nand U9287 (N_9287,N_3021,N_4328);
nor U9288 (N_9288,N_1476,N_3148);
or U9289 (N_9289,N_323,N_4591);
or U9290 (N_9290,N_2459,N_3379);
nand U9291 (N_9291,N_88,N_4957);
xor U9292 (N_9292,N_1888,N_1349);
nand U9293 (N_9293,N_3918,N_3654);
nand U9294 (N_9294,N_1505,N_2315);
and U9295 (N_9295,N_763,N_733);
nor U9296 (N_9296,N_4494,N_4536);
and U9297 (N_9297,N_4078,N_2991);
xnor U9298 (N_9298,N_851,N_4806);
or U9299 (N_9299,N_3900,N_2981);
nor U9300 (N_9300,N_1556,N_3794);
nand U9301 (N_9301,N_4439,N_3963);
xor U9302 (N_9302,N_667,N_3174);
nand U9303 (N_9303,N_2555,N_4468);
xor U9304 (N_9304,N_3825,N_2616);
nand U9305 (N_9305,N_113,N_1477);
nand U9306 (N_9306,N_3181,N_4514);
and U9307 (N_9307,N_2217,N_2459);
or U9308 (N_9308,N_4471,N_2593);
and U9309 (N_9309,N_2708,N_1220);
or U9310 (N_9310,N_3094,N_3396);
nand U9311 (N_9311,N_4294,N_4841);
xnor U9312 (N_9312,N_3521,N_664);
xor U9313 (N_9313,N_2424,N_2373);
or U9314 (N_9314,N_2178,N_1636);
nand U9315 (N_9315,N_3815,N_1175);
nor U9316 (N_9316,N_1279,N_4907);
xnor U9317 (N_9317,N_4983,N_1169);
nor U9318 (N_9318,N_3339,N_3301);
and U9319 (N_9319,N_1306,N_3041);
xnor U9320 (N_9320,N_4020,N_2554);
and U9321 (N_9321,N_197,N_3955);
or U9322 (N_9322,N_2927,N_1582);
or U9323 (N_9323,N_2228,N_4691);
nand U9324 (N_9324,N_2517,N_4540);
and U9325 (N_9325,N_4110,N_2950);
or U9326 (N_9326,N_1845,N_3155);
nand U9327 (N_9327,N_1800,N_1889);
or U9328 (N_9328,N_2430,N_2742);
or U9329 (N_9329,N_783,N_2433);
and U9330 (N_9330,N_3982,N_1789);
nor U9331 (N_9331,N_1884,N_3055);
and U9332 (N_9332,N_1204,N_3944);
and U9333 (N_9333,N_98,N_1089);
or U9334 (N_9334,N_285,N_553);
xnor U9335 (N_9335,N_3899,N_2398);
nand U9336 (N_9336,N_352,N_3842);
nand U9337 (N_9337,N_3234,N_35);
nand U9338 (N_9338,N_2618,N_4977);
nor U9339 (N_9339,N_1907,N_3358);
or U9340 (N_9340,N_598,N_3218);
nand U9341 (N_9341,N_1972,N_916);
xnor U9342 (N_9342,N_4593,N_2803);
or U9343 (N_9343,N_1986,N_4731);
or U9344 (N_9344,N_1684,N_587);
nand U9345 (N_9345,N_1425,N_3428);
and U9346 (N_9346,N_1605,N_1677);
xor U9347 (N_9347,N_1099,N_1990);
xnor U9348 (N_9348,N_4474,N_4801);
xor U9349 (N_9349,N_2049,N_1612);
or U9350 (N_9350,N_1901,N_4043);
nor U9351 (N_9351,N_470,N_4299);
nor U9352 (N_9352,N_770,N_4219);
xnor U9353 (N_9353,N_1763,N_1080);
nand U9354 (N_9354,N_4034,N_3860);
or U9355 (N_9355,N_870,N_1885);
and U9356 (N_9356,N_3493,N_2529);
nor U9357 (N_9357,N_335,N_1929);
nand U9358 (N_9358,N_3678,N_2063);
nand U9359 (N_9359,N_4229,N_1124);
nor U9360 (N_9360,N_4300,N_2275);
nand U9361 (N_9361,N_824,N_4330);
nand U9362 (N_9362,N_4853,N_1080);
xor U9363 (N_9363,N_2332,N_3812);
xnor U9364 (N_9364,N_4615,N_3568);
and U9365 (N_9365,N_410,N_2040);
nand U9366 (N_9366,N_1185,N_4642);
nor U9367 (N_9367,N_3381,N_4752);
nand U9368 (N_9368,N_203,N_3526);
or U9369 (N_9369,N_1490,N_323);
or U9370 (N_9370,N_3840,N_4553);
and U9371 (N_9371,N_1759,N_326);
xnor U9372 (N_9372,N_1188,N_771);
xnor U9373 (N_9373,N_4452,N_2885);
and U9374 (N_9374,N_748,N_1393);
nor U9375 (N_9375,N_3872,N_676);
or U9376 (N_9376,N_2803,N_3713);
nor U9377 (N_9377,N_136,N_4493);
xnor U9378 (N_9378,N_4813,N_4728);
nand U9379 (N_9379,N_1887,N_3956);
nor U9380 (N_9380,N_1602,N_1391);
and U9381 (N_9381,N_4069,N_2409);
xor U9382 (N_9382,N_1251,N_1672);
or U9383 (N_9383,N_3584,N_56);
nor U9384 (N_9384,N_3533,N_3282);
xor U9385 (N_9385,N_4614,N_4246);
nand U9386 (N_9386,N_720,N_1958);
xor U9387 (N_9387,N_2983,N_971);
xor U9388 (N_9388,N_427,N_3189);
or U9389 (N_9389,N_1171,N_2764);
xnor U9390 (N_9390,N_1140,N_1754);
xor U9391 (N_9391,N_4304,N_3167);
nand U9392 (N_9392,N_2629,N_693);
and U9393 (N_9393,N_1642,N_351);
and U9394 (N_9394,N_3551,N_3591);
or U9395 (N_9395,N_1139,N_3085);
nand U9396 (N_9396,N_262,N_3200);
nor U9397 (N_9397,N_3851,N_2236);
nor U9398 (N_9398,N_4057,N_3052);
xnor U9399 (N_9399,N_4859,N_781);
and U9400 (N_9400,N_3832,N_3462);
and U9401 (N_9401,N_3115,N_3074);
or U9402 (N_9402,N_1214,N_4280);
nor U9403 (N_9403,N_4908,N_1016);
xnor U9404 (N_9404,N_2213,N_3248);
or U9405 (N_9405,N_3082,N_628);
xnor U9406 (N_9406,N_4132,N_4530);
and U9407 (N_9407,N_785,N_2499);
or U9408 (N_9408,N_124,N_2682);
and U9409 (N_9409,N_1102,N_4841);
xor U9410 (N_9410,N_2215,N_1021);
or U9411 (N_9411,N_1702,N_2774);
nor U9412 (N_9412,N_4929,N_1710);
nor U9413 (N_9413,N_93,N_2546);
nor U9414 (N_9414,N_3441,N_2363);
or U9415 (N_9415,N_509,N_4852);
nand U9416 (N_9416,N_23,N_2443);
nor U9417 (N_9417,N_4159,N_986);
or U9418 (N_9418,N_10,N_1385);
nor U9419 (N_9419,N_4518,N_3977);
nand U9420 (N_9420,N_2620,N_3926);
nor U9421 (N_9421,N_4647,N_3885);
and U9422 (N_9422,N_3629,N_2647);
and U9423 (N_9423,N_256,N_1049);
or U9424 (N_9424,N_1257,N_2298);
nand U9425 (N_9425,N_2768,N_2872);
or U9426 (N_9426,N_4004,N_4772);
xnor U9427 (N_9427,N_2120,N_3267);
xnor U9428 (N_9428,N_2840,N_2894);
nand U9429 (N_9429,N_276,N_509);
xnor U9430 (N_9430,N_4279,N_2028);
and U9431 (N_9431,N_865,N_3689);
nor U9432 (N_9432,N_2643,N_242);
and U9433 (N_9433,N_4887,N_4356);
nor U9434 (N_9434,N_328,N_1769);
xor U9435 (N_9435,N_3890,N_3571);
nor U9436 (N_9436,N_3208,N_3778);
nand U9437 (N_9437,N_4939,N_2051);
nand U9438 (N_9438,N_3646,N_2863);
or U9439 (N_9439,N_1717,N_2568);
and U9440 (N_9440,N_3792,N_1695);
nand U9441 (N_9441,N_1546,N_3166);
or U9442 (N_9442,N_1684,N_3754);
xor U9443 (N_9443,N_121,N_850);
nand U9444 (N_9444,N_1374,N_4120);
and U9445 (N_9445,N_1607,N_1263);
or U9446 (N_9446,N_2184,N_2334);
and U9447 (N_9447,N_1501,N_1564);
nand U9448 (N_9448,N_2539,N_1661);
and U9449 (N_9449,N_1132,N_1537);
and U9450 (N_9450,N_502,N_2287);
nand U9451 (N_9451,N_957,N_445);
and U9452 (N_9452,N_96,N_4521);
and U9453 (N_9453,N_242,N_860);
nor U9454 (N_9454,N_338,N_674);
xnor U9455 (N_9455,N_4950,N_2496);
nand U9456 (N_9456,N_263,N_3166);
nor U9457 (N_9457,N_3867,N_755);
or U9458 (N_9458,N_213,N_4185);
nand U9459 (N_9459,N_1815,N_1299);
nand U9460 (N_9460,N_4386,N_2099);
nor U9461 (N_9461,N_1393,N_249);
nor U9462 (N_9462,N_3945,N_2983);
nand U9463 (N_9463,N_409,N_3560);
and U9464 (N_9464,N_3913,N_4802);
and U9465 (N_9465,N_3354,N_3544);
and U9466 (N_9466,N_4912,N_2374);
nor U9467 (N_9467,N_3723,N_4694);
and U9468 (N_9468,N_3100,N_3737);
nor U9469 (N_9469,N_1500,N_4629);
nor U9470 (N_9470,N_1136,N_3789);
and U9471 (N_9471,N_331,N_4171);
nand U9472 (N_9472,N_41,N_3511);
or U9473 (N_9473,N_1216,N_2496);
nand U9474 (N_9474,N_2085,N_150);
nor U9475 (N_9475,N_1504,N_1758);
nand U9476 (N_9476,N_1769,N_3947);
nand U9477 (N_9477,N_3132,N_4631);
and U9478 (N_9478,N_2028,N_1544);
nor U9479 (N_9479,N_2061,N_3253);
nand U9480 (N_9480,N_4481,N_732);
or U9481 (N_9481,N_814,N_2514);
or U9482 (N_9482,N_4706,N_2462);
nor U9483 (N_9483,N_4441,N_2527);
or U9484 (N_9484,N_3159,N_2577);
nand U9485 (N_9485,N_2128,N_2020);
or U9486 (N_9486,N_2493,N_4816);
or U9487 (N_9487,N_3959,N_3021);
nand U9488 (N_9488,N_397,N_2313);
and U9489 (N_9489,N_462,N_1459);
xor U9490 (N_9490,N_1477,N_4072);
nand U9491 (N_9491,N_847,N_4410);
xor U9492 (N_9492,N_3724,N_4336);
nor U9493 (N_9493,N_2981,N_838);
nand U9494 (N_9494,N_4894,N_4612);
nand U9495 (N_9495,N_1461,N_2945);
xnor U9496 (N_9496,N_1217,N_4005);
nor U9497 (N_9497,N_1933,N_4152);
or U9498 (N_9498,N_94,N_504);
nor U9499 (N_9499,N_3794,N_4912);
and U9500 (N_9500,N_1833,N_1188);
xor U9501 (N_9501,N_975,N_895);
nand U9502 (N_9502,N_1950,N_4044);
nor U9503 (N_9503,N_4791,N_650);
and U9504 (N_9504,N_2425,N_2533);
and U9505 (N_9505,N_4060,N_3565);
nand U9506 (N_9506,N_3628,N_1710);
xnor U9507 (N_9507,N_4895,N_1237);
nand U9508 (N_9508,N_1187,N_4941);
or U9509 (N_9509,N_668,N_3643);
nor U9510 (N_9510,N_4739,N_4435);
and U9511 (N_9511,N_4965,N_2261);
nand U9512 (N_9512,N_831,N_69);
xnor U9513 (N_9513,N_1728,N_1753);
nand U9514 (N_9514,N_1132,N_3697);
nand U9515 (N_9515,N_3700,N_1406);
and U9516 (N_9516,N_843,N_3195);
nor U9517 (N_9517,N_469,N_1530);
or U9518 (N_9518,N_4280,N_4429);
nand U9519 (N_9519,N_4782,N_2843);
nor U9520 (N_9520,N_186,N_1009);
or U9521 (N_9521,N_4334,N_3055);
or U9522 (N_9522,N_2924,N_1704);
or U9523 (N_9523,N_471,N_4385);
nand U9524 (N_9524,N_2933,N_1390);
xnor U9525 (N_9525,N_3859,N_2464);
or U9526 (N_9526,N_201,N_3115);
nand U9527 (N_9527,N_1547,N_3906);
xor U9528 (N_9528,N_3719,N_3228);
or U9529 (N_9529,N_4169,N_4111);
or U9530 (N_9530,N_744,N_3395);
and U9531 (N_9531,N_4429,N_173);
or U9532 (N_9532,N_2228,N_2423);
and U9533 (N_9533,N_4222,N_3416);
and U9534 (N_9534,N_4953,N_4197);
and U9535 (N_9535,N_3595,N_642);
or U9536 (N_9536,N_2245,N_2004);
xor U9537 (N_9537,N_1944,N_3256);
xnor U9538 (N_9538,N_174,N_3287);
xnor U9539 (N_9539,N_3340,N_2534);
nor U9540 (N_9540,N_2575,N_2336);
nand U9541 (N_9541,N_1586,N_1062);
nand U9542 (N_9542,N_2278,N_2586);
nor U9543 (N_9543,N_4286,N_910);
or U9544 (N_9544,N_1532,N_4512);
and U9545 (N_9545,N_340,N_66);
nor U9546 (N_9546,N_223,N_3804);
and U9547 (N_9547,N_4710,N_4762);
nand U9548 (N_9548,N_442,N_1832);
xor U9549 (N_9549,N_1365,N_4134);
nand U9550 (N_9550,N_1403,N_1491);
and U9551 (N_9551,N_1491,N_1365);
nor U9552 (N_9552,N_2177,N_3090);
xor U9553 (N_9553,N_1344,N_3660);
nor U9554 (N_9554,N_1693,N_1098);
and U9555 (N_9555,N_4655,N_3484);
nor U9556 (N_9556,N_1908,N_4845);
nand U9557 (N_9557,N_633,N_4283);
nor U9558 (N_9558,N_934,N_1325);
or U9559 (N_9559,N_491,N_3942);
and U9560 (N_9560,N_4009,N_3727);
or U9561 (N_9561,N_447,N_2445);
or U9562 (N_9562,N_1999,N_1752);
nor U9563 (N_9563,N_2630,N_852);
nor U9564 (N_9564,N_3502,N_411);
xnor U9565 (N_9565,N_22,N_3617);
and U9566 (N_9566,N_4344,N_4849);
nor U9567 (N_9567,N_170,N_1597);
nand U9568 (N_9568,N_4029,N_2037);
or U9569 (N_9569,N_2072,N_3500);
nor U9570 (N_9570,N_1049,N_272);
nor U9571 (N_9571,N_847,N_3267);
nand U9572 (N_9572,N_2232,N_2289);
and U9573 (N_9573,N_4275,N_193);
nor U9574 (N_9574,N_1789,N_4918);
nand U9575 (N_9575,N_249,N_2001);
and U9576 (N_9576,N_1013,N_4017);
nor U9577 (N_9577,N_2332,N_1740);
xnor U9578 (N_9578,N_3646,N_913);
nor U9579 (N_9579,N_760,N_4074);
and U9580 (N_9580,N_1129,N_628);
nand U9581 (N_9581,N_3723,N_3410);
nand U9582 (N_9582,N_4396,N_3244);
xor U9583 (N_9583,N_818,N_103);
nor U9584 (N_9584,N_27,N_3221);
xnor U9585 (N_9585,N_337,N_240);
nand U9586 (N_9586,N_2024,N_1463);
nand U9587 (N_9587,N_3050,N_4076);
and U9588 (N_9588,N_416,N_4344);
or U9589 (N_9589,N_1250,N_2623);
and U9590 (N_9590,N_3018,N_3901);
nand U9591 (N_9591,N_144,N_2550);
or U9592 (N_9592,N_4356,N_1693);
and U9593 (N_9593,N_1446,N_3189);
nor U9594 (N_9594,N_3308,N_711);
nor U9595 (N_9595,N_309,N_4065);
xnor U9596 (N_9596,N_87,N_1229);
nor U9597 (N_9597,N_3858,N_272);
or U9598 (N_9598,N_532,N_2116);
xnor U9599 (N_9599,N_1069,N_3111);
nor U9600 (N_9600,N_3879,N_34);
nand U9601 (N_9601,N_4801,N_1207);
nand U9602 (N_9602,N_3741,N_2947);
or U9603 (N_9603,N_3013,N_2783);
or U9604 (N_9604,N_198,N_455);
nor U9605 (N_9605,N_2086,N_3531);
nand U9606 (N_9606,N_3346,N_2348);
xnor U9607 (N_9607,N_3363,N_2504);
nor U9608 (N_9608,N_134,N_3214);
xnor U9609 (N_9609,N_2419,N_1487);
nand U9610 (N_9610,N_2415,N_4061);
and U9611 (N_9611,N_528,N_2679);
xor U9612 (N_9612,N_2160,N_3625);
or U9613 (N_9613,N_2139,N_2805);
or U9614 (N_9614,N_1901,N_4670);
nand U9615 (N_9615,N_4386,N_3839);
xor U9616 (N_9616,N_1887,N_4967);
and U9617 (N_9617,N_1454,N_3615);
nor U9618 (N_9618,N_1467,N_2648);
nand U9619 (N_9619,N_1065,N_2074);
and U9620 (N_9620,N_4146,N_4275);
xnor U9621 (N_9621,N_2963,N_4567);
or U9622 (N_9622,N_1573,N_493);
nor U9623 (N_9623,N_1338,N_4086);
and U9624 (N_9624,N_2295,N_1986);
xnor U9625 (N_9625,N_3909,N_3311);
nand U9626 (N_9626,N_3366,N_2418);
nand U9627 (N_9627,N_3248,N_3361);
and U9628 (N_9628,N_2638,N_380);
or U9629 (N_9629,N_2625,N_403);
or U9630 (N_9630,N_3858,N_4941);
or U9631 (N_9631,N_4359,N_4154);
xnor U9632 (N_9632,N_4022,N_3447);
xor U9633 (N_9633,N_892,N_1599);
xnor U9634 (N_9634,N_145,N_1364);
xnor U9635 (N_9635,N_1458,N_2117);
and U9636 (N_9636,N_3609,N_3717);
nand U9637 (N_9637,N_4003,N_1581);
and U9638 (N_9638,N_1923,N_1396);
nand U9639 (N_9639,N_4690,N_1097);
nor U9640 (N_9640,N_2779,N_4416);
nor U9641 (N_9641,N_1115,N_4797);
or U9642 (N_9642,N_868,N_1333);
and U9643 (N_9643,N_4287,N_208);
nor U9644 (N_9644,N_3254,N_4860);
xnor U9645 (N_9645,N_2111,N_1099);
or U9646 (N_9646,N_3331,N_655);
and U9647 (N_9647,N_3152,N_2792);
xnor U9648 (N_9648,N_2628,N_3646);
nor U9649 (N_9649,N_4307,N_3138);
and U9650 (N_9650,N_3693,N_1073);
xnor U9651 (N_9651,N_726,N_784);
nand U9652 (N_9652,N_4281,N_226);
nor U9653 (N_9653,N_711,N_162);
xnor U9654 (N_9654,N_774,N_4426);
xnor U9655 (N_9655,N_156,N_2300);
nor U9656 (N_9656,N_447,N_4958);
and U9657 (N_9657,N_4873,N_2067);
xnor U9658 (N_9658,N_241,N_227);
nor U9659 (N_9659,N_4859,N_2850);
xor U9660 (N_9660,N_2100,N_165);
xnor U9661 (N_9661,N_1010,N_3352);
xnor U9662 (N_9662,N_2113,N_4662);
nand U9663 (N_9663,N_3657,N_1699);
nand U9664 (N_9664,N_3612,N_2026);
xor U9665 (N_9665,N_1632,N_2166);
and U9666 (N_9666,N_3460,N_1274);
nor U9667 (N_9667,N_3482,N_1099);
nand U9668 (N_9668,N_122,N_4148);
and U9669 (N_9669,N_1155,N_2886);
nand U9670 (N_9670,N_3659,N_3745);
and U9671 (N_9671,N_2538,N_4290);
nand U9672 (N_9672,N_3380,N_1568);
and U9673 (N_9673,N_1210,N_3946);
xor U9674 (N_9674,N_954,N_1674);
xnor U9675 (N_9675,N_1895,N_3835);
nor U9676 (N_9676,N_4409,N_4928);
nor U9677 (N_9677,N_4829,N_541);
nor U9678 (N_9678,N_247,N_1528);
nor U9679 (N_9679,N_3155,N_1560);
or U9680 (N_9680,N_4007,N_1159);
nor U9681 (N_9681,N_1407,N_4034);
or U9682 (N_9682,N_983,N_2534);
xnor U9683 (N_9683,N_3825,N_2477);
xnor U9684 (N_9684,N_4408,N_1276);
nor U9685 (N_9685,N_4436,N_71);
nor U9686 (N_9686,N_906,N_293);
nor U9687 (N_9687,N_325,N_3813);
and U9688 (N_9688,N_1750,N_685);
nor U9689 (N_9689,N_3400,N_4430);
nor U9690 (N_9690,N_2277,N_3716);
nand U9691 (N_9691,N_4130,N_3193);
nand U9692 (N_9692,N_3165,N_4086);
and U9693 (N_9693,N_4762,N_1546);
and U9694 (N_9694,N_309,N_4688);
nand U9695 (N_9695,N_3066,N_3324);
xor U9696 (N_9696,N_253,N_4392);
xor U9697 (N_9697,N_678,N_4598);
xnor U9698 (N_9698,N_361,N_3250);
xor U9699 (N_9699,N_923,N_2457);
xnor U9700 (N_9700,N_4008,N_1092);
nor U9701 (N_9701,N_414,N_1980);
nand U9702 (N_9702,N_4599,N_2595);
nand U9703 (N_9703,N_1124,N_2972);
and U9704 (N_9704,N_3629,N_32);
and U9705 (N_9705,N_2173,N_609);
or U9706 (N_9706,N_3786,N_3945);
and U9707 (N_9707,N_2438,N_3486);
xnor U9708 (N_9708,N_2957,N_1340);
xor U9709 (N_9709,N_539,N_2470);
xnor U9710 (N_9710,N_4104,N_1729);
xor U9711 (N_9711,N_3163,N_3318);
nor U9712 (N_9712,N_491,N_3372);
and U9713 (N_9713,N_3113,N_1335);
or U9714 (N_9714,N_4515,N_4431);
xor U9715 (N_9715,N_1303,N_4208);
or U9716 (N_9716,N_1560,N_2302);
and U9717 (N_9717,N_4193,N_4561);
nand U9718 (N_9718,N_1059,N_842);
or U9719 (N_9719,N_385,N_621);
nor U9720 (N_9720,N_3651,N_1135);
and U9721 (N_9721,N_3504,N_2398);
and U9722 (N_9722,N_664,N_4233);
or U9723 (N_9723,N_649,N_1948);
xor U9724 (N_9724,N_3673,N_1743);
nor U9725 (N_9725,N_4093,N_2269);
nor U9726 (N_9726,N_2428,N_2826);
and U9727 (N_9727,N_4342,N_3340);
xor U9728 (N_9728,N_937,N_751);
xor U9729 (N_9729,N_1239,N_4100);
and U9730 (N_9730,N_4027,N_4489);
xnor U9731 (N_9731,N_2270,N_3550);
and U9732 (N_9732,N_4256,N_4958);
or U9733 (N_9733,N_1245,N_1620);
xor U9734 (N_9734,N_3702,N_1523);
xnor U9735 (N_9735,N_2760,N_1808);
or U9736 (N_9736,N_1655,N_4926);
nor U9737 (N_9737,N_1026,N_1827);
nand U9738 (N_9738,N_4643,N_1877);
xor U9739 (N_9739,N_1369,N_2216);
or U9740 (N_9740,N_4633,N_4705);
or U9741 (N_9741,N_480,N_4210);
xor U9742 (N_9742,N_4257,N_2560);
xor U9743 (N_9743,N_4730,N_3083);
and U9744 (N_9744,N_1922,N_2255);
and U9745 (N_9745,N_3093,N_3343);
or U9746 (N_9746,N_1577,N_845);
xnor U9747 (N_9747,N_4395,N_3941);
or U9748 (N_9748,N_2666,N_2347);
xor U9749 (N_9749,N_2063,N_4768);
and U9750 (N_9750,N_601,N_2628);
or U9751 (N_9751,N_3760,N_3070);
or U9752 (N_9752,N_2074,N_1019);
xor U9753 (N_9753,N_2584,N_1498);
xor U9754 (N_9754,N_832,N_200);
or U9755 (N_9755,N_1712,N_3970);
xor U9756 (N_9756,N_3817,N_2112);
xnor U9757 (N_9757,N_3764,N_2751);
xor U9758 (N_9758,N_4066,N_4383);
xnor U9759 (N_9759,N_417,N_2618);
nand U9760 (N_9760,N_483,N_1970);
nand U9761 (N_9761,N_1872,N_2365);
xor U9762 (N_9762,N_232,N_1737);
nand U9763 (N_9763,N_1001,N_845);
nand U9764 (N_9764,N_3595,N_2026);
and U9765 (N_9765,N_4511,N_4340);
nand U9766 (N_9766,N_2633,N_1730);
and U9767 (N_9767,N_228,N_3463);
nand U9768 (N_9768,N_3430,N_3964);
xnor U9769 (N_9769,N_1495,N_113);
nor U9770 (N_9770,N_1562,N_3393);
xor U9771 (N_9771,N_135,N_577);
and U9772 (N_9772,N_4907,N_13);
or U9773 (N_9773,N_4281,N_3354);
xor U9774 (N_9774,N_4124,N_888);
or U9775 (N_9775,N_606,N_2745);
and U9776 (N_9776,N_3955,N_276);
xnor U9777 (N_9777,N_4026,N_4736);
nor U9778 (N_9778,N_2026,N_587);
xor U9779 (N_9779,N_3350,N_1929);
nor U9780 (N_9780,N_981,N_1428);
nand U9781 (N_9781,N_1471,N_4182);
and U9782 (N_9782,N_3201,N_3255);
nor U9783 (N_9783,N_3149,N_3032);
xor U9784 (N_9784,N_3873,N_390);
nand U9785 (N_9785,N_1877,N_3104);
and U9786 (N_9786,N_1269,N_1531);
or U9787 (N_9787,N_387,N_1642);
or U9788 (N_9788,N_28,N_2037);
and U9789 (N_9789,N_3063,N_3030);
nor U9790 (N_9790,N_542,N_1934);
nor U9791 (N_9791,N_3232,N_2970);
xor U9792 (N_9792,N_576,N_4207);
xnor U9793 (N_9793,N_3463,N_4484);
and U9794 (N_9794,N_1273,N_1677);
nand U9795 (N_9795,N_2970,N_4734);
nand U9796 (N_9796,N_2087,N_2411);
or U9797 (N_9797,N_2260,N_1397);
and U9798 (N_9798,N_2812,N_3278);
nand U9799 (N_9799,N_1880,N_3339);
and U9800 (N_9800,N_2537,N_1918);
or U9801 (N_9801,N_1470,N_1405);
xnor U9802 (N_9802,N_140,N_2951);
nand U9803 (N_9803,N_3396,N_755);
and U9804 (N_9804,N_4531,N_892);
nor U9805 (N_9805,N_2052,N_2545);
and U9806 (N_9806,N_2922,N_3704);
or U9807 (N_9807,N_3299,N_1033);
xor U9808 (N_9808,N_3427,N_4922);
nand U9809 (N_9809,N_686,N_4361);
nand U9810 (N_9810,N_2409,N_1892);
and U9811 (N_9811,N_2353,N_1413);
xnor U9812 (N_9812,N_2821,N_2004);
or U9813 (N_9813,N_4414,N_3755);
and U9814 (N_9814,N_2676,N_2461);
xor U9815 (N_9815,N_2278,N_3087);
nand U9816 (N_9816,N_3346,N_1077);
nand U9817 (N_9817,N_4782,N_3558);
xor U9818 (N_9818,N_4078,N_3823);
or U9819 (N_9819,N_1703,N_1901);
nand U9820 (N_9820,N_4190,N_2668);
or U9821 (N_9821,N_2946,N_3140);
nand U9822 (N_9822,N_3372,N_3404);
nor U9823 (N_9823,N_2943,N_3057);
or U9824 (N_9824,N_2742,N_4040);
or U9825 (N_9825,N_2335,N_2862);
or U9826 (N_9826,N_1881,N_2793);
and U9827 (N_9827,N_4231,N_1835);
nand U9828 (N_9828,N_2242,N_2725);
nand U9829 (N_9829,N_4273,N_1299);
or U9830 (N_9830,N_668,N_1738);
nor U9831 (N_9831,N_1835,N_4905);
xor U9832 (N_9832,N_1220,N_243);
or U9833 (N_9833,N_2633,N_240);
and U9834 (N_9834,N_3009,N_1273);
and U9835 (N_9835,N_1515,N_2801);
xor U9836 (N_9836,N_2478,N_1045);
nand U9837 (N_9837,N_1984,N_2053);
and U9838 (N_9838,N_3680,N_2783);
xnor U9839 (N_9839,N_3791,N_3725);
nand U9840 (N_9840,N_1804,N_1026);
and U9841 (N_9841,N_1951,N_2080);
nand U9842 (N_9842,N_2463,N_942);
and U9843 (N_9843,N_1592,N_3985);
and U9844 (N_9844,N_3991,N_892);
nor U9845 (N_9845,N_3473,N_1184);
nor U9846 (N_9846,N_4822,N_1478);
or U9847 (N_9847,N_3964,N_2186);
xor U9848 (N_9848,N_1455,N_3757);
nand U9849 (N_9849,N_4329,N_428);
nor U9850 (N_9850,N_643,N_477);
nor U9851 (N_9851,N_3823,N_351);
nand U9852 (N_9852,N_1308,N_1212);
nor U9853 (N_9853,N_1284,N_4194);
xnor U9854 (N_9854,N_920,N_4825);
nand U9855 (N_9855,N_333,N_3810);
xor U9856 (N_9856,N_73,N_3134);
or U9857 (N_9857,N_1473,N_1086);
or U9858 (N_9858,N_1671,N_1950);
xor U9859 (N_9859,N_658,N_4547);
nor U9860 (N_9860,N_4958,N_1487);
or U9861 (N_9861,N_1378,N_2149);
or U9862 (N_9862,N_1672,N_1402);
and U9863 (N_9863,N_1700,N_1388);
xor U9864 (N_9864,N_1866,N_3051);
and U9865 (N_9865,N_2621,N_3242);
and U9866 (N_9866,N_4286,N_566);
xor U9867 (N_9867,N_3383,N_3390);
or U9868 (N_9868,N_1944,N_3306);
or U9869 (N_9869,N_4159,N_4051);
or U9870 (N_9870,N_2041,N_2821);
and U9871 (N_9871,N_2005,N_4988);
nand U9872 (N_9872,N_1116,N_2257);
nand U9873 (N_9873,N_4869,N_4097);
nand U9874 (N_9874,N_3029,N_4818);
nor U9875 (N_9875,N_191,N_2831);
and U9876 (N_9876,N_3066,N_1839);
xor U9877 (N_9877,N_2581,N_2217);
xnor U9878 (N_9878,N_2171,N_1142);
and U9879 (N_9879,N_3633,N_450);
xor U9880 (N_9880,N_574,N_1021);
and U9881 (N_9881,N_278,N_3720);
or U9882 (N_9882,N_1184,N_2011);
xor U9883 (N_9883,N_671,N_1410);
xnor U9884 (N_9884,N_1225,N_3685);
nand U9885 (N_9885,N_1458,N_1439);
nand U9886 (N_9886,N_696,N_4266);
and U9887 (N_9887,N_2816,N_4772);
and U9888 (N_9888,N_3000,N_4114);
nand U9889 (N_9889,N_551,N_368);
nor U9890 (N_9890,N_768,N_4332);
or U9891 (N_9891,N_65,N_3318);
xor U9892 (N_9892,N_2498,N_4734);
nand U9893 (N_9893,N_4531,N_2261);
or U9894 (N_9894,N_4302,N_745);
and U9895 (N_9895,N_494,N_4167);
nor U9896 (N_9896,N_2548,N_898);
or U9897 (N_9897,N_2382,N_554);
nor U9898 (N_9898,N_4494,N_3806);
nand U9899 (N_9899,N_1791,N_2357);
nor U9900 (N_9900,N_1416,N_4125);
nand U9901 (N_9901,N_4186,N_3081);
nand U9902 (N_9902,N_4306,N_2472);
nand U9903 (N_9903,N_36,N_576);
xor U9904 (N_9904,N_4920,N_241);
and U9905 (N_9905,N_4830,N_2363);
and U9906 (N_9906,N_2524,N_2299);
nor U9907 (N_9907,N_3841,N_1061);
xor U9908 (N_9908,N_4362,N_4618);
nor U9909 (N_9909,N_50,N_2104);
nor U9910 (N_9910,N_4149,N_881);
and U9911 (N_9911,N_4896,N_4516);
and U9912 (N_9912,N_590,N_3829);
nor U9913 (N_9913,N_3678,N_4001);
or U9914 (N_9914,N_215,N_1589);
xor U9915 (N_9915,N_4951,N_2814);
nor U9916 (N_9916,N_4422,N_3846);
xnor U9917 (N_9917,N_232,N_4083);
and U9918 (N_9918,N_3312,N_3949);
and U9919 (N_9919,N_691,N_535);
xnor U9920 (N_9920,N_2518,N_1290);
and U9921 (N_9921,N_1670,N_327);
or U9922 (N_9922,N_3778,N_4405);
nor U9923 (N_9923,N_3038,N_616);
nor U9924 (N_9924,N_3027,N_3004);
or U9925 (N_9925,N_4936,N_3624);
and U9926 (N_9926,N_2301,N_837);
nand U9927 (N_9927,N_1472,N_608);
or U9928 (N_9928,N_2551,N_4690);
xor U9929 (N_9929,N_1052,N_148);
xnor U9930 (N_9930,N_660,N_2818);
xnor U9931 (N_9931,N_3736,N_3481);
nor U9932 (N_9932,N_3137,N_439);
nor U9933 (N_9933,N_43,N_1771);
or U9934 (N_9934,N_872,N_3475);
xnor U9935 (N_9935,N_2332,N_4609);
nand U9936 (N_9936,N_58,N_1067);
nand U9937 (N_9937,N_2033,N_785);
nor U9938 (N_9938,N_1724,N_455);
nor U9939 (N_9939,N_2601,N_4016);
and U9940 (N_9940,N_2340,N_4883);
xor U9941 (N_9941,N_3692,N_3095);
xnor U9942 (N_9942,N_3446,N_4515);
or U9943 (N_9943,N_4120,N_4192);
nor U9944 (N_9944,N_481,N_27);
and U9945 (N_9945,N_831,N_4565);
nand U9946 (N_9946,N_3342,N_3220);
or U9947 (N_9947,N_1637,N_4146);
xor U9948 (N_9948,N_3794,N_3220);
or U9949 (N_9949,N_4373,N_4483);
xnor U9950 (N_9950,N_235,N_3729);
and U9951 (N_9951,N_3048,N_386);
and U9952 (N_9952,N_4662,N_3308);
nand U9953 (N_9953,N_2220,N_280);
and U9954 (N_9954,N_1650,N_1984);
nand U9955 (N_9955,N_3589,N_1069);
and U9956 (N_9956,N_4593,N_486);
and U9957 (N_9957,N_3044,N_2844);
or U9958 (N_9958,N_236,N_1496);
nor U9959 (N_9959,N_2809,N_2980);
nand U9960 (N_9960,N_2023,N_3084);
nor U9961 (N_9961,N_2876,N_1404);
and U9962 (N_9962,N_4164,N_148);
and U9963 (N_9963,N_4091,N_3559);
and U9964 (N_9964,N_3218,N_689);
and U9965 (N_9965,N_547,N_2109);
or U9966 (N_9966,N_149,N_393);
nor U9967 (N_9967,N_2503,N_4883);
xnor U9968 (N_9968,N_3766,N_1700);
nand U9969 (N_9969,N_4796,N_469);
or U9970 (N_9970,N_3100,N_2158);
nor U9971 (N_9971,N_3506,N_2357);
nand U9972 (N_9972,N_2772,N_241);
nand U9973 (N_9973,N_52,N_3706);
nor U9974 (N_9974,N_510,N_4352);
nor U9975 (N_9975,N_4601,N_490);
nor U9976 (N_9976,N_2865,N_3702);
xnor U9977 (N_9977,N_4838,N_1598);
nor U9978 (N_9978,N_4273,N_2996);
nor U9979 (N_9979,N_1071,N_163);
nand U9980 (N_9980,N_1478,N_209);
nand U9981 (N_9981,N_2277,N_4529);
and U9982 (N_9982,N_2223,N_4269);
xnor U9983 (N_9983,N_2079,N_4104);
or U9984 (N_9984,N_2404,N_3596);
or U9985 (N_9985,N_4531,N_3782);
xor U9986 (N_9986,N_195,N_4281);
nand U9987 (N_9987,N_2712,N_294);
or U9988 (N_9988,N_4910,N_1330);
and U9989 (N_9989,N_3471,N_4085);
xnor U9990 (N_9990,N_708,N_483);
and U9991 (N_9991,N_3912,N_1855);
nand U9992 (N_9992,N_4443,N_3535);
xnor U9993 (N_9993,N_2308,N_3543);
nand U9994 (N_9994,N_4179,N_4039);
and U9995 (N_9995,N_3973,N_1547);
nand U9996 (N_9996,N_2476,N_607);
nand U9997 (N_9997,N_4975,N_4607);
xnor U9998 (N_9998,N_3364,N_3619);
nand U9999 (N_9999,N_2765,N_2376);
nor U10000 (N_10000,N_7769,N_5809);
nand U10001 (N_10001,N_8662,N_6428);
xnor U10002 (N_10002,N_7449,N_8930);
or U10003 (N_10003,N_8255,N_7230);
nand U10004 (N_10004,N_7245,N_5953);
or U10005 (N_10005,N_8869,N_9065);
nor U10006 (N_10006,N_5643,N_5424);
or U10007 (N_10007,N_6817,N_6830);
nand U10008 (N_10008,N_9063,N_9184);
xor U10009 (N_10009,N_5281,N_8514);
nand U10010 (N_10010,N_7857,N_6400);
and U10011 (N_10011,N_9246,N_9967);
and U10012 (N_10012,N_9887,N_7674);
xnor U10013 (N_10013,N_5466,N_8069);
xnor U10014 (N_10014,N_5129,N_6944);
nor U10015 (N_10015,N_7711,N_6484);
nor U10016 (N_10016,N_6735,N_9103);
nor U10017 (N_10017,N_9002,N_7429);
or U10018 (N_10018,N_8620,N_9274);
nand U10019 (N_10019,N_7794,N_7334);
and U10020 (N_10020,N_8455,N_5137);
and U10021 (N_10021,N_9347,N_7069);
nand U10022 (N_10022,N_5050,N_6551);
nand U10023 (N_10023,N_7903,N_8827);
nor U10024 (N_10024,N_6713,N_9912);
nor U10025 (N_10025,N_7930,N_5936);
nor U10026 (N_10026,N_9699,N_8442);
and U10027 (N_10027,N_7056,N_6811);
and U10028 (N_10028,N_6905,N_9484);
and U10029 (N_10029,N_8368,N_5387);
and U10030 (N_10030,N_5413,N_7477);
nor U10031 (N_10031,N_7292,N_5013);
xnor U10032 (N_10032,N_7510,N_8879);
xor U10033 (N_10033,N_6542,N_5333);
or U10034 (N_10034,N_9426,N_5390);
and U10035 (N_10035,N_6034,N_5046);
and U10036 (N_10036,N_9676,N_6559);
nor U10037 (N_10037,N_9503,N_5716);
nand U10038 (N_10038,N_9144,N_5527);
or U10039 (N_10039,N_9383,N_9437);
xnor U10040 (N_10040,N_8886,N_9166);
nand U10041 (N_10041,N_8502,N_8062);
and U10042 (N_10042,N_8139,N_8240);
and U10043 (N_10043,N_9129,N_7094);
and U10044 (N_10044,N_7518,N_6437);
nor U10045 (N_10045,N_5010,N_6798);
nand U10046 (N_10046,N_5986,N_9348);
or U10047 (N_10047,N_9499,N_9464);
xnor U10048 (N_10048,N_5200,N_7084);
nand U10049 (N_10049,N_9090,N_8802);
xnor U10050 (N_10050,N_6614,N_5829);
or U10051 (N_10051,N_6216,N_5488);
nor U10052 (N_10052,N_8756,N_8916);
and U10053 (N_10053,N_7490,N_9283);
xnor U10054 (N_10054,N_9584,N_9543);
xor U10055 (N_10055,N_5025,N_5127);
and U10056 (N_10056,N_6083,N_7091);
xor U10057 (N_10057,N_7832,N_8887);
xor U10058 (N_10058,N_6898,N_9877);
and U10059 (N_10059,N_5246,N_5041);
xor U10060 (N_10060,N_5168,N_9577);
or U10061 (N_10061,N_7482,N_9731);
xnor U10062 (N_10062,N_8909,N_5341);
or U10063 (N_10063,N_7238,N_5812);
xor U10064 (N_10064,N_5225,N_5991);
nor U10065 (N_10065,N_5315,N_8675);
nand U10066 (N_10066,N_6116,N_7578);
or U10067 (N_10067,N_8285,N_8454);
xor U10068 (N_10068,N_5566,N_6543);
nand U10069 (N_10069,N_6653,N_7552);
nor U10070 (N_10070,N_8427,N_9972);
nand U10071 (N_10071,N_8633,N_8892);
xor U10072 (N_10072,N_9918,N_9336);
nand U10073 (N_10073,N_7335,N_8969);
xnor U10074 (N_10074,N_6991,N_9329);
xnor U10075 (N_10075,N_9636,N_5144);
or U10076 (N_10076,N_9349,N_5957);
and U10077 (N_10077,N_8720,N_8176);
or U10078 (N_10078,N_9496,N_5051);
and U10079 (N_10079,N_5079,N_7059);
nand U10080 (N_10080,N_6256,N_6609);
nor U10081 (N_10081,N_5021,N_9169);
nand U10082 (N_10082,N_8051,N_8725);
and U10083 (N_10083,N_7534,N_6884);
nor U10084 (N_10084,N_9368,N_5234);
xnor U10085 (N_10085,N_8395,N_8746);
and U10086 (N_10086,N_6536,N_7563);
or U10087 (N_10087,N_9644,N_7648);
or U10088 (N_10088,N_8371,N_7286);
xnor U10089 (N_10089,N_9334,N_5714);
or U10090 (N_10090,N_8966,N_7182);
or U10091 (N_10091,N_5139,N_9792);
xor U10092 (N_10092,N_6629,N_8537);
xor U10093 (N_10093,N_7822,N_7480);
and U10094 (N_10094,N_6397,N_5628);
and U10095 (N_10095,N_7602,N_7263);
nand U10096 (N_10096,N_5211,N_7498);
xor U10097 (N_10097,N_6937,N_9844);
and U10098 (N_10098,N_8790,N_5340);
and U10099 (N_10099,N_5810,N_5295);
or U10100 (N_10100,N_6195,N_9981);
or U10101 (N_10101,N_9305,N_6700);
xor U10102 (N_10102,N_5892,N_7894);
xor U10103 (N_10103,N_8083,N_9658);
nor U10104 (N_10104,N_6917,N_9915);
nor U10105 (N_10105,N_8761,N_8276);
nor U10106 (N_10106,N_5405,N_9740);
and U10107 (N_10107,N_7907,N_6483);
and U10108 (N_10108,N_8902,N_8170);
nor U10109 (N_10109,N_8159,N_6855);
or U10110 (N_10110,N_7651,N_6273);
xnor U10111 (N_10111,N_7496,N_7437);
nand U10112 (N_10112,N_8772,N_8666);
nand U10113 (N_10113,N_5406,N_8302);
xor U10114 (N_10114,N_7675,N_5368);
nor U10115 (N_10115,N_7111,N_6237);
nand U10116 (N_10116,N_8222,N_8940);
xnor U10117 (N_10117,N_6761,N_9038);
xor U10118 (N_10118,N_8534,N_5393);
xor U10119 (N_10119,N_7078,N_8810);
nor U10120 (N_10120,N_7953,N_9082);
or U10121 (N_10121,N_9021,N_5993);
and U10122 (N_10122,N_6411,N_7555);
nor U10123 (N_10123,N_5596,N_7764);
nor U10124 (N_10124,N_7246,N_8536);
or U10125 (N_10125,N_8331,N_6520);
nor U10126 (N_10126,N_6595,N_7910);
nand U10127 (N_10127,N_7573,N_6436);
xnor U10128 (N_10128,N_5784,N_9939);
or U10129 (N_10129,N_5088,N_9277);
nand U10130 (N_10130,N_5223,N_7233);
and U10131 (N_10131,N_7671,N_7195);
nand U10132 (N_10132,N_8858,N_9811);
and U10133 (N_10133,N_9935,N_8861);
nor U10134 (N_10134,N_5448,N_7279);
nor U10135 (N_10135,N_7556,N_8671);
or U10136 (N_10136,N_5635,N_6841);
nor U10137 (N_10137,N_7854,N_7974);
xnor U10138 (N_10138,N_6247,N_5155);
nand U10139 (N_10139,N_8158,N_8438);
and U10140 (N_10140,N_5302,N_7736);
and U10141 (N_10141,N_9363,N_8364);
xnor U10142 (N_10142,N_8608,N_6077);
nor U10143 (N_10143,N_7714,N_9473);
nor U10144 (N_10144,N_5577,N_9052);
xnor U10145 (N_10145,N_9051,N_5715);
xor U10146 (N_10146,N_6205,N_8722);
and U10147 (N_10147,N_6152,N_7349);
nor U10148 (N_10148,N_9493,N_5774);
and U10149 (N_10149,N_6580,N_8961);
nand U10150 (N_10150,N_7739,N_8372);
or U10151 (N_10151,N_8094,N_9855);
nor U10152 (N_10152,N_7402,N_8496);
nand U10153 (N_10153,N_9869,N_8248);
nand U10154 (N_10154,N_8263,N_8360);
or U10155 (N_10155,N_7244,N_6788);
xnor U10156 (N_10156,N_7257,N_9903);
or U10157 (N_10157,N_8140,N_7462);
nand U10158 (N_10158,N_8901,N_8224);
and U10159 (N_10159,N_7696,N_5650);
or U10160 (N_10160,N_8737,N_6210);
or U10161 (N_10161,N_8813,N_5181);
and U10162 (N_10162,N_8125,N_6674);
nor U10163 (N_10163,N_9888,N_5251);
nor U10164 (N_10164,N_5286,N_9727);
nor U10165 (N_10165,N_8845,N_6581);
or U10166 (N_10166,N_6959,N_5889);
and U10167 (N_10167,N_7049,N_5349);
xnor U10168 (N_10168,N_5569,N_8112);
xor U10169 (N_10169,N_5588,N_6045);
and U10170 (N_10170,N_7283,N_7274);
and U10171 (N_10171,N_7684,N_9088);
nand U10172 (N_10172,N_8218,N_9562);
nor U10173 (N_10173,N_5170,N_7422);
and U10174 (N_10174,N_8279,N_9900);
or U10175 (N_10175,N_7299,N_5813);
xnor U10176 (N_10176,N_7366,N_9551);
xor U10177 (N_10177,N_9718,N_9535);
or U10178 (N_10178,N_6987,N_6507);
or U10179 (N_10179,N_8403,N_6321);
and U10180 (N_10180,N_5480,N_5749);
and U10181 (N_10181,N_6492,N_6856);
nand U10182 (N_10182,N_7616,N_5007);
nor U10183 (N_10183,N_6862,N_9949);
nand U10184 (N_10184,N_9863,N_6327);
nand U10185 (N_10185,N_5497,N_5854);
or U10186 (N_10186,N_8997,N_9695);
or U10187 (N_10187,N_9650,N_5922);
xnor U10188 (N_10188,N_7594,N_6197);
or U10189 (N_10189,N_6339,N_6166);
xnor U10190 (N_10190,N_6225,N_5262);
and U10191 (N_10191,N_9081,N_5012);
xor U10192 (N_10192,N_9100,N_7989);
or U10193 (N_10193,N_8038,N_5549);
nand U10194 (N_10194,N_8043,N_9353);
nand U10195 (N_10195,N_8503,N_5827);
and U10196 (N_10196,N_7317,N_8658);
nand U10197 (N_10197,N_7083,N_6505);
nor U10198 (N_10198,N_6930,N_7791);
xnor U10199 (N_10199,N_5180,N_9569);
and U10200 (N_10200,N_6943,N_9954);
nand U10201 (N_10201,N_7087,N_7810);
nor U10202 (N_10202,N_9269,N_9756);
or U10203 (N_10203,N_7288,N_5726);
and U10204 (N_10204,N_9064,N_9250);
or U10205 (N_10205,N_7300,N_5456);
xnor U10206 (N_10206,N_5027,N_9494);
nand U10207 (N_10207,N_9848,N_9640);
or U10208 (N_10208,N_6230,N_8924);
and U10209 (N_10209,N_7312,N_8651);
or U10210 (N_10210,N_5967,N_6669);
nand U10211 (N_10211,N_5968,N_5376);
or U10212 (N_10212,N_6773,N_9627);
xnor U10213 (N_10213,N_5469,N_6717);
and U10214 (N_10214,N_6560,N_8749);
nor U10215 (N_10215,N_5781,N_9549);
nand U10216 (N_10216,N_7881,N_6528);
nor U10217 (N_10217,N_5288,N_5342);
and U10218 (N_10218,N_5339,N_8053);
and U10219 (N_10219,N_8102,N_6851);
xnor U10220 (N_10220,N_8303,N_8617);
xnor U10221 (N_10221,N_8817,N_6600);
nor U10222 (N_10222,N_6740,N_6885);
and U10223 (N_10223,N_6092,N_6497);
nor U10224 (N_10224,N_7136,N_6940);
nand U10225 (N_10225,N_5943,N_9476);
and U10226 (N_10226,N_5990,N_9053);
nor U10227 (N_10227,N_7662,N_8831);
xnor U10228 (N_10228,N_6963,N_9587);
xnor U10229 (N_10229,N_9456,N_9730);
nand U10230 (N_10230,N_5183,N_8079);
xor U10231 (N_10231,N_8359,N_9254);
nand U10232 (N_10232,N_8922,N_7319);
nand U10233 (N_10233,N_9242,N_8153);
xor U10234 (N_10234,N_7050,N_9001);
and U10235 (N_10235,N_5189,N_6202);
nor U10236 (N_10236,N_9359,N_5780);
and U10237 (N_10237,N_7514,N_8678);
nor U10238 (N_10238,N_6526,N_9582);
nand U10239 (N_10239,N_9298,N_8167);
and U10240 (N_10240,N_6458,N_7060);
or U10241 (N_10241,N_5850,N_8217);
nand U10242 (N_10242,N_7611,N_5910);
nand U10243 (N_10243,N_5103,N_6553);
nand U10244 (N_10244,N_6519,N_7768);
and U10245 (N_10245,N_9030,N_9106);
and U10246 (N_10246,N_9435,N_5840);
nand U10247 (N_10247,N_9634,N_9501);
xor U10248 (N_10248,N_6596,N_9055);
nor U10249 (N_10249,N_5230,N_5049);
nand U10250 (N_10250,N_6795,N_7887);
nor U10251 (N_10251,N_8311,N_7085);
xor U10252 (N_10252,N_8573,N_7729);
or U10253 (N_10253,N_5503,N_7596);
nand U10254 (N_10254,N_7682,N_6270);
and U10255 (N_10255,N_5517,N_8814);
or U10256 (N_10256,N_6741,N_7499);
nand U10257 (N_10257,N_5553,N_8721);
nor U10258 (N_10258,N_8424,N_5075);
nand U10259 (N_10259,N_6659,N_5821);
or U10260 (N_10260,N_9107,N_6163);
nand U10261 (N_10261,N_7398,N_5842);
or U10262 (N_10262,N_7475,N_8391);
nand U10263 (N_10263,N_9571,N_8650);
and U10264 (N_10264,N_8466,N_8387);
xnor U10265 (N_10265,N_5932,N_8733);
or U10266 (N_10266,N_6957,N_7450);
xor U10267 (N_10267,N_9137,N_7090);
nor U10268 (N_10268,N_7034,N_8266);
or U10269 (N_10269,N_9952,N_7329);
xnor U10270 (N_10270,N_8705,N_5818);
xor U10271 (N_10271,N_8127,N_8314);
nor U10272 (N_10272,N_9333,N_5559);
and U10273 (N_10273,N_6575,N_7524);
and U10274 (N_10274,N_6103,N_9238);
and U10275 (N_10275,N_5008,N_9817);
nor U10276 (N_10276,N_8184,N_8398);
nand U10277 (N_10277,N_5598,N_8479);
and U10278 (N_10278,N_7224,N_8273);
or U10279 (N_10279,N_7753,N_7957);
xnor U10280 (N_10280,N_7842,N_5835);
or U10281 (N_10281,N_6141,N_9362);
and U10282 (N_10282,N_9157,N_9414);
nand U10283 (N_10283,N_9358,N_8039);
nor U10284 (N_10284,N_9071,N_6696);
and U10285 (N_10285,N_7723,N_7618);
and U10286 (N_10286,N_5169,N_8646);
xnor U10287 (N_10287,N_6775,N_5490);
nor U10288 (N_10288,N_6387,N_8807);
and U10289 (N_10289,N_8407,N_6467);
nand U10290 (N_10290,N_5601,N_9560);
or U10291 (N_10291,N_9762,N_7567);
or U10292 (N_10292,N_6755,N_8553);
xor U10293 (N_10293,N_6405,N_6768);
nand U10294 (N_10294,N_5004,N_7442);
and U10295 (N_10295,N_5475,N_8147);
nand U10296 (N_10296,N_9694,N_6335);
nor U10297 (N_10297,N_7793,N_9755);
nor U10298 (N_10298,N_9592,N_6843);
and U10299 (N_10299,N_6514,N_9774);
nand U10300 (N_10300,N_5580,N_9315);
nand U10301 (N_10301,N_7859,N_6683);
and U10302 (N_10302,N_7620,N_5348);
and U10303 (N_10303,N_8082,N_7527);
nor U10304 (N_10304,N_5055,N_6232);
nor U10305 (N_10305,N_6810,N_7585);
xor U10306 (N_10306,N_6971,N_7321);
xor U10307 (N_10307,N_6353,N_8459);
nand U10308 (N_10308,N_5114,N_8647);
nor U10309 (N_10309,N_9712,N_5930);
nor U10310 (N_10310,N_7964,N_7874);
nand U10311 (N_10311,N_5542,N_5186);
nor U10312 (N_10312,N_9508,N_7021);
or U10313 (N_10313,N_5844,N_5064);
xnor U10314 (N_10314,N_7763,N_8097);
xor U10315 (N_10315,N_9264,N_5972);
xor U10316 (N_10316,N_7837,N_9294);
nand U10317 (N_10317,N_6350,N_5603);
or U10318 (N_10318,N_7659,N_8264);
xnor U10319 (N_10319,N_7472,N_6178);
nand U10320 (N_10320,N_8088,N_8340);
and U10321 (N_10321,N_8137,N_6376);
nand U10322 (N_10322,N_6089,N_8771);
nor U10323 (N_10323,N_8815,N_6969);
xor U10324 (N_10324,N_7082,N_9003);
xor U10325 (N_10325,N_8483,N_8660);
nand U10326 (N_10326,N_9777,N_5963);
or U10327 (N_10327,N_6236,N_5401);
or U10328 (N_10328,N_5353,N_5575);
and U10329 (N_10329,N_6510,N_7403);
xor U10330 (N_10330,N_6509,N_6714);
or U10331 (N_10331,N_9374,N_5274);
or U10332 (N_10332,N_8577,N_6607);
or U10333 (N_10333,N_8609,N_6567);
and U10334 (N_10334,N_9345,N_9632);
and U10335 (N_10335,N_8192,N_8524);
or U10336 (N_10336,N_8832,N_9432);
nor U10337 (N_10337,N_6794,N_9164);
nand U10338 (N_10338,N_9706,N_9173);
nor U10339 (N_10339,N_7470,N_8563);
nor U10340 (N_10340,N_6299,N_5875);
or U10341 (N_10341,N_7013,N_5450);
or U10342 (N_10342,N_6495,N_9791);
nor U10343 (N_10343,N_7064,N_6086);
xnor U10344 (N_10344,N_6782,N_8766);
xnor U10345 (N_10345,N_7562,N_7841);
nand U10346 (N_10346,N_6970,N_6455);
nor U10347 (N_10347,N_5940,N_5950);
nand U10348 (N_10348,N_6468,N_8952);
xnor U10349 (N_10349,N_9075,N_5748);
nand U10350 (N_10350,N_6379,N_9602);
xor U10351 (N_10351,N_8580,N_7588);
nor U10352 (N_10352,N_8282,N_6874);
nor U10353 (N_10353,N_8745,N_7077);
xnor U10354 (N_10354,N_7479,N_7191);
and U10355 (N_10355,N_8358,N_6573);
xor U10356 (N_10356,N_7173,N_9293);
nor U10357 (N_10357,N_9225,N_5113);
or U10358 (N_10358,N_9297,N_8541);
xor U10359 (N_10359,N_6274,N_6785);
or U10360 (N_10360,N_5623,N_5671);
xnor U10361 (N_10361,N_5941,N_9880);
and U10362 (N_10362,N_5023,N_5193);
nand U10363 (N_10363,N_8863,N_5266);
nor U10364 (N_10364,N_7044,N_7550);
nand U10365 (N_10365,N_7447,N_7985);
or U10366 (N_10366,N_6887,N_7650);
nor U10367 (N_10367,N_8474,N_9319);
nand U10368 (N_10368,N_8588,N_5960);
nor U10369 (N_10369,N_9971,N_9621);
or U10370 (N_10370,N_7625,N_9529);
or U10371 (N_10371,N_8382,N_5664);
nor U10372 (N_10372,N_5746,N_6754);
nor U10373 (N_10373,N_5526,N_5319);
and U10374 (N_10374,N_5775,N_7967);
and U10375 (N_10375,N_7253,N_6287);
nand U10376 (N_10376,N_9341,N_8181);
nand U10377 (N_10377,N_9603,N_9911);
nor U10378 (N_10378,N_6946,N_5773);
and U10379 (N_10379,N_8385,N_9457);
nor U10380 (N_10380,N_9470,N_9490);
nor U10381 (N_10381,N_6876,N_6984);
xor U10382 (N_10382,N_5111,N_9400);
nor U10383 (N_10383,N_6144,N_6921);
nor U10384 (N_10384,N_6283,N_6312);
or U10385 (N_10385,N_5045,N_9876);
nor U10386 (N_10386,N_6017,N_6477);
nand U10387 (N_10387,N_6566,N_8974);
or U10388 (N_10388,N_7008,N_9896);
or U10389 (N_10389,N_5839,N_9946);
nand U10390 (N_10390,N_9940,N_6470);
xnor U10391 (N_10391,N_9851,N_6814);
or U10392 (N_10392,N_7733,N_9502);
or U10393 (N_10393,N_9633,N_9486);
or U10394 (N_10394,N_7661,N_7564);
nor U10395 (N_10395,N_8219,N_6544);
xor U10396 (N_10396,N_7853,N_8175);
nand U10397 (N_10397,N_6156,N_7901);
or U10398 (N_10398,N_6114,N_5529);
or U10399 (N_10399,N_8014,N_5060);
nor U10400 (N_10400,N_5188,N_9488);
xor U10401 (N_10401,N_7189,N_7131);
and U10402 (N_10402,N_5481,N_8927);
or U10403 (N_10403,N_8226,N_5192);
nand U10404 (N_10404,N_9957,N_5639);
or U10405 (N_10405,N_7344,N_9881);
or U10406 (N_10406,N_9084,N_9096);
xor U10407 (N_10407,N_8730,N_6125);
nor U10408 (N_10408,N_9380,N_7958);
xnor U10409 (N_10409,N_7395,N_6488);
xnor U10410 (N_10410,N_7710,N_6222);
xnor U10411 (N_10411,N_7055,N_5567);
or U10412 (N_10412,N_5620,N_8999);
xnor U10413 (N_10413,N_7147,N_6252);
xor U10414 (N_10414,N_6562,N_9203);
nand U10415 (N_10415,N_8995,N_5868);
xnor U10416 (N_10416,N_6968,N_6266);
xnor U10417 (N_10417,N_8769,N_7115);
xor U10418 (N_10418,N_8185,N_9990);
xnor U10419 (N_10419,N_6693,N_7241);
nand U10420 (N_10420,N_9759,N_5116);
nand U10421 (N_10421,N_8934,N_9482);
nor U10422 (N_10422,N_7818,N_9691);
and U10423 (N_10423,N_8001,N_6952);
xor U10424 (N_10424,N_7549,N_6039);
nor U10425 (N_10425,N_8971,N_6842);
or U10426 (N_10426,N_6618,N_8275);
nor U10427 (N_10427,N_5110,N_9258);
nand U10428 (N_10428,N_7201,N_6981);
and U10429 (N_10429,N_9642,N_5328);
and U10430 (N_10430,N_6269,N_5356);
nor U10431 (N_10431,N_7000,N_9121);
and U10432 (N_10432,N_6155,N_5420);
and U10433 (N_10433,N_8623,N_8031);
and U10434 (N_10434,N_6158,N_7608);
nor U10435 (N_10435,N_6336,N_5062);
nor U10436 (N_10436,N_7266,N_5792);
and U10437 (N_10437,N_5999,N_7963);
and U10438 (N_10438,N_9651,N_7797);
or U10439 (N_10439,N_5325,N_5727);
nand U10440 (N_10440,N_6464,N_9689);
nor U10441 (N_10441,N_5730,N_6199);
nand U10442 (N_10442,N_7929,N_7852);
or U10443 (N_10443,N_7346,N_5306);
nor U10444 (N_10444,N_5425,N_7051);
nor U10445 (N_10445,N_9748,N_9149);
nor U10446 (N_10446,N_9641,N_9239);
xnor U10447 (N_10447,N_7574,N_9853);
or U10448 (N_10448,N_7599,N_8200);
and U10449 (N_10449,N_5956,N_7681);
and U10450 (N_10450,N_8527,N_9520);
and U10451 (N_10451,N_5179,N_5618);
xor U10452 (N_10452,N_8659,N_6028);
xor U10453 (N_10453,N_5757,N_6005);
nand U10454 (N_10454,N_9776,N_5300);
nand U10455 (N_10455,N_6190,N_5296);
xor U10456 (N_10456,N_5962,N_9110);
or U10457 (N_10457,N_8124,N_9454);
nand U10458 (N_10458,N_8050,N_5787);
xnor U10459 (N_10459,N_5489,N_9466);
nor U10460 (N_10460,N_9802,N_7664);
nand U10461 (N_10461,N_9237,N_9767);
nand U10462 (N_10462,N_6844,N_7481);
and U10463 (N_10463,N_9816,N_5560);
xnor U10464 (N_10464,N_9145,N_8690);
or U10465 (N_10465,N_5059,N_7746);
nand U10466 (N_10466,N_9089,N_7047);
nand U10467 (N_10467,N_9404,N_8341);
xor U10468 (N_10468,N_5440,N_9991);
or U10469 (N_10469,N_8067,N_8674);
or U10470 (N_10470,N_6621,N_8028);
and U10471 (N_10471,N_8595,N_5283);
and U10472 (N_10472,N_7787,N_6018);
nor U10473 (N_10473,N_9840,N_7775);
or U10474 (N_10474,N_9527,N_9317);
and U10475 (N_10475,N_5675,N_6719);
and U10476 (N_10476,N_8880,N_9492);
nor U10477 (N_10477,N_5254,N_5697);
xor U10478 (N_10478,N_5166,N_8173);
or U10479 (N_10479,N_6238,N_7502);
nand U10480 (N_10480,N_6284,N_9010);
xnor U10481 (N_10481,N_5444,N_6623);
xor U10482 (N_10482,N_9323,N_7235);
nand U10483 (N_10483,N_6245,N_9530);
or U10484 (N_10484,N_9583,N_5092);
nor U10485 (N_10485,N_6722,N_6352);
and U10486 (N_10486,N_8792,N_8419);
nor U10487 (N_10487,N_8768,N_7698);
nand U10488 (N_10488,N_5754,N_5446);
and U10489 (N_10489,N_5629,N_5001);
xnor U10490 (N_10490,N_7871,N_8521);
and U10491 (N_10491,N_6332,N_8325);
xnor U10492 (N_10492,N_8317,N_9878);
nor U10493 (N_10493,N_5142,N_7328);
xor U10494 (N_10494,N_5634,N_6863);
nand U10495 (N_10495,N_8783,N_5885);
and U10496 (N_10496,N_7135,N_7298);
nor U10497 (N_10497,N_9673,N_8431);
or U10498 (N_10498,N_5708,N_9916);
nand U10499 (N_10499,N_9872,N_9847);
nand U10500 (N_10500,N_7215,N_6800);
xor U10501 (N_10501,N_6820,N_5633);
xnor U10502 (N_10502,N_9284,N_5701);
xor U10503 (N_10503,N_5135,N_6302);
or U10504 (N_10504,N_9407,N_7913);
nor U10505 (N_10505,N_6165,N_8708);
or U10506 (N_10506,N_6254,N_6777);
and U10507 (N_10507,N_6478,N_5778);
or U10508 (N_10508,N_6167,N_9652);
nor U10509 (N_10509,N_5574,N_8236);
nor U10510 (N_10510,N_7965,N_7583);
and U10511 (N_10511,N_5033,N_9648);
nand U10512 (N_10512,N_7258,N_9472);
and U10513 (N_10513,N_9643,N_8828);
and U10514 (N_10514,N_6774,N_6698);
nand U10515 (N_10515,N_6311,N_6857);
xor U10516 (N_10516,N_7046,N_8283);
nand U10517 (N_10517,N_8294,N_6320);
nor U10518 (N_10518,N_8315,N_8357);
xor U10519 (N_10519,N_5790,N_5253);
nor U10520 (N_10520,N_5445,N_6110);
nor U10521 (N_10521,N_7706,N_9536);
nor U10522 (N_10522,N_6701,N_5298);
xor U10523 (N_10523,N_6260,N_8444);
nor U10524 (N_10524,N_8374,N_6825);
or U10525 (N_10525,N_8602,N_5750);
nor U10526 (N_10526,N_9423,N_7336);
nand U10527 (N_10527,N_6385,N_8247);
or U10528 (N_10528,N_9890,N_8008);
and U10529 (N_10529,N_8838,N_5160);
nand U10530 (N_10530,N_9000,N_6682);
or U10531 (N_10531,N_6511,N_5370);
or U10532 (N_10532,N_5533,N_5530);
xnor U10533 (N_10533,N_9188,N_7914);
or U10534 (N_10534,N_9119,N_7700);
nor U10535 (N_10535,N_9728,N_5120);
nor U10536 (N_10536,N_7971,N_9028);
or U10537 (N_10537,N_8132,N_8090);
nor U10538 (N_10538,N_8904,N_7081);
or U10539 (N_10539,N_8187,N_5418);
nand U10540 (N_10540,N_7998,N_7935);
and U10541 (N_10541,N_9963,N_5824);
xnor U10542 (N_10542,N_8943,N_6752);
and U10543 (N_10543,N_8443,N_8686);
and U10544 (N_10544,N_7032,N_7105);
or U10545 (N_10545,N_6890,N_8033);
nor U10546 (N_10546,N_6160,N_9248);
and U10547 (N_10547,N_5699,N_6815);
nand U10548 (N_10548,N_9376,N_5037);
nor U10549 (N_10549,N_9961,N_6404);
xnor U10550 (N_10550,N_6715,N_5357);
nand U10551 (N_10551,N_6627,N_9760);
or U10552 (N_10552,N_9240,N_8253);
and U10553 (N_10553,N_8923,N_7001);
and U10554 (N_10554,N_8500,N_7384);
and U10555 (N_10555,N_8926,N_9161);
and U10556 (N_10556,N_6218,N_6063);
nand U10557 (N_10557,N_9754,N_7825);
nand U10558 (N_10558,N_5121,N_5858);
xnor U10559 (N_10559,N_8677,N_9210);
and U10560 (N_10560,N_8267,N_7738);
and U10561 (N_10561,N_7351,N_5165);
and U10562 (N_10562,N_9775,N_5378);
and U10563 (N_10563,N_5082,N_8918);
or U10564 (N_10564,N_6911,N_8672);
nor U10565 (N_10565,N_5908,N_7007);
nor U10566 (N_10566,N_9440,N_5516);
nor U10567 (N_10567,N_8401,N_5038);
and U10568 (N_10568,N_5721,N_5873);
nand U10569 (N_10569,N_6134,N_8826);
and U10570 (N_10570,N_6781,N_7396);
or U10571 (N_10571,N_8973,N_5496);
and U10572 (N_10572,N_7080,N_8960);
or U10573 (N_10573,N_9076,N_9937);
nor U10574 (N_10574,N_8329,N_5670);
or U10575 (N_10575,N_6891,N_6101);
nand U10576 (N_10576,N_8522,N_7024);
xor U10577 (N_10577,N_8323,N_9458);
or U10578 (N_10578,N_5294,N_6564);
nor U10579 (N_10579,N_5646,N_5336);
or U10580 (N_10580,N_7656,N_9593);
nor U10581 (N_10581,N_5720,N_9524);
xor U10582 (N_10582,N_7058,N_9279);
or U10583 (N_10583,N_8320,N_6318);
or U10584 (N_10584,N_5913,N_8959);
or U10585 (N_10585,N_9975,N_5769);
nor U10586 (N_10586,N_8316,N_8074);
and U10587 (N_10587,N_5649,N_5866);
nand U10588 (N_10588,N_6624,N_8687);
nor U10589 (N_10589,N_6903,N_7461);
xor U10590 (N_10590,N_5545,N_5191);
xnor U10591 (N_10591,N_8936,N_5355);
and U10592 (N_10592,N_6291,N_5066);
xnor U10593 (N_10593,N_9183,N_9958);
nor U10594 (N_10594,N_5995,N_7086);
xnor U10595 (N_10595,N_9309,N_6915);
nor U10596 (N_10596,N_9864,N_9693);
or U10597 (N_10597,N_5236,N_5346);
nor U10598 (N_10598,N_6285,N_6657);
nor U10599 (N_10599,N_8489,N_8414);
xnor U10600 (N_10600,N_7119,N_5026);
or U10601 (N_10601,N_5123,N_9057);
xor U10602 (N_10602,N_5942,N_5557);
nor U10603 (N_10603,N_6871,N_6384);
nand U10604 (N_10604,N_8873,N_5162);
xor U10605 (N_10605,N_6177,N_6792);
or U10606 (N_10606,N_8797,N_6220);
or U10607 (N_10607,N_9385,N_7673);
nor U10608 (N_10608,N_9011,N_8697);
and U10609 (N_10609,N_6646,N_6852);
nor U10610 (N_10610,N_9459,N_7864);
or U10611 (N_10611,N_9966,N_5725);
and U10612 (N_10612,N_6742,N_8152);
xnor U10613 (N_10613,N_5916,N_6334);
nor U10614 (N_10614,N_6496,N_9998);
nor U10615 (N_10615,N_7375,N_8344);
xnor U10616 (N_10616,N_9992,N_6150);
and U10617 (N_10617,N_5705,N_5194);
xor U10618 (N_10618,N_7506,N_8877);
nand U10619 (N_10619,N_5884,N_9430);
nand U10620 (N_10620,N_5388,N_5586);
xnor U10621 (N_10621,N_9252,N_8844);
nor U10622 (N_10622,N_7634,N_7928);
and U10623 (N_10623,N_8699,N_9780);
nand U10624 (N_10624,N_9697,N_5073);
xor U10625 (N_10625,N_9153,N_5964);
xor U10626 (N_10626,N_8946,N_9101);
nand U10627 (N_10627,N_5642,N_8568);
xor U10628 (N_10628,N_7848,N_8113);
xnor U10629 (N_10629,N_5287,N_5918);
nor U10630 (N_10630,N_7315,N_5126);
xor U10631 (N_10631,N_7483,N_5805);
or U10632 (N_10632,N_9793,N_5693);
xnor U10633 (N_10633,N_9513,N_5602);
xnor U10634 (N_10634,N_8293,N_5978);
nand U10635 (N_10635,N_7424,N_6571);
nand U10636 (N_10636,N_7548,N_8951);
nor U10637 (N_10637,N_7211,N_8469);
nor U10638 (N_10638,N_8723,N_8308);
or U10639 (N_10639,N_5293,N_6136);
nor U10640 (N_10640,N_6490,N_7271);
xor U10641 (N_10641,N_5044,N_5119);
or U10642 (N_10642,N_8509,N_6226);
nor U10643 (N_10643,N_8476,N_6329);
and U10644 (N_10644,N_7504,N_9127);
nand U10645 (N_10645,N_5091,N_6130);
nor U10646 (N_10646,N_6960,N_8481);
nand U10647 (N_10647,N_8242,N_8468);
nor U10648 (N_10648,N_5927,N_9698);
nand U10649 (N_10649,N_8432,N_9312);
or U10650 (N_10650,N_9046,N_6389);
nand U10651 (N_10651,N_8421,N_6985);
and U10652 (N_10652,N_8882,N_6709);
nand U10653 (N_10653,N_7460,N_7207);
nor U10654 (N_10654,N_6296,N_5779);
nand U10655 (N_10655,N_9512,N_7560);
or U10656 (N_10656,N_9735,N_5572);
or U10657 (N_10657,N_6322,N_9953);
or U10658 (N_10658,N_5439,N_7603);
and U10659 (N_10659,N_9865,N_8780);
nor U10660 (N_10660,N_7613,N_6622);
nor U10661 (N_10661,N_6860,N_9226);
xor U10662 (N_10662,N_5305,N_6516);
xor U10663 (N_10663,N_5143,N_5925);
and U10664 (N_10664,N_9843,N_8446);
xnor U10665 (N_10665,N_8406,N_7255);
nor U10666 (N_10666,N_7692,N_6821);
nor U10667 (N_10667,N_9744,N_7751);
and U10668 (N_10668,N_7401,N_9232);
or U10669 (N_10669,N_7256,N_6524);
and U10670 (N_10670,N_8994,N_9007);
nand U10671 (N_10671,N_7325,N_5463);
xnor U10672 (N_10672,N_8622,N_8229);
nor U10673 (N_10673,N_8913,N_7902);
or U10674 (N_10674,N_7219,N_8865);
xnor U10675 (N_10675,N_6605,N_5024);
and U10676 (N_10676,N_7765,N_8231);
nand U10677 (N_10677,N_6235,N_5876);
nor U10678 (N_10678,N_8355,N_6889);
xnor U10679 (N_10679,N_8691,N_6042);
nand U10680 (N_10680,N_6878,N_5961);
or U10681 (N_10681,N_5825,N_6325);
or U10682 (N_10682,N_8155,N_7925);
and U10683 (N_10683,N_5719,N_6660);
and U10684 (N_10684,N_5455,N_5381);
or U10685 (N_10685,N_8441,N_9628);
or U10686 (N_10686,N_9061,N_8767);
nor U10687 (N_10687,N_8517,N_8840);
and U10688 (N_10688,N_9684,N_6349);
and U10689 (N_10689,N_8533,N_7730);
nor U10690 (N_10690,N_6793,N_9343);
or U10691 (N_10691,N_6359,N_7089);
or U10692 (N_10692,N_9964,N_9316);
xor U10693 (N_10693,N_8084,N_7206);
and U10694 (N_10694,N_5257,N_6574);
nor U10695 (N_10695,N_6179,N_9229);
nor U10696 (N_10696,N_9931,N_7337);
xor U10697 (N_10697,N_6787,N_6050);
nand U10698 (N_10698,N_8763,N_6345);
nor U10699 (N_10699,N_7154,N_6219);
or U10700 (N_10700,N_6839,N_8848);
xor U10701 (N_10701,N_9649,N_7416);
xor U10702 (N_10702,N_7529,N_8162);
nor U10703 (N_10703,N_9540,N_8654);
nor U10704 (N_10704,N_8907,N_7679);
and U10705 (N_10705,N_7517,N_9122);
xnor U10706 (N_10706,N_7847,N_8872);
nor U10707 (N_10707,N_8004,N_7978);
xor U10708 (N_10708,N_5227,N_8296);
and U10709 (N_10709,N_8692,N_9442);
or U10710 (N_10710,N_8569,N_9068);
and U10711 (N_10711,N_8025,N_8804);
or U10712 (N_10712,N_5808,N_7626);
xor U10713 (N_10713,N_6196,N_5722);
or U10714 (N_10714,N_8350,N_9823);
or U10715 (N_10715,N_5157,N_8567);
xnor U10716 (N_10716,N_9436,N_8643);
xor U10717 (N_10717,N_5133,N_7627);
or U10718 (N_10718,N_7485,N_9941);
and U10719 (N_10719,N_7614,N_5703);
nor U10720 (N_10720,N_9328,N_5612);
nor U10721 (N_10721,N_8174,N_7242);
xor U10722 (N_10722,N_5472,N_8965);
or U10723 (N_10723,N_6778,N_6712);
nor U10724 (N_10724,N_9616,N_7306);
and U10725 (N_10725,N_6370,N_9812);
nor U10726 (N_10726,N_6818,N_9711);
nand U10727 (N_10727,N_8758,N_7088);
nor U10728 (N_10728,N_9799,N_7382);
xor U10729 (N_10729,N_7121,N_8682);
nand U10730 (N_10730,N_5652,N_6882);
and U10731 (N_10731,N_6021,N_5627);
nor U10732 (N_10732,N_7017,N_9405);
and U10733 (N_10733,N_5134,N_7523);
nand U10734 (N_10734,N_5043,N_8732);
and U10735 (N_10735,N_5147,N_6161);
nor U10736 (N_10736,N_5926,N_6308);
xor U10737 (N_10737,N_6108,N_7067);
and U10738 (N_10738,N_7511,N_8376);
or U10739 (N_10739,N_7036,N_6973);
or U10740 (N_10740,N_5806,N_8963);
nand U10741 (N_10741,N_5656,N_9017);
and U10742 (N_10742,N_7354,N_5237);
xor U10743 (N_10743,N_6003,N_7497);
nand U10744 (N_10744,N_5905,N_6850);
nor U10745 (N_10745,N_8847,N_8390);
xnor U10746 (N_10746,N_8508,N_9805);
or U10747 (N_10747,N_6087,N_7737);
nor U10748 (N_10748,N_8412,N_9989);
xor U10749 (N_10749,N_6681,N_8549);
nor U10750 (N_10750,N_9599,N_5511);
nand U10751 (N_10751,N_5676,N_8035);
xnor U10752 (N_10752,N_9441,N_9771);
xor U10753 (N_10753,N_6515,N_5581);
nand U10754 (N_10754,N_6934,N_7972);
or U10755 (N_10755,N_9399,N_8520);
xor U10756 (N_10756,N_7026,N_9922);
nand U10757 (N_10757,N_6586,N_9986);
nand U10758 (N_10758,N_8205,N_9810);
xor U10759 (N_10759,N_7165,N_5535);
and U10760 (N_10760,N_8110,N_6294);
nor U10761 (N_10761,N_5637,N_8759);
and U10762 (N_10762,N_5877,N_9970);
or U10763 (N_10763,N_6888,N_6678);
and U10764 (N_10764,N_8061,N_6610);
nand U10765 (N_10765,N_7647,N_7959);
and U10766 (N_10766,N_9555,N_9257);
nor U10767 (N_10767,N_6950,N_5919);
xnor U10768 (N_10768,N_9255,N_9299);
and U10769 (N_10769,N_8193,N_7747);
and U10770 (N_10770,N_6718,N_5462);
and U10771 (N_10771,N_7566,N_9322);
nand U10772 (N_10772,N_6081,N_7757);
or U10773 (N_10773,N_7268,N_6757);
or U10774 (N_10774,N_9686,N_7851);
nand U10775 (N_10775,N_6881,N_9526);
xor U10776 (N_10776,N_5870,N_6859);
xor U10777 (N_10777,N_7466,N_9814);
or U10778 (N_10778,N_5297,N_7421);
and U10779 (N_10779,N_9568,N_9690);
and U10780 (N_10780,N_7582,N_6344);
xor U10781 (N_10781,N_7702,N_8005);
nor U10782 (N_10782,N_6323,N_9033);
xor U10783 (N_10783,N_9703,N_6670);
or U10784 (N_10784,N_5534,N_6651);
and U10785 (N_10785,N_9443,N_6214);
and U10786 (N_10786,N_7033,N_8754);
nor U10787 (N_10787,N_8566,N_9308);
or U10788 (N_10788,N_8049,N_5731);
or U10789 (N_10789,N_9902,N_7559);
nand U10790 (N_10790,N_8397,N_5292);
and U10791 (N_10791,N_7758,N_5329);
xor U10792 (N_10792,N_7889,N_5389);
nand U10793 (N_10793,N_5521,N_8834);
xor U10794 (N_10794,N_6633,N_5175);
nor U10795 (N_10795,N_6868,N_9837);
xnor U10796 (N_10796,N_7113,N_6418);
and U10797 (N_10797,N_5770,N_5924);
or U10798 (N_10798,N_8546,N_5228);
nand U10799 (N_10799,N_8632,N_8777);
xnor U10800 (N_10800,N_9723,N_8223);
or U10801 (N_10801,N_7886,N_6686);
and U10802 (N_10802,N_8189,N_9477);
nand U10803 (N_10803,N_8396,N_6012);
xor U10804 (N_10804,N_8955,N_8141);
xor U10805 (N_10805,N_9854,N_9291);
or U10806 (N_10806,N_5056,N_5138);
and U10807 (N_10807,N_5582,N_8906);
nand U10808 (N_10808,N_5600,N_8178);
xnor U10809 (N_10809,N_7920,N_7308);
or U10810 (N_10810,N_9742,N_8998);
nand U10811 (N_10811,N_8893,N_6918);
or U10812 (N_10812,N_6303,N_9741);
and U10813 (N_10813,N_9196,N_5214);
xor U10814 (N_10814,N_8823,N_9175);
or U10815 (N_10815,N_5931,N_9313);
and U10816 (N_10816,N_6480,N_6013);
xor U10817 (N_10817,N_5984,N_7019);
nor U10818 (N_10818,N_5920,N_8232);
and U10819 (N_10819,N_7152,N_7530);
nor U10820 (N_10820,N_8741,N_8410);
nand U10821 (N_10821,N_7425,N_5226);
and U10822 (N_10822,N_7619,N_5303);
and U10823 (N_10823,N_7441,N_7622);
and U10824 (N_10824,N_8839,N_8701);
xor U10825 (N_10825,N_9700,N_8299);
nand U10826 (N_10826,N_9132,N_6826);
xnor U10827 (N_10827,N_6052,N_8449);
nor U10828 (N_10828,N_7697,N_8346);
or U10829 (N_10829,N_5979,N_8484);
xnor U10830 (N_10830,N_5476,N_5863);
xor U10831 (N_10831,N_5578,N_9516);
or U10832 (N_10832,N_8225,N_6085);
and U10833 (N_10833,N_8362,N_6563);
or U10834 (N_10834,N_8369,N_9367);
or U10835 (N_10835,N_5679,N_6289);
nand U10836 (N_10836,N_9675,N_6807);
xnor U10837 (N_10837,N_8931,N_6043);
nor U10838 (N_10838,N_6685,N_9509);
nand U10839 (N_10839,N_5685,N_9142);
nand U10840 (N_10840,N_7839,N_7637);
nand U10841 (N_10841,N_8875,N_8297);
nand U10842 (N_10842,N_5657,N_9419);
and U10843 (N_10843,N_8237,N_6277);
xnor U10844 (N_10844,N_8183,N_9955);
nand U10845 (N_10845,N_9781,N_5971);
nand U10846 (N_10846,N_8416,N_6955);
nand U10847 (N_10847,N_8268,N_8846);
nor U10848 (N_10848,N_9671,N_5422);
or U10849 (N_10849,N_5912,N_5430);
nand U10850 (N_10850,N_5408,N_5299);
xnor U10851 (N_10851,N_7473,N_7022);
nand U10852 (N_10852,N_6132,N_7932);
nand U10853 (N_10853,N_5969,N_8798);
or U10854 (N_10854,N_9763,N_8289);
xor U10855 (N_10855,N_5800,N_9666);
nand U10856 (N_10856,N_6606,N_9249);
and U10857 (N_10857,N_7660,N_5256);
or U10858 (N_10858,N_6636,N_8430);
nor U10859 (N_10859,N_5289,N_5735);
or U10860 (N_10860,N_5063,N_8386);
nand U10861 (N_10861,N_6549,N_5814);
xor U10862 (N_10862,N_8962,N_5611);
nand U10863 (N_10863,N_6060,N_7813);
nand U10864 (N_10864,N_7800,N_6023);
nor U10865 (N_10865,N_5118,N_6424);
nand U10866 (N_10866,N_9831,N_7565);
nor U10867 (N_10867,N_9406,N_5006);
xor U10868 (N_10868,N_8899,N_8626);
nand U10869 (N_10869,N_8774,N_5592);
xnor U10870 (N_10870,N_7405,N_9795);
nand U10871 (N_10871,N_9984,N_5261);
nor U10872 (N_10872,N_5945,N_8058);
and U10873 (N_10873,N_7748,N_7906);
xnor U10874 (N_10874,N_7703,N_6748);
and U10875 (N_10875,N_5382,N_6875);
nand U10876 (N_10876,N_5832,N_5753);
nor U10877 (N_10877,N_7786,N_5187);
xnor U10878 (N_10878,N_9337,N_5402);
or U10879 (N_10879,N_8668,N_7214);
nor U10880 (N_10880,N_5864,N_6255);
xnor U10881 (N_10881,N_8188,N_5845);
or U10882 (N_10882,N_8119,N_9734);
or U10883 (N_10883,N_5648,N_7685);
nor U10884 (N_10884,N_6095,N_5585);
nor U10885 (N_10885,N_9525,N_6989);
and U10886 (N_10886,N_9152,N_8096);
and U10887 (N_10887,N_7833,N_9136);
or U10888 (N_10888,N_7544,N_5109);
and U10889 (N_10889,N_6002,N_7488);
and U10890 (N_10890,N_8743,N_9709);
or U10891 (N_10891,N_6928,N_8642);
nor U10892 (N_10892,N_8629,N_7689);
nand U10893 (N_10893,N_5512,N_7812);
nand U10894 (N_10894,N_8542,N_5786);
and U10895 (N_10895,N_8042,N_5255);
xnor U10896 (N_10896,N_6751,N_6394);
or U10897 (N_10897,N_9014,N_7609);
xnor U10898 (N_10898,N_9923,N_7924);
or U10899 (N_10899,N_7184,N_5558);
or U10900 (N_10900,N_7893,N_6186);
and U10901 (N_10901,N_8518,N_9914);
or U10902 (N_10902,N_7943,N_6124);
and U10903 (N_10903,N_5732,N_5343);
nor U10904 (N_10904,N_6797,N_7824);
and U10905 (N_10905,N_8244,N_8649);
nand U10906 (N_10906,N_8213,N_6756);
nor U10907 (N_10907,N_9427,N_9455);
xnor U10908 (N_10908,N_5543,N_5252);
nand U10909 (N_10909,N_6479,N_5568);
nand U10910 (N_10910,N_7232,N_5802);
or U10911 (N_10911,N_8980,N_6730);
nand U10912 (N_10912,N_9109,N_8322);
nand U10913 (N_10913,N_7428,N_8007);
nand U10914 (N_10914,N_5531,N_5065);
nor U10915 (N_10915,N_5665,N_6182);
nand U10916 (N_10916,N_7210,N_8335);
and U10917 (N_10917,N_6295,N_9202);
nor U10918 (N_10918,N_7997,N_5163);
or U10919 (N_10919,N_7476,N_8448);
and U10920 (N_10920,N_7939,N_9043);
xnor U10921 (N_10921,N_5607,N_6962);
xnor U10922 (N_10922,N_7216,N_6547);
nand U10923 (N_10923,N_9985,N_7640);
nand U10924 (N_10924,N_5599,N_9408);
or U10925 (N_10925,N_8808,N_5794);
nor U10926 (N_10926,N_6708,N_7125);
and U10927 (N_10927,N_5374,N_7052);
or U10928 (N_10928,N_7468,N_8197);
or U10929 (N_10929,N_6395,N_8683);
nor U10930 (N_10930,N_9830,N_9669);
nand U10931 (N_10931,N_9114,N_8439);
and U10932 (N_10932,N_8286,N_7223);
nand U10933 (N_10933,N_9600,N_7572);
xor U10934 (N_10934,N_9092,N_9223);
xnor U10935 (N_10935,N_9702,N_9511);
nor U10936 (N_10936,N_7705,N_5323);
nand U10937 (N_10937,N_9772,N_5752);
nor U10938 (N_10938,N_6961,N_9828);
or U10939 (N_10939,N_5217,N_7187);
nor U10940 (N_10940,N_5921,N_6427);
nand U10941 (N_10941,N_7172,N_6634);
or U10942 (N_10942,N_7116,N_5843);
or U10943 (N_10943,N_6530,N_8238);
xnor U10944 (N_10944,N_5443,N_9211);
and U10945 (N_10945,N_9314,N_6153);
nand U10946 (N_10946,N_6175,N_5606);
and U10947 (N_10947,N_9008,N_7140);
nand U10948 (N_10948,N_7386,N_6425);
nand U10949 (N_10949,N_6442,N_5167);
or U10950 (N_10950,N_5974,N_8306);
or U10951 (N_10951,N_7879,N_6923);
xor U10952 (N_10952,N_6789,N_8993);
nand U10953 (N_10953,N_9838,N_8133);
nand U10954 (N_10954,N_7861,N_5487);
or U10955 (N_10955,N_9517,N_5617);
and U10956 (N_10956,N_5077,N_7071);
xnor U10957 (N_10957,N_5819,N_6974);
and U10958 (N_10958,N_8291,N_7296);
or U10959 (N_10959,N_9751,N_8435);
and U10960 (N_10960,N_6664,N_9667);
or U10961 (N_10961,N_7761,N_7717);
and U10962 (N_10962,N_7944,N_6729);
or U10963 (N_10963,N_8281,N_7708);
nor U10964 (N_10964,N_9126,N_6486);
or U10965 (N_10965,N_9969,N_7727);
or U10966 (N_10966,N_5247,N_8819);
or U10967 (N_10967,N_5002,N_9335);
and U10968 (N_10968,N_8154,N_7387);
xor U10969 (N_10969,N_7843,N_9639);
and U10970 (N_10970,N_6615,N_5717);
nor U10971 (N_10971,N_8859,N_9532);
and U10972 (N_10972,N_5479,N_8560);
and U10973 (N_10973,N_9234,N_6084);
nor U10974 (N_10974,N_7672,N_6743);
xor U10975 (N_10975,N_6500,N_5396);
or U10976 (N_10976,N_9024,N_6958);
nor U10977 (N_10977,N_8064,N_6286);
and U10978 (N_10978,N_6119,N_8348);
and U10979 (N_10979,N_9475,N_8679);
nand U10980 (N_10980,N_8203,N_8099);
xor U10981 (N_10981,N_8172,N_5125);
xor U10982 (N_10982,N_9959,N_5684);
or U10983 (N_10983,N_7979,N_5958);
nand U10984 (N_10984,N_7341,N_8160);
nor U10985 (N_10985,N_8929,N_9162);
or U10986 (N_10986,N_6272,N_5667);
nor U10987 (N_10987,N_8572,N_5148);
or U10988 (N_10988,N_6587,N_6187);
nor U10989 (N_10989,N_8715,N_6319);
and U10990 (N_10990,N_8556,N_9999);
nand U10991 (N_10991,N_7303,N_6176);
nor U10992 (N_10992,N_6173,N_9789);
nand U10993 (N_10993,N_5783,N_7217);
nor U10994 (N_10994,N_8399,N_5367);
nand U10995 (N_10995,N_6009,N_7988);
or U10996 (N_10996,N_7863,N_9072);
xor U10997 (N_10997,N_6126,N_7029);
xnor U10998 (N_10998,N_9227,N_5804);
xnor U10999 (N_10999,N_6517,N_7505);
nand U11000 (N_11000,N_8227,N_6038);
xnor U11001 (N_11001,N_9386,N_5208);
and U11002 (N_11002,N_8949,N_7635);
and U11003 (N_11003,N_9429,N_9994);
and U11004 (N_11004,N_7836,N_8779);
nor U11005 (N_11005,N_5360,N_9893);
nand U11006 (N_11006,N_9968,N_8107);
nor U11007 (N_11007,N_8148,N_5403);
or U11008 (N_11008,N_9561,N_7539);
nor U11009 (N_11009,N_7474,N_6240);
or U11010 (N_11010,N_8040,N_7333);
xor U11011 (N_11011,N_6603,N_6423);
nor U11012 (N_11012,N_6552,N_7691);
and U11013 (N_11013,N_7267,N_8128);
nand U11014 (N_11014,N_9190,N_6749);
nand U11015 (N_11015,N_6877,N_5763);
nor U11016 (N_11016,N_5171,N_9646);
or U11017 (N_11017,N_7073,N_7667);
xor U11018 (N_11018,N_9265,N_8078);
xnor U11019 (N_11019,N_7551,N_8451);
or U11020 (N_11020,N_9006,N_8933);
and U11021 (N_11021,N_6011,N_5154);
nand U11022 (N_11022,N_5740,N_5564);
nand U11023 (N_11023,N_8809,N_8712);
or U11024 (N_11024,N_5394,N_6739);
nor U11025 (N_11025,N_5500,N_5904);
xnor U11026 (N_11026,N_7420,N_7109);
and U11027 (N_11027,N_5996,N_6358);
and U11028 (N_11028,N_8978,N_5326);
and U11029 (N_11029,N_6501,N_5830);
nand U11030 (N_11030,N_7937,N_5218);
nor U11031 (N_11031,N_8343,N_9354);
nand U11032 (N_11032,N_6861,N_9910);
and U11033 (N_11033,N_6941,N_9199);
and U11034 (N_11034,N_9747,N_9463);
xnor U11035 (N_11035,N_5944,N_8408);
xnor U11036 (N_11036,N_5150,N_7446);
xor U11037 (N_11037,N_7668,N_9219);
or U11038 (N_11038,N_8206,N_8757);
nand U11039 (N_11039,N_9733,N_5683);
or U11040 (N_11040,N_5788,N_7663);
and U11041 (N_11041,N_9797,N_6667);
xnor U11042 (N_11042,N_7597,N_5655);
nand U11043 (N_11043,N_9614,N_7631);
nand U11044 (N_11044,N_6804,N_9630);
xnor U11045 (N_11045,N_8136,N_6929);
nand U11046 (N_11046,N_5826,N_9505);
nor U11047 (N_11047,N_9498,N_9987);
or U11048 (N_11048,N_5433,N_8233);
nor U11049 (N_11049,N_9453,N_6532);
nor U11050 (N_11050,N_7642,N_8301);
xor U11051 (N_11051,N_9598,N_7304);
and U11052 (N_11052,N_5363,N_6692);
and U11053 (N_11053,N_6261,N_5071);
nor U11054 (N_11054,N_7670,N_7870);
or U11055 (N_11055,N_9310,N_9588);
or U11056 (N_11056,N_5985,N_9807);
and U11057 (N_11057,N_8867,N_6725);
nand U11058 (N_11058,N_9301,N_7819);
xor U11059 (N_11059,N_7157,N_6976);
or U11060 (N_11060,N_7860,N_8345);
and U11061 (N_11061,N_7970,N_6512);
nand U11062 (N_11062,N_8612,N_7816);
nor U11063 (N_11063,N_6115,N_8216);
nand U11064 (N_11064,N_7749,N_6630);
and U11065 (N_11065,N_8023,N_7297);
nand U11066 (N_11066,N_8681,N_9491);
nor U11067 (N_11067,N_7122,N_7883);
and U11068 (N_11068,N_9926,N_5700);
or U11069 (N_11069,N_6707,N_8816);
xor U11070 (N_11070,N_7003,N_5759);
or U11071 (N_11071,N_7057,N_7591);
xnor U11072 (N_11072,N_5562,N_6658);
and U11073 (N_11073,N_5681,N_6896);
xnor U11074 (N_11074,N_8585,N_9595);
or U11075 (N_11075,N_6784,N_8259);
or U11076 (N_11076,N_5604,N_9995);
xnor U11077 (N_11077,N_7951,N_5537);
nand U11078 (N_11078,N_7391,N_9874);
nand U11079 (N_11079,N_6020,N_5871);
and U11080 (N_11080,N_5020,N_8535);
nand U11081 (N_11081,N_8793,N_5654);
and U11082 (N_11082,N_5838,N_9894);
nor U11083 (N_11083,N_5085,N_5706);
nand U11084 (N_11084,N_7610,N_6233);
and U11085 (N_11085,N_6513,N_8958);
xnor U11086 (N_11086,N_7720,N_8539);
nand U11087 (N_11087,N_7347,N_9141);
or U11088 (N_11088,N_6297,N_8150);
and U11089 (N_11089,N_8470,N_8689);
or U11090 (N_11090,N_5501,N_9631);
nor U11091 (N_11091,N_8849,N_7365);
nor U11092 (N_11092,N_7276,N_7467);
xnor U11093 (N_11093,N_8710,N_8850);
nor U11094 (N_11094,N_8037,N_8900);
nor U11095 (N_11095,N_6809,N_8639);
or U11096 (N_11096,N_7213,N_7409);
or U11097 (N_11097,N_6687,N_8377);
and U11098 (N_11098,N_5235,N_5036);
nor U11099 (N_11099,N_6188,N_8736);
nand U11100 (N_11100,N_8003,N_5309);
nor U11101 (N_11101,N_8006,N_6309);
nand U11102 (N_11102,N_7407,N_9025);
nor U11103 (N_11103,N_9339,N_8310);
xnor U11104 (N_11104,N_6939,N_6638);
or U11105 (N_11105,N_8778,N_9370);
or U11106 (N_11106,N_6031,N_7803);
nor U11107 (N_11107,N_5005,N_6977);
xnor U11108 (N_11108,N_9044,N_9824);
and U11109 (N_11109,N_6100,N_5178);
nand U11110 (N_11110,N_7792,N_7882);
or U11111 (N_11111,N_7916,N_7742);
or U11112 (N_11112,N_6131,N_8030);
or U11113 (N_11113,N_8252,N_5338);
xor U11114 (N_11114,N_6033,N_9556);
and U11115 (N_11115,N_9668,N_9474);
and U11116 (N_11116,N_5421,N_9221);
and U11117 (N_11117,N_9059,N_6760);
or U11118 (N_11118,N_6001,N_8891);
xnor U11119 (N_11119,N_5856,N_9565);
nand U11120 (N_11120,N_6326,N_9012);
nand U11121 (N_11121,N_6239,N_9942);
or U11122 (N_11122,N_9895,N_8381);
xnor U11123 (N_11123,N_6328,N_8575);
xor U11124 (N_11124,N_5758,N_6184);
nor U11125 (N_11125,N_5264,N_9819);
or U11126 (N_11126,N_9779,N_9947);
nor U11127 (N_11127,N_9715,N_8657);
and U11128 (N_11128,N_8624,N_5039);
nand U11129 (N_11129,N_6275,N_5124);
or U11130 (N_11130,N_5414,N_9875);
xor U11131 (N_11131,N_7414,N_9155);
or U11132 (N_11132,N_5644,N_8009);
xnor U11133 (N_11133,N_6816,N_9327);
or U11134 (N_11134,N_8836,N_7099);
xor U11135 (N_11135,N_9764,N_5687);
nor U11136 (N_11136,N_7796,N_8000);
nor U11137 (N_11137,N_8388,N_5395);
nand U11138 (N_11138,N_8057,N_9332);
nand U11139 (N_11139,N_7278,N_6048);
and U11140 (N_11140,N_8925,N_9753);
xnor U11141 (N_11141,N_7815,N_7075);
or U11142 (N_11142,N_9189,N_7781);
nand U11143 (N_11143,N_6263,N_8365);
or U11144 (N_11144,N_9653,N_7068);
nor U11145 (N_11145,N_7171,N_5158);
and U11146 (N_11146,N_6300,N_5797);
or U11147 (N_11147,N_8676,N_8636);
and U11148 (N_11148,N_5099,N_9548);
xor U11149 (N_11149,N_7507,N_9019);
xnor U11150 (N_11150,N_8165,N_5896);
nand U11151 (N_11151,N_7554,N_9163);
xor U11152 (N_11152,N_6215,N_8478);
nor U11153 (N_11153,N_6460,N_7338);
nand U11154 (N_11154,N_9060,N_9263);
and U11155 (N_11155,N_8447,N_9519);
or U11156 (N_11156,N_9539,N_8948);
nand U11157 (N_11157,N_5053,N_7209);
and U11158 (N_11158,N_9213,N_7732);
or U11159 (N_11159,N_7367,N_6554);
or U11160 (N_11160,N_9719,N_7954);
nand U11161 (N_11161,N_8202,N_9861);
and U11162 (N_11162,N_8304,N_5219);
nor U11163 (N_11163,N_5933,N_7227);
nand U11164 (N_11164,N_6769,N_9095);
nor U11165 (N_11165,N_9187,N_6383);
or U11166 (N_11166,N_8789,N_5207);
nor U11167 (N_11167,N_7418,N_6454);
xor U11168 (N_11168,N_9412,N_6453);
or U11169 (N_11169,N_9611,N_8488);
nor U11170 (N_11170,N_7532,N_6555);
xor U11171 (N_11171,N_5659,N_5893);
xnor U11172 (N_11172,N_7629,N_6066);
or U11173 (N_11173,N_5076,N_5364);
or U11174 (N_11174,N_7869,N_8796);
nand U11175 (N_11175,N_5074,N_7353);
and U11176 (N_11176,N_9150,N_6369);
or U11177 (N_11177,N_6895,N_6594);
nand U11178 (N_11178,N_6090,N_8897);
nor U11179 (N_11179,N_5492,N_7443);
nand U11180 (N_11180,N_7074,N_5841);
and U11181 (N_11181,N_6914,N_7445);
or U11182 (N_11182,N_8246,N_7145);
nand U11183 (N_11183,N_8239,N_7079);
or U11184 (N_11184,N_9567,N_5594);
xor U11185 (N_11185,N_9721,N_6908);
nor U11186 (N_11186,N_7439,N_5250);
nand U11187 (N_11187,N_8947,N_9206);
xor U11188 (N_11188,N_7411,N_7987);
xnor U11189 (N_11189,N_6223,N_8020);
nand U11190 (N_11190,N_5608,N_8941);
or U11191 (N_11191,N_6766,N_7713);
nor U11192 (N_11192,N_8752,N_8312);
nor U11193 (N_11193,N_6440,N_9460);
or U11194 (N_11194,N_9079,N_5316);
or U11195 (N_11195,N_9917,N_5738);
nor U11196 (N_11196,N_7129,N_8460);
xnor U11197 (N_11197,N_7137,N_7575);
xnor U11198 (N_11198,N_5452,N_7712);
xor U11199 (N_11199,N_5107,N_9559);
and U11200 (N_11200,N_9619,N_5240);
and U11201 (N_11201,N_5471,N_7170);
and U11202 (N_11202,N_8032,N_8835);
xor U11203 (N_11203,N_8581,N_7875);
xnor U11204 (N_11204,N_8169,N_5478);
nor U11205 (N_11205,N_9397,N_5546);
and U11206 (N_11206,N_5976,N_6572);
xnor U11207 (N_11207,N_7345,N_7962);
nand U11208 (N_11208,N_6406,N_7669);
or U11209 (N_11209,N_9597,N_5973);
or U11210 (N_11210,N_5795,N_5210);
xnor U11211 (N_11211,N_5159,N_9402);
nor U11212 (N_11212,N_6726,N_5669);
or U11213 (N_11213,N_9036,N_9609);
xor U11214 (N_11214,N_9410,N_6576);
and U11215 (N_11215,N_9821,N_9047);
nor U11216 (N_11216,N_6697,N_7435);
and U11217 (N_11217,N_8313,N_8103);
nor U11218 (N_11218,N_9296,N_6644);
or U11219 (N_11219,N_6372,N_5277);
nand U11220 (N_11220,N_9682,N_8550);
xor U11221 (N_11221,N_5556,N_9424);
nand U11222 (N_11222,N_7940,N_5199);
xor U11223 (N_11223,N_6068,N_8592);
and U11224 (N_11224,N_9231,N_8597);
xnor U11225 (N_11225,N_7273,N_6396);
nand U11226 (N_11226,N_7364,N_7174);
xor U11227 (N_11227,N_6612,N_7831);
xor U11228 (N_11228,N_5391,N_5742);
and U11229 (N_11229,N_9664,N_9198);
and U11230 (N_11230,N_6242,N_5638);
nor U11231 (N_11231,N_5442,N_6410);
xnor U11232 (N_11232,N_9270,N_8652);
nand U11233 (N_11233,N_7827,N_9495);
xnor U11234 (N_11234,N_6978,N_8970);
nand U11235 (N_11235,N_5468,N_6143);
or U11236 (N_11236,N_8467,N_5878);
or U11237 (N_11237,N_6632,N_9041);
or U11238 (N_11238,N_7630,N_9612);
nand U11239 (N_11239,N_5837,N_6584);
nand U11240 (N_11240,N_6313,N_5351);
xnor U11241 (N_11241,N_8548,N_6639);
xnor U11242 (N_11242,N_7830,N_6192);
or U11243 (N_11243,N_8795,N_8932);
nand U11244 (N_11244,N_7128,N_7726);
nand U11245 (N_11245,N_7992,N_9428);
xor U11246 (N_11246,N_5280,N_7724);
xnor U11247 (N_11247,N_9062,N_5573);
or U11248 (N_11248,N_7880,N_8392);
xnor U11249 (N_11249,N_8063,N_7410);
nor U11250 (N_11250,N_5816,N_7324);
nand U11251 (N_11251,N_8254,N_7092);
and U11252 (N_11252,N_6151,N_9085);
or U11253 (N_11253,N_5833,N_7981);
xor U11254 (N_11254,N_8499,N_8885);
nand U11255 (N_11255,N_8221,N_7589);
or U11256 (N_11256,N_5347,N_9138);
xnor U11257 (N_11257,N_5164,N_5270);
nor U11258 (N_11258,N_7666,N_8319);
or U11259 (N_11259,N_5354,N_7540);
xor U11260 (N_11260,N_6067,N_8300);
nor U11261 (N_11261,N_7114,N_7655);
nor U11262 (N_11262,N_8728,N_5377);
nand U11263 (N_11263,N_6228,N_9770);
nand U11264 (N_11264,N_5959,N_6652);
nand U11265 (N_11265,N_5470,N_8111);
nor U11266 (N_11266,N_9905,N_5507);
nor U11267 (N_11267,N_9624,N_6886);
xnor U11268 (N_11268,N_5197,N_5031);
nand U11269 (N_11269,N_5713,N_9286);
nor U11270 (N_11270,N_8166,N_9067);
or U11271 (N_11271,N_9856,N_9845);
nor U11272 (N_11272,N_8822,N_6662);
nor U11273 (N_11273,N_8422,N_9977);
or U11274 (N_11274,N_9176,N_7876);
or U11275 (N_11275,N_8515,N_5828);
nand U11276 (N_11276,N_9659,N_9104);
or U11277 (N_11277,N_8601,N_7043);
and U11278 (N_11278,N_5929,N_8896);
or U11279 (N_11279,N_6805,N_8287);
nor U11280 (N_11280,N_7343,N_7829);
nor U11281 (N_11281,N_6541,N_5040);
nand U11282 (N_11282,N_8305,N_6037);
nand U11283 (N_11283,N_7516,N_6391);
nand U11284 (N_11284,N_6901,N_6986);
xor U11285 (N_11285,N_8404,N_9720);
and U11286 (N_11286,N_8915,N_5086);
nand U11287 (N_11287,N_8803,N_6282);
and U11288 (N_11288,N_7108,N_8791);
nor U11289 (N_11289,N_6439,N_8256);
or U11290 (N_11290,N_7149,N_5184);
nand U11291 (N_11291,N_5042,N_9504);
nand U11292 (N_11292,N_6171,N_5524);
and U11293 (N_11293,N_5886,N_5729);
or U11294 (N_11294,N_7785,N_9444);
nor U11295 (N_11295,N_9461,N_6348);
and U11296 (N_11296,N_7101,N_7359);
nand U11297 (N_11297,N_6316,N_8118);
nand U11298 (N_11298,N_8610,N_8120);
or U11299 (N_11299,N_9818,N_5474);
and U11300 (N_11300,N_8002,N_5030);
or U11301 (N_11301,N_6399,N_6916);
xor U11302 (N_11302,N_9447,N_9832);
nor U11303 (N_11303,N_9207,N_7601);
nand U11304 (N_11304,N_8898,N_7054);
or U11305 (N_11305,N_8409,N_5108);
xor U11306 (N_11306,N_7433,N_5486);
nor U11307 (N_11307,N_8307,N_9425);
or U11308 (N_11308,N_6430,N_8837);
nor U11309 (N_11309,N_5874,N_9233);
xor U11310 (N_11310,N_8171,N_5563);
and U11311 (N_11311,N_9366,N_7911);
nor U11312 (N_11312,N_7249,N_5994);
nand U11313 (N_11313,N_7835,N_7181);
xor U11314 (N_11314,N_7352,N_7686);
and U11315 (N_11315,N_7677,N_5291);
nor U11316 (N_11316,N_5231,N_9373);
and U11317 (N_11317,N_8786,N_5407);
or U11318 (N_11318,N_9467,N_5888);
or U11319 (N_11319,N_9304,N_8089);
and U11320 (N_11320,N_7103,N_9151);
xnor U11321 (N_11321,N_7448,N_9886);
nand U11322 (N_11322,N_5429,N_7598);
and U11323 (N_11323,N_9256,N_6533);
nand U11324 (N_11324,N_8434,N_6854);
nor U11325 (N_11325,N_6949,N_8284);
nand U11326 (N_11326,N_6213,N_6123);
nand U11327 (N_11327,N_5437,N_5438);
nor U11328 (N_11328,N_8773,N_6374);
nand U11329 (N_11329,N_8024,N_8630);
nand U11330 (N_11330,N_7356,N_9662);
nand U11331 (N_11331,N_5615,N_9280);
nor U11332 (N_11332,N_9268,N_5484);
xnor U11333 (N_11333,N_6504,N_8251);
xnor U11334 (N_11334,N_9128,N_6094);
nor U11335 (N_11335,N_5680,N_8423);
or U11336 (N_11336,N_6138,N_5822);
or U11337 (N_11337,N_5954,N_9708);
or U11338 (N_11338,N_5736,N_9147);
and U11339 (N_11339,N_7728,N_9352);
or U11340 (N_11340,N_6364,N_6838);
or U11341 (N_11341,N_9143,N_8471);
and U11342 (N_11342,N_7546,N_7984);
or U11343 (N_11343,N_7168,N_9550);
nor U11344 (N_11344,N_8829,N_7584);
or U11345 (N_11345,N_7638,N_9537);
and U11346 (N_11346,N_5243,N_6062);
or U11347 (N_11347,N_7855,N_6461);
and U11348 (N_11348,N_9661,N_7202);
and U11349 (N_11349,N_8985,N_5259);
xor U11350 (N_11350,N_6763,N_6105);
nand U11351 (N_11351,N_9564,N_6080);
nor U11352 (N_11352,N_7716,N_5590);
nor U11353 (N_11353,N_5260,N_7009);
and U11354 (N_11354,N_6836,N_7838);
or U11355 (N_11355,N_6169,N_6745);
nor U11356 (N_11356,N_9446,N_6942);
xor U11357 (N_11357,N_8440,N_5301);
and U11358 (N_11358,N_8644,N_5561);
and U11359 (N_11359,N_5409,N_8108);
or U11360 (N_11360,N_8910,N_7680);
nand U11361 (N_11361,N_8582,N_9331);
or U11362 (N_11362,N_7991,N_8463);
or U11363 (N_11363,N_6919,N_6791);
or U11364 (N_11364,N_6010,N_9913);
nor U11365 (N_11365,N_9413,N_8091);
or U11366 (N_11366,N_9288,N_8680);
nor U11367 (N_11367,N_7066,N_9302);
or U11368 (N_11368,N_8280,N_7722);
and U11369 (N_11369,N_6290,N_8191);
xor U11370 (N_11370,N_5851,N_8356);
nor U11371 (N_11371,N_5579,N_5220);
or U11372 (N_11372,N_6337,N_9330);
xor U11373 (N_11373,N_8426,N_6648);
and U11374 (N_11374,N_8022,N_9186);
xnor U11375 (N_11375,N_6835,N_7065);
nor U11376 (N_11376,N_7163,N_5101);
xor U11377 (N_11377,N_7112,N_7076);
nand U11378 (N_11378,N_7715,N_5937);
nor U11379 (N_11379,N_6071,N_6873);
nor U11380 (N_11380,N_7491,N_6865);
and U11381 (N_11381,N_5022,N_5457);
nor U11382 (N_11382,N_6620,N_8513);
nand U11383 (N_11383,N_9670,N_6172);
nor U11384 (N_11384,N_5156,N_8071);
xnor U11385 (N_11385,N_8353,N_6343);
nand U11386 (N_11386,N_8122,N_8760);
xor U11387 (N_11387,N_5515,N_7178);
and U11388 (N_11388,N_5249,N_5153);
or U11389 (N_11389,N_7397,N_6072);
xor U11390 (N_11390,N_8095,N_6951);
nand U11391 (N_11391,N_8230,N_7100);
and U11392 (N_11392,N_6661,N_8116);
nor U11393 (N_11393,N_8199,N_6491);
or U11394 (N_11394,N_9739,N_6450);
xnor U11395 (N_11395,N_8328,N_9899);
xnor U11396 (N_11396,N_5798,N_8794);
xor U11397 (N_11397,N_9355,N_5811);
and U11398 (N_11398,N_6926,N_7814);
nand U11399 (N_11399,N_6481,N_8070);
xnor U11400 (N_11400,N_6317,N_8950);
and U11401 (N_11401,N_9311,N_9552);
xor U11402 (N_11402,N_9783,N_5939);
nand U11403 (N_11403,N_6767,N_6476);
or U11404 (N_11404,N_8673,N_6990);
and U11405 (N_11405,N_8787,N_6414);
and U11406 (N_11406,N_5514,N_6408);
nand U11407 (N_11407,N_9806,N_9118);
nor U11408 (N_11408,N_8986,N_6931);
and U11409 (N_11409,N_9804,N_8603);
nor U11410 (N_11410,N_6598,N_6208);
nand U11411 (N_11411,N_6556,N_6466);
nor U11412 (N_11412,N_5454,N_9262);
nand U11413 (N_11413,N_9185,N_7262);
nand U11414 (N_11414,N_8594,N_6765);
xor U11415 (N_11415,N_7688,N_9159);
nand U11416 (N_11416,N_7873,N_8507);
and U11417 (N_11417,N_7117,N_9825);
and U11418 (N_11418,N_9483,N_5767);
or U11419 (N_11419,N_9253,N_7368);
nor U11420 (N_11420,N_8618,N_8805);
or U11421 (N_11421,N_7027,N_7969);
nand U11422 (N_11422,N_6819,N_9575);
nor U11423 (N_11423,N_5149,N_8528);
nor U11424 (N_11424,N_7915,N_6447);
nand U11425 (N_11425,N_8077,N_7392);
xor U11426 (N_11426,N_7896,N_9182);
and U11427 (N_11427,N_6354,N_8457);
and U11428 (N_11428,N_9112,N_8044);
and U11429 (N_11429,N_9415,N_9168);
or U11430 (N_11430,N_5796,N_7798);
nor U11431 (N_11431,N_6054,N_7899);
nor U11432 (N_11432,N_9097,N_9098);
xnor U11433 (N_11433,N_6088,N_6257);
nor U11434 (N_11434,N_6832,N_8277);
nand U11435 (N_11435,N_9542,N_9391);
nand U11436 (N_11436,N_8425,N_5965);
xor U11437 (N_11437,N_6672,N_8543);
or U11438 (N_11438,N_8516,N_9165);
nand U11439 (N_11439,N_5061,N_6704);
and U11440 (N_11440,N_5386,N_5263);
or U11441 (N_11441,N_9139,N_7357);
nand U11442 (N_11442,N_6361,N_7531);
xor U11443 (N_11443,N_9222,N_8638);
nand U11444 (N_11444,N_5862,N_6122);
nand U11445 (N_11445,N_6705,N_7205);
xnor U11446 (N_11446,N_9438,N_7327);
or U11447 (N_11447,N_5704,N_9901);
xor U11448 (N_11448,N_8352,N_9950);
nand U11449 (N_11449,N_6750,N_7146);
xnor U11450 (N_11450,N_9077,N_9220);
or U11451 (N_11451,N_9236,N_7821);
and U11452 (N_11452,N_8905,N_6422);
and U11453 (N_11453,N_5015,N_6892);
nand U11454 (N_11454,N_9820,N_5369);
and U11455 (N_11455,N_7451,N_8613);
nor U11456 (N_11456,N_6997,N_9086);
nand U11457 (N_11457,N_7167,N_9906);
nor U11458 (N_11458,N_8485,N_7945);
xnor U11459 (N_11459,N_6137,N_9216);
and U11460 (N_11460,N_6207,N_9800);
nor U11461 (N_11461,N_8019,N_8076);
xor U11462 (N_11462,N_6954,N_8830);
nor U11463 (N_11463,N_5460,N_5106);
nor U11464 (N_11464,N_8726,N_6443);
or U11465 (N_11465,N_8704,N_9395);
nand U11466 (N_11466,N_6880,N_6142);
and U11467 (N_11467,N_8393,N_6503);
nor U11468 (N_11468,N_6040,N_7947);
nand U11469 (N_11469,N_7175,N_5311);
or U11470 (N_11470,N_8209,N_6869);
nand U11471 (N_11471,N_5131,N_5799);
nand U11472 (N_11472,N_6355,N_7525);
nand U11473 (N_11473,N_6008,N_5385);
xor U11474 (N_11474,N_5682,N_5881);
or U11475 (N_11475,N_6241,N_9290);
nand U11476 (N_11476,N_6527,N_7900);
nand U11477 (N_11477,N_5506,N_9172);
nand U11478 (N_11478,N_5267,N_7624);
nand U11479 (N_11479,N_6059,N_7143);
nor U11480 (N_11480,N_6540,N_7133);
nand U11481 (N_11481,N_7623,N_6276);
nand U11482 (N_11482,N_7676,N_8245);
nand U11483 (N_11483,N_8755,N_5897);
and U11484 (N_11484,N_7371,N_5431);
nor U11485 (N_11485,N_7636,N_5902);
nand U11486 (N_11486,N_6899,N_9993);
and U11487 (N_11487,N_5576,N_7176);
nand U11488 (N_11488,N_5080,N_6631);
nand U11489 (N_11489,N_9921,N_6107);
and U11490 (N_11490,N_9480,N_5947);
or U11491 (N_11491,N_8857,N_6112);
nand U11492 (N_11492,N_5185,N_5098);
or U11493 (N_11493,N_6966,N_9205);
and U11494 (N_11494,N_7690,N_9835);
and U11495 (N_11495,N_6611,N_7096);
nand U11496 (N_11496,N_6140,N_9070);
nor U11497 (N_11497,N_5689,N_6212);
and U11498 (N_11498,N_8744,N_5083);
nor U11499 (N_11499,N_7196,N_7261);
nand U11500 (N_11500,N_7222,N_8298);
nor U11501 (N_11501,N_5691,N_5093);
or U11502 (N_11502,N_8866,N_7234);
xor U11503 (N_11503,N_6046,N_9364);
nand U11504 (N_11504,N_5711,N_8811);
and U11505 (N_11505,N_5335,N_9528);
nand U11506 (N_11506,N_8878,N_6375);
or U11507 (N_11507,N_6243,N_8383);
nand U11508 (N_11508,N_6035,N_8201);
and U11509 (N_11509,N_9932,N_9009);
or U11510 (N_11510,N_8168,N_6227);
xnor U11511 (N_11511,N_7938,N_7789);
nand U11512 (N_11512,N_9978,N_7801);
nand U11513 (N_11513,N_5122,N_7607);
nand U11514 (N_11514,N_5946,N_8269);
or U11515 (N_11515,N_6412,N_6912);
or U11516 (N_11516,N_8117,N_7247);
and U11517 (N_11517,N_9179,N_9146);
nand U11518 (N_11518,N_6229,N_8501);
or U11519 (N_11519,N_6680,N_6602);
nor U11520 (N_11520,N_7048,N_5491);
nor U11521 (N_11521,N_9204,N_5321);
xnor U11522 (N_11522,N_6168,N_9620);
or U11523 (N_11523,N_7070,N_7487);
nor U11524 (N_11524,N_7917,N_9411);
xor U11525 (N_11525,N_9276,N_5464);
or U11526 (N_11526,N_6340,N_5268);
and U11527 (N_11527,N_7612,N_7290);
xor U11528 (N_11528,N_9087,N_7994);
xor U11529 (N_11529,N_7185,N_6502);
nand U11530 (N_11530,N_9573,N_6590);
or U11531 (N_11531,N_6641,N_9523);
nand U11532 (N_11532,N_9048,N_8073);
or U11533 (N_11533,N_6988,N_6833);
and U11534 (N_11534,N_5550,N_8186);
nor U11535 (N_11535,N_9500,N_6902);
nand U11536 (N_11536,N_5145,N_9960);
and U11537 (N_11537,N_9852,N_9123);
nand U11538 (N_11538,N_7404,N_6585);
or U11539 (N_11539,N_5894,N_5284);
and U11540 (N_11540,N_5570,N_5728);
or U11541 (N_11541,N_7118,N_7996);
and U11542 (N_11542,N_5483,N_6829);
xor U11543 (N_11543,N_7486,N_6569);
nor U11544 (N_11544,N_8234,N_9069);
nand U11545 (N_11545,N_8093,N_9037);
nor U11546 (N_11546,N_6924,N_5308);
or U11547 (N_11547,N_6849,N_6047);
nand U11548 (N_11548,N_6786,N_8864);
nand U11549 (N_11549,N_6953,N_8487);
or U11550 (N_11550,N_6231,N_5756);
nor U11551 (N_11551,N_8718,N_6772);
and U11552 (N_11552,N_9859,N_6534);
or U11553 (N_11553,N_6894,N_6643);
xnor U11554 (N_11554,N_7281,N_7975);
and U11555 (N_11555,N_7432,N_7977);
or U11556 (N_11556,N_5273,N_5209);
or U11557 (N_11557,N_8727,N_9889);
nor U11558 (N_11558,N_5350,N_8599);
or U11559 (N_11559,N_6264,N_7494);
nor U11560 (N_11560,N_7621,N_9757);
or U11561 (N_11561,N_7144,N_5626);
or U11562 (N_11562,N_7020,N_5428);
or U11563 (N_11563,N_6927,N_5761);
xor U11564 (N_11564,N_8706,N_7774);
or U11565 (N_11565,N_7350,N_7632);
nand U11566 (N_11566,N_9891,N_9647);
xor U11567 (N_11567,N_8349,N_6967);
or U11568 (N_11568,N_9342,N_8605);
or U11569 (N_11569,N_6293,N_6732);
or U11570 (N_11570,N_9058,N_7220);
or U11571 (N_11571,N_8338,N_7006);
and U11572 (N_11572,N_7802,N_5105);
or U11573 (N_11573,N_6529,N_5625);
or U11574 (N_11574,N_8862,N_7541);
or U11575 (N_11575,N_5069,N_8625);
nand U11576 (N_11576,N_5935,N_6711);
nand U11577 (N_11577,N_6780,N_9839);
and U11578 (N_11578,N_8519,N_8131);
and U11579 (N_11579,N_5980,N_5379);
and U11580 (N_11580,N_9732,N_9710);
nand U11581 (N_11581,N_8041,N_6493);
or U11582 (N_11582,N_8526,N_7665);
nor U11583 (N_11583,N_6737,N_7394);
or U11584 (N_11584,N_6824,N_8871);
nand U11585 (N_11585,N_6980,N_6462);
xnor U11586 (N_11586,N_8655,N_7884);
xor U11587 (N_11587,N_5966,N_6499);
xor U11588 (N_11588,N_6879,N_8121);
xor U11589 (N_11589,N_6073,N_6764);
xnor U11590 (N_11590,N_7141,N_7740);
and U11591 (N_11591,N_8018,N_6162);
nand U11592 (N_11592,N_9722,N_7039);
and U11593 (N_11593,N_6204,N_7061);
and U11594 (N_11594,N_6758,N_9576);
or U11595 (N_11595,N_5640,N_7888);
and U11596 (N_11596,N_6147,N_9547);
or U11597 (N_11597,N_7980,N_5096);
and U11598 (N_11598,N_9974,N_6994);
xor U11599 (N_11599,N_9829,N_7868);
or U11600 (N_11600,N_8324,N_5593);
xnor U11601 (N_11601,N_5698,N_5265);
xnor U11602 (N_11602,N_8587,N_8984);
and U11603 (N_11603,N_7805,N_9389);
nor U11604 (N_11604,N_9827,N_7495);
nor U11605 (N_11605,N_7993,N_8332);
xnor U11606 (N_11606,N_7400,N_8992);
nand U11607 (N_11607,N_7440,N_8106);
and U11608 (N_11608,N_7095,N_7295);
nor U11609 (N_11609,N_6341,N_5190);
and U11610 (N_11610,N_9350,N_5987);
and U11611 (N_11611,N_8693,N_7465);
nor U11612 (N_11612,N_5248,N_5823);
or U11613 (N_11613,N_7719,N_9927);
or U11614 (N_11614,N_6111,N_8684);
and U11615 (N_11615,N_8523,N_7809);
nand U11616 (N_11616,N_6535,N_5605);
or U11617 (N_11617,N_5686,N_9765);
xnor U11618 (N_11618,N_8367,N_5502);
or U11619 (N_11619,N_9108,N_5399);
or U11620 (N_11620,N_5327,N_7877);
nand U11621 (N_11621,N_6146,N_9135);
nand U11622 (N_11622,N_5899,N_8336);
nand U11623 (N_11623,N_5318,N_9381);
xor U11624 (N_11624,N_9356,N_7919);
nand U11625 (N_11625,N_8884,N_7307);
nor U11626 (N_11626,N_9289,N_8801);
nand U11627 (N_11627,N_8198,N_9178);
nor U11628 (N_11628,N_9032,N_6268);
and U11629 (N_11629,N_8333,N_8260);
xnor U11630 (N_11630,N_6677,N_9870);
or U11631 (N_11631,N_8821,N_8667);
and U11632 (N_11632,N_7139,N_6362);
xor U11633 (N_11633,N_5417,N_5555);
nand U11634 (N_11634,N_9369,N_7653);
or U11635 (N_11635,N_7850,N_9113);
nand U11636 (N_11636,N_7817,N_5216);
and U11637 (N_11637,N_9416,N_5970);
nand U11638 (N_11638,N_6253,N_7348);
and U11639 (N_11639,N_8512,N_5791);
and U11640 (N_11640,N_8881,N_9324);
nand U11641 (N_11641,N_9956,N_6452);
or U11642 (N_11642,N_6733,N_6806);
and U11643 (N_11643,N_8015,N_8740);
nand U11644 (N_11644,N_7767,N_7322);
nor U11645 (N_11645,N_5747,N_7866);
xor U11646 (N_11646,N_9860,N_9907);
or U11647 (N_11647,N_7699,N_9752);
nand U11648 (N_11648,N_7127,N_9988);
and U11649 (N_11649,N_6314,N_9857);
xnor U11650 (N_11650,N_5435,N_6463);
and U11651 (N_11651,N_9729,N_8402);
nand U11652 (N_11652,N_5906,N_8852);
and U11653 (N_11653,N_8616,N_7208);
xnor U11654 (N_11654,N_6434,N_5229);
or U11655 (N_11655,N_5658,N_6900);
xnor U11656 (N_11656,N_8607,N_5380);
nand U11657 (N_11657,N_6473,N_9716);
nand U11658 (N_11658,N_7921,N_8641);
nor U11659 (N_11659,N_8271,N_9388);
xnor U11660 (N_11660,N_7361,N_9133);
xor U11661 (N_11661,N_9544,N_9379);
and U11662 (N_11662,N_8579,N_7936);
or U11663 (N_11663,N_7926,N_6117);
or U11664 (N_11664,N_7399,N_8855);
or U11665 (N_11665,N_5352,N_8784);
nor U11666 (N_11666,N_5447,N_7455);
xor U11667 (N_11667,N_8735,N_5883);
xnor U11668 (N_11668,N_9705,N_7535);
xor U11669 (N_11669,N_9773,N_5453);
and U11670 (N_11670,N_8606,N_6301);
and U11671 (N_11671,N_6831,N_9679);
xor U11672 (N_11672,N_5909,N_5755);
nor U11673 (N_11673,N_8968,N_6305);
nand U11674 (N_11674,N_5744,N_8052);
nor U11675 (N_11675,N_6055,N_8180);
and U11676 (N_11676,N_9450,N_7393);
xor U11677 (N_11677,N_9192,N_8987);
or U11678 (N_11678,N_7721,N_5272);
and U11679 (N_11679,N_5734,N_5494);
nor U11680 (N_11680,N_9538,N_7193);
xor U11681 (N_11681,N_9726,N_5117);
or U11682 (N_11682,N_9674,N_8161);
or U11683 (N_11683,N_8462,N_8129);
nand U11684 (N_11684,N_9224,N_8048);
or U11685 (N_11685,N_6506,N_9558);
nor U11686 (N_11686,N_7406,N_9360);
nand U11687 (N_11687,N_8631,N_7153);
nor U11688 (N_11688,N_8554,N_6292);
xor U11689 (N_11689,N_6625,N_8983);
or U11690 (N_11690,N_6956,N_9557);
nand U11691 (N_11691,N_5411,N_6738);
or U11692 (N_11692,N_5058,N_8799);
or U11693 (N_11693,N_6082,N_7200);
and U11694 (N_11694,N_5449,N_9579);
nand U11695 (N_11695,N_5047,N_7707);
xor U11696 (N_11696,N_8619,N_7646);
xnor U11697 (N_11697,N_5702,N_9241);
and U11698 (N_11698,N_8917,N_7369);
nor U11699 (N_11699,N_6121,N_8510);
nand U11700 (N_11700,N_6813,N_9235);
and U11701 (N_11701,N_6053,N_8989);
nor U11702 (N_11702,N_9124,N_6822);
or U11703 (N_11703,N_6357,N_8290);
nand U11704 (N_11704,N_9099,N_8562);
nand U11705 (N_11705,N_6799,N_6548);
xnor U11706 (N_11706,N_8967,N_7106);
nand U11707 (N_11707,N_7293,N_5366);
nor U11708 (N_11708,N_7493,N_6840);
nor U11709 (N_11709,N_6078,N_7251);
nor U11710 (N_11710,N_5928,N_8895);
nand U11711 (N_11711,N_7500,N_8921);
nor U11712 (N_11712,N_8696,N_8196);
xnor U11713 (N_11713,N_6538,N_9761);
nand U11714 (N_11714,N_8493,N_6181);
nand U11715 (N_11715,N_9531,N_9074);
and U11716 (N_11716,N_9850,N_5801);
nor U11717 (N_11717,N_7586,N_7615);
nand U11718 (N_11718,N_6578,N_6026);
nand U11719 (N_11719,N_9338,N_8453);
and U11720 (N_11720,N_9271,N_8663);
and U11721 (N_11721,N_6993,N_8195);
nand U11722 (N_11722,N_5345,N_9083);
and U11723 (N_11723,N_6945,N_6617);
or U11724 (N_11724,N_5203,N_8868);
or U11725 (N_11725,N_9193,N_8498);
nor U11726 (N_11726,N_7569,N_9174);
nor U11727 (N_11727,N_6194,N_8559);
and U11728 (N_11728,N_6027,N_5451);
nand U11729 (N_11729,N_9045,N_5882);
nand U11730 (N_11730,N_6539,N_6673);
or U11731 (N_11731,N_9717,N_7342);
or U11732 (N_11732,N_6827,N_7633);
nand U11733 (N_11733,N_7438,N_5115);
nor U11734 (N_11734,N_9244,N_7452);
nand U11735 (N_11735,N_7934,N_7282);
and U11736 (N_11736,N_5362,N_7385);
xnor U11737 (N_11737,N_5412,N_6074);
nor U11738 (N_11738,N_7946,N_7035);
and U11739 (N_11739,N_8751,N_5419);
or U11740 (N_11740,N_6420,N_9004);
nor U11741 (N_11741,N_7326,N_5551);
xnor U11742 (N_11742,N_7961,N_6925);
nor U11743 (N_11743,N_9862,N_7045);
nor U11744 (N_11744,N_8716,N_6803);
nand U11745 (N_11745,N_7430,N_6642);
xnor U11746 (N_11746,N_7030,N_5128);
and U11747 (N_11747,N_6064,N_8688);
nand U11748 (N_11748,N_9465,N_7231);
nand U11749 (N_11749,N_5198,N_8016);
nor U11750 (N_11750,N_6537,N_5860);
and U11751 (N_11751,N_5583,N_9042);
and U11752 (N_11752,N_9434,N_6024);
nor U11753 (N_11753,N_5745,N_6593);
nor U11754 (N_11754,N_6947,N_5949);
nand U11755 (N_11755,N_9623,N_5951);
nand U11756 (N_11756,N_8506,N_9326);
nor U11757 (N_11757,N_5891,N_9403);
nor U11758 (N_11758,N_6419,N_5477);
xor U11759 (N_11759,N_6666,N_9479);
or U11760 (N_11760,N_5215,N_5322);
nor U11761 (N_11761,N_8731,N_9195);
and U11762 (N_11762,N_6561,N_6995);
nor U11763 (N_11763,N_6058,N_6382);
xor U11764 (N_11764,N_9884,N_7931);
or U11765 (N_11765,N_6867,N_9361);
and U11766 (N_11766,N_7002,N_5140);
or U11767 (N_11767,N_5307,N_7259);
xor U11768 (N_11768,N_7203,N_6601);
nor U11769 (N_11769,N_8996,N_6398);
or U11770 (N_11770,N_7897,N_6174);
and U11771 (N_11771,N_9156,N_5029);
nor U11772 (N_11772,N_6545,N_8841);
nor U11773 (N_11773,N_5662,N_7617);
nor U11774 (N_11774,N_7427,N_6079);
and U11775 (N_11775,N_5094,N_5397);
xor U11776 (N_11776,N_8982,N_9979);
or U11777 (N_11777,N_5536,N_9521);
xor U11778 (N_11778,N_6265,N_8270);
xor U11779 (N_11779,N_6069,N_7016);
xor U11780 (N_11780,N_7908,N_6706);
nor U11781 (N_11781,N_8571,N_8045);
and U11782 (N_11782,N_8208,N_9833);
or U11783 (N_11783,N_6935,N_9570);
nand U11784 (N_11784,N_8976,N_9340);
or U11785 (N_11785,N_5330,N_9451);
and U11786 (N_11786,N_7845,N_9983);
xor U11787 (N_11787,N_7005,N_8782);
xor U11788 (N_11788,N_8486,N_5034);
xnor U11789 (N_11789,N_5392,N_6036);
xor U11790 (N_11790,N_6721,N_7062);
nor U11791 (N_11791,N_5400,N_8370);
xor U11792 (N_11792,N_6441,N_5495);
nand U11793 (N_11793,N_8818,N_7891);
xor U11794 (N_11794,N_7973,N_6096);
or U11795 (N_11795,N_8964,N_8555);
nand U11796 (N_11796,N_5741,N_5917);
xnor U11797 (N_11797,N_5100,N_5332);
nor U11798 (N_11798,N_9615,N_6206);
or U11799 (N_11799,N_5624,N_8800);
or U11800 (N_11800,N_9287,N_7484);
and U11801 (N_11801,N_9259,N_5696);
and U11802 (N_11802,N_5815,N_9417);
or U11803 (N_11803,N_6846,N_7520);
or U11804 (N_11804,N_9796,N_8257);
nor U11805 (N_11805,N_7999,N_9724);
or U11806 (N_11806,N_5173,N_7148);
xnor U11807 (N_11807,N_8123,N_5365);
nand U11808 (N_11808,N_8068,N_9409);
xnor U11809 (N_11809,N_6583,N_6866);
nor U11810 (N_11810,N_7155,N_6897);
and U11811 (N_11811,N_8748,N_8378);
xor U11812 (N_11812,N_6120,N_5525);
nand U11813 (N_11813,N_9768,N_5314);
xnor U11814 (N_11814,N_8211,N_7415);
and U11815 (N_11815,N_9080,N_9487);
nor U11816 (N_11816,N_5232,N_8711);
xor U11817 (N_11817,N_9545,N_8146);
nand U11818 (N_11818,N_5275,N_7536);
nand U11819 (N_11819,N_7381,N_5887);
nor U11820 (N_11820,N_7104,N_9813);
and U11821 (N_11821,N_8142,N_9769);
and U11822 (N_11822,N_6979,N_7252);
nor U11823 (N_11823,N_6702,N_7072);
or U11824 (N_11824,N_6244,N_8614);
nand U11825 (N_11825,N_6377,N_6342);
nand U11826 (N_11826,N_7657,N_7683);
nand U11827 (N_11827,N_9866,N_9965);
xnor U11828 (N_11828,N_9637,N_7454);
nand U11829 (N_11829,N_6720,N_6691);
xor U11830 (N_11830,N_7734,N_8326);
and U11831 (N_11831,N_8991,N_5224);
nand U11832 (N_11832,N_5631,N_8477);
or U11833 (N_11833,N_7890,N_8975);
or U11834 (N_11834,N_8557,N_9449);
nor U11835 (N_11835,N_6139,N_5934);
xor U11836 (N_11836,N_9626,N_8220);
and U11837 (N_11837,N_8363,N_6592);
nand U11838 (N_11838,N_7358,N_5672);
nor U11839 (N_11839,N_9933,N_8903);
and U11840 (N_11840,N_7380,N_7557);
or U11841 (N_11841,N_8204,N_8384);
nor U11842 (N_11842,N_5900,N_7856);
or U11843 (N_11843,N_7950,N_5258);
nor U11844 (N_11844,N_6380,N_6589);
nor U11845 (N_11845,N_7788,N_8318);
and U11846 (N_11846,N_7731,N_9050);
xor U11847 (N_11847,N_7459,N_5054);
nand U11848 (N_11848,N_7362,N_7311);
nand U11849 (N_11849,N_7776,N_5743);
and U11850 (N_11850,N_8738,N_8429);
and U11851 (N_11851,N_6367,N_9514);
or U11852 (N_11852,N_8648,N_7704);
nand U11853 (N_11853,N_6099,N_7457);
nor U11854 (N_11854,N_8475,N_5771);
nor U11855 (N_11855,N_9117,N_8190);
nand U11856 (N_11856,N_7956,N_7955);
xor U11857 (N_11857,N_7501,N_9266);
nor U11858 (N_11858,N_9879,N_6922);
nor U11859 (N_11859,N_9606,N_5852);
or U11860 (N_11860,N_8405,N_5373);
nor U11861 (N_11861,N_7313,N_5890);
and U11862 (N_11862,N_9478,N_8911);
nand U11863 (N_11863,N_6211,N_9704);
nand U11864 (N_11864,N_6671,N_5867);
or U11865 (N_11865,N_8373,N_7652);
or U11866 (N_11866,N_8529,N_5102);
xor U11867 (N_11867,N_6368,N_8241);
and U11868 (N_11868,N_6694,N_5271);
nor U11869 (N_11869,N_5847,N_6475);
nor U11870 (N_11870,N_6753,N_8104);
and U11871 (N_11871,N_9023,N_9714);
nand U11872 (N_11872,N_6936,N_8228);
nand U11873 (N_11873,N_5436,N_7040);
or U11874 (N_11874,N_5614,N_9951);
xor U11875 (N_11875,N_6429,N_5383);
and U11876 (N_11876,N_8544,N_6417);
xor U11877 (N_11877,N_6893,N_8920);
and U11878 (N_11878,N_8411,N_6075);
nand U11879 (N_11879,N_7107,N_5647);
and U11880 (N_11880,N_9282,N_9384);
and U11881 (N_11881,N_6746,N_7339);
or U11882 (N_11882,N_7772,N_7360);
nand U11883 (N_11883,N_6456,N_6663);
and U11884 (N_11884,N_7909,N_8027);
nand U11885 (N_11885,N_9749,N_7379);
or U11886 (N_11886,N_5552,N_6982);
nand U11887 (N_11887,N_6703,N_6262);
and U11888 (N_11888,N_7028,N_7849);
xor U11889 (N_11889,N_6315,N_5584);
and U11890 (N_11890,N_5337,N_6330);
nand U11891 (N_11891,N_6148,N_6065);
nor U11892 (N_11892,N_9078,N_7645);
and U11893 (N_11893,N_6438,N_6056);
nand U11894 (N_11894,N_7221,N_5694);
nand U11895 (N_11895,N_5312,N_7784);
nor U11896 (N_11896,N_8445,N_5136);
or U11897 (N_11897,N_8914,N_9645);
nand U11898 (N_11898,N_8452,N_6118);
nand U11899 (N_11899,N_6845,N_5766);
xnor U11900 (N_11900,N_8695,N_8635);
xor U11901 (N_11901,N_5269,N_7898);
or U11902 (N_11902,N_7037,N_5846);
nor U11903 (N_11903,N_9601,N_8812);
or U11904 (N_11904,N_7604,N_6834);
or U11905 (N_11905,N_6185,N_8145);
nor U11906 (N_11906,N_5636,N_8525);
nand U11907 (N_11907,N_5095,N_6409);
and U11908 (N_11908,N_7790,N_6485);
nor U11909 (N_11909,N_7426,N_9925);
nor U11910 (N_11910,N_7332,N_7519);
nor U11911 (N_11911,N_5003,N_6776);
nand U11912 (N_11912,N_8596,N_7600);
nor U11913 (N_11913,N_6070,N_9581);
nand U11914 (N_11914,N_7509,N_8860);
nand U11915 (N_11915,N_7151,N_5988);
and U11916 (N_11916,N_6498,N_8214);
nor U11917 (N_11917,N_7204,N_8394);
nor U11918 (N_11918,N_5776,N_7197);
nand U11919 (N_11919,N_8420,N_7186);
and U11920 (N_11920,N_8458,N_6853);
xnor U11921 (N_11921,N_6920,N_6258);
nand U11922 (N_11922,N_9822,N_9111);
or U11923 (N_11923,N_8729,N_8080);
xor U11924 (N_11924,N_9608,N_9510);
nor U11925 (N_11925,N_6004,N_5459);
nand U11926 (N_11926,N_8776,N_5666);
xor U11927 (N_11927,N_8825,N_8889);
or U11928 (N_11928,N_6619,N_7628);
or U11929 (N_11929,N_8762,N_7579);
nand U11930 (N_11930,N_9629,N_5660);
nand U11931 (N_11931,N_9158,N_7053);
nand U11932 (N_11932,N_5410,N_8105);
and U11933 (N_11933,N_5621,N_9871);
or U11934 (N_11934,N_7872,N_9701);
nor U11935 (N_11935,N_8417,N_7779);
nor U11936 (N_11936,N_6157,N_5849);
nand U11937 (N_11937,N_5404,N_7595);
and U11938 (N_11938,N_9421,N_8309);
or U11939 (N_11939,N_6728,N_6351);
nand U11940 (N_11940,N_9120,N_8552);
and U11941 (N_11941,N_8750,N_9841);
or U11942 (N_11942,N_9215,N_7553);
nand U11943 (N_11943,N_6546,N_7545);
or U11944 (N_11944,N_8977,N_7160);
or U11945 (N_11945,N_7492,N_5653);
or U11946 (N_11946,N_8724,N_8151);
nor U11947 (N_11947,N_6964,N_9996);
nand U11948 (N_11948,N_9815,N_8856);
or U11949 (N_11949,N_5712,N_9737);
and U11950 (N_11950,N_9344,N_6487);
xor U11951 (N_11951,N_5344,N_5610);
or U11952 (N_11952,N_8988,N_8292);
or U11953 (N_11953,N_6338,N_6907);
xor U11954 (N_11954,N_5078,N_8883);
nand U11955 (N_11955,N_7041,N_7990);
or U11956 (N_11956,N_9394,N_7199);
or U11957 (N_11957,N_7150,N_9553);
and U11958 (N_11958,N_8707,N_5239);
nand U11959 (N_11959,N_8979,N_7777);
xor U11960 (N_11960,N_5528,N_9656);
and U11961 (N_11961,N_6724,N_7811);
nor U11962 (N_11962,N_6448,N_7015);
and U11963 (N_11963,N_9292,N_6801);
and U11964 (N_11964,N_6044,N_8182);
and U11965 (N_11965,N_7735,N_7537);
or U11966 (N_11966,N_7949,N_7782);
nand U11967 (N_11967,N_9766,N_8854);
nand U11968 (N_11968,N_7161,N_9973);
nor U11969 (N_11969,N_5313,N_8021);
nor U11970 (N_11970,N_6201,N_6459);
or U11971 (N_11971,N_5310,N_7269);
xor U11972 (N_11972,N_9093,N_7038);
nor U11973 (N_11973,N_7063,N_9026);
nor U11974 (N_11974,N_6465,N_8492);
and U11975 (N_11975,N_5048,N_5903);
and U11976 (N_11976,N_7264,N_9073);
or U11977 (N_11977,N_8366,N_9898);
nand U11978 (N_11978,N_9787,N_8135);
nand U11979 (N_11979,N_6278,N_7521);
nand U11980 (N_11980,N_9507,N_9580);
or U11981 (N_11981,N_9418,N_7412);
or U11982 (N_11982,N_9892,N_6591);
and U11983 (N_11983,N_8482,N_9261);
or U11984 (N_11984,N_7458,N_7294);
or U11985 (N_11985,N_8085,N_5737);
nor U11986 (N_11986,N_6159,N_8143);
xnor U11987 (N_11987,N_6445,N_8919);
and U11988 (N_11988,N_8656,N_7948);
nand U11989 (N_11989,N_9725,N_6127);
nor U11990 (N_11990,N_6451,N_6381);
or U11991 (N_11991,N_7280,N_9707);
and U11992 (N_11992,N_5789,N_6628);
or U11993 (N_11993,N_6482,N_6699);
xnor U11994 (N_11994,N_9245,N_9515);
nand U11995 (N_11995,N_6684,N_7577);
and U11996 (N_11996,N_8944,N_9591);
xnor U11997 (N_11997,N_8637,N_5848);
nor U11998 (N_11998,N_7478,N_8437);
nand U11999 (N_11999,N_9858,N_7302);
xnor U12000 (N_12000,N_6025,N_9578);
nor U12001 (N_12001,N_6649,N_9105);
and U12002 (N_12002,N_7927,N_5324);
nor U12003 (N_12003,N_6471,N_8890);
xnor U12004 (N_12004,N_5090,N_6446);
xor U12005 (N_12005,N_8473,N_5522);
nor U12006 (N_12006,N_6762,N_7547);
or U12007 (N_12007,N_6790,N_7918);
nand U12008 (N_12008,N_9635,N_9307);
xnor U12009 (N_12009,N_5202,N_5938);
nand U12010 (N_12010,N_8179,N_7194);
nand U12011 (N_12011,N_9908,N_6637);
or U12012 (N_12012,N_6635,N_8586);
and U12013 (N_12013,N_8942,N_6654);
nor U12014 (N_12014,N_6093,N_6234);
nor U12015 (N_12015,N_6049,N_5245);
nand U12016 (N_12016,N_8156,N_6690);
xnor U12017 (N_12017,N_9610,N_8109);
xor U12018 (N_12018,N_7658,N_6489);
xnor U12019 (N_12019,N_9638,N_6731);
nor U12020 (N_12020,N_5765,N_8565);
nor U12021 (N_12021,N_8702,N_6421);
nor U12022 (N_12022,N_8753,N_7654);
or U12023 (N_12023,N_5880,N_9125);
nor U12024 (N_12024,N_8545,N_9306);
nand U12025 (N_12025,N_9928,N_6014);
nor U12026 (N_12026,N_8531,N_9934);
or U12027 (N_12027,N_6783,N_6154);
or U12028 (N_12028,N_8351,N_9809);
nor U12029 (N_12029,N_5834,N_9230);
or U12030 (N_12030,N_9803,N_8465);
or U12031 (N_12031,N_5014,N_5182);
or U12032 (N_12032,N_8628,N_8098);
or U12033 (N_12033,N_7042,N_9377);
or U12034 (N_12034,N_7905,N_6932);
nand U12035 (N_12035,N_9962,N_7515);
xor U12036 (N_12036,N_9382,N_5241);
or U12037 (N_12037,N_6910,N_5019);
and U12038 (N_12038,N_9303,N_5674);
xor U12039 (N_12039,N_9212,N_8060);
nand U12040 (N_12040,N_8700,N_9672);
xnor U12041 (N_12041,N_7807,N_6872);
xnor U12042 (N_12042,N_6200,N_7179);
xor U12043 (N_12043,N_9713,N_6558);
or U12044 (N_12044,N_5869,N_7799);
and U12045 (N_12045,N_8075,N_8389);
or U12046 (N_12046,N_9938,N_7743);
or U12047 (N_12047,N_8072,N_9736);
and U12048 (N_12048,N_6393,N_5426);
nor U12049 (N_12049,N_7389,N_5785);
nand U12050 (N_12050,N_5632,N_7942);
nor U12051 (N_12051,N_5718,N_7456);
nor U12052 (N_12052,N_8327,N_6613);
xor U12053 (N_12053,N_8945,N_5361);
nor U12054 (N_12054,N_5467,N_8491);
nor U12055 (N_12055,N_5544,N_9201);
xor U12056 (N_12056,N_5710,N_6170);
nor U12057 (N_12057,N_6904,N_8908);
and U12058 (N_12058,N_6149,N_7316);
nand U12059 (N_12059,N_8621,N_5622);
and U12060 (N_12060,N_9834,N_5663);
and U12061 (N_12061,N_7701,N_9267);
or U12062 (N_12062,N_7228,N_8742);
xor U12063 (N_12063,N_5504,N_7528);
xnor U12064 (N_12064,N_5975,N_8551);
and U12065 (N_12065,N_6999,N_8972);
nand U12066 (N_12066,N_8764,N_5651);
and U12067 (N_12067,N_9758,N_8717);
or U12068 (N_12068,N_7542,N_9040);
and U12069 (N_12069,N_7463,N_6250);
nand U12070 (N_12070,N_6525,N_9945);
or U12071 (N_12071,N_5571,N_8149);
nand U12072 (N_12072,N_8436,N_6135);
nor U12073 (N_12073,N_7098,N_6864);
and U12074 (N_12074,N_7248,N_7130);
and U12075 (N_12075,N_8634,N_9943);
or U12076 (N_12076,N_5989,N_9919);
and U12077 (N_12077,N_5195,N_5510);
and U12078 (N_12078,N_9617,N_7229);
or U12079 (N_12079,N_9836,N_6771);
xnor U12080 (N_12080,N_9148,N_9607);
nor U12081 (N_12081,N_8126,N_5505);
nor U12082 (N_12082,N_7649,N_6906);
nand U12083 (N_12083,N_5057,N_7287);
and U12084 (N_12084,N_7858,N_6550);
xor U12085 (N_12085,N_5104,N_9281);
and U12086 (N_12086,N_8450,N_5359);
xor U12087 (N_12087,N_6248,N_7587);
or U12088 (N_12088,N_5011,N_5724);
nor U12089 (N_12089,N_9015,N_6057);
nor U12090 (N_12090,N_7218,N_7976);
xnor U12091 (N_12091,N_5709,N_5375);
nor U12092 (N_12092,N_8591,N_9167);
and U12093 (N_12093,N_8842,N_8956);
nor U12094 (N_12094,N_5196,N_6006);
nand U12095 (N_12095,N_6582,N_8574);
and U12096 (N_12096,N_5955,N_6416);
nand U12097 (N_12097,N_7933,N_8532);
nor U12098 (N_12098,N_7533,N_7755);
nor U12099 (N_12099,N_5415,N_7120);
and U12100 (N_12100,N_7571,N_8935);
xnor U12101 (N_12101,N_5807,N_8347);
nor U12102 (N_12102,N_8461,N_7808);
xnor U12103 (N_12103,N_7320,N_6518);
and U12104 (N_12104,N_6938,N_5416);
xor U12105 (N_12105,N_8611,N_6676);
and U12106 (N_12106,N_5089,N_5221);
nand U12107 (N_12107,N_6431,N_6193);
xnor U12108 (N_12108,N_5914,N_8456);
or U12109 (N_12109,N_7752,N_8990);
nand U12110 (N_12110,N_5677,N_8065);
or U12111 (N_12111,N_7923,N_9217);
nand U12112 (N_12112,N_9448,N_5762);
or U12113 (N_12113,N_6689,N_9140);
nand U12114 (N_12114,N_9171,N_9920);
and U12115 (N_12115,N_9177,N_9318);
nor U12116 (N_12116,N_8939,N_8494);
or U12117 (N_12117,N_7718,N_5609);
or U12118 (N_12118,N_7374,N_6449);
nand U12119 (N_12119,N_9018,N_6823);
or U12120 (N_12120,N_6847,N_6407);
and U12121 (N_12121,N_6716,N_7804);
or U12122 (N_12122,N_8495,N_8578);
nor U12123 (N_12123,N_5518,N_8615);
xnor U12124 (N_12124,N_9039,N_7725);
nand U12125 (N_12125,N_7754,N_7378);
and U12126 (N_12126,N_7922,N_8194);
nand U12127 (N_12127,N_8215,N_5132);
nor U12128 (N_12128,N_8258,N_8661);
nor U12129 (N_12129,N_7318,N_8339);
and U12130 (N_12130,N_5641,N_8134);
or U12131 (N_12131,N_6675,N_7986);
or U12132 (N_12132,N_9589,N_8055);
xnor U12133 (N_12133,N_7004,N_5948);
or U12134 (N_12134,N_5513,N_7904);
or U12135 (N_12135,N_8010,N_8719);
xor U12136 (N_12136,N_5587,N_9005);
and U12137 (N_12137,N_9533,N_9365);
xor U12138 (N_12138,N_6061,N_5836);
nand U12139 (N_12139,N_9622,N_9285);
and U12140 (N_12140,N_6948,N_6647);
xor U12141 (N_12141,N_6770,N_9849);
nand U12142 (N_12142,N_9585,N_9909);
nand U12143 (N_12143,N_8235,N_5859);
nand U12144 (N_12144,N_8806,N_6104);
xor U12145 (N_12145,N_6030,N_5565);
and U12146 (N_12146,N_7198,N_7590);
xor U12147 (N_12147,N_7169,N_5591);
xnor U12148 (N_12148,N_9398,N_7641);
nor U12149 (N_12149,N_7778,N_7826);
or U12150 (N_12150,N_7960,N_6759);
or U12151 (N_12151,N_8540,N_7166);
xnor U12152 (N_12152,N_9746,N_9351);
nor U12153 (N_12153,N_8288,N_6828);
nor U12154 (N_12154,N_5434,N_5130);
and U12155 (N_12155,N_9745,N_5523);
nand U12156 (N_12156,N_9750,N_7593);
or U12157 (N_12157,N_7372,N_6616);
and U12158 (N_12158,N_9034,N_9586);
and U12159 (N_12159,N_9431,N_9180);
or U12160 (N_12160,N_7862,N_9439);
and U12161 (N_12161,N_6133,N_7126);
nor U12162 (N_12162,N_7291,N_7694);
nand U12163 (N_12163,N_8059,N_7687);
nor U12164 (N_12164,N_8210,N_5678);
nor U12165 (N_12165,N_7983,N_6109);
or U12166 (N_12166,N_9375,N_7693);
nand U12167 (N_12167,N_6198,N_8380);
and U12168 (N_12168,N_8981,N_7012);
and U12169 (N_12169,N_7912,N_8330);
nand U12170 (N_12170,N_7453,N_8714);
nand U12171 (N_12171,N_9605,N_8272);
nor U12172 (N_12172,N_6883,N_8627);
nor U12173 (N_12173,N_6022,N_8558);
or U12174 (N_12174,N_9371,N_8164);
or U12175 (N_12175,N_5764,N_7237);
and U12176 (N_12176,N_6378,N_5174);
or U12177 (N_12177,N_7018,N_9170);
xor U12178 (N_12178,N_8278,N_9275);
nand U12179 (N_12179,N_5067,N_5238);
nor U12180 (N_12180,N_8589,N_5009);
nor U12181 (N_12181,N_7592,N_5981);
nor U12182 (N_12182,N_6933,N_9251);
xor U12183 (N_12183,N_5733,N_9541);
xor U12184 (N_12184,N_5233,N_6267);
nand U12185 (N_12185,N_7301,N_9433);
nand U12186 (N_12186,N_7309,N_8709);
and U12187 (N_12187,N_7123,N_9685);
nor U12188 (N_12188,N_5911,N_7820);
xnor U12189 (N_12189,N_6608,N_9247);
or U12190 (N_12190,N_7526,N_5097);
nor U12191 (N_12191,N_8138,N_7561);
nand U12192 (N_12192,N_6688,N_6279);
xor U12193 (N_12193,N_7419,N_7952);
nor U12194 (N_12194,N_7885,N_8177);
xor U12195 (N_12195,N_5432,N_9625);
nor U12196 (N_12196,N_6281,N_5084);
xor U12197 (N_12197,N_5372,N_5760);
nand U12198 (N_12198,N_9794,N_6640);
nor U12199 (N_12199,N_9534,N_8036);
nand U12200 (N_12200,N_9016,N_7236);
and U12201 (N_12201,N_8472,N_6565);
nand U12202 (N_12202,N_6304,N_8876);
and U12203 (N_12203,N_8354,N_5423);
nand U12204 (N_12204,N_6128,N_8584);
or U12205 (N_12205,N_6747,N_7275);
or U12206 (N_12206,N_9743,N_5952);
or U12207 (N_12207,N_8505,N_9997);
or U12208 (N_12208,N_5212,N_6656);
xnor U12209 (N_12209,N_9897,N_7413);
nand U12210 (N_12210,N_8870,N_5595);
and U12211 (N_12211,N_9944,N_9066);
xor U12212 (N_12212,N_7132,N_9208);
nand U12213 (N_12213,N_8561,N_6779);
or U12214 (N_12214,N_7305,N_6796);
nor U12215 (N_12215,N_9116,N_7941);
xor U12216 (N_12216,N_9594,N_9785);
and U12217 (N_12217,N_9462,N_6259);
nand U12218 (N_12218,N_8497,N_6097);
xnor U12219 (N_12219,N_9091,N_5222);
nand U12220 (N_12220,N_5597,N_8928);
nand U12221 (N_12221,N_6029,N_9660);
and U12222 (N_12222,N_7759,N_5898);
or U12223 (N_12223,N_5017,N_6599);
nor U12224 (N_12224,N_5072,N_6909);
or U12225 (N_12225,N_9295,N_9013);
or U12226 (N_12226,N_8115,N_7695);
xor U12227 (N_12227,N_7766,N_8564);
xor U12228 (N_12228,N_7323,N_5172);
and U12229 (N_12229,N_6180,N_5461);
and U12230 (N_12230,N_7183,N_7741);
and U12231 (N_12231,N_7376,N_9022);
xor U12232 (N_12232,N_5613,N_6802);
nand U12233 (N_12233,N_6522,N_8249);
nand U12234 (N_12234,N_9102,N_5803);
and U12235 (N_12235,N_8747,N_6402);
nand U12236 (N_12236,N_9372,N_9497);
nor U12237 (N_12237,N_6521,N_5279);
and U12238 (N_12238,N_9790,N_9692);
nor U12239 (N_12239,N_6679,N_9445);
and U12240 (N_12240,N_9272,N_7744);
and U12241 (N_12241,N_8011,N_9798);
nand U12242 (N_12242,N_9396,N_8953);
nor U12243 (N_12243,N_6346,N_7188);
or U12244 (N_12244,N_7124,N_7471);
and U12245 (N_12245,N_8433,N_8086);
or U12246 (N_12246,N_9160,N_9094);
nor U12247 (N_12247,N_6366,N_7162);
or U12248 (N_12248,N_6106,N_9930);
nand U12249 (N_12249,N_5879,N_6577);
nand U12250 (N_12250,N_6251,N_5923);
nand U12251 (N_12251,N_7750,N_9677);
or U12252 (N_12252,N_5112,N_5028);
xnor U12253 (N_12253,N_7503,N_6837);
nor U12254 (N_12254,N_7709,N_5141);
xnor U12255 (N_12255,N_9300,N_5176);
or U12256 (N_12256,N_9654,N_5151);
or U12257 (N_12257,N_9563,N_5384);
nor U12258 (N_12258,N_6579,N_9842);
and U12259 (N_12259,N_8054,N_9214);
nand U12260 (N_12260,N_5018,N_6812);
xor U12261 (N_12261,N_8047,N_5630);
nor U12262 (N_12262,N_7464,N_5541);
and U12263 (N_12263,N_7760,N_7982);
xor U12264 (N_12264,N_7164,N_9401);
and U12265 (N_12265,N_5499,N_7330);
xnor U12266 (N_12266,N_6494,N_5161);
xor U12267 (N_12267,N_6209,N_9134);
and U12268 (N_12268,N_9655,N_8775);
nand U12269 (N_12269,N_5146,N_5538);
nand U12270 (N_12270,N_6668,N_9392);
or U12271 (N_12271,N_9688,N_6032);
nor U12272 (N_12272,N_8157,N_8938);
nor U12273 (N_12273,N_9663,N_9786);
xor U12274 (N_12274,N_8480,N_5661);
or U12275 (N_12275,N_7289,N_9572);
or U12276 (N_12276,N_6347,N_6744);
xnor U12277 (N_12277,N_6388,N_7390);
and U12278 (N_12278,N_5983,N_8937);
and U12279 (N_12279,N_7639,N_7014);
nand U12280 (N_12280,N_8765,N_5278);
nand U12281 (N_12281,N_7844,N_8698);
nor U12282 (N_12282,N_7783,N_5520);
xor U12283 (N_12283,N_9422,N_8590);
nor U12284 (N_12284,N_8295,N_9197);
nor U12285 (N_12285,N_6371,N_8418);
xnor U12286 (N_12286,N_9181,N_9471);
xnor U12287 (N_12287,N_7867,N_5244);
and U12288 (N_12288,N_7780,N_7469);
nor U12289 (N_12289,N_9696,N_9566);
nand U12290 (N_12290,N_8415,N_9683);
or U12291 (N_12291,N_6386,N_8670);
or U12292 (N_12292,N_5465,N_8653);
nor U12293 (N_12293,N_7995,N_5493);
or U12294 (N_12294,N_5539,N_8664);
nand U12295 (N_12295,N_8342,N_6432);
and U12296 (N_12296,N_5977,N_7331);
and U12297 (N_12297,N_9590,N_8703);
xnor U12298 (N_12298,N_8665,N_9056);
nand U12299 (N_12299,N_9873,N_8547);
xnor U12300 (N_12300,N_8604,N_7159);
nand U12301 (N_12301,N_5695,N_7363);
nor U12302 (N_12302,N_9130,N_6324);
nor U12303 (N_12303,N_9485,N_6189);
nor U12304 (N_12304,N_9604,N_8853);
or U12305 (N_12305,N_6415,N_5547);
xor U12306 (N_12306,N_6433,N_5982);
xor U12307 (N_12307,N_9982,N_7138);
nor U12308 (N_12308,N_5692,N_5304);
and U12309 (N_12309,N_8954,N_9452);
xor U12310 (N_12310,N_7192,N_7240);
or U12311 (N_12311,N_7190,N_6015);
or U12312 (N_12312,N_9393,N_5201);
nor U12313 (N_12313,N_8379,N_9320);
or U12314 (N_12314,N_9194,N_9420);
nand U12315 (N_12315,N_5782,N_8029);
nand U12316 (N_12316,N_8101,N_8820);
nand U12317 (N_12317,N_8262,N_7158);
or U12318 (N_12318,N_6129,N_9924);
xnor U12319 (N_12319,N_7383,N_7031);
and U12320 (N_12320,N_8600,N_7846);
nand U12321 (N_12321,N_7434,N_7773);
or U12322 (N_12322,N_8013,N_8100);
nand U12323 (N_12323,N_7272,N_8739);
or U12324 (N_12324,N_6403,N_7806);
nand U12325 (N_12325,N_6310,N_6604);
nor U12326 (N_12326,N_7102,N_5831);
and U12327 (N_12327,N_5482,N_8130);
or U12328 (N_12328,N_9390,N_5016);
nand U12329 (N_12329,N_9154,N_8012);
nand U12330 (N_12330,N_7417,N_8243);
xnor U12331 (N_12331,N_8788,N_7097);
and U12332 (N_12332,N_9678,N_7260);
nand U12333 (N_12333,N_8321,N_8770);
nand U12334 (N_12334,N_6246,N_5668);
or U12335 (N_12335,N_7444,N_6870);
nor U12336 (N_12336,N_5861,N_7110);
xnor U12337 (N_12337,N_7093,N_7795);
nand U12338 (N_12338,N_9936,N_5589);
and U12339 (N_12339,N_5768,N_5508);
xnor U12340 (N_12340,N_7431,N_6373);
nor U12341 (N_12341,N_5997,N_5690);
or U12342 (N_12342,N_7265,N_5872);
xor U12343 (N_12343,N_9387,N_7226);
nand U12344 (N_12344,N_8713,N_6307);
and U12345 (N_12345,N_7340,N_9115);
nand U12346 (N_12346,N_8092,N_5317);
nor U12347 (N_12347,N_7678,N_6975);
nor U12348 (N_12348,N_6469,N_7314);
xor U12349 (N_12349,N_9209,N_8114);
nor U12350 (N_12350,N_5276,N_5688);
xor U12351 (N_12351,N_9618,N_8026);
and U12352 (N_12352,N_6102,N_6164);
nor U12353 (N_12353,N_7250,N_7834);
and U12354 (N_12354,N_9784,N_6597);
or U12355 (N_12355,N_7489,N_5793);
nand U12356 (N_12356,N_9489,N_9029);
xor U12357 (N_12357,N_8144,N_9846);
and U12358 (N_12358,N_9882,N_9469);
or U12359 (N_12359,N_6858,N_9522);
or U12360 (N_12360,N_7643,N_9357);
nand U12361 (N_12361,N_5035,N_7512);
nor U12362 (N_12362,N_8087,N_7180);
or U12363 (N_12363,N_8511,N_8888);
nand U12364 (N_12364,N_7225,N_8538);
xor U12365 (N_12365,N_7011,N_6626);
nor U12366 (N_12366,N_6965,N_9868);
nor U12367 (N_12367,N_6736,N_7895);
nand U12368 (N_12368,N_8337,N_7966);
and U12369 (N_12369,N_7580,N_6363);
xnor U12370 (N_12370,N_8583,N_6145);
and U12371 (N_12371,N_6972,N_5532);
xor U12372 (N_12372,N_9027,N_6992);
or U12373 (N_12373,N_5206,N_6365);
xor U12374 (N_12374,N_5358,N_9885);
nand U12375 (N_12375,N_8066,N_9681);
and U12376 (N_12376,N_6508,N_7570);
nor U12377 (N_12377,N_7023,N_6570);
xnor U12378 (N_12378,N_5285,N_9049);
or U12379 (N_12379,N_5290,N_5865);
or U12380 (N_12380,N_5473,N_8851);
and U12381 (N_12381,N_6568,N_8504);
nand U12382 (N_12382,N_8081,N_7270);
and U12383 (N_12383,N_5320,N_5540);
nor U12384 (N_12384,N_5901,N_5855);
or U12385 (N_12385,N_9680,N_7581);
and U12386 (N_12386,N_5857,N_7370);
or U12387 (N_12387,N_6390,N_5152);
nand U12388 (N_12388,N_6183,N_6306);
nand U12389 (N_12389,N_9976,N_6734);
nor U12390 (N_12390,N_9325,N_8734);
nand U12391 (N_12391,N_6203,N_5068);
xnor U12392 (N_12392,N_8400,N_7892);
and U12393 (N_12393,N_5458,N_7508);
nand U12394 (N_12394,N_8645,N_6221);
or U12395 (N_12395,N_5052,N_7243);
nand U12396 (N_12396,N_8957,N_6401);
nor U12397 (N_12397,N_7134,N_6523);
nor U12398 (N_12398,N_8250,N_9782);
nand U12399 (N_12399,N_5548,N_6360);
nand U12400 (N_12400,N_5081,N_9665);
nand U12401 (N_12401,N_7377,N_7408);
or U12402 (N_12402,N_9788,N_5616);
nor U12403 (N_12403,N_8207,N_7436);
nor U12404 (N_12404,N_8490,N_5204);
nor U12405 (N_12405,N_6113,N_6695);
and U12406 (N_12406,N_5509,N_8428);
nand U12407 (N_12407,N_5334,N_6356);
nor U12408 (N_12408,N_8669,N_6007);
xnor U12409 (N_12409,N_7355,N_5554);
and U12410 (N_12410,N_9613,N_9260);
or U12411 (N_12411,N_8694,N_9929);
nand U12412 (N_12412,N_7284,N_7277);
xnor U12413 (N_12413,N_5907,N_5992);
or U12414 (N_12414,N_6041,N_9506);
nor U12415 (N_12415,N_6016,N_8034);
xor U12416 (N_12416,N_7576,N_7025);
nor U12417 (N_12417,N_7177,N_7823);
nor U12418 (N_12418,N_6457,N_6426);
nor U12419 (N_12419,N_5645,N_8912);
or U12420 (N_12420,N_5087,N_7568);
xnor U12421 (N_12421,N_6288,N_7756);
nor U12422 (N_12422,N_7558,N_7538);
nor U12423 (N_12423,N_5751,N_9778);
and U12424 (N_12424,N_9035,N_6645);
nand U12425 (N_12425,N_5817,N_9054);
and U12426 (N_12426,N_7771,N_9904);
nand U12427 (N_12427,N_8265,N_6557);
xnor U12428 (N_12428,N_5398,N_6650);
nand U12429 (N_12429,N_6848,N_6413);
and U12430 (N_12430,N_8413,N_7543);
nand U12431 (N_12431,N_6333,N_5673);
or U12432 (N_12432,N_7605,N_8894);
and U12433 (N_12433,N_6331,N_5371);
nand U12434 (N_12434,N_6098,N_6051);
nor U12435 (N_12435,N_8785,N_7840);
nor U12436 (N_12436,N_7388,N_5485);
and U12437 (N_12437,N_8824,N_7373);
xnor U12438 (N_12438,N_8576,N_7968);
nor U12439 (N_12439,N_8530,N_9867);
or U12440 (N_12440,N_6280,N_9218);
nand U12441 (N_12441,N_5707,N_6271);
nor U12442 (N_12442,N_6000,N_9546);
or U12443 (N_12443,N_9468,N_7878);
nor U12444 (N_12444,N_5032,N_8640);
nand U12445 (N_12445,N_5853,N_5915);
nand U12446 (N_12446,N_9518,N_6655);
nand U12447 (N_12447,N_9574,N_9801);
nand U12448 (N_12448,N_8017,N_5519);
or U12449 (N_12449,N_9554,N_5619);
nor U12450 (N_12450,N_7865,N_5998);
xnor U12451 (N_12451,N_9228,N_5000);
and U12452 (N_12452,N_9980,N_5427);
and U12453 (N_12453,N_7239,N_9321);
xor U12454 (N_12454,N_8163,N_5441);
or U12455 (N_12455,N_6249,N_7644);
nand U12456 (N_12456,N_6191,N_7828);
xor U12457 (N_12457,N_8261,N_8464);
or U12458 (N_12458,N_7522,N_7762);
nor U12459 (N_12459,N_7513,N_9738);
and U12460 (N_12460,N_6998,N_5205);
or U12461 (N_12461,N_6808,N_8593);
nand U12462 (N_12462,N_9378,N_8833);
nor U12463 (N_12463,N_6531,N_8598);
nor U12464 (N_12464,N_8274,N_6472);
nand U12465 (N_12465,N_6435,N_9883);
xor U12466 (N_12466,N_7770,N_9200);
xor U12467 (N_12467,N_5777,N_5820);
or U12468 (N_12468,N_5772,N_9346);
or U12469 (N_12469,N_9131,N_5242);
and U12470 (N_12470,N_5895,N_6076);
and U12471 (N_12471,N_9481,N_9596);
or U12472 (N_12472,N_9808,N_7745);
nand U12473 (N_12473,N_9031,N_8334);
nor U12474 (N_12474,N_8375,N_6723);
or U12475 (N_12475,N_6983,N_9191);
and U12476 (N_12476,N_6217,N_6091);
nand U12477 (N_12477,N_9826,N_5177);
nand U12478 (N_12478,N_6588,N_8570);
nand U12479 (N_12479,N_9273,N_7310);
nand U12480 (N_12480,N_6710,N_8874);
nor U12481 (N_12481,N_7423,N_9657);
nor U12482 (N_12482,N_7142,N_6727);
nor U12483 (N_12483,N_8046,N_7212);
or U12484 (N_12484,N_6474,N_6665);
nand U12485 (N_12485,N_9243,N_7010);
or U12486 (N_12486,N_5498,N_9948);
nor U12487 (N_12487,N_8212,N_6996);
nand U12488 (N_12488,N_6913,N_8843);
nand U12489 (N_12489,N_5282,N_7285);
xnor U12490 (N_12490,N_9020,N_7156);
and U12491 (N_12491,N_7606,N_6444);
nor U12492 (N_12492,N_8685,N_8056);
nand U12493 (N_12493,N_9687,N_7254);
nor U12494 (N_12494,N_5331,N_5739);
xnor U12495 (N_12495,N_6392,N_5070);
nand U12496 (N_12496,N_5213,N_6298);
nand U12497 (N_12497,N_8361,N_9278);
and U12498 (N_12498,N_8781,N_5723);
nor U12499 (N_12499,N_6019,N_6224);
or U12500 (N_12500,N_6609,N_9153);
or U12501 (N_12501,N_5225,N_5511);
or U12502 (N_12502,N_8083,N_5236);
nor U12503 (N_12503,N_6946,N_9018);
xnor U12504 (N_12504,N_9658,N_5148);
xnor U12505 (N_12505,N_5115,N_6342);
nand U12506 (N_12506,N_8318,N_6932);
and U12507 (N_12507,N_8030,N_9308);
nor U12508 (N_12508,N_8597,N_8341);
or U12509 (N_12509,N_8884,N_9477);
or U12510 (N_12510,N_7698,N_5271);
nor U12511 (N_12511,N_6254,N_7517);
or U12512 (N_12512,N_9497,N_5533);
nand U12513 (N_12513,N_6360,N_8408);
or U12514 (N_12514,N_8494,N_9634);
or U12515 (N_12515,N_9229,N_9306);
nor U12516 (N_12516,N_8289,N_8029);
xnor U12517 (N_12517,N_7650,N_8770);
nor U12518 (N_12518,N_7653,N_5443);
nor U12519 (N_12519,N_9995,N_9259);
and U12520 (N_12520,N_7103,N_8095);
xnor U12521 (N_12521,N_7227,N_8133);
nor U12522 (N_12522,N_8473,N_8107);
xnor U12523 (N_12523,N_6616,N_9951);
nand U12524 (N_12524,N_6288,N_6955);
or U12525 (N_12525,N_9413,N_5874);
nor U12526 (N_12526,N_7360,N_5731);
and U12527 (N_12527,N_7060,N_8684);
and U12528 (N_12528,N_7452,N_8893);
nor U12529 (N_12529,N_7950,N_7170);
nor U12530 (N_12530,N_7016,N_7950);
nor U12531 (N_12531,N_5462,N_5204);
nor U12532 (N_12532,N_6122,N_7887);
nor U12533 (N_12533,N_5612,N_6904);
nand U12534 (N_12534,N_8811,N_9558);
nor U12535 (N_12535,N_8831,N_9630);
nand U12536 (N_12536,N_6433,N_5925);
nor U12537 (N_12537,N_5259,N_6309);
nand U12538 (N_12538,N_9129,N_8618);
or U12539 (N_12539,N_9244,N_5592);
and U12540 (N_12540,N_8595,N_6315);
nor U12541 (N_12541,N_6768,N_9950);
nand U12542 (N_12542,N_5646,N_5028);
or U12543 (N_12543,N_7896,N_5286);
or U12544 (N_12544,N_8493,N_8199);
xnor U12545 (N_12545,N_5200,N_5240);
xor U12546 (N_12546,N_5763,N_5202);
and U12547 (N_12547,N_7006,N_6641);
or U12548 (N_12548,N_8737,N_6679);
and U12549 (N_12549,N_6688,N_7181);
and U12550 (N_12550,N_9601,N_7192);
or U12551 (N_12551,N_7161,N_8734);
nand U12552 (N_12552,N_8201,N_7782);
xnor U12553 (N_12553,N_8168,N_8418);
or U12554 (N_12554,N_7565,N_9521);
and U12555 (N_12555,N_5692,N_9240);
xnor U12556 (N_12556,N_5941,N_8512);
or U12557 (N_12557,N_5568,N_8308);
and U12558 (N_12558,N_8853,N_8075);
xnor U12559 (N_12559,N_8002,N_8479);
nor U12560 (N_12560,N_5688,N_5018);
and U12561 (N_12561,N_8067,N_5477);
or U12562 (N_12562,N_5722,N_9663);
and U12563 (N_12563,N_8080,N_6311);
xnor U12564 (N_12564,N_7932,N_5705);
xnor U12565 (N_12565,N_9504,N_6626);
or U12566 (N_12566,N_6923,N_8807);
or U12567 (N_12567,N_8722,N_5876);
or U12568 (N_12568,N_7043,N_9722);
and U12569 (N_12569,N_6405,N_7648);
xnor U12570 (N_12570,N_8671,N_7990);
xnor U12571 (N_12571,N_8838,N_7249);
and U12572 (N_12572,N_6148,N_5815);
and U12573 (N_12573,N_7007,N_5170);
and U12574 (N_12574,N_9938,N_6678);
nand U12575 (N_12575,N_8327,N_7512);
or U12576 (N_12576,N_5321,N_6072);
nor U12577 (N_12577,N_5701,N_8524);
and U12578 (N_12578,N_9609,N_5355);
nor U12579 (N_12579,N_8114,N_7213);
xnor U12580 (N_12580,N_9990,N_5371);
nand U12581 (N_12581,N_5687,N_5241);
and U12582 (N_12582,N_7742,N_6094);
nor U12583 (N_12583,N_8915,N_7391);
nor U12584 (N_12584,N_6940,N_9424);
nor U12585 (N_12585,N_6672,N_9311);
and U12586 (N_12586,N_8519,N_9562);
and U12587 (N_12587,N_9534,N_9204);
and U12588 (N_12588,N_5983,N_5377);
xor U12589 (N_12589,N_8435,N_9532);
xnor U12590 (N_12590,N_5241,N_5540);
or U12591 (N_12591,N_9008,N_9010);
nand U12592 (N_12592,N_6182,N_8692);
xor U12593 (N_12593,N_6265,N_9683);
and U12594 (N_12594,N_8584,N_8554);
xor U12595 (N_12595,N_6272,N_9425);
nor U12596 (N_12596,N_5687,N_7049);
or U12597 (N_12597,N_8949,N_7300);
nor U12598 (N_12598,N_8993,N_6784);
xor U12599 (N_12599,N_8597,N_9589);
and U12600 (N_12600,N_8102,N_5108);
nand U12601 (N_12601,N_9390,N_9338);
xnor U12602 (N_12602,N_6783,N_9659);
xnor U12603 (N_12603,N_8960,N_9046);
or U12604 (N_12604,N_7831,N_9738);
or U12605 (N_12605,N_9717,N_7359);
xnor U12606 (N_12606,N_8292,N_7367);
and U12607 (N_12607,N_6601,N_8981);
xor U12608 (N_12608,N_8170,N_9115);
and U12609 (N_12609,N_5066,N_6624);
xnor U12610 (N_12610,N_6462,N_8833);
or U12611 (N_12611,N_9655,N_8434);
and U12612 (N_12612,N_9120,N_8304);
xnor U12613 (N_12613,N_5370,N_8059);
nor U12614 (N_12614,N_9663,N_6740);
xor U12615 (N_12615,N_5350,N_9319);
xnor U12616 (N_12616,N_6705,N_5547);
and U12617 (N_12617,N_9154,N_7312);
nand U12618 (N_12618,N_5894,N_9310);
and U12619 (N_12619,N_8455,N_9386);
nand U12620 (N_12620,N_7142,N_7245);
or U12621 (N_12621,N_7487,N_8760);
or U12622 (N_12622,N_8192,N_7134);
and U12623 (N_12623,N_6025,N_5579);
or U12624 (N_12624,N_9052,N_7263);
xnor U12625 (N_12625,N_9665,N_5516);
and U12626 (N_12626,N_8859,N_8224);
nor U12627 (N_12627,N_8938,N_8768);
and U12628 (N_12628,N_6645,N_7342);
nand U12629 (N_12629,N_9044,N_8531);
and U12630 (N_12630,N_5709,N_7906);
xor U12631 (N_12631,N_5792,N_5372);
and U12632 (N_12632,N_7405,N_5690);
nor U12633 (N_12633,N_5609,N_7253);
and U12634 (N_12634,N_9344,N_7950);
nand U12635 (N_12635,N_5110,N_8444);
xnor U12636 (N_12636,N_5015,N_6813);
xnor U12637 (N_12637,N_8403,N_8423);
or U12638 (N_12638,N_9440,N_6394);
and U12639 (N_12639,N_8168,N_5035);
or U12640 (N_12640,N_7824,N_6610);
nand U12641 (N_12641,N_6633,N_8468);
nand U12642 (N_12642,N_6131,N_5974);
nand U12643 (N_12643,N_9997,N_8487);
nand U12644 (N_12644,N_9421,N_6532);
and U12645 (N_12645,N_5447,N_9712);
xnor U12646 (N_12646,N_6343,N_8697);
nor U12647 (N_12647,N_6672,N_7599);
xnor U12648 (N_12648,N_8490,N_6566);
or U12649 (N_12649,N_6941,N_9684);
and U12650 (N_12650,N_6277,N_5893);
nor U12651 (N_12651,N_8406,N_6694);
or U12652 (N_12652,N_5091,N_9108);
and U12653 (N_12653,N_7998,N_5488);
xnor U12654 (N_12654,N_6860,N_7546);
or U12655 (N_12655,N_7195,N_8302);
xor U12656 (N_12656,N_9335,N_9276);
nor U12657 (N_12657,N_5313,N_5771);
xor U12658 (N_12658,N_7603,N_5806);
nor U12659 (N_12659,N_7625,N_8387);
and U12660 (N_12660,N_6586,N_6547);
or U12661 (N_12661,N_9741,N_8025);
or U12662 (N_12662,N_9642,N_5253);
and U12663 (N_12663,N_9392,N_7663);
nand U12664 (N_12664,N_8965,N_8929);
and U12665 (N_12665,N_6870,N_7164);
and U12666 (N_12666,N_8633,N_8557);
nor U12667 (N_12667,N_8339,N_9892);
xor U12668 (N_12668,N_7208,N_6478);
nor U12669 (N_12669,N_5715,N_8911);
nor U12670 (N_12670,N_6567,N_8513);
nand U12671 (N_12671,N_6236,N_6182);
and U12672 (N_12672,N_7416,N_9706);
nor U12673 (N_12673,N_5386,N_6296);
and U12674 (N_12674,N_8195,N_9059);
nor U12675 (N_12675,N_5770,N_8503);
xnor U12676 (N_12676,N_7225,N_8039);
or U12677 (N_12677,N_8641,N_5456);
and U12678 (N_12678,N_9473,N_5641);
xor U12679 (N_12679,N_7957,N_8338);
or U12680 (N_12680,N_9696,N_9564);
nor U12681 (N_12681,N_7787,N_9804);
or U12682 (N_12682,N_8865,N_8194);
and U12683 (N_12683,N_8072,N_6666);
or U12684 (N_12684,N_5991,N_6992);
or U12685 (N_12685,N_7820,N_6974);
nor U12686 (N_12686,N_6424,N_9912);
nand U12687 (N_12687,N_5932,N_9799);
and U12688 (N_12688,N_5795,N_5282);
nand U12689 (N_12689,N_6066,N_7841);
or U12690 (N_12690,N_7188,N_5138);
or U12691 (N_12691,N_5085,N_8967);
or U12692 (N_12692,N_6571,N_8962);
and U12693 (N_12693,N_7192,N_9715);
xor U12694 (N_12694,N_9454,N_8153);
or U12695 (N_12695,N_9320,N_6688);
and U12696 (N_12696,N_6621,N_7674);
xor U12697 (N_12697,N_6076,N_7910);
nand U12698 (N_12698,N_9873,N_5393);
or U12699 (N_12699,N_5612,N_7699);
and U12700 (N_12700,N_9683,N_7265);
nor U12701 (N_12701,N_6655,N_6552);
xnor U12702 (N_12702,N_9652,N_9867);
nand U12703 (N_12703,N_6610,N_5218);
and U12704 (N_12704,N_7485,N_5856);
nand U12705 (N_12705,N_9237,N_6666);
and U12706 (N_12706,N_7287,N_8984);
nor U12707 (N_12707,N_7731,N_6437);
xor U12708 (N_12708,N_9369,N_7926);
xor U12709 (N_12709,N_5756,N_6106);
and U12710 (N_12710,N_6641,N_6648);
and U12711 (N_12711,N_8960,N_9827);
xor U12712 (N_12712,N_9169,N_8868);
xnor U12713 (N_12713,N_9023,N_9410);
or U12714 (N_12714,N_5952,N_7851);
nand U12715 (N_12715,N_9304,N_7523);
xor U12716 (N_12716,N_9174,N_6732);
and U12717 (N_12717,N_8035,N_9547);
nand U12718 (N_12718,N_8533,N_9271);
or U12719 (N_12719,N_7990,N_6275);
or U12720 (N_12720,N_8888,N_5344);
nor U12721 (N_12721,N_8239,N_6717);
xor U12722 (N_12722,N_9778,N_8937);
and U12723 (N_12723,N_9448,N_5503);
xnor U12724 (N_12724,N_7021,N_6396);
or U12725 (N_12725,N_5899,N_5484);
or U12726 (N_12726,N_9096,N_7533);
and U12727 (N_12727,N_5506,N_8324);
and U12728 (N_12728,N_9880,N_7222);
or U12729 (N_12729,N_5675,N_7619);
and U12730 (N_12730,N_5819,N_6637);
and U12731 (N_12731,N_5948,N_5850);
nor U12732 (N_12732,N_9127,N_9853);
or U12733 (N_12733,N_9075,N_8284);
nand U12734 (N_12734,N_8405,N_8397);
or U12735 (N_12735,N_7655,N_9378);
nand U12736 (N_12736,N_5452,N_8401);
nand U12737 (N_12737,N_9718,N_6045);
and U12738 (N_12738,N_5950,N_7007);
and U12739 (N_12739,N_9717,N_9270);
nand U12740 (N_12740,N_6422,N_6313);
xnor U12741 (N_12741,N_6826,N_7006);
nor U12742 (N_12742,N_7569,N_9331);
nand U12743 (N_12743,N_7956,N_9981);
nand U12744 (N_12744,N_9587,N_7020);
xnor U12745 (N_12745,N_8829,N_8338);
xor U12746 (N_12746,N_5106,N_5909);
nor U12747 (N_12747,N_8105,N_5364);
nor U12748 (N_12748,N_6455,N_7687);
nand U12749 (N_12749,N_6781,N_8411);
and U12750 (N_12750,N_8533,N_9054);
or U12751 (N_12751,N_6480,N_9664);
and U12752 (N_12752,N_5137,N_9378);
nand U12753 (N_12753,N_9209,N_6124);
nand U12754 (N_12754,N_8612,N_6633);
xnor U12755 (N_12755,N_9906,N_8990);
nand U12756 (N_12756,N_6546,N_7402);
xor U12757 (N_12757,N_7125,N_9290);
xnor U12758 (N_12758,N_6439,N_6203);
or U12759 (N_12759,N_5726,N_9783);
nand U12760 (N_12760,N_7031,N_9245);
nand U12761 (N_12761,N_9509,N_9142);
or U12762 (N_12762,N_9244,N_7367);
and U12763 (N_12763,N_6930,N_7107);
xnor U12764 (N_12764,N_7328,N_5874);
xor U12765 (N_12765,N_7217,N_9363);
nor U12766 (N_12766,N_7156,N_9484);
nand U12767 (N_12767,N_5747,N_5697);
or U12768 (N_12768,N_7394,N_6389);
or U12769 (N_12769,N_9393,N_6152);
or U12770 (N_12770,N_5346,N_6797);
or U12771 (N_12771,N_8672,N_9883);
or U12772 (N_12772,N_7401,N_9609);
nor U12773 (N_12773,N_8038,N_5409);
nand U12774 (N_12774,N_9906,N_9872);
and U12775 (N_12775,N_7865,N_7263);
xor U12776 (N_12776,N_5750,N_9124);
or U12777 (N_12777,N_6934,N_5552);
xor U12778 (N_12778,N_5731,N_7548);
nor U12779 (N_12779,N_7185,N_9308);
nand U12780 (N_12780,N_5439,N_8569);
nor U12781 (N_12781,N_5563,N_9688);
nor U12782 (N_12782,N_6737,N_5397);
nor U12783 (N_12783,N_5048,N_5086);
or U12784 (N_12784,N_7363,N_5060);
xnor U12785 (N_12785,N_6316,N_9787);
nor U12786 (N_12786,N_7133,N_5682);
nor U12787 (N_12787,N_9167,N_8200);
nand U12788 (N_12788,N_6913,N_7822);
or U12789 (N_12789,N_9557,N_9083);
nor U12790 (N_12790,N_6004,N_8277);
nor U12791 (N_12791,N_6746,N_5165);
nor U12792 (N_12792,N_9302,N_8698);
and U12793 (N_12793,N_5312,N_5421);
or U12794 (N_12794,N_5266,N_8987);
nor U12795 (N_12795,N_8953,N_5501);
nor U12796 (N_12796,N_8765,N_5039);
nand U12797 (N_12797,N_9059,N_9775);
or U12798 (N_12798,N_5653,N_5783);
nor U12799 (N_12799,N_8719,N_6158);
nand U12800 (N_12800,N_9863,N_7878);
nor U12801 (N_12801,N_9803,N_6670);
and U12802 (N_12802,N_9128,N_5290);
and U12803 (N_12803,N_8132,N_7938);
nor U12804 (N_12804,N_6505,N_8965);
or U12805 (N_12805,N_9713,N_7333);
or U12806 (N_12806,N_9652,N_7282);
xnor U12807 (N_12807,N_6388,N_7324);
or U12808 (N_12808,N_5196,N_7021);
and U12809 (N_12809,N_5762,N_8220);
or U12810 (N_12810,N_6291,N_5205);
or U12811 (N_12811,N_8747,N_8245);
nand U12812 (N_12812,N_5640,N_6786);
nor U12813 (N_12813,N_6993,N_8033);
or U12814 (N_12814,N_6089,N_7129);
nand U12815 (N_12815,N_6518,N_8226);
nor U12816 (N_12816,N_6910,N_6189);
nand U12817 (N_12817,N_7394,N_7334);
and U12818 (N_12818,N_7751,N_5907);
nand U12819 (N_12819,N_6273,N_9212);
xor U12820 (N_12820,N_7779,N_5390);
or U12821 (N_12821,N_7235,N_9610);
and U12822 (N_12822,N_5052,N_6613);
nor U12823 (N_12823,N_7176,N_8209);
and U12824 (N_12824,N_9323,N_5833);
or U12825 (N_12825,N_5152,N_5435);
or U12826 (N_12826,N_5489,N_9982);
xor U12827 (N_12827,N_6444,N_9923);
or U12828 (N_12828,N_8157,N_6718);
xor U12829 (N_12829,N_5939,N_7992);
xnor U12830 (N_12830,N_8368,N_6014);
nor U12831 (N_12831,N_7840,N_9277);
and U12832 (N_12832,N_8812,N_8045);
and U12833 (N_12833,N_8037,N_7603);
or U12834 (N_12834,N_8024,N_9309);
nor U12835 (N_12835,N_6815,N_7515);
or U12836 (N_12836,N_8118,N_5849);
nor U12837 (N_12837,N_5144,N_5594);
xnor U12838 (N_12838,N_9214,N_8343);
nand U12839 (N_12839,N_8184,N_5851);
nor U12840 (N_12840,N_5632,N_6050);
nor U12841 (N_12841,N_5293,N_9385);
and U12842 (N_12842,N_5561,N_8926);
xor U12843 (N_12843,N_7368,N_9942);
or U12844 (N_12844,N_8778,N_8662);
nor U12845 (N_12845,N_7072,N_5198);
nand U12846 (N_12846,N_6775,N_5925);
nand U12847 (N_12847,N_6063,N_7125);
and U12848 (N_12848,N_9304,N_5963);
or U12849 (N_12849,N_9812,N_8543);
and U12850 (N_12850,N_7767,N_8263);
nand U12851 (N_12851,N_9882,N_8918);
or U12852 (N_12852,N_6515,N_9963);
nor U12853 (N_12853,N_7332,N_9872);
nand U12854 (N_12854,N_7579,N_7353);
nand U12855 (N_12855,N_7762,N_6595);
and U12856 (N_12856,N_9390,N_7601);
nor U12857 (N_12857,N_8443,N_8754);
nor U12858 (N_12858,N_6976,N_6397);
nand U12859 (N_12859,N_5932,N_5718);
xor U12860 (N_12860,N_8926,N_7699);
and U12861 (N_12861,N_9004,N_9882);
and U12862 (N_12862,N_9069,N_7129);
nor U12863 (N_12863,N_6888,N_5240);
nor U12864 (N_12864,N_7527,N_6862);
nor U12865 (N_12865,N_8608,N_5832);
nand U12866 (N_12866,N_5493,N_9454);
xnor U12867 (N_12867,N_5341,N_7629);
or U12868 (N_12868,N_8485,N_6898);
and U12869 (N_12869,N_7059,N_7051);
xor U12870 (N_12870,N_6759,N_6963);
nand U12871 (N_12871,N_9828,N_9847);
or U12872 (N_12872,N_7674,N_5852);
or U12873 (N_12873,N_9465,N_9817);
and U12874 (N_12874,N_6131,N_9990);
or U12875 (N_12875,N_9290,N_6258);
and U12876 (N_12876,N_5818,N_6943);
nor U12877 (N_12877,N_9125,N_8925);
or U12878 (N_12878,N_9321,N_8173);
xor U12879 (N_12879,N_6596,N_9686);
nand U12880 (N_12880,N_6785,N_7274);
and U12881 (N_12881,N_9612,N_8868);
and U12882 (N_12882,N_7158,N_6578);
nor U12883 (N_12883,N_5202,N_8307);
or U12884 (N_12884,N_5152,N_9832);
and U12885 (N_12885,N_5277,N_5858);
xnor U12886 (N_12886,N_5439,N_6158);
or U12887 (N_12887,N_8461,N_6687);
nor U12888 (N_12888,N_9081,N_7756);
or U12889 (N_12889,N_5375,N_6702);
nor U12890 (N_12890,N_8065,N_5005);
and U12891 (N_12891,N_8406,N_5346);
or U12892 (N_12892,N_7790,N_6490);
nand U12893 (N_12893,N_7045,N_9775);
or U12894 (N_12894,N_9753,N_5917);
or U12895 (N_12895,N_9563,N_7796);
and U12896 (N_12896,N_7010,N_5753);
nand U12897 (N_12897,N_5875,N_7374);
xor U12898 (N_12898,N_7513,N_8253);
or U12899 (N_12899,N_8412,N_6899);
or U12900 (N_12900,N_6811,N_5946);
or U12901 (N_12901,N_5477,N_5661);
nor U12902 (N_12902,N_9712,N_5464);
or U12903 (N_12903,N_8327,N_6307);
nor U12904 (N_12904,N_6208,N_8807);
or U12905 (N_12905,N_9132,N_8264);
nand U12906 (N_12906,N_5862,N_8436);
or U12907 (N_12907,N_5767,N_7874);
xnor U12908 (N_12908,N_8400,N_8543);
nand U12909 (N_12909,N_7695,N_7930);
and U12910 (N_12910,N_5733,N_6130);
and U12911 (N_12911,N_9692,N_9608);
and U12912 (N_12912,N_7453,N_7019);
or U12913 (N_12913,N_5803,N_7027);
and U12914 (N_12914,N_7575,N_8120);
or U12915 (N_12915,N_5499,N_5339);
and U12916 (N_12916,N_9258,N_6608);
xnor U12917 (N_12917,N_9075,N_7282);
nor U12918 (N_12918,N_8912,N_5816);
nor U12919 (N_12919,N_7034,N_9310);
xor U12920 (N_12920,N_6652,N_6932);
nor U12921 (N_12921,N_5955,N_7705);
or U12922 (N_12922,N_7221,N_6504);
or U12923 (N_12923,N_5538,N_8183);
and U12924 (N_12924,N_6811,N_6302);
nor U12925 (N_12925,N_8145,N_7764);
and U12926 (N_12926,N_5258,N_6047);
or U12927 (N_12927,N_9575,N_8353);
xnor U12928 (N_12928,N_8692,N_5412);
or U12929 (N_12929,N_6517,N_7594);
xnor U12930 (N_12930,N_7083,N_9488);
or U12931 (N_12931,N_7260,N_5088);
nand U12932 (N_12932,N_7533,N_6958);
nand U12933 (N_12933,N_5787,N_8958);
xor U12934 (N_12934,N_6572,N_5934);
nor U12935 (N_12935,N_6699,N_7952);
or U12936 (N_12936,N_9124,N_6515);
and U12937 (N_12937,N_6726,N_9727);
nor U12938 (N_12938,N_5667,N_5498);
nor U12939 (N_12939,N_9592,N_6120);
nand U12940 (N_12940,N_8181,N_7334);
nor U12941 (N_12941,N_7156,N_8826);
nor U12942 (N_12942,N_5421,N_5693);
xor U12943 (N_12943,N_5480,N_6274);
xnor U12944 (N_12944,N_5205,N_5668);
nand U12945 (N_12945,N_7541,N_5660);
nand U12946 (N_12946,N_7235,N_5472);
nand U12947 (N_12947,N_7033,N_5180);
or U12948 (N_12948,N_5269,N_8745);
nor U12949 (N_12949,N_6729,N_8244);
or U12950 (N_12950,N_7298,N_7325);
or U12951 (N_12951,N_9266,N_8147);
and U12952 (N_12952,N_7367,N_8329);
or U12953 (N_12953,N_5151,N_5866);
or U12954 (N_12954,N_7563,N_6149);
or U12955 (N_12955,N_9530,N_5666);
xor U12956 (N_12956,N_8546,N_7649);
and U12957 (N_12957,N_9421,N_6135);
or U12958 (N_12958,N_6284,N_6334);
xor U12959 (N_12959,N_8876,N_9303);
or U12960 (N_12960,N_7777,N_9839);
xnor U12961 (N_12961,N_8503,N_6335);
or U12962 (N_12962,N_9545,N_9426);
xnor U12963 (N_12963,N_5989,N_8361);
nor U12964 (N_12964,N_5808,N_5085);
nand U12965 (N_12965,N_8161,N_8622);
xor U12966 (N_12966,N_6594,N_5205);
and U12967 (N_12967,N_6398,N_9683);
nand U12968 (N_12968,N_8946,N_8646);
or U12969 (N_12969,N_9278,N_5632);
nand U12970 (N_12970,N_9621,N_6214);
and U12971 (N_12971,N_9973,N_7691);
and U12972 (N_12972,N_8572,N_9203);
xor U12973 (N_12973,N_6069,N_5927);
xnor U12974 (N_12974,N_6430,N_8646);
xnor U12975 (N_12975,N_5851,N_9137);
nor U12976 (N_12976,N_9282,N_5354);
or U12977 (N_12977,N_7546,N_8577);
nor U12978 (N_12978,N_8023,N_9535);
nor U12979 (N_12979,N_8273,N_8536);
xnor U12980 (N_12980,N_8382,N_9369);
and U12981 (N_12981,N_6840,N_8890);
nor U12982 (N_12982,N_8561,N_5777);
nor U12983 (N_12983,N_9154,N_9854);
nand U12984 (N_12984,N_7325,N_5244);
xor U12985 (N_12985,N_9600,N_8041);
or U12986 (N_12986,N_7223,N_7236);
xor U12987 (N_12987,N_9208,N_9456);
nor U12988 (N_12988,N_5920,N_6260);
nor U12989 (N_12989,N_6621,N_5182);
and U12990 (N_12990,N_6489,N_5443);
xor U12991 (N_12991,N_5867,N_9199);
or U12992 (N_12992,N_8727,N_7110);
xnor U12993 (N_12993,N_8670,N_5976);
nand U12994 (N_12994,N_7219,N_5431);
xor U12995 (N_12995,N_6516,N_9618);
nor U12996 (N_12996,N_8581,N_5966);
xnor U12997 (N_12997,N_9484,N_5844);
nand U12998 (N_12998,N_9055,N_7394);
xor U12999 (N_12999,N_6967,N_7916);
xor U13000 (N_13000,N_6464,N_7961);
xnor U13001 (N_13001,N_5716,N_8741);
nor U13002 (N_13002,N_5686,N_6870);
or U13003 (N_13003,N_6365,N_8331);
nor U13004 (N_13004,N_7787,N_8592);
nand U13005 (N_13005,N_9685,N_5306);
or U13006 (N_13006,N_7371,N_7409);
or U13007 (N_13007,N_6462,N_6786);
nand U13008 (N_13008,N_8720,N_5907);
or U13009 (N_13009,N_6477,N_9191);
xor U13010 (N_13010,N_6829,N_9724);
nand U13011 (N_13011,N_5165,N_9515);
nand U13012 (N_13012,N_8737,N_9374);
nor U13013 (N_13013,N_5803,N_6940);
nand U13014 (N_13014,N_9601,N_7910);
and U13015 (N_13015,N_7849,N_5641);
and U13016 (N_13016,N_8044,N_8251);
xnor U13017 (N_13017,N_8958,N_5294);
nor U13018 (N_13018,N_6225,N_7941);
nand U13019 (N_13019,N_5960,N_9725);
and U13020 (N_13020,N_5892,N_5882);
nand U13021 (N_13021,N_7274,N_5025);
nand U13022 (N_13022,N_7941,N_8779);
or U13023 (N_13023,N_5181,N_8360);
nand U13024 (N_13024,N_9074,N_8641);
nand U13025 (N_13025,N_7793,N_5435);
nor U13026 (N_13026,N_6098,N_9621);
and U13027 (N_13027,N_7327,N_6160);
xor U13028 (N_13028,N_9775,N_5465);
xnor U13029 (N_13029,N_7632,N_6105);
and U13030 (N_13030,N_9713,N_7411);
and U13031 (N_13031,N_6440,N_8717);
xor U13032 (N_13032,N_9914,N_9540);
nand U13033 (N_13033,N_7611,N_8664);
nor U13034 (N_13034,N_5026,N_7181);
nand U13035 (N_13035,N_6086,N_5881);
and U13036 (N_13036,N_6710,N_6184);
nand U13037 (N_13037,N_6526,N_6646);
nand U13038 (N_13038,N_6771,N_6563);
nand U13039 (N_13039,N_5688,N_7435);
xor U13040 (N_13040,N_8543,N_9231);
and U13041 (N_13041,N_6951,N_9057);
nor U13042 (N_13042,N_9130,N_5606);
and U13043 (N_13043,N_5548,N_5894);
nor U13044 (N_13044,N_8476,N_8938);
nand U13045 (N_13045,N_6066,N_7563);
or U13046 (N_13046,N_6119,N_8134);
and U13047 (N_13047,N_5929,N_8364);
nor U13048 (N_13048,N_9081,N_7519);
or U13049 (N_13049,N_9000,N_6975);
and U13050 (N_13050,N_7408,N_9367);
nand U13051 (N_13051,N_6779,N_9463);
xor U13052 (N_13052,N_7417,N_8371);
nor U13053 (N_13053,N_6153,N_8491);
nand U13054 (N_13054,N_6277,N_8861);
or U13055 (N_13055,N_9731,N_8014);
xor U13056 (N_13056,N_5622,N_5462);
or U13057 (N_13057,N_7237,N_9946);
and U13058 (N_13058,N_5858,N_6135);
xnor U13059 (N_13059,N_8745,N_5021);
and U13060 (N_13060,N_5193,N_8723);
nor U13061 (N_13061,N_7351,N_8789);
xor U13062 (N_13062,N_9789,N_7498);
nand U13063 (N_13063,N_7802,N_6169);
xor U13064 (N_13064,N_5413,N_9559);
xnor U13065 (N_13065,N_9719,N_9546);
and U13066 (N_13066,N_6570,N_5735);
nor U13067 (N_13067,N_6754,N_5486);
and U13068 (N_13068,N_6525,N_8789);
or U13069 (N_13069,N_8970,N_9388);
nor U13070 (N_13070,N_9759,N_9178);
nor U13071 (N_13071,N_6417,N_9425);
nor U13072 (N_13072,N_6595,N_6043);
or U13073 (N_13073,N_8706,N_6478);
nor U13074 (N_13074,N_7948,N_8976);
or U13075 (N_13075,N_5002,N_7008);
xor U13076 (N_13076,N_8910,N_6591);
or U13077 (N_13077,N_7872,N_8983);
and U13078 (N_13078,N_9442,N_8085);
nand U13079 (N_13079,N_8810,N_9787);
nand U13080 (N_13080,N_9477,N_7812);
or U13081 (N_13081,N_5620,N_9013);
or U13082 (N_13082,N_7615,N_8340);
nand U13083 (N_13083,N_8788,N_8532);
nor U13084 (N_13084,N_7441,N_5500);
nand U13085 (N_13085,N_9789,N_9213);
xor U13086 (N_13086,N_9502,N_6902);
and U13087 (N_13087,N_8987,N_7390);
or U13088 (N_13088,N_9821,N_8596);
and U13089 (N_13089,N_6688,N_7484);
xor U13090 (N_13090,N_9141,N_8362);
and U13091 (N_13091,N_7861,N_9388);
nand U13092 (N_13092,N_7904,N_6778);
nor U13093 (N_13093,N_8640,N_6162);
nor U13094 (N_13094,N_5588,N_5973);
xnor U13095 (N_13095,N_9329,N_8990);
xnor U13096 (N_13096,N_5399,N_6744);
nor U13097 (N_13097,N_7630,N_5694);
xnor U13098 (N_13098,N_9422,N_5721);
or U13099 (N_13099,N_5629,N_5526);
and U13100 (N_13100,N_9140,N_9908);
and U13101 (N_13101,N_6151,N_9982);
and U13102 (N_13102,N_7793,N_5233);
xor U13103 (N_13103,N_5521,N_7395);
nand U13104 (N_13104,N_7069,N_8074);
and U13105 (N_13105,N_5588,N_7950);
nand U13106 (N_13106,N_8834,N_8689);
or U13107 (N_13107,N_5369,N_6370);
xnor U13108 (N_13108,N_5869,N_6753);
nor U13109 (N_13109,N_6521,N_6729);
and U13110 (N_13110,N_7998,N_9677);
nand U13111 (N_13111,N_5837,N_7147);
and U13112 (N_13112,N_6559,N_9452);
nor U13113 (N_13113,N_6622,N_7467);
nor U13114 (N_13114,N_6810,N_8874);
or U13115 (N_13115,N_7876,N_6750);
nand U13116 (N_13116,N_7511,N_9877);
or U13117 (N_13117,N_6915,N_8542);
or U13118 (N_13118,N_8250,N_7715);
xnor U13119 (N_13119,N_5643,N_9351);
xor U13120 (N_13120,N_8238,N_9605);
nor U13121 (N_13121,N_8278,N_5063);
nand U13122 (N_13122,N_7789,N_8365);
nand U13123 (N_13123,N_5101,N_9913);
nand U13124 (N_13124,N_8094,N_5884);
or U13125 (N_13125,N_8141,N_8188);
and U13126 (N_13126,N_7132,N_8747);
and U13127 (N_13127,N_7944,N_9806);
or U13128 (N_13128,N_7495,N_6382);
nand U13129 (N_13129,N_5074,N_8175);
or U13130 (N_13130,N_8915,N_8399);
xor U13131 (N_13131,N_6244,N_7813);
xor U13132 (N_13132,N_9346,N_9806);
or U13133 (N_13133,N_6941,N_5056);
nand U13134 (N_13134,N_7107,N_6100);
or U13135 (N_13135,N_7521,N_6490);
xor U13136 (N_13136,N_8883,N_5798);
nor U13137 (N_13137,N_6936,N_8143);
xnor U13138 (N_13138,N_8638,N_9762);
and U13139 (N_13139,N_5577,N_5709);
or U13140 (N_13140,N_5326,N_5536);
nor U13141 (N_13141,N_8025,N_9970);
and U13142 (N_13142,N_5840,N_9533);
or U13143 (N_13143,N_5500,N_9489);
xnor U13144 (N_13144,N_9244,N_5234);
or U13145 (N_13145,N_9719,N_7598);
and U13146 (N_13146,N_7237,N_5372);
nor U13147 (N_13147,N_5199,N_5443);
nor U13148 (N_13148,N_7067,N_5280);
xnor U13149 (N_13149,N_9045,N_7518);
or U13150 (N_13150,N_9790,N_9623);
nor U13151 (N_13151,N_8199,N_8658);
or U13152 (N_13152,N_6145,N_9739);
nor U13153 (N_13153,N_8097,N_9777);
nor U13154 (N_13154,N_6809,N_5734);
nand U13155 (N_13155,N_8268,N_6259);
or U13156 (N_13156,N_6339,N_7168);
nor U13157 (N_13157,N_5052,N_8140);
nand U13158 (N_13158,N_9450,N_7910);
and U13159 (N_13159,N_9235,N_7752);
nor U13160 (N_13160,N_8441,N_5944);
xnor U13161 (N_13161,N_8614,N_5990);
nand U13162 (N_13162,N_8584,N_9713);
nand U13163 (N_13163,N_9340,N_8541);
xor U13164 (N_13164,N_5930,N_8793);
or U13165 (N_13165,N_7969,N_8305);
xor U13166 (N_13166,N_8933,N_9686);
nor U13167 (N_13167,N_6154,N_6598);
and U13168 (N_13168,N_8104,N_6123);
xnor U13169 (N_13169,N_9345,N_6348);
nand U13170 (N_13170,N_6890,N_7487);
nor U13171 (N_13171,N_9498,N_6828);
xnor U13172 (N_13172,N_9882,N_9132);
nand U13173 (N_13173,N_8920,N_8318);
and U13174 (N_13174,N_9601,N_9790);
or U13175 (N_13175,N_9680,N_8113);
nor U13176 (N_13176,N_5586,N_9205);
or U13177 (N_13177,N_9044,N_6619);
nor U13178 (N_13178,N_6128,N_7512);
nand U13179 (N_13179,N_8345,N_8699);
xnor U13180 (N_13180,N_7511,N_7233);
and U13181 (N_13181,N_9564,N_8153);
or U13182 (N_13182,N_5681,N_5607);
nand U13183 (N_13183,N_8939,N_5401);
nand U13184 (N_13184,N_6747,N_6378);
and U13185 (N_13185,N_8953,N_5201);
and U13186 (N_13186,N_8108,N_8789);
and U13187 (N_13187,N_6368,N_7164);
nand U13188 (N_13188,N_9956,N_9650);
or U13189 (N_13189,N_7383,N_5628);
or U13190 (N_13190,N_5322,N_5325);
xnor U13191 (N_13191,N_5114,N_5299);
xor U13192 (N_13192,N_8167,N_7817);
nand U13193 (N_13193,N_5083,N_5062);
nand U13194 (N_13194,N_8778,N_6563);
and U13195 (N_13195,N_8201,N_9856);
nand U13196 (N_13196,N_7158,N_9724);
or U13197 (N_13197,N_9474,N_5039);
nand U13198 (N_13198,N_6932,N_9352);
xnor U13199 (N_13199,N_7205,N_9727);
xnor U13200 (N_13200,N_9406,N_5601);
and U13201 (N_13201,N_8498,N_8387);
nor U13202 (N_13202,N_5252,N_8760);
nor U13203 (N_13203,N_8104,N_8326);
or U13204 (N_13204,N_7187,N_8574);
xnor U13205 (N_13205,N_9798,N_6179);
nand U13206 (N_13206,N_8692,N_9897);
xor U13207 (N_13207,N_5507,N_7901);
and U13208 (N_13208,N_6155,N_9316);
xnor U13209 (N_13209,N_7616,N_7471);
or U13210 (N_13210,N_6099,N_7482);
or U13211 (N_13211,N_9289,N_6753);
xor U13212 (N_13212,N_7026,N_8649);
nor U13213 (N_13213,N_8055,N_5533);
or U13214 (N_13214,N_7634,N_6399);
and U13215 (N_13215,N_6812,N_8590);
and U13216 (N_13216,N_8235,N_5254);
nor U13217 (N_13217,N_9490,N_6398);
nand U13218 (N_13218,N_5264,N_7045);
and U13219 (N_13219,N_6178,N_5722);
nor U13220 (N_13220,N_9077,N_8247);
or U13221 (N_13221,N_8937,N_6910);
nand U13222 (N_13222,N_9848,N_7048);
nand U13223 (N_13223,N_6460,N_5779);
nand U13224 (N_13224,N_7243,N_8750);
nand U13225 (N_13225,N_7448,N_8531);
and U13226 (N_13226,N_8410,N_7147);
and U13227 (N_13227,N_7302,N_9796);
xor U13228 (N_13228,N_9805,N_6338);
xor U13229 (N_13229,N_8277,N_5784);
xor U13230 (N_13230,N_7925,N_6410);
xnor U13231 (N_13231,N_9288,N_7563);
and U13232 (N_13232,N_8273,N_9221);
xnor U13233 (N_13233,N_6325,N_7154);
nor U13234 (N_13234,N_9037,N_5913);
and U13235 (N_13235,N_7770,N_8649);
and U13236 (N_13236,N_8127,N_8039);
nand U13237 (N_13237,N_5289,N_6601);
xor U13238 (N_13238,N_5278,N_7737);
nand U13239 (N_13239,N_8529,N_9960);
nor U13240 (N_13240,N_8012,N_7252);
and U13241 (N_13241,N_6190,N_8765);
nand U13242 (N_13242,N_9764,N_5471);
nand U13243 (N_13243,N_5598,N_9425);
nand U13244 (N_13244,N_6286,N_9364);
nand U13245 (N_13245,N_7300,N_8025);
xor U13246 (N_13246,N_6336,N_6295);
xnor U13247 (N_13247,N_5570,N_5999);
xor U13248 (N_13248,N_9144,N_6509);
or U13249 (N_13249,N_5643,N_6069);
nor U13250 (N_13250,N_8424,N_7521);
or U13251 (N_13251,N_5166,N_5159);
or U13252 (N_13252,N_5455,N_8704);
or U13253 (N_13253,N_7569,N_7180);
and U13254 (N_13254,N_9844,N_8426);
nor U13255 (N_13255,N_6067,N_8709);
xnor U13256 (N_13256,N_7088,N_6359);
nand U13257 (N_13257,N_5867,N_9803);
nor U13258 (N_13258,N_6338,N_8467);
xor U13259 (N_13259,N_6644,N_9654);
nand U13260 (N_13260,N_8704,N_9785);
nand U13261 (N_13261,N_7527,N_6133);
nor U13262 (N_13262,N_9837,N_7688);
nand U13263 (N_13263,N_6684,N_5891);
xor U13264 (N_13264,N_8842,N_6598);
xor U13265 (N_13265,N_7959,N_9889);
nor U13266 (N_13266,N_6121,N_7352);
nand U13267 (N_13267,N_8108,N_9263);
or U13268 (N_13268,N_8573,N_8823);
and U13269 (N_13269,N_9506,N_8132);
xnor U13270 (N_13270,N_7059,N_5870);
xor U13271 (N_13271,N_9590,N_9458);
xnor U13272 (N_13272,N_6461,N_5922);
nor U13273 (N_13273,N_7315,N_8660);
xor U13274 (N_13274,N_8357,N_7383);
nand U13275 (N_13275,N_6287,N_6724);
nor U13276 (N_13276,N_6766,N_6219);
or U13277 (N_13277,N_9672,N_9806);
or U13278 (N_13278,N_6382,N_7237);
nand U13279 (N_13279,N_7115,N_7060);
nand U13280 (N_13280,N_8494,N_6254);
and U13281 (N_13281,N_6525,N_7323);
or U13282 (N_13282,N_7218,N_9790);
xnor U13283 (N_13283,N_7712,N_6813);
and U13284 (N_13284,N_9715,N_9931);
and U13285 (N_13285,N_6414,N_5887);
or U13286 (N_13286,N_7260,N_8622);
xor U13287 (N_13287,N_7840,N_7237);
or U13288 (N_13288,N_7039,N_7044);
nor U13289 (N_13289,N_9367,N_6057);
nor U13290 (N_13290,N_6734,N_6472);
or U13291 (N_13291,N_8730,N_9329);
and U13292 (N_13292,N_7901,N_7603);
or U13293 (N_13293,N_7203,N_7674);
nand U13294 (N_13294,N_9311,N_5060);
and U13295 (N_13295,N_6245,N_6010);
nand U13296 (N_13296,N_8927,N_5192);
nand U13297 (N_13297,N_8495,N_6331);
xnor U13298 (N_13298,N_5201,N_5621);
nor U13299 (N_13299,N_6939,N_7845);
or U13300 (N_13300,N_8363,N_9855);
nor U13301 (N_13301,N_8429,N_6266);
or U13302 (N_13302,N_7030,N_9070);
and U13303 (N_13303,N_5243,N_8437);
nand U13304 (N_13304,N_6178,N_8936);
nand U13305 (N_13305,N_8055,N_9566);
and U13306 (N_13306,N_5886,N_6237);
xnor U13307 (N_13307,N_5096,N_7603);
xor U13308 (N_13308,N_6803,N_8253);
xor U13309 (N_13309,N_7607,N_5517);
nand U13310 (N_13310,N_7389,N_7739);
nor U13311 (N_13311,N_8561,N_7594);
or U13312 (N_13312,N_7988,N_7935);
xor U13313 (N_13313,N_7661,N_6213);
xnor U13314 (N_13314,N_8795,N_9978);
nand U13315 (N_13315,N_8329,N_5107);
and U13316 (N_13316,N_9968,N_5585);
or U13317 (N_13317,N_6367,N_6799);
xnor U13318 (N_13318,N_9809,N_7570);
xor U13319 (N_13319,N_5899,N_6382);
or U13320 (N_13320,N_7342,N_9699);
and U13321 (N_13321,N_6914,N_8678);
nor U13322 (N_13322,N_9518,N_5969);
xor U13323 (N_13323,N_5198,N_7051);
nand U13324 (N_13324,N_5338,N_6332);
nor U13325 (N_13325,N_6187,N_8004);
nand U13326 (N_13326,N_9577,N_6677);
xnor U13327 (N_13327,N_7335,N_7732);
or U13328 (N_13328,N_5044,N_9508);
xor U13329 (N_13329,N_9908,N_9145);
nor U13330 (N_13330,N_9199,N_7469);
or U13331 (N_13331,N_7993,N_5821);
nor U13332 (N_13332,N_5122,N_9560);
or U13333 (N_13333,N_9218,N_7170);
nand U13334 (N_13334,N_5483,N_9027);
or U13335 (N_13335,N_7348,N_6491);
xor U13336 (N_13336,N_7514,N_8608);
nand U13337 (N_13337,N_8054,N_5263);
xnor U13338 (N_13338,N_9705,N_7718);
xor U13339 (N_13339,N_6497,N_9082);
nor U13340 (N_13340,N_7324,N_5188);
and U13341 (N_13341,N_6850,N_8995);
xor U13342 (N_13342,N_9452,N_8729);
nor U13343 (N_13343,N_7157,N_8198);
or U13344 (N_13344,N_6509,N_9350);
or U13345 (N_13345,N_7447,N_6472);
xor U13346 (N_13346,N_9974,N_7092);
or U13347 (N_13347,N_8925,N_7301);
and U13348 (N_13348,N_6448,N_8950);
nand U13349 (N_13349,N_5697,N_9147);
nand U13350 (N_13350,N_5025,N_5988);
nor U13351 (N_13351,N_5790,N_5687);
or U13352 (N_13352,N_6463,N_9391);
or U13353 (N_13353,N_6452,N_7438);
and U13354 (N_13354,N_5574,N_9739);
or U13355 (N_13355,N_5273,N_5632);
or U13356 (N_13356,N_8228,N_5819);
and U13357 (N_13357,N_7393,N_8109);
or U13358 (N_13358,N_7052,N_8649);
xor U13359 (N_13359,N_7636,N_9193);
nor U13360 (N_13360,N_9858,N_5443);
nor U13361 (N_13361,N_8018,N_9837);
xor U13362 (N_13362,N_8892,N_9840);
nand U13363 (N_13363,N_5973,N_7108);
and U13364 (N_13364,N_9806,N_9475);
nand U13365 (N_13365,N_7478,N_7282);
nand U13366 (N_13366,N_9083,N_6501);
and U13367 (N_13367,N_5088,N_9933);
and U13368 (N_13368,N_9632,N_5291);
xor U13369 (N_13369,N_9561,N_9258);
xnor U13370 (N_13370,N_6159,N_7056);
nor U13371 (N_13371,N_8714,N_8418);
or U13372 (N_13372,N_7270,N_8978);
or U13373 (N_13373,N_6609,N_5228);
and U13374 (N_13374,N_8036,N_9137);
or U13375 (N_13375,N_6110,N_5331);
and U13376 (N_13376,N_6927,N_6525);
nand U13377 (N_13377,N_7183,N_8473);
xor U13378 (N_13378,N_9624,N_7350);
and U13379 (N_13379,N_7444,N_6209);
or U13380 (N_13380,N_8090,N_8585);
nand U13381 (N_13381,N_5540,N_5104);
nand U13382 (N_13382,N_9070,N_7338);
and U13383 (N_13383,N_9179,N_7732);
nor U13384 (N_13384,N_7344,N_8328);
nor U13385 (N_13385,N_8045,N_5524);
or U13386 (N_13386,N_7566,N_7326);
xor U13387 (N_13387,N_9617,N_9994);
nand U13388 (N_13388,N_7419,N_5190);
nand U13389 (N_13389,N_5984,N_8853);
nand U13390 (N_13390,N_9964,N_5706);
nor U13391 (N_13391,N_5654,N_7174);
nor U13392 (N_13392,N_9207,N_7064);
nand U13393 (N_13393,N_9854,N_8803);
and U13394 (N_13394,N_6192,N_8721);
xor U13395 (N_13395,N_7149,N_5612);
xor U13396 (N_13396,N_5086,N_7857);
xnor U13397 (N_13397,N_9041,N_9847);
nor U13398 (N_13398,N_5196,N_7359);
and U13399 (N_13399,N_8401,N_5676);
xnor U13400 (N_13400,N_9329,N_6711);
nor U13401 (N_13401,N_9211,N_8286);
or U13402 (N_13402,N_9358,N_6692);
xor U13403 (N_13403,N_8893,N_8150);
xor U13404 (N_13404,N_7578,N_6654);
or U13405 (N_13405,N_6885,N_6193);
or U13406 (N_13406,N_9862,N_6699);
nor U13407 (N_13407,N_5358,N_9976);
nand U13408 (N_13408,N_6432,N_9163);
xor U13409 (N_13409,N_7144,N_8304);
nor U13410 (N_13410,N_7165,N_6583);
and U13411 (N_13411,N_6731,N_5703);
nor U13412 (N_13412,N_7332,N_6582);
or U13413 (N_13413,N_8317,N_7981);
nor U13414 (N_13414,N_7140,N_5750);
nor U13415 (N_13415,N_7879,N_6973);
nor U13416 (N_13416,N_8576,N_7644);
nand U13417 (N_13417,N_5989,N_8013);
nor U13418 (N_13418,N_7774,N_9585);
xor U13419 (N_13419,N_7904,N_8779);
xor U13420 (N_13420,N_8321,N_6702);
and U13421 (N_13421,N_5229,N_7128);
xnor U13422 (N_13422,N_6243,N_9078);
nor U13423 (N_13423,N_6299,N_7562);
xor U13424 (N_13424,N_8587,N_8432);
nor U13425 (N_13425,N_5932,N_5653);
nor U13426 (N_13426,N_6321,N_8552);
nor U13427 (N_13427,N_7337,N_6722);
or U13428 (N_13428,N_8680,N_8371);
nor U13429 (N_13429,N_6241,N_8671);
xnor U13430 (N_13430,N_9416,N_9885);
nand U13431 (N_13431,N_6898,N_6785);
and U13432 (N_13432,N_5410,N_8701);
nor U13433 (N_13433,N_6883,N_6312);
or U13434 (N_13434,N_7297,N_9305);
nor U13435 (N_13435,N_6550,N_8675);
nand U13436 (N_13436,N_5298,N_9450);
xnor U13437 (N_13437,N_5580,N_8228);
nand U13438 (N_13438,N_6560,N_8520);
xor U13439 (N_13439,N_9629,N_6463);
xor U13440 (N_13440,N_6285,N_9460);
and U13441 (N_13441,N_9403,N_9790);
nor U13442 (N_13442,N_9741,N_7183);
xor U13443 (N_13443,N_9201,N_5803);
nand U13444 (N_13444,N_5824,N_8321);
nor U13445 (N_13445,N_7480,N_9443);
nor U13446 (N_13446,N_5203,N_6484);
or U13447 (N_13447,N_5617,N_7797);
or U13448 (N_13448,N_9988,N_6483);
and U13449 (N_13449,N_6094,N_9028);
xor U13450 (N_13450,N_7561,N_9413);
nand U13451 (N_13451,N_9723,N_8265);
or U13452 (N_13452,N_6097,N_6344);
xor U13453 (N_13453,N_9116,N_9631);
nor U13454 (N_13454,N_9224,N_6546);
xnor U13455 (N_13455,N_9406,N_6953);
xnor U13456 (N_13456,N_6796,N_9790);
nor U13457 (N_13457,N_9968,N_9419);
or U13458 (N_13458,N_9724,N_5596);
and U13459 (N_13459,N_9575,N_8137);
and U13460 (N_13460,N_7084,N_7715);
nor U13461 (N_13461,N_9016,N_5504);
and U13462 (N_13462,N_9751,N_5335);
nor U13463 (N_13463,N_9500,N_7892);
nand U13464 (N_13464,N_6039,N_9759);
xnor U13465 (N_13465,N_7755,N_6524);
xnor U13466 (N_13466,N_8431,N_5960);
and U13467 (N_13467,N_6824,N_5836);
nand U13468 (N_13468,N_8524,N_6860);
nand U13469 (N_13469,N_5133,N_6918);
or U13470 (N_13470,N_6543,N_7873);
xor U13471 (N_13471,N_9752,N_7165);
or U13472 (N_13472,N_5185,N_9920);
nor U13473 (N_13473,N_6369,N_8376);
or U13474 (N_13474,N_8453,N_6410);
and U13475 (N_13475,N_6682,N_5868);
nor U13476 (N_13476,N_7437,N_9388);
or U13477 (N_13477,N_7924,N_6553);
nor U13478 (N_13478,N_8396,N_9410);
nand U13479 (N_13479,N_8466,N_7013);
xor U13480 (N_13480,N_8347,N_6043);
or U13481 (N_13481,N_9201,N_5496);
nand U13482 (N_13482,N_6735,N_9009);
nor U13483 (N_13483,N_6900,N_9180);
or U13484 (N_13484,N_6615,N_7783);
and U13485 (N_13485,N_8099,N_8450);
nand U13486 (N_13486,N_8659,N_9595);
or U13487 (N_13487,N_5256,N_8330);
and U13488 (N_13488,N_5718,N_5073);
xnor U13489 (N_13489,N_5424,N_8326);
xnor U13490 (N_13490,N_5878,N_5548);
and U13491 (N_13491,N_5590,N_5960);
xor U13492 (N_13492,N_9286,N_7905);
or U13493 (N_13493,N_5787,N_9302);
nand U13494 (N_13494,N_9929,N_7675);
and U13495 (N_13495,N_6960,N_5617);
nand U13496 (N_13496,N_8395,N_9913);
nand U13497 (N_13497,N_5095,N_5929);
nand U13498 (N_13498,N_6588,N_7465);
nor U13499 (N_13499,N_5998,N_7101);
and U13500 (N_13500,N_7194,N_7073);
nor U13501 (N_13501,N_8654,N_7630);
nor U13502 (N_13502,N_6706,N_7993);
or U13503 (N_13503,N_8847,N_7328);
and U13504 (N_13504,N_5304,N_6811);
nand U13505 (N_13505,N_9137,N_9542);
nand U13506 (N_13506,N_8095,N_5887);
nor U13507 (N_13507,N_9759,N_9547);
nand U13508 (N_13508,N_7055,N_9718);
and U13509 (N_13509,N_7057,N_7835);
and U13510 (N_13510,N_6252,N_6251);
nor U13511 (N_13511,N_8203,N_6642);
or U13512 (N_13512,N_7712,N_9824);
nor U13513 (N_13513,N_9521,N_7800);
or U13514 (N_13514,N_8707,N_5810);
nand U13515 (N_13515,N_5423,N_6725);
and U13516 (N_13516,N_5560,N_9133);
nand U13517 (N_13517,N_7313,N_9138);
and U13518 (N_13518,N_8526,N_7169);
nand U13519 (N_13519,N_7250,N_8361);
nand U13520 (N_13520,N_9884,N_6033);
or U13521 (N_13521,N_6929,N_5228);
xnor U13522 (N_13522,N_9311,N_9678);
nand U13523 (N_13523,N_8118,N_7272);
or U13524 (N_13524,N_8407,N_6183);
nor U13525 (N_13525,N_9257,N_6951);
xor U13526 (N_13526,N_7186,N_8507);
or U13527 (N_13527,N_5715,N_7707);
and U13528 (N_13528,N_5365,N_7018);
and U13529 (N_13529,N_5857,N_5692);
nor U13530 (N_13530,N_7131,N_6174);
xor U13531 (N_13531,N_8865,N_7053);
nand U13532 (N_13532,N_5492,N_7832);
and U13533 (N_13533,N_9808,N_6758);
or U13534 (N_13534,N_5869,N_7923);
xor U13535 (N_13535,N_8688,N_5513);
nor U13536 (N_13536,N_7951,N_6523);
xnor U13537 (N_13537,N_9288,N_8569);
and U13538 (N_13538,N_5607,N_5626);
xor U13539 (N_13539,N_6425,N_6500);
and U13540 (N_13540,N_7478,N_9819);
or U13541 (N_13541,N_5741,N_6234);
xnor U13542 (N_13542,N_9569,N_9190);
or U13543 (N_13543,N_5645,N_6131);
or U13544 (N_13544,N_8927,N_8419);
nor U13545 (N_13545,N_5699,N_9678);
nor U13546 (N_13546,N_7563,N_7946);
nor U13547 (N_13547,N_5732,N_7026);
nand U13548 (N_13548,N_7928,N_5119);
nor U13549 (N_13549,N_8965,N_5505);
xnor U13550 (N_13550,N_8846,N_6773);
and U13551 (N_13551,N_5268,N_8033);
xor U13552 (N_13552,N_7977,N_9092);
xor U13553 (N_13553,N_6642,N_6423);
xor U13554 (N_13554,N_8893,N_7140);
nor U13555 (N_13555,N_9346,N_8048);
nor U13556 (N_13556,N_8730,N_8467);
and U13557 (N_13557,N_5927,N_5820);
or U13558 (N_13558,N_9462,N_6824);
nand U13559 (N_13559,N_5740,N_7677);
xor U13560 (N_13560,N_5038,N_8390);
nand U13561 (N_13561,N_9512,N_8205);
nor U13562 (N_13562,N_9113,N_9497);
nand U13563 (N_13563,N_9842,N_8463);
or U13564 (N_13564,N_7484,N_6437);
nand U13565 (N_13565,N_7959,N_9669);
xnor U13566 (N_13566,N_8644,N_8896);
nor U13567 (N_13567,N_6601,N_6183);
or U13568 (N_13568,N_9388,N_7274);
nor U13569 (N_13569,N_9168,N_7832);
xor U13570 (N_13570,N_7567,N_5881);
or U13571 (N_13571,N_5170,N_9408);
nand U13572 (N_13572,N_8455,N_5333);
nand U13573 (N_13573,N_8884,N_5913);
or U13574 (N_13574,N_5663,N_5678);
and U13575 (N_13575,N_7189,N_5302);
xor U13576 (N_13576,N_5271,N_9218);
xor U13577 (N_13577,N_5470,N_7867);
nor U13578 (N_13578,N_8657,N_5318);
nand U13579 (N_13579,N_5336,N_5709);
xor U13580 (N_13580,N_9067,N_6768);
or U13581 (N_13581,N_9174,N_7997);
nand U13582 (N_13582,N_6256,N_9189);
nand U13583 (N_13583,N_9334,N_8348);
nand U13584 (N_13584,N_7839,N_6320);
and U13585 (N_13585,N_7882,N_9521);
and U13586 (N_13586,N_8708,N_7615);
nand U13587 (N_13587,N_6200,N_8894);
or U13588 (N_13588,N_6644,N_7150);
xor U13589 (N_13589,N_6429,N_9427);
or U13590 (N_13590,N_9197,N_6632);
or U13591 (N_13591,N_8935,N_7408);
or U13592 (N_13592,N_6426,N_9972);
xor U13593 (N_13593,N_5369,N_5769);
or U13594 (N_13594,N_9707,N_5553);
nor U13595 (N_13595,N_9382,N_6769);
xnor U13596 (N_13596,N_7467,N_7201);
or U13597 (N_13597,N_6336,N_6981);
nor U13598 (N_13598,N_7234,N_6339);
or U13599 (N_13599,N_5434,N_6623);
or U13600 (N_13600,N_6604,N_9947);
or U13601 (N_13601,N_5458,N_8874);
xnor U13602 (N_13602,N_9495,N_8614);
xor U13603 (N_13603,N_8730,N_9004);
nand U13604 (N_13604,N_8084,N_5927);
nor U13605 (N_13605,N_6480,N_5773);
xor U13606 (N_13606,N_5407,N_5997);
and U13607 (N_13607,N_7368,N_9984);
nand U13608 (N_13608,N_7794,N_5893);
nand U13609 (N_13609,N_8927,N_9090);
and U13610 (N_13610,N_6322,N_7269);
nor U13611 (N_13611,N_6145,N_7817);
and U13612 (N_13612,N_8676,N_9283);
xor U13613 (N_13613,N_8557,N_7316);
nor U13614 (N_13614,N_6883,N_6514);
or U13615 (N_13615,N_9451,N_5693);
or U13616 (N_13616,N_9327,N_6930);
nor U13617 (N_13617,N_6771,N_5451);
xor U13618 (N_13618,N_9454,N_9370);
nor U13619 (N_13619,N_9091,N_5087);
xor U13620 (N_13620,N_6998,N_9980);
nor U13621 (N_13621,N_5398,N_9520);
nand U13622 (N_13622,N_9011,N_8836);
and U13623 (N_13623,N_5226,N_9346);
nand U13624 (N_13624,N_9965,N_6103);
xnor U13625 (N_13625,N_6301,N_7816);
xor U13626 (N_13626,N_8556,N_9574);
xnor U13627 (N_13627,N_5148,N_8067);
nor U13628 (N_13628,N_7269,N_8304);
or U13629 (N_13629,N_8276,N_7673);
or U13630 (N_13630,N_7858,N_7901);
and U13631 (N_13631,N_8600,N_9139);
xnor U13632 (N_13632,N_7036,N_5391);
xnor U13633 (N_13633,N_5390,N_5233);
and U13634 (N_13634,N_5884,N_7350);
xor U13635 (N_13635,N_6011,N_6074);
nor U13636 (N_13636,N_7819,N_5160);
nor U13637 (N_13637,N_5763,N_8190);
xor U13638 (N_13638,N_9355,N_5313);
or U13639 (N_13639,N_6176,N_5319);
xor U13640 (N_13640,N_9539,N_5214);
nand U13641 (N_13641,N_8711,N_8308);
and U13642 (N_13642,N_8502,N_8320);
or U13643 (N_13643,N_6232,N_8142);
and U13644 (N_13644,N_6948,N_6352);
nor U13645 (N_13645,N_9351,N_9110);
or U13646 (N_13646,N_5017,N_7914);
and U13647 (N_13647,N_5912,N_6053);
nand U13648 (N_13648,N_5760,N_9960);
and U13649 (N_13649,N_8911,N_9048);
nor U13650 (N_13650,N_5249,N_5973);
or U13651 (N_13651,N_5917,N_9296);
xor U13652 (N_13652,N_8687,N_8657);
or U13653 (N_13653,N_6224,N_6010);
or U13654 (N_13654,N_5393,N_6276);
or U13655 (N_13655,N_9845,N_9934);
or U13656 (N_13656,N_5621,N_6346);
or U13657 (N_13657,N_8021,N_8497);
and U13658 (N_13658,N_8563,N_7985);
xnor U13659 (N_13659,N_7385,N_7124);
or U13660 (N_13660,N_5161,N_6834);
xnor U13661 (N_13661,N_9173,N_5798);
and U13662 (N_13662,N_9626,N_5094);
or U13663 (N_13663,N_6124,N_5830);
and U13664 (N_13664,N_7964,N_8591);
or U13665 (N_13665,N_6297,N_7353);
nor U13666 (N_13666,N_7680,N_7630);
and U13667 (N_13667,N_8715,N_7782);
or U13668 (N_13668,N_5425,N_8272);
xor U13669 (N_13669,N_8473,N_9942);
nor U13670 (N_13670,N_7092,N_7985);
and U13671 (N_13671,N_8595,N_7051);
xor U13672 (N_13672,N_6680,N_6173);
or U13673 (N_13673,N_7061,N_6784);
nor U13674 (N_13674,N_6477,N_5887);
nor U13675 (N_13675,N_5790,N_9254);
nor U13676 (N_13676,N_5973,N_6434);
nand U13677 (N_13677,N_5653,N_8009);
xor U13678 (N_13678,N_6113,N_8347);
xnor U13679 (N_13679,N_8569,N_7331);
nand U13680 (N_13680,N_5461,N_7753);
nor U13681 (N_13681,N_8126,N_6058);
and U13682 (N_13682,N_6363,N_9953);
nor U13683 (N_13683,N_9472,N_6448);
xnor U13684 (N_13684,N_7330,N_6715);
and U13685 (N_13685,N_6695,N_7700);
and U13686 (N_13686,N_8263,N_9383);
xnor U13687 (N_13687,N_6093,N_6282);
xor U13688 (N_13688,N_8296,N_8760);
or U13689 (N_13689,N_9735,N_5071);
or U13690 (N_13690,N_9385,N_9387);
xnor U13691 (N_13691,N_5420,N_5842);
and U13692 (N_13692,N_6726,N_7274);
nor U13693 (N_13693,N_8987,N_5821);
and U13694 (N_13694,N_7324,N_7000);
xor U13695 (N_13695,N_8344,N_8777);
xor U13696 (N_13696,N_8709,N_7856);
xor U13697 (N_13697,N_7358,N_6496);
nand U13698 (N_13698,N_9206,N_8439);
or U13699 (N_13699,N_7689,N_7969);
nor U13700 (N_13700,N_7032,N_9263);
nand U13701 (N_13701,N_9098,N_6030);
nor U13702 (N_13702,N_9932,N_5578);
and U13703 (N_13703,N_9649,N_8548);
nand U13704 (N_13704,N_5037,N_5684);
and U13705 (N_13705,N_8819,N_6963);
xor U13706 (N_13706,N_5319,N_9926);
nor U13707 (N_13707,N_5223,N_5728);
nand U13708 (N_13708,N_7393,N_9309);
or U13709 (N_13709,N_7461,N_8444);
nor U13710 (N_13710,N_7566,N_5108);
nor U13711 (N_13711,N_9246,N_5396);
nand U13712 (N_13712,N_5810,N_6196);
or U13713 (N_13713,N_9320,N_5541);
nor U13714 (N_13714,N_7473,N_7511);
or U13715 (N_13715,N_9924,N_8023);
xor U13716 (N_13716,N_5075,N_6473);
nand U13717 (N_13717,N_8188,N_8499);
or U13718 (N_13718,N_7536,N_5927);
xor U13719 (N_13719,N_7221,N_9647);
nand U13720 (N_13720,N_9707,N_5924);
xor U13721 (N_13721,N_7319,N_5483);
nand U13722 (N_13722,N_5856,N_8328);
nor U13723 (N_13723,N_8446,N_5689);
nand U13724 (N_13724,N_6841,N_8533);
and U13725 (N_13725,N_5455,N_8467);
xnor U13726 (N_13726,N_8981,N_7250);
nor U13727 (N_13727,N_7533,N_7597);
xor U13728 (N_13728,N_9617,N_7400);
and U13729 (N_13729,N_8776,N_6212);
nor U13730 (N_13730,N_9105,N_5678);
and U13731 (N_13731,N_5074,N_7232);
nor U13732 (N_13732,N_5255,N_8688);
and U13733 (N_13733,N_5071,N_9010);
nor U13734 (N_13734,N_6926,N_8849);
or U13735 (N_13735,N_5927,N_7709);
nand U13736 (N_13736,N_9486,N_7970);
or U13737 (N_13737,N_6491,N_9813);
nor U13738 (N_13738,N_7416,N_6305);
nor U13739 (N_13739,N_8807,N_5681);
nor U13740 (N_13740,N_5145,N_5239);
or U13741 (N_13741,N_5760,N_9701);
nand U13742 (N_13742,N_6572,N_6258);
nor U13743 (N_13743,N_9333,N_8040);
or U13744 (N_13744,N_9953,N_7351);
and U13745 (N_13745,N_8531,N_8436);
nor U13746 (N_13746,N_9401,N_6506);
nor U13747 (N_13747,N_7092,N_5276);
nor U13748 (N_13748,N_8776,N_5890);
and U13749 (N_13749,N_9868,N_6864);
nand U13750 (N_13750,N_7278,N_9387);
nand U13751 (N_13751,N_5357,N_9859);
nand U13752 (N_13752,N_7957,N_6904);
and U13753 (N_13753,N_7123,N_6216);
and U13754 (N_13754,N_5530,N_6355);
nand U13755 (N_13755,N_7379,N_7929);
or U13756 (N_13756,N_9819,N_7768);
nand U13757 (N_13757,N_7230,N_9059);
nand U13758 (N_13758,N_7276,N_7635);
and U13759 (N_13759,N_5894,N_9370);
or U13760 (N_13760,N_9570,N_6735);
and U13761 (N_13761,N_5883,N_7529);
nand U13762 (N_13762,N_5849,N_8809);
and U13763 (N_13763,N_9241,N_7514);
nand U13764 (N_13764,N_6375,N_9557);
and U13765 (N_13765,N_8848,N_7973);
and U13766 (N_13766,N_8211,N_7988);
xor U13767 (N_13767,N_8601,N_6800);
and U13768 (N_13768,N_7768,N_7343);
nand U13769 (N_13769,N_6126,N_6872);
xor U13770 (N_13770,N_5525,N_5857);
and U13771 (N_13771,N_5769,N_8601);
or U13772 (N_13772,N_7416,N_5477);
nor U13773 (N_13773,N_7402,N_8649);
xnor U13774 (N_13774,N_9909,N_9516);
xor U13775 (N_13775,N_6959,N_9626);
xnor U13776 (N_13776,N_7935,N_6820);
nand U13777 (N_13777,N_7606,N_6236);
xnor U13778 (N_13778,N_7877,N_7006);
or U13779 (N_13779,N_9671,N_8082);
and U13780 (N_13780,N_5514,N_7593);
or U13781 (N_13781,N_9189,N_9187);
nand U13782 (N_13782,N_6599,N_5257);
or U13783 (N_13783,N_9321,N_5821);
or U13784 (N_13784,N_9898,N_5410);
or U13785 (N_13785,N_8816,N_8009);
or U13786 (N_13786,N_5558,N_7320);
and U13787 (N_13787,N_6812,N_8464);
xnor U13788 (N_13788,N_8358,N_7777);
nor U13789 (N_13789,N_9725,N_5485);
or U13790 (N_13790,N_6879,N_7064);
and U13791 (N_13791,N_5290,N_8555);
nand U13792 (N_13792,N_8174,N_7386);
and U13793 (N_13793,N_7245,N_8034);
or U13794 (N_13794,N_8269,N_9072);
nand U13795 (N_13795,N_6692,N_5905);
nand U13796 (N_13796,N_9715,N_9468);
nand U13797 (N_13797,N_6638,N_7040);
xor U13798 (N_13798,N_5098,N_8859);
nand U13799 (N_13799,N_8674,N_6103);
nor U13800 (N_13800,N_7743,N_6271);
nand U13801 (N_13801,N_9665,N_8112);
and U13802 (N_13802,N_9763,N_8495);
or U13803 (N_13803,N_5101,N_6004);
nor U13804 (N_13804,N_6444,N_7695);
nor U13805 (N_13805,N_5889,N_5595);
or U13806 (N_13806,N_6073,N_7024);
nor U13807 (N_13807,N_9784,N_7674);
nor U13808 (N_13808,N_9105,N_6236);
nand U13809 (N_13809,N_7880,N_8764);
and U13810 (N_13810,N_5495,N_7532);
or U13811 (N_13811,N_5147,N_9552);
nand U13812 (N_13812,N_9582,N_5656);
nand U13813 (N_13813,N_9915,N_5290);
and U13814 (N_13814,N_9583,N_9294);
nor U13815 (N_13815,N_9147,N_6780);
nand U13816 (N_13816,N_5620,N_9891);
or U13817 (N_13817,N_8567,N_6579);
nand U13818 (N_13818,N_6778,N_7678);
xor U13819 (N_13819,N_7662,N_9248);
nand U13820 (N_13820,N_5988,N_5977);
or U13821 (N_13821,N_7290,N_8004);
or U13822 (N_13822,N_6319,N_7837);
or U13823 (N_13823,N_6954,N_6657);
or U13824 (N_13824,N_9479,N_5846);
nand U13825 (N_13825,N_9996,N_6400);
and U13826 (N_13826,N_8172,N_6768);
nor U13827 (N_13827,N_7531,N_5755);
xor U13828 (N_13828,N_7511,N_8031);
xor U13829 (N_13829,N_5082,N_6271);
or U13830 (N_13830,N_5979,N_7746);
and U13831 (N_13831,N_5736,N_5556);
and U13832 (N_13832,N_5105,N_7137);
or U13833 (N_13833,N_6657,N_9989);
or U13834 (N_13834,N_6533,N_7988);
and U13835 (N_13835,N_7833,N_8519);
nand U13836 (N_13836,N_9864,N_9476);
or U13837 (N_13837,N_7137,N_6425);
nand U13838 (N_13838,N_5288,N_7152);
xnor U13839 (N_13839,N_5135,N_6387);
xnor U13840 (N_13840,N_7353,N_9431);
nand U13841 (N_13841,N_5890,N_8334);
nand U13842 (N_13842,N_9773,N_9326);
or U13843 (N_13843,N_6211,N_7056);
and U13844 (N_13844,N_7344,N_5171);
and U13845 (N_13845,N_7398,N_7127);
nor U13846 (N_13846,N_5998,N_9146);
or U13847 (N_13847,N_6057,N_5344);
nand U13848 (N_13848,N_7669,N_9679);
or U13849 (N_13849,N_9511,N_8420);
and U13850 (N_13850,N_7761,N_7815);
or U13851 (N_13851,N_8170,N_8685);
nand U13852 (N_13852,N_9537,N_7976);
or U13853 (N_13853,N_6123,N_8398);
nand U13854 (N_13854,N_5815,N_9032);
or U13855 (N_13855,N_7372,N_9984);
and U13856 (N_13856,N_9320,N_7498);
or U13857 (N_13857,N_7147,N_5158);
nand U13858 (N_13858,N_6944,N_6379);
xnor U13859 (N_13859,N_9328,N_9716);
xnor U13860 (N_13860,N_6908,N_7635);
nor U13861 (N_13861,N_6487,N_5933);
or U13862 (N_13862,N_6289,N_5446);
or U13863 (N_13863,N_9412,N_9096);
or U13864 (N_13864,N_6504,N_5197);
nand U13865 (N_13865,N_6385,N_7914);
or U13866 (N_13866,N_7102,N_9007);
nor U13867 (N_13867,N_9231,N_7057);
nor U13868 (N_13868,N_8825,N_9028);
and U13869 (N_13869,N_7916,N_9354);
nand U13870 (N_13870,N_7273,N_8320);
or U13871 (N_13871,N_9446,N_9206);
nand U13872 (N_13872,N_8871,N_8908);
nor U13873 (N_13873,N_8204,N_6029);
nor U13874 (N_13874,N_8735,N_8199);
or U13875 (N_13875,N_8827,N_9095);
xnor U13876 (N_13876,N_6678,N_7080);
or U13877 (N_13877,N_6151,N_6379);
and U13878 (N_13878,N_9010,N_6185);
or U13879 (N_13879,N_7342,N_9023);
nor U13880 (N_13880,N_8534,N_9268);
and U13881 (N_13881,N_6519,N_7832);
or U13882 (N_13882,N_9894,N_6810);
xor U13883 (N_13883,N_7651,N_6833);
xnor U13884 (N_13884,N_8231,N_5449);
nand U13885 (N_13885,N_7204,N_8704);
xnor U13886 (N_13886,N_8418,N_7174);
and U13887 (N_13887,N_5242,N_5858);
xor U13888 (N_13888,N_9361,N_7668);
xnor U13889 (N_13889,N_7218,N_6225);
nand U13890 (N_13890,N_5553,N_7643);
and U13891 (N_13891,N_5562,N_7432);
or U13892 (N_13892,N_5067,N_9491);
or U13893 (N_13893,N_9313,N_6069);
xor U13894 (N_13894,N_9062,N_7762);
and U13895 (N_13895,N_6259,N_5922);
or U13896 (N_13896,N_8774,N_9766);
xor U13897 (N_13897,N_5884,N_5309);
nor U13898 (N_13898,N_6137,N_6334);
and U13899 (N_13899,N_9595,N_7763);
and U13900 (N_13900,N_8496,N_6514);
xnor U13901 (N_13901,N_8165,N_7571);
and U13902 (N_13902,N_9216,N_7247);
nand U13903 (N_13903,N_9188,N_5004);
nor U13904 (N_13904,N_9120,N_9207);
xor U13905 (N_13905,N_6233,N_9607);
or U13906 (N_13906,N_7792,N_9313);
and U13907 (N_13907,N_8053,N_5164);
or U13908 (N_13908,N_8306,N_6408);
or U13909 (N_13909,N_8989,N_7481);
and U13910 (N_13910,N_5942,N_9426);
xor U13911 (N_13911,N_8472,N_6708);
nor U13912 (N_13912,N_8533,N_5462);
nor U13913 (N_13913,N_6100,N_5784);
xor U13914 (N_13914,N_7125,N_6589);
xor U13915 (N_13915,N_8803,N_8399);
xnor U13916 (N_13916,N_5462,N_5357);
xor U13917 (N_13917,N_8578,N_8782);
nand U13918 (N_13918,N_5283,N_7878);
xor U13919 (N_13919,N_6453,N_6652);
or U13920 (N_13920,N_7215,N_5913);
nand U13921 (N_13921,N_5035,N_6412);
xor U13922 (N_13922,N_5379,N_5312);
nand U13923 (N_13923,N_5635,N_8073);
nand U13924 (N_13924,N_6688,N_5239);
xor U13925 (N_13925,N_5081,N_6874);
nand U13926 (N_13926,N_7826,N_7972);
and U13927 (N_13927,N_7934,N_7221);
or U13928 (N_13928,N_9559,N_8377);
xnor U13929 (N_13929,N_8689,N_7618);
or U13930 (N_13930,N_9500,N_8671);
xnor U13931 (N_13931,N_7264,N_7722);
nor U13932 (N_13932,N_5024,N_8382);
or U13933 (N_13933,N_5012,N_7723);
xnor U13934 (N_13934,N_7608,N_6635);
xor U13935 (N_13935,N_6560,N_9713);
or U13936 (N_13936,N_8970,N_8495);
or U13937 (N_13937,N_7438,N_7419);
nor U13938 (N_13938,N_7629,N_5108);
xnor U13939 (N_13939,N_6642,N_8856);
and U13940 (N_13940,N_6106,N_6703);
and U13941 (N_13941,N_6707,N_5904);
nor U13942 (N_13942,N_8228,N_5934);
nand U13943 (N_13943,N_6172,N_6177);
xor U13944 (N_13944,N_8737,N_9617);
or U13945 (N_13945,N_8147,N_7736);
nor U13946 (N_13946,N_9218,N_5721);
or U13947 (N_13947,N_8171,N_7824);
and U13948 (N_13948,N_5457,N_8614);
nand U13949 (N_13949,N_6411,N_9517);
and U13950 (N_13950,N_8414,N_6742);
nand U13951 (N_13951,N_7386,N_7925);
and U13952 (N_13952,N_9475,N_6080);
nand U13953 (N_13953,N_9009,N_6450);
nand U13954 (N_13954,N_6000,N_7759);
or U13955 (N_13955,N_6007,N_8529);
or U13956 (N_13956,N_5520,N_6853);
and U13957 (N_13957,N_9873,N_6514);
nand U13958 (N_13958,N_7774,N_7028);
nor U13959 (N_13959,N_5541,N_9278);
xor U13960 (N_13960,N_7658,N_7083);
nor U13961 (N_13961,N_5017,N_9772);
nand U13962 (N_13962,N_8923,N_5325);
or U13963 (N_13963,N_8972,N_8395);
nor U13964 (N_13964,N_6935,N_6582);
nand U13965 (N_13965,N_9158,N_7592);
nor U13966 (N_13966,N_9956,N_5025);
xnor U13967 (N_13967,N_6632,N_5213);
nor U13968 (N_13968,N_6403,N_9114);
and U13969 (N_13969,N_6339,N_5130);
nand U13970 (N_13970,N_6407,N_7619);
nor U13971 (N_13971,N_9033,N_6969);
nor U13972 (N_13972,N_8228,N_5848);
and U13973 (N_13973,N_8392,N_9433);
nor U13974 (N_13974,N_9270,N_7874);
and U13975 (N_13975,N_5728,N_5991);
nor U13976 (N_13976,N_9204,N_6535);
or U13977 (N_13977,N_7981,N_9268);
nand U13978 (N_13978,N_6353,N_7406);
xor U13979 (N_13979,N_6560,N_6145);
and U13980 (N_13980,N_9172,N_6984);
nand U13981 (N_13981,N_8027,N_6694);
xnor U13982 (N_13982,N_9854,N_8854);
or U13983 (N_13983,N_9382,N_6990);
nand U13984 (N_13984,N_8671,N_7906);
xor U13985 (N_13985,N_7074,N_7073);
or U13986 (N_13986,N_7521,N_5939);
or U13987 (N_13987,N_8299,N_9426);
nor U13988 (N_13988,N_7941,N_8809);
and U13989 (N_13989,N_6832,N_5969);
and U13990 (N_13990,N_5624,N_7388);
xnor U13991 (N_13991,N_6951,N_9289);
or U13992 (N_13992,N_8216,N_5185);
nor U13993 (N_13993,N_6390,N_9842);
nand U13994 (N_13994,N_6772,N_7581);
and U13995 (N_13995,N_9848,N_9268);
and U13996 (N_13996,N_8556,N_9774);
nand U13997 (N_13997,N_7861,N_9439);
or U13998 (N_13998,N_7698,N_9661);
nand U13999 (N_13999,N_5963,N_9904);
and U14000 (N_14000,N_8642,N_8637);
nand U14001 (N_14001,N_7485,N_6028);
xnor U14002 (N_14002,N_9771,N_7806);
nand U14003 (N_14003,N_5459,N_5393);
xor U14004 (N_14004,N_6050,N_6873);
xnor U14005 (N_14005,N_5821,N_8480);
nor U14006 (N_14006,N_9482,N_8704);
nand U14007 (N_14007,N_7377,N_6433);
or U14008 (N_14008,N_5119,N_8634);
nor U14009 (N_14009,N_6899,N_9240);
nor U14010 (N_14010,N_8968,N_6431);
nor U14011 (N_14011,N_5567,N_8861);
or U14012 (N_14012,N_5518,N_7951);
nand U14013 (N_14013,N_5155,N_9691);
nand U14014 (N_14014,N_7168,N_9273);
and U14015 (N_14015,N_6231,N_8161);
nor U14016 (N_14016,N_9971,N_9511);
and U14017 (N_14017,N_9707,N_5338);
nand U14018 (N_14018,N_7535,N_9988);
xor U14019 (N_14019,N_8922,N_9530);
or U14020 (N_14020,N_8150,N_8585);
nor U14021 (N_14021,N_6294,N_5223);
xor U14022 (N_14022,N_8850,N_8759);
and U14023 (N_14023,N_5278,N_6138);
nand U14024 (N_14024,N_5249,N_6549);
nand U14025 (N_14025,N_6886,N_8391);
and U14026 (N_14026,N_8442,N_6492);
xnor U14027 (N_14027,N_7490,N_7896);
nor U14028 (N_14028,N_8913,N_6143);
nor U14029 (N_14029,N_9363,N_7296);
nor U14030 (N_14030,N_5627,N_6081);
and U14031 (N_14031,N_9767,N_8309);
nand U14032 (N_14032,N_6009,N_8961);
or U14033 (N_14033,N_8955,N_7104);
nor U14034 (N_14034,N_5280,N_5276);
nand U14035 (N_14035,N_7438,N_9138);
or U14036 (N_14036,N_8967,N_6440);
and U14037 (N_14037,N_5150,N_6498);
or U14038 (N_14038,N_9477,N_7814);
xor U14039 (N_14039,N_5327,N_6597);
or U14040 (N_14040,N_9929,N_6953);
nor U14041 (N_14041,N_5046,N_7763);
and U14042 (N_14042,N_8326,N_6473);
and U14043 (N_14043,N_9046,N_9829);
or U14044 (N_14044,N_7242,N_6375);
nand U14045 (N_14045,N_6324,N_6656);
xor U14046 (N_14046,N_8495,N_7240);
nor U14047 (N_14047,N_6605,N_5020);
nand U14048 (N_14048,N_7674,N_5876);
or U14049 (N_14049,N_7379,N_6104);
nor U14050 (N_14050,N_6179,N_8237);
nor U14051 (N_14051,N_7292,N_6591);
and U14052 (N_14052,N_9195,N_9460);
or U14053 (N_14053,N_5567,N_6981);
nor U14054 (N_14054,N_9525,N_8409);
nand U14055 (N_14055,N_8342,N_5012);
nand U14056 (N_14056,N_8701,N_7872);
nand U14057 (N_14057,N_5526,N_5884);
or U14058 (N_14058,N_9481,N_7701);
nor U14059 (N_14059,N_7148,N_8110);
nor U14060 (N_14060,N_6786,N_5364);
nand U14061 (N_14061,N_5055,N_7028);
or U14062 (N_14062,N_7390,N_8389);
nand U14063 (N_14063,N_8453,N_9221);
or U14064 (N_14064,N_9263,N_5469);
nand U14065 (N_14065,N_6497,N_8939);
nand U14066 (N_14066,N_7095,N_5832);
nand U14067 (N_14067,N_6259,N_5499);
nand U14068 (N_14068,N_9437,N_8292);
nor U14069 (N_14069,N_7209,N_6541);
nand U14070 (N_14070,N_7468,N_8368);
xor U14071 (N_14071,N_5533,N_8006);
and U14072 (N_14072,N_6250,N_9080);
xnor U14073 (N_14073,N_7114,N_5707);
and U14074 (N_14074,N_7327,N_7874);
xnor U14075 (N_14075,N_5383,N_5756);
nand U14076 (N_14076,N_7427,N_8546);
and U14077 (N_14077,N_7822,N_6328);
or U14078 (N_14078,N_7613,N_9806);
or U14079 (N_14079,N_5524,N_5623);
or U14080 (N_14080,N_9784,N_7308);
nor U14081 (N_14081,N_5708,N_6847);
nand U14082 (N_14082,N_9784,N_8927);
or U14083 (N_14083,N_7168,N_9553);
and U14084 (N_14084,N_9941,N_7056);
xnor U14085 (N_14085,N_5162,N_8046);
and U14086 (N_14086,N_7771,N_5436);
xor U14087 (N_14087,N_8576,N_5705);
nor U14088 (N_14088,N_6331,N_7877);
or U14089 (N_14089,N_9910,N_7170);
nor U14090 (N_14090,N_7634,N_7622);
or U14091 (N_14091,N_8485,N_6423);
nor U14092 (N_14092,N_7854,N_8416);
nor U14093 (N_14093,N_6310,N_9691);
nand U14094 (N_14094,N_7617,N_5835);
xor U14095 (N_14095,N_6591,N_8442);
or U14096 (N_14096,N_7795,N_9609);
and U14097 (N_14097,N_7305,N_9298);
nand U14098 (N_14098,N_6500,N_7048);
nor U14099 (N_14099,N_6174,N_5590);
nand U14100 (N_14100,N_6123,N_9999);
nor U14101 (N_14101,N_6862,N_6316);
nand U14102 (N_14102,N_9796,N_5479);
or U14103 (N_14103,N_8818,N_7254);
and U14104 (N_14104,N_7937,N_8879);
nor U14105 (N_14105,N_9157,N_6548);
and U14106 (N_14106,N_9906,N_8691);
xor U14107 (N_14107,N_5809,N_9750);
and U14108 (N_14108,N_9399,N_5749);
xnor U14109 (N_14109,N_6815,N_5167);
and U14110 (N_14110,N_6510,N_9276);
xor U14111 (N_14111,N_8416,N_5295);
or U14112 (N_14112,N_8635,N_8969);
or U14113 (N_14113,N_9214,N_6996);
nor U14114 (N_14114,N_9309,N_9449);
nand U14115 (N_14115,N_6950,N_5514);
xor U14116 (N_14116,N_5025,N_9622);
nor U14117 (N_14117,N_8359,N_9122);
and U14118 (N_14118,N_7991,N_6435);
or U14119 (N_14119,N_5836,N_5202);
xnor U14120 (N_14120,N_8566,N_5938);
or U14121 (N_14121,N_8752,N_6130);
nor U14122 (N_14122,N_5662,N_5380);
or U14123 (N_14123,N_9391,N_6892);
and U14124 (N_14124,N_6442,N_6969);
nor U14125 (N_14125,N_5451,N_7775);
nand U14126 (N_14126,N_6337,N_5220);
and U14127 (N_14127,N_7592,N_9292);
nor U14128 (N_14128,N_6528,N_7966);
xnor U14129 (N_14129,N_7670,N_8692);
or U14130 (N_14130,N_9704,N_9502);
and U14131 (N_14131,N_7713,N_9760);
nand U14132 (N_14132,N_9414,N_9816);
xnor U14133 (N_14133,N_5331,N_9589);
nor U14134 (N_14134,N_6528,N_6879);
nor U14135 (N_14135,N_9629,N_5532);
xor U14136 (N_14136,N_5718,N_7268);
or U14137 (N_14137,N_9406,N_5931);
nand U14138 (N_14138,N_6554,N_7897);
nand U14139 (N_14139,N_7227,N_8169);
nor U14140 (N_14140,N_9720,N_9668);
nand U14141 (N_14141,N_9886,N_9602);
and U14142 (N_14142,N_5906,N_5825);
nand U14143 (N_14143,N_5555,N_6907);
or U14144 (N_14144,N_6630,N_5857);
xor U14145 (N_14145,N_5209,N_5865);
xor U14146 (N_14146,N_9037,N_7538);
or U14147 (N_14147,N_7122,N_8229);
nand U14148 (N_14148,N_6820,N_5765);
nor U14149 (N_14149,N_8138,N_7940);
xor U14150 (N_14150,N_5937,N_5930);
nor U14151 (N_14151,N_5110,N_9681);
nor U14152 (N_14152,N_8290,N_5254);
xor U14153 (N_14153,N_6390,N_8576);
xor U14154 (N_14154,N_8781,N_9386);
xnor U14155 (N_14155,N_6347,N_7979);
xor U14156 (N_14156,N_6303,N_5592);
or U14157 (N_14157,N_6497,N_5152);
or U14158 (N_14158,N_8460,N_5264);
or U14159 (N_14159,N_7257,N_9617);
nand U14160 (N_14160,N_7150,N_6459);
and U14161 (N_14161,N_7129,N_6888);
nand U14162 (N_14162,N_7055,N_8449);
and U14163 (N_14163,N_6308,N_7370);
nand U14164 (N_14164,N_8307,N_9220);
or U14165 (N_14165,N_9931,N_5825);
and U14166 (N_14166,N_6102,N_5256);
and U14167 (N_14167,N_7805,N_5239);
and U14168 (N_14168,N_8490,N_9445);
xnor U14169 (N_14169,N_6846,N_7464);
nand U14170 (N_14170,N_5515,N_6617);
nor U14171 (N_14171,N_5098,N_7800);
nor U14172 (N_14172,N_9641,N_8333);
or U14173 (N_14173,N_9252,N_5532);
and U14174 (N_14174,N_8885,N_9172);
xor U14175 (N_14175,N_6076,N_5279);
nor U14176 (N_14176,N_6808,N_6492);
nand U14177 (N_14177,N_9394,N_5536);
and U14178 (N_14178,N_9665,N_9553);
or U14179 (N_14179,N_7836,N_8731);
and U14180 (N_14180,N_5005,N_9097);
or U14181 (N_14181,N_6454,N_9354);
nor U14182 (N_14182,N_7912,N_5029);
nor U14183 (N_14183,N_9862,N_5028);
nor U14184 (N_14184,N_6469,N_8251);
nor U14185 (N_14185,N_9504,N_5273);
nand U14186 (N_14186,N_8613,N_5338);
nor U14187 (N_14187,N_8967,N_8676);
or U14188 (N_14188,N_7459,N_8257);
nor U14189 (N_14189,N_8011,N_8488);
and U14190 (N_14190,N_6282,N_8327);
or U14191 (N_14191,N_5554,N_5542);
nand U14192 (N_14192,N_6610,N_7237);
nand U14193 (N_14193,N_8768,N_8828);
xnor U14194 (N_14194,N_5149,N_7985);
nor U14195 (N_14195,N_5782,N_7164);
nor U14196 (N_14196,N_9662,N_8014);
and U14197 (N_14197,N_5439,N_5524);
and U14198 (N_14198,N_5395,N_7416);
or U14199 (N_14199,N_8290,N_9663);
nor U14200 (N_14200,N_5120,N_5385);
nor U14201 (N_14201,N_8541,N_8545);
xnor U14202 (N_14202,N_9082,N_7385);
nand U14203 (N_14203,N_8270,N_7557);
and U14204 (N_14204,N_8029,N_6598);
xor U14205 (N_14205,N_6111,N_8029);
xnor U14206 (N_14206,N_5106,N_7344);
nand U14207 (N_14207,N_5910,N_9862);
nand U14208 (N_14208,N_8230,N_5142);
or U14209 (N_14209,N_8612,N_9374);
xor U14210 (N_14210,N_5494,N_7336);
or U14211 (N_14211,N_7472,N_7535);
and U14212 (N_14212,N_9387,N_5358);
nand U14213 (N_14213,N_9584,N_8165);
or U14214 (N_14214,N_5828,N_5854);
nand U14215 (N_14215,N_5440,N_7670);
xnor U14216 (N_14216,N_8542,N_8640);
and U14217 (N_14217,N_5029,N_7322);
and U14218 (N_14218,N_8433,N_9720);
nor U14219 (N_14219,N_6337,N_6712);
and U14220 (N_14220,N_8257,N_8031);
and U14221 (N_14221,N_9397,N_7692);
nand U14222 (N_14222,N_5130,N_7483);
and U14223 (N_14223,N_6276,N_7308);
nor U14224 (N_14224,N_6480,N_7054);
xnor U14225 (N_14225,N_8072,N_6912);
nor U14226 (N_14226,N_7367,N_5092);
or U14227 (N_14227,N_6694,N_8158);
and U14228 (N_14228,N_9730,N_7996);
nor U14229 (N_14229,N_5182,N_8911);
nor U14230 (N_14230,N_7821,N_7253);
or U14231 (N_14231,N_5569,N_8911);
xnor U14232 (N_14232,N_9010,N_6512);
nor U14233 (N_14233,N_8376,N_6353);
nor U14234 (N_14234,N_7186,N_9306);
xor U14235 (N_14235,N_7858,N_9475);
xor U14236 (N_14236,N_8481,N_5756);
nor U14237 (N_14237,N_5190,N_8338);
nor U14238 (N_14238,N_5351,N_9467);
nand U14239 (N_14239,N_5822,N_9437);
or U14240 (N_14240,N_8204,N_5420);
or U14241 (N_14241,N_9319,N_6762);
nand U14242 (N_14242,N_9378,N_8842);
or U14243 (N_14243,N_7676,N_9738);
or U14244 (N_14244,N_6000,N_7909);
and U14245 (N_14245,N_7974,N_9957);
and U14246 (N_14246,N_6560,N_8352);
and U14247 (N_14247,N_8585,N_8490);
and U14248 (N_14248,N_9401,N_5693);
xnor U14249 (N_14249,N_6943,N_6666);
nand U14250 (N_14250,N_7874,N_5656);
and U14251 (N_14251,N_9601,N_5780);
and U14252 (N_14252,N_9406,N_5284);
and U14253 (N_14253,N_6053,N_7630);
and U14254 (N_14254,N_5225,N_6642);
xnor U14255 (N_14255,N_8661,N_5657);
or U14256 (N_14256,N_9311,N_7803);
nand U14257 (N_14257,N_6057,N_6469);
xnor U14258 (N_14258,N_6633,N_7808);
or U14259 (N_14259,N_9107,N_5251);
or U14260 (N_14260,N_8858,N_7756);
or U14261 (N_14261,N_6058,N_6974);
nor U14262 (N_14262,N_7722,N_8783);
and U14263 (N_14263,N_9307,N_5665);
nor U14264 (N_14264,N_8140,N_7409);
or U14265 (N_14265,N_6811,N_7329);
and U14266 (N_14266,N_8270,N_5385);
nand U14267 (N_14267,N_7238,N_8233);
or U14268 (N_14268,N_6758,N_8266);
and U14269 (N_14269,N_6049,N_5688);
or U14270 (N_14270,N_7183,N_7577);
nand U14271 (N_14271,N_9500,N_6357);
nand U14272 (N_14272,N_5735,N_7783);
nor U14273 (N_14273,N_7660,N_9072);
xor U14274 (N_14274,N_9632,N_7407);
and U14275 (N_14275,N_6482,N_5175);
nor U14276 (N_14276,N_8535,N_6822);
or U14277 (N_14277,N_8078,N_8123);
nor U14278 (N_14278,N_8366,N_7482);
xnor U14279 (N_14279,N_7161,N_6992);
and U14280 (N_14280,N_9644,N_7750);
xnor U14281 (N_14281,N_8394,N_8136);
or U14282 (N_14282,N_7881,N_8223);
xor U14283 (N_14283,N_9411,N_6906);
or U14284 (N_14284,N_8316,N_5244);
nand U14285 (N_14285,N_6903,N_9556);
and U14286 (N_14286,N_8116,N_9268);
or U14287 (N_14287,N_9171,N_9276);
and U14288 (N_14288,N_7942,N_6167);
xor U14289 (N_14289,N_7877,N_7532);
or U14290 (N_14290,N_9791,N_6268);
or U14291 (N_14291,N_9457,N_7117);
nand U14292 (N_14292,N_5792,N_7621);
nand U14293 (N_14293,N_8057,N_9210);
and U14294 (N_14294,N_6453,N_7396);
or U14295 (N_14295,N_9280,N_6578);
or U14296 (N_14296,N_9785,N_7199);
and U14297 (N_14297,N_9073,N_7312);
xor U14298 (N_14298,N_9873,N_5524);
xnor U14299 (N_14299,N_5812,N_9465);
xnor U14300 (N_14300,N_7924,N_5542);
and U14301 (N_14301,N_5588,N_9771);
or U14302 (N_14302,N_9493,N_9507);
nand U14303 (N_14303,N_9874,N_6032);
or U14304 (N_14304,N_5202,N_7962);
nand U14305 (N_14305,N_9564,N_7887);
xor U14306 (N_14306,N_9163,N_7038);
nor U14307 (N_14307,N_5510,N_6957);
xnor U14308 (N_14308,N_6492,N_5687);
nand U14309 (N_14309,N_7227,N_5660);
or U14310 (N_14310,N_6679,N_9700);
and U14311 (N_14311,N_9942,N_6646);
xnor U14312 (N_14312,N_6157,N_6155);
and U14313 (N_14313,N_9707,N_9030);
xnor U14314 (N_14314,N_7169,N_5407);
xor U14315 (N_14315,N_9540,N_7816);
nand U14316 (N_14316,N_8672,N_7700);
nor U14317 (N_14317,N_7496,N_5199);
and U14318 (N_14318,N_5924,N_6491);
xnor U14319 (N_14319,N_7736,N_9621);
nor U14320 (N_14320,N_9422,N_7342);
xnor U14321 (N_14321,N_7335,N_9618);
xor U14322 (N_14322,N_9070,N_7581);
nand U14323 (N_14323,N_8031,N_8419);
and U14324 (N_14324,N_7208,N_7254);
nor U14325 (N_14325,N_6672,N_5808);
xor U14326 (N_14326,N_6426,N_9473);
xnor U14327 (N_14327,N_7752,N_7930);
or U14328 (N_14328,N_6560,N_5872);
and U14329 (N_14329,N_9922,N_5053);
or U14330 (N_14330,N_8720,N_8147);
or U14331 (N_14331,N_8209,N_7685);
xor U14332 (N_14332,N_7685,N_8593);
nor U14333 (N_14333,N_5623,N_6771);
or U14334 (N_14334,N_6822,N_9780);
or U14335 (N_14335,N_8581,N_5104);
nor U14336 (N_14336,N_9005,N_7915);
nor U14337 (N_14337,N_7002,N_6518);
or U14338 (N_14338,N_5432,N_7178);
xnor U14339 (N_14339,N_9773,N_9333);
or U14340 (N_14340,N_5566,N_7610);
or U14341 (N_14341,N_8410,N_6295);
or U14342 (N_14342,N_7252,N_8568);
or U14343 (N_14343,N_5137,N_8862);
xor U14344 (N_14344,N_9773,N_7870);
or U14345 (N_14345,N_9699,N_5895);
xnor U14346 (N_14346,N_7920,N_6002);
and U14347 (N_14347,N_6070,N_9537);
nor U14348 (N_14348,N_9276,N_8270);
nor U14349 (N_14349,N_8710,N_8773);
and U14350 (N_14350,N_7110,N_7005);
xor U14351 (N_14351,N_9482,N_5548);
nand U14352 (N_14352,N_7566,N_8344);
xnor U14353 (N_14353,N_9377,N_7085);
and U14354 (N_14354,N_8012,N_6171);
and U14355 (N_14355,N_9258,N_9232);
xor U14356 (N_14356,N_6283,N_6194);
and U14357 (N_14357,N_9246,N_9540);
or U14358 (N_14358,N_5248,N_5164);
nor U14359 (N_14359,N_7842,N_9748);
and U14360 (N_14360,N_8651,N_8326);
nand U14361 (N_14361,N_6355,N_7327);
nor U14362 (N_14362,N_6034,N_9534);
xor U14363 (N_14363,N_6902,N_6234);
nand U14364 (N_14364,N_8797,N_6134);
nand U14365 (N_14365,N_9175,N_5093);
xor U14366 (N_14366,N_5615,N_7299);
nor U14367 (N_14367,N_7187,N_8578);
nand U14368 (N_14368,N_8387,N_5195);
xnor U14369 (N_14369,N_5794,N_9160);
and U14370 (N_14370,N_9312,N_6620);
xnor U14371 (N_14371,N_9356,N_6717);
xor U14372 (N_14372,N_9146,N_8444);
nand U14373 (N_14373,N_6523,N_6772);
nand U14374 (N_14374,N_6906,N_8895);
and U14375 (N_14375,N_7728,N_6900);
nand U14376 (N_14376,N_8670,N_9541);
or U14377 (N_14377,N_5106,N_6591);
and U14378 (N_14378,N_5911,N_6855);
xnor U14379 (N_14379,N_8180,N_6165);
and U14380 (N_14380,N_6736,N_8857);
and U14381 (N_14381,N_7552,N_5861);
nand U14382 (N_14382,N_7109,N_8711);
nor U14383 (N_14383,N_8754,N_8013);
xnor U14384 (N_14384,N_7958,N_6811);
xnor U14385 (N_14385,N_5796,N_9818);
xor U14386 (N_14386,N_5864,N_6137);
xnor U14387 (N_14387,N_5646,N_5184);
xor U14388 (N_14388,N_6990,N_7114);
and U14389 (N_14389,N_7578,N_5833);
or U14390 (N_14390,N_9185,N_7632);
nor U14391 (N_14391,N_8519,N_5629);
and U14392 (N_14392,N_7740,N_9512);
xor U14393 (N_14393,N_6769,N_9812);
nand U14394 (N_14394,N_9296,N_6660);
nor U14395 (N_14395,N_6173,N_5404);
or U14396 (N_14396,N_8227,N_5247);
and U14397 (N_14397,N_6738,N_7594);
or U14398 (N_14398,N_9971,N_8826);
and U14399 (N_14399,N_8614,N_9137);
nor U14400 (N_14400,N_8888,N_8334);
or U14401 (N_14401,N_8830,N_6223);
nor U14402 (N_14402,N_8372,N_9369);
xnor U14403 (N_14403,N_9493,N_5790);
nand U14404 (N_14404,N_9589,N_9954);
nand U14405 (N_14405,N_6471,N_6561);
and U14406 (N_14406,N_5391,N_7524);
xor U14407 (N_14407,N_7596,N_5673);
nor U14408 (N_14408,N_8002,N_6397);
nor U14409 (N_14409,N_5048,N_8870);
nand U14410 (N_14410,N_7866,N_8498);
or U14411 (N_14411,N_5981,N_7084);
nor U14412 (N_14412,N_5394,N_9455);
nor U14413 (N_14413,N_5275,N_7258);
and U14414 (N_14414,N_7468,N_7783);
and U14415 (N_14415,N_9007,N_5995);
nand U14416 (N_14416,N_5061,N_6223);
and U14417 (N_14417,N_7237,N_7949);
or U14418 (N_14418,N_7953,N_5096);
nand U14419 (N_14419,N_6397,N_7430);
xor U14420 (N_14420,N_7671,N_8762);
and U14421 (N_14421,N_6940,N_8950);
or U14422 (N_14422,N_7077,N_7004);
and U14423 (N_14423,N_8787,N_7253);
nor U14424 (N_14424,N_8204,N_5715);
nor U14425 (N_14425,N_6128,N_8726);
or U14426 (N_14426,N_9041,N_5060);
xor U14427 (N_14427,N_9495,N_9864);
xor U14428 (N_14428,N_7107,N_9085);
nor U14429 (N_14429,N_9475,N_8427);
or U14430 (N_14430,N_9497,N_9472);
nor U14431 (N_14431,N_5049,N_8421);
or U14432 (N_14432,N_7998,N_7785);
xor U14433 (N_14433,N_7077,N_6191);
nand U14434 (N_14434,N_9536,N_6309);
xor U14435 (N_14435,N_5650,N_5459);
nor U14436 (N_14436,N_9622,N_7800);
and U14437 (N_14437,N_9739,N_6238);
or U14438 (N_14438,N_6415,N_5059);
or U14439 (N_14439,N_6496,N_9732);
nor U14440 (N_14440,N_9339,N_6190);
or U14441 (N_14441,N_7193,N_9574);
or U14442 (N_14442,N_7617,N_6775);
and U14443 (N_14443,N_5287,N_7242);
or U14444 (N_14444,N_9322,N_5065);
nand U14445 (N_14445,N_6694,N_6969);
nor U14446 (N_14446,N_9014,N_5695);
nand U14447 (N_14447,N_7155,N_7124);
or U14448 (N_14448,N_7080,N_9594);
and U14449 (N_14449,N_5759,N_7730);
and U14450 (N_14450,N_9623,N_6530);
or U14451 (N_14451,N_8957,N_8399);
nand U14452 (N_14452,N_9693,N_9945);
xor U14453 (N_14453,N_7833,N_7544);
or U14454 (N_14454,N_7010,N_5344);
nand U14455 (N_14455,N_7210,N_6362);
and U14456 (N_14456,N_7762,N_8482);
and U14457 (N_14457,N_6240,N_9259);
or U14458 (N_14458,N_7531,N_8314);
nor U14459 (N_14459,N_5047,N_5157);
nor U14460 (N_14460,N_9874,N_5894);
nand U14461 (N_14461,N_7568,N_6342);
xor U14462 (N_14462,N_5046,N_7962);
nand U14463 (N_14463,N_5689,N_9591);
xnor U14464 (N_14464,N_7982,N_7540);
xor U14465 (N_14465,N_5365,N_7706);
or U14466 (N_14466,N_8065,N_6112);
or U14467 (N_14467,N_8399,N_7177);
xnor U14468 (N_14468,N_5230,N_6429);
and U14469 (N_14469,N_7794,N_7032);
and U14470 (N_14470,N_6403,N_7627);
and U14471 (N_14471,N_8563,N_5060);
xor U14472 (N_14472,N_5222,N_7708);
xor U14473 (N_14473,N_7021,N_9418);
nor U14474 (N_14474,N_5084,N_8502);
nor U14475 (N_14475,N_9453,N_9875);
nor U14476 (N_14476,N_6770,N_7299);
nand U14477 (N_14477,N_6329,N_8153);
nand U14478 (N_14478,N_6559,N_9050);
or U14479 (N_14479,N_7292,N_5683);
and U14480 (N_14480,N_7061,N_5144);
nor U14481 (N_14481,N_7195,N_6118);
nand U14482 (N_14482,N_7064,N_9835);
and U14483 (N_14483,N_5108,N_7903);
and U14484 (N_14484,N_9645,N_9203);
nor U14485 (N_14485,N_9593,N_7509);
or U14486 (N_14486,N_8120,N_5347);
xor U14487 (N_14487,N_8197,N_5394);
xnor U14488 (N_14488,N_5255,N_6619);
nand U14489 (N_14489,N_8229,N_7690);
or U14490 (N_14490,N_5430,N_9939);
or U14491 (N_14491,N_7276,N_5998);
or U14492 (N_14492,N_5259,N_5368);
and U14493 (N_14493,N_8764,N_7262);
nor U14494 (N_14494,N_5866,N_8552);
or U14495 (N_14495,N_5762,N_6236);
nor U14496 (N_14496,N_5102,N_6995);
or U14497 (N_14497,N_9163,N_6791);
and U14498 (N_14498,N_5114,N_9084);
xnor U14499 (N_14499,N_9837,N_5272);
nand U14500 (N_14500,N_5956,N_6647);
or U14501 (N_14501,N_8584,N_7566);
or U14502 (N_14502,N_5713,N_9155);
nor U14503 (N_14503,N_5943,N_5614);
nor U14504 (N_14504,N_5936,N_9796);
xnor U14505 (N_14505,N_6109,N_7095);
xnor U14506 (N_14506,N_8663,N_5784);
nand U14507 (N_14507,N_7618,N_8105);
nand U14508 (N_14508,N_9016,N_7672);
or U14509 (N_14509,N_8668,N_7802);
xor U14510 (N_14510,N_8048,N_5665);
or U14511 (N_14511,N_8639,N_6106);
or U14512 (N_14512,N_8760,N_7083);
xnor U14513 (N_14513,N_5393,N_6324);
xor U14514 (N_14514,N_9425,N_6212);
xnor U14515 (N_14515,N_9965,N_5923);
xor U14516 (N_14516,N_8845,N_8241);
and U14517 (N_14517,N_9434,N_5345);
or U14518 (N_14518,N_9458,N_6585);
nand U14519 (N_14519,N_8103,N_8844);
or U14520 (N_14520,N_6566,N_5537);
xnor U14521 (N_14521,N_9597,N_9799);
xnor U14522 (N_14522,N_5707,N_9735);
xor U14523 (N_14523,N_9216,N_7546);
and U14524 (N_14524,N_7512,N_5825);
nand U14525 (N_14525,N_8987,N_9963);
nor U14526 (N_14526,N_8183,N_9995);
nand U14527 (N_14527,N_8897,N_5442);
nor U14528 (N_14528,N_7630,N_9290);
nor U14529 (N_14529,N_7382,N_5961);
or U14530 (N_14530,N_9001,N_6698);
nand U14531 (N_14531,N_9170,N_5290);
nand U14532 (N_14532,N_7582,N_6593);
nor U14533 (N_14533,N_9612,N_7740);
nor U14534 (N_14534,N_9854,N_9728);
and U14535 (N_14535,N_6468,N_6803);
nand U14536 (N_14536,N_9939,N_6452);
and U14537 (N_14537,N_5123,N_7353);
or U14538 (N_14538,N_7400,N_6086);
or U14539 (N_14539,N_6963,N_5380);
and U14540 (N_14540,N_6865,N_9945);
nand U14541 (N_14541,N_5785,N_7393);
and U14542 (N_14542,N_5170,N_9809);
nand U14543 (N_14543,N_9814,N_9463);
nand U14544 (N_14544,N_8336,N_9759);
or U14545 (N_14545,N_6283,N_8857);
and U14546 (N_14546,N_5309,N_7797);
or U14547 (N_14547,N_9776,N_7298);
nand U14548 (N_14548,N_6424,N_9218);
and U14549 (N_14549,N_5399,N_9865);
nand U14550 (N_14550,N_8271,N_5407);
xor U14551 (N_14551,N_8147,N_5881);
or U14552 (N_14552,N_7470,N_8657);
or U14553 (N_14553,N_7659,N_6328);
nand U14554 (N_14554,N_5767,N_9721);
nor U14555 (N_14555,N_6543,N_7306);
nor U14556 (N_14556,N_6339,N_8105);
xor U14557 (N_14557,N_9151,N_9556);
nor U14558 (N_14558,N_5466,N_7110);
nor U14559 (N_14559,N_6660,N_9013);
nand U14560 (N_14560,N_7250,N_9539);
or U14561 (N_14561,N_6261,N_9583);
nand U14562 (N_14562,N_8849,N_8418);
and U14563 (N_14563,N_9517,N_7793);
nand U14564 (N_14564,N_9339,N_9505);
nor U14565 (N_14565,N_9663,N_7637);
and U14566 (N_14566,N_7115,N_7581);
xnor U14567 (N_14567,N_8776,N_8022);
nor U14568 (N_14568,N_5802,N_7424);
or U14569 (N_14569,N_5513,N_5905);
or U14570 (N_14570,N_9790,N_8074);
xnor U14571 (N_14571,N_8668,N_5679);
and U14572 (N_14572,N_8176,N_8223);
or U14573 (N_14573,N_5229,N_7799);
xnor U14574 (N_14574,N_8733,N_7723);
nand U14575 (N_14575,N_8639,N_6411);
and U14576 (N_14576,N_9927,N_6885);
xnor U14577 (N_14577,N_7321,N_5582);
or U14578 (N_14578,N_5846,N_8351);
and U14579 (N_14579,N_5089,N_7288);
xnor U14580 (N_14580,N_9905,N_8220);
xor U14581 (N_14581,N_7552,N_7352);
or U14582 (N_14582,N_8228,N_9501);
nor U14583 (N_14583,N_6222,N_9729);
or U14584 (N_14584,N_5595,N_6319);
or U14585 (N_14585,N_9721,N_6427);
nor U14586 (N_14586,N_6200,N_9327);
and U14587 (N_14587,N_7393,N_7784);
and U14588 (N_14588,N_9175,N_5393);
and U14589 (N_14589,N_5415,N_6317);
or U14590 (N_14590,N_7433,N_8917);
nor U14591 (N_14591,N_6907,N_8431);
xnor U14592 (N_14592,N_7869,N_7855);
and U14593 (N_14593,N_6763,N_6494);
nor U14594 (N_14594,N_5377,N_7857);
xor U14595 (N_14595,N_7509,N_9525);
nand U14596 (N_14596,N_6273,N_6477);
nand U14597 (N_14597,N_8778,N_6313);
or U14598 (N_14598,N_7619,N_5238);
or U14599 (N_14599,N_5847,N_8035);
or U14600 (N_14600,N_7127,N_8970);
nor U14601 (N_14601,N_6363,N_9562);
xor U14602 (N_14602,N_6977,N_8336);
or U14603 (N_14603,N_8081,N_9328);
and U14604 (N_14604,N_6543,N_8560);
nor U14605 (N_14605,N_7486,N_5946);
nand U14606 (N_14606,N_9340,N_7787);
xor U14607 (N_14607,N_5566,N_8418);
nor U14608 (N_14608,N_8442,N_7849);
or U14609 (N_14609,N_6695,N_9144);
and U14610 (N_14610,N_6338,N_5926);
and U14611 (N_14611,N_5183,N_7848);
xor U14612 (N_14612,N_6171,N_9626);
nor U14613 (N_14613,N_8820,N_6279);
and U14614 (N_14614,N_7903,N_9607);
or U14615 (N_14615,N_8170,N_7598);
nand U14616 (N_14616,N_9938,N_6760);
xnor U14617 (N_14617,N_7586,N_6856);
or U14618 (N_14618,N_9211,N_9774);
and U14619 (N_14619,N_6077,N_8592);
and U14620 (N_14620,N_9620,N_8996);
or U14621 (N_14621,N_5855,N_6658);
nor U14622 (N_14622,N_7161,N_6730);
nand U14623 (N_14623,N_5994,N_9758);
and U14624 (N_14624,N_6860,N_6499);
or U14625 (N_14625,N_8473,N_7442);
and U14626 (N_14626,N_9398,N_7634);
nor U14627 (N_14627,N_5791,N_8063);
nand U14628 (N_14628,N_8125,N_9612);
nor U14629 (N_14629,N_6824,N_9238);
xor U14630 (N_14630,N_6613,N_8462);
and U14631 (N_14631,N_8982,N_8199);
nand U14632 (N_14632,N_7871,N_8257);
nor U14633 (N_14633,N_5177,N_7946);
and U14634 (N_14634,N_9266,N_8348);
and U14635 (N_14635,N_7526,N_9761);
xor U14636 (N_14636,N_7278,N_6562);
nor U14637 (N_14637,N_5681,N_8029);
and U14638 (N_14638,N_8809,N_9496);
or U14639 (N_14639,N_9495,N_5734);
xor U14640 (N_14640,N_5466,N_5011);
or U14641 (N_14641,N_8865,N_5028);
nor U14642 (N_14642,N_7722,N_5330);
or U14643 (N_14643,N_5980,N_9837);
xor U14644 (N_14644,N_5357,N_7295);
xnor U14645 (N_14645,N_5400,N_6622);
nor U14646 (N_14646,N_5770,N_6329);
xor U14647 (N_14647,N_8330,N_5875);
nor U14648 (N_14648,N_8592,N_7279);
nor U14649 (N_14649,N_5334,N_8071);
and U14650 (N_14650,N_9958,N_7852);
xnor U14651 (N_14651,N_8313,N_6942);
nor U14652 (N_14652,N_5419,N_5596);
nor U14653 (N_14653,N_8958,N_5376);
and U14654 (N_14654,N_5748,N_7932);
nor U14655 (N_14655,N_7594,N_5921);
nand U14656 (N_14656,N_9513,N_8358);
and U14657 (N_14657,N_7511,N_9496);
xnor U14658 (N_14658,N_7089,N_9480);
or U14659 (N_14659,N_5550,N_7336);
or U14660 (N_14660,N_6119,N_5019);
or U14661 (N_14661,N_5528,N_8045);
nand U14662 (N_14662,N_5774,N_9957);
nand U14663 (N_14663,N_6099,N_6164);
nand U14664 (N_14664,N_6961,N_7823);
or U14665 (N_14665,N_9715,N_7854);
and U14666 (N_14666,N_8582,N_5855);
and U14667 (N_14667,N_5597,N_7559);
and U14668 (N_14668,N_5202,N_5099);
nand U14669 (N_14669,N_7360,N_9898);
nand U14670 (N_14670,N_6326,N_7370);
and U14671 (N_14671,N_6687,N_8814);
or U14672 (N_14672,N_7286,N_7293);
nand U14673 (N_14673,N_5354,N_9416);
xnor U14674 (N_14674,N_7682,N_5614);
or U14675 (N_14675,N_7982,N_9317);
or U14676 (N_14676,N_5277,N_9347);
nand U14677 (N_14677,N_9128,N_7705);
nand U14678 (N_14678,N_7306,N_8230);
nor U14679 (N_14679,N_7257,N_6641);
nand U14680 (N_14680,N_6055,N_9185);
nor U14681 (N_14681,N_7744,N_9061);
or U14682 (N_14682,N_9123,N_8170);
and U14683 (N_14683,N_5555,N_7184);
nor U14684 (N_14684,N_6745,N_5890);
nand U14685 (N_14685,N_6771,N_8442);
nor U14686 (N_14686,N_7012,N_6160);
or U14687 (N_14687,N_8783,N_6793);
and U14688 (N_14688,N_9464,N_8976);
nor U14689 (N_14689,N_7071,N_5269);
and U14690 (N_14690,N_6904,N_5214);
nand U14691 (N_14691,N_5566,N_8186);
xor U14692 (N_14692,N_6805,N_8891);
or U14693 (N_14693,N_7736,N_7433);
nor U14694 (N_14694,N_5284,N_6053);
nor U14695 (N_14695,N_8438,N_5284);
or U14696 (N_14696,N_7587,N_9236);
nor U14697 (N_14697,N_7296,N_9840);
or U14698 (N_14698,N_7869,N_9374);
nand U14699 (N_14699,N_5482,N_9856);
or U14700 (N_14700,N_7814,N_9820);
nor U14701 (N_14701,N_5886,N_6503);
or U14702 (N_14702,N_7723,N_6477);
xor U14703 (N_14703,N_9064,N_7174);
and U14704 (N_14704,N_9538,N_5905);
or U14705 (N_14705,N_8408,N_5388);
nand U14706 (N_14706,N_8487,N_6801);
nand U14707 (N_14707,N_9531,N_6042);
and U14708 (N_14708,N_7946,N_6081);
and U14709 (N_14709,N_5466,N_6265);
nor U14710 (N_14710,N_7386,N_5509);
nor U14711 (N_14711,N_6887,N_8539);
xnor U14712 (N_14712,N_6111,N_7097);
and U14713 (N_14713,N_6057,N_9199);
and U14714 (N_14714,N_8072,N_6443);
nand U14715 (N_14715,N_5046,N_7085);
xor U14716 (N_14716,N_6290,N_9709);
nand U14717 (N_14717,N_7046,N_6800);
and U14718 (N_14718,N_8497,N_5446);
nor U14719 (N_14719,N_5093,N_9202);
or U14720 (N_14720,N_8531,N_7879);
or U14721 (N_14721,N_8189,N_9268);
nor U14722 (N_14722,N_9513,N_9519);
nand U14723 (N_14723,N_7977,N_7253);
nand U14724 (N_14724,N_8103,N_9883);
and U14725 (N_14725,N_6360,N_9194);
nor U14726 (N_14726,N_7580,N_5761);
nand U14727 (N_14727,N_8791,N_8570);
and U14728 (N_14728,N_6282,N_8065);
and U14729 (N_14729,N_5652,N_9473);
and U14730 (N_14730,N_9877,N_9367);
xor U14731 (N_14731,N_8644,N_5177);
or U14732 (N_14732,N_9043,N_9632);
xor U14733 (N_14733,N_6633,N_9516);
and U14734 (N_14734,N_6826,N_7043);
and U14735 (N_14735,N_5712,N_9512);
xor U14736 (N_14736,N_5933,N_9920);
or U14737 (N_14737,N_9284,N_5618);
nand U14738 (N_14738,N_6799,N_5432);
or U14739 (N_14739,N_9908,N_9450);
xor U14740 (N_14740,N_8204,N_7770);
and U14741 (N_14741,N_6420,N_7151);
xor U14742 (N_14742,N_8260,N_6243);
nor U14743 (N_14743,N_5957,N_7058);
or U14744 (N_14744,N_7639,N_6491);
nand U14745 (N_14745,N_5924,N_7298);
and U14746 (N_14746,N_6011,N_8025);
nand U14747 (N_14747,N_5488,N_7613);
or U14748 (N_14748,N_9848,N_5502);
xnor U14749 (N_14749,N_6896,N_5792);
nand U14750 (N_14750,N_9475,N_8395);
and U14751 (N_14751,N_7571,N_7091);
xor U14752 (N_14752,N_9196,N_5017);
and U14753 (N_14753,N_7718,N_8509);
nand U14754 (N_14754,N_7311,N_6265);
xor U14755 (N_14755,N_6003,N_5178);
or U14756 (N_14756,N_6564,N_6949);
xor U14757 (N_14757,N_9522,N_7910);
xnor U14758 (N_14758,N_8785,N_6630);
xor U14759 (N_14759,N_6365,N_5339);
nor U14760 (N_14760,N_5806,N_6102);
nand U14761 (N_14761,N_5375,N_5354);
or U14762 (N_14762,N_8078,N_7106);
or U14763 (N_14763,N_5980,N_5945);
nor U14764 (N_14764,N_5048,N_8394);
xnor U14765 (N_14765,N_8156,N_7334);
nor U14766 (N_14766,N_6087,N_6563);
or U14767 (N_14767,N_5388,N_5913);
nand U14768 (N_14768,N_7991,N_8110);
and U14769 (N_14769,N_7277,N_7713);
or U14770 (N_14770,N_8924,N_5467);
xor U14771 (N_14771,N_6845,N_8348);
nor U14772 (N_14772,N_7592,N_5810);
nor U14773 (N_14773,N_9726,N_7083);
and U14774 (N_14774,N_5116,N_9780);
nor U14775 (N_14775,N_9267,N_7207);
or U14776 (N_14776,N_5854,N_8047);
nand U14777 (N_14777,N_7194,N_9588);
nor U14778 (N_14778,N_9787,N_9154);
nand U14779 (N_14779,N_8532,N_9080);
nand U14780 (N_14780,N_7740,N_8349);
and U14781 (N_14781,N_8023,N_9330);
and U14782 (N_14782,N_8726,N_9594);
nor U14783 (N_14783,N_7582,N_7152);
nand U14784 (N_14784,N_6049,N_9050);
nand U14785 (N_14785,N_8279,N_6340);
or U14786 (N_14786,N_5511,N_8201);
nor U14787 (N_14787,N_8583,N_9800);
and U14788 (N_14788,N_9978,N_7738);
or U14789 (N_14789,N_6779,N_9571);
nor U14790 (N_14790,N_5349,N_7944);
nand U14791 (N_14791,N_5585,N_7576);
and U14792 (N_14792,N_6326,N_8046);
and U14793 (N_14793,N_5606,N_5185);
xor U14794 (N_14794,N_6421,N_8995);
and U14795 (N_14795,N_6210,N_9252);
or U14796 (N_14796,N_6688,N_5581);
nor U14797 (N_14797,N_5812,N_5357);
xor U14798 (N_14798,N_5953,N_7317);
nand U14799 (N_14799,N_8881,N_7912);
and U14800 (N_14800,N_5064,N_7109);
or U14801 (N_14801,N_9778,N_7521);
and U14802 (N_14802,N_6361,N_9347);
nand U14803 (N_14803,N_5161,N_5565);
nand U14804 (N_14804,N_9529,N_9712);
nor U14805 (N_14805,N_9016,N_9873);
nand U14806 (N_14806,N_7592,N_8116);
and U14807 (N_14807,N_6841,N_9306);
or U14808 (N_14808,N_5376,N_6878);
nand U14809 (N_14809,N_7548,N_8131);
and U14810 (N_14810,N_5469,N_7497);
nor U14811 (N_14811,N_8970,N_9394);
nor U14812 (N_14812,N_7704,N_7046);
nand U14813 (N_14813,N_6177,N_9416);
nor U14814 (N_14814,N_7739,N_6572);
or U14815 (N_14815,N_8993,N_7918);
xor U14816 (N_14816,N_9512,N_5647);
xor U14817 (N_14817,N_6140,N_6616);
nor U14818 (N_14818,N_5155,N_7171);
nand U14819 (N_14819,N_9426,N_9612);
nand U14820 (N_14820,N_8924,N_6481);
and U14821 (N_14821,N_8939,N_9484);
nor U14822 (N_14822,N_5511,N_7455);
nor U14823 (N_14823,N_9329,N_9179);
nand U14824 (N_14824,N_8178,N_8535);
nor U14825 (N_14825,N_7015,N_9144);
nand U14826 (N_14826,N_8850,N_8825);
nand U14827 (N_14827,N_6080,N_5671);
or U14828 (N_14828,N_9814,N_9308);
nand U14829 (N_14829,N_9536,N_5374);
and U14830 (N_14830,N_8720,N_6242);
or U14831 (N_14831,N_9651,N_5590);
or U14832 (N_14832,N_5458,N_5370);
xnor U14833 (N_14833,N_7235,N_7402);
nand U14834 (N_14834,N_5625,N_9370);
or U14835 (N_14835,N_6140,N_8423);
or U14836 (N_14836,N_5783,N_5478);
xor U14837 (N_14837,N_7671,N_5246);
or U14838 (N_14838,N_7886,N_6607);
xor U14839 (N_14839,N_9604,N_8520);
nand U14840 (N_14840,N_5241,N_8557);
nand U14841 (N_14841,N_6729,N_5377);
and U14842 (N_14842,N_7871,N_5962);
xor U14843 (N_14843,N_7746,N_6816);
nand U14844 (N_14844,N_7345,N_6916);
nand U14845 (N_14845,N_5855,N_5420);
nand U14846 (N_14846,N_8693,N_6484);
xor U14847 (N_14847,N_8105,N_6684);
or U14848 (N_14848,N_9250,N_8190);
and U14849 (N_14849,N_6844,N_5334);
or U14850 (N_14850,N_9262,N_8192);
xnor U14851 (N_14851,N_8950,N_5598);
xor U14852 (N_14852,N_6795,N_8633);
nor U14853 (N_14853,N_7422,N_9179);
xor U14854 (N_14854,N_7296,N_5137);
xor U14855 (N_14855,N_7997,N_8435);
xnor U14856 (N_14856,N_7057,N_8600);
nand U14857 (N_14857,N_6174,N_6744);
or U14858 (N_14858,N_9662,N_8284);
xnor U14859 (N_14859,N_6067,N_6249);
nor U14860 (N_14860,N_9698,N_6790);
nand U14861 (N_14861,N_6372,N_6021);
xor U14862 (N_14862,N_9853,N_9087);
xor U14863 (N_14863,N_5043,N_9319);
or U14864 (N_14864,N_7199,N_6599);
and U14865 (N_14865,N_8577,N_8244);
nor U14866 (N_14866,N_9158,N_9414);
xor U14867 (N_14867,N_5410,N_8575);
or U14868 (N_14868,N_6722,N_8845);
nor U14869 (N_14869,N_5207,N_5749);
or U14870 (N_14870,N_8897,N_9550);
xor U14871 (N_14871,N_8887,N_6714);
or U14872 (N_14872,N_9429,N_6198);
nand U14873 (N_14873,N_7447,N_8134);
nor U14874 (N_14874,N_8883,N_7610);
nand U14875 (N_14875,N_7431,N_6413);
and U14876 (N_14876,N_5468,N_6443);
nor U14877 (N_14877,N_5847,N_5000);
xor U14878 (N_14878,N_7730,N_8984);
nor U14879 (N_14879,N_7234,N_6912);
nor U14880 (N_14880,N_8136,N_7785);
or U14881 (N_14881,N_6242,N_5999);
or U14882 (N_14882,N_9625,N_7777);
and U14883 (N_14883,N_6486,N_8225);
xor U14884 (N_14884,N_6729,N_5009);
xor U14885 (N_14885,N_5891,N_7605);
or U14886 (N_14886,N_6526,N_5274);
nand U14887 (N_14887,N_8880,N_6239);
or U14888 (N_14888,N_5718,N_8167);
nor U14889 (N_14889,N_7576,N_5684);
nand U14890 (N_14890,N_8924,N_7023);
or U14891 (N_14891,N_5353,N_8618);
or U14892 (N_14892,N_7138,N_6003);
and U14893 (N_14893,N_9825,N_5177);
xor U14894 (N_14894,N_8780,N_6988);
xnor U14895 (N_14895,N_6521,N_8852);
nand U14896 (N_14896,N_7650,N_9996);
xnor U14897 (N_14897,N_9994,N_6083);
and U14898 (N_14898,N_9178,N_7810);
xnor U14899 (N_14899,N_8880,N_9866);
xnor U14900 (N_14900,N_6337,N_9920);
nor U14901 (N_14901,N_6028,N_9277);
nand U14902 (N_14902,N_8088,N_8338);
nand U14903 (N_14903,N_5501,N_6042);
xor U14904 (N_14904,N_8351,N_9407);
nor U14905 (N_14905,N_9338,N_5509);
or U14906 (N_14906,N_5346,N_9346);
or U14907 (N_14907,N_5502,N_5164);
or U14908 (N_14908,N_5815,N_9371);
nand U14909 (N_14909,N_7985,N_5392);
or U14910 (N_14910,N_8327,N_6511);
nor U14911 (N_14911,N_5248,N_9021);
or U14912 (N_14912,N_6740,N_5161);
nor U14913 (N_14913,N_6768,N_5379);
nand U14914 (N_14914,N_8549,N_8366);
nand U14915 (N_14915,N_6116,N_5235);
nor U14916 (N_14916,N_7745,N_8409);
and U14917 (N_14917,N_7431,N_6466);
xor U14918 (N_14918,N_6735,N_9079);
or U14919 (N_14919,N_8201,N_8362);
and U14920 (N_14920,N_5563,N_5499);
and U14921 (N_14921,N_7802,N_6103);
and U14922 (N_14922,N_5582,N_5838);
nor U14923 (N_14923,N_9750,N_9305);
or U14924 (N_14924,N_6507,N_7921);
xor U14925 (N_14925,N_5471,N_8067);
xnor U14926 (N_14926,N_9877,N_6730);
or U14927 (N_14927,N_8058,N_7040);
or U14928 (N_14928,N_7748,N_8624);
xnor U14929 (N_14929,N_5102,N_5361);
xnor U14930 (N_14930,N_7653,N_8486);
xnor U14931 (N_14931,N_8384,N_9499);
xnor U14932 (N_14932,N_6219,N_9915);
or U14933 (N_14933,N_7838,N_9580);
xor U14934 (N_14934,N_7689,N_7090);
nand U14935 (N_14935,N_7278,N_8812);
nand U14936 (N_14936,N_5209,N_5861);
nor U14937 (N_14937,N_9289,N_6710);
xor U14938 (N_14938,N_8339,N_9180);
or U14939 (N_14939,N_6771,N_9449);
nor U14940 (N_14940,N_5046,N_5731);
and U14941 (N_14941,N_8054,N_5972);
xor U14942 (N_14942,N_5525,N_9990);
or U14943 (N_14943,N_9774,N_5871);
or U14944 (N_14944,N_9667,N_5310);
nand U14945 (N_14945,N_7265,N_8063);
xor U14946 (N_14946,N_5980,N_8859);
nor U14947 (N_14947,N_5480,N_5939);
and U14948 (N_14948,N_8859,N_7917);
nand U14949 (N_14949,N_8536,N_5487);
nor U14950 (N_14950,N_8144,N_5510);
xor U14951 (N_14951,N_8158,N_8577);
or U14952 (N_14952,N_9682,N_7752);
xor U14953 (N_14953,N_8119,N_6130);
xnor U14954 (N_14954,N_7040,N_8208);
and U14955 (N_14955,N_8160,N_8961);
nor U14956 (N_14956,N_7643,N_5742);
nor U14957 (N_14957,N_7067,N_7011);
or U14958 (N_14958,N_7235,N_6701);
nand U14959 (N_14959,N_8859,N_8072);
and U14960 (N_14960,N_9174,N_6583);
nor U14961 (N_14961,N_5015,N_5792);
xor U14962 (N_14962,N_5522,N_8159);
nor U14963 (N_14963,N_9227,N_8739);
nor U14964 (N_14964,N_6839,N_6832);
or U14965 (N_14965,N_6603,N_9819);
nand U14966 (N_14966,N_8035,N_7432);
nand U14967 (N_14967,N_5312,N_6999);
nand U14968 (N_14968,N_7055,N_8337);
nand U14969 (N_14969,N_6554,N_9115);
or U14970 (N_14970,N_7968,N_6933);
nor U14971 (N_14971,N_8684,N_5067);
nor U14972 (N_14972,N_7511,N_6166);
nand U14973 (N_14973,N_9014,N_8494);
or U14974 (N_14974,N_7088,N_9545);
or U14975 (N_14975,N_9100,N_8388);
nand U14976 (N_14976,N_5417,N_6537);
xnor U14977 (N_14977,N_8677,N_5002);
nor U14978 (N_14978,N_6014,N_6495);
or U14979 (N_14979,N_5678,N_6347);
and U14980 (N_14980,N_8765,N_5254);
and U14981 (N_14981,N_6254,N_8324);
and U14982 (N_14982,N_7789,N_8349);
nand U14983 (N_14983,N_6949,N_6347);
and U14984 (N_14984,N_6864,N_5117);
nor U14985 (N_14985,N_8134,N_9727);
nor U14986 (N_14986,N_7615,N_5137);
nor U14987 (N_14987,N_8003,N_9844);
nor U14988 (N_14988,N_8124,N_9705);
or U14989 (N_14989,N_6170,N_8892);
xnor U14990 (N_14990,N_7091,N_9954);
or U14991 (N_14991,N_9494,N_8662);
and U14992 (N_14992,N_8023,N_5820);
or U14993 (N_14993,N_9547,N_8404);
and U14994 (N_14994,N_8181,N_5258);
nor U14995 (N_14995,N_9769,N_9681);
nand U14996 (N_14996,N_7907,N_9054);
and U14997 (N_14997,N_6978,N_6712);
xnor U14998 (N_14998,N_6624,N_7582);
nand U14999 (N_14999,N_5960,N_9468);
and U15000 (N_15000,N_13941,N_13169);
xnor U15001 (N_15001,N_12372,N_13140);
xnor U15002 (N_15002,N_12949,N_14017);
nand U15003 (N_15003,N_13062,N_12108);
nand U15004 (N_15004,N_13255,N_12672);
and U15005 (N_15005,N_12758,N_14263);
xnor U15006 (N_15006,N_12141,N_12289);
or U15007 (N_15007,N_10846,N_13238);
or U15008 (N_15008,N_13813,N_13240);
nand U15009 (N_15009,N_14175,N_13551);
and U15010 (N_15010,N_12168,N_10905);
nand U15011 (N_15011,N_14166,N_10779);
and U15012 (N_15012,N_11284,N_14875);
xnor U15013 (N_15013,N_14781,N_11109);
xnor U15014 (N_15014,N_13418,N_11854);
and U15015 (N_15015,N_13113,N_11601);
nand U15016 (N_15016,N_14709,N_13907);
xnor U15017 (N_15017,N_14458,N_10300);
or U15018 (N_15018,N_11505,N_13381);
and U15019 (N_15019,N_10099,N_11356);
nand U15020 (N_15020,N_10222,N_10490);
or U15021 (N_15021,N_11479,N_12238);
or U15022 (N_15022,N_10205,N_10096);
or U15023 (N_15023,N_10928,N_14176);
nor U15024 (N_15024,N_13477,N_10083);
or U15025 (N_15025,N_13825,N_11676);
or U15026 (N_15026,N_11001,N_13281);
nand U15027 (N_15027,N_11228,N_10832);
nand U15028 (N_15028,N_13469,N_14472);
nor U15029 (N_15029,N_13713,N_13965);
and U15030 (N_15030,N_13883,N_14305);
or U15031 (N_15031,N_14287,N_12216);
xnor U15032 (N_15032,N_13319,N_13804);
and U15033 (N_15033,N_12553,N_12480);
nor U15034 (N_15034,N_13518,N_14122);
and U15035 (N_15035,N_11937,N_10898);
xor U15036 (N_15036,N_10526,N_11891);
nand U15037 (N_15037,N_13686,N_12091);
xor U15038 (N_15038,N_12605,N_11757);
xnor U15039 (N_15039,N_13051,N_13337);
or U15040 (N_15040,N_13647,N_13746);
or U15041 (N_15041,N_12412,N_13996);
xnor U15042 (N_15042,N_10834,N_13975);
nor U15043 (N_15043,N_11899,N_13787);
or U15044 (N_15044,N_13884,N_12516);
nor U15045 (N_15045,N_14089,N_13642);
xor U15046 (N_15046,N_14269,N_10502);
xnor U15047 (N_15047,N_13373,N_11207);
and U15048 (N_15048,N_14370,N_13376);
xnor U15049 (N_15049,N_12433,N_11821);
nand U15050 (N_15050,N_14828,N_10101);
and U15051 (N_15051,N_12648,N_13680);
xnor U15052 (N_15052,N_12470,N_14173);
xnor U15053 (N_15053,N_11088,N_11996);
and U15054 (N_15054,N_14824,N_12835);
and U15055 (N_15055,N_14502,N_11585);
or U15056 (N_15056,N_14628,N_12531);
nand U15057 (N_15057,N_10460,N_11923);
nor U15058 (N_15058,N_10001,N_10376);
and U15059 (N_15059,N_10111,N_13390);
and U15060 (N_15060,N_10066,N_13993);
nor U15061 (N_15061,N_13872,N_12966);
or U15062 (N_15062,N_13425,N_13944);
or U15063 (N_15063,N_12101,N_11355);
nor U15064 (N_15064,N_12662,N_10295);
and U15065 (N_15065,N_11464,N_14994);
xor U15066 (N_15066,N_11111,N_10687);
nand U15067 (N_15067,N_14038,N_10173);
xnor U15068 (N_15068,N_13606,N_11625);
and U15069 (N_15069,N_11940,N_14174);
and U15070 (N_15070,N_10613,N_14009);
or U15071 (N_15071,N_11262,N_11221);
xor U15072 (N_15072,N_12765,N_10631);
nand U15073 (N_15073,N_14219,N_11906);
xnor U15074 (N_15074,N_10944,N_10864);
and U15075 (N_15075,N_10984,N_12431);
nand U15076 (N_15076,N_13502,N_13397);
xor U15077 (N_15077,N_11208,N_14001);
nor U15078 (N_15078,N_13249,N_10799);
xor U15079 (N_15079,N_13657,N_10122);
nand U15080 (N_15080,N_11860,N_12554);
nand U15081 (N_15081,N_11881,N_11481);
xnor U15082 (N_15082,N_11919,N_14278);
and U15083 (N_15083,N_12533,N_14304);
nor U15084 (N_15084,N_13192,N_12088);
nor U15085 (N_15085,N_13517,N_13268);
nor U15086 (N_15086,N_12436,N_12171);
xor U15087 (N_15087,N_10869,N_13382);
xnor U15088 (N_15088,N_12185,N_13478);
or U15089 (N_15089,N_12539,N_14046);
nand U15090 (N_15090,N_11289,N_10575);
xnor U15091 (N_15091,N_10335,N_10593);
or U15092 (N_15092,N_12110,N_11984);
and U15093 (N_15093,N_13842,N_13457);
nor U15094 (N_15094,N_10394,N_11810);
or U15095 (N_15095,N_13850,N_11368);
xnor U15096 (N_15096,N_14244,N_11204);
nand U15097 (N_15097,N_10647,N_11418);
nand U15098 (N_15098,N_12203,N_10450);
nand U15099 (N_15099,N_10621,N_13714);
and U15100 (N_15100,N_14598,N_13495);
nand U15101 (N_15101,N_10091,N_10492);
or U15102 (N_15102,N_12059,N_11801);
and U15103 (N_15103,N_10219,N_11215);
nand U15104 (N_15104,N_13359,N_11823);
nor U15105 (N_15105,N_10202,N_13733);
and U15106 (N_15106,N_12679,N_13404);
and U15107 (N_15107,N_13898,N_11133);
nor U15108 (N_15108,N_10074,N_13492);
xor U15109 (N_15109,N_14470,N_12428);
xnor U15110 (N_15110,N_12955,N_14109);
or U15111 (N_15111,N_14921,N_13383);
or U15112 (N_15112,N_11933,N_14876);
xor U15113 (N_15113,N_14347,N_14158);
and U15114 (N_15114,N_14185,N_14044);
nor U15115 (N_15115,N_14378,N_13563);
nand U15116 (N_15116,N_14388,N_13650);
and U15117 (N_15117,N_13833,N_13393);
and U15118 (N_15118,N_11931,N_13443);
xor U15119 (N_15119,N_14357,N_14084);
or U15120 (N_15120,N_13429,N_13945);
and U15121 (N_15121,N_10899,N_13936);
and U15122 (N_15122,N_14982,N_12705);
xnor U15123 (N_15123,N_14292,N_10155);
and U15124 (N_15124,N_14484,N_14005);
nor U15125 (N_15125,N_13147,N_11834);
xor U15126 (N_15126,N_11503,N_10212);
xnor U15127 (N_15127,N_12871,N_12286);
or U15128 (N_15128,N_13829,N_11077);
or U15129 (N_15129,N_11292,N_10599);
nor U15130 (N_15130,N_11312,N_11826);
nor U15131 (N_15131,N_11648,N_10038);
nor U15132 (N_15132,N_13776,N_14637);
xor U15133 (N_15133,N_10512,N_12330);
or U15134 (N_15134,N_11381,N_12825);
nand U15135 (N_15135,N_11715,N_13632);
nor U15136 (N_15136,N_14478,N_10058);
and U15137 (N_15137,N_12862,N_11236);
nand U15138 (N_15138,N_11015,N_12838);
or U15139 (N_15139,N_13835,N_10130);
xor U15140 (N_15140,N_11908,N_12696);
and U15141 (N_15141,N_12598,N_10589);
nor U15142 (N_15142,N_11402,N_14389);
nor U15143 (N_15143,N_13475,N_11622);
nand U15144 (N_15144,N_11125,N_11574);
nand U15145 (N_15145,N_11283,N_10748);
or U15146 (N_15146,N_13957,N_12063);
nor U15147 (N_15147,N_13282,N_13056);
or U15148 (N_15148,N_14755,N_14245);
or U15149 (N_15149,N_10031,N_12085);
nand U15150 (N_15150,N_12906,N_10412);
xnor U15151 (N_15151,N_14604,N_10851);
xnor U15152 (N_15152,N_12848,N_12034);
nor U15153 (N_15153,N_14178,N_13375);
xnor U15154 (N_15154,N_12723,N_12604);
nand U15155 (N_15155,N_14130,N_10178);
nand U15156 (N_15156,N_14193,N_10347);
and U15157 (N_15157,N_11305,N_12830);
nand U15158 (N_15158,N_11978,N_12644);
or U15159 (N_15159,N_13233,N_14400);
nand U15160 (N_15160,N_13782,N_10439);
and U15161 (N_15161,N_10041,N_14862);
and U15162 (N_15162,N_10642,N_11139);
xnor U15163 (N_15163,N_12469,N_13239);
xnor U15164 (N_15164,N_14640,N_11615);
nor U15165 (N_15165,N_11963,N_13914);
and U15166 (N_15166,N_14534,N_11980);
xnor U15167 (N_15167,N_11595,N_13866);
and U15168 (N_15168,N_11530,N_12146);
or U15169 (N_15169,N_14874,N_10800);
and U15170 (N_15170,N_13433,N_10257);
xnor U15171 (N_15171,N_10032,N_14566);
nand U15172 (N_15172,N_12288,N_11203);
nor U15173 (N_15173,N_14426,N_13926);
or U15174 (N_15174,N_14000,N_12664);
and U15175 (N_15175,N_10025,N_12131);
xnor U15176 (N_15176,N_11059,N_11918);
or U15177 (N_15177,N_14679,N_13274);
xor U15178 (N_15178,N_13560,N_12383);
nor U15179 (N_15179,N_13566,N_13507);
or U15180 (N_15180,N_13799,N_12150);
nand U15181 (N_15181,N_14843,N_14855);
nand U15182 (N_15182,N_10777,N_13174);
nor U15183 (N_15183,N_13949,N_11112);
or U15184 (N_15184,N_14354,N_14814);
xnor U15185 (N_15185,N_13540,N_11490);
nor U15186 (N_15186,N_12017,N_11375);
or U15187 (N_15187,N_12075,N_11778);
xor U15188 (N_15188,N_14528,N_13612);
and U15189 (N_15189,N_11995,N_12317);
or U15190 (N_15190,N_10005,N_12828);
and U15191 (N_15191,N_10421,N_13075);
nor U15192 (N_15192,N_14218,N_13868);
nor U15193 (N_15193,N_14999,N_12213);
nor U15194 (N_15194,N_14030,N_11451);
xnor U15195 (N_15195,N_13974,N_10540);
nand U15196 (N_15196,N_10209,N_14236);
and U15197 (N_15197,N_11539,N_14481);
nand U15198 (N_15198,N_10919,N_11831);
nor U15199 (N_15199,N_10780,N_13635);
xnor U15200 (N_15200,N_13526,N_13784);
and U15201 (N_15201,N_10420,N_14333);
nand U15202 (N_15202,N_13536,N_11740);
or U15203 (N_15203,N_13687,N_14976);
nor U15204 (N_15204,N_14054,N_12273);
or U15205 (N_15205,N_12635,N_12967);
xnor U15206 (N_15206,N_13942,N_14731);
xor U15207 (N_15207,N_12886,N_14662);
or U15208 (N_15208,N_14799,N_14606);
or U15209 (N_15209,N_11085,N_13508);
or U15210 (N_15210,N_12432,N_12524);
xnor U15211 (N_15211,N_10885,N_10211);
and U15212 (N_15212,N_13439,N_10027);
nor U15213 (N_15213,N_14264,N_14677);
nand U15214 (N_15214,N_12822,N_13740);
or U15215 (N_15215,N_10579,N_10226);
xor U15216 (N_15216,N_11813,N_10148);
and U15217 (N_15217,N_12087,N_10560);
nor U15218 (N_15218,N_13143,N_11020);
nand U15219 (N_15219,N_12167,N_14061);
or U15220 (N_15220,N_12728,N_12000);
xnor U15221 (N_15221,N_13882,N_12260);
nor U15222 (N_15222,N_10600,N_12360);
nor U15223 (N_15223,N_12242,N_14237);
and U15224 (N_15224,N_11158,N_12205);
xor U15225 (N_15225,N_14404,N_14319);
nor U15226 (N_15226,N_10391,N_11165);
or U15227 (N_15227,N_14942,N_12234);
xnor U15228 (N_15228,N_13937,N_13963);
or U15229 (N_15229,N_12509,N_12742);
nand U15230 (N_15230,N_10020,N_13100);
or U15231 (N_15231,N_10999,N_12441);
xor U15232 (N_15232,N_11745,N_13830);
xor U15233 (N_15233,N_12715,N_14406);
or U15234 (N_15234,N_13743,N_11030);
or U15235 (N_15235,N_14878,N_14747);
xnor U15236 (N_15236,N_13483,N_14527);
nand U15237 (N_15237,N_10217,N_12549);
and U15238 (N_15238,N_13771,N_13023);
nand U15239 (N_15239,N_10602,N_12423);
or U15240 (N_15240,N_14719,N_11930);
or U15241 (N_15241,N_12003,N_11633);
nor U15242 (N_15242,N_11532,N_12202);
xnor U15243 (N_15243,N_10986,N_10204);
nor U15244 (N_15244,N_10089,N_11383);
nand U15245 (N_15245,N_10625,N_12178);
xnor U15246 (N_15246,N_10723,N_13160);
nor U15247 (N_15247,N_10484,N_11150);
nand U15248 (N_15248,N_12404,N_12126);
xnor U15249 (N_15249,N_12977,N_13641);
nor U15250 (N_15250,N_14833,N_13759);
xor U15251 (N_15251,N_13086,N_10705);
nor U15252 (N_15252,N_14341,N_10789);
or U15253 (N_15253,N_13278,N_11176);
and U15254 (N_15254,N_11956,N_13946);
and U15255 (N_15255,N_13628,N_12435);
nor U15256 (N_15256,N_12631,N_14373);
nor U15257 (N_15257,N_13119,N_11518);
or U15258 (N_15258,N_13739,N_14672);
and U15259 (N_15259,N_14392,N_11107);
nand U15260 (N_15260,N_13108,N_10056);
xor U15261 (N_15261,N_12558,N_10225);
or U15262 (N_15262,N_14112,N_11679);
xor U15263 (N_15263,N_10021,N_13082);
nor U15264 (N_15264,N_10532,N_10877);
nor U15265 (N_15265,N_10109,N_13311);
and U15266 (N_15266,N_14854,N_11256);
and U15267 (N_15267,N_11626,N_10641);
nor U15268 (N_15268,N_12961,N_12225);
nand U15269 (N_15269,N_12466,N_11607);
xnor U15270 (N_15270,N_12111,N_14629);
nand U15271 (N_15271,N_14969,N_14845);
and U15272 (N_15272,N_12037,N_12287);
nor U15273 (N_15273,N_13610,N_14091);
nor U15274 (N_15274,N_10646,N_10659);
or U15275 (N_15275,N_11042,N_14523);
and U15276 (N_15276,N_12726,N_14530);
nand U15277 (N_15277,N_12251,N_14049);
or U15278 (N_15278,N_11145,N_11507);
or U15279 (N_15279,N_12935,N_10232);
xnor U15280 (N_15280,N_12725,N_11987);
xnor U15281 (N_15281,N_10845,N_10182);
nor U15282 (N_15282,N_13665,N_14499);
nand U15283 (N_15283,N_14079,N_13725);
and U15284 (N_15284,N_10678,N_12921);
and U15285 (N_15285,N_13213,N_11581);
nor U15286 (N_15286,N_13807,N_11371);
xor U15287 (N_15287,N_11596,N_14327);
xor U15288 (N_15288,N_10585,N_13790);
xnor U15289 (N_15289,N_12744,N_11017);
nand U15290 (N_15290,N_11719,N_11295);
nor U15291 (N_15291,N_10924,N_13742);
xor U15292 (N_15292,N_10966,N_14806);
nand U15293 (N_15293,N_12724,N_10437);
and U15294 (N_15294,N_11678,N_12622);
nor U15295 (N_15295,N_13316,N_14593);
and U15296 (N_15296,N_12446,N_10783);
or U15297 (N_15297,N_12910,N_14362);
xnor U15298 (N_15298,N_11340,N_11773);
or U15299 (N_15299,N_13146,N_14568);
nand U15300 (N_15300,N_14192,N_14172);
nand U15301 (N_15301,N_14184,N_10732);
nand U15302 (N_15302,N_10298,N_10317);
xor U15303 (N_15303,N_12236,N_12380);
xnor U15304 (N_15304,N_11102,N_13910);
or U15305 (N_15305,N_12066,N_13925);
nand U15306 (N_15306,N_14664,N_10922);
and U15307 (N_15307,N_10988,N_10766);
nand U15308 (N_15308,N_12313,N_11709);
nand U15309 (N_15309,N_14989,N_13840);
nand U15310 (N_15310,N_13902,N_11866);
nand U15311 (N_15311,N_13172,N_14216);
nor U15312 (N_15312,N_13248,N_14159);
and U15313 (N_15313,N_12782,N_10793);
and U15314 (N_15314,N_13034,N_13050);
xor U15315 (N_15315,N_13654,N_14577);
nand U15316 (N_15316,N_11192,N_12453);
nor U15317 (N_15317,N_11062,N_10906);
nor U15318 (N_15318,N_10138,N_13852);
or U15319 (N_15319,N_12253,N_13301);
xor U15320 (N_15320,N_12299,N_10088);
nor U15321 (N_15321,N_11119,N_13116);
xnor U15322 (N_15322,N_11226,N_10392);
and U15323 (N_15323,N_14567,N_10474);
and U15324 (N_15324,N_13235,N_11515);
nand U15325 (N_15325,N_10082,N_14718);
or U15326 (N_15326,N_12552,N_10653);
and U15327 (N_15327,N_11384,N_13021);
or U15328 (N_15328,N_13250,N_10008);
and U15329 (N_15329,N_13493,N_14587);
or U15330 (N_15330,N_12505,N_12760);
or U15331 (N_15331,N_11056,N_13028);
and U15332 (N_15332,N_11041,N_10655);
nor U15333 (N_15333,N_12323,N_14898);
nand U15334 (N_15334,N_13094,N_14221);
nand U15335 (N_15335,N_13621,N_12937);
and U15336 (N_15336,N_13747,N_10912);
nand U15337 (N_15337,N_12866,N_11774);
and U15338 (N_15338,N_10131,N_14710);
and U15339 (N_15339,N_12142,N_10398);
nand U15340 (N_15340,N_11482,N_11696);
or U15341 (N_15341,N_14111,N_10565);
and U15342 (N_15342,N_12581,N_14151);
and U15343 (N_15343,N_14098,N_14302);
xnor U15344 (N_15344,N_13726,N_14934);
xnor U15345 (N_15345,N_10343,N_11019);
and U15346 (N_15346,N_10037,N_11943);
and U15347 (N_15347,N_14285,N_10824);
and U15348 (N_15348,N_11270,N_11833);
and U15349 (N_15349,N_14343,N_10338);
nand U15350 (N_15350,N_14461,N_14213);
and U15351 (N_15351,N_13121,N_12856);
or U15352 (N_15352,N_10276,N_14101);
xnor U15353 (N_15353,N_11863,N_12256);
and U15354 (N_15354,N_13327,N_11267);
xor U15355 (N_15355,N_13285,N_14047);
and U15356 (N_15356,N_12162,N_12915);
and U15357 (N_15357,N_12709,N_11962);
or U15358 (N_15358,N_12132,N_10751);
xnor U15359 (N_15359,N_10471,N_13838);
and U15360 (N_15360,N_13355,N_12953);
or U15361 (N_15361,N_13753,N_10545);
xor U15362 (N_15362,N_10690,N_14561);
and U15363 (N_15363,N_12576,N_10324);
nand U15364 (N_15364,N_11422,N_14889);
or U15365 (N_15365,N_12095,N_10941);
nand U15366 (N_15366,N_10369,N_13229);
xor U15367 (N_15367,N_13745,N_12876);
nor U15368 (N_15368,N_14361,N_13573);
xor U15369 (N_15369,N_14246,N_12402);
nor U15370 (N_15370,N_11855,N_11793);
and U15371 (N_15371,N_11791,N_11724);
nor U15372 (N_15372,N_12702,N_14582);
and U15373 (N_15373,N_14090,N_13959);
nand U15374 (N_15374,N_11559,N_14043);
xnor U15375 (N_15375,N_10821,N_13353);
or U15376 (N_15376,N_13730,N_10520);
nor U15377 (N_15377,N_11718,N_11332);
nor U15378 (N_15378,N_12395,N_13603);
nor U15379 (N_15379,N_13844,N_14202);
or U15380 (N_15380,N_13164,N_10516);
or U15381 (N_15381,N_14475,N_13361);
nand U15382 (N_15382,N_10273,N_10361);
and U15383 (N_15383,N_11462,N_13369);
and U15384 (N_15384,N_14137,N_14456);
nand U15385 (N_15385,N_13916,N_11373);
or U15386 (N_15386,N_14663,N_11972);
nor U15387 (N_15387,N_12668,N_11474);
or U15388 (N_15388,N_12817,N_10657);
or U15389 (N_15389,N_14313,N_13841);
xor U15390 (N_15390,N_13499,N_10566);
nand U15391 (N_15391,N_12860,N_14991);
or U15392 (N_15392,N_11729,N_13110);
nor U15393 (N_15393,N_10431,N_12422);
nand U15394 (N_15394,N_12829,N_13038);
nand U15395 (N_15395,N_12704,N_12337);
and U15396 (N_15396,N_13474,N_14698);
or U15397 (N_15397,N_12461,N_13177);
nor U15398 (N_15398,N_11438,N_12941);
xor U15399 (N_15399,N_12547,N_10830);
and U15400 (N_15400,N_11419,N_12858);
nor U15401 (N_15401,N_11843,N_13436);
nand U15402 (N_15402,N_10255,N_12889);
xnor U15403 (N_15403,N_10077,N_13045);
nand U15404 (N_15404,N_10648,N_12462);
and U15405 (N_15405,N_14438,N_11363);
nor U15406 (N_15406,N_14035,N_11443);
or U15407 (N_15407,N_13703,N_14635);
or U15408 (N_15408,N_14376,N_11146);
and U15409 (N_15409,N_13903,N_12184);
or U15410 (N_15410,N_10910,N_12770);
nor U15411 (N_15411,N_12487,N_14225);
and U15412 (N_15412,N_10169,N_14867);
and U15413 (N_15413,N_10836,N_14424);
and U15414 (N_15414,N_11924,N_10064);
or U15415 (N_15415,N_14031,N_11327);
nand U15416 (N_15416,N_11921,N_10674);
xor U15417 (N_15417,N_12094,N_11242);
nand U15418 (N_15418,N_14838,N_10619);
xor U15419 (N_15419,N_14778,N_13862);
nor U15420 (N_15420,N_11320,N_12943);
nor U15421 (N_15421,N_11222,N_10993);
nand U15422 (N_15422,N_11348,N_14564);
nand U15423 (N_15423,N_10345,N_10592);
nand U15424 (N_15424,N_10923,N_14517);
nor U15425 (N_15425,N_11889,N_11733);
nor U15426 (N_15426,N_11105,N_12048);
or U15427 (N_15427,N_13630,N_14670);
and U15428 (N_15428,N_13998,N_12310);
nand U15429 (N_15429,N_11100,N_10557);
xnor U15430 (N_15430,N_11661,N_14762);
and U15431 (N_15431,N_12786,N_14542);
nand U15432 (N_15432,N_10531,N_12948);
or U15433 (N_15433,N_10442,N_14965);
or U15434 (N_15434,N_11321,N_11926);
and U15435 (N_15435,N_12143,N_14256);
nor U15436 (N_15436,N_10110,N_14684);
nor U15437 (N_15437,N_10253,N_14384);
or U15438 (N_15438,N_14791,N_10603);
nor U15439 (N_15439,N_12761,N_14544);
nand U15440 (N_15440,N_10665,N_11720);
xor U15441 (N_15441,N_14634,N_10573);
and U15442 (N_15442,N_12615,N_10584);
xnor U15443 (N_15443,N_11786,N_10835);
nor U15444 (N_15444,N_10661,N_11417);
or U15445 (N_15445,N_14708,N_14108);
xor U15446 (N_15446,N_11732,N_12322);
or U15447 (N_15447,N_11334,N_10543);
nor U15448 (N_15448,N_12827,N_10453);
or U15449 (N_15449,N_11436,N_10039);
nor U15450 (N_15450,N_14655,N_11091);
and U15451 (N_15451,N_13717,N_14220);
nor U15452 (N_15452,N_11768,N_10995);
nor U15453 (N_15453,N_14575,N_12654);
nor U15454 (N_15454,N_10294,N_11517);
nor U15455 (N_15455,N_14701,N_13869);
and U15456 (N_15456,N_12529,N_14686);
nand U15457 (N_15457,N_12204,N_14641);
xnor U15458 (N_15458,N_10792,N_10179);
nor U15459 (N_15459,N_10805,N_12619);
nor U15460 (N_15460,N_10380,N_13848);
nand U15461 (N_15461,N_13215,N_13450);
nand U15462 (N_15462,N_11654,N_13580);
xor U15463 (N_15463,N_11586,N_10165);
nand U15464 (N_15464,N_10362,N_12276);
xnor U15465 (N_15465,N_11021,N_12525);
or U15466 (N_15466,N_12607,N_13581);
xor U15467 (N_15467,N_13245,N_10272);
and U15468 (N_15468,N_10546,N_12179);
and U15469 (N_15469,N_12837,N_11263);
nand U15470 (N_15470,N_14441,N_13952);
nor U15471 (N_15471,N_14590,N_12389);
and U15472 (N_15472,N_13490,N_13468);
or U15473 (N_15473,N_10360,N_13105);
nand U15474 (N_15474,N_10203,N_14647);
nor U15475 (N_15475,N_12170,N_10574);
nand U15476 (N_15476,N_10292,N_14657);
nand U15477 (N_15477,N_13637,N_12769);
nand U15478 (N_15478,N_13693,N_12475);
or U15479 (N_15479,N_10081,N_11308);
or U15480 (N_15480,N_10019,N_11531);
nor U15481 (N_15481,N_13823,N_14687);
nand U15482 (N_15482,N_14074,N_10011);
nor U15483 (N_15483,N_13938,N_11990);
nor U15484 (N_15484,N_11913,N_13906);
xor U15485 (N_15485,N_12646,N_10727);
and U15486 (N_15486,N_14842,N_11160);
nand U15487 (N_15487,N_10880,N_12897);
nand U15488 (N_15488,N_10978,N_13762);
nor U15489 (N_15489,N_10628,N_12010);
and U15490 (N_15490,N_14180,N_14531);
nand U15491 (N_15491,N_14076,N_12028);
and U15492 (N_15492,N_11947,N_11702);
xnor U15493 (N_15493,N_13542,N_13428);
nor U15494 (N_15494,N_10314,N_12434);
nor U15495 (N_15495,N_11509,N_10833);
and U15496 (N_15496,N_11526,N_10873);
or U15497 (N_15497,N_10850,N_13210);
or U15498 (N_15498,N_10134,N_13484);
nand U15499 (N_15499,N_11841,N_12346);
nand U15500 (N_15500,N_11703,N_12078);
and U15501 (N_15501,N_11421,N_13756);
or U15502 (N_15502,N_12358,N_14469);
nand U15503 (N_15503,N_12677,N_11883);
and U15504 (N_15504,N_12972,N_14467);
or U15505 (N_15505,N_11471,N_11483);
or U15506 (N_15506,N_14179,N_12777);
xor U15507 (N_15507,N_11149,N_11023);
nand U15508 (N_15508,N_11434,N_13166);
nand U15509 (N_15509,N_11856,N_10463);
or U15510 (N_15510,N_11359,N_12147);
or U15511 (N_15511,N_10920,N_14829);
xnor U15512 (N_15512,N_12057,N_12384);
xnor U15513 (N_15513,N_12149,N_14696);
nand U15514 (N_15514,N_14535,N_10983);
or U15515 (N_15515,N_12873,N_11337);
and U15516 (N_15516,N_10583,N_10710);
and U15517 (N_15517,N_14849,N_10570);
nor U15518 (N_15518,N_12510,N_11639);
xnor U15519 (N_15519,N_10514,N_14676);
and U15520 (N_15520,N_12022,N_14546);
nor U15521 (N_15521,N_10215,N_12350);
or U15522 (N_15522,N_13261,N_13130);
and U15523 (N_15523,N_10527,N_12869);
and U15524 (N_15524,N_11298,N_11599);
and U15525 (N_15525,N_11424,N_14730);
xnor U15526 (N_15526,N_12474,N_12232);
nor U15527 (N_15527,N_10100,N_10996);
nor U15528 (N_15528,N_12512,N_12640);
xor U15529 (N_15529,N_14445,N_10580);
or U15530 (N_15530,N_14412,N_11961);
or U15531 (N_15531,N_14066,N_14087);
nor U15532 (N_15532,N_11191,N_13003);
and U15533 (N_15533,N_13257,N_10753);
nor U15534 (N_15534,N_12120,N_12691);
nor U15535 (N_15535,N_12351,N_11372);
nand U15536 (N_15536,N_10759,N_10156);
and U15537 (N_15537,N_11890,N_13206);
xnor U15538 (N_15538,N_12884,N_10430);
and U15539 (N_15539,N_10237,N_14737);
nand U15540 (N_15540,N_11430,N_14800);
nor U15541 (N_15541,N_10511,N_14015);
xnor U15542 (N_15542,N_13435,N_11074);
or U15543 (N_15543,N_11920,N_14608);
or U15544 (N_15544,N_11075,N_10427);
xnor U15545 (N_15545,N_12138,N_11668);
nor U15546 (N_15546,N_12818,N_10491);
and U15547 (N_15547,N_12840,N_11808);
nor U15548 (N_15548,N_10216,N_10210);
nor U15549 (N_15549,N_10414,N_14036);
nand U15550 (N_15550,N_13738,N_13999);
nor U15551 (N_15551,N_13063,N_10494);
xor U15552 (N_15552,N_14959,N_14295);
xnor U15553 (N_15553,N_12816,N_11764);
or U15554 (N_15554,N_14879,N_14363);
xnor U15555 (N_15555,N_14039,N_10889);
nand U15556 (N_15556,N_14451,N_10688);
xnor U15557 (N_15557,N_14848,N_11538);
xor U15558 (N_15558,N_12439,N_13374);
or U15559 (N_15559,N_13048,N_10519);
and U15560 (N_15560,N_11240,N_13377);
or U15561 (N_15561,N_10861,N_13977);
nand U15562 (N_15562,N_14462,N_14533);
nand U15563 (N_15563,N_12784,N_10501);
nor U15564 (N_15564,N_10413,N_12720);
xnor U15565 (N_15565,N_13636,N_10128);
nand U15566 (N_15566,N_10578,N_12574);
nand U15567 (N_15567,N_11052,N_13251);
or U15568 (N_15568,N_10240,N_14153);
nand U15569 (N_15569,N_10040,N_13181);
or U15570 (N_15570,N_11812,N_14987);
nor U15571 (N_15571,N_12708,N_12283);
or U15572 (N_15572,N_13964,N_11343);
and U15573 (N_15573,N_10868,N_10826);
xor U15574 (N_15574,N_11024,N_11958);
nand U15575 (N_15575,N_14133,N_11113);
and U15576 (N_15576,N_12975,N_12023);
nor U15577 (N_15577,N_13372,N_11649);
or U15578 (N_15578,N_13480,N_12130);
and U15579 (N_15579,N_14364,N_11083);
and U15580 (N_15580,N_14757,N_10016);
nor U15581 (N_15581,N_11201,N_11945);
or U15582 (N_15582,N_12220,N_11012);
or U15583 (N_15583,N_11859,N_11050);
xor U15584 (N_15584,N_10092,N_10954);
nand U15585 (N_15585,N_10669,N_14396);
and U15586 (N_15586,N_13047,N_11301);
nor U15587 (N_15587,N_10670,N_10250);
or U15588 (N_15588,N_14359,N_14435);
and U15589 (N_15589,N_10365,N_13201);
nor U15590 (N_15590,N_10699,N_11618);
nor U15591 (N_15591,N_13666,N_13315);
xnor U15592 (N_15592,N_14768,N_14749);
nor U15593 (N_15593,N_13587,N_14489);
nor U15594 (N_15594,N_13664,N_12671);
nor U15595 (N_15595,N_14086,N_12764);
or U15596 (N_15596,N_13676,N_14277);
nor U15597 (N_15597,N_12307,N_12917);
and U15598 (N_15598,N_13901,N_12732);
nand U15599 (N_15599,N_12849,N_12667);
nand U15600 (N_15600,N_10103,N_14513);
nand U15601 (N_15601,N_11876,N_13534);
or U15602 (N_15602,N_10544,N_11911);
and U15603 (N_15603,N_10624,N_12112);
and U15604 (N_15604,N_11631,N_11093);
xnor U15605 (N_15605,N_12268,N_12235);
or U15606 (N_15606,N_10781,N_10395);
nand U15607 (N_15607,N_12653,N_12985);
and U15608 (N_15608,N_10513,N_13917);
nand U15609 (N_15609,N_10310,N_11965);
xor U15610 (N_15610,N_12033,N_12410);
or U15611 (N_15611,N_10595,N_13357);
or U15612 (N_15612,N_14807,N_13658);
or U15613 (N_15613,N_13058,N_14583);
or U15614 (N_15614,N_13156,N_12052);
or U15615 (N_15615,N_10318,N_13027);
nor U15616 (N_15616,N_14464,N_12748);
xor U15617 (N_15617,N_12391,N_13449);
nand U15618 (N_15618,N_13191,N_10078);
xor U15619 (N_15619,N_10930,N_14715);
and U15620 (N_15620,N_10524,N_11617);
nand U15621 (N_15621,N_12246,N_10990);
or U15622 (N_15622,N_14139,N_13889);
nor U15623 (N_15623,N_14058,N_14443);
and U15624 (N_15624,N_10499,N_13036);
nand U15625 (N_15625,N_13184,N_13982);
and U15626 (N_15626,N_10319,N_14688);
nand U15627 (N_15627,N_14260,N_11609);
and U15628 (N_15628,N_13792,N_14745);
or U15629 (N_15629,N_10087,N_10946);
or U15630 (N_15630,N_11776,N_14656);
xnor U15631 (N_15631,N_11140,N_14181);
or U15632 (N_15632,N_12096,N_10243);
or U15633 (N_15633,N_14104,N_10508);
or U15634 (N_15634,N_14764,N_11864);
xnor U15635 (N_15635,N_13219,N_11246);
nand U15636 (N_15636,N_14621,N_10476);
or U15637 (N_15637,N_12187,N_14680);
xor U15638 (N_15638,N_10191,N_14006);
nor U15639 (N_15639,N_13934,N_12665);
nor U15640 (N_15640,N_14482,N_12859);
and U15641 (N_15641,N_14630,N_14189);
nand U15642 (N_15642,N_12097,N_10902);
or U15643 (N_15643,N_14563,N_10926);
and U15644 (N_15644,N_13077,N_14100);
and U15645 (N_15645,N_11783,N_11034);
or U15646 (N_15646,N_12751,N_11588);
or U15647 (N_15647,N_14899,N_12946);
nand U15648 (N_15648,N_14140,N_10523);
nand U15649 (N_15649,N_12329,N_13099);
nor U15650 (N_15650,N_11397,N_13865);
or U15651 (N_15651,N_12308,N_12880);
or U15652 (N_15652,N_11606,N_10937);
xnor U15653 (N_15653,N_12065,N_10416);
xnor U15654 (N_15654,N_10894,N_11707);
or U15655 (N_15655,N_14669,N_13434);
xnor U15656 (N_15656,N_10904,N_10720);
nand U15657 (N_15657,N_13575,N_11488);
nor U15658 (N_15658,N_11142,N_11877);
or U15659 (N_15659,N_11550,N_10183);
and U15660 (N_15660,N_12309,N_13719);
and U15661 (N_15661,N_14970,N_13333);
or U15662 (N_15662,N_10997,N_12409);
and U15663 (N_15663,N_14041,N_12006);
nor U15664 (N_15664,N_10073,N_13853);
nand U15665 (N_15665,N_10788,N_14826);
nor U15666 (N_15666,N_10466,N_12734);
nand U15667 (N_15667,N_14892,N_14099);
nand U15668 (N_15668,N_10948,N_12796);
xnor U15669 (N_15669,N_14871,N_14146);
or U15670 (N_15670,N_14619,N_12980);
nand U15671 (N_15671,N_12438,N_13897);
nor U15672 (N_15672,N_14483,N_12228);
or U15673 (N_15673,N_13197,N_12020);
xnor U15674 (N_15674,N_13527,N_14600);
or U15675 (N_15675,N_14685,N_13515);
xor U15676 (N_15676,N_11805,N_10473);
and U15677 (N_15677,N_12666,N_12506);
and U15678 (N_15678,N_14816,N_12923);
nor U15679 (N_15679,N_13292,N_13103);
and U15680 (N_15680,N_14736,N_12743);
and U15681 (N_15681,N_11591,N_11551);
nor U15682 (N_15682,N_14082,N_14095);
nor U15683 (N_15683,N_13295,N_10662);
and U15684 (N_15684,N_11306,N_14819);
xnor U15685 (N_15685,N_11470,N_13639);
xnor U15686 (N_15686,N_11840,N_10115);
nand U15687 (N_15687,N_14233,N_12145);
nor U15688 (N_15688,N_13283,N_12767);
xnor U15689 (N_15689,N_14311,N_14155);
nor U15690 (N_15690,N_11896,N_14721);
nor U15691 (N_15691,N_11184,N_14760);
or U15692 (N_15692,N_11031,N_13055);
and U15693 (N_15693,N_14485,N_12277);
or U15694 (N_15694,N_14584,N_14667);
nand U15695 (N_15695,N_13682,N_12163);
and U15696 (N_15696,N_14134,N_10486);
or U15697 (N_15697,N_10495,N_14261);
nor U15698 (N_15698,N_14742,N_14380);
and U15699 (N_15699,N_14350,N_14627);
or U15700 (N_15700,N_14321,N_12991);
nor U15701 (N_15701,N_10837,N_10778);
xor U15702 (N_15702,N_13422,N_10139);
xnor U15703 (N_15703,N_13565,N_13243);
xor U15704 (N_15704,N_14303,N_12104);
and U15705 (N_15705,N_11117,N_14008);
xnor U15706 (N_15706,N_13424,N_11328);
xor U15707 (N_15707,N_14228,N_13208);
xor U15708 (N_15708,N_11345,N_11563);
or U15709 (N_15709,N_10745,N_14241);
and U15710 (N_15710,N_12736,N_10377);
xnor U15711 (N_15711,N_11459,N_11174);
nand U15712 (N_15712,N_12540,N_10972);
nand U15713 (N_15713,N_11888,N_13699);
xor U15714 (N_15714,N_10963,N_11759);
xnor U15715 (N_15715,N_13660,N_10776);
and U15716 (N_15716,N_12182,N_10321);
and U15717 (N_15717,N_13007,N_14042);
or U15718 (N_15718,N_14916,N_10454);
nand U15719 (N_15719,N_12074,N_10287);
xor U15720 (N_15720,N_13705,N_13777);
or U15721 (N_15721,N_12129,N_11029);
or U15722 (N_15722,N_12301,N_11623);
nor U15723 (N_15723,N_11828,N_12321);
nand U15724 (N_15724,N_14733,N_14811);
or U15725 (N_15725,N_13117,N_14349);
nor U15726 (N_15726,N_13124,N_14858);
and U15727 (N_15727,N_13622,N_10677);
nand U15728 (N_15728,N_13000,N_14580);
and U15729 (N_15729,N_13976,N_13796);
xor U15730 (N_15730,N_12488,N_13498);
nor U15731 (N_15731,N_13202,N_13887);
and U15732 (N_15732,N_13576,N_10747);
nor U15733 (N_15733,N_13109,N_10440);
or U15734 (N_15734,N_12661,N_14940);
nor U15735 (N_15735,N_14385,N_10224);
nor U15736 (N_15736,N_12452,N_14840);
nor U15737 (N_15737,N_13004,N_10775);
or U15738 (N_15738,N_12250,N_12971);
xor U15739 (N_15739,N_11739,N_12226);
and U15740 (N_15740,N_10932,N_11455);
nor U15741 (N_15741,N_14425,N_13867);
nand U15742 (N_15742,N_12545,N_12804);
xor U15743 (N_15743,N_12832,N_14480);
nor U15744 (N_15744,N_10612,N_13440);
xnor U15745 (N_15745,N_14573,N_11374);
and U15746 (N_15746,N_13800,N_12633);
or U15747 (N_15747,N_13571,N_14196);
and U15748 (N_15748,N_14067,N_14594);
xor U15749 (N_15749,N_10193,N_10451);
xnor U15750 (N_15750,N_13371,N_14129);
or U15751 (N_15751,N_13864,N_12357);
nor U15752 (N_15752,N_10332,N_14556);
nand U15753 (N_15753,N_14881,N_11281);
or U15754 (N_15754,N_12685,N_10563);
xor U15755 (N_15755,N_12537,N_14453);
nand U15756 (N_15756,N_12364,N_12593);
nand U15757 (N_15757,N_12419,N_14825);
xor U15758 (N_15758,N_12503,N_11442);
and U15759 (N_15759,N_12318,N_11644);
or U15760 (N_15760,N_10146,N_13231);
and U15761 (N_15761,N_11562,N_14200);
xnor U15762 (N_15762,N_12824,N_11068);
nor U15763 (N_15763,N_14992,N_10804);
nor U15764 (N_15764,N_11820,N_14941);
xor U15765 (N_15765,N_13984,N_12519);
or U15766 (N_15766,N_11971,N_14801);
xor U15767 (N_15767,N_13096,N_14342);
nor U15768 (N_15768,N_11792,N_14660);
xor U15769 (N_15769,N_10246,N_13989);
nand U15770 (N_15770,N_13948,N_11404);
nand U15771 (N_15771,N_11974,N_14518);
and U15772 (N_15772,N_12393,N_11447);
nor U15773 (N_15773,N_12655,N_13463);
xor U15774 (N_15774,N_12627,N_13709);
or U15775 (N_15775,N_10279,N_14787);
nand U15776 (N_15776,N_11695,N_13317);
nand U15777 (N_15777,N_10679,N_10701);
and U15778 (N_15778,N_14997,N_12909);
or U15779 (N_15779,N_13801,N_13360);
or U15780 (N_15780,N_10013,N_14059);
or U15781 (N_15781,N_13854,N_12368);
nor U15782 (N_15782,N_12390,N_14907);
and U15783 (N_15783,N_14020,N_11121);
and U15784 (N_15784,N_10251,N_12284);
and U15785 (N_15785,N_10848,N_11460);
xnor U15786 (N_15786,N_10504,N_11403);
xnor U15787 (N_15787,N_11714,N_14886);
and U15788 (N_15788,N_14032,N_10840);
xor U15789 (N_15789,N_11845,N_13803);
nor U15790 (N_15790,N_12154,N_12151);
or U15791 (N_15791,N_12934,N_14746);
nor U15792 (N_15792,N_10525,N_12885);
and U15793 (N_15793,N_13927,N_12737);
xor U15794 (N_15794,N_10807,N_14665);
and U15795 (N_15795,N_12984,N_13165);
nor U15796 (N_15796,N_12706,N_14869);
xor U15797 (N_15797,N_13167,N_12541);
nor U15798 (N_15798,N_13851,N_14397);
or U15799 (N_15799,N_11565,N_13267);
nand U15800 (N_15800,N_14492,N_10396);
xnor U15801 (N_15801,N_11814,N_12514);
or U15802 (N_15802,N_14248,N_11975);
nor U15803 (N_15803,N_13735,N_10664);
xor U15804 (N_15804,N_11053,N_12511);
xnor U15805 (N_15805,N_10639,N_14675);
xor U15806 (N_15806,N_11469,N_10576);
xnor U15807 (N_15807,N_13920,N_11035);
and U15808 (N_15808,N_13546,N_13557);
and U15809 (N_15809,N_13857,N_11795);
and U15810 (N_15810,N_12814,N_12166);
nand U15811 (N_15811,N_11300,N_10921);
nand U15812 (N_15812,N_11463,N_10060);
nand U15813 (N_15813,N_14379,N_12939);
nand U15814 (N_15814,N_14559,N_11173);
or U15815 (N_15815,N_12291,N_10616);
nand U15816 (N_15816,N_14975,N_13260);
and U15817 (N_15817,N_14063,N_14813);
nand U15818 (N_15818,N_14332,N_10419);
nor U15819 (N_15819,N_13423,N_12442);
xnor U15820 (N_15820,N_14545,N_11018);
or U15821 (N_15821,N_12920,N_12902);
xnor U15822 (N_15822,N_11060,N_11590);
xor U15823 (N_15823,N_14118,N_11660);
xnor U15824 (N_15824,N_14979,N_14974);
xnor U15825 (N_15825,N_11457,N_12681);
and U15826 (N_15826,N_12378,N_13481);
xnor U15827 (N_15827,N_12940,N_12944);
nand U15828 (N_15828,N_12739,N_14457);
xor U15829 (N_15829,N_13005,N_10614);
nand U15830 (N_15830,N_13710,N_10634);
or U15831 (N_15831,N_14274,N_12602);
nand U15832 (N_15832,N_11147,N_12850);
xor U15833 (N_15833,N_12618,N_11078);
and U15834 (N_15834,N_10541,N_10949);
nand U15835 (N_15835,N_14741,N_14169);
and U15836 (N_15836,N_10187,N_12707);
nor U15837 (N_15837,N_10444,N_12195);
xnor U15838 (N_15838,N_11016,N_14356);
nand U15839 (N_15839,N_14788,N_13821);
or U15840 (N_15840,N_14748,N_14446);
nand U15841 (N_15841,N_11804,N_10327);
nand U15842 (N_15842,N_14692,N_11401);
and U15843 (N_15843,N_12161,N_12408);
xor U15844 (N_15844,N_12089,N_14860);
and U15845 (N_15845,N_14045,N_12123);
xor U15846 (N_15846,N_11037,N_10185);
xnor U15847 (N_15847,N_10897,N_13894);
xor U15848 (N_15848,N_10663,N_11072);
nand U15849 (N_15849,N_12491,N_13523);
or U15850 (N_15850,N_14064,N_10892);
nand U15851 (N_15851,N_14930,N_10098);
nor U15852 (N_15852,N_11620,N_14423);
and U15853 (N_15853,N_11441,N_12054);
or U15854 (N_15854,N_10964,N_13950);
and U15855 (N_15855,N_10643,N_13528);
and U15856 (N_15856,N_13438,N_11022);
and U15857 (N_15857,N_11602,N_12752);
nor U15858 (N_15858,N_10291,N_11275);
nor U15859 (N_15859,N_13328,N_10236);
nand U15860 (N_15860,N_10974,N_14334);
or U15861 (N_15861,N_11453,N_13137);
or U15862 (N_15862,N_12272,N_12675);
or U15863 (N_15863,N_14883,N_12219);
nand U15864 (N_15864,N_11027,N_14508);
or U15865 (N_15865,N_12883,N_11431);
xor U15866 (N_15866,N_11155,N_11991);
xnor U15867 (N_15867,N_10241,N_14494);
or U15868 (N_15868,N_14943,N_10180);
nand U15869 (N_15869,N_10124,N_11428);
xnor U15870 (N_15870,N_13880,N_11662);
or U15871 (N_15871,N_13768,N_12172);
and U15872 (N_15872,N_14851,N_14936);
xor U15873 (N_15873,N_12997,N_11756);
nor U15874 (N_15874,N_11797,N_13242);
xor U15875 (N_15875,N_11749,N_13849);
xor U15876 (N_15876,N_11073,N_12407);
nor U15877 (N_15877,N_13304,N_12741);
and U15878 (N_15878,N_13627,N_11494);
nor U15879 (N_15879,N_14013,N_12678);
xor U15880 (N_15880,N_14501,N_13395);
or U15881 (N_15881,N_11276,N_14521);
nor U15882 (N_15882,N_13026,N_10105);
nand U15883 (N_15883,N_14937,N_11868);
xnor U15884 (N_15884,N_10893,N_11164);
nor U15885 (N_15885,N_10582,N_13885);
xnor U15886 (N_15886,N_11985,N_10282);
nor U15887 (N_15887,N_12521,N_12485);
and U15888 (N_15888,N_13269,N_12614);
nand U15889 (N_15889,N_13277,N_13625);
nand U15890 (N_15890,N_10827,N_10722);
xor U15891 (N_15891,N_13831,N_10304);
or U15892 (N_15892,N_12297,N_11346);
nand U15893 (N_15893,N_14652,N_11592);
nand U15894 (N_15894,N_10459,N_12382);
nand U15895 (N_15895,N_14432,N_13347);
nand U15896 (N_15896,N_13037,N_10724);
nor U15897 (N_15897,N_12669,N_12247);
nand U15898 (N_15898,N_10957,N_11489);
xor U15899 (N_15899,N_10606,N_11344);
nand U15900 (N_15900,N_12766,N_11688);
nand U15901 (N_15901,N_13516,N_14348);
nor U15902 (N_15902,N_10229,N_10729);
xnor U15903 (N_15903,N_12798,N_10895);
or U15904 (N_15904,N_13981,N_12918);
nor U15905 (N_15905,N_10465,N_14252);
or U15906 (N_15906,N_13017,N_11377);
nor U15907 (N_15907,N_11594,N_11934);
xor U15908 (N_15908,N_13645,N_14836);
and U15909 (N_15909,N_12212,N_11241);
xnor U15910 (N_15910,N_12617,N_13893);
xor U15911 (N_15911,N_14157,N_11156);
nand U15912 (N_15912,N_10389,N_10015);
or U15913 (N_15913,N_10953,N_10706);
xor U15914 (N_15914,N_11364,N_11225);
xnor U15915 (N_15915,N_13539,N_10388);
and U15916 (N_15916,N_14312,N_14442);
and U15917 (N_15917,N_14300,N_14403);
nor U15918 (N_15918,N_11516,N_12535);
xnor U15919 (N_15919,N_10239,N_14037);
xnor U15920 (N_15920,N_12083,N_13624);
nor U15921 (N_15921,N_10691,N_10685);
or U15922 (N_15922,N_12269,N_12561);
nor U15923 (N_15923,N_11352,N_14276);
xor U15924 (N_15924,N_13509,N_14765);
nand U15925 (N_15925,N_11635,N_10323);
and U15926 (N_15926,N_12749,N_11893);
xor U15927 (N_15927,N_14344,N_13115);
nand U15928 (N_15928,N_13362,N_12926);
nor U15929 (N_15929,N_10554,N_12312);
and U15930 (N_15930,N_10053,N_12201);
xor U15931 (N_15931,N_11082,N_14609);
or U15932 (N_15932,N_11170,N_11977);
nand U15933 (N_15933,N_13049,N_12701);
xnor U15934 (N_15934,N_12938,N_13313);
nand U15935 (N_15935,N_13106,N_12156);
nand U15936 (N_15936,N_13749,N_13655);
xor U15937 (N_15937,N_12261,N_10461);
and U15938 (N_15938,N_13198,N_14847);
nor U15939 (N_15939,N_12610,N_14234);
nor U15940 (N_15940,N_10355,N_10915);
xor U15941 (N_15941,N_12007,N_13590);
nand U15942 (N_15942,N_13700,N_10797);
nor U15943 (N_15943,N_14863,N_10284);
nor U15944 (N_15944,N_13180,N_14324);
nand U15945 (N_15945,N_14779,N_12630);
and U15946 (N_15946,N_14360,N_11912);
xnor U15947 (N_15947,N_13512,N_14428);
nand U15948 (N_15948,N_10968,N_11186);
nand U15949 (N_15949,N_13114,N_11008);
nor U15950 (N_15950,N_11725,N_14212);
xnor U15951 (N_15951,N_11541,N_10927);
and U15952 (N_15952,N_12047,N_14913);
nand U15953 (N_15953,N_13479,N_12468);
xor U15954 (N_15954,N_11433,N_12998);
nor U15955 (N_15955,N_10671,N_12306);
and U15956 (N_15956,N_14268,N_13545);
nor U15957 (N_15957,N_12427,N_14810);
xnor U15958 (N_15958,N_14106,N_11941);
nand U15959 (N_15959,N_14625,N_13895);
or U15960 (N_15960,N_11875,N_11342);
nand U15961 (N_15961,N_12118,N_14251);
or U15962 (N_15962,N_14281,N_13227);
and U15963 (N_15963,N_11650,N_10756);
xor U15964 (N_15964,N_12044,N_14644);
and U15965 (N_15965,N_11385,N_10931);
xnor U15966 (N_15966,N_12173,N_11838);
or U15967 (N_15967,N_13111,N_11787);
nor U15968 (N_15968,N_13988,N_12069);
nand U15969 (N_15969,N_13615,N_12585);
nand U15970 (N_15970,N_13586,N_13737);
nor U15971 (N_15971,N_13960,N_11183);
or U15972 (N_15972,N_10816,N_12136);
nor U15973 (N_15973,N_11878,N_10564);
or U15974 (N_15974,N_13253,N_11852);
nor U15975 (N_15975,N_13716,N_12797);
nor U15976 (N_15976,N_14182,N_13548);
or U15977 (N_15977,N_13644,N_11261);
and U15978 (N_15978,N_10509,N_11904);
or U15979 (N_15979,N_11521,N_11712);
nand U15980 (N_15980,N_12449,N_10708);
nand U15981 (N_15981,N_10743,N_13672);
nand U15982 (N_15982,N_11303,N_10366);
nand U15983 (N_15983,N_12406,N_12628);
nor U15984 (N_15984,N_11540,N_11399);
or U15985 (N_15985,N_11135,N_11040);
and U15986 (N_15986,N_13379,N_14596);
nor U15987 (N_15987,N_14977,N_11816);
and U15988 (N_15988,N_13600,N_14386);
and U15989 (N_15989,N_11988,N_10808);
xor U15990 (N_15990,N_10967,N_12543);
nand U15991 (N_15991,N_14250,N_14771);
and U15992 (N_15992,N_10887,N_10478);
and U15993 (N_15993,N_11089,N_14919);
nand U15994 (N_15994,N_12016,N_12353);
nand U15995 (N_15995,N_12638,N_12032);
or U15996 (N_15996,N_12241,N_10363);
nor U15997 (N_15997,N_10112,N_14306);
or U15998 (N_15998,N_13971,N_11857);
xnor U15999 (N_15999,N_12077,N_13335);
xor U16000 (N_16000,N_14383,N_12682);
nor U16001 (N_16001,N_10280,N_12262);
and U16002 (N_16002,N_13419,N_13089);
and U16003 (N_16003,N_12155,N_14078);
nor U16004 (N_16004,N_14818,N_12626);
nand U16005 (N_16005,N_10132,N_12305);
and U16006 (N_16006,N_13670,N_11185);
and U16007 (N_16007,N_10432,N_12694);
nor U16008 (N_16008,N_11873,N_13403);
xnor U16009 (N_16009,N_13322,N_11498);
or U16010 (N_16010,N_12218,N_13300);
nand U16011 (N_16011,N_11561,N_13947);
nand U16012 (N_16012,N_14177,N_11099);
or U16013 (N_16013,N_11009,N_12050);
and U16014 (N_16014,N_14171,N_11473);
nand U16015 (N_16015,N_14290,N_13727);
nor U16016 (N_16016,N_13983,N_11286);
nor U16017 (N_16017,N_11524,N_12068);
and U16018 (N_16018,N_12870,N_14900);
or U16019 (N_16019,N_13176,N_10769);
xor U16020 (N_16020,N_14585,N_11229);
nor U16021 (N_16021,N_11508,N_12444);
xnor U16022 (N_16022,N_14603,N_13958);
nand U16023 (N_16023,N_14183,N_13723);
xor U16024 (N_16024,N_11955,N_13426);
and U16025 (N_16025,N_14448,N_12459);
nand U16026 (N_16026,N_12564,N_13462);
or U16027 (N_16027,N_13162,N_11477);
and U16028 (N_16028,N_10309,N_12637);
xor U16029 (N_16029,N_14463,N_10802);
or U16030 (N_16030,N_13558,N_11476);
xor U16031 (N_16031,N_10341,N_14422);
or U16032 (N_16032,N_14330,N_11693);
nor U16033 (N_16033,N_10443,N_14444);
nor U16034 (N_16034,N_10438,N_13607);
nor U16035 (N_16035,N_14170,N_14094);
xor U16036 (N_16036,N_14516,N_12504);
nand U16037 (N_16037,N_13915,N_12051);
xor U16038 (N_16038,N_13183,N_11067);
xnor U16039 (N_16039,N_14612,N_11694);
nor U16040 (N_16040,N_12756,N_12625);
and U16041 (N_16041,N_12113,N_11730);
nand U16042 (N_16042,N_14387,N_10260);
nand U16043 (N_16043,N_11556,N_12546);
and U16044 (N_16044,N_14639,N_13951);
xor U16045 (N_16045,N_12379,N_12258);
nor U16046 (N_16046,N_11090,N_14345);
nand U16047 (N_16047,N_14823,N_12616);
xor U16048 (N_16048,N_14691,N_13011);
and U16049 (N_16049,N_13870,N_11612);
or U16050 (N_16050,N_10962,N_13453);
or U16051 (N_16051,N_12819,N_11642);
and U16052 (N_16052,N_13349,N_14549);
or U16053 (N_16053,N_14022,N_13861);
or U16054 (N_16054,N_14870,N_12335);
xnor U16055 (N_16055,N_11175,N_11218);
and U16056 (N_16056,N_14822,N_14658);
xnor U16057 (N_16057,N_14352,N_14188);
nor U16058 (N_16058,N_11582,N_14722);
nor U16059 (N_16059,N_13708,N_13380);
or U16060 (N_16060,N_14754,N_13334);
xor U16061 (N_16061,N_13366,N_12865);
nand U16062 (N_16062,N_11335,N_10166);
nor U16063 (N_16063,N_14650,N_12995);
nand U16064 (N_16064,N_13170,N_13554);
nor U16065 (N_16065,N_14034,N_11500);
and U16066 (N_16066,N_12019,N_13221);
nor U16067 (N_16067,N_12343,N_10375);
nand U16068 (N_16068,N_10761,N_11766);
nand U16069 (N_16069,N_13284,N_14273);
nand U16070 (N_16070,N_12043,N_11674);
nand U16071 (N_16071,N_13846,N_13185);
nand U16072 (N_16072,N_11126,N_12810);
or U16073 (N_16073,N_12191,N_13129);
nand U16074 (N_16074,N_10734,N_12430);
nand U16075 (N_16075,N_14928,N_11354);
xor U16076 (N_16076,N_12314,N_12252);
xor U16077 (N_16077,N_12958,N_10740);
nand U16078 (N_16078,N_13318,N_14541);
and U16079 (N_16079,N_13266,N_12566);
nor U16080 (N_16080,N_11775,N_14374);
nor U16081 (N_16081,N_14646,N_11981);
and U16082 (N_16082,N_12060,N_14926);
or U16083 (N_16083,N_10036,N_13520);
and U16084 (N_16084,N_11571,N_10561);
xnor U16085 (N_16085,N_11554,N_10457);
xor U16086 (N_16086,N_12746,N_10046);
or U16087 (N_16087,N_11392,N_14693);
nor U16088 (N_16088,N_10145,N_10029);
or U16089 (N_16089,N_14150,N_12624);
nor U16090 (N_16090,N_14011,N_10858);
nand U16091 (N_16091,N_12490,N_14507);
and U16092 (N_16092,N_12964,N_10551);
and U16093 (N_16093,N_12979,N_14803);
or U16094 (N_16094,N_12649,N_14707);
nand U16095 (N_16095,N_14266,N_12963);
or U16096 (N_16096,N_10693,N_10617);
nand U16097 (N_16097,N_12875,N_10881);
nor U16098 (N_16098,N_12515,N_10333);
xor U16099 (N_16099,N_12639,N_13298);
and U16100 (N_16100,N_10530,N_13290);
nor U16101 (N_16101,N_12344,N_12534);
xor U16102 (N_16102,N_11692,N_11901);
xor U16103 (N_16103,N_10611,N_14040);
nand U16104 (N_16104,N_11163,N_12952);
or U16105 (N_16105,N_13272,N_10143);
or U16106 (N_16106,N_12304,N_14756);
xnor U16107 (N_16107,N_11885,N_10133);
xor U16108 (N_16108,N_10487,N_11049);
nor U16109 (N_16109,N_10518,N_11199);
and U16110 (N_16110,N_10865,N_11497);
nor U16111 (N_16111,N_14558,N_11254);
nor U16112 (N_16112,N_12575,N_13505);
xor U16113 (N_16113,N_10249,N_10752);
nor U16114 (N_16114,N_13421,N_12092);
xnor U16115 (N_16115,N_11123,N_14586);
xnor U16116 (N_16116,N_12255,N_12542);
nand U16117 (N_16117,N_13979,N_14703);
nor U16118 (N_16118,N_13519,N_12562);
and U16119 (N_16119,N_14767,N_14025);
nor U16120 (N_16120,N_14119,N_13406);
nand U16121 (N_16121,N_10917,N_10831);
or U16122 (N_16122,N_10507,N_14632);
nor U16123 (N_16123,N_10876,N_13299);
nor U16124 (N_16124,N_11624,N_14514);
or U16125 (N_16125,N_14211,N_10571);
or U16126 (N_16126,N_11608,N_13510);
or U16127 (N_16127,N_12592,N_14859);
or U16128 (N_16128,N_12418,N_12703);
or U16129 (N_16129,N_10980,N_11288);
and U16130 (N_16130,N_11851,N_12611);
nand U16131 (N_16131,N_13415,N_10689);
nand U16132 (N_16132,N_14714,N_13455);
xnor U16133 (N_16133,N_11407,N_13256);
nor U16134 (N_16134,N_13513,N_14935);
nor U16135 (N_16135,N_12855,N_14752);
nand U16136 (N_16136,N_10632,N_11744);
nand U16137 (N_16137,N_13793,N_10528);
or U16138 (N_16138,N_13002,N_10399);
and U16139 (N_16139,N_13040,N_14618);
and U16140 (N_16140,N_11865,N_14776);
nand U16141 (N_16141,N_10506,N_10270);
nor U16142 (N_16142,N_10233,N_13836);
and U16143 (N_16143,N_13400,N_14607);
nor U16144 (N_16144,N_11084,N_13271);
and U16145 (N_16145,N_12100,N_14540);
xor U16146 (N_16146,N_12080,N_12279);
nand U16147 (N_16147,N_12300,N_13697);
or U16148 (N_16148,N_12500,N_11637);
xor U16149 (N_16149,N_11449,N_14168);
or U16150 (N_16150,N_12947,N_11426);
nand U16151 (N_16151,N_13721,N_12341);
and U16152 (N_16152,N_11743,N_11903);
and U16153 (N_16153,N_11272,N_11220);
nor U16154 (N_16154,N_11928,N_11915);
and U16155 (N_16155,N_10533,N_12388);
xor U16156 (N_16156,N_10106,N_11755);
xnor U16157 (N_16157,N_14016,N_11706);
or U16158 (N_16158,N_14995,N_11997);
nor U16159 (N_16159,N_10422,N_11728);
xor U16160 (N_16160,N_10434,N_10556);
nor U16161 (N_16161,N_12570,N_14224);
and U16162 (N_16162,N_10762,N_12397);
xor U16163 (N_16163,N_14550,N_14053);
xnor U16164 (N_16164,N_10860,N_11827);
nand U16165 (N_16165,N_13544,N_11378);
nand U16166 (N_16166,N_14529,N_14486);
nor U16167 (N_16167,N_10289,N_12989);
nand U16168 (N_16168,N_11051,N_14966);
xnor U16169 (N_16169,N_13559,N_12890);
and U16170 (N_16170,N_11738,N_12900);
nand U16171 (N_16171,N_11916,N_12927);
and U16172 (N_16172,N_12290,N_14242);
or U16173 (N_16173,N_12718,N_11512);
and U16174 (N_16174,N_10329,N_13452);
and U16175 (N_16175,N_10080,N_13370);
or U16176 (N_16176,N_14500,N_13629);
nor U16177 (N_16177,N_13459,N_14128);
xnor U16178 (N_16178,N_14065,N_13154);
nor U16179 (N_16179,N_11159,N_10464);
or U16180 (N_16180,N_12013,N_10108);
nor U16181 (N_16181,N_11652,N_11528);
and U16182 (N_16182,N_13204,N_11318);
xnor U16183 (N_16183,N_12538,N_12580);
nor U16184 (N_16184,N_12951,N_11966);
or U16185 (N_16185,N_13652,N_10736);
or U16186 (N_16186,N_12658,N_11347);
and U16187 (N_16187,N_11291,N_14953);
nor U16188 (N_16188,N_13780,N_14897);
or U16189 (N_16189,N_10152,N_14610);
and U16190 (N_16190,N_13653,N_12071);
nor U16191 (N_16191,N_12275,N_14455);
nand U16192 (N_16192,N_13015,N_13923);
and U16193 (N_16193,N_13543,N_11669);
or U16194 (N_16194,N_11627,N_14487);
nor U16195 (N_16195,N_10048,N_10660);
nor U16196 (N_16196,N_14077,N_11762);
nand U16197 (N_16197,N_11953,N_14856);
nor U16198 (N_16198,N_10119,N_13132);
xor U16199 (N_16199,N_10405,N_11231);
and U16200 (N_16200,N_10994,N_11905);
or U16201 (N_16201,N_12854,N_13524);
or U16202 (N_16202,N_11080,N_11491);
and U16203 (N_16203,N_14659,N_13309);
nand U16204 (N_16204,N_14967,N_10050);
nand U16205 (N_16205,N_13553,N_12898);
nor U16206 (N_16206,N_11326,N_12755);
and U16207 (N_16207,N_10859,N_10231);
nor U16208 (N_16208,N_11954,N_10055);
or U16209 (N_16209,N_11874,N_14476);
or U16210 (N_16210,N_14792,N_11922);
xnor U16211 (N_16211,N_10950,N_14739);
nand U16212 (N_16212,N_14240,N_10975);
nand U16213 (N_16213,N_12231,N_10247);
or U16214 (N_16214,N_10194,N_12930);
or U16215 (N_16215,N_14337,N_10320);
nand U16216 (N_16216,N_10730,N_14613);
nand U16217 (N_16217,N_10741,N_12015);
or U16218 (N_16218,N_13112,N_13572);
xor U16219 (N_16219,N_14437,N_12609);
nand U16220 (N_16220,N_12676,N_14798);
or U16221 (N_16221,N_14834,N_13626);
and U16222 (N_16222,N_13363,N_12176);
xor U16223 (N_16223,N_12278,N_14391);
nor U16224 (N_16224,N_14275,N_12465);
or U16225 (N_16225,N_14459,N_14088);
xor U16226 (N_16226,N_14410,N_14981);
xnor U16227 (N_16227,N_10770,N_11110);
nor U16228 (N_16228,N_12548,N_14877);
and U16229 (N_16229,N_10505,N_11233);
and U16230 (N_16230,N_10998,N_13503);
or U16231 (N_16231,N_14050,N_13384);
nor U16232 (N_16232,N_11545,N_10346);
and U16233 (N_16233,N_10286,N_14294);
nand U16234 (N_16234,N_11092,N_12976);
xor U16235 (N_16235,N_14167,N_11789);
nand U16236 (N_16236,N_11949,N_13997);
or U16237 (N_16237,N_14857,N_14068);
nor U16238 (N_16238,N_14257,N_10951);
and U16239 (N_16239,N_10559,N_10267);
xnor U16240 (N_16240,N_13681,N_14963);
or U16241 (N_16241,N_12194,N_14191);
or U16242 (N_16242,N_14732,N_11168);
nand U16243 (N_16243,N_12904,N_13032);
nand U16244 (N_16244,N_10572,N_13704);
xor U16245 (N_16245,N_11255,N_12134);
xnor U16246 (N_16246,N_14651,N_14335);
and U16247 (N_16247,N_12799,N_13305);
xnor U16248 (N_16248,N_11807,N_11583);
xor U16249 (N_16249,N_14591,N_12747);
nand U16250 (N_16250,N_14920,N_12334);
and U16251 (N_16251,N_13420,N_12879);
xnor U16252 (N_16252,N_11390,N_13409);
xor U16253 (N_16253,N_12785,N_13365);
xnor U16254 (N_16254,N_14931,N_10339);
and U16255 (N_16255,N_14548,N_11269);
nand U16256 (N_16256,N_14002,N_12636);
xor U16257 (N_16257,N_14852,N_10598);
nor U16258 (N_16258,N_13648,N_10900);
xor U16259 (N_16259,N_11558,N_12414);
or U16260 (N_16260,N_12070,N_14908);
nand U16261 (N_16261,N_10086,N_14579);
and U16262 (N_16262,N_12029,N_10023);
and U16263 (N_16263,N_10801,N_13228);
xor U16264 (N_16264,N_13731,N_12486);
or U16265 (N_16265,N_14543,N_14204);
and U16266 (N_16266,N_14595,N_12530);
nor U16267 (N_16267,N_12222,N_10230);
xor U16268 (N_16268,N_10174,N_13057);
nor U16269 (N_16269,N_14532,N_11043);
nor U16270 (N_16270,N_13312,N_10258);
nand U16271 (N_16271,N_14365,N_13832);
nand U16272 (N_16272,N_11646,N_10330);
or U16273 (N_16273,N_11380,N_10254);
xor U16274 (N_16274,N_12293,N_10790);
and U16275 (N_16275,N_14206,N_10539);
xnor U16276 (N_16276,N_10242,N_14918);
xnor U16277 (N_16277,N_13131,N_11772);
nor U16278 (N_16278,N_14689,N_14198);
nor U16279 (N_16279,N_10383,N_10313);
nor U16280 (N_16280,N_12331,N_11527);
nor U16281 (N_16281,N_10043,N_11414);
or U16282 (N_16282,N_10955,N_14293);
nand U16283 (N_16283,N_11848,N_13961);
or U16284 (N_16284,N_12660,N_12105);
nand U16285 (N_16285,N_12990,N_11700);
nand U16286 (N_16286,N_11673,N_12657);
nor U16287 (N_16287,N_13150,N_12957);
nand U16288 (N_16288,N_13955,N_11735);
nand U16289 (N_16289,N_13843,N_13814);
or U16290 (N_16290,N_11809,N_11317);
or U16291 (N_16291,N_11710,N_12757);
nor U16292 (N_16292,N_13767,N_11761);
nand U16293 (N_16293,N_12093,N_14262);
xnor U16294 (N_16294,N_13601,N_12371);
nor U16295 (N_16295,N_13135,N_12518);
and U16296 (N_16296,N_10702,N_11573);
nand U16297 (N_16297,N_11011,N_13765);
xnor U16298 (N_16298,N_11361,N_13120);
nand U16299 (N_16299,N_11248,N_10676);
nor U16300 (N_16300,N_13161,N_13496);
nand U16301 (N_16301,N_13616,N_13995);
xor U16302 (N_16302,N_10626,N_14417);
nand U16303 (N_16303,N_10553,N_14298);
and U16304 (N_16304,N_10735,N_11324);
xnor U16305 (N_16305,N_12999,N_12729);
and U16306 (N_16306,N_13052,N_12400);
xnor U16307 (N_16307,N_11484,N_12181);
nand U16308 (N_16308,N_11153,N_13568);
xor U16309 (N_16309,N_14113,N_13659);
xnor U16310 (N_16310,N_11869,N_11629);
nand U16311 (N_16311,N_13583,N_13605);
and U16312 (N_16312,N_11684,N_14683);
xor U16313 (N_16313,N_14143,N_11069);
or U16314 (N_16314,N_10481,N_12789);
nand U16315 (N_16315,N_13035,N_10035);
and U16316 (N_16316,N_11323,N_12420);
nand U16317 (N_16317,N_13339,N_10009);
xor U16318 (N_16318,N_13389,N_10977);
nor U16319 (N_16319,N_13155,N_14465);
nand U16320 (N_16320,N_13921,N_11294);
nor U16321 (N_16321,N_13044,N_11698);
nand U16322 (N_16322,N_10934,N_10269);
or U16323 (N_16323,N_12294,N_11546);
or U16324 (N_16324,N_13688,N_12842);
xnor U16325 (N_16325,N_11935,N_10896);
or U16326 (N_16326,N_11213,N_14557);
and U16327 (N_16327,N_11760,N_11495);
and U16328 (N_16328,N_12210,N_12582);
xnor U16329 (N_16329,N_13461,N_10340);
nand U16330 (N_16330,N_10825,N_11597);
nor U16331 (N_16331,N_14901,N_14812);
nand U16332 (N_16332,N_11611,N_14555);
and U16333 (N_16333,N_10649,N_13391);
xor U16334 (N_16334,N_12960,N_13592);
nand U16335 (N_16335,N_11274,N_14431);
or U16336 (N_16336,N_10301,N_10911);
and U16337 (N_16337,N_10164,N_10749);
nor U16338 (N_16338,N_11450,N_11437);
xnor U16339 (N_16339,N_13090,N_10618);
nor U16340 (N_16340,N_13649,N_10757);
nor U16341 (N_16341,N_12908,N_11446);
and U16342 (N_16342,N_10549,N_10409);
and U16343 (N_16343,N_14839,N_11726);
or U16344 (N_16344,N_10142,N_10093);
nor U16345 (N_16345,N_10739,N_11806);
or U16346 (N_16346,N_13098,N_13211);
or U16347 (N_16347,N_13286,N_11493);
or U16348 (N_16348,N_13613,N_11765);
or U16349 (N_16349,N_12791,N_11055);
nand U16350 (N_16350,N_12109,N_10640);
and U16351 (N_16351,N_14267,N_11750);
and U16352 (N_16352,N_12455,N_14322);
or U16353 (N_16353,N_13695,N_14751);
and U16354 (N_16354,N_13667,N_10436);
nor U16355 (N_16355,N_11047,N_13663);
xnor U16356 (N_16356,N_10918,N_13820);
and U16357 (N_16357,N_14141,N_12090);
nand U16358 (N_16358,N_14750,N_14537);
xor U16359 (N_16359,N_14317,N_10003);
or U16360 (N_16360,N_10415,N_13394);
nand U16361 (N_16361,N_11861,N_10728);
xor U16362 (N_16362,N_13432,N_14780);
and U16363 (N_16363,N_14789,N_13019);
and U16364 (N_16364,N_10813,N_14460);
nor U16365 (N_16365,N_13448,N_11045);
or U16366 (N_16366,N_12413,N_12456);
nand U16367 (N_16367,N_11871,N_12738);
xnor U16368 (N_16368,N_14581,N_10006);
nor U16369 (N_16369,N_11280,N_10534);
nor U16370 (N_16370,N_14466,N_14110);
or U16371 (N_16371,N_12778,N_10223);
xor U16372 (N_16372,N_14326,N_14735);
nor U16373 (N_16373,N_13345,N_14283);
or U16374 (N_16374,N_11357,N_14371);
nand U16375 (N_16375,N_13786,N_10961);
or U16376 (N_16376,N_14144,N_10856);
nand U16377 (N_16377,N_11395,N_10261);
xnor U16378 (N_16378,N_12103,N_14488);
or U16379 (N_16379,N_10299,N_13863);
nand U16380 (N_16380,N_14366,N_11502);
and U16381 (N_16381,N_14939,N_11560);
nor U16382 (N_16382,N_12844,N_10987);
nor U16383 (N_16383,N_14145,N_14978);
nor U16384 (N_16384,N_12772,N_12919);
xnor U16385 (N_16385,N_10981,N_12603);
nand U16386 (N_16386,N_13531,N_12690);
and U16387 (N_16387,N_10871,N_13095);
and U16388 (N_16388,N_14372,N_10969);
nand U16389 (N_16389,N_14509,N_14611);
nor U16390 (N_16390,N_13476,N_10630);
and U16391 (N_16391,N_10186,N_10448);
nor U16392 (N_16392,N_14449,N_11134);
or U16393 (N_16393,N_13431,N_12374);
and U16394 (N_16394,N_12352,N_14888);
nand U16395 (N_16395,N_13962,N_14562);
and U16396 (N_16396,N_13031,N_10116);
or U16397 (N_16397,N_12596,N_14214);
nor U16398 (N_16398,N_13972,N_10137);
nor U16399 (N_16399,N_10697,N_11862);
xnor U16400 (N_16400,N_10028,N_10510);
nor U16401 (N_16401,N_14249,N_10517);
nand U16402 (N_16402,N_11197,N_10627);
nand U16403 (N_16403,N_12556,N_14904);
or U16404 (N_16404,N_13598,N_13778);
nand U16405 (N_16405,N_14782,N_13012);
or U16406 (N_16406,N_12632,N_11211);
nor U16407 (N_16407,N_10707,N_11007);
or U16408 (N_16408,N_11690,N_11683);
and U16409 (N_16409,N_14547,N_14226);
nor U16410 (N_16410,N_10785,N_12712);
xor U16411 (N_16411,N_13087,N_12845);
xnor U16412 (N_16412,N_11699,N_13722);
nand U16413 (N_16413,N_12472,N_13067);
or U16414 (N_16414,N_12735,N_12867);
nand U16415 (N_16415,N_14430,N_10387);
xnor U16416 (N_16416,N_14473,N_13398);
nand U16417 (N_16417,N_11237,N_11999);
and U16418 (N_16418,N_11737,N_12591);
and U16419 (N_16419,N_11182,N_11982);
nand U16420 (N_16420,N_11552,N_10379);
xor U16421 (N_16421,N_10654,N_10909);
nand U16422 (N_16422,N_10367,N_14468);
xnor U16423 (N_16423,N_13173,N_13411);
nor U16424 (N_16424,N_11501,N_11663);
nand U16425 (N_16425,N_12572,N_11205);
xnor U16426 (N_16426,N_13593,N_13386);
nand U16427 (N_16427,N_14436,N_10141);
xnor U16428 (N_16428,N_13696,N_11141);
or U16429 (N_16429,N_14681,N_14743);
xor U16430 (N_16430,N_14419,N_10297);
or U16431 (N_16431,N_12727,N_14479);
and U16432 (N_16432,N_11895,N_14927);
nand U16433 (N_16433,N_11026,N_10428);
xor U16434 (N_16434,N_12722,N_12983);
xnor U16435 (N_16435,N_10349,N_14447);
nor U16436 (N_16436,N_14832,N_12978);
nor U16437 (N_16437,N_13331,N_10771);
and U16438 (N_16438,N_13689,N_11496);
xor U16439 (N_16439,N_13350,N_10811);
nor U16440 (N_16440,N_11010,N_11576);
nor U16441 (N_16441,N_12803,N_11647);
nand U16442 (N_16442,N_11705,N_13225);
or U16443 (N_16443,N_13860,N_13223);
and U16444 (N_16444,N_13276,N_14716);
nand U16445 (N_16445,N_14944,N_10828);
and U16446 (N_16446,N_13200,N_10075);
or U16447 (N_16447,N_14408,N_14835);
nand U16448 (N_16448,N_11124,N_11330);
nand U16449 (N_16449,N_12137,N_14414);
and U16450 (N_16450,N_10374,N_10010);
nor U16451 (N_16451,N_14394,N_10404);
and U16452 (N_16452,N_10485,N_11161);
xnor U16453 (N_16453,N_14496,N_10373);
xnor U16454 (N_16454,N_10248,N_14097);
or U16455 (N_16455,N_13467,N_12753);
and U16456 (N_16456,N_10590,N_13187);
nand U16457 (N_16457,N_12650,N_11081);
nor U16458 (N_16458,N_14571,N_14504);
xnor U16459 (N_16459,N_13990,N_14026);
nor U16460 (N_16460,N_13153,N_11533);
nor U16461 (N_16461,N_13473,N_11353);
nor U16462 (N_16462,N_14631,N_11731);
nor U16463 (N_16463,N_13899,N_11104);
nand U16464 (N_16464,N_14952,N_10992);
or U16465 (N_16465,N_10577,N_11458);
xor U16466 (N_16466,N_12974,N_12986);
nor U16467 (N_16467,N_12768,N_12240);
xor U16468 (N_16468,N_10842,N_11986);
and U16469 (N_16469,N_12440,N_11299);
xor U16470 (N_16470,N_10853,N_13008);
and U16471 (N_16471,N_12479,N_11499);
and U16472 (N_16472,N_10681,N_10929);
and U16473 (N_16473,N_10004,N_10268);
and U16474 (N_16474,N_14615,N_12501);
nor U16475 (N_16475,N_14288,N_10875);
nor U16476 (N_16476,N_11167,N_12698);
xor U16477 (N_16477,N_10633,N_12623);
and U16478 (N_16478,N_10275,N_14804);
and U16479 (N_16479,N_11537,N_10787);
xor U16480 (N_16480,N_13489,N_14339);
or U16481 (N_16481,N_10357,N_14850);
xnor U16482 (N_16482,N_13186,N_12513);
nor U16483 (N_16483,N_13078,N_12244);
nor U16484 (N_16484,N_11079,N_14643);
nand U16485 (N_16485,N_14021,N_12387);
and U16486 (N_16486,N_13458,N_13413);
nor U16487 (N_16487,N_13412,N_11054);
or U16488 (N_16488,N_14491,N_11391);
nand U16489 (N_16489,N_11794,N_10315);
nand U16490 (N_16490,N_14702,N_11936);
xnor U16491 (N_16491,N_12347,N_14841);
or U16492 (N_16492,N_13538,N_13447);
and U16493 (N_16493,N_13329,N_13270);
and U16494 (N_16494,N_10316,N_11544);
and U16495 (N_16495,N_10754,N_14668);
nand U16496 (N_16496,N_11687,N_13224);
nor U16497 (N_16497,N_10158,N_11120);
nand U16498 (N_16498,N_10063,N_14375);
xnor U16499 (N_16499,N_12652,N_14539);
or U16500 (N_16500,N_11171,N_10024);
xor U16501 (N_16501,N_10400,N_10733);
xor U16502 (N_16502,N_10252,N_13881);
and U16503 (N_16503,N_14010,N_14784);
xor U16504 (N_16504,N_11252,N_12874);
xor U16505 (N_16505,N_13074,N_12221);
xor U16506 (N_16506,N_10854,N_12730);
nor U16507 (N_16507,N_11388,N_14299);
or U16508 (N_16508,N_12073,N_13465);
nor U16509 (N_16509,N_13097,N_12492);
xor U16510 (N_16510,N_14830,N_12333);
or U16511 (N_16511,N_11070,N_11425);
and U16512 (N_16512,N_14648,N_10411);
nor U16513 (N_16513,N_10488,N_10447);
xnor U16514 (N_16514,N_12081,N_12211);
nand U16515 (N_16515,N_10874,N_13567);
or U16516 (N_16516,N_14846,N_10651);
nor U16517 (N_16517,N_12710,N_11967);
nor U16518 (N_16518,N_11096,N_10072);
nand U16519 (N_16519,N_11086,N_13638);
nand U16520 (N_16520,N_11114,N_10337);
nor U16521 (N_16521,N_12174,N_12852);
xor U16522 (N_16522,N_13102,N_11439);
xor U16523 (N_16523,N_12336,N_13511);
nor U16524 (N_16524,N_11358,N_11002);
or U16525 (N_16525,N_13341,N_14817);
nor U16526 (N_16526,N_13246,N_13059);
xnor U16527 (N_16527,N_10192,N_10810);
and U16528 (N_16528,N_12224,N_13774);
nand U16529 (N_16529,N_11767,N_11331);
xor U16530 (N_16530,N_12328,N_12237);
or U16531 (N_16531,N_10587,N_12692);
nor U16532 (N_16532,N_10814,N_11492);
or U16533 (N_16533,N_13579,N_14138);
xor U16534 (N_16534,N_11187,N_12002);
nand U16535 (N_16535,N_10569,N_13752);
or U16536 (N_16536,N_10263,N_10719);
nand U16537 (N_16537,N_10000,N_14207);
or U16538 (N_16538,N_14187,N_14238);
or U16539 (N_16539,N_13678,N_12559);
or U16540 (N_16540,N_12362,N_11557);
nand U16541 (N_16541,N_12820,N_11870);
and U16542 (N_16542,N_14060,N_11957);
xor U16543 (N_16543,N_13163,N_10847);
or U16544 (N_16544,N_13340,N_13446);
or U16545 (N_16545,N_11837,N_13471);
or U16546 (N_16546,N_12613,N_11983);
xor U16547 (N_16547,N_10493,N_14195);
xnor U16548 (N_16548,N_12588,N_11653);
or U16549 (N_16549,N_13220,N_14402);
nand U16550 (N_16550,N_12206,N_12928);
xor U16551 (N_16551,N_10094,N_13310);
nand U16552 (N_16552,N_11389,N_12099);
and U16553 (N_16553,N_13750,N_12932);
xnor U16554 (N_16554,N_12731,N_11587);
xor U16555 (N_16555,N_13326,N_11366);
nand U16556 (N_16556,N_12773,N_10982);
or U16557 (N_16557,N_10424,N_11101);
nor U16558 (N_16558,N_11456,N_10538);
and U16559 (N_16559,N_11614,N_12064);
xnor U16560 (N_16560,N_12041,N_12847);
nand U16561 (N_16561,N_11641,N_12416);
or U16562 (N_16562,N_10445,N_10548);
xnor U16563 (N_16563,N_13441,N_12169);
xnor U16564 (N_16564,N_12021,N_13158);
xnor U16565 (N_16565,N_14642,N_13755);
and U16566 (N_16566,N_10057,N_10171);
nor U16567 (N_16567,N_13847,N_11722);
or U16568 (N_16568,N_11747,N_13247);
nor U16569 (N_16569,N_12959,N_13128);
xnor U16570 (N_16570,N_11879,N_11932);
nor U16571 (N_16571,N_13808,N_11382);
and U16572 (N_16572,N_14820,N_11271);
xor U16573 (N_16573,N_14903,N_10959);
nor U16574 (N_16574,N_14429,N_13795);
nand U16575 (N_16575,N_11836,N_14124);
or U16576 (N_16576,N_14980,N_12056);
and U16577 (N_16577,N_11902,N_10503);
or U16578 (N_16578,N_11440,N_12683);
xnor U16579 (N_16579,N_12058,N_11746);
and U16580 (N_16580,N_12319,N_10070);
xor U16581 (N_16581,N_12868,N_12084);
nor U16582 (N_16582,N_14057,N_12494);
xor U16583 (N_16583,N_12590,N_14720);
or U16584 (N_16584,N_12356,N_13416);
or U16585 (N_16585,N_14924,N_11198);
nor U16586 (N_16586,N_13874,N_11711);
nor U16587 (N_16587,N_11790,N_14592);
and U16588 (N_16588,N_13296,N_13179);
and U16589 (N_16589,N_12193,N_10772);
or U16590 (N_16590,N_10208,N_11942);
nor U16591 (N_16591,N_11206,N_12527);
nor U16592 (N_16592,N_11118,N_10952);
and U16593 (N_16593,N_12721,N_13222);
or U16594 (N_16594,N_14270,N_10552);
and U16595 (N_16595,N_11387,N_13562);
and U16596 (N_16596,N_13043,N_12282);
or U16597 (N_16597,N_14837,N_10601);
xor U16598 (N_16598,N_13679,N_12924);
nand U16599 (N_16599,N_11259,N_11238);
nor U16600 (N_16600,N_14259,N_14713);
or U16601 (N_16601,N_11535,N_10199);
nand U16602 (N_16602,N_12836,N_13501);
nand U16603 (N_16603,N_12348,N_10629);
or U16604 (N_16604,N_14232,N_10672);
nor U16605 (N_16605,N_11992,N_11189);
and U16606 (N_16606,N_11033,N_13142);
and U16607 (N_16607,N_12839,N_11769);
nand U16608 (N_16608,N_12831,N_13757);
and U16609 (N_16609,N_13619,N_13585);
or U16610 (N_16610,N_13303,N_12815);
xor U16611 (N_16611,N_10456,N_11897);
and U16612 (N_16612,N_10342,N_14307);
nand U16613 (N_16613,N_11970,N_13789);
or U16614 (N_16614,N_14205,N_13354);
and U16615 (N_16615,N_14209,N_10429);
or U16616 (N_16616,N_10149,N_11290);
nand U16617 (N_16617,N_12577,N_14474);
nand U16618 (N_16618,N_11264,N_12482);
and U16619 (N_16619,N_12805,N_11394);
xor U16620 (N_16620,N_14697,N_13216);
nor U16621 (N_16621,N_12801,N_13053);
xnor U16622 (N_16622,N_14853,N_11835);
or U16623 (N_16623,N_12759,N_10136);
nor U16624 (N_16624,N_13970,N_10188);
xor U16625 (N_16625,N_13071,N_11333);
xor U16626 (N_16626,N_14409,N_10358);
nand U16627 (N_16627,N_12780,N_11413);
or U16628 (N_16628,N_14636,N_10113);
xor U16629 (N_16629,N_12477,N_13207);
nor U16630 (N_16630,N_13410,N_11643);
nand U16631 (N_16631,N_13824,N_11853);
nand U16632 (N_16632,N_13330,N_10151);
and U16633 (N_16633,N_12489,N_11819);
xor U16634 (N_16634,N_13085,N_12114);
or U16635 (N_16635,N_14399,N_14623);
and U16636 (N_16636,N_11032,N_13046);
or U16637 (N_16637,N_10973,N_12369);
or U16638 (N_16638,N_14958,N_11844);
xnor U16639 (N_16639,N_13402,N_10738);
nand U16640 (N_16640,N_11234,N_12851);
xnor U16641 (N_16641,N_10482,N_11628);
xor U16642 (N_16642,N_13346,N_10065);
and U16643 (N_16643,N_14891,N_11046);
and U16644 (N_16644,N_11842,N_13486);
xor U16645 (N_16645,N_12600,N_12656);
and U16646 (N_16646,N_14390,N_12217);
nand U16647 (N_16647,N_12415,N_14769);
or U16648 (N_16648,N_10030,N_14440);
nand U16649 (N_16649,N_14601,N_12933);
nor U16650 (N_16650,N_13715,N_11886);
nor U16651 (N_16651,N_11468,N_10668);
xor U16652 (N_16652,N_12259,N_14203);
xor U16653 (N_16653,N_11224,N_14777);
or U16654 (N_16654,N_13321,N_14323);
nor U16655 (N_16655,N_11670,N_10170);
nand U16656 (N_16656,N_11763,N_13264);
nand U16657 (N_16657,N_12673,N_13020);
xor U16658 (N_16658,N_13291,N_12573);
and U16659 (N_16659,N_13025,N_11910);
nand U16660 (N_16660,N_10033,N_12912);
and U16661 (N_16661,N_12394,N_14519);
nand U16662 (N_16662,N_10916,N_10054);
and U16663 (N_16663,N_10985,N_13992);
nor U16664 (N_16664,N_13148,N_12532);
nor U16665 (N_16665,N_13466,N_13414);
nor U16666 (N_16666,N_11682,N_12471);
or U16667 (N_16667,N_10886,N_12248);
xor U16668 (N_16668,N_10758,N_11365);
nor U16669 (N_16669,N_14023,N_10866);
xnor U16670 (N_16670,N_12823,N_14126);
xnor U16671 (N_16671,N_11103,N_10265);
or U16672 (N_16672,N_10562,N_11568);
xnor U16673 (N_16673,N_12005,N_14793);
xnor U16674 (N_16674,N_10666,N_10638);
and U16675 (N_16675,N_14790,N_14948);
nand U16676 (N_16676,N_13039,N_14766);
xnor U16677 (N_16677,N_10198,N_11376);
or U16678 (N_16678,N_11172,N_13351);
or U16679 (N_16679,N_10888,N_11993);
xnor U16680 (N_16680,N_12249,N_14673);
nand U16681 (N_16681,N_13604,N_12793);
or U16682 (N_16682,N_14080,N_11944);
and U16683 (N_16683,N_13042,N_14654);
nor U16684 (N_16684,N_10034,N_13574);
nand U16685 (N_16685,N_10244,N_11671);
nor U16686 (N_16686,N_14115,N_11362);
or U16687 (N_16687,N_12053,N_14725);
and U16688 (N_16688,N_13911,N_12517);
xnor U16689 (N_16689,N_14149,N_10596);
and U16690 (N_16690,N_11815,N_10472);
xnor U16691 (N_16691,N_14338,N_10062);
nand U16692 (N_16692,N_11681,N_14620);
nor U16693 (N_16693,N_11122,N_10586);
nor U16694 (N_16694,N_12292,N_13194);
nand U16695 (N_16695,N_13118,N_12327);
or U16696 (N_16696,N_10344,N_12606);
and U16697 (N_16697,N_12714,N_13878);
nand U16698 (N_16698,N_11325,N_14271);
or U16699 (N_16699,N_13009,N_12956);
and U16700 (N_16700,N_14738,N_13521);
and U16701 (N_16701,N_10692,N_12443);
or U16702 (N_16702,N_13815,N_13307);
or U16703 (N_16703,N_14915,N_11579);
or U16704 (N_16704,N_11882,N_12316);
nor U16705 (N_16705,N_14729,N_12363);
or U16706 (N_16706,N_11632,N_13364);
xnor U16707 (N_16707,N_12473,N_10277);
nand U16708 (N_16708,N_12700,N_13623);
nand U16709 (N_16709,N_12208,N_10938);
or U16710 (N_16710,N_11386,N_12144);
xor U16711 (N_16711,N_11338,N_13967);
nand U16712 (N_16712,N_14553,N_13646);
and U16713 (N_16713,N_10283,N_10410);
nand U16714 (N_16714,N_12342,N_14986);
nand U16715 (N_16715,N_13837,N_11339);
xnor U16716 (N_16716,N_12263,N_14633);
nand U16717 (N_16717,N_12424,N_10125);
xor U16718 (N_16718,N_12199,N_10195);
nor U16719 (N_16719,N_10791,N_10568);
or U16720 (N_16720,N_11445,N_12882);
or U16721 (N_16721,N_11800,N_12124);
and U16722 (N_16722,N_10716,N_13408);
nor U16723 (N_16723,N_14774,N_11504);
and U16724 (N_16724,N_11645,N_12965);
nor U16725 (N_16725,N_12326,N_10385);
and U16726 (N_16726,N_14135,N_10245);
nor U16727 (N_16727,N_10441,N_13275);
nor U16728 (N_16728,N_10597,N_10153);
nor U16729 (N_16729,N_12405,N_11780);
nand U16730 (N_16730,N_12888,N_12027);
nand U16731 (N_16731,N_13810,N_11406);
xnor U16732 (N_16732,N_12740,N_10555);
and U16733 (N_16733,N_13126,N_10849);
or U16734 (N_16734,N_12448,N_11000);
xnor U16735 (N_16735,N_11057,N_14355);
and U16736 (N_16736,N_10403,N_10475);
and U16737 (N_16737,N_13662,N_12597);
or U16738 (N_16738,N_13891,N_11351);
xor U16739 (N_16739,N_14493,N_14450);
and U16740 (N_16740,N_13706,N_14522);
and U16741 (N_16741,N_10372,N_13770);
or U16742 (N_16742,N_11066,N_14955);
and U16743 (N_16743,N_12599,N_14165);
nor U16744 (N_16744,N_10118,N_12229);
nor U16745 (N_16745,N_12280,N_12067);
nand U16746 (N_16746,N_12813,N_12040);
and U16747 (N_16747,N_10903,N_14208);
and U16748 (N_16748,N_13259,N_13561);
and U16749 (N_16749,N_14505,N_14572);
nand U16750 (N_16750,N_13084,N_10764);
and U16751 (N_16751,N_11144,N_10947);
nand U16752 (N_16752,N_13931,N_13643);
or U16753 (N_16753,N_10207,N_12994);
nand U16754 (N_16754,N_10547,N_11227);
nand U16755 (N_16755,N_12082,N_14968);
nand U16756 (N_16756,N_11555,N_12076);
and U16757 (N_16757,N_14512,N_14405);
or U16758 (N_16758,N_14815,N_10712);
nor U16759 (N_16759,N_13855,N_12670);
xor U16760 (N_16760,N_11370,N_14072);
nor U16761 (N_16761,N_13488,N_11410);
or U16762 (N_16762,N_13994,N_11667);
or U16763 (N_16763,N_10378,N_12680);
nand U16764 (N_16764,N_12857,N_10773);
or U16765 (N_16765,N_10307,N_14565);
nor U16766 (N_16766,N_13491,N_11850);
or U16767 (N_16767,N_10238,N_10620);
xor U16768 (N_16768,N_10742,N_10843);
nor U16769 (N_16769,N_11006,N_11665);
nand U16770 (N_16770,N_14301,N_13064);
or U16771 (N_16771,N_12152,N_11553);
nor U16772 (N_16772,N_11398,N_12877);
nand U16773 (N_16773,N_14223,N_11279);
or U16774 (N_16774,N_12795,N_13876);
xnor U16775 (N_16775,N_10489,N_14954);
or U16776 (N_16776,N_14983,N_13924);
and U16777 (N_16777,N_14526,N_14199);
and U16778 (N_16778,N_10175,N_10870);
or U16779 (N_16779,N_13273,N_14227);
nor U16780 (N_16780,N_13913,N_11600);
and U16781 (N_16781,N_12429,N_10610);
nand U16782 (N_16782,N_13073,N_10163);
or U16783 (N_16783,N_12651,N_13968);
xor U16784 (N_16784,N_10857,N_10259);
xor U16785 (N_16785,N_11216,N_11784);
and U16786 (N_16786,N_12555,N_12266);
and U16787 (N_16787,N_14990,N_13728);
or U16788 (N_16788,N_10477,N_11448);
nor U16789 (N_16789,N_12689,N_13905);
or U16790 (N_16790,N_12787,N_12568);
nand U16791 (N_16791,N_14551,N_11950);
nor U16792 (N_16792,N_12079,N_10235);
or U16793 (N_16793,N_13802,N_13712);
and U16794 (N_16794,N_14477,N_13072);
nor U16795 (N_16795,N_13834,N_13061);
and U16796 (N_16796,N_13633,N_14367);
nand U16797 (N_16797,N_14984,N_14439);
and U16798 (N_16798,N_11824,N_10190);
nor U16799 (N_16799,N_13134,N_14314);
nor U16800 (N_16800,N_14103,N_11887);
or U16801 (N_16801,N_11307,N_12569);
xnor U16802 (N_16802,N_13029,N_10200);
nor U16803 (N_16803,N_13980,N_12045);
and U16804 (N_16804,N_14734,N_11127);
nor U16805 (N_16805,N_11115,N_14230);
xor U16806 (N_16806,N_13209,N_14092);
xnor U16807 (N_16807,N_11846,N_11638);
nand U16808 (N_16808,N_13368,N_14772);
nand U16809 (N_16809,N_12189,N_12642);
nor U16810 (N_16810,N_13237,N_14497);
nor U16811 (N_16811,N_13485,N_11044);
nor U16812 (N_16812,N_11058,N_10913);
or U16813 (N_16813,N_12687,N_14998);
nand U16814 (N_16814,N_11979,N_12004);
and U16815 (N_16815,N_14706,N_14320);
and U16816 (N_16816,N_12520,N_10206);
nor U16817 (N_16817,N_11655,N_10855);
xnor U16818 (N_16818,N_12403,N_12645);
nand U16819 (N_16819,N_11580,N_13859);
nand U16820 (N_16820,N_12157,N_10390);
nor U16821 (N_16821,N_13729,N_10423);
or U16822 (N_16822,N_14160,N_12907);
xnor U16823 (N_16823,N_11666,N_10022);
and U16824 (N_16824,N_10786,N_13252);
and U16825 (N_16825,N_10406,N_14960);
and U16826 (N_16826,N_14217,N_14674);
nor U16827 (N_16827,N_14887,N_11781);
nand U16828 (N_16828,N_14971,N_10296);
xor U16829 (N_16829,N_14996,N_11898);
and U16830 (N_16830,N_14310,N_13858);
nor U16831 (N_16831,N_14525,N_11610);
nand U16832 (N_16832,N_12175,N_11566);
or U16833 (N_16833,N_14905,N_13070);
and U16834 (N_16834,N_10468,N_10076);
xnor U16835 (N_16835,N_13487,N_11265);
and U16836 (N_16836,N_14235,N_11529);
nand U16837 (N_16837,N_10750,N_13596);
or U16838 (N_16838,N_14018,N_11454);
and U16839 (N_16839,N_13856,N_11946);
or U16840 (N_16840,N_10822,N_12454);
or U16841 (N_16841,N_11179,N_12046);
nor U16842 (N_16842,N_11960,N_12872);
and U16843 (N_16843,N_10370,N_14597);
and U16844 (N_16844,N_13817,N_14956);
or U16845 (N_16845,N_14411,N_13263);
or U16846 (N_16846,N_12036,N_10278);
nand U16847 (N_16847,N_13758,N_11570);
xnor U16848 (N_16848,N_13262,N_12281);
xor U16849 (N_16849,N_11938,N_11603);
or U16850 (N_16850,N_10452,N_10550);
nor U16851 (N_16851,N_13724,N_10709);
or U16852 (N_16852,N_12467,N_13280);
and U16853 (N_16853,N_11411,N_10829);
and U16854 (N_16854,N_10127,N_14988);
nor U16855 (N_16855,N_12688,N_10935);
and U16856 (N_16856,N_12711,N_10622);
nand U16857 (N_16857,N_13497,N_13577);
or U16858 (N_16858,N_10220,N_11190);
and U16859 (N_16859,N_14578,N_12159);
nor U16860 (N_16860,N_12381,N_13602);
xor U16861 (N_16861,N_11830,N_11247);
xor U16862 (N_16862,N_10839,N_10939);
or U16863 (N_16863,N_13529,N_11212);
nor U16864 (N_16864,N_13407,N_13954);
and U16865 (N_16865,N_10049,N_13336);
xnor U16866 (N_16866,N_11880,N_13683);
nor U16867 (N_16867,N_12207,N_11039);
nand U16868 (N_16868,N_12062,N_13845);
or U16869 (N_16869,N_10529,N_10401);
nand U16870 (N_16870,N_11475,N_11480);
nor U16871 (N_16871,N_14062,N_14433);
and U16872 (N_16872,N_10045,N_12349);
nand U16873 (N_16873,N_10945,N_10189);
nor U16874 (N_16874,N_14626,N_12507);
nor U16875 (N_16875,N_10196,N_10942);
and U16876 (N_16876,N_14071,N_14407);
or U16877 (N_16877,N_11316,N_11686);
or U16878 (N_16878,N_11071,N_11169);
nand U16879 (N_16879,N_13640,N_13555);
nor U16880 (N_16880,N_12496,N_14121);
nor U16881 (N_16881,N_10891,N_10435);
xor U16882 (N_16882,N_12119,N_12802);
nand U16883 (N_16883,N_11154,N_14156);
or U16884 (N_16884,N_13685,N_13241);
nor U16885 (N_16885,N_11884,N_10455);
and U16886 (N_16886,N_11548,N_12843);
or U16887 (N_16887,N_12140,N_11194);
nor U16888 (N_16888,N_10368,N_12035);
and U16889 (N_16889,N_12895,N_13014);
xnor U16890 (N_16890,N_10407,N_10588);
and U16891 (N_16891,N_10774,N_10704);
and U16892 (N_16892,N_13760,N_14239);
xor U16893 (N_16893,N_14132,N_14325);
nand U16894 (N_16894,N_11753,N_11578);
nand U16895 (N_16895,N_14985,N_13953);
nor U16896 (N_16896,N_14552,N_11640);
or U16897 (N_16897,N_12038,N_14506);
and U16898 (N_16898,N_13764,N_14289);
or U16899 (N_16899,N_11605,N_14576);
xor U16900 (N_16900,N_10713,N_11613);
nand U16901 (N_16901,N_14704,N_12557);
xnor U16902 (N_16902,N_12807,N_12950);
xor U16903 (N_16903,N_11969,N_11137);
nand U16904 (N_16904,N_10607,N_10218);
nand U16905 (N_16905,N_12421,N_12811);
xnor U16906 (N_16906,N_12121,N_14911);
or U16907 (N_16907,N_11245,N_13797);
nor U16908 (N_16908,N_13614,N_12257);
nand U16909 (N_16909,N_11777,N_14929);
and U16910 (N_16910,N_11063,N_14081);
nor U16911 (N_16911,N_14511,N_13987);
or U16912 (N_16912,N_13691,N_11964);
or U16913 (N_16913,N_14004,N_12899);
nand U16914 (N_16914,N_10497,N_12905);
nand U16915 (N_16915,N_13556,N_11758);
or U16916 (N_16916,N_14127,N_12345);
and U16917 (N_16917,N_14027,N_10879);
xnor U16918 (N_16918,N_12893,N_12922);
nor U16919 (N_16919,N_11409,N_12133);
or U16920 (N_16920,N_13552,N_11188);
nor U16921 (N_16921,N_14515,N_14033);
xnor U16922 (N_16922,N_13482,N_14638);
and U16923 (N_16923,N_10970,N_11485);
xor U16924 (N_16924,N_14802,N_11892);
or U16925 (N_16925,N_10908,N_14554);
or U16926 (N_16926,N_12579,N_14666);
or U16927 (N_16927,N_13217,N_10120);
and U16928 (N_16928,N_11959,N_14917);
or U16929 (N_16929,N_13671,N_10334);
or U16930 (N_16930,N_13873,N_13791);
nor U16931 (N_16931,N_11867,N_12153);
nor U16932 (N_16932,N_12338,N_12265);
xor U16933 (N_16933,N_14694,N_14029);
xor U16934 (N_16934,N_10782,N_13589);
nand U16935 (N_16935,N_10303,N_13904);
nand U16936 (N_16936,N_13888,N_11486);
and U16937 (N_16937,N_13504,N_14932);
or U16938 (N_16938,N_12864,N_14574);
or U16939 (N_16939,N_11511,N_13595);
or U16940 (N_16940,N_10637,N_11296);
xnor U16941 (N_16941,N_14286,N_13769);
nand U16942 (N_16942,N_12026,N_14377);
xor U16943 (N_16943,N_13582,N_14329);
or U16944 (N_16944,N_12612,N_14434);
or U16945 (N_16945,N_13900,N_12399);
nor U16946 (N_16946,N_11634,N_11025);
or U16947 (N_16947,N_12853,N_14152);
or U16948 (N_16948,N_13444,N_13702);
or U16949 (N_16949,N_10581,N_11701);
or U16950 (N_16950,N_11604,N_14699);
xor U16951 (N_16951,N_12011,N_12750);
and U16952 (N_16952,N_10172,N_13588);
nor U16953 (N_16953,N_14012,N_14398);
and U16954 (N_16954,N_10958,N_13522);
and U16955 (N_16955,N_13966,N_12565);
nand U16956 (N_16956,N_13244,N_14695);
nand U16957 (N_16957,N_12177,N_10256);
or U16958 (N_16958,N_14728,N_13338);
nand U16959 (N_16959,N_10007,N_12914);
or U16960 (N_16960,N_11005,N_13711);
nor U16961 (N_16961,N_12550,N_12846);
nand U16962 (N_16962,N_10167,N_14125);
nand U16963 (N_16963,N_14520,N_14821);
and U16964 (N_16964,N_14700,N_11736);
and U16965 (N_16965,N_10815,N_11651);
or U16966 (N_16966,N_10397,N_11547);
or U16967 (N_16967,N_11277,N_13734);
nand U16968 (N_16968,N_10262,N_11575);
and U16969 (N_16969,N_13550,N_11549);
or U16970 (N_16970,N_12776,N_12484);
or U16971 (N_16971,N_12693,N_12783);
or U16972 (N_16972,N_10536,N_10234);
or U16973 (N_16973,N_13532,N_12502);
xnor U16974 (N_16974,N_12892,N_14893);
nand U16975 (N_16975,N_10635,N_11872);
nor U16976 (N_16976,N_11685,N_11829);
or U16977 (N_16977,N_10479,N_13773);
or U16978 (N_16978,N_10393,N_13081);
and U16979 (N_16979,N_10809,N_12982);
xor U16980 (N_16980,N_14950,N_11543);
and U16981 (N_16981,N_10213,N_11734);
and U16982 (N_16982,N_14906,N_11210);
and U16983 (N_16983,N_14827,N_11244);
or U16984 (N_16984,N_11251,N_10795);
or U16985 (N_16985,N_10384,N_10470);
or U16986 (N_16986,N_11567,N_12139);
nor U16987 (N_16987,N_12107,N_10121);
nand U16988 (N_16988,N_12833,N_11065);
xor U16989 (N_16989,N_12699,N_11148);
xor U16990 (N_16990,N_13609,N_12806);
and U16991 (N_16991,N_11619,N_12931);
and U16992 (N_16992,N_14864,N_14912);
nor U16993 (N_16993,N_12320,N_13289);
xor U16994 (N_16994,N_12499,N_14873);
xor U16995 (N_16995,N_14454,N_11968);
and U16996 (N_16996,N_13320,N_12165);
and U16997 (N_16997,N_13494,N_11742);
xnor U16998 (N_16998,N_10976,N_11542);
nand U16999 (N_16999,N_13294,N_11181);
or U17000 (N_17000,N_14711,N_10971);
nand U17001 (N_17001,N_10684,N_12332);
nand U17002 (N_17002,N_12643,N_10161);
or U17003 (N_17003,N_12271,N_14186);
nor U17004 (N_17004,N_12411,N_10726);
or U17005 (N_17005,N_12775,N_14210);
xor U17006 (N_17006,N_13692,N_12526);
nor U17007 (N_17007,N_13928,N_12587);
and U17008 (N_17008,N_12634,N_12697);
xnor U17009 (N_17009,N_11721,N_12270);
and U17010 (N_17010,N_12135,N_13230);
nand U17011 (N_17011,N_11367,N_11003);
nor U17012 (N_17012,N_12302,N_10943);
or U17013 (N_17013,N_10351,N_14809);
nand U17014 (N_17014,N_14247,N_11152);
nand U17015 (N_17015,N_11432,N_12359);
nor U17016 (N_17016,N_12115,N_13437);
and U17017 (N_17017,N_11180,N_14922);
xnor U17018 (N_17018,N_11202,N_12008);
nand U17019 (N_17019,N_14761,N_13618);
and U17020 (N_17020,N_14649,N_10718);
nor U17021 (N_17021,N_11350,N_14382);
or U17022 (N_17022,N_13634,N_10176);
or U17023 (N_17023,N_11788,N_13065);
nor U17024 (N_17024,N_14880,N_12792);
or U17025 (N_17025,N_14882,N_11522);
and U17026 (N_17026,N_10181,N_10695);
xor U17027 (N_17027,N_14055,N_12401);
nand U17028 (N_17028,N_14589,N_13935);
or U17029 (N_17029,N_10890,N_14052);
xor U17030 (N_17030,N_12039,N_12376);
or U17031 (N_17031,N_13798,N_12164);
xor U17032 (N_17032,N_14723,N_14381);
and U17033 (N_17033,N_13912,N_14868);
and U17034 (N_17034,N_11680,N_13104);
xor U17035 (N_17035,N_11948,N_11393);
or U17036 (N_17036,N_11193,N_14560);
nor U17037 (N_17037,N_14427,N_10271);
nor U17038 (N_17038,N_13066,N_11825);
xor U17039 (N_17039,N_11466,N_13030);
nor U17040 (N_17040,N_12298,N_13022);
xor U17041 (N_17041,N_10535,N_13871);
xor U17042 (N_17042,N_12903,N_12493);
nand U17043 (N_17043,N_13189,N_12878);
xor U17044 (N_17044,N_10760,N_12560);
and U17045 (N_17045,N_14085,N_14413);
nand U17046 (N_17046,N_13430,N_10418);
xor U17047 (N_17047,N_12988,N_12295);
nor U17048 (N_17048,N_10940,N_12463);
and U17049 (N_17049,N_14616,N_14471);
nor U17050 (N_17050,N_10933,N_10308);
and U17051 (N_17051,N_11412,N_10979);
or U17052 (N_17052,N_13342,N_14773);
and U17053 (N_17053,N_14895,N_11094);
xor U17054 (N_17054,N_11822,N_12508);
nand U17055 (N_17055,N_12800,N_12745);
nor U17056 (N_17056,N_13929,N_11478);
nand U17057 (N_17057,N_10467,N_10721);
nor U17058 (N_17058,N_11349,N_14162);
and U17059 (N_17059,N_11243,N_11268);
xor U17060 (N_17060,N_11396,N_12425);
nand U17061 (N_17061,N_11973,N_11909);
or U17062 (N_17062,N_11839,N_11506);
nand U17063 (N_17063,N_13356,N_12621);
or U17064 (N_17064,N_10312,N_10841);
or U17065 (N_17065,N_11952,N_11658);
xor U17066 (N_17066,N_10852,N_13149);
nor U17067 (N_17067,N_12188,N_12719);
nand U17068 (N_17068,N_12072,N_13775);
or U17069 (N_17069,N_12629,N_10114);
or U17070 (N_17070,N_14770,N_14945);
xor U17071 (N_17071,N_13736,N_12024);
or U17072 (N_17072,N_14351,N_12160);
nand U17073 (N_17073,N_14415,N_12996);
nor U17074 (N_17074,N_10266,N_13677);
or U17075 (N_17075,N_13107,N_14093);
and U17076 (N_17076,N_11832,N_13690);
nand U17077 (N_17077,N_11196,N_14759);
and U17078 (N_17078,N_10737,N_11427);
xor U17079 (N_17079,N_11219,N_13578);
and U17080 (N_17080,N_12426,N_13218);
nand U17081 (N_17081,N_11452,N_13344);
or U17082 (N_17082,N_10820,N_12993);
nor U17083 (N_17083,N_12663,N_13392);
and U17084 (N_17084,N_11048,N_13720);
xnor U17085 (N_17085,N_14369,N_11487);
nor U17086 (N_17086,N_11659,N_13387);
nand U17087 (N_17087,N_13054,N_10123);
or U17088 (N_17088,N_10129,N_11467);
and U17089 (N_17089,N_12215,N_10154);
and U17090 (N_17090,N_11796,N_11004);
nand U17091 (N_17091,N_14368,N_10542);
xnor U17092 (N_17092,N_12325,N_10696);
or U17093 (N_17093,N_13943,N_10026);
or U17094 (N_17094,N_11803,N_13088);
nand U17095 (N_17095,N_13828,N_12197);
and U17096 (N_17096,N_13991,N_11038);
nand U17097 (N_17097,N_14024,N_11230);
or U17098 (N_17098,N_11847,N_12214);
and U17099 (N_17099,N_14614,N_10052);
or U17100 (N_17100,N_13175,N_11095);
xnor U17101 (N_17101,N_10144,N_12464);
nand U17102 (N_17102,N_13352,N_13199);
or U17103 (N_17103,N_11013,N_13886);
and U17104 (N_17104,N_13076,N_14861);
and U17105 (N_17105,N_12127,N_13591);
xor U17106 (N_17106,N_11209,N_12183);
and U17107 (N_17107,N_11129,N_11704);
or U17108 (N_17108,N_14190,N_13288);
nand U17109 (N_17109,N_14418,N_10498);
and U17110 (N_17110,N_12373,N_12274);
nand U17111 (N_17111,N_13205,N_10862);
nor U17112 (N_17112,N_10703,N_10160);
or U17113 (N_17113,N_12367,N_14114);
xnor U17114 (N_17114,N_11689,N_11132);
and U17115 (N_17115,N_12771,N_10147);
xnor U17116 (N_17116,N_10838,N_14885);
nor U17117 (N_17117,N_11927,N_10960);
or U17118 (N_17118,N_13919,N_10079);
and U17119 (N_17119,N_11336,N_14896);
nor U17120 (N_17120,N_12913,N_14538);
xor U17121 (N_17121,N_13918,N_14105);
and U17122 (N_17122,N_13013,N_13367);
nor U17123 (N_17123,N_14925,N_13141);
nor U17124 (N_17124,N_13940,N_10500);
nand U17125 (N_17125,N_10591,N_11811);
nand U17126 (N_17126,N_10991,N_11329);
nand U17127 (N_17127,N_11098,N_10567);
and U17128 (N_17128,N_10107,N_14075);
and U17129 (N_17129,N_10907,N_12478);
or U17130 (N_17130,N_12476,N_10157);
nor U17131 (N_17131,N_10558,N_10767);
or U17132 (N_17132,N_12968,N_10274);
and U17133 (N_17133,N_13306,N_14255);
nand U17134 (N_17134,N_14336,N_11664);
and U17135 (N_17135,N_13212,N_13399);
or U17136 (N_17136,N_13839,N_11717);
xor U17137 (N_17137,N_12243,N_10522);
and U17138 (N_17138,N_14624,N_13506);
nand U17139 (N_17139,N_13427,N_14951);
nand U17140 (N_17140,N_11131,N_11472);
xor U17141 (N_17141,N_13809,N_10818);
xor U17142 (N_17142,N_10867,N_13514);
xnor U17143 (N_17143,N_12528,N_13324);
and U17144 (N_17144,N_11116,N_14705);
and U17145 (N_17145,N_12794,N_10197);
xor U17146 (N_17146,N_12460,N_11151);
xor U17147 (N_17147,N_13232,N_11672);
xor U17148 (N_17148,N_10675,N_11420);
xnor U17149 (N_17149,N_11097,N_10796);
nor U17150 (N_17150,N_13287,N_13751);
nor U17151 (N_17151,N_13541,N_13136);
nand U17152 (N_17152,N_11166,N_13785);
nor U17153 (N_17153,N_11177,N_13631);
xnor U17154 (N_17154,N_11108,N_12398);
nand U17155 (N_17155,N_14421,N_14865);
nand U17156 (N_17156,N_13297,N_12375);
nand U17157 (N_17157,N_12495,N_12774);
nand U17158 (N_17158,N_10537,N_14120);
xor U17159 (N_17159,N_14346,N_13569);
and U17160 (N_17160,N_13549,N_10047);
or U17161 (N_17161,N_12544,N_14744);
or U17162 (N_17162,N_13500,N_14510);
nor U17163 (N_17163,N_14353,N_14296);
xor U17164 (N_17164,N_14653,N_14602);
nand U17165 (N_17165,N_12018,N_13006);
nand U17166 (N_17166,N_12451,N_14096);
xnor U17167 (N_17167,N_10002,N_11998);
nand U17168 (N_17168,N_14902,N_11416);
nor U17169 (N_17169,N_10817,N_13805);
xor U17170 (N_17170,N_10768,N_10449);
nand U17171 (N_17171,N_13608,N_13816);
xnor U17172 (N_17172,N_10012,N_11564);
or U17173 (N_17173,N_10214,N_10381);
or U17174 (N_17174,N_11297,N_14569);
or U17175 (N_17175,N_12042,N_12324);
nand U17176 (N_17176,N_14051,N_14231);
xnor U17177 (N_17177,N_14726,N_14910);
and U17178 (N_17178,N_10496,N_11799);
xnor U17179 (N_17179,N_13939,N_10925);
xnor U17180 (N_17180,N_10480,N_11273);
xor U17181 (N_17181,N_13417,N_13388);
xor U17182 (N_17182,N_10615,N_10717);
xor U17183 (N_17183,N_12861,N_13196);
or U17184 (N_17184,N_11239,N_13754);
nand U17185 (N_17185,N_14194,N_11314);
xor U17186 (N_17186,N_10306,N_10458);
nand U17187 (N_17187,N_10059,N_12821);
and U17188 (N_17188,N_13783,N_12826);
nand U17189 (N_17189,N_14957,N_13060);
and U17190 (N_17190,N_11519,N_11525);
and U17191 (N_17191,N_11217,N_10068);
xnor U17192 (N_17192,N_12125,N_14358);
and U17193 (N_17193,N_11465,N_10402);
or U17194 (N_17194,N_10715,N_14617);
and U17195 (N_17195,N_14308,N_13254);
nand U17196 (N_17196,N_10285,N_12365);
nor U17197 (N_17197,N_12589,N_14786);
xnor U17198 (N_17198,N_13732,N_14671);
nand U17199 (N_17199,N_13877,N_10784);
or U17200 (N_17200,N_13537,N_10356);
xnor U17201 (N_17201,N_12945,N_12031);
nand U17202 (N_17202,N_14116,N_14972);
xnor U17203 (N_17203,N_11621,N_13460);
xor U17204 (N_17204,N_11258,N_14946);
nand U17205 (N_17205,N_11577,N_11162);
xnor U17206 (N_17206,N_12659,N_12417);
or U17207 (N_17207,N_10042,N_14536);
and U17208 (N_17208,N_14923,N_13472);
and U17209 (N_17209,N_11369,N_13033);
or U17210 (N_17210,N_14395,N_10014);
and U17211 (N_17211,N_10844,N_11322);
xor U17212 (N_17212,N_13265,N_14279);
xnor U17213 (N_17213,N_13978,N_13741);
nor U17214 (N_17214,N_11951,N_11514);
and U17215 (N_17215,N_11232,N_14588);
or U17216 (N_17216,N_13879,N_11076);
xor U17217 (N_17217,N_11520,N_11282);
xnor U17218 (N_17218,N_14599,N_13812);
nor U17219 (N_17219,N_14645,N_14964);
nor U17220 (N_17220,N_14678,N_13080);
nor U17221 (N_17221,N_12916,N_12809);
nor U17222 (N_17222,N_10352,N_12594);
or U17223 (N_17223,N_12571,N_11572);
and U17224 (N_17224,N_11818,N_11315);
nand U17225 (N_17225,N_11028,N_13779);
xor U17226 (N_17226,N_13788,N_13564);
nand U17227 (N_17227,N_11195,N_13675);
xnor U17228 (N_17228,N_11751,N_13001);
and U17229 (N_17229,N_11782,N_13348);
nand U17230 (N_17230,N_13308,N_12117);
nor U17231 (N_17231,N_14048,N_14712);
nand U17232 (N_17232,N_12973,N_14717);
nand U17233 (N_17233,N_10328,N_12523);
and U17234 (N_17234,N_10636,N_13358);
xnor U17235 (N_17235,N_12200,N_14690);
xnor U17236 (N_17236,N_11849,N_11616);
nor U17237 (N_17237,N_14142,N_14401);
and U17238 (N_17238,N_10652,N_13145);
and U17239 (N_17239,N_14831,N_13133);
nor U17240 (N_17240,N_11589,N_13168);
nand U17241 (N_17241,N_14197,N_14265);
xor U17242 (N_17242,N_13673,N_13293);
nand U17243 (N_17243,N_12264,N_10798);
and U17244 (N_17244,N_13234,N_12481);
or U17245 (N_17245,N_11415,N_12396);
nand U17246 (N_17246,N_10882,N_14073);
and U17247 (N_17247,N_12122,N_14117);
nand U17248 (N_17248,N_13772,N_12209);
or U17249 (N_17249,N_11405,N_10989);
and U17250 (N_17250,N_14284,N_12445);
nor U17251 (N_17251,N_14393,N_12102);
nor U17252 (N_17252,N_13811,N_14215);
or U17253 (N_17253,N_11697,N_12595);
xnor U17254 (N_17254,N_11994,N_11513);
xnor U17255 (N_17255,N_10290,N_12970);
and U17256 (N_17256,N_12695,N_10515);
or U17257 (N_17257,N_10126,N_13651);
nor U17258 (N_17258,N_10746,N_11656);
or U17259 (N_17259,N_11304,N_12303);
nor U17260 (N_17260,N_12227,N_12551);
xor U17261 (N_17261,N_12498,N_10102);
nand U17262 (N_17262,N_10359,N_12881);
and U17263 (N_17263,N_10264,N_11907);
nand U17264 (N_17264,N_13611,N_14282);
nand U17265 (N_17265,N_13822,N_12790);
xor U17266 (N_17266,N_11598,N_13018);
nor U17267 (N_17267,N_13401,N_10228);
or U17268 (N_17268,N_12733,N_10806);
xnor U17269 (N_17269,N_14783,N_10878);
or U17270 (N_17270,N_12925,N_13985);
xnor U17271 (N_17271,N_12641,N_14147);
and U17272 (N_17272,N_13969,N_13701);
nor U17273 (N_17273,N_10104,N_12969);
or U17274 (N_17274,N_13661,N_10067);
nor U17275 (N_17275,N_10744,N_11802);
nor U17276 (N_17276,N_10819,N_10162);
nand U17277 (N_17277,N_10044,N_12458);
xnor U17278 (N_17278,N_12686,N_12929);
xnor U17279 (N_17279,N_12339,N_13584);
or U17280 (N_17280,N_13442,N_10803);
and U17281 (N_17281,N_10354,N_14570);
and U17282 (N_17282,N_14131,N_11727);
nor U17283 (N_17283,N_13378,N_13279);
xor U17284 (N_17284,N_12025,N_13396);
nor U17285 (N_17285,N_11087,N_12942);
nand U17286 (N_17286,N_11287,N_10090);
and U17287 (N_17287,N_13171,N_11310);
xnor U17288 (N_17288,N_12315,N_11925);
nor U17289 (N_17289,N_14796,N_14914);
xor U17290 (N_17290,N_11929,N_14070);
or U17291 (N_17291,N_11817,N_14740);
xor U17292 (N_17292,N_10763,N_10348);
xnor U17293 (N_17293,N_14280,N_13083);
or U17294 (N_17294,N_12457,N_11798);
and U17295 (N_17295,N_14201,N_13093);
nand U17296 (N_17296,N_12601,N_14933);
xnor U17297 (N_17297,N_11536,N_10095);
or U17298 (N_17298,N_14622,N_10150);
or U17299 (N_17299,N_12447,N_10794);
xnor U17300 (N_17300,N_12863,N_13127);
nor U17301 (N_17301,N_12285,N_12296);
and U17302 (N_17302,N_12086,N_13933);
and U17303 (N_17303,N_13470,N_12812);
xor U17304 (N_17304,N_14775,N_14243);
nor U17305 (N_17305,N_13781,N_11741);
nor U17306 (N_17306,N_10683,N_11523);
nand U17307 (N_17307,N_14318,N_11713);
and U17308 (N_17308,N_10469,N_13454);
nor U17309 (N_17309,N_10293,N_11534);
xnor U17310 (N_17310,N_12887,N_12536);
nand U17311 (N_17311,N_13091,N_10382);
nand U17312 (N_17312,N_10605,N_11136);
nand U17313 (N_17313,N_13188,N_13193);
nor U17314 (N_17314,N_10281,N_11157);
and U17315 (N_17315,N_13684,N_12896);
nor U17316 (N_17316,N_14605,N_13079);
xnor U17317 (N_17317,N_13763,N_13385);
nand U17318 (N_17318,N_11914,N_10682);
nor U17319 (N_17319,N_13909,N_13674);
and U17320 (N_17320,N_13896,N_14331);
nand U17321 (N_17321,N_12483,N_11379);
or U17322 (N_17322,N_12014,N_12098);
nand U17323 (N_17323,N_10288,N_13157);
xor U17324 (N_17324,N_11293,N_12267);
or U17325 (N_17325,N_13144,N_10331);
or U17326 (N_17326,N_12563,N_13748);
or U17327 (N_17327,N_12717,N_13101);
nand U17328 (N_17328,N_12713,N_10350);
and U17329 (N_17329,N_11752,N_14083);
nor U17330 (N_17330,N_12674,N_12584);
nand U17331 (N_17331,N_10965,N_10872);
nor U17332 (N_17332,N_13258,N_13190);
or U17333 (N_17333,N_13323,N_10658);
or U17334 (N_17334,N_14340,N_12049);
nand U17335 (N_17335,N_12128,N_10322);
nor U17336 (N_17336,N_12196,N_10901);
and U17337 (N_17337,N_13122,N_12954);
xnor U17338 (N_17338,N_10051,N_12788);
xnor U17339 (N_17339,N_13892,N_12192);
nor U17340 (N_17340,N_14993,N_10159);
nor U17341 (N_17341,N_11309,N_14254);
nor U17342 (N_17342,N_11278,N_11302);
and U17343 (N_17343,N_13236,N_13152);
or U17344 (N_17344,N_14328,N_10069);
nand U17345 (N_17345,N_12377,N_13761);
or U17346 (N_17346,N_10604,N_12385);
or U17347 (N_17347,N_11214,N_12233);
or U17348 (N_17348,N_14884,N_11677);
xnor U17349 (N_17349,N_12522,N_10177);
and U17350 (N_17350,N_11260,N_11200);
nand U17351 (N_17351,N_10426,N_13214);
nor U17352 (N_17352,N_10680,N_12981);
nand U17353 (N_17353,N_13818,N_11408);
or U17354 (N_17354,N_12620,N_14102);
nand U17355 (N_17355,N_12009,N_11064);
and U17356 (N_17356,N_11510,N_14872);
nor U17357 (N_17357,N_11785,N_13620);
and U17358 (N_17358,N_11061,N_13707);
nor U17359 (N_17359,N_11657,N_14490);
or U17360 (N_17360,N_10417,N_11400);
nor U17361 (N_17361,N_13178,N_11319);
xor U17362 (N_17362,N_13890,N_14028);
and U17363 (N_17363,N_10731,N_12230);
nor U17364 (N_17364,N_12901,N_10863);
and U17365 (N_17365,N_10302,N_13794);
and U17366 (N_17366,N_13182,N_14107);
nor U17367 (N_17367,N_14161,N_12311);
nor U17368 (N_17368,N_10936,N_13159);
and U17369 (N_17369,N_10521,N_11771);
nor U17370 (N_17370,N_11917,N_13151);
nand U17371 (N_17371,N_13445,N_14056);
and U17372 (N_17372,N_14148,N_13617);
nor U17373 (N_17373,N_13226,N_10623);
nand U17374 (N_17374,N_12684,N_11249);
or U17375 (N_17375,N_10694,N_12987);
and U17376 (N_17376,N_13570,N_10645);
nand U17377 (N_17377,N_11250,N_13986);
and U17378 (N_17378,N_14309,N_14973);
nor U17379 (N_17379,N_10686,N_12962);
nand U17380 (N_17380,N_14909,N_13010);
and U17381 (N_17381,N_11939,N_11106);
nor U17382 (N_17382,N_10135,N_11636);
xor U17383 (N_17383,N_12647,N_10914);
nand U17384 (N_17384,N_12392,N_12158);
or U17385 (N_17385,N_10667,N_14164);
or U17386 (N_17386,N_10326,N_10336);
nand U17387 (N_17387,N_14258,N_13125);
xnor U17388 (N_17388,N_11779,N_10017);
xnor U17389 (N_17389,N_10812,N_10184);
nand U17390 (N_17390,N_14007,N_13694);
nor U17391 (N_17391,N_14794,N_11723);
nor U17392 (N_17392,N_12608,N_14503);
nand U17393 (N_17393,N_11036,N_10644);
or U17394 (N_17394,N_14727,N_14123);
nand U17395 (N_17395,N_13302,N_13826);
and U17396 (N_17396,N_13456,N_13908);
xor U17397 (N_17397,N_12578,N_11894);
nor U17398 (N_17398,N_13123,N_11143);
nand U17399 (N_17399,N_11584,N_11235);
nand U17400 (N_17400,N_13718,N_12198);
and U17401 (N_17401,N_10061,N_14797);
nor U17402 (N_17402,N_13973,N_10725);
xnor U17403 (N_17403,N_11285,N_12012);
xor U17404 (N_17404,N_12936,N_12841);
nand U17405 (N_17405,N_12190,N_12354);
and U17406 (N_17406,N_14452,N_13325);
or U17407 (N_17407,N_14947,N_10765);
and U17408 (N_17408,N_10673,N_10698);
nor U17409 (N_17409,N_13405,N_14890);
nor U17410 (N_17410,N_14416,N_13930);
xor U17411 (N_17411,N_11360,N_11266);
nand U17412 (N_17412,N_13875,N_13314);
nand U17413 (N_17413,N_13332,N_12763);
and U17414 (N_17414,N_14253,N_12754);
nand U17415 (N_17415,N_12497,N_11989);
xor U17416 (N_17416,N_13932,N_10227);
xor U17417 (N_17417,N_10311,N_11178);
nand U17418 (N_17418,N_14003,N_10700);
and U17419 (N_17419,N_13024,N_12355);
nand U17420 (N_17420,N_10755,N_11858);
xor U17421 (N_17421,N_11128,N_10608);
nand U17422 (N_17422,N_14763,N_11976);
nand U17423 (N_17423,N_10140,N_13599);
or U17424 (N_17424,N_12116,N_12891);
and U17425 (N_17425,N_14272,N_12180);
xor U17426 (N_17426,N_13597,N_10305);
xor U17427 (N_17427,N_10711,N_14753);
nand U17428 (N_17428,N_11593,N_14961);
xor U17429 (N_17429,N_14682,N_12808);
xor U17430 (N_17430,N_12245,N_13547);
nand U17431 (N_17431,N_12361,N_10462);
or U17432 (N_17432,N_14524,N_10956);
nand U17433 (N_17433,N_10433,N_10097);
nor U17434 (N_17434,N_12223,N_12583);
xnor U17435 (N_17435,N_14894,N_13525);
xnor U17436 (N_17436,N_11748,N_10085);
or U17437 (N_17437,N_13069,N_12186);
xnor U17438 (N_17438,N_12716,N_10656);
or U17439 (N_17439,N_11708,N_12386);
and U17440 (N_17440,N_10883,N_12239);
or U17441 (N_17441,N_12834,N_13092);
nor U17442 (N_17442,N_10609,N_14291);
xor U17443 (N_17443,N_13464,N_12779);
or U17444 (N_17444,N_12030,N_14069);
nor U17445 (N_17445,N_13533,N_11770);
nand U17446 (N_17446,N_13668,N_12370);
nor U17447 (N_17447,N_12340,N_12762);
nor U17448 (N_17448,N_10353,N_12254);
nand U17449 (N_17449,N_12894,N_10201);
nor U17450 (N_17450,N_14795,N_13766);
and U17451 (N_17451,N_10221,N_10650);
xnor U17452 (N_17452,N_12106,N_12055);
nor U17453 (N_17453,N_10325,N_14758);
or U17454 (N_17454,N_11223,N_14297);
and U17455 (N_17455,N_11691,N_12781);
nand U17456 (N_17456,N_14019,N_11716);
xor U17457 (N_17457,N_12911,N_11754);
nand U17458 (N_17458,N_14844,N_12567);
xor U17459 (N_17459,N_10371,N_11569);
nor U17460 (N_17460,N_13139,N_14136);
nor U17461 (N_17461,N_13451,N_11675);
nand U17462 (N_17462,N_10117,N_14420);
xnor U17463 (N_17463,N_13806,N_13068);
xor U17464 (N_17464,N_13819,N_12148);
nor U17465 (N_17465,N_10594,N_14229);
and U17466 (N_17466,N_12061,N_14808);
nor U17467 (N_17467,N_13922,N_14014);
nand U17468 (N_17468,N_10446,N_12586);
or U17469 (N_17469,N_10386,N_13195);
nor U17470 (N_17470,N_10483,N_10018);
xnor U17471 (N_17471,N_14724,N_14661);
xor U17472 (N_17472,N_10168,N_10364);
xor U17473 (N_17473,N_13138,N_14785);
nand U17474 (N_17474,N_13827,N_10425);
nand U17475 (N_17475,N_14962,N_14805);
nor U17476 (N_17476,N_10884,N_12366);
and U17477 (N_17477,N_11630,N_14495);
xnor U17478 (N_17478,N_12450,N_13041);
nand U17479 (N_17479,N_14222,N_11461);
nor U17480 (N_17480,N_13744,N_11341);
xnor U17481 (N_17481,N_11257,N_10408);
nand U17482 (N_17482,N_14163,N_14498);
nand U17483 (N_17483,N_11138,N_13530);
and U17484 (N_17484,N_14866,N_14316);
nor U17485 (N_17485,N_11429,N_14315);
nor U17486 (N_17486,N_11313,N_11311);
nor U17487 (N_17487,N_13669,N_13343);
nor U17488 (N_17488,N_13698,N_11444);
and U17489 (N_17489,N_11014,N_10714);
nor U17490 (N_17490,N_13656,N_14938);
nand U17491 (N_17491,N_11423,N_13956);
nand U17492 (N_17492,N_12001,N_11253);
xnor U17493 (N_17493,N_13535,N_12437);
nor U17494 (N_17494,N_10823,N_13203);
or U17495 (N_17495,N_11900,N_11130);
xor U17496 (N_17496,N_12992,N_13016);
xor U17497 (N_17497,N_10084,N_10071);
or U17498 (N_17498,N_13594,N_14949);
nand U17499 (N_17499,N_11435,N_14154);
nor U17500 (N_17500,N_14036,N_11149);
or U17501 (N_17501,N_10270,N_14728);
xor U17502 (N_17502,N_10336,N_14086);
xor U17503 (N_17503,N_10923,N_11294);
or U17504 (N_17504,N_10198,N_13213);
or U17505 (N_17505,N_14712,N_14644);
and U17506 (N_17506,N_12000,N_12019);
xor U17507 (N_17507,N_12335,N_13482);
nand U17508 (N_17508,N_14054,N_13739);
xnor U17509 (N_17509,N_12115,N_14544);
nor U17510 (N_17510,N_12244,N_14170);
and U17511 (N_17511,N_13074,N_13036);
and U17512 (N_17512,N_14920,N_13528);
nor U17513 (N_17513,N_14006,N_13026);
nor U17514 (N_17514,N_10015,N_13467);
xor U17515 (N_17515,N_13212,N_12625);
nor U17516 (N_17516,N_12248,N_13740);
and U17517 (N_17517,N_10992,N_13757);
nand U17518 (N_17518,N_11381,N_13496);
or U17519 (N_17519,N_14505,N_11985);
nand U17520 (N_17520,N_13972,N_10737);
or U17521 (N_17521,N_12292,N_10342);
and U17522 (N_17522,N_14839,N_10659);
and U17523 (N_17523,N_10739,N_13128);
nor U17524 (N_17524,N_12053,N_12217);
or U17525 (N_17525,N_10716,N_14777);
xnor U17526 (N_17526,N_12419,N_12069);
and U17527 (N_17527,N_14100,N_13274);
nand U17528 (N_17528,N_13638,N_10200);
nand U17529 (N_17529,N_10138,N_12364);
or U17530 (N_17530,N_14181,N_12196);
or U17531 (N_17531,N_10929,N_11716);
or U17532 (N_17532,N_10825,N_11694);
or U17533 (N_17533,N_14777,N_10481);
xnor U17534 (N_17534,N_14017,N_13885);
nand U17535 (N_17535,N_14501,N_12488);
nor U17536 (N_17536,N_13840,N_12603);
xor U17537 (N_17537,N_11348,N_12567);
or U17538 (N_17538,N_13056,N_10143);
xor U17539 (N_17539,N_12747,N_11036);
xor U17540 (N_17540,N_11259,N_14895);
and U17541 (N_17541,N_13608,N_10315);
nand U17542 (N_17542,N_10094,N_11368);
nand U17543 (N_17543,N_13343,N_10543);
or U17544 (N_17544,N_12183,N_13963);
or U17545 (N_17545,N_13340,N_13014);
xnor U17546 (N_17546,N_13713,N_13513);
xor U17547 (N_17547,N_14736,N_12754);
and U17548 (N_17548,N_13788,N_14507);
nand U17549 (N_17549,N_10679,N_13549);
or U17550 (N_17550,N_11446,N_13224);
and U17551 (N_17551,N_10023,N_14961);
and U17552 (N_17552,N_11692,N_12622);
or U17553 (N_17553,N_11270,N_11376);
or U17554 (N_17554,N_11983,N_11897);
xnor U17555 (N_17555,N_14120,N_13281);
nand U17556 (N_17556,N_10383,N_10944);
and U17557 (N_17557,N_12133,N_13576);
or U17558 (N_17558,N_10933,N_13522);
xnor U17559 (N_17559,N_14028,N_12058);
and U17560 (N_17560,N_13400,N_10073);
and U17561 (N_17561,N_11316,N_11579);
nor U17562 (N_17562,N_11873,N_10020);
nand U17563 (N_17563,N_14839,N_13316);
nand U17564 (N_17564,N_12846,N_12286);
and U17565 (N_17565,N_13313,N_14388);
nand U17566 (N_17566,N_13928,N_13590);
nor U17567 (N_17567,N_12439,N_12852);
nand U17568 (N_17568,N_14420,N_11019);
nor U17569 (N_17569,N_13006,N_12843);
and U17570 (N_17570,N_10424,N_13713);
and U17571 (N_17571,N_10680,N_13081);
or U17572 (N_17572,N_14846,N_11975);
nand U17573 (N_17573,N_12504,N_14432);
nor U17574 (N_17574,N_10681,N_11980);
xor U17575 (N_17575,N_11305,N_10411);
and U17576 (N_17576,N_11955,N_13119);
and U17577 (N_17577,N_12409,N_10801);
xnor U17578 (N_17578,N_12322,N_11843);
and U17579 (N_17579,N_10898,N_14575);
and U17580 (N_17580,N_11499,N_10891);
xor U17581 (N_17581,N_13866,N_13056);
or U17582 (N_17582,N_12965,N_11008);
xnor U17583 (N_17583,N_10361,N_14129);
or U17584 (N_17584,N_12630,N_13132);
nand U17585 (N_17585,N_11929,N_13340);
nor U17586 (N_17586,N_13421,N_13172);
nand U17587 (N_17587,N_12209,N_10232);
nor U17588 (N_17588,N_14256,N_14021);
nand U17589 (N_17589,N_12576,N_10877);
or U17590 (N_17590,N_13903,N_13265);
nor U17591 (N_17591,N_13751,N_10643);
nand U17592 (N_17592,N_13227,N_10036);
or U17593 (N_17593,N_11006,N_13620);
nand U17594 (N_17594,N_11561,N_13633);
and U17595 (N_17595,N_14785,N_12362);
and U17596 (N_17596,N_14045,N_12490);
nand U17597 (N_17597,N_10470,N_14258);
or U17598 (N_17598,N_11766,N_13514);
and U17599 (N_17599,N_11450,N_10833);
xnor U17600 (N_17600,N_14925,N_10335);
nand U17601 (N_17601,N_13629,N_14044);
and U17602 (N_17602,N_11802,N_12278);
xor U17603 (N_17603,N_12236,N_10235);
nand U17604 (N_17604,N_10913,N_14730);
nand U17605 (N_17605,N_13555,N_11076);
or U17606 (N_17606,N_14482,N_12842);
or U17607 (N_17607,N_12462,N_13987);
and U17608 (N_17608,N_12042,N_12571);
xor U17609 (N_17609,N_10368,N_13101);
or U17610 (N_17610,N_12511,N_13800);
nor U17611 (N_17611,N_10797,N_11823);
or U17612 (N_17612,N_13486,N_14588);
xnor U17613 (N_17613,N_14301,N_14028);
nand U17614 (N_17614,N_14685,N_13764);
nor U17615 (N_17615,N_14540,N_14451);
or U17616 (N_17616,N_14076,N_12335);
and U17617 (N_17617,N_12291,N_14827);
xnor U17618 (N_17618,N_10159,N_10042);
or U17619 (N_17619,N_13880,N_12106);
nand U17620 (N_17620,N_13087,N_10945);
nor U17621 (N_17621,N_14374,N_11711);
or U17622 (N_17622,N_14362,N_13916);
nand U17623 (N_17623,N_12624,N_13683);
xnor U17624 (N_17624,N_11370,N_10400);
nand U17625 (N_17625,N_13249,N_13671);
and U17626 (N_17626,N_14313,N_11732);
and U17627 (N_17627,N_14823,N_10317);
and U17628 (N_17628,N_11451,N_10285);
or U17629 (N_17629,N_13033,N_13952);
or U17630 (N_17630,N_13170,N_11543);
or U17631 (N_17631,N_11276,N_13511);
and U17632 (N_17632,N_11926,N_12913);
nor U17633 (N_17633,N_12784,N_10596);
and U17634 (N_17634,N_10304,N_11714);
xnor U17635 (N_17635,N_13106,N_13323);
and U17636 (N_17636,N_13399,N_12443);
nor U17637 (N_17637,N_13063,N_12743);
or U17638 (N_17638,N_14819,N_10599);
nor U17639 (N_17639,N_10028,N_12560);
nand U17640 (N_17640,N_11426,N_11193);
or U17641 (N_17641,N_13171,N_12171);
or U17642 (N_17642,N_11388,N_10402);
and U17643 (N_17643,N_14257,N_10684);
nand U17644 (N_17644,N_10994,N_12065);
xnor U17645 (N_17645,N_10716,N_12749);
or U17646 (N_17646,N_11719,N_10985);
nand U17647 (N_17647,N_10415,N_13133);
nor U17648 (N_17648,N_12631,N_10621);
xnor U17649 (N_17649,N_13090,N_14933);
or U17650 (N_17650,N_13755,N_12580);
and U17651 (N_17651,N_11106,N_13526);
xnor U17652 (N_17652,N_10555,N_12373);
or U17653 (N_17653,N_10111,N_14599);
nor U17654 (N_17654,N_13157,N_12151);
or U17655 (N_17655,N_13664,N_14845);
xor U17656 (N_17656,N_14292,N_14220);
or U17657 (N_17657,N_12640,N_10324);
nor U17658 (N_17658,N_11825,N_14412);
nand U17659 (N_17659,N_13784,N_11609);
and U17660 (N_17660,N_14002,N_13649);
or U17661 (N_17661,N_12729,N_13289);
nor U17662 (N_17662,N_11765,N_14496);
xor U17663 (N_17663,N_12975,N_13080);
nand U17664 (N_17664,N_12961,N_10646);
nor U17665 (N_17665,N_11426,N_13529);
nor U17666 (N_17666,N_10042,N_11265);
nand U17667 (N_17667,N_10238,N_11718);
xnor U17668 (N_17668,N_14478,N_13754);
xnor U17669 (N_17669,N_14873,N_13932);
xor U17670 (N_17670,N_12822,N_13131);
nor U17671 (N_17671,N_12980,N_11940);
or U17672 (N_17672,N_14975,N_14862);
nand U17673 (N_17673,N_12834,N_13236);
and U17674 (N_17674,N_12722,N_11356);
or U17675 (N_17675,N_13412,N_13869);
and U17676 (N_17676,N_12937,N_14615);
nand U17677 (N_17677,N_14611,N_11499);
xor U17678 (N_17678,N_12338,N_14488);
xor U17679 (N_17679,N_14822,N_14032);
and U17680 (N_17680,N_10757,N_11394);
and U17681 (N_17681,N_14387,N_14165);
and U17682 (N_17682,N_14726,N_14851);
xnor U17683 (N_17683,N_14835,N_11313);
nor U17684 (N_17684,N_14067,N_11439);
and U17685 (N_17685,N_13776,N_13686);
xnor U17686 (N_17686,N_12653,N_11461);
xor U17687 (N_17687,N_13508,N_14233);
nor U17688 (N_17688,N_13646,N_11006);
xnor U17689 (N_17689,N_11960,N_14308);
xor U17690 (N_17690,N_12255,N_10487);
xnor U17691 (N_17691,N_13040,N_11599);
or U17692 (N_17692,N_11507,N_13071);
and U17693 (N_17693,N_12393,N_10751);
nand U17694 (N_17694,N_10098,N_12261);
or U17695 (N_17695,N_14936,N_13978);
or U17696 (N_17696,N_10205,N_12043);
or U17697 (N_17697,N_13873,N_14206);
nor U17698 (N_17698,N_13676,N_12715);
or U17699 (N_17699,N_10026,N_13076);
and U17700 (N_17700,N_11701,N_11798);
nor U17701 (N_17701,N_12017,N_10171);
nand U17702 (N_17702,N_12610,N_10487);
nand U17703 (N_17703,N_10086,N_10443);
nand U17704 (N_17704,N_10999,N_11875);
and U17705 (N_17705,N_12203,N_11410);
nor U17706 (N_17706,N_10488,N_12827);
xnor U17707 (N_17707,N_10616,N_13469);
nand U17708 (N_17708,N_14119,N_10319);
nor U17709 (N_17709,N_11322,N_10305);
or U17710 (N_17710,N_14550,N_14003);
nand U17711 (N_17711,N_11452,N_11774);
xor U17712 (N_17712,N_13203,N_12736);
nand U17713 (N_17713,N_13803,N_10466);
nor U17714 (N_17714,N_11501,N_13989);
nand U17715 (N_17715,N_14632,N_11634);
and U17716 (N_17716,N_11142,N_10770);
nor U17717 (N_17717,N_12857,N_11067);
and U17718 (N_17718,N_14658,N_11203);
or U17719 (N_17719,N_13932,N_14829);
nand U17720 (N_17720,N_12465,N_14517);
or U17721 (N_17721,N_14545,N_13382);
or U17722 (N_17722,N_14589,N_11745);
nor U17723 (N_17723,N_12295,N_13586);
and U17724 (N_17724,N_11764,N_13259);
or U17725 (N_17725,N_13753,N_11241);
and U17726 (N_17726,N_13556,N_13537);
nand U17727 (N_17727,N_10962,N_12096);
or U17728 (N_17728,N_14663,N_13091);
or U17729 (N_17729,N_10073,N_14019);
and U17730 (N_17730,N_12232,N_13504);
xor U17731 (N_17731,N_13681,N_11645);
nand U17732 (N_17732,N_13697,N_11347);
or U17733 (N_17733,N_14170,N_11451);
nand U17734 (N_17734,N_14365,N_13768);
or U17735 (N_17735,N_12538,N_10866);
and U17736 (N_17736,N_10063,N_11027);
nand U17737 (N_17737,N_10895,N_14244);
nand U17738 (N_17738,N_14781,N_14851);
xnor U17739 (N_17739,N_14382,N_13860);
nor U17740 (N_17740,N_12091,N_14294);
xor U17741 (N_17741,N_11436,N_14826);
xor U17742 (N_17742,N_13144,N_11232);
xor U17743 (N_17743,N_14045,N_14263);
and U17744 (N_17744,N_12102,N_11717);
or U17745 (N_17745,N_10110,N_14566);
or U17746 (N_17746,N_13577,N_13117);
nor U17747 (N_17747,N_11624,N_13334);
xnor U17748 (N_17748,N_13169,N_12769);
xor U17749 (N_17749,N_10834,N_14852);
nor U17750 (N_17750,N_14000,N_14183);
nand U17751 (N_17751,N_14370,N_11867);
and U17752 (N_17752,N_13116,N_10275);
or U17753 (N_17753,N_10691,N_13695);
nor U17754 (N_17754,N_14054,N_14831);
nand U17755 (N_17755,N_10929,N_13140);
nor U17756 (N_17756,N_14356,N_14504);
nor U17757 (N_17757,N_10210,N_10717);
or U17758 (N_17758,N_14294,N_11184);
xnor U17759 (N_17759,N_11705,N_12839);
and U17760 (N_17760,N_13104,N_10354);
xnor U17761 (N_17761,N_10822,N_14804);
or U17762 (N_17762,N_11817,N_11831);
nor U17763 (N_17763,N_14593,N_10955);
nand U17764 (N_17764,N_10113,N_13651);
nand U17765 (N_17765,N_12891,N_13505);
and U17766 (N_17766,N_11906,N_10980);
and U17767 (N_17767,N_10345,N_12845);
or U17768 (N_17768,N_11351,N_10578);
xor U17769 (N_17769,N_12773,N_14313);
xnor U17770 (N_17770,N_11256,N_10099);
and U17771 (N_17771,N_12799,N_10451);
nand U17772 (N_17772,N_11060,N_11054);
and U17773 (N_17773,N_11909,N_13607);
or U17774 (N_17774,N_13197,N_12019);
xnor U17775 (N_17775,N_14961,N_13481);
xnor U17776 (N_17776,N_11818,N_10090);
nand U17777 (N_17777,N_10731,N_14297);
nor U17778 (N_17778,N_13831,N_10818);
nand U17779 (N_17779,N_12983,N_11397);
or U17780 (N_17780,N_13087,N_12388);
nor U17781 (N_17781,N_14138,N_14962);
nor U17782 (N_17782,N_12690,N_13747);
nor U17783 (N_17783,N_13876,N_11909);
xor U17784 (N_17784,N_11955,N_10072);
or U17785 (N_17785,N_13799,N_14731);
nand U17786 (N_17786,N_10429,N_13045);
nor U17787 (N_17787,N_10992,N_10786);
nor U17788 (N_17788,N_11256,N_12006);
and U17789 (N_17789,N_11129,N_10891);
and U17790 (N_17790,N_10166,N_10498);
xnor U17791 (N_17791,N_14703,N_11597);
nand U17792 (N_17792,N_11771,N_13755);
or U17793 (N_17793,N_12571,N_14137);
nor U17794 (N_17794,N_10766,N_13789);
nand U17795 (N_17795,N_10079,N_14234);
or U17796 (N_17796,N_13219,N_11174);
nor U17797 (N_17797,N_12157,N_14284);
or U17798 (N_17798,N_14487,N_14376);
nor U17799 (N_17799,N_14710,N_10059);
or U17800 (N_17800,N_14837,N_10132);
xnor U17801 (N_17801,N_11147,N_14957);
and U17802 (N_17802,N_13522,N_11162);
nand U17803 (N_17803,N_10966,N_12963);
xnor U17804 (N_17804,N_14989,N_14736);
or U17805 (N_17805,N_11832,N_12043);
nor U17806 (N_17806,N_14345,N_11847);
or U17807 (N_17807,N_14795,N_14741);
xor U17808 (N_17808,N_11671,N_13280);
nor U17809 (N_17809,N_13983,N_10648);
and U17810 (N_17810,N_11229,N_10015);
and U17811 (N_17811,N_12150,N_14858);
nor U17812 (N_17812,N_14084,N_10351);
xor U17813 (N_17813,N_10703,N_11397);
xor U17814 (N_17814,N_14633,N_12936);
xnor U17815 (N_17815,N_10239,N_13162);
xor U17816 (N_17816,N_11507,N_13505);
and U17817 (N_17817,N_14537,N_14012);
nor U17818 (N_17818,N_11674,N_11331);
nor U17819 (N_17819,N_10069,N_14812);
nand U17820 (N_17820,N_14755,N_11824);
and U17821 (N_17821,N_12205,N_10677);
and U17822 (N_17822,N_14748,N_14940);
nor U17823 (N_17823,N_10237,N_11519);
nand U17824 (N_17824,N_13071,N_10655);
xnor U17825 (N_17825,N_10076,N_14438);
nand U17826 (N_17826,N_14190,N_11210);
and U17827 (N_17827,N_13931,N_13889);
nand U17828 (N_17828,N_10464,N_14543);
or U17829 (N_17829,N_14221,N_10482);
xnor U17830 (N_17830,N_13405,N_10055);
nand U17831 (N_17831,N_10053,N_14975);
and U17832 (N_17832,N_10654,N_13657);
and U17833 (N_17833,N_11933,N_12211);
or U17834 (N_17834,N_14888,N_13381);
xor U17835 (N_17835,N_10660,N_13020);
or U17836 (N_17836,N_13110,N_13236);
or U17837 (N_17837,N_12487,N_12346);
and U17838 (N_17838,N_12005,N_12211);
or U17839 (N_17839,N_10483,N_12797);
nand U17840 (N_17840,N_12639,N_11272);
nand U17841 (N_17841,N_11484,N_11676);
nand U17842 (N_17842,N_12669,N_13025);
xnor U17843 (N_17843,N_10648,N_12775);
and U17844 (N_17844,N_10998,N_11458);
or U17845 (N_17845,N_10522,N_10848);
or U17846 (N_17846,N_11514,N_11221);
and U17847 (N_17847,N_13201,N_12347);
nand U17848 (N_17848,N_11154,N_14975);
nor U17849 (N_17849,N_10344,N_13636);
xor U17850 (N_17850,N_12359,N_14089);
and U17851 (N_17851,N_12654,N_11527);
nor U17852 (N_17852,N_14009,N_10402);
nor U17853 (N_17853,N_10954,N_11914);
nand U17854 (N_17854,N_13266,N_13409);
xor U17855 (N_17855,N_10605,N_11945);
or U17856 (N_17856,N_11567,N_11246);
or U17857 (N_17857,N_12680,N_14662);
nand U17858 (N_17858,N_14620,N_14014);
xor U17859 (N_17859,N_11182,N_13441);
or U17860 (N_17860,N_13887,N_13978);
and U17861 (N_17861,N_12565,N_11294);
xor U17862 (N_17862,N_10745,N_13572);
nand U17863 (N_17863,N_13171,N_13719);
and U17864 (N_17864,N_10154,N_12006);
and U17865 (N_17865,N_12416,N_11442);
xnor U17866 (N_17866,N_13958,N_10742);
nand U17867 (N_17867,N_13151,N_10844);
nand U17868 (N_17868,N_14791,N_11472);
nand U17869 (N_17869,N_12146,N_10103);
or U17870 (N_17870,N_13833,N_11657);
or U17871 (N_17871,N_13867,N_13438);
nor U17872 (N_17872,N_13953,N_10765);
and U17873 (N_17873,N_14719,N_13302);
and U17874 (N_17874,N_11092,N_13086);
xor U17875 (N_17875,N_11447,N_10879);
nor U17876 (N_17876,N_12233,N_13826);
nor U17877 (N_17877,N_14536,N_14270);
nor U17878 (N_17878,N_13588,N_12459);
nand U17879 (N_17879,N_13349,N_13276);
or U17880 (N_17880,N_12992,N_10194);
and U17881 (N_17881,N_14771,N_13556);
nand U17882 (N_17882,N_13539,N_12322);
nand U17883 (N_17883,N_12719,N_10444);
or U17884 (N_17884,N_14959,N_12593);
nand U17885 (N_17885,N_10778,N_13298);
nor U17886 (N_17886,N_13637,N_14703);
xor U17887 (N_17887,N_14187,N_12246);
or U17888 (N_17888,N_14320,N_13863);
nor U17889 (N_17889,N_14979,N_13451);
or U17890 (N_17890,N_14959,N_13653);
nor U17891 (N_17891,N_12497,N_13492);
nor U17892 (N_17892,N_12990,N_12607);
nand U17893 (N_17893,N_13698,N_11241);
and U17894 (N_17894,N_13287,N_13961);
or U17895 (N_17895,N_14719,N_11921);
nand U17896 (N_17896,N_11470,N_12598);
or U17897 (N_17897,N_10006,N_13031);
and U17898 (N_17898,N_12347,N_10185);
xor U17899 (N_17899,N_13657,N_11930);
nand U17900 (N_17900,N_12429,N_13850);
nand U17901 (N_17901,N_11448,N_12653);
xor U17902 (N_17902,N_12586,N_14230);
and U17903 (N_17903,N_11926,N_14899);
or U17904 (N_17904,N_12124,N_12985);
xnor U17905 (N_17905,N_14917,N_14334);
nor U17906 (N_17906,N_13259,N_10077);
nand U17907 (N_17907,N_13944,N_13676);
xor U17908 (N_17908,N_11019,N_10331);
and U17909 (N_17909,N_13762,N_14256);
xnor U17910 (N_17910,N_11146,N_12440);
xor U17911 (N_17911,N_14272,N_12926);
xor U17912 (N_17912,N_12173,N_14449);
xnor U17913 (N_17913,N_11621,N_12681);
nor U17914 (N_17914,N_12780,N_12228);
nor U17915 (N_17915,N_10889,N_13402);
nand U17916 (N_17916,N_10852,N_11297);
nor U17917 (N_17917,N_13605,N_12996);
or U17918 (N_17918,N_14266,N_14273);
nand U17919 (N_17919,N_10627,N_11876);
and U17920 (N_17920,N_13710,N_11867);
nand U17921 (N_17921,N_14604,N_12896);
or U17922 (N_17922,N_14682,N_12831);
nand U17923 (N_17923,N_13487,N_12274);
xnor U17924 (N_17924,N_14124,N_14195);
nand U17925 (N_17925,N_14789,N_10414);
and U17926 (N_17926,N_11666,N_13815);
nor U17927 (N_17927,N_13858,N_14565);
or U17928 (N_17928,N_14412,N_12530);
or U17929 (N_17929,N_14806,N_13992);
nor U17930 (N_17930,N_14003,N_13102);
and U17931 (N_17931,N_13063,N_14157);
nand U17932 (N_17932,N_13073,N_14823);
nor U17933 (N_17933,N_11614,N_11605);
nor U17934 (N_17934,N_11577,N_12336);
and U17935 (N_17935,N_10701,N_11014);
or U17936 (N_17936,N_14516,N_13513);
or U17937 (N_17937,N_12728,N_12011);
nand U17938 (N_17938,N_12685,N_11952);
xor U17939 (N_17939,N_13997,N_11753);
nor U17940 (N_17940,N_11823,N_14307);
nand U17941 (N_17941,N_13043,N_11344);
nor U17942 (N_17942,N_14845,N_12073);
and U17943 (N_17943,N_12932,N_14696);
and U17944 (N_17944,N_12203,N_14350);
or U17945 (N_17945,N_11388,N_13193);
or U17946 (N_17946,N_12951,N_10094);
or U17947 (N_17947,N_11569,N_12862);
and U17948 (N_17948,N_12668,N_11567);
nor U17949 (N_17949,N_11189,N_13334);
nand U17950 (N_17950,N_12048,N_14494);
nand U17951 (N_17951,N_12659,N_12354);
nor U17952 (N_17952,N_13261,N_11437);
and U17953 (N_17953,N_13938,N_12327);
xnor U17954 (N_17954,N_12500,N_12039);
or U17955 (N_17955,N_12357,N_10808);
or U17956 (N_17956,N_14934,N_11195);
or U17957 (N_17957,N_13615,N_10096);
or U17958 (N_17958,N_12709,N_10014);
nand U17959 (N_17959,N_11966,N_13391);
and U17960 (N_17960,N_14784,N_11774);
nand U17961 (N_17961,N_10782,N_12416);
xor U17962 (N_17962,N_14774,N_12895);
nor U17963 (N_17963,N_14329,N_14814);
nor U17964 (N_17964,N_12400,N_12080);
nor U17965 (N_17965,N_14685,N_12150);
or U17966 (N_17966,N_13834,N_11199);
nor U17967 (N_17967,N_14873,N_11532);
nand U17968 (N_17968,N_10004,N_13997);
or U17969 (N_17969,N_13976,N_11577);
or U17970 (N_17970,N_11963,N_11251);
and U17971 (N_17971,N_13261,N_14932);
xnor U17972 (N_17972,N_13209,N_11367);
xor U17973 (N_17973,N_12336,N_13299);
and U17974 (N_17974,N_13907,N_12342);
and U17975 (N_17975,N_12295,N_13867);
or U17976 (N_17976,N_11295,N_12952);
and U17977 (N_17977,N_11490,N_11028);
and U17978 (N_17978,N_13453,N_14133);
nand U17979 (N_17979,N_11053,N_10058);
or U17980 (N_17980,N_14225,N_14665);
nand U17981 (N_17981,N_10158,N_12601);
or U17982 (N_17982,N_13036,N_10208);
or U17983 (N_17983,N_11351,N_14777);
xor U17984 (N_17984,N_12542,N_11107);
nand U17985 (N_17985,N_11857,N_14858);
and U17986 (N_17986,N_13165,N_10584);
nand U17987 (N_17987,N_14194,N_14814);
nor U17988 (N_17988,N_12772,N_11468);
nor U17989 (N_17989,N_11101,N_12786);
and U17990 (N_17990,N_12148,N_12346);
or U17991 (N_17991,N_12407,N_12372);
nor U17992 (N_17992,N_14336,N_11596);
nor U17993 (N_17993,N_11619,N_14925);
nand U17994 (N_17994,N_13003,N_14738);
nand U17995 (N_17995,N_11059,N_13355);
or U17996 (N_17996,N_11173,N_13923);
xnor U17997 (N_17997,N_13017,N_13614);
nand U17998 (N_17998,N_13424,N_12463);
nand U17999 (N_17999,N_11203,N_13064);
nor U18000 (N_18000,N_14420,N_14418);
nor U18001 (N_18001,N_10009,N_10537);
xnor U18002 (N_18002,N_11874,N_13324);
nor U18003 (N_18003,N_13856,N_10028);
nand U18004 (N_18004,N_12520,N_10372);
nand U18005 (N_18005,N_10118,N_12878);
or U18006 (N_18006,N_11003,N_10466);
nor U18007 (N_18007,N_14204,N_10565);
xnor U18008 (N_18008,N_13805,N_10610);
and U18009 (N_18009,N_11530,N_14576);
nand U18010 (N_18010,N_10880,N_13345);
nor U18011 (N_18011,N_12507,N_12271);
nor U18012 (N_18012,N_12907,N_10619);
or U18013 (N_18013,N_11337,N_12997);
or U18014 (N_18014,N_14633,N_10964);
nand U18015 (N_18015,N_14759,N_13802);
or U18016 (N_18016,N_10438,N_11034);
or U18017 (N_18017,N_12494,N_14139);
xnor U18018 (N_18018,N_12474,N_12154);
nand U18019 (N_18019,N_14448,N_12589);
nor U18020 (N_18020,N_14685,N_12517);
and U18021 (N_18021,N_10631,N_11990);
or U18022 (N_18022,N_13115,N_12287);
nand U18023 (N_18023,N_11519,N_11319);
nor U18024 (N_18024,N_13797,N_14653);
nor U18025 (N_18025,N_13098,N_11346);
xnor U18026 (N_18026,N_12523,N_10924);
and U18027 (N_18027,N_14825,N_12728);
xnor U18028 (N_18028,N_14584,N_13340);
and U18029 (N_18029,N_13958,N_10265);
nor U18030 (N_18030,N_12014,N_14352);
or U18031 (N_18031,N_13002,N_10228);
xnor U18032 (N_18032,N_14725,N_14295);
and U18033 (N_18033,N_14951,N_12368);
nand U18034 (N_18034,N_10000,N_13809);
and U18035 (N_18035,N_14903,N_14336);
xor U18036 (N_18036,N_12308,N_11723);
xor U18037 (N_18037,N_12503,N_10585);
or U18038 (N_18038,N_10803,N_13284);
nor U18039 (N_18039,N_10952,N_11292);
nand U18040 (N_18040,N_14568,N_12446);
nand U18041 (N_18041,N_14177,N_10698);
and U18042 (N_18042,N_10855,N_11646);
and U18043 (N_18043,N_11325,N_11067);
nor U18044 (N_18044,N_10912,N_12445);
or U18045 (N_18045,N_10375,N_11734);
nor U18046 (N_18046,N_14518,N_11767);
xnor U18047 (N_18047,N_11132,N_13978);
and U18048 (N_18048,N_13656,N_14496);
and U18049 (N_18049,N_10156,N_14831);
xor U18050 (N_18050,N_13195,N_13900);
and U18051 (N_18051,N_14658,N_10163);
xor U18052 (N_18052,N_11281,N_13694);
or U18053 (N_18053,N_10538,N_10099);
nand U18054 (N_18054,N_13474,N_12312);
nand U18055 (N_18055,N_10828,N_11468);
or U18056 (N_18056,N_14983,N_13698);
nor U18057 (N_18057,N_13605,N_14899);
nand U18058 (N_18058,N_10249,N_12469);
nand U18059 (N_18059,N_10907,N_11229);
xnor U18060 (N_18060,N_13061,N_10643);
or U18061 (N_18061,N_12220,N_11258);
xor U18062 (N_18062,N_12176,N_11689);
nor U18063 (N_18063,N_13634,N_13839);
nand U18064 (N_18064,N_12743,N_10911);
or U18065 (N_18065,N_14858,N_11636);
xnor U18066 (N_18066,N_13913,N_11880);
nor U18067 (N_18067,N_12648,N_10948);
nor U18068 (N_18068,N_10390,N_10139);
xnor U18069 (N_18069,N_11476,N_10628);
nor U18070 (N_18070,N_11715,N_12674);
nor U18071 (N_18071,N_11519,N_10795);
nor U18072 (N_18072,N_11133,N_10919);
xor U18073 (N_18073,N_11139,N_13207);
xnor U18074 (N_18074,N_14453,N_14301);
nor U18075 (N_18075,N_14619,N_12380);
nand U18076 (N_18076,N_12115,N_10532);
nor U18077 (N_18077,N_14707,N_12106);
or U18078 (N_18078,N_13207,N_13224);
or U18079 (N_18079,N_14190,N_14261);
nand U18080 (N_18080,N_10390,N_12594);
nand U18081 (N_18081,N_12966,N_14207);
nor U18082 (N_18082,N_10135,N_11890);
nor U18083 (N_18083,N_10732,N_14384);
nor U18084 (N_18084,N_12507,N_11950);
nor U18085 (N_18085,N_12128,N_12514);
or U18086 (N_18086,N_12048,N_10466);
and U18087 (N_18087,N_13088,N_10679);
xor U18088 (N_18088,N_13980,N_14585);
nand U18089 (N_18089,N_14149,N_11271);
xor U18090 (N_18090,N_13600,N_10903);
and U18091 (N_18091,N_12472,N_13763);
nor U18092 (N_18092,N_11434,N_13668);
or U18093 (N_18093,N_13558,N_10609);
xnor U18094 (N_18094,N_10882,N_12748);
and U18095 (N_18095,N_14616,N_13064);
xnor U18096 (N_18096,N_11349,N_11579);
nor U18097 (N_18097,N_10317,N_13254);
nand U18098 (N_18098,N_10213,N_13551);
or U18099 (N_18099,N_12769,N_13355);
nand U18100 (N_18100,N_10876,N_12530);
xor U18101 (N_18101,N_12421,N_13338);
xnor U18102 (N_18102,N_11840,N_12684);
and U18103 (N_18103,N_11605,N_13325);
and U18104 (N_18104,N_10957,N_11064);
xor U18105 (N_18105,N_12566,N_14369);
nand U18106 (N_18106,N_12759,N_11904);
and U18107 (N_18107,N_10751,N_10418);
and U18108 (N_18108,N_13857,N_14068);
or U18109 (N_18109,N_12611,N_10308);
xor U18110 (N_18110,N_14270,N_12510);
nor U18111 (N_18111,N_12873,N_10838);
xor U18112 (N_18112,N_13930,N_13669);
or U18113 (N_18113,N_11005,N_13917);
xor U18114 (N_18114,N_11342,N_11357);
xnor U18115 (N_18115,N_12655,N_14174);
or U18116 (N_18116,N_13497,N_12289);
and U18117 (N_18117,N_12092,N_14826);
or U18118 (N_18118,N_11383,N_10211);
nand U18119 (N_18119,N_12018,N_14808);
xnor U18120 (N_18120,N_13016,N_14283);
nand U18121 (N_18121,N_11558,N_14899);
nor U18122 (N_18122,N_10238,N_11639);
nand U18123 (N_18123,N_11262,N_13540);
or U18124 (N_18124,N_13275,N_12550);
or U18125 (N_18125,N_10485,N_11280);
and U18126 (N_18126,N_13757,N_14113);
nor U18127 (N_18127,N_14617,N_11265);
xnor U18128 (N_18128,N_12746,N_13380);
nor U18129 (N_18129,N_11289,N_13072);
nor U18130 (N_18130,N_14598,N_11146);
and U18131 (N_18131,N_11885,N_10471);
nor U18132 (N_18132,N_11888,N_12683);
nor U18133 (N_18133,N_10728,N_14695);
or U18134 (N_18134,N_13544,N_10260);
nand U18135 (N_18135,N_11134,N_11756);
and U18136 (N_18136,N_12576,N_12173);
and U18137 (N_18137,N_13690,N_11672);
or U18138 (N_18138,N_11493,N_14093);
nor U18139 (N_18139,N_11743,N_13383);
and U18140 (N_18140,N_13226,N_11656);
nor U18141 (N_18141,N_12548,N_14624);
nand U18142 (N_18142,N_11933,N_11068);
nand U18143 (N_18143,N_12336,N_10418);
nor U18144 (N_18144,N_11305,N_12727);
nor U18145 (N_18145,N_10937,N_14255);
nor U18146 (N_18146,N_13862,N_12336);
nand U18147 (N_18147,N_14929,N_14977);
or U18148 (N_18148,N_12652,N_13497);
nor U18149 (N_18149,N_12869,N_10608);
nor U18150 (N_18150,N_13416,N_11314);
or U18151 (N_18151,N_10771,N_13933);
and U18152 (N_18152,N_14473,N_12336);
nor U18153 (N_18153,N_12335,N_12405);
or U18154 (N_18154,N_11969,N_14253);
or U18155 (N_18155,N_12206,N_10320);
nand U18156 (N_18156,N_12500,N_12125);
or U18157 (N_18157,N_13214,N_10248);
xnor U18158 (N_18158,N_13027,N_10752);
or U18159 (N_18159,N_13558,N_11835);
and U18160 (N_18160,N_13652,N_14126);
xnor U18161 (N_18161,N_13882,N_13642);
and U18162 (N_18162,N_13480,N_14661);
and U18163 (N_18163,N_10841,N_14270);
xnor U18164 (N_18164,N_10207,N_12234);
nand U18165 (N_18165,N_10536,N_10551);
or U18166 (N_18166,N_13925,N_10427);
xor U18167 (N_18167,N_12193,N_14741);
and U18168 (N_18168,N_14518,N_10163);
nand U18169 (N_18169,N_10614,N_12484);
xnor U18170 (N_18170,N_12856,N_11174);
or U18171 (N_18171,N_10298,N_13183);
and U18172 (N_18172,N_11972,N_13191);
nand U18173 (N_18173,N_14537,N_13632);
nor U18174 (N_18174,N_14529,N_12995);
xor U18175 (N_18175,N_12913,N_14384);
and U18176 (N_18176,N_12964,N_11101);
nor U18177 (N_18177,N_11617,N_14409);
xnor U18178 (N_18178,N_10301,N_11359);
xor U18179 (N_18179,N_13293,N_11980);
or U18180 (N_18180,N_10112,N_10575);
or U18181 (N_18181,N_12540,N_11250);
nor U18182 (N_18182,N_11445,N_10706);
or U18183 (N_18183,N_12245,N_10310);
or U18184 (N_18184,N_10252,N_11558);
and U18185 (N_18185,N_12870,N_14555);
nor U18186 (N_18186,N_14173,N_14846);
nor U18187 (N_18187,N_12743,N_12395);
xnor U18188 (N_18188,N_10051,N_13191);
nor U18189 (N_18189,N_14799,N_10178);
xnor U18190 (N_18190,N_14094,N_12558);
xor U18191 (N_18191,N_11188,N_12393);
nor U18192 (N_18192,N_10782,N_14425);
nand U18193 (N_18193,N_11182,N_14849);
nor U18194 (N_18194,N_10297,N_13852);
or U18195 (N_18195,N_14185,N_11062);
nor U18196 (N_18196,N_10066,N_10809);
and U18197 (N_18197,N_11033,N_12793);
or U18198 (N_18198,N_12569,N_10185);
and U18199 (N_18199,N_14097,N_10206);
and U18200 (N_18200,N_10614,N_13417);
nor U18201 (N_18201,N_12383,N_10950);
xor U18202 (N_18202,N_13486,N_11569);
nor U18203 (N_18203,N_11304,N_10819);
xor U18204 (N_18204,N_12596,N_10522);
nor U18205 (N_18205,N_14758,N_14829);
and U18206 (N_18206,N_12307,N_10073);
nand U18207 (N_18207,N_10208,N_13158);
nand U18208 (N_18208,N_12828,N_12893);
xnor U18209 (N_18209,N_11999,N_12573);
nand U18210 (N_18210,N_10874,N_13641);
and U18211 (N_18211,N_14074,N_10409);
or U18212 (N_18212,N_14098,N_10853);
or U18213 (N_18213,N_11689,N_10209);
nor U18214 (N_18214,N_11700,N_11432);
xnor U18215 (N_18215,N_13062,N_11238);
nor U18216 (N_18216,N_10401,N_14325);
nand U18217 (N_18217,N_13446,N_11007);
xor U18218 (N_18218,N_13943,N_11709);
nor U18219 (N_18219,N_13451,N_14899);
xnor U18220 (N_18220,N_13862,N_10843);
or U18221 (N_18221,N_13309,N_13333);
and U18222 (N_18222,N_14295,N_12969);
xnor U18223 (N_18223,N_11772,N_10767);
and U18224 (N_18224,N_14016,N_13370);
or U18225 (N_18225,N_12252,N_14210);
and U18226 (N_18226,N_11978,N_10904);
or U18227 (N_18227,N_11411,N_13780);
or U18228 (N_18228,N_13623,N_11335);
nor U18229 (N_18229,N_12043,N_10220);
or U18230 (N_18230,N_12321,N_10082);
or U18231 (N_18231,N_12514,N_13448);
xor U18232 (N_18232,N_11725,N_14555);
xor U18233 (N_18233,N_12073,N_12974);
xnor U18234 (N_18234,N_13448,N_10671);
and U18235 (N_18235,N_14373,N_13750);
or U18236 (N_18236,N_11177,N_10985);
xnor U18237 (N_18237,N_10792,N_13040);
or U18238 (N_18238,N_11617,N_10645);
and U18239 (N_18239,N_10763,N_14300);
and U18240 (N_18240,N_13011,N_11003);
xnor U18241 (N_18241,N_12410,N_14383);
xnor U18242 (N_18242,N_10577,N_12531);
and U18243 (N_18243,N_12703,N_11416);
nand U18244 (N_18244,N_11061,N_12241);
nor U18245 (N_18245,N_11991,N_10515);
xor U18246 (N_18246,N_10231,N_11649);
and U18247 (N_18247,N_13318,N_13892);
and U18248 (N_18248,N_12759,N_12037);
or U18249 (N_18249,N_13085,N_11064);
nand U18250 (N_18250,N_11321,N_11306);
and U18251 (N_18251,N_11076,N_12707);
or U18252 (N_18252,N_13863,N_10025);
and U18253 (N_18253,N_12108,N_13079);
or U18254 (N_18254,N_14700,N_10611);
or U18255 (N_18255,N_13922,N_14613);
nand U18256 (N_18256,N_10360,N_10404);
nor U18257 (N_18257,N_13958,N_12257);
or U18258 (N_18258,N_11156,N_12940);
and U18259 (N_18259,N_10247,N_12697);
or U18260 (N_18260,N_11864,N_10015);
xnor U18261 (N_18261,N_10770,N_12757);
xnor U18262 (N_18262,N_10826,N_10299);
or U18263 (N_18263,N_13416,N_11794);
and U18264 (N_18264,N_12462,N_12083);
nand U18265 (N_18265,N_14987,N_10700);
nor U18266 (N_18266,N_10835,N_12870);
nor U18267 (N_18267,N_13686,N_12381);
and U18268 (N_18268,N_14022,N_10767);
and U18269 (N_18269,N_10963,N_12436);
xor U18270 (N_18270,N_12034,N_12922);
or U18271 (N_18271,N_11735,N_10277);
xnor U18272 (N_18272,N_10575,N_14685);
nor U18273 (N_18273,N_10926,N_11319);
nor U18274 (N_18274,N_13954,N_11735);
nor U18275 (N_18275,N_14642,N_14867);
nand U18276 (N_18276,N_12116,N_13902);
xnor U18277 (N_18277,N_10012,N_11170);
or U18278 (N_18278,N_14642,N_11797);
and U18279 (N_18279,N_14615,N_10921);
xnor U18280 (N_18280,N_12247,N_14217);
nand U18281 (N_18281,N_13271,N_14853);
and U18282 (N_18282,N_13599,N_10310);
nand U18283 (N_18283,N_11496,N_11802);
nor U18284 (N_18284,N_11918,N_11461);
xor U18285 (N_18285,N_13872,N_14031);
xnor U18286 (N_18286,N_14048,N_12646);
nor U18287 (N_18287,N_13651,N_13794);
nand U18288 (N_18288,N_11220,N_13926);
and U18289 (N_18289,N_10636,N_11947);
nand U18290 (N_18290,N_12473,N_12096);
nand U18291 (N_18291,N_13009,N_13864);
or U18292 (N_18292,N_12115,N_10474);
nor U18293 (N_18293,N_10218,N_14141);
xnor U18294 (N_18294,N_14416,N_10361);
and U18295 (N_18295,N_11556,N_10279);
xnor U18296 (N_18296,N_10434,N_12083);
and U18297 (N_18297,N_11751,N_10248);
nand U18298 (N_18298,N_11267,N_11078);
nand U18299 (N_18299,N_10901,N_14901);
nor U18300 (N_18300,N_13826,N_13593);
nor U18301 (N_18301,N_12075,N_11601);
nand U18302 (N_18302,N_14297,N_12270);
nand U18303 (N_18303,N_11454,N_10340);
nand U18304 (N_18304,N_14459,N_14355);
nor U18305 (N_18305,N_12357,N_13943);
nor U18306 (N_18306,N_10480,N_13804);
nand U18307 (N_18307,N_12579,N_14779);
nor U18308 (N_18308,N_12590,N_14196);
nand U18309 (N_18309,N_14188,N_10441);
nor U18310 (N_18310,N_13749,N_12981);
nor U18311 (N_18311,N_12398,N_12754);
xor U18312 (N_18312,N_14627,N_11161);
nor U18313 (N_18313,N_12664,N_13137);
and U18314 (N_18314,N_14583,N_11267);
nand U18315 (N_18315,N_10371,N_12113);
and U18316 (N_18316,N_10741,N_11904);
and U18317 (N_18317,N_12064,N_10071);
nor U18318 (N_18318,N_13037,N_12513);
nor U18319 (N_18319,N_14970,N_13484);
or U18320 (N_18320,N_10277,N_11553);
and U18321 (N_18321,N_12662,N_13190);
and U18322 (N_18322,N_10744,N_13515);
and U18323 (N_18323,N_13628,N_11070);
or U18324 (N_18324,N_10450,N_12299);
and U18325 (N_18325,N_11231,N_11357);
and U18326 (N_18326,N_14004,N_11241);
xnor U18327 (N_18327,N_11299,N_13657);
or U18328 (N_18328,N_10013,N_11562);
xnor U18329 (N_18329,N_13281,N_13825);
nand U18330 (N_18330,N_10278,N_11202);
nand U18331 (N_18331,N_10276,N_12689);
nor U18332 (N_18332,N_13567,N_12249);
nand U18333 (N_18333,N_10303,N_12685);
or U18334 (N_18334,N_10434,N_13085);
or U18335 (N_18335,N_10556,N_11639);
nand U18336 (N_18336,N_11025,N_11288);
and U18337 (N_18337,N_10197,N_10296);
nand U18338 (N_18338,N_14668,N_14808);
or U18339 (N_18339,N_13256,N_14741);
nand U18340 (N_18340,N_10587,N_13222);
xor U18341 (N_18341,N_10511,N_14099);
nand U18342 (N_18342,N_13607,N_11711);
and U18343 (N_18343,N_13088,N_12933);
and U18344 (N_18344,N_13558,N_11071);
nand U18345 (N_18345,N_14910,N_13794);
xnor U18346 (N_18346,N_10654,N_10532);
or U18347 (N_18347,N_10255,N_12498);
nor U18348 (N_18348,N_10783,N_13761);
and U18349 (N_18349,N_10506,N_13708);
nor U18350 (N_18350,N_11675,N_13166);
nor U18351 (N_18351,N_14395,N_12517);
nor U18352 (N_18352,N_12021,N_10246);
nor U18353 (N_18353,N_13855,N_12413);
or U18354 (N_18354,N_12159,N_14594);
and U18355 (N_18355,N_10915,N_13524);
nor U18356 (N_18356,N_13596,N_10777);
or U18357 (N_18357,N_14951,N_12438);
and U18358 (N_18358,N_12644,N_13420);
and U18359 (N_18359,N_12819,N_10554);
xor U18360 (N_18360,N_12573,N_12983);
and U18361 (N_18361,N_14363,N_12152);
xnor U18362 (N_18362,N_10213,N_10991);
xnor U18363 (N_18363,N_10812,N_10880);
nand U18364 (N_18364,N_10448,N_12220);
and U18365 (N_18365,N_14712,N_10492);
nor U18366 (N_18366,N_11500,N_11949);
or U18367 (N_18367,N_12321,N_10176);
nor U18368 (N_18368,N_13077,N_14823);
nand U18369 (N_18369,N_11973,N_13088);
nor U18370 (N_18370,N_13458,N_13147);
xor U18371 (N_18371,N_12539,N_11639);
nor U18372 (N_18372,N_13787,N_11789);
nor U18373 (N_18373,N_13218,N_13081);
nand U18374 (N_18374,N_11183,N_11427);
and U18375 (N_18375,N_11036,N_11838);
nor U18376 (N_18376,N_13923,N_12456);
or U18377 (N_18377,N_13450,N_11171);
nor U18378 (N_18378,N_14391,N_11459);
and U18379 (N_18379,N_10644,N_13100);
nor U18380 (N_18380,N_10847,N_12474);
or U18381 (N_18381,N_14523,N_12765);
nor U18382 (N_18382,N_10536,N_14143);
xnor U18383 (N_18383,N_12546,N_11229);
nor U18384 (N_18384,N_14924,N_12888);
or U18385 (N_18385,N_13938,N_13202);
nor U18386 (N_18386,N_11536,N_11210);
or U18387 (N_18387,N_11172,N_10578);
nor U18388 (N_18388,N_12492,N_10891);
and U18389 (N_18389,N_11851,N_12730);
nor U18390 (N_18390,N_11353,N_11834);
or U18391 (N_18391,N_12046,N_10939);
and U18392 (N_18392,N_10768,N_12238);
nand U18393 (N_18393,N_11594,N_10439);
xor U18394 (N_18394,N_12407,N_11252);
nand U18395 (N_18395,N_10255,N_11022);
xor U18396 (N_18396,N_12364,N_11917);
and U18397 (N_18397,N_11029,N_10441);
and U18398 (N_18398,N_14387,N_14422);
or U18399 (N_18399,N_13210,N_12969);
nor U18400 (N_18400,N_12777,N_12670);
and U18401 (N_18401,N_11634,N_14681);
or U18402 (N_18402,N_11270,N_10487);
nand U18403 (N_18403,N_14983,N_12948);
and U18404 (N_18404,N_12422,N_13313);
or U18405 (N_18405,N_10618,N_12596);
nand U18406 (N_18406,N_10709,N_10838);
and U18407 (N_18407,N_13324,N_12091);
or U18408 (N_18408,N_14761,N_10611);
xnor U18409 (N_18409,N_10508,N_12491);
nand U18410 (N_18410,N_12994,N_10766);
nand U18411 (N_18411,N_10321,N_10909);
and U18412 (N_18412,N_11114,N_11435);
and U18413 (N_18413,N_12346,N_13542);
or U18414 (N_18414,N_13608,N_13108);
and U18415 (N_18415,N_10582,N_14394);
nor U18416 (N_18416,N_12201,N_12401);
nor U18417 (N_18417,N_13107,N_14018);
and U18418 (N_18418,N_14751,N_10143);
nor U18419 (N_18419,N_13992,N_12718);
nand U18420 (N_18420,N_12241,N_11805);
nor U18421 (N_18421,N_13878,N_12787);
xnor U18422 (N_18422,N_14535,N_13730);
nor U18423 (N_18423,N_10572,N_14962);
nand U18424 (N_18424,N_13915,N_14672);
or U18425 (N_18425,N_14386,N_11054);
and U18426 (N_18426,N_10379,N_12371);
or U18427 (N_18427,N_12403,N_10717);
xor U18428 (N_18428,N_14991,N_11315);
or U18429 (N_18429,N_10291,N_14680);
and U18430 (N_18430,N_14734,N_12826);
xnor U18431 (N_18431,N_11799,N_11685);
nor U18432 (N_18432,N_14256,N_11801);
xor U18433 (N_18433,N_10113,N_13920);
xor U18434 (N_18434,N_10372,N_13602);
nand U18435 (N_18435,N_11595,N_10044);
or U18436 (N_18436,N_11887,N_14806);
nand U18437 (N_18437,N_10648,N_13223);
nor U18438 (N_18438,N_12793,N_12932);
xor U18439 (N_18439,N_11092,N_12814);
nor U18440 (N_18440,N_10641,N_11687);
or U18441 (N_18441,N_10746,N_11296);
nor U18442 (N_18442,N_12630,N_14449);
nand U18443 (N_18443,N_13432,N_10914);
xnor U18444 (N_18444,N_14570,N_11675);
nor U18445 (N_18445,N_13559,N_12984);
nand U18446 (N_18446,N_10550,N_10324);
nor U18447 (N_18447,N_10967,N_14970);
nor U18448 (N_18448,N_11096,N_11442);
xor U18449 (N_18449,N_12548,N_13700);
nand U18450 (N_18450,N_11916,N_14171);
nand U18451 (N_18451,N_10576,N_10020);
or U18452 (N_18452,N_12002,N_11646);
xor U18453 (N_18453,N_12958,N_11882);
and U18454 (N_18454,N_11035,N_14286);
or U18455 (N_18455,N_12903,N_13724);
nor U18456 (N_18456,N_10767,N_13951);
nor U18457 (N_18457,N_14183,N_12863);
and U18458 (N_18458,N_11199,N_11289);
nor U18459 (N_18459,N_10437,N_10562);
and U18460 (N_18460,N_13139,N_13214);
nand U18461 (N_18461,N_14878,N_11583);
xnor U18462 (N_18462,N_14699,N_14656);
or U18463 (N_18463,N_13508,N_10827);
or U18464 (N_18464,N_11166,N_12791);
nand U18465 (N_18465,N_13190,N_13572);
nor U18466 (N_18466,N_11807,N_14903);
nor U18467 (N_18467,N_11387,N_14661);
xnor U18468 (N_18468,N_10666,N_10066);
xnor U18469 (N_18469,N_14818,N_14017);
xnor U18470 (N_18470,N_11929,N_14741);
and U18471 (N_18471,N_10277,N_10050);
or U18472 (N_18472,N_14367,N_12136);
nand U18473 (N_18473,N_11609,N_14149);
xnor U18474 (N_18474,N_10795,N_13452);
nand U18475 (N_18475,N_14621,N_10819);
or U18476 (N_18476,N_10049,N_14057);
nand U18477 (N_18477,N_12939,N_12006);
xnor U18478 (N_18478,N_11217,N_12451);
xnor U18479 (N_18479,N_10736,N_12065);
nor U18480 (N_18480,N_10974,N_12978);
nor U18481 (N_18481,N_14333,N_10586);
xnor U18482 (N_18482,N_10682,N_10535);
or U18483 (N_18483,N_14693,N_13593);
xor U18484 (N_18484,N_12006,N_12304);
and U18485 (N_18485,N_10447,N_11956);
nand U18486 (N_18486,N_11018,N_14054);
or U18487 (N_18487,N_10295,N_12285);
nand U18488 (N_18488,N_14849,N_13458);
nor U18489 (N_18489,N_12849,N_14694);
or U18490 (N_18490,N_12493,N_13281);
nand U18491 (N_18491,N_10705,N_14853);
xnor U18492 (N_18492,N_11009,N_11640);
or U18493 (N_18493,N_12948,N_13842);
nor U18494 (N_18494,N_14621,N_14667);
xor U18495 (N_18495,N_13339,N_10919);
or U18496 (N_18496,N_14526,N_14995);
or U18497 (N_18497,N_14444,N_11446);
nor U18498 (N_18498,N_12929,N_11271);
and U18499 (N_18499,N_13127,N_14188);
and U18500 (N_18500,N_10739,N_14104);
and U18501 (N_18501,N_13209,N_10119);
and U18502 (N_18502,N_14331,N_13944);
nand U18503 (N_18503,N_11103,N_12293);
nor U18504 (N_18504,N_10330,N_10000);
or U18505 (N_18505,N_14984,N_13384);
or U18506 (N_18506,N_14525,N_13139);
nand U18507 (N_18507,N_11801,N_10092);
nor U18508 (N_18508,N_12813,N_11537);
or U18509 (N_18509,N_11673,N_11679);
and U18510 (N_18510,N_14603,N_13311);
xnor U18511 (N_18511,N_14862,N_11532);
or U18512 (N_18512,N_14947,N_10184);
nor U18513 (N_18513,N_13300,N_10556);
xnor U18514 (N_18514,N_10031,N_11410);
nand U18515 (N_18515,N_11982,N_10393);
nor U18516 (N_18516,N_14350,N_13368);
and U18517 (N_18517,N_13434,N_10954);
nor U18518 (N_18518,N_14733,N_12761);
xnor U18519 (N_18519,N_14136,N_14516);
and U18520 (N_18520,N_14651,N_10434);
nor U18521 (N_18521,N_13850,N_12228);
nor U18522 (N_18522,N_10937,N_13091);
xor U18523 (N_18523,N_14028,N_12028);
xnor U18524 (N_18524,N_14219,N_12260);
xnor U18525 (N_18525,N_11882,N_13369);
or U18526 (N_18526,N_12872,N_11057);
and U18527 (N_18527,N_13441,N_13294);
or U18528 (N_18528,N_13211,N_14108);
or U18529 (N_18529,N_13202,N_11311);
nor U18530 (N_18530,N_13685,N_12513);
nor U18531 (N_18531,N_10723,N_12010);
and U18532 (N_18532,N_11180,N_10640);
or U18533 (N_18533,N_12555,N_10435);
nand U18534 (N_18534,N_10313,N_14420);
xor U18535 (N_18535,N_13688,N_10464);
nor U18536 (N_18536,N_13662,N_11198);
and U18537 (N_18537,N_11452,N_12422);
xnor U18538 (N_18538,N_10148,N_14270);
or U18539 (N_18539,N_13066,N_13692);
nand U18540 (N_18540,N_12380,N_12051);
or U18541 (N_18541,N_11693,N_12349);
nor U18542 (N_18542,N_12739,N_12865);
nor U18543 (N_18543,N_11587,N_14982);
or U18544 (N_18544,N_10632,N_10905);
nor U18545 (N_18545,N_14951,N_14912);
nand U18546 (N_18546,N_10997,N_14033);
or U18547 (N_18547,N_14633,N_11402);
and U18548 (N_18548,N_11218,N_10748);
and U18549 (N_18549,N_10393,N_12645);
nand U18550 (N_18550,N_11757,N_13431);
or U18551 (N_18551,N_12780,N_13524);
nand U18552 (N_18552,N_13613,N_11576);
xnor U18553 (N_18553,N_13895,N_13815);
or U18554 (N_18554,N_11793,N_13766);
and U18555 (N_18555,N_11828,N_12820);
nor U18556 (N_18556,N_11386,N_14252);
and U18557 (N_18557,N_14399,N_10063);
nor U18558 (N_18558,N_12815,N_11481);
nand U18559 (N_18559,N_13227,N_13920);
nand U18560 (N_18560,N_11622,N_10985);
and U18561 (N_18561,N_14666,N_11828);
nor U18562 (N_18562,N_14520,N_11423);
or U18563 (N_18563,N_13149,N_14411);
or U18564 (N_18564,N_13314,N_10673);
nor U18565 (N_18565,N_12425,N_14392);
nor U18566 (N_18566,N_14820,N_13449);
or U18567 (N_18567,N_11839,N_10124);
xor U18568 (N_18568,N_10304,N_14349);
nor U18569 (N_18569,N_14462,N_12009);
xnor U18570 (N_18570,N_11870,N_10996);
nor U18571 (N_18571,N_14711,N_13750);
xnor U18572 (N_18572,N_10306,N_11198);
nor U18573 (N_18573,N_11065,N_12937);
and U18574 (N_18574,N_13568,N_11242);
nor U18575 (N_18575,N_13502,N_10446);
nor U18576 (N_18576,N_11473,N_12681);
and U18577 (N_18577,N_12925,N_10018);
nand U18578 (N_18578,N_13627,N_10558);
nor U18579 (N_18579,N_11579,N_13827);
xnor U18580 (N_18580,N_12288,N_14929);
nand U18581 (N_18581,N_11096,N_11013);
and U18582 (N_18582,N_13847,N_12722);
xnor U18583 (N_18583,N_13660,N_10523);
or U18584 (N_18584,N_14031,N_12845);
xnor U18585 (N_18585,N_14151,N_12830);
nand U18586 (N_18586,N_10806,N_12519);
xor U18587 (N_18587,N_14589,N_13105);
xor U18588 (N_18588,N_12492,N_11892);
or U18589 (N_18589,N_14531,N_11921);
or U18590 (N_18590,N_12900,N_10261);
or U18591 (N_18591,N_12994,N_11928);
nand U18592 (N_18592,N_14898,N_11315);
nor U18593 (N_18593,N_13419,N_13386);
or U18594 (N_18594,N_12056,N_14230);
xor U18595 (N_18595,N_13633,N_13575);
or U18596 (N_18596,N_10508,N_12588);
nor U18597 (N_18597,N_11307,N_14660);
and U18598 (N_18598,N_12281,N_13743);
and U18599 (N_18599,N_11759,N_14159);
xor U18600 (N_18600,N_10541,N_11263);
nor U18601 (N_18601,N_12048,N_11100);
nand U18602 (N_18602,N_12610,N_13085);
xnor U18603 (N_18603,N_12679,N_11591);
xnor U18604 (N_18604,N_11099,N_14238);
xor U18605 (N_18605,N_12252,N_13660);
nor U18606 (N_18606,N_14701,N_10697);
and U18607 (N_18607,N_14041,N_11564);
xor U18608 (N_18608,N_14110,N_14335);
nor U18609 (N_18609,N_12524,N_11486);
or U18610 (N_18610,N_10640,N_10039);
or U18611 (N_18611,N_12128,N_12889);
xnor U18612 (N_18612,N_13600,N_12916);
and U18613 (N_18613,N_12668,N_14423);
and U18614 (N_18614,N_11888,N_14231);
and U18615 (N_18615,N_11200,N_10490);
and U18616 (N_18616,N_10444,N_13859);
xnor U18617 (N_18617,N_12727,N_11226);
and U18618 (N_18618,N_13739,N_11953);
xor U18619 (N_18619,N_10886,N_14389);
xnor U18620 (N_18620,N_11071,N_11293);
or U18621 (N_18621,N_14681,N_14336);
nor U18622 (N_18622,N_11089,N_14943);
nor U18623 (N_18623,N_14720,N_13844);
xnor U18624 (N_18624,N_12756,N_10185);
nand U18625 (N_18625,N_14218,N_10894);
nor U18626 (N_18626,N_11186,N_14330);
xor U18627 (N_18627,N_10924,N_14865);
xor U18628 (N_18628,N_10290,N_10663);
xnor U18629 (N_18629,N_14375,N_12418);
nor U18630 (N_18630,N_12535,N_14583);
and U18631 (N_18631,N_11254,N_10743);
xnor U18632 (N_18632,N_13255,N_12074);
nand U18633 (N_18633,N_11618,N_10924);
xor U18634 (N_18634,N_14611,N_14038);
xnor U18635 (N_18635,N_13727,N_13159);
nor U18636 (N_18636,N_12980,N_11762);
xor U18637 (N_18637,N_10253,N_11340);
nand U18638 (N_18638,N_13127,N_14918);
xor U18639 (N_18639,N_11466,N_13465);
nor U18640 (N_18640,N_13458,N_14327);
and U18641 (N_18641,N_10596,N_11944);
and U18642 (N_18642,N_11965,N_14053);
xnor U18643 (N_18643,N_14941,N_11696);
nor U18644 (N_18644,N_14665,N_10969);
or U18645 (N_18645,N_12745,N_11643);
or U18646 (N_18646,N_14608,N_12376);
or U18647 (N_18647,N_13124,N_11977);
xnor U18648 (N_18648,N_11598,N_14691);
and U18649 (N_18649,N_11568,N_13547);
nor U18650 (N_18650,N_12059,N_12664);
nand U18651 (N_18651,N_10568,N_11811);
and U18652 (N_18652,N_13465,N_12506);
xor U18653 (N_18653,N_14639,N_10793);
xor U18654 (N_18654,N_10121,N_10837);
or U18655 (N_18655,N_10859,N_12938);
and U18656 (N_18656,N_14884,N_12540);
nand U18657 (N_18657,N_12283,N_12192);
nor U18658 (N_18658,N_14940,N_14345);
nand U18659 (N_18659,N_11290,N_14143);
nand U18660 (N_18660,N_10665,N_12177);
nand U18661 (N_18661,N_12626,N_12333);
xor U18662 (N_18662,N_14901,N_13333);
or U18663 (N_18663,N_10455,N_12201);
or U18664 (N_18664,N_10204,N_14848);
xor U18665 (N_18665,N_11195,N_12772);
xnor U18666 (N_18666,N_11883,N_12478);
and U18667 (N_18667,N_13718,N_10203);
nand U18668 (N_18668,N_10624,N_14233);
and U18669 (N_18669,N_14509,N_14219);
nor U18670 (N_18670,N_13066,N_13891);
nor U18671 (N_18671,N_14065,N_11929);
xor U18672 (N_18672,N_13658,N_14622);
or U18673 (N_18673,N_10318,N_12146);
nand U18674 (N_18674,N_11979,N_11632);
or U18675 (N_18675,N_13198,N_10509);
or U18676 (N_18676,N_13057,N_11637);
nor U18677 (N_18677,N_11721,N_13518);
or U18678 (N_18678,N_10325,N_13511);
nor U18679 (N_18679,N_14093,N_13911);
nor U18680 (N_18680,N_12010,N_11225);
xnor U18681 (N_18681,N_13029,N_14665);
xor U18682 (N_18682,N_11664,N_14489);
or U18683 (N_18683,N_10335,N_12775);
and U18684 (N_18684,N_11452,N_10437);
nand U18685 (N_18685,N_14045,N_12673);
xnor U18686 (N_18686,N_12702,N_13800);
or U18687 (N_18687,N_14443,N_13030);
nor U18688 (N_18688,N_10296,N_11419);
nor U18689 (N_18689,N_10869,N_14532);
nand U18690 (N_18690,N_14256,N_14876);
and U18691 (N_18691,N_10528,N_10479);
or U18692 (N_18692,N_11075,N_12929);
nor U18693 (N_18693,N_10737,N_14441);
or U18694 (N_18694,N_11230,N_14699);
xnor U18695 (N_18695,N_10697,N_14492);
nand U18696 (N_18696,N_14831,N_11705);
and U18697 (N_18697,N_11792,N_11753);
nor U18698 (N_18698,N_14259,N_12910);
nor U18699 (N_18699,N_10551,N_11404);
nor U18700 (N_18700,N_11941,N_11277);
or U18701 (N_18701,N_11736,N_12125);
xor U18702 (N_18702,N_13002,N_11122);
or U18703 (N_18703,N_12945,N_11024);
nor U18704 (N_18704,N_10728,N_13759);
nand U18705 (N_18705,N_12248,N_13157);
nor U18706 (N_18706,N_14839,N_11513);
nand U18707 (N_18707,N_14517,N_11420);
nor U18708 (N_18708,N_11243,N_13051);
nor U18709 (N_18709,N_12003,N_12214);
or U18710 (N_18710,N_11842,N_10945);
nand U18711 (N_18711,N_13163,N_10035);
nor U18712 (N_18712,N_14044,N_12057);
or U18713 (N_18713,N_11830,N_12915);
nor U18714 (N_18714,N_10911,N_11827);
xor U18715 (N_18715,N_12731,N_14523);
nor U18716 (N_18716,N_13640,N_12708);
nor U18717 (N_18717,N_13261,N_12854);
or U18718 (N_18718,N_10083,N_11616);
nor U18719 (N_18719,N_13218,N_13484);
xnor U18720 (N_18720,N_10778,N_10021);
xnor U18721 (N_18721,N_12002,N_13943);
nor U18722 (N_18722,N_14500,N_13324);
xnor U18723 (N_18723,N_13396,N_13621);
nand U18724 (N_18724,N_10144,N_13391);
xor U18725 (N_18725,N_13528,N_13650);
nand U18726 (N_18726,N_11666,N_12323);
nand U18727 (N_18727,N_14390,N_10809);
nor U18728 (N_18728,N_11281,N_13209);
nor U18729 (N_18729,N_14768,N_14801);
nand U18730 (N_18730,N_12764,N_14518);
and U18731 (N_18731,N_12497,N_13064);
nand U18732 (N_18732,N_13513,N_14293);
nor U18733 (N_18733,N_13492,N_13105);
xnor U18734 (N_18734,N_11255,N_10593);
or U18735 (N_18735,N_12806,N_12551);
or U18736 (N_18736,N_13738,N_13982);
or U18737 (N_18737,N_11999,N_11646);
and U18738 (N_18738,N_10545,N_13164);
xnor U18739 (N_18739,N_11233,N_10907);
and U18740 (N_18740,N_13760,N_11299);
and U18741 (N_18741,N_12763,N_14774);
nand U18742 (N_18742,N_10433,N_10315);
or U18743 (N_18743,N_13107,N_11587);
nand U18744 (N_18744,N_10353,N_13072);
nor U18745 (N_18745,N_14791,N_12521);
and U18746 (N_18746,N_11620,N_13874);
and U18747 (N_18747,N_12564,N_12116);
nor U18748 (N_18748,N_10255,N_10469);
nand U18749 (N_18749,N_10409,N_13619);
and U18750 (N_18750,N_10732,N_13275);
and U18751 (N_18751,N_10999,N_12826);
nor U18752 (N_18752,N_14392,N_14447);
nor U18753 (N_18753,N_12118,N_13640);
and U18754 (N_18754,N_11312,N_12692);
nand U18755 (N_18755,N_14160,N_10574);
nor U18756 (N_18756,N_13603,N_11656);
nand U18757 (N_18757,N_11817,N_10294);
nor U18758 (N_18758,N_13135,N_14470);
or U18759 (N_18759,N_11211,N_13010);
or U18760 (N_18760,N_11522,N_12271);
nor U18761 (N_18761,N_10845,N_14448);
or U18762 (N_18762,N_13718,N_11606);
nor U18763 (N_18763,N_10780,N_14051);
nand U18764 (N_18764,N_11895,N_11316);
and U18765 (N_18765,N_10996,N_14934);
nor U18766 (N_18766,N_13578,N_13569);
nor U18767 (N_18767,N_12754,N_14153);
xnor U18768 (N_18768,N_14960,N_12521);
nor U18769 (N_18769,N_10510,N_11058);
or U18770 (N_18770,N_12129,N_10536);
xnor U18771 (N_18771,N_10016,N_14752);
nor U18772 (N_18772,N_10509,N_13788);
nor U18773 (N_18773,N_14596,N_11587);
nand U18774 (N_18774,N_11356,N_13155);
xor U18775 (N_18775,N_13467,N_14429);
or U18776 (N_18776,N_13459,N_14414);
and U18777 (N_18777,N_11488,N_14982);
nor U18778 (N_18778,N_11297,N_12635);
or U18779 (N_18779,N_12405,N_10348);
and U18780 (N_18780,N_10670,N_14322);
xor U18781 (N_18781,N_10455,N_11472);
nand U18782 (N_18782,N_13760,N_11637);
nand U18783 (N_18783,N_13067,N_11908);
or U18784 (N_18784,N_12168,N_13400);
or U18785 (N_18785,N_10061,N_10545);
nor U18786 (N_18786,N_14220,N_14135);
nand U18787 (N_18787,N_11265,N_11898);
nand U18788 (N_18788,N_14524,N_13897);
xor U18789 (N_18789,N_10903,N_14335);
nor U18790 (N_18790,N_12891,N_14746);
nand U18791 (N_18791,N_12887,N_13519);
or U18792 (N_18792,N_13306,N_12921);
or U18793 (N_18793,N_13914,N_10101);
and U18794 (N_18794,N_12409,N_14544);
nor U18795 (N_18795,N_13710,N_11585);
xnor U18796 (N_18796,N_13998,N_10396);
and U18797 (N_18797,N_12189,N_13713);
and U18798 (N_18798,N_13929,N_10991);
xnor U18799 (N_18799,N_12782,N_13818);
or U18800 (N_18800,N_12884,N_12012);
and U18801 (N_18801,N_14802,N_12642);
xor U18802 (N_18802,N_13013,N_10587);
and U18803 (N_18803,N_10475,N_14628);
and U18804 (N_18804,N_14875,N_11209);
nand U18805 (N_18805,N_13284,N_12186);
xor U18806 (N_18806,N_10508,N_14717);
or U18807 (N_18807,N_10838,N_10330);
xor U18808 (N_18808,N_12165,N_11127);
xor U18809 (N_18809,N_13064,N_13364);
nand U18810 (N_18810,N_13241,N_13974);
or U18811 (N_18811,N_11896,N_14218);
or U18812 (N_18812,N_11346,N_14666);
and U18813 (N_18813,N_11481,N_11262);
and U18814 (N_18814,N_14642,N_11508);
xnor U18815 (N_18815,N_12846,N_11176);
nor U18816 (N_18816,N_13171,N_13912);
or U18817 (N_18817,N_12167,N_12003);
xnor U18818 (N_18818,N_13296,N_13343);
nand U18819 (N_18819,N_10107,N_12540);
or U18820 (N_18820,N_11567,N_11751);
xor U18821 (N_18821,N_14567,N_12222);
nand U18822 (N_18822,N_10051,N_13405);
or U18823 (N_18823,N_11636,N_11512);
nand U18824 (N_18824,N_10132,N_10554);
nand U18825 (N_18825,N_11891,N_10436);
or U18826 (N_18826,N_10236,N_10702);
nand U18827 (N_18827,N_13154,N_11126);
nor U18828 (N_18828,N_13151,N_11647);
and U18829 (N_18829,N_11629,N_14778);
or U18830 (N_18830,N_11482,N_12930);
and U18831 (N_18831,N_12921,N_11075);
or U18832 (N_18832,N_13584,N_11147);
nor U18833 (N_18833,N_13374,N_12377);
and U18834 (N_18834,N_12550,N_11825);
and U18835 (N_18835,N_10860,N_12589);
and U18836 (N_18836,N_10591,N_14286);
or U18837 (N_18837,N_13562,N_13440);
nand U18838 (N_18838,N_11640,N_14467);
and U18839 (N_18839,N_12592,N_12283);
nor U18840 (N_18840,N_10528,N_10146);
nor U18841 (N_18841,N_13831,N_13391);
nor U18842 (N_18842,N_13635,N_14263);
nor U18843 (N_18843,N_13361,N_13063);
nor U18844 (N_18844,N_14102,N_10004);
or U18845 (N_18845,N_10466,N_11678);
or U18846 (N_18846,N_14831,N_12405);
nand U18847 (N_18847,N_10891,N_10680);
nor U18848 (N_18848,N_13666,N_12983);
xor U18849 (N_18849,N_11054,N_10441);
and U18850 (N_18850,N_12451,N_12086);
xor U18851 (N_18851,N_12803,N_10588);
nand U18852 (N_18852,N_12773,N_14210);
nor U18853 (N_18853,N_10440,N_12515);
or U18854 (N_18854,N_10807,N_11244);
or U18855 (N_18855,N_14389,N_11023);
or U18856 (N_18856,N_10121,N_14799);
nand U18857 (N_18857,N_13596,N_11108);
xor U18858 (N_18858,N_11976,N_11037);
nand U18859 (N_18859,N_11295,N_11699);
xnor U18860 (N_18860,N_14801,N_13867);
or U18861 (N_18861,N_11305,N_13130);
nor U18862 (N_18862,N_11803,N_10724);
and U18863 (N_18863,N_10975,N_12924);
xor U18864 (N_18864,N_11588,N_13982);
or U18865 (N_18865,N_11276,N_13400);
nor U18866 (N_18866,N_13216,N_10940);
nand U18867 (N_18867,N_14117,N_11088);
nand U18868 (N_18868,N_13225,N_14571);
nor U18869 (N_18869,N_12287,N_12773);
xnor U18870 (N_18870,N_10115,N_12557);
or U18871 (N_18871,N_12238,N_13612);
or U18872 (N_18872,N_14763,N_14476);
xor U18873 (N_18873,N_12623,N_12894);
nor U18874 (N_18874,N_11867,N_11833);
nand U18875 (N_18875,N_13081,N_14625);
nand U18876 (N_18876,N_12383,N_14255);
and U18877 (N_18877,N_12057,N_10776);
nand U18878 (N_18878,N_11964,N_12447);
xnor U18879 (N_18879,N_12422,N_12371);
xnor U18880 (N_18880,N_14842,N_10347);
or U18881 (N_18881,N_10266,N_13698);
nor U18882 (N_18882,N_11594,N_10775);
xor U18883 (N_18883,N_13030,N_12863);
nor U18884 (N_18884,N_12739,N_10936);
xor U18885 (N_18885,N_12867,N_14883);
nand U18886 (N_18886,N_13414,N_12323);
nor U18887 (N_18887,N_10891,N_13354);
and U18888 (N_18888,N_12067,N_14848);
and U18889 (N_18889,N_13969,N_12281);
nor U18890 (N_18890,N_12167,N_12084);
and U18891 (N_18891,N_11117,N_12557);
nand U18892 (N_18892,N_13921,N_13867);
and U18893 (N_18893,N_13658,N_12218);
nand U18894 (N_18894,N_10581,N_11491);
or U18895 (N_18895,N_11893,N_14352);
or U18896 (N_18896,N_10370,N_13310);
nor U18897 (N_18897,N_10865,N_10657);
nor U18898 (N_18898,N_12160,N_12292);
and U18899 (N_18899,N_13771,N_13783);
or U18900 (N_18900,N_14425,N_10888);
and U18901 (N_18901,N_10635,N_10260);
xnor U18902 (N_18902,N_11377,N_12371);
nand U18903 (N_18903,N_14312,N_11780);
nor U18904 (N_18904,N_14409,N_12170);
nor U18905 (N_18905,N_12246,N_11469);
nor U18906 (N_18906,N_10249,N_14716);
xor U18907 (N_18907,N_14390,N_14658);
nand U18908 (N_18908,N_14210,N_14223);
nand U18909 (N_18909,N_10436,N_12487);
nor U18910 (N_18910,N_13580,N_10983);
or U18911 (N_18911,N_12375,N_11862);
and U18912 (N_18912,N_11941,N_14718);
xnor U18913 (N_18913,N_11236,N_11616);
and U18914 (N_18914,N_14519,N_14524);
nor U18915 (N_18915,N_13515,N_13395);
xnor U18916 (N_18916,N_14338,N_10507);
and U18917 (N_18917,N_12651,N_13264);
nand U18918 (N_18918,N_13106,N_12206);
nor U18919 (N_18919,N_14926,N_10899);
nor U18920 (N_18920,N_12824,N_12003);
nand U18921 (N_18921,N_10388,N_11529);
xor U18922 (N_18922,N_13967,N_12932);
or U18923 (N_18923,N_10763,N_12990);
nor U18924 (N_18924,N_12181,N_12402);
and U18925 (N_18925,N_12809,N_11591);
nand U18926 (N_18926,N_10586,N_10448);
nor U18927 (N_18927,N_12202,N_10168);
nand U18928 (N_18928,N_13501,N_14632);
nor U18929 (N_18929,N_12604,N_10225);
nand U18930 (N_18930,N_10000,N_10138);
or U18931 (N_18931,N_10189,N_10295);
xor U18932 (N_18932,N_11967,N_13779);
and U18933 (N_18933,N_13496,N_14234);
or U18934 (N_18934,N_13163,N_12877);
nand U18935 (N_18935,N_11084,N_13590);
xor U18936 (N_18936,N_11873,N_10015);
and U18937 (N_18937,N_10109,N_10688);
nor U18938 (N_18938,N_12757,N_12503);
nand U18939 (N_18939,N_10231,N_10379);
and U18940 (N_18940,N_12584,N_13556);
and U18941 (N_18941,N_14299,N_13654);
and U18942 (N_18942,N_14476,N_11798);
nand U18943 (N_18943,N_10316,N_14295);
or U18944 (N_18944,N_10577,N_13883);
or U18945 (N_18945,N_14566,N_13034);
or U18946 (N_18946,N_10807,N_13555);
or U18947 (N_18947,N_10875,N_14555);
xor U18948 (N_18948,N_13570,N_10211);
nand U18949 (N_18949,N_13575,N_14444);
or U18950 (N_18950,N_12022,N_12027);
xor U18951 (N_18951,N_13628,N_11548);
and U18952 (N_18952,N_12194,N_14311);
or U18953 (N_18953,N_10131,N_14906);
and U18954 (N_18954,N_13670,N_11765);
nor U18955 (N_18955,N_13575,N_11646);
or U18956 (N_18956,N_14000,N_10958);
xnor U18957 (N_18957,N_11950,N_13057);
nand U18958 (N_18958,N_13339,N_12457);
xor U18959 (N_18959,N_10036,N_14260);
nand U18960 (N_18960,N_11269,N_14452);
nand U18961 (N_18961,N_13255,N_13849);
xnor U18962 (N_18962,N_10524,N_14673);
and U18963 (N_18963,N_14430,N_14453);
or U18964 (N_18964,N_14199,N_12032);
nor U18965 (N_18965,N_10840,N_11000);
nor U18966 (N_18966,N_14524,N_13255);
and U18967 (N_18967,N_13307,N_10768);
nand U18968 (N_18968,N_14687,N_11384);
nor U18969 (N_18969,N_12771,N_12418);
xor U18970 (N_18970,N_13023,N_14749);
nand U18971 (N_18971,N_13355,N_10541);
and U18972 (N_18972,N_13281,N_13059);
or U18973 (N_18973,N_13810,N_13486);
xor U18974 (N_18974,N_14152,N_12540);
nor U18975 (N_18975,N_11706,N_13726);
nor U18976 (N_18976,N_12650,N_12911);
or U18977 (N_18977,N_14753,N_12965);
nand U18978 (N_18978,N_11140,N_14153);
xor U18979 (N_18979,N_11685,N_12648);
and U18980 (N_18980,N_12530,N_12251);
xnor U18981 (N_18981,N_12531,N_12440);
or U18982 (N_18982,N_13679,N_11894);
and U18983 (N_18983,N_11174,N_12241);
nand U18984 (N_18984,N_14033,N_10005);
or U18985 (N_18985,N_12551,N_14403);
and U18986 (N_18986,N_13031,N_11958);
xor U18987 (N_18987,N_14674,N_14522);
or U18988 (N_18988,N_12397,N_11916);
or U18989 (N_18989,N_11970,N_14479);
xnor U18990 (N_18990,N_12410,N_10546);
and U18991 (N_18991,N_12494,N_13292);
xnor U18992 (N_18992,N_14332,N_14738);
or U18993 (N_18993,N_11161,N_10530);
nor U18994 (N_18994,N_10646,N_10900);
and U18995 (N_18995,N_11493,N_12113);
nor U18996 (N_18996,N_11264,N_14758);
and U18997 (N_18997,N_11555,N_14553);
xnor U18998 (N_18998,N_14972,N_13737);
or U18999 (N_18999,N_14622,N_11968);
xor U19000 (N_19000,N_10622,N_13522);
nand U19001 (N_19001,N_13884,N_11980);
and U19002 (N_19002,N_13966,N_10971);
nor U19003 (N_19003,N_13338,N_11915);
xnor U19004 (N_19004,N_14141,N_13038);
xor U19005 (N_19005,N_11200,N_13687);
and U19006 (N_19006,N_13321,N_14081);
or U19007 (N_19007,N_13786,N_11926);
xnor U19008 (N_19008,N_10861,N_13588);
xnor U19009 (N_19009,N_11496,N_13216);
and U19010 (N_19010,N_11446,N_12447);
or U19011 (N_19011,N_10688,N_12124);
and U19012 (N_19012,N_10721,N_11114);
nor U19013 (N_19013,N_12086,N_13362);
xor U19014 (N_19014,N_13066,N_10643);
or U19015 (N_19015,N_12242,N_11993);
nand U19016 (N_19016,N_11964,N_14636);
nand U19017 (N_19017,N_11054,N_11802);
nand U19018 (N_19018,N_14453,N_14196);
nand U19019 (N_19019,N_11673,N_11936);
and U19020 (N_19020,N_10922,N_11429);
nor U19021 (N_19021,N_14414,N_14566);
xnor U19022 (N_19022,N_12533,N_14639);
and U19023 (N_19023,N_13701,N_10685);
or U19024 (N_19024,N_11623,N_10346);
nor U19025 (N_19025,N_11673,N_10569);
and U19026 (N_19026,N_14710,N_10032);
and U19027 (N_19027,N_11978,N_14481);
nor U19028 (N_19028,N_14941,N_12449);
nand U19029 (N_19029,N_13279,N_13494);
or U19030 (N_19030,N_12299,N_13395);
xor U19031 (N_19031,N_10041,N_10406);
or U19032 (N_19032,N_12798,N_13405);
and U19033 (N_19033,N_14784,N_14864);
nand U19034 (N_19034,N_14461,N_13667);
nor U19035 (N_19035,N_12014,N_11931);
nor U19036 (N_19036,N_12639,N_12790);
nand U19037 (N_19037,N_13926,N_11663);
and U19038 (N_19038,N_13545,N_14835);
nor U19039 (N_19039,N_10083,N_13275);
xnor U19040 (N_19040,N_11060,N_14137);
and U19041 (N_19041,N_14551,N_10684);
nand U19042 (N_19042,N_13080,N_11198);
or U19043 (N_19043,N_11969,N_14833);
nand U19044 (N_19044,N_10922,N_13606);
or U19045 (N_19045,N_10919,N_13129);
nand U19046 (N_19046,N_13791,N_11163);
xor U19047 (N_19047,N_13628,N_10744);
nand U19048 (N_19048,N_11482,N_11436);
and U19049 (N_19049,N_13181,N_10563);
and U19050 (N_19050,N_10951,N_12807);
or U19051 (N_19051,N_14632,N_12954);
or U19052 (N_19052,N_13277,N_14766);
nor U19053 (N_19053,N_13214,N_11761);
nand U19054 (N_19054,N_11376,N_11067);
and U19055 (N_19055,N_11659,N_12800);
nor U19056 (N_19056,N_11379,N_13835);
xor U19057 (N_19057,N_13248,N_11369);
nor U19058 (N_19058,N_10823,N_11212);
and U19059 (N_19059,N_10170,N_12115);
or U19060 (N_19060,N_14252,N_14403);
and U19061 (N_19061,N_13600,N_13401);
or U19062 (N_19062,N_11755,N_11033);
nor U19063 (N_19063,N_12578,N_11523);
xor U19064 (N_19064,N_12798,N_12663);
xnor U19065 (N_19065,N_11241,N_10423);
nor U19066 (N_19066,N_12019,N_11942);
and U19067 (N_19067,N_14805,N_11554);
nand U19068 (N_19068,N_14549,N_12863);
xnor U19069 (N_19069,N_12653,N_10379);
and U19070 (N_19070,N_11814,N_14100);
xor U19071 (N_19071,N_10918,N_11689);
or U19072 (N_19072,N_12813,N_10566);
and U19073 (N_19073,N_14916,N_13795);
nor U19074 (N_19074,N_13854,N_11170);
nand U19075 (N_19075,N_12408,N_14060);
or U19076 (N_19076,N_12560,N_11968);
xor U19077 (N_19077,N_10167,N_14917);
or U19078 (N_19078,N_10561,N_10220);
or U19079 (N_19079,N_11352,N_12470);
and U19080 (N_19080,N_10480,N_10652);
nor U19081 (N_19081,N_11735,N_12519);
nor U19082 (N_19082,N_12984,N_14708);
or U19083 (N_19083,N_13207,N_10237);
or U19084 (N_19084,N_10570,N_14470);
nand U19085 (N_19085,N_14729,N_11452);
xnor U19086 (N_19086,N_10317,N_13688);
and U19087 (N_19087,N_13585,N_13565);
and U19088 (N_19088,N_14468,N_12540);
nand U19089 (N_19089,N_10143,N_13602);
or U19090 (N_19090,N_10012,N_10878);
and U19091 (N_19091,N_13966,N_13409);
or U19092 (N_19092,N_11222,N_13664);
or U19093 (N_19093,N_14236,N_12045);
or U19094 (N_19094,N_14185,N_14813);
or U19095 (N_19095,N_12565,N_11778);
xnor U19096 (N_19096,N_10007,N_12012);
nor U19097 (N_19097,N_13399,N_13255);
xnor U19098 (N_19098,N_13600,N_12124);
xor U19099 (N_19099,N_11614,N_13461);
nor U19100 (N_19100,N_12007,N_12526);
nand U19101 (N_19101,N_14640,N_10447);
or U19102 (N_19102,N_13826,N_10112);
nor U19103 (N_19103,N_14529,N_10570);
and U19104 (N_19104,N_14298,N_10284);
nand U19105 (N_19105,N_13242,N_13274);
or U19106 (N_19106,N_10240,N_13728);
nand U19107 (N_19107,N_13401,N_13468);
nor U19108 (N_19108,N_12276,N_14219);
nand U19109 (N_19109,N_14045,N_11715);
and U19110 (N_19110,N_11656,N_13776);
or U19111 (N_19111,N_13431,N_13329);
and U19112 (N_19112,N_10770,N_14227);
nor U19113 (N_19113,N_13440,N_11686);
and U19114 (N_19114,N_12129,N_13359);
xnor U19115 (N_19115,N_14530,N_12587);
nor U19116 (N_19116,N_14779,N_10809);
xnor U19117 (N_19117,N_11939,N_13070);
nor U19118 (N_19118,N_14940,N_14031);
nand U19119 (N_19119,N_12268,N_11542);
nor U19120 (N_19120,N_11660,N_12881);
nor U19121 (N_19121,N_12016,N_14534);
and U19122 (N_19122,N_14053,N_13449);
xor U19123 (N_19123,N_11878,N_12297);
nor U19124 (N_19124,N_12558,N_14763);
and U19125 (N_19125,N_10867,N_12391);
or U19126 (N_19126,N_13033,N_10027);
nor U19127 (N_19127,N_13530,N_14135);
and U19128 (N_19128,N_12384,N_12320);
or U19129 (N_19129,N_12315,N_14980);
or U19130 (N_19130,N_12882,N_14483);
or U19131 (N_19131,N_13556,N_12266);
and U19132 (N_19132,N_11290,N_14764);
or U19133 (N_19133,N_14496,N_11784);
xnor U19134 (N_19134,N_14378,N_14259);
nand U19135 (N_19135,N_11120,N_11093);
nor U19136 (N_19136,N_14996,N_12234);
and U19137 (N_19137,N_11041,N_12348);
nor U19138 (N_19138,N_12841,N_13616);
nor U19139 (N_19139,N_12702,N_10905);
nand U19140 (N_19140,N_10607,N_13576);
and U19141 (N_19141,N_12057,N_11027);
nand U19142 (N_19142,N_12657,N_10122);
nand U19143 (N_19143,N_10815,N_13426);
nand U19144 (N_19144,N_14527,N_14809);
nor U19145 (N_19145,N_11510,N_14605);
nand U19146 (N_19146,N_13387,N_12153);
and U19147 (N_19147,N_12890,N_11862);
xnor U19148 (N_19148,N_12173,N_14198);
and U19149 (N_19149,N_10608,N_14617);
and U19150 (N_19150,N_14786,N_12356);
and U19151 (N_19151,N_14680,N_13159);
xnor U19152 (N_19152,N_12159,N_11116);
or U19153 (N_19153,N_10197,N_13418);
nor U19154 (N_19154,N_10411,N_10389);
nor U19155 (N_19155,N_11462,N_14328);
xor U19156 (N_19156,N_13450,N_10087);
xor U19157 (N_19157,N_14315,N_13363);
xor U19158 (N_19158,N_13287,N_12722);
nand U19159 (N_19159,N_11467,N_12866);
nor U19160 (N_19160,N_12299,N_13038);
and U19161 (N_19161,N_12249,N_10726);
nor U19162 (N_19162,N_11522,N_12103);
or U19163 (N_19163,N_11282,N_10862);
nor U19164 (N_19164,N_12317,N_14667);
nor U19165 (N_19165,N_14083,N_12796);
nor U19166 (N_19166,N_12713,N_12096);
and U19167 (N_19167,N_14117,N_12993);
nor U19168 (N_19168,N_10678,N_12224);
nand U19169 (N_19169,N_10006,N_13379);
xnor U19170 (N_19170,N_13514,N_12047);
nand U19171 (N_19171,N_13738,N_14832);
nor U19172 (N_19172,N_13402,N_11215);
or U19173 (N_19173,N_10901,N_13061);
and U19174 (N_19174,N_10113,N_14831);
and U19175 (N_19175,N_11832,N_10944);
nand U19176 (N_19176,N_10962,N_10336);
or U19177 (N_19177,N_12119,N_13391);
nor U19178 (N_19178,N_11053,N_14640);
xnor U19179 (N_19179,N_14969,N_11519);
xor U19180 (N_19180,N_11563,N_12146);
nand U19181 (N_19181,N_11069,N_11450);
xnor U19182 (N_19182,N_11019,N_10151);
and U19183 (N_19183,N_14982,N_12497);
nand U19184 (N_19184,N_10125,N_14434);
nand U19185 (N_19185,N_13429,N_10163);
nand U19186 (N_19186,N_10317,N_12084);
nor U19187 (N_19187,N_14480,N_12431);
nor U19188 (N_19188,N_14415,N_13656);
xnor U19189 (N_19189,N_11232,N_12174);
xor U19190 (N_19190,N_14472,N_13123);
nor U19191 (N_19191,N_14015,N_10307);
nor U19192 (N_19192,N_11097,N_10961);
or U19193 (N_19193,N_14603,N_13949);
xor U19194 (N_19194,N_10843,N_14702);
nor U19195 (N_19195,N_12049,N_14507);
or U19196 (N_19196,N_12387,N_11501);
and U19197 (N_19197,N_10226,N_13283);
nand U19198 (N_19198,N_11392,N_10363);
and U19199 (N_19199,N_11988,N_13960);
nor U19200 (N_19200,N_13653,N_12931);
nor U19201 (N_19201,N_14542,N_11251);
or U19202 (N_19202,N_14959,N_14310);
xor U19203 (N_19203,N_14734,N_12758);
nand U19204 (N_19204,N_13619,N_11971);
nor U19205 (N_19205,N_12716,N_11463);
or U19206 (N_19206,N_12822,N_14737);
and U19207 (N_19207,N_10088,N_12065);
nand U19208 (N_19208,N_10885,N_12396);
nand U19209 (N_19209,N_13197,N_11693);
or U19210 (N_19210,N_12572,N_13832);
nand U19211 (N_19211,N_13846,N_14530);
nand U19212 (N_19212,N_13612,N_13660);
nand U19213 (N_19213,N_12529,N_10620);
and U19214 (N_19214,N_10494,N_11628);
nor U19215 (N_19215,N_11311,N_13994);
or U19216 (N_19216,N_12292,N_14179);
nor U19217 (N_19217,N_11501,N_11522);
nor U19218 (N_19218,N_10678,N_13141);
and U19219 (N_19219,N_12275,N_14567);
or U19220 (N_19220,N_14673,N_11184);
or U19221 (N_19221,N_14652,N_10962);
nand U19222 (N_19222,N_13899,N_14015);
nand U19223 (N_19223,N_14127,N_12972);
nand U19224 (N_19224,N_10401,N_12987);
xor U19225 (N_19225,N_13431,N_10846);
and U19226 (N_19226,N_12576,N_12501);
nand U19227 (N_19227,N_13927,N_10232);
or U19228 (N_19228,N_12822,N_11504);
nand U19229 (N_19229,N_11838,N_13734);
nor U19230 (N_19230,N_11987,N_12811);
nand U19231 (N_19231,N_12708,N_11418);
and U19232 (N_19232,N_11594,N_10078);
nand U19233 (N_19233,N_11384,N_13998);
or U19234 (N_19234,N_11612,N_12268);
and U19235 (N_19235,N_12407,N_11164);
and U19236 (N_19236,N_13547,N_14614);
or U19237 (N_19237,N_14868,N_12852);
or U19238 (N_19238,N_11452,N_13159);
and U19239 (N_19239,N_10849,N_10730);
and U19240 (N_19240,N_10080,N_11136);
nand U19241 (N_19241,N_14472,N_10672);
nor U19242 (N_19242,N_10434,N_14888);
xnor U19243 (N_19243,N_13993,N_10873);
xnor U19244 (N_19244,N_12442,N_12169);
nand U19245 (N_19245,N_14953,N_14911);
nor U19246 (N_19246,N_14036,N_14402);
xnor U19247 (N_19247,N_11799,N_14877);
and U19248 (N_19248,N_11699,N_12059);
or U19249 (N_19249,N_13351,N_11874);
nor U19250 (N_19250,N_11224,N_11943);
and U19251 (N_19251,N_14916,N_11223);
or U19252 (N_19252,N_13191,N_12398);
xnor U19253 (N_19253,N_11674,N_14715);
and U19254 (N_19254,N_14311,N_11835);
nor U19255 (N_19255,N_12779,N_11295);
xor U19256 (N_19256,N_14068,N_13577);
and U19257 (N_19257,N_10720,N_13602);
nor U19258 (N_19258,N_10813,N_11545);
xor U19259 (N_19259,N_12824,N_12012);
xnor U19260 (N_19260,N_12692,N_14512);
nand U19261 (N_19261,N_11118,N_13710);
xor U19262 (N_19262,N_13366,N_14151);
and U19263 (N_19263,N_11718,N_13838);
nor U19264 (N_19264,N_13389,N_11406);
nand U19265 (N_19265,N_12166,N_13295);
nand U19266 (N_19266,N_14630,N_12449);
nand U19267 (N_19267,N_12027,N_14505);
xor U19268 (N_19268,N_12921,N_13062);
nand U19269 (N_19269,N_10752,N_13905);
nand U19270 (N_19270,N_14087,N_11276);
nor U19271 (N_19271,N_11711,N_13146);
nand U19272 (N_19272,N_12868,N_10358);
xor U19273 (N_19273,N_14923,N_13845);
xnor U19274 (N_19274,N_13815,N_13892);
nor U19275 (N_19275,N_12584,N_10912);
nor U19276 (N_19276,N_11134,N_14680);
and U19277 (N_19277,N_10863,N_12008);
or U19278 (N_19278,N_14403,N_12073);
and U19279 (N_19279,N_14989,N_14495);
nor U19280 (N_19280,N_14039,N_12354);
xor U19281 (N_19281,N_13922,N_12439);
nand U19282 (N_19282,N_10006,N_14778);
nor U19283 (N_19283,N_12667,N_10514);
and U19284 (N_19284,N_11688,N_14878);
xnor U19285 (N_19285,N_13623,N_11585);
xnor U19286 (N_19286,N_12242,N_11014);
nor U19287 (N_19287,N_12723,N_12133);
nor U19288 (N_19288,N_12306,N_13767);
xor U19289 (N_19289,N_10201,N_10314);
nor U19290 (N_19290,N_14141,N_11896);
xnor U19291 (N_19291,N_10849,N_13868);
nand U19292 (N_19292,N_14456,N_13752);
and U19293 (N_19293,N_11003,N_10229);
and U19294 (N_19294,N_12035,N_13258);
and U19295 (N_19295,N_14529,N_10520);
xor U19296 (N_19296,N_14252,N_13624);
or U19297 (N_19297,N_11741,N_10056);
and U19298 (N_19298,N_11742,N_11514);
or U19299 (N_19299,N_13564,N_10698);
nor U19300 (N_19300,N_13913,N_12803);
or U19301 (N_19301,N_10690,N_12470);
xor U19302 (N_19302,N_10875,N_14093);
or U19303 (N_19303,N_13970,N_13411);
nand U19304 (N_19304,N_14466,N_13655);
or U19305 (N_19305,N_13172,N_14194);
nor U19306 (N_19306,N_13216,N_13162);
and U19307 (N_19307,N_10092,N_14351);
xor U19308 (N_19308,N_14467,N_13129);
or U19309 (N_19309,N_12087,N_12775);
xor U19310 (N_19310,N_12917,N_13590);
or U19311 (N_19311,N_11204,N_12411);
nand U19312 (N_19312,N_12104,N_12714);
nor U19313 (N_19313,N_12021,N_10095);
and U19314 (N_19314,N_13223,N_13913);
nand U19315 (N_19315,N_11353,N_12249);
and U19316 (N_19316,N_10349,N_11015);
and U19317 (N_19317,N_10092,N_10205);
or U19318 (N_19318,N_14961,N_10669);
nand U19319 (N_19319,N_11555,N_10026);
and U19320 (N_19320,N_14730,N_10708);
nand U19321 (N_19321,N_14588,N_10553);
and U19322 (N_19322,N_12173,N_12505);
nor U19323 (N_19323,N_12596,N_14367);
and U19324 (N_19324,N_10177,N_11498);
or U19325 (N_19325,N_13170,N_11574);
xor U19326 (N_19326,N_13826,N_10071);
nor U19327 (N_19327,N_13396,N_12042);
nand U19328 (N_19328,N_10525,N_14266);
nor U19329 (N_19329,N_11118,N_10414);
xnor U19330 (N_19330,N_12011,N_13383);
or U19331 (N_19331,N_12318,N_10332);
xnor U19332 (N_19332,N_12540,N_14657);
nor U19333 (N_19333,N_11994,N_14971);
or U19334 (N_19334,N_11808,N_12523);
xor U19335 (N_19335,N_14973,N_14923);
and U19336 (N_19336,N_14984,N_13553);
xnor U19337 (N_19337,N_14619,N_13340);
or U19338 (N_19338,N_13705,N_14830);
nor U19339 (N_19339,N_13280,N_11722);
and U19340 (N_19340,N_12472,N_14061);
xor U19341 (N_19341,N_10146,N_14002);
nor U19342 (N_19342,N_11887,N_14775);
xnor U19343 (N_19343,N_11924,N_10678);
or U19344 (N_19344,N_10764,N_12320);
nor U19345 (N_19345,N_14658,N_14866);
nor U19346 (N_19346,N_12028,N_13420);
or U19347 (N_19347,N_11487,N_10922);
and U19348 (N_19348,N_10058,N_10939);
nor U19349 (N_19349,N_12586,N_10650);
nand U19350 (N_19350,N_12406,N_11770);
nor U19351 (N_19351,N_14272,N_10941);
nand U19352 (N_19352,N_12792,N_13685);
and U19353 (N_19353,N_12146,N_12686);
nor U19354 (N_19354,N_10263,N_11456);
xor U19355 (N_19355,N_11199,N_11931);
xnor U19356 (N_19356,N_13258,N_13251);
xor U19357 (N_19357,N_13517,N_13817);
nand U19358 (N_19358,N_12968,N_13590);
nand U19359 (N_19359,N_14229,N_13691);
or U19360 (N_19360,N_12448,N_10376);
or U19361 (N_19361,N_14846,N_10965);
xor U19362 (N_19362,N_12609,N_10569);
xnor U19363 (N_19363,N_10137,N_12134);
nor U19364 (N_19364,N_12027,N_13960);
nor U19365 (N_19365,N_10555,N_12091);
or U19366 (N_19366,N_14518,N_11042);
nor U19367 (N_19367,N_11455,N_12368);
or U19368 (N_19368,N_14121,N_13923);
nor U19369 (N_19369,N_11140,N_13360);
nand U19370 (N_19370,N_12180,N_10947);
or U19371 (N_19371,N_10565,N_12895);
or U19372 (N_19372,N_13995,N_12391);
xnor U19373 (N_19373,N_12146,N_13750);
or U19374 (N_19374,N_11221,N_13318);
nor U19375 (N_19375,N_13427,N_13458);
or U19376 (N_19376,N_10747,N_12341);
nor U19377 (N_19377,N_13775,N_10216);
xnor U19378 (N_19378,N_12326,N_12242);
and U19379 (N_19379,N_14383,N_11940);
and U19380 (N_19380,N_13938,N_12983);
xor U19381 (N_19381,N_14779,N_13940);
or U19382 (N_19382,N_10832,N_11894);
and U19383 (N_19383,N_11034,N_11975);
xor U19384 (N_19384,N_10634,N_13199);
nand U19385 (N_19385,N_14778,N_14893);
nand U19386 (N_19386,N_13684,N_14157);
nor U19387 (N_19387,N_13193,N_13278);
xnor U19388 (N_19388,N_10837,N_10672);
nand U19389 (N_19389,N_11727,N_10459);
xor U19390 (N_19390,N_12021,N_14911);
nand U19391 (N_19391,N_13890,N_11715);
nor U19392 (N_19392,N_14894,N_12738);
nor U19393 (N_19393,N_10301,N_13599);
and U19394 (N_19394,N_13924,N_11042);
or U19395 (N_19395,N_10368,N_14406);
nor U19396 (N_19396,N_10455,N_10677);
xor U19397 (N_19397,N_14214,N_12767);
or U19398 (N_19398,N_13829,N_12179);
xor U19399 (N_19399,N_14737,N_14837);
and U19400 (N_19400,N_12175,N_13446);
and U19401 (N_19401,N_12895,N_14676);
nand U19402 (N_19402,N_14391,N_13129);
xnor U19403 (N_19403,N_11707,N_12955);
or U19404 (N_19404,N_10299,N_14049);
nor U19405 (N_19405,N_10403,N_14125);
or U19406 (N_19406,N_11194,N_13550);
and U19407 (N_19407,N_13999,N_13809);
or U19408 (N_19408,N_13412,N_12112);
nand U19409 (N_19409,N_14272,N_10939);
and U19410 (N_19410,N_13978,N_13701);
or U19411 (N_19411,N_10545,N_13129);
and U19412 (N_19412,N_11426,N_14010);
and U19413 (N_19413,N_14849,N_11672);
xnor U19414 (N_19414,N_10203,N_14212);
nor U19415 (N_19415,N_14204,N_13034);
or U19416 (N_19416,N_13022,N_12975);
xnor U19417 (N_19417,N_11850,N_13010);
or U19418 (N_19418,N_13209,N_12565);
nor U19419 (N_19419,N_11926,N_10887);
or U19420 (N_19420,N_14879,N_10610);
and U19421 (N_19421,N_10678,N_13012);
nor U19422 (N_19422,N_14478,N_10158);
or U19423 (N_19423,N_13063,N_11366);
xor U19424 (N_19424,N_12381,N_12298);
xor U19425 (N_19425,N_10998,N_12948);
nand U19426 (N_19426,N_11180,N_14755);
nor U19427 (N_19427,N_11334,N_11923);
or U19428 (N_19428,N_11886,N_13785);
nor U19429 (N_19429,N_13784,N_13890);
nor U19430 (N_19430,N_12191,N_11481);
nand U19431 (N_19431,N_14518,N_13730);
or U19432 (N_19432,N_10609,N_13502);
or U19433 (N_19433,N_14347,N_14105);
and U19434 (N_19434,N_13898,N_11069);
or U19435 (N_19435,N_13810,N_12702);
xor U19436 (N_19436,N_14750,N_12136);
nor U19437 (N_19437,N_13106,N_14928);
nand U19438 (N_19438,N_12064,N_10847);
and U19439 (N_19439,N_14374,N_12648);
xor U19440 (N_19440,N_11351,N_12728);
and U19441 (N_19441,N_12567,N_13919);
nor U19442 (N_19442,N_10091,N_12539);
or U19443 (N_19443,N_11355,N_11834);
nand U19444 (N_19444,N_10174,N_14889);
and U19445 (N_19445,N_14212,N_11321);
or U19446 (N_19446,N_13772,N_11895);
xnor U19447 (N_19447,N_12930,N_14113);
xor U19448 (N_19448,N_11735,N_10389);
and U19449 (N_19449,N_13458,N_13068);
or U19450 (N_19450,N_11137,N_12693);
or U19451 (N_19451,N_11796,N_13142);
nor U19452 (N_19452,N_12692,N_11474);
nand U19453 (N_19453,N_14844,N_14672);
or U19454 (N_19454,N_10404,N_12892);
and U19455 (N_19455,N_11597,N_12619);
or U19456 (N_19456,N_11817,N_10473);
or U19457 (N_19457,N_13974,N_12614);
or U19458 (N_19458,N_12899,N_12504);
and U19459 (N_19459,N_14716,N_14826);
or U19460 (N_19460,N_10849,N_14210);
and U19461 (N_19461,N_11724,N_14597);
nor U19462 (N_19462,N_12353,N_11030);
nand U19463 (N_19463,N_13014,N_13704);
xnor U19464 (N_19464,N_10445,N_12100);
nand U19465 (N_19465,N_14222,N_13339);
or U19466 (N_19466,N_13733,N_12737);
xnor U19467 (N_19467,N_11514,N_12040);
nand U19468 (N_19468,N_14187,N_12021);
nand U19469 (N_19469,N_13927,N_14674);
nor U19470 (N_19470,N_11061,N_14418);
xnor U19471 (N_19471,N_14957,N_13727);
xor U19472 (N_19472,N_14191,N_10969);
xnor U19473 (N_19473,N_13026,N_12295);
or U19474 (N_19474,N_14924,N_13763);
and U19475 (N_19475,N_14815,N_10957);
or U19476 (N_19476,N_11287,N_13598);
or U19477 (N_19477,N_12939,N_12165);
nand U19478 (N_19478,N_10932,N_13899);
or U19479 (N_19479,N_12653,N_13572);
or U19480 (N_19480,N_13272,N_11712);
and U19481 (N_19481,N_14860,N_14784);
nand U19482 (N_19482,N_12057,N_14342);
xor U19483 (N_19483,N_10376,N_10315);
xnor U19484 (N_19484,N_13386,N_14865);
xnor U19485 (N_19485,N_11054,N_13127);
nand U19486 (N_19486,N_10405,N_12289);
nor U19487 (N_19487,N_12798,N_13522);
and U19488 (N_19488,N_13945,N_10451);
and U19489 (N_19489,N_13621,N_13628);
nor U19490 (N_19490,N_13701,N_13853);
nor U19491 (N_19491,N_11793,N_14814);
or U19492 (N_19492,N_14228,N_12916);
nor U19493 (N_19493,N_11591,N_14436);
or U19494 (N_19494,N_12281,N_13426);
or U19495 (N_19495,N_13907,N_12710);
xor U19496 (N_19496,N_13826,N_13540);
nor U19497 (N_19497,N_14860,N_11950);
xnor U19498 (N_19498,N_12699,N_10486);
xnor U19499 (N_19499,N_10451,N_13921);
or U19500 (N_19500,N_12576,N_11724);
and U19501 (N_19501,N_13162,N_10181);
or U19502 (N_19502,N_12058,N_14539);
nand U19503 (N_19503,N_12937,N_12121);
xor U19504 (N_19504,N_11268,N_11932);
or U19505 (N_19505,N_14159,N_11203);
xnor U19506 (N_19506,N_14122,N_14130);
xnor U19507 (N_19507,N_10990,N_11339);
or U19508 (N_19508,N_12664,N_13822);
xor U19509 (N_19509,N_10694,N_14801);
xnor U19510 (N_19510,N_11539,N_11995);
xor U19511 (N_19511,N_11515,N_14285);
and U19512 (N_19512,N_11089,N_13860);
nor U19513 (N_19513,N_12981,N_13790);
xor U19514 (N_19514,N_14355,N_13971);
and U19515 (N_19515,N_14580,N_10538);
and U19516 (N_19516,N_11062,N_12145);
xor U19517 (N_19517,N_10227,N_10289);
nand U19518 (N_19518,N_10291,N_14446);
or U19519 (N_19519,N_14538,N_12131);
or U19520 (N_19520,N_10377,N_11348);
nor U19521 (N_19521,N_12309,N_14969);
nor U19522 (N_19522,N_13126,N_13865);
or U19523 (N_19523,N_12339,N_14754);
or U19524 (N_19524,N_14091,N_12545);
and U19525 (N_19525,N_13311,N_13847);
nand U19526 (N_19526,N_10010,N_11300);
nor U19527 (N_19527,N_11450,N_11183);
xnor U19528 (N_19528,N_11609,N_14938);
nor U19529 (N_19529,N_11894,N_14207);
nand U19530 (N_19530,N_14510,N_12248);
and U19531 (N_19531,N_11318,N_10847);
and U19532 (N_19532,N_10294,N_11425);
and U19533 (N_19533,N_12096,N_13642);
or U19534 (N_19534,N_13575,N_13603);
nand U19535 (N_19535,N_14280,N_14355);
nand U19536 (N_19536,N_10238,N_12998);
and U19537 (N_19537,N_13132,N_14363);
nand U19538 (N_19538,N_10686,N_12519);
xor U19539 (N_19539,N_13754,N_13704);
nor U19540 (N_19540,N_11588,N_10857);
and U19541 (N_19541,N_13375,N_11391);
nor U19542 (N_19542,N_10060,N_10824);
nand U19543 (N_19543,N_14917,N_12863);
nand U19544 (N_19544,N_13964,N_13403);
nand U19545 (N_19545,N_14818,N_12668);
and U19546 (N_19546,N_14108,N_11652);
nand U19547 (N_19547,N_13186,N_10691);
xnor U19548 (N_19548,N_10468,N_10623);
nor U19549 (N_19549,N_14283,N_10564);
or U19550 (N_19550,N_13636,N_13282);
xor U19551 (N_19551,N_10978,N_14560);
and U19552 (N_19552,N_14431,N_10867);
nand U19553 (N_19553,N_11714,N_13793);
and U19554 (N_19554,N_11491,N_10343);
nand U19555 (N_19555,N_11867,N_10904);
nand U19556 (N_19556,N_13062,N_13056);
or U19557 (N_19557,N_11536,N_10750);
nand U19558 (N_19558,N_13442,N_10996);
xor U19559 (N_19559,N_12745,N_11746);
xor U19560 (N_19560,N_14957,N_13298);
nand U19561 (N_19561,N_13449,N_14487);
or U19562 (N_19562,N_11606,N_11113);
xnor U19563 (N_19563,N_11648,N_10500);
and U19564 (N_19564,N_14356,N_13858);
nor U19565 (N_19565,N_13949,N_12143);
nand U19566 (N_19566,N_10524,N_13657);
nand U19567 (N_19567,N_12608,N_11443);
nand U19568 (N_19568,N_10214,N_14300);
and U19569 (N_19569,N_14714,N_12091);
and U19570 (N_19570,N_13327,N_13650);
xnor U19571 (N_19571,N_12106,N_14535);
nand U19572 (N_19572,N_12420,N_11080);
and U19573 (N_19573,N_11499,N_11492);
nand U19574 (N_19574,N_12151,N_10396);
and U19575 (N_19575,N_10389,N_10579);
nor U19576 (N_19576,N_10900,N_14677);
nor U19577 (N_19577,N_11156,N_12732);
nor U19578 (N_19578,N_11371,N_14391);
xor U19579 (N_19579,N_11088,N_14397);
or U19580 (N_19580,N_10794,N_13482);
or U19581 (N_19581,N_13458,N_14232);
nand U19582 (N_19582,N_14221,N_12712);
nor U19583 (N_19583,N_11201,N_12698);
and U19584 (N_19584,N_13006,N_13837);
nor U19585 (N_19585,N_14237,N_12964);
or U19586 (N_19586,N_12882,N_14749);
nand U19587 (N_19587,N_11519,N_10064);
and U19588 (N_19588,N_13340,N_13148);
and U19589 (N_19589,N_12899,N_13193);
xnor U19590 (N_19590,N_14833,N_14899);
or U19591 (N_19591,N_14246,N_14242);
or U19592 (N_19592,N_11580,N_14582);
xor U19593 (N_19593,N_10752,N_12933);
nand U19594 (N_19594,N_11751,N_14183);
nor U19595 (N_19595,N_11891,N_13352);
xor U19596 (N_19596,N_12908,N_14438);
nand U19597 (N_19597,N_14594,N_14085);
xnor U19598 (N_19598,N_13081,N_12451);
and U19599 (N_19599,N_11543,N_11111);
xnor U19600 (N_19600,N_14606,N_12498);
xor U19601 (N_19601,N_14332,N_14223);
and U19602 (N_19602,N_11504,N_12726);
xnor U19603 (N_19603,N_13453,N_12100);
and U19604 (N_19604,N_12791,N_10427);
nor U19605 (N_19605,N_12512,N_11313);
xor U19606 (N_19606,N_11697,N_13514);
and U19607 (N_19607,N_14971,N_13924);
or U19608 (N_19608,N_11686,N_14369);
and U19609 (N_19609,N_14855,N_14077);
nor U19610 (N_19610,N_14887,N_12935);
nand U19611 (N_19611,N_12131,N_11875);
and U19612 (N_19612,N_14670,N_11406);
or U19613 (N_19613,N_12955,N_13355);
nor U19614 (N_19614,N_13183,N_11112);
and U19615 (N_19615,N_14791,N_12690);
or U19616 (N_19616,N_14911,N_11357);
nor U19617 (N_19617,N_14783,N_11088);
nand U19618 (N_19618,N_11482,N_14242);
nand U19619 (N_19619,N_13516,N_11910);
xor U19620 (N_19620,N_13650,N_12279);
nor U19621 (N_19621,N_12049,N_11158);
xor U19622 (N_19622,N_10064,N_12538);
nor U19623 (N_19623,N_12795,N_12824);
or U19624 (N_19624,N_10874,N_13199);
and U19625 (N_19625,N_10559,N_13636);
or U19626 (N_19626,N_11155,N_13268);
and U19627 (N_19627,N_14404,N_11000);
and U19628 (N_19628,N_12704,N_11627);
nor U19629 (N_19629,N_11335,N_14898);
nor U19630 (N_19630,N_12137,N_13210);
nand U19631 (N_19631,N_10784,N_10207);
nand U19632 (N_19632,N_13440,N_14703);
or U19633 (N_19633,N_13603,N_13591);
and U19634 (N_19634,N_12679,N_14718);
and U19635 (N_19635,N_11462,N_11960);
nand U19636 (N_19636,N_14891,N_11125);
nor U19637 (N_19637,N_12678,N_12174);
nor U19638 (N_19638,N_11297,N_11478);
and U19639 (N_19639,N_12335,N_14071);
nand U19640 (N_19640,N_13041,N_14648);
and U19641 (N_19641,N_10908,N_14411);
or U19642 (N_19642,N_12530,N_12023);
nor U19643 (N_19643,N_12641,N_11083);
nand U19644 (N_19644,N_10551,N_11962);
nor U19645 (N_19645,N_12600,N_13301);
nand U19646 (N_19646,N_11496,N_13666);
or U19647 (N_19647,N_12706,N_11965);
or U19648 (N_19648,N_12011,N_10882);
xor U19649 (N_19649,N_14662,N_12112);
nor U19650 (N_19650,N_10446,N_13682);
or U19651 (N_19651,N_10962,N_10631);
xor U19652 (N_19652,N_11654,N_12933);
xor U19653 (N_19653,N_13329,N_12725);
nor U19654 (N_19654,N_14990,N_10919);
nor U19655 (N_19655,N_12781,N_13287);
or U19656 (N_19656,N_13147,N_11632);
or U19657 (N_19657,N_14928,N_13170);
nand U19658 (N_19658,N_10523,N_12811);
xnor U19659 (N_19659,N_11927,N_12679);
nand U19660 (N_19660,N_12208,N_13884);
and U19661 (N_19661,N_12027,N_10220);
xor U19662 (N_19662,N_11739,N_10341);
or U19663 (N_19663,N_10901,N_14717);
and U19664 (N_19664,N_13421,N_10270);
and U19665 (N_19665,N_10029,N_11921);
xor U19666 (N_19666,N_10933,N_10895);
nor U19667 (N_19667,N_10739,N_12337);
nand U19668 (N_19668,N_12434,N_11705);
xnor U19669 (N_19669,N_10066,N_14812);
nand U19670 (N_19670,N_11914,N_14957);
and U19671 (N_19671,N_10634,N_11372);
xor U19672 (N_19672,N_12352,N_14951);
nor U19673 (N_19673,N_13868,N_14551);
and U19674 (N_19674,N_14667,N_10742);
nor U19675 (N_19675,N_13460,N_12570);
and U19676 (N_19676,N_10708,N_10556);
xor U19677 (N_19677,N_13023,N_10995);
or U19678 (N_19678,N_13743,N_14717);
nor U19679 (N_19679,N_13776,N_12624);
and U19680 (N_19680,N_11608,N_12408);
or U19681 (N_19681,N_13804,N_13708);
nor U19682 (N_19682,N_12293,N_13308);
nor U19683 (N_19683,N_13105,N_10498);
or U19684 (N_19684,N_10966,N_11120);
xor U19685 (N_19685,N_12486,N_11010);
and U19686 (N_19686,N_12417,N_13705);
or U19687 (N_19687,N_10898,N_12025);
or U19688 (N_19688,N_13118,N_11289);
and U19689 (N_19689,N_14707,N_12747);
xnor U19690 (N_19690,N_14698,N_13690);
xnor U19691 (N_19691,N_12422,N_13432);
and U19692 (N_19692,N_12137,N_11035);
nand U19693 (N_19693,N_14290,N_10990);
and U19694 (N_19694,N_13049,N_12583);
or U19695 (N_19695,N_11799,N_14309);
nand U19696 (N_19696,N_10718,N_12109);
nor U19697 (N_19697,N_12304,N_10333);
nand U19698 (N_19698,N_11912,N_13357);
and U19699 (N_19699,N_11126,N_10188);
nor U19700 (N_19700,N_14842,N_12753);
nor U19701 (N_19701,N_13048,N_10791);
nand U19702 (N_19702,N_13028,N_10519);
and U19703 (N_19703,N_10501,N_12163);
nor U19704 (N_19704,N_11014,N_11017);
nor U19705 (N_19705,N_11683,N_14464);
xor U19706 (N_19706,N_12371,N_12442);
nor U19707 (N_19707,N_10816,N_12877);
nand U19708 (N_19708,N_14684,N_10879);
xnor U19709 (N_19709,N_10686,N_14137);
nor U19710 (N_19710,N_13743,N_10955);
nand U19711 (N_19711,N_12537,N_10850);
nor U19712 (N_19712,N_14083,N_14984);
or U19713 (N_19713,N_11249,N_12515);
nand U19714 (N_19714,N_10316,N_14005);
or U19715 (N_19715,N_12295,N_12039);
and U19716 (N_19716,N_11224,N_10462);
nand U19717 (N_19717,N_14101,N_11789);
nand U19718 (N_19718,N_14313,N_14543);
nor U19719 (N_19719,N_14681,N_13130);
nand U19720 (N_19720,N_13867,N_12156);
nand U19721 (N_19721,N_10348,N_13478);
nor U19722 (N_19722,N_11502,N_14407);
nand U19723 (N_19723,N_14597,N_11128);
nand U19724 (N_19724,N_11222,N_12680);
and U19725 (N_19725,N_11568,N_10752);
or U19726 (N_19726,N_13836,N_12213);
nor U19727 (N_19727,N_10810,N_14782);
nor U19728 (N_19728,N_11547,N_11435);
xor U19729 (N_19729,N_12995,N_10469);
nand U19730 (N_19730,N_10242,N_12587);
nand U19731 (N_19731,N_13631,N_10342);
nor U19732 (N_19732,N_14894,N_11352);
nor U19733 (N_19733,N_10737,N_13854);
xnor U19734 (N_19734,N_13651,N_11150);
nand U19735 (N_19735,N_12917,N_14983);
nor U19736 (N_19736,N_10213,N_13963);
or U19737 (N_19737,N_11023,N_10074);
xor U19738 (N_19738,N_12991,N_11215);
nor U19739 (N_19739,N_10339,N_12139);
xnor U19740 (N_19740,N_12409,N_10789);
and U19741 (N_19741,N_12890,N_12173);
nor U19742 (N_19742,N_10112,N_13475);
or U19743 (N_19743,N_12787,N_12695);
and U19744 (N_19744,N_10102,N_11832);
or U19745 (N_19745,N_10735,N_11422);
and U19746 (N_19746,N_13790,N_11881);
and U19747 (N_19747,N_14671,N_11003);
xor U19748 (N_19748,N_10597,N_13415);
and U19749 (N_19749,N_13949,N_12275);
and U19750 (N_19750,N_13125,N_11846);
or U19751 (N_19751,N_10861,N_13531);
nand U19752 (N_19752,N_11880,N_14963);
xnor U19753 (N_19753,N_10240,N_13070);
or U19754 (N_19754,N_11104,N_13367);
nand U19755 (N_19755,N_11272,N_12635);
nor U19756 (N_19756,N_12831,N_13174);
nor U19757 (N_19757,N_12162,N_13687);
nor U19758 (N_19758,N_11166,N_11830);
nor U19759 (N_19759,N_11039,N_14771);
nor U19760 (N_19760,N_10309,N_11371);
and U19761 (N_19761,N_10876,N_11508);
and U19762 (N_19762,N_10236,N_11959);
and U19763 (N_19763,N_14868,N_10769);
xnor U19764 (N_19764,N_13576,N_11523);
xor U19765 (N_19765,N_10704,N_12737);
or U19766 (N_19766,N_10304,N_10115);
and U19767 (N_19767,N_13541,N_10450);
and U19768 (N_19768,N_12682,N_12080);
nand U19769 (N_19769,N_11995,N_14167);
nor U19770 (N_19770,N_10936,N_14974);
and U19771 (N_19771,N_12974,N_10685);
or U19772 (N_19772,N_12719,N_12633);
and U19773 (N_19773,N_12860,N_11536);
nor U19774 (N_19774,N_13199,N_12667);
xnor U19775 (N_19775,N_11818,N_12612);
nand U19776 (N_19776,N_10545,N_12694);
nand U19777 (N_19777,N_12642,N_11055);
xor U19778 (N_19778,N_13858,N_13345);
and U19779 (N_19779,N_13337,N_10320);
xnor U19780 (N_19780,N_11305,N_14402);
nor U19781 (N_19781,N_14018,N_11739);
or U19782 (N_19782,N_12407,N_12745);
nand U19783 (N_19783,N_14048,N_12864);
nor U19784 (N_19784,N_10150,N_11659);
nor U19785 (N_19785,N_13658,N_10054);
nor U19786 (N_19786,N_10568,N_11285);
nor U19787 (N_19787,N_13887,N_10464);
or U19788 (N_19788,N_12298,N_10805);
and U19789 (N_19789,N_11659,N_10333);
nor U19790 (N_19790,N_13712,N_11624);
nor U19791 (N_19791,N_11281,N_14385);
or U19792 (N_19792,N_14268,N_12125);
nor U19793 (N_19793,N_10864,N_11249);
nand U19794 (N_19794,N_14501,N_10201);
and U19795 (N_19795,N_13857,N_13220);
xnor U19796 (N_19796,N_13593,N_13097);
xor U19797 (N_19797,N_11156,N_13343);
xor U19798 (N_19798,N_12273,N_14011);
nand U19799 (N_19799,N_10418,N_14404);
nand U19800 (N_19800,N_11915,N_14248);
xnor U19801 (N_19801,N_11560,N_13509);
and U19802 (N_19802,N_14001,N_12654);
nand U19803 (N_19803,N_13967,N_11347);
xnor U19804 (N_19804,N_11192,N_10948);
or U19805 (N_19805,N_13679,N_10529);
and U19806 (N_19806,N_10415,N_12659);
or U19807 (N_19807,N_11250,N_11766);
and U19808 (N_19808,N_13738,N_14765);
nand U19809 (N_19809,N_13033,N_13024);
nor U19810 (N_19810,N_11885,N_14887);
nor U19811 (N_19811,N_11053,N_14794);
xnor U19812 (N_19812,N_11487,N_11113);
and U19813 (N_19813,N_13259,N_10815);
nor U19814 (N_19814,N_13178,N_10512);
nor U19815 (N_19815,N_11407,N_11330);
or U19816 (N_19816,N_14307,N_13459);
nand U19817 (N_19817,N_10297,N_14727);
xnor U19818 (N_19818,N_11443,N_14995);
nor U19819 (N_19819,N_13500,N_11835);
nand U19820 (N_19820,N_14411,N_12172);
or U19821 (N_19821,N_14271,N_13382);
nor U19822 (N_19822,N_14007,N_14073);
xnor U19823 (N_19823,N_10382,N_11442);
nor U19824 (N_19824,N_14089,N_13227);
or U19825 (N_19825,N_14559,N_12766);
nor U19826 (N_19826,N_11277,N_12730);
nand U19827 (N_19827,N_13325,N_11291);
and U19828 (N_19828,N_11883,N_14712);
and U19829 (N_19829,N_11690,N_13047);
and U19830 (N_19830,N_13200,N_10592);
nand U19831 (N_19831,N_14547,N_10392);
or U19832 (N_19832,N_12014,N_12464);
and U19833 (N_19833,N_13969,N_10382);
xor U19834 (N_19834,N_10294,N_13537);
nand U19835 (N_19835,N_10198,N_11675);
nand U19836 (N_19836,N_13383,N_13133);
and U19837 (N_19837,N_11762,N_10664);
nor U19838 (N_19838,N_14972,N_10492);
or U19839 (N_19839,N_11465,N_11652);
nor U19840 (N_19840,N_12711,N_13478);
or U19841 (N_19841,N_13650,N_10363);
nand U19842 (N_19842,N_11372,N_12156);
nand U19843 (N_19843,N_12929,N_13707);
nor U19844 (N_19844,N_14938,N_11474);
or U19845 (N_19845,N_13488,N_12052);
and U19846 (N_19846,N_11351,N_10892);
nor U19847 (N_19847,N_10743,N_10873);
xor U19848 (N_19848,N_12398,N_12168);
nor U19849 (N_19849,N_10445,N_12168);
nand U19850 (N_19850,N_10750,N_10919);
nor U19851 (N_19851,N_12907,N_11703);
or U19852 (N_19852,N_10286,N_11474);
and U19853 (N_19853,N_12739,N_12536);
nand U19854 (N_19854,N_14158,N_10421);
and U19855 (N_19855,N_14916,N_10901);
nor U19856 (N_19856,N_14663,N_13784);
and U19857 (N_19857,N_12566,N_11438);
nand U19858 (N_19858,N_13119,N_13198);
or U19859 (N_19859,N_10219,N_14380);
nand U19860 (N_19860,N_11531,N_12657);
and U19861 (N_19861,N_10998,N_10498);
xnor U19862 (N_19862,N_10420,N_10402);
or U19863 (N_19863,N_12211,N_13100);
and U19864 (N_19864,N_13841,N_12575);
nand U19865 (N_19865,N_10910,N_13499);
nor U19866 (N_19866,N_13480,N_12413);
and U19867 (N_19867,N_11020,N_14735);
nor U19868 (N_19868,N_14730,N_13756);
or U19869 (N_19869,N_13568,N_11922);
or U19870 (N_19870,N_11121,N_14291);
nand U19871 (N_19871,N_14807,N_13059);
xnor U19872 (N_19872,N_14482,N_10965);
nand U19873 (N_19873,N_11143,N_11834);
and U19874 (N_19874,N_12580,N_13031);
xnor U19875 (N_19875,N_10258,N_12719);
nor U19876 (N_19876,N_14606,N_10414);
or U19877 (N_19877,N_14696,N_11265);
xnor U19878 (N_19878,N_10350,N_14339);
xor U19879 (N_19879,N_10688,N_14852);
and U19880 (N_19880,N_11640,N_12639);
nand U19881 (N_19881,N_10432,N_14534);
nor U19882 (N_19882,N_13090,N_11770);
xnor U19883 (N_19883,N_14884,N_14634);
xnor U19884 (N_19884,N_11166,N_12282);
nand U19885 (N_19885,N_10522,N_14035);
nand U19886 (N_19886,N_13362,N_12051);
xor U19887 (N_19887,N_10513,N_13373);
and U19888 (N_19888,N_11093,N_12789);
or U19889 (N_19889,N_13674,N_14439);
or U19890 (N_19890,N_11228,N_14486);
xnor U19891 (N_19891,N_13074,N_10516);
or U19892 (N_19892,N_14313,N_14546);
xor U19893 (N_19893,N_14855,N_14681);
and U19894 (N_19894,N_11353,N_12469);
nand U19895 (N_19895,N_10158,N_11247);
or U19896 (N_19896,N_11500,N_13960);
nand U19897 (N_19897,N_13484,N_14060);
xnor U19898 (N_19898,N_13772,N_14458);
xor U19899 (N_19899,N_10521,N_11514);
xor U19900 (N_19900,N_10783,N_10720);
nand U19901 (N_19901,N_11108,N_13010);
or U19902 (N_19902,N_10306,N_11560);
or U19903 (N_19903,N_12522,N_10465);
and U19904 (N_19904,N_11433,N_13624);
nor U19905 (N_19905,N_14419,N_12597);
xnor U19906 (N_19906,N_12890,N_10660);
or U19907 (N_19907,N_14224,N_14816);
or U19908 (N_19908,N_10965,N_13455);
xnor U19909 (N_19909,N_12106,N_10318);
nor U19910 (N_19910,N_10615,N_13631);
or U19911 (N_19911,N_12404,N_11003);
and U19912 (N_19912,N_10580,N_13540);
nand U19913 (N_19913,N_13841,N_13599);
xnor U19914 (N_19914,N_10416,N_13445);
nor U19915 (N_19915,N_11557,N_11229);
and U19916 (N_19916,N_12714,N_10348);
or U19917 (N_19917,N_12697,N_13485);
xnor U19918 (N_19918,N_11620,N_12804);
or U19919 (N_19919,N_10913,N_12089);
xnor U19920 (N_19920,N_12488,N_14672);
or U19921 (N_19921,N_12380,N_11959);
nand U19922 (N_19922,N_11216,N_10525);
nand U19923 (N_19923,N_10894,N_11719);
nand U19924 (N_19924,N_11467,N_13330);
or U19925 (N_19925,N_11699,N_14660);
nor U19926 (N_19926,N_13096,N_11446);
nand U19927 (N_19927,N_13148,N_11117);
and U19928 (N_19928,N_10572,N_10946);
xor U19929 (N_19929,N_12527,N_14539);
nand U19930 (N_19930,N_11926,N_11936);
xor U19931 (N_19931,N_14661,N_13065);
nand U19932 (N_19932,N_12779,N_14406);
xnor U19933 (N_19933,N_13025,N_13951);
and U19934 (N_19934,N_13568,N_11119);
nor U19935 (N_19935,N_10302,N_14747);
xnor U19936 (N_19936,N_14421,N_10569);
nand U19937 (N_19937,N_14420,N_12245);
and U19938 (N_19938,N_10724,N_12020);
and U19939 (N_19939,N_13024,N_14520);
nor U19940 (N_19940,N_13965,N_13615);
xnor U19941 (N_19941,N_10624,N_10346);
or U19942 (N_19942,N_10613,N_14504);
or U19943 (N_19943,N_11409,N_12987);
xor U19944 (N_19944,N_11318,N_12895);
xnor U19945 (N_19945,N_14923,N_12330);
or U19946 (N_19946,N_12553,N_13339);
or U19947 (N_19947,N_12939,N_12166);
or U19948 (N_19948,N_11246,N_11624);
and U19949 (N_19949,N_11733,N_14163);
xor U19950 (N_19950,N_10341,N_13322);
xnor U19951 (N_19951,N_11296,N_13408);
nand U19952 (N_19952,N_10283,N_12668);
nor U19953 (N_19953,N_13616,N_11004);
nor U19954 (N_19954,N_13974,N_11979);
xor U19955 (N_19955,N_14410,N_12665);
nand U19956 (N_19956,N_10340,N_11342);
nand U19957 (N_19957,N_13849,N_10135);
nand U19958 (N_19958,N_10329,N_10383);
xor U19959 (N_19959,N_11782,N_11712);
nand U19960 (N_19960,N_11772,N_14938);
nand U19961 (N_19961,N_10506,N_14671);
nand U19962 (N_19962,N_13565,N_12111);
or U19963 (N_19963,N_13887,N_13126);
and U19964 (N_19964,N_13842,N_10399);
nor U19965 (N_19965,N_11861,N_11789);
nand U19966 (N_19966,N_13102,N_10538);
nand U19967 (N_19967,N_13160,N_10935);
or U19968 (N_19968,N_12089,N_11834);
and U19969 (N_19969,N_12878,N_12998);
or U19970 (N_19970,N_10129,N_10445);
or U19971 (N_19971,N_10939,N_13906);
nand U19972 (N_19972,N_13492,N_12971);
and U19973 (N_19973,N_11958,N_14263);
xor U19974 (N_19974,N_12762,N_11170);
nor U19975 (N_19975,N_14880,N_10498);
xnor U19976 (N_19976,N_14553,N_10451);
or U19977 (N_19977,N_12208,N_12352);
nor U19978 (N_19978,N_12502,N_14187);
xnor U19979 (N_19979,N_10627,N_14330);
or U19980 (N_19980,N_14736,N_10106);
or U19981 (N_19981,N_14997,N_14940);
and U19982 (N_19982,N_13122,N_12401);
and U19983 (N_19983,N_11992,N_10262);
and U19984 (N_19984,N_14796,N_13973);
or U19985 (N_19985,N_11003,N_13848);
or U19986 (N_19986,N_13468,N_13150);
and U19987 (N_19987,N_13104,N_14319);
nand U19988 (N_19988,N_13437,N_13388);
nand U19989 (N_19989,N_11726,N_10801);
nand U19990 (N_19990,N_10728,N_11274);
or U19991 (N_19991,N_10804,N_10193);
xor U19992 (N_19992,N_14855,N_10399);
or U19993 (N_19993,N_14868,N_11913);
nor U19994 (N_19994,N_14888,N_13228);
nor U19995 (N_19995,N_14685,N_10372);
xnor U19996 (N_19996,N_12915,N_14143);
xor U19997 (N_19997,N_13368,N_14995);
nand U19998 (N_19998,N_13216,N_12184);
nand U19999 (N_19999,N_10379,N_13947);
nand UO_0 (O_0,N_18555,N_16174);
and UO_1 (O_1,N_15097,N_17459);
nor UO_2 (O_2,N_19427,N_16010);
and UO_3 (O_3,N_17996,N_16664);
or UO_4 (O_4,N_15078,N_16107);
and UO_5 (O_5,N_16096,N_17074);
or UO_6 (O_6,N_15352,N_19802);
xor UO_7 (O_7,N_16713,N_17222);
and UO_8 (O_8,N_18173,N_17934);
and UO_9 (O_9,N_17643,N_16592);
or UO_10 (O_10,N_18243,N_15554);
and UO_11 (O_11,N_19444,N_16387);
nor UO_12 (O_12,N_18284,N_19624);
nor UO_13 (O_13,N_17630,N_17507);
and UO_14 (O_14,N_18864,N_19907);
or UO_15 (O_15,N_18915,N_16746);
nand UO_16 (O_16,N_15831,N_19918);
or UO_17 (O_17,N_18129,N_16864);
and UO_18 (O_18,N_18247,N_19042);
and UO_19 (O_19,N_18704,N_15779);
or UO_20 (O_20,N_18404,N_15059);
or UO_21 (O_21,N_19975,N_15308);
nor UO_22 (O_22,N_15798,N_19549);
xor UO_23 (O_23,N_17777,N_19872);
nor UO_24 (O_24,N_16776,N_18605);
or UO_25 (O_25,N_15667,N_19262);
and UO_26 (O_26,N_15626,N_19877);
nor UO_27 (O_27,N_16011,N_19919);
nand UO_28 (O_28,N_18447,N_16788);
xor UO_29 (O_29,N_16656,N_15482);
xor UO_30 (O_30,N_16636,N_17456);
nand UO_31 (O_31,N_16936,N_16228);
and UO_32 (O_32,N_17875,N_19789);
nand UO_33 (O_33,N_16185,N_18524);
and UO_34 (O_34,N_19479,N_15011);
or UO_35 (O_35,N_18719,N_19947);
xor UO_36 (O_36,N_16618,N_17712);
xor UO_37 (O_37,N_19951,N_19509);
and UO_38 (O_38,N_18171,N_17056);
nand UO_39 (O_39,N_15280,N_17055);
xor UO_40 (O_40,N_16529,N_16497);
or UO_41 (O_41,N_19803,N_16873);
xor UO_42 (O_42,N_17268,N_16832);
xnor UO_43 (O_43,N_19359,N_16837);
or UO_44 (O_44,N_16694,N_18700);
or UO_45 (O_45,N_15868,N_15670);
nand UO_46 (O_46,N_19871,N_15760);
or UO_47 (O_47,N_17967,N_15620);
nand UO_48 (O_48,N_19633,N_18885);
or UO_49 (O_49,N_15811,N_18633);
and UO_50 (O_50,N_18701,N_17231);
nand UO_51 (O_51,N_18015,N_16934);
and UO_52 (O_52,N_18220,N_19041);
or UO_53 (O_53,N_15592,N_18723);
or UO_54 (O_54,N_18169,N_15141);
nor UO_55 (O_55,N_18384,N_16124);
or UO_56 (O_56,N_19632,N_18549);
and UO_57 (O_57,N_18465,N_15134);
xnor UO_58 (O_58,N_19358,N_16225);
or UO_59 (O_59,N_18735,N_16749);
nand UO_60 (O_60,N_15999,N_16483);
or UO_61 (O_61,N_19010,N_15107);
nor UO_62 (O_62,N_19648,N_16119);
or UO_63 (O_63,N_16649,N_19527);
nor UO_64 (O_64,N_18232,N_17285);
nor UO_65 (O_65,N_15653,N_17527);
nor UO_66 (O_66,N_15187,N_18974);
nor UO_67 (O_67,N_16783,N_19916);
nand UO_68 (O_68,N_18867,N_15402);
and UO_69 (O_69,N_17157,N_18536);
xnor UO_70 (O_70,N_15710,N_18373);
or UO_71 (O_71,N_15629,N_16814);
nor UO_72 (O_72,N_19826,N_19206);
xnor UO_73 (O_73,N_17890,N_17506);
and UO_74 (O_74,N_19581,N_17894);
xnor UO_75 (O_75,N_18418,N_16449);
nand UO_76 (O_76,N_18755,N_19099);
xor UO_77 (O_77,N_18027,N_15053);
xnor UO_78 (O_78,N_18592,N_16210);
nand UO_79 (O_79,N_19917,N_19959);
nor UO_80 (O_80,N_17541,N_17327);
and UO_81 (O_81,N_19596,N_16580);
nand UO_82 (O_82,N_16233,N_19186);
xor UO_83 (O_83,N_18625,N_17363);
nand UO_84 (O_84,N_18250,N_19412);
and UO_85 (O_85,N_18399,N_15627);
and UO_86 (O_86,N_19554,N_18050);
xor UO_87 (O_87,N_18333,N_15062);
nand UO_88 (O_88,N_15372,N_16921);
and UO_89 (O_89,N_19120,N_17435);
nor UO_90 (O_90,N_16595,N_19171);
nand UO_91 (O_91,N_17917,N_17679);
or UO_92 (O_92,N_16614,N_17431);
or UO_93 (O_93,N_17426,N_18789);
or UO_94 (O_94,N_19403,N_18416);
and UO_95 (O_95,N_15228,N_15919);
nor UO_96 (O_96,N_19642,N_16028);
or UO_97 (O_97,N_17633,N_16950);
nor UO_98 (O_98,N_19183,N_17622);
nand UO_99 (O_99,N_19004,N_18034);
or UO_100 (O_100,N_18068,N_19921);
and UO_101 (O_101,N_17878,N_19544);
xor UO_102 (O_102,N_15431,N_18726);
nand UO_103 (O_103,N_16286,N_18016);
and UO_104 (O_104,N_15874,N_15366);
xor UO_105 (O_105,N_16771,N_18803);
or UO_106 (O_106,N_19843,N_15476);
or UO_107 (O_107,N_19279,N_15600);
nand UO_108 (O_108,N_16520,N_16253);
or UO_109 (O_109,N_19822,N_15736);
xnor UO_110 (O_110,N_17012,N_15396);
xnor UO_111 (O_111,N_18707,N_18586);
and UO_112 (O_112,N_17753,N_18550);
nand UO_113 (O_113,N_18215,N_19708);
nand UO_114 (O_114,N_15878,N_18811);
and UO_115 (O_115,N_19253,N_17690);
or UO_116 (O_116,N_18074,N_15698);
and UO_117 (O_117,N_16082,N_19266);
or UO_118 (O_118,N_16710,N_15666);
or UO_119 (O_119,N_16019,N_18998);
nor UO_120 (O_120,N_16725,N_15504);
and UO_121 (O_121,N_18358,N_18347);
or UO_122 (O_122,N_18329,N_18795);
or UO_123 (O_123,N_19376,N_15944);
or UO_124 (O_124,N_19326,N_19053);
xnor UO_125 (O_125,N_16365,N_17422);
xor UO_126 (O_126,N_19553,N_15037);
nand UO_127 (O_127,N_16163,N_19863);
or UO_128 (O_128,N_17707,N_17427);
xnor UO_129 (O_129,N_16468,N_15392);
xor UO_130 (O_130,N_19059,N_18679);
or UO_131 (O_131,N_17759,N_17884);
xnor UO_132 (O_132,N_19345,N_18944);
nor UO_133 (O_133,N_17742,N_15624);
or UO_134 (O_134,N_15573,N_16973);
and UO_135 (O_135,N_16275,N_16659);
or UO_136 (O_136,N_15112,N_16963);
nor UO_137 (O_137,N_17142,N_15935);
nor UO_138 (O_138,N_15942,N_18315);
and UO_139 (O_139,N_19374,N_17810);
and UO_140 (O_140,N_18466,N_17519);
xor UO_141 (O_141,N_15481,N_15010);
nor UO_142 (O_142,N_15799,N_16277);
nor UO_143 (O_143,N_19067,N_19923);
and UO_144 (O_144,N_17616,N_15315);
nor UO_145 (O_145,N_18023,N_18834);
nand UO_146 (O_146,N_17562,N_16232);
xnor UO_147 (O_147,N_16142,N_18567);
xor UO_148 (O_148,N_16915,N_15379);
xnor UO_149 (O_149,N_16889,N_18890);
and UO_150 (O_150,N_15047,N_16698);
nand UO_151 (O_151,N_15892,N_19626);
and UO_152 (O_152,N_19770,N_18102);
nand UO_153 (O_153,N_16573,N_18619);
nor UO_154 (O_154,N_17662,N_16866);
and UO_155 (O_155,N_18649,N_19050);
nand UO_156 (O_156,N_17105,N_16782);
nor UO_157 (O_157,N_19566,N_19697);
xor UO_158 (O_158,N_19208,N_16371);
and UO_159 (O_159,N_16463,N_15715);
and UO_160 (O_160,N_19720,N_17156);
nand UO_161 (O_161,N_19893,N_16406);
nor UO_162 (O_162,N_16103,N_19982);
nor UO_163 (O_163,N_18281,N_19800);
xnor UO_164 (O_164,N_18519,N_18797);
nor UO_165 (O_165,N_15483,N_18954);
or UO_166 (O_166,N_16125,N_16147);
nor UO_167 (O_167,N_15227,N_18613);
nor UO_168 (O_168,N_17444,N_19338);
xnor UO_169 (O_169,N_16536,N_19833);
nand UO_170 (O_170,N_19997,N_19013);
xor UO_171 (O_171,N_15336,N_16421);
xnor UO_172 (O_172,N_17388,N_19523);
nor UO_173 (O_173,N_16440,N_16385);
xor UO_174 (O_174,N_17607,N_19560);
nand UO_175 (O_175,N_18694,N_17325);
or UO_176 (O_176,N_17714,N_17596);
xor UO_177 (O_177,N_16744,N_17301);
or UO_178 (O_178,N_15310,N_17460);
and UO_179 (O_179,N_15035,N_17711);
nand UO_180 (O_180,N_18893,N_17956);
or UO_181 (O_181,N_17385,N_15327);
nand UO_182 (O_182,N_15883,N_19330);
nand UO_183 (O_183,N_18774,N_15344);
xnor UO_184 (O_184,N_15536,N_17017);
and UO_185 (O_185,N_18033,N_17421);
and UO_186 (O_186,N_15996,N_18073);
and UO_187 (O_187,N_16803,N_19768);
nor UO_188 (O_188,N_17628,N_18515);
and UO_189 (O_189,N_16789,N_17389);
or UO_190 (O_190,N_19033,N_16550);
and UO_191 (O_191,N_17634,N_17371);
nand UO_192 (O_192,N_19504,N_17829);
or UO_193 (O_193,N_16352,N_16653);
nand UO_194 (O_194,N_16216,N_15155);
and UO_195 (O_195,N_19943,N_17529);
xor UO_196 (O_196,N_16677,N_19933);
nand UO_197 (O_197,N_15085,N_16917);
and UO_198 (O_198,N_18455,N_19589);
xor UO_199 (O_199,N_19847,N_18327);
xor UO_200 (O_200,N_16894,N_15314);
and UO_201 (O_201,N_17227,N_15075);
or UO_202 (O_202,N_17042,N_15083);
nand UO_203 (O_203,N_15837,N_16999);
xnor UO_204 (O_204,N_18963,N_18420);
or UO_205 (O_205,N_17936,N_15603);
nor UO_206 (O_206,N_19468,N_18158);
or UO_207 (O_207,N_17754,N_15928);
and UO_208 (O_208,N_15304,N_15196);
and UO_209 (O_209,N_17481,N_18681);
and UO_210 (O_210,N_19868,N_15915);
xnor UO_211 (O_211,N_19119,N_15478);
xnor UO_212 (O_212,N_19732,N_18246);
and UO_213 (O_213,N_18394,N_15084);
and UO_214 (O_214,N_17287,N_18752);
or UO_215 (O_215,N_17785,N_16637);
and UO_216 (O_216,N_18288,N_19144);
nor UO_217 (O_217,N_17373,N_18110);
nand UO_218 (O_218,N_16538,N_18037);
nor UO_219 (O_219,N_18135,N_15466);
xor UO_220 (O_220,N_15091,N_19252);
nand UO_221 (O_221,N_19239,N_17136);
or UO_222 (O_222,N_19673,N_19836);
nor UO_223 (O_223,N_17603,N_18643);
nand UO_224 (O_224,N_16646,N_15370);
or UO_225 (O_225,N_16150,N_15044);
xnor UO_226 (O_226,N_15726,N_17534);
nand UO_227 (O_227,N_18209,N_15279);
nand UO_228 (O_228,N_16102,N_17284);
and UO_229 (O_229,N_15998,N_15087);
nor UO_230 (O_230,N_19852,N_17366);
xnor UO_231 (O_231,N_17896,N_16402);
nor UO_232 (O_232,N_18172,N_15976);
xor UO_233 (O_233,N_16162,N_18879);
nand UO_234 (O_234,N_17262,N_19618);
nand UO_235 (O_235,N_17729,N_18968);
and UO_236 (O_236,N_18262,N_16647);
nor UO_237 (O_237,N_18386,N_16242);
nor UO_238 (O_238,N_19324,N_16109);
xor UO_239 (O_239,N_16711,N_19762);
nor UO_240 (O_240,N_18510,N_18067);
nor UO_241 (O_241,N_17434,N_16527);
and UO_242 (O_242,N_16063,N_16346);
nor UO_243 (O_243,N_19623,N_19363);
xor UO_244 (O_244,N_17642,N_16298);
nand UO_245 (O_245,N_19078,N_19988);
nor UO_246 (O_246,N_19857,N_15444);
and UO_247 (O_247,N_16904,N_15008);
nor UO_248 (O_248,N_15438,N_19433);
or UO_249 (O_249,N_15079,N_15411);
and UO_250 (O_250,N_16422,N_19277);
nor UO_251 (O_251,N_17577,N_18750);
nand UO_252 (O_252,N_15341,N_17860);
nand UO_253 (O_253,N_15572,N_18545);
nand UO_254 (O_254,N_15198,N_16762);
xor UO_255 (O_255,N_18588,N_19023);
nand UO_256 (O_256,N_16015,N_15386);
and UO_257 (O_257,N_17584,N_16675);
or UO_258 (O_258,N_17764,N_17469);
xnor UO_259 (O_259,N_18622,N_16716);
xnor UO_260 (O_260,N_17033,N_18433);
nor UO_261 (O_261,N_17653,N_17300);
nand UO_262 (O_262,N_19325,N_16770);
nor UO_263 (O_263,N_19986,N_17874);
or UO_264 (O_264,N_17597,N_17181);
xnor UO_265 (O_265,N_19411,N_19094);
or UO_266 (O_266,N_16196,N_16414);
nand UO_267 (O_267,N_15284,N_17407);
and UO_268 (O_268,N_19726,N_18140);
xnor UO_269 (O_269,N_17220,N_17044);
and UO_270 (O_270,N_19440,N_19488);
xnor UO_271 (O_271,N_18261,N_16420);
or UO_272 (O_272,N_15317,N_15166);
or UO_273 (O_273,N_15525,N_18159);
and UO_274 (O_274,N_18663,N_16207);
or UO_275 (O_275,N_19556,N_16736);
xnor UO_276 (O_276,N_18430,N_17261);
nor UO_277 (O_277,N_16479,N_19601);
and UO_278 (O_278,N_19090,N_19713);
nand UO_279 (O_279,N_17818,N_17304);
nand UO_280 (O_280,N_16672,N_19804);
nand UO_281 (O_281,N_16415,N_19670);
nand UO_282 (O_282,N_18297,N_16035);
nand UO_283 (O_283,N_19141,N_18423);
and UO_284 (O_284,N_18448,N_16978);
nor UO_285 (O_285,N_18504,N_17492);
xnor UO_286 (O_286,N_17416,N_19929);
nor UO_287 (O_287,N_16087,N_18579);
xor UO_288 (O_288,N_18277,N_15383);
or UO_289 (O_289,N_18117,N_19784);
nor UO_290 (O_290,N_18636,N_18665);
xor UO_291 (O_291,N_18478,N_16780);
or UO_292 (O_292,N_19228,N_16938);
xnor UO_293 (O_293,N_19920,N_19678);
nand UO_294 (O_294,N_16053,N_16942);
nand UO_295 (O_295,N_18689,N_18730);
nand UO_296 (O_296,N_15510,N_15565);
nor UO_297 (O_297,N_16160,N_17931);
and UO_298 (O_298,N_15730,N_18930);
or UO_299 (O_299,N_15556,N_15321);
and UO_300 (O_300,N_18398,N_16624);
xor UO_301 (O_301,N_19038,N_17848);
nand UO_302 (O_302,N_17491,N_19952);
and UO_303 (O_303,N_18513,N_16733);
nand UO_304 (O_304,N_18532,N_16608);
and UO_305 (O_305,N_17945,N_16327);
xor UO_306 (O_306,N_16926,N_17194);
or UO_307 (O_307,N_19323,N_19408);
nor UO_308 (O_308,N_15029,N_17820);
nand UO_309 (O_309,N_17216,N_19735);
xnor UO_310 (O_310,N_17219,N_18467);
nand UO_311 (O_311,N_18990,N_17163);
or UO_312 (O_312,N_16123,N_17836);
or UO_313 (O_313,N_15890,N_18363);
or UO_314 (O_314,N_15003,N_18417);
nor UO_315 (O_315,N_16979,N_19382);
nand UO_316 (O_316,N_19774,N_15328);
and UO_317 (O_317,N_18630,N_15407);
or UO_318 (O_318,N_15113,N_18842);
xor UO_319 (O_319,N_18731,N_19514);
nor UO_320 (O_320,N_19970,N_18717);
or UO_321 (O_321,N_18094,N_19234);
nand UO_322 (O_322,N_16471,N_18598);
nor UO_323 (O_323,N_19453,N_18419);
nor UO_324 (O_324,N_15264,N_15121);
xor UO_325 (O_325,N_15448,N_15738);
or UO_326 (O_326,N_15032,N_18537);
xnor UO_327 (O_327,N_16001,N_18236);
nor UO_328 (O_328,N_18368,N_15540);
or UO_329 (O_329,N_15244,N_18491);
nor UO_330 (O_330,N_17828,N_17992);
xnor UO_331 (O_331,N_19602,N_17257);
xnor UO_332 (O_332,N_18224,N_16845);
and UO_333 (O_333,N_17661,N_19992);
nor UO_334 (O_334,N_15982,N_16436);
nand UO_335 (O_335,N_16296,N_15122);
or UO_336 (O_336,N_16351,N_15302);
and UO_337 (O_337,N_19664,N_18383);
nor UO_338 (O_338,N_17240,N_17508);
and UO_339 (O_339,N_16335,N_16775);
and UO_340 (O_340,N_18995,N_18911);
or UO_341 (O_341,N_19261,N_16029);
and UO_342 (O_342,N_17799,N_19035);
xor UO_343 (O_343,N_18366,N_15455);
or UO_344 (O_344,N_15421,N_19763);
nor UO_345 (O_345,N_16732,N_16093);
and UO_346 (O_346,N_16720,N_18624);
or UO_347 (O_347,N_19818,N_17648);
nand UO_348 (O_348,N_19892,N_18364);
nor UO_349 (O_349,N_17530,N_15329);
nor UO_350 (O_350,N_16060,N_16642);
and UO_351 (O_351,N_17104,N_19350);
nand UO_352 (O_352,N_17516,N_17817);
nand UO_353 (O_353,N_19257,N_16426);
or UO_354 (O_354,N_19162,N_16175);
nor UO_355 (O_355,N_15414,N_19701);
xnor UO_356 (O_356,N_19361,N_15972);
nor UO_357 (O_357,N_18566,N_19793);
or UO_358 (O_358,N_15991,N_19728);
and UO_359 (O_359,N_19398,N_19927);
and UO_360 (O_360,N_17573,N_17182);
and UO_361 (O_361,N_19886,N_17564);
nand UO_362 (O_362,N_18156,N_16126);
nand UO_363 (O_363,N_17167,N_18035);
and UO_364 (O_364,N_18044,N_16772);
or UO_365 (O_365,N_19675,N_15225);
nor UO_366 (O_366,N_15686,N_17709);
xnor UO_367 (O_367,N_15619,N_17950);
and UO_368 (O_368,N_18179,N_18442);
nor UO_369 (O_369,N_15849,N_19354);
nor UO_370 (O_370,N_18746,N_17805);
or UO_371 (O_371,N_18502,N_15115);
and UO_372 (O_372,N_15384,N_19238);
and UO_373 (O_373,N_19771,N_18562);
nor UO_374 (O_374,N_16234,N_19295);
and UO_375 (O_375,N_17706,N_15722);
nand UO_376 (O_376,N_15790,N_18675);
xnor UO_377 (O_377,N_19574,N_15827);
nor UO_378 (O_378,N_19034,N_16553);
or UO_379 (O_379,N_16157,N_17187);
nand UO_380 (O_380,N_18472,N_15480);
xor UO_381 (O_381,N_17451,N_19087);
or UO_382 (O_382,N_18326,N_17265);
nand UO_383 (O_383,N_17612,N_15777);
nor UO_384 (O_384,N_17344,N_18943);
nor UO_385 (O_385,N_18484,N_18907);
and UO_386 (O_386,N_16899,N_19658);
or UO_387 (O_387,N_17927,N_16180);
and UO_388 (O_388,N_17358,N_18047);
or UO_389 (O_389,N_19582,N_19368);
xor UO_390 (O_390,N_16472,N_19968);
or UO_391 (O_391,N_16236,N_19397);
and UO_392 (O_392,N_17682,N_19765);
or UO_393 (O_393,N_15145,N_16222);
or UO_394 (O_394,N_19093,N_15829);
or UO_395 (O_395,N_19320,N_19605);
xnor UO_396 (O_396,N_18111,N_18964);
and UO_397 (O_397,N_19296,N_17401);
and UO_398 (O_398,N_18408,N_17380);
xnor UO_399 (O_399,N_15348,N_16954);
nor UO_400 (O_400,N_15541,N_16676);
nor UO_401 (O_401,N_18798,N_18107);
and UO_402 (O_402,N_16517,N_17600);
xor UO_403 (O_403,N_17310,N_18053);
or UO_404 (O_404,N_17217,N_18535);
or UO_405 (O_405,N_15013,N_16360);
xnor UO_406 (O_406,N_19275,N_18350);
or UO_407 (O_407,N_19798,N_18662);
and UO_408 (O_408,N_17790,N_17062);
nor UO_409 (O_409,N_16765,N_17998);
nand UO_410 (O_410,N_17567,N_16598);
and UO_411 (O_411,N_19445,N_18984);
or UO_412 (O_412,N_17740,N_15903);
nand UO_413 (O_413,N_17502,N_17767);
xor UO_414 (O_414,N_15521,N_18606);
nor UO_415 (O_415,N_17346,N_16095);
nand UO_416 (O_416,N_18621,N_17902);
xor UO_417 (O_417,N_19475,N_16247);
nor UO_418 (O_418,N_19215,N_18608);
or UO_419 (O_419,N_19052,N_15439);
nand UO_420 (O_420,N_15498,N_19245);
nand UO_421 (O_421,N_15707,N_16952);
xor UO_422 (O_422,N_17239,N_17542);
or UO_423 (O_423,N_16840,N_16545);
or UO_424 (O_424,N_19015,N_19799);
nand UO_425 (O_425,N_16369,N_15989);
nor UO_426 (O_426,N_16968,N_19967);
xnor UO_427 (O_427,N_19645,N_18096);
xnor UO_428 (O_428,N_15733,N_16910);
nor UO_429 (O_429,N_18590,N_17132);
nand UO_430 (O_430,N_17649,N_18794);
and UO_431 (O_431,N_15485,N_19101);
or UO_432 (O_432,N_17910,N_15207);
xnor UO_433 (O_433,N_15009,N_17505);
or UO_434 (O_434,N_17968,N_16502);
and UO_435 (O_435,N_16961,N_18301);
or UO_436 (O_436,N_15248,N_16975);
and UO_437 (O_437,N_16081,N_16092);
and UO_438 (O_438,N_16416,N_17453);
nand UO_439 (O_439,N_19410,N_17798);
nor UO_440 (O_440,N_17585,N_18713);
or UO_441 (O_441,N_17771,N_15019);
xor UO_442 (O_442,N_19938,N_15608);
nand UO_443 (O_443,N_17765,N_17851);
or UO_444 (O_444,N_19704,N_18387);
and UO_445 (O_445,N_16184,N_16108);
and UO_446 (O_446,N_19932,N_17166);
or UO_447 (O_447,N_16700,N_18312);
or UO_448 (O_448,N_18201,N_17440);
nand UO_449 (O_449,N_18884,N_17842);
nor UO_450 (O_450,N_17420,N_16674);
xnor UO_451 (O_451,N_19724,N_18542);
or UO_452 (O_452,N_16717,N_17233);
and UO_453 (O_453,N_16356,N_19526);
or UO_454 (O_454,N_17856,N_19996);
nor UO_455 (O_455,N_15168,N_15066);
or UO_456 (O_456,N_17034,N_16893);
nor UO_457 (O_457,N_18365,N_19519);
nand UO_458 (O_458,N_15233,N_16843);
or UO_459 (O_459,N_18607,N_19842);
nand UO_460 (O_460,N_18471,N_19168);
or UO_461 (O_461,N_19205,N_16524);
or UO_462 (O_462,N_19106,N_17922);
nand UO_463 (O_463,N_16606,N_16578);
nand UO_464 (O_464,N_15410,N_19231);
nand UO_465 (O_465,N_18290,N_18126);
nor UO_466 (O_466,N_19901,N_18677);
and UO_467 (O_467,N_17164,N_18775);
xor UO_468 (O_468,N_19734,N_15997);
xor UO_469 (O_469,N_17908,N_15508);
xnor UO_470 (O_470,N_16164,N_16829);
nand UO_471 (O_471,N_19156,N_18060);
xnor UO_472 (O_472,N_17117,N_18934);
xor UO_473 (O_473,N_19191,N_19585);
nand UO_474 (O_474,N_15948,N_15735);
nor UO_475 (O_475,N_19219,N_17667);
and UO_476 (O_476,N_17303,N_19969);
xor UO_477 (O_477,N_17755,N_15387);
and UO_478 (O_478,N_18935,N_17354);
nand UO_479 (O_479,N_19429,N_18083);
nor UO_480 (O_480,N_19117,N_17887);
nand UO_481 (O_481,N_17343,N_19853);
nand UO_482 (O_482,N_19603,N_18596);
xor UO_483 (O_483,N_16226,N_18889);
and UO_484 (O_484,N_19511,N_15358);
or UO_485 (O_485,N_15263,N_19471);
nand UO_486 (O_486,N_15893,N_18492);
xor UO_487 (O_487,N_18428,N_18054);
nand UO_488 (O_488,N_17943,N_17028);
xor UO_489 (O_489,N_16302,N_19114);
nand UO_490 (O_490,N_18881,N_17395);
xnor UO_491 (O_491,N_19881,N_18918);
xor UO_492 (O_492,N_16445,N_16355);
or UO_493 (O_493,N_15203,N_17610);
nand UO_494 (O_494,N_19964,N_18085);
and UO_495 (O_495,N_17009,N_16359);
and UO_496 (O_496,N_19913,N_18520);
xor UO_497 (O_497,N_19360,N_18882);
xor UO_498 (O_498,N_16061,N_19812);
nor UO_499 (O_499,N_15428,N_19532);
xor UO_500 (O_500,N_18199,N_15217);
or UO_501 (O_501,N_18604,N_16533);
nand UO_502 (O_502,N_16325,N_17669);
nor UO_503 (O_503,N_18320,N_18287);
and UO_504 (O_504,N_15356,N_16344);
or UO_505 (O_505,N_17885,N_19729);
and UO_506 (O_506,N_15371,N_19570);
nor UO_507 (O_507,N_15323,N_16202);
or UO_508 (O_508,N_15130,N_16542);
nor UO_509 (O_509,N_18256,N_15992);
or UO_510 (O_510,N_15369,N_19819);
nand UO_511 (O_511,N_18791,N_17356);
xnor UO_512 (O_512,N_16178,N_18474);
nor UO_513 (O_513,N_19346,N_16807);
nor UO_514 (O_514,N_15434,N_19031);
xnor UO_515 (O_515,N_18644,N_17589);
nand UO_516 (O_516,N_17093,N_16551);
nand UO_517 (O_517,N_16278,N_16340);
xor UO_518 (O_518,N_18062,N_16380);
or UO_519 (O_519,N_17879,N_19256);
nor UO_520 (O_520,N_17543,N_17443);
nor UO_521 (O_521,N_17883,N_17384);
and UO_522 (O_522,N_17417,N_16328);
nand UO_523 (O_523,N_19578,N_18876);
or UO_524 (O_524,N_19794,N_16867);
and UO_525 (O_525,N_18196,N_15192);
nor UO_526 (O_526,N_18696,N_17605);
nor UO_527 (O_527,N_17226,N_17832);
or UO_528 (O_528,N_16409,N_15473);
nand UO_529 (O_529,N_18498,N_18177);
nand UO_530 (O_530,N_15869,N_18210);
xnor UO_531 (O_531,N_16179,N_19264);
or UO_532 (O_532,N_17704,N_19493);
xor UO_533 (O_533,N_16094,N_17313);
or UO_534 (O_534,N_15191,N_17839);
or UO_535 (O_535,N_15936,N_19143);
nor UO_536 (O_536,N_18506,N_19305);
nor UO_537 (O_537,N_17857,N_18600);
nand UO_538 (O_538,N_15157,N_18453);
and UO_539 (O_539,N_17901,N_18868);
xnor UO_540 (O_540,N_19515,N_19148);
nand UO_541 (O_541,N_17705,N_18923);
nand UO_542 (O_542,N_18572,N_17695);
or UO_543 (O_543,N_17763,N_15979);
nor UO_544 (O_544,N_15324,N_19902);
or UO_545 (O_545,N_16182,N_18850);
or UO_546 (O_546,N_18988,N_16072);
nor UO_547 (O_547,N_17847,N_17550);
nor UO_548 (O_548,N_17770,N_16381);
and UO_549 (O_549,N_17073,N_17168);
or UO_550 (O_550,N_17576,N_19108);
and UO_551 (O_551,N_18711,N_15361);
or UO_552 (O_552,N_17248,N_16276);
nor UO_553 (O_553,N_15290,N_15949);
or UO_554 (O_554,N_17861,N_18145);
nand UO_555 (O_555,N_16321,N_16515);
or UO_556 (O_556,N_19250,N_19421);
and UO_557 (O_557,N_19599,N_16303);
xor UO_558 (O_558,N_16571,N_15836);
nor UO_559 (O_559,N_16049,N_18950);
and UO_560 (O_560,N_19116,N_18105);
and UO_561 (O_561,N_16265,N_19150);
nand UO_562 (O_562,N_19291,N_16922);
nand UO_563 (O_563,N_18828,N_19155);
and UO_564 (O_564,N_17381,N_17904);
and UO_565 (O_565,N_17685,N_17914);
and UO_566 (O_566,N_17038,N_19054);
nor UO_567 (O_567,N_16332,N_18254);
xnor UO_568 (O_568,N_16858,N_17719);
and UO_569 (O_569,N_19809,N_17930);
nand UO_570 (O_570,N_18438,N_16752);
or UO_571 (O_571,N_19334,N_17893);
and UO_572 (O_572,N_15295,N_16575);
or UO_573 (O_573,N_19441,N_19776);
nor UO_574 (O_574,N_16892,N_19367);
nor UO_575 (O_575,N_15640,N_18962);
or UO_576 (O_576,N_17961,N_19008);
xnor UO_577 (O_577,N_15177,N_18229);
or UO_578 (O_578,N_16432,N_16870);
or UO_579 (O_579,N_15813,N_18091);
xor UO_580 (O_580,N_16727,N_18330);
and UO_581 (O_581,N_15232,N_19169);
nor UO_582 (O_582,N_16407,N_17415);
nand UO_583 (O_583,N_18112,N_15787);
nor UO_584 (O_584,N_19159,N_17170);
xor UO_585 (O_585,N_15891,N_15389);
or UO_586 (O_586,N_19832,N_18334);
or UO_587 (O_587,N_18002,N_16288);
or UO_588 (O_588,N_16790,N_19751);
xnor UO_589 (O_589,N_15757,N_16104);
or UO_590 (O_590,N_17243,N_17863);
xor UO_591 (O_591,N_18877,N_19752);
nand UO_592 (O_592,N_18059,N_15126);
or UO_593 (O_593,N_15172,N_18257);
or UO_594 (O_594,N_15804,N_18991);
or UO_595 (O_595,N_16745,N_17159);
xnor UO_596 (O_596,N_17873,N_15974);
or UO_597 (O_597,N_16946,N_19267);
and UO_598 (O_598,N_16259,N_17405);
or UO_599 (O_599,N_18522,N_18977);
nand UO_600 (O_600,N_15658,N_19687);
nand UO_601 (O_601,N_17213,N_16494);
nor UO_602 (O_602,N_15486,N_18339);
xnor UO_603 (O_603,N_18431,N_16537);
or UO_604 (O_604,N_17061,N_17656);
or UO_605 (O_605,N_17247,N_17374);
and UO_606 (O_606,N_17666,N_17185);
nand UO_607 (O_607,N_18792,N_17035);
xor UO_608 (O_608,N_15380,N_15253);
xor UO_609 (O_609,N_16006,N_18787);
nand UO_610 (O_610,N_15704,N_16261);
nor UO_611 (O_611,N_15440,N_15353);
xor UO_612 (O_612,N_16833,N_15491);
and UO_613 (O_613,N_17973,N_15423);
and UO_614 (O_614,N_17521,N_16512);
nand UO_615 (O_615,N_15254,N_16684);
nand UO_616 (O_616,N_15981,N_15006);
nor UO_617 (O_617,N_19955,N_17155);
xnor UO_618 (O_618,N_16742,N_19564);
nand UO_619 (O_619,N_18260,N_16523);
nand UO_620 (O_620,N_17811,N_19772);
nor UO_621 (O_621,N_16281,N_18058);
and UO_622 (O_622,N_19494,N_16918);
or UO_623 (O_623,N_19513,N_18010);
and UO_624 (O_624,N_15294,N_17466);
nand UO_625 (O_625,N_15306,N_17414);
nand UO_626 (O_626,N_17497,N_17958);
and UO_627 (O_627,N_17555,N_18426);
or UO_628 (O_628,N_18282,N_19142);
xor UO_629 (O_629,N_16971,N_16042);
and UO_630 (O_630,N_15394,N_19580);
nor UO_631 (O_631,N_15870,N_17057);
or UO_632 (O_632,N_17544,N_16490);
or UO_633 (O_633,N_18009,N_15450);
and UO_634 (O_634,N_18829,N_15454);
and UO_635 (O_635,N_17476,N_15218);
and UO_636 (O_636,N_18994,N_18610);
or UO_637 (O_637,N_17907,N_17436);
and UO_638 (O_638,N_17402,N_16322);
and UO_639 (O_639,N_17269,N_18843);
xnor UO_640 (O_640,N_16213,N_16813);
nand UO_641 (O_641,N_19195,N_16648);
xnor UO_642 (O_642,N_19399,N_16404);
or UO_643 (O_643,N_19060,N_18558);
and UO_644 (O_644,N_16777,N_16129);
and UO_645 (O_645,N_16331,N_19721);
or UO_646 (O_646,N_16574,N_16341);
nor UO_647 (O_647,N_17060,N_15144);
xor UO_648 (O_648,N_18680,N_15100);
nand UO_649 (O_649,N_16956,N_15477);
xnor UO_650 (O_650,N_17047,N_15834);
nor UO_651 (O_651,N_16263,N_17253);
and UO_652 (O_652,N_16584,N_18344);
xnor UO_653 (O_653,N_16827,N_16547);
xor UO_654 (O_654,N_19512,N_19387);
xnor UO_655 (O_655,N_19930,N_18902);
nand UO_656 (O_656,N_15731,N_16014);
nor UO_657 (O_657,N_16992,N_17458);
and UO_658 (O_658,N_16375,N_17862);
nand UO_659 (O_659,N_18155,N_18862);
nand UO_660 (O_660,N_19714,N_17691);
xnor UO_661 (O_661,N_17001,N_19301);
xor UO_662 (O_662,N_18580,N_19025);
and UO_663 (O_663,N_18582,N_15339);
or UO_664 (O_664,N_16132,N_17315);
or UO_665 (O_665,N_17470,N_18148);
nor UO_666 (O_666,N_16903,N_17846);
nand UO_667 (O_667,N_16683,N_19133);
xnor UO_668 (O_668,N_15591,N_19529);
nand UO_669 (O_669,N_15301,N_16787);
and UO_670 (O_670,N_19173,N_15634);
nand UO_671 (O_671,N_15583,N_16928);
and UO_672 (O_672,N_18457,N_18161);
xor UO_673 (O_673,N_17983,N_18221);
nor UO_674 (O_674,N_18866,N_15178);
nand UO_675 (O_675,N_16484,N_15840);
or UO_676 (O_676,N_19547,N_15775);
and UO_677 (O_677,N_18040,N_15795);
and UO_678 (O_678,N_15563,N_16556);
and UO_679 (O_679,N_19125,N_19655);
or UO_680 (O_680,N_15119,N_15672);
and UO_681 (O_681,N_18230,N_17207);
xor UO_682 (O_682,N_18556,N_16729);
and UO_683 (O_683,N_15680,N_15500);
nand UO_684 (O_684,N_19828,N_17548);
and UO_685 (O_685,N_17064,N_15801);
or UO_686 (O_686,N_15727,N_18683);
and UO_687 (O_687,N_16590,N_18518);
nand UO_688 (O_688,N_15266,N_17412);
and UO_689 (O_689,N_17094,N_17872);
or UO_690 (O_690,N_15616,N_16304);
xor UO_691 (O_691,N_16844,N_18920);
or UO_692 (O_692,N_17593,N_18768);
xnor UO_693 (O_693,N_17728,N_17118);
xnor UO_694 (O_694,N_16881,N_17457);
xor UO_695 (O_695,N_17978,N_18898);
nor UO_696 (O_696,N_16431,N_18661);
xnor UO_697 (O_697,N_17102,N_17095);
nand UO_698 (O_698,N_18439,N_15692);
nand UO_699 (O_699,N_15946,N_15060);
nor UO_700 (O_700,N_19680,N_16037);
or UO_701 (O_701,N_17951,N_19674);
nor UO_702 (O_702,N_17146,N_15520);
and UO_703 (O_703,N_18204,N_17722);
nor UO_704 (O_704,N_18933,N_19147);
xor UO_705 (O_705,N_17424,N_16521);
or UO_706 (O_706,N_18092,N_16661);
xor UO_707 (O_707,N_15319,N_19958);
or UO_708 (O_708,N_17556,N_19122);
xor UO_709 (O_709,N_16991,N_16250);
nand UO_710 (O_710,N_18184,N_15269);
xnor UO_711 (O_711,N_17318,N_19859);
xnor UO_712 (O_712,N_18367,N_18784);
nor UO_713 (O_713,N_19285,N_19703);
or UO_714 (O_714,N_16419,N_16701);
xnor UO_715 (O_715,N_16924,N_15676);
or UO_716 (O_716,N_19331,N_18629);
nand UO_717 (O_717,N_15663,N_19531);
xnor UO_718 (O_718,N_15409,N_18845);
and UO_719 (O_719,N_19679,N_19196);
nand UO_720 (O_720,N_17204,N_18021);
or UO_721 (O_721,N_15199,N_16203);
or UO_722 (O_722,N_16383,N_19370);
and UO_723 (O_723,N_15912,N_17149);
or UO_724 (O_724,N_18846,N_17067);
and UO_725 (O_725,N_16805,N_15960);
and UO_726 (O_726,N_18182,N_16411);
nor UO_727 (O_727,N_15151,N_19999);
and UO_728 (O_728,N_17235,N_18006);
or UO_729 (O_729,N_17640,N_17926);
or UO_730 (O_730,N_17328,N_15743);
or UO_731 (O_731,N_19095,N_15830);
xor UO_732 (O_732,N_15633,N_19153);
nand UO_733 (O_733,N_19681,N_16144);
or UO_734 (O_734,N_16013,N_15424);
or UO_735 (O_735,N_18456,N_15293);
nor UO_736 (O_736,N_16972,N_18166);
nor UO_737 (O_737,N_19823,N_19838);
nand UO_738 (O_738,N_15004,N_16667);
xor UO_739 (O_739,N_15190,N_15971);
xnor UO_740 (O_740,N_16268,N_16249);
nor UO_741 (O_741,N_17377,N_15182);
nand UO_742 (O_742,N_15355,N_19273);
xor UO_743 (O_743,N_15229,N_18553);
or UO_744 (O_744,N_17403,N_18913);
and UO_745 (O_745,N_16778,N_16318);
and UO_746 (O_746,N_18319,N_18706);
and UO_747 (O_747,N_15577,N_16198);
or UO_748 (O_748,N_18796,N_18987);
xor UO_749 (O_749,N_15274,N_15842);
nor UO_750 (O_750,N_15288,N_17128);
nand UO_751 (O_751,N_15506,N_19057);
and UO_752 (O_752,N_15399,N_15511);
or UO_753 (O_753,N_17059,N_15068);
nor UO_754 (O_754,N_17224,N_19889);
nor UO_755 (O_755,N_17841,N_18217);
or UO_756 (O_756,N_18815,N_17096);
or UO_757 (O_757,N_16681,N_19414);
and UO_758 (O_758,N_18275,N_17337);
nand UO_759 (O_759,N_16818,N_16173);
or UO_760 (O_760,N_16927,N_19805);
nand UO_761 (O_761,N_19230,N_17808);
nor UO_762 (O_762,N_15557,N_17258);
and UO_763 (O_763,N_17700,N_17158);
xnor UO_764 (O_764,N_15041,N_19562);
nand UO_765 (O_765,N_16603,N_16835);
or UO_766 (O_766,N_16386,N_19481);
nand UO_767 (O_767,N_16320,N_15705);
or UO_768 (O_768,N_19380,N_17522);
nand UO_769 (O_769,N_15251,N_17739);
xnor UO_770 (O_770,N_16859,N_17749);
nand UO_771 (O_771,N_15544,N_19344);
or UO_772 (O_772,N_15001,N_15530);
nand UO_773 (O_773,N_19584,N_16994);
nor UO_774 (O_774,N_19251,N_15547);
nor UO_775 (O_775,N_16631,N_19341);
and UO_776 (O_776,N_17909,N_18130);
nor UO_777 (O_777,N_19020,N_18324);
nor UO_778 (O_778,N_19037,N_18570);
xor UO_779 (O_779,N_19625,N_17330);
xor UO_780 (O_780,N_17608,N_15111);
nand UO_781 (O_781,N_18736,N_17831);
or UO_782 (O_782,N_18989,N_18512);
or UO_783 (O_783,N_16678,N_15247);
xnor UO_784 (O_784,N_18897,N_18258);
nor UO_785 (O_785,N_17751,N_15391);
xor UO_786 (O_786,N_16412,N_16806);
nor UO_787 (O_787,N_17398,N_19573);
nand UO_788 (O_788,N_18724,N_15025);
nor UO_789 (O_789,N_15906,N_17234);
nor UO_790 (O_790,N_18693,N_15305);
and UO_791 (O_791,N_17572,N_15957);
or UO_792 (O_792,N_16243,N_15590);
nor UO_793 (O_793,N_16071,N_15459);
nand UO_794 (O_794,N_17254,N_17448);
nand UO_795 (O_795,N_19644,N_15281);
xor UO_796 (O_796,N_17480,N_18651);
xnor UO_797 (O_797,N_17355,N_17058);
xor UO_798 (O_798,N_17976,N_19606);
and UO_799 (O_799,N_16937,N_15758);
and UO_800 (O_800,N_17553,N_16682);
xor UO_801 (O_801,N_17625,N_19446);
or UO_802 (O_802,N_18965,N_19563);
xnor UO_803 (O_803,N_17379,N_18773);
xnor UO_804 (O_804,N_17986,N_18543);
nor UO_805 (O_805,N_16865,N_16655);
xor UO_806 (O_806,N_15651,N_18595);
nor UO_807 (O_807,N_18432,N_18657);
nand UO_808 (O_808,N_18374,N_16947);
or UO_809 (O_809,N_15617,N_17246);
and UO_810 (O_810,N_19436,N_19555);
or UO_811 (O_811,N_15807,N_18781);
and UO_812 (O_812,N_16781,N_19293);
and UO_813 (O_813,N_15895,N_15994);
or UO_814 (O_814,N_16586,N_15907);
or UO_815 (O_815,N_19476,N_19972);
nor UO_816 (O_816,N_19146,N_15240);
nand UO_817 (O_817,N_17792,N_19299);
xnor UO_818 (O_818,N_19072,N_15398);
nor UO_819 (O_819,N_18772,N_16401);
or UO_820 (O_820,N_15962,N_18628);
nor UO_821 (O_821,N_16112,N_17833);
or UO_822 (O_822,N_15533,N_19977);
xnor UO_823 (O_823,N_15039,N_15772);
nor UO_824 (O_824,N_19520,N_19069);
nand UO_825 (O_825,N_17816,N_19831);
or UO_826 (O_826,N_16605,N_17399);
xor UO_827 (O_827,N_15390,N_19613);
and UO_828 (O_828,N_18808,N_16046);
and UO_829 (O_829,N_16183,N_18372);
or UO_830 (O_830,N_19525,N_18511);
xor UO_831 (O_831,N_16424,N_19702);
nor UO_832 (O_832,N_18355,N_18200);
xor UO_833 (O_833,N_16974,N_18079);
nor UO_834 (O_834,N_15442,N_18078);
or UO_835 (O_835,N_16612,N_16283);
and UO_836 (O_836,N_15559,N_17693);
nor UO_837 (O_837,N_15258,N_18462);
xnor UO_838 (O_838,N_19647,N_16003);
and UO_839 (O_839,N_15678,N_18503);
xnor UO_840 (O_840,N_17201,N_18069);
and UO_841 (O_841,N_15625,N_15679);
xor UO_842 (O_842,N_18632,N_15154);
xor UO_843 (O_843,N_15513,N_17675);
or UO_844 (O_844,N_15761,N_15497);
xnor UO_845 (O_845,N_17899,N_19941);
nor UO_846 (O_846,N_19939,N_18435);
and UO_847 (O_847,N_18487,N_16139);
and UO_848 (O_848,N_15861,N_16237);
and UO_849 (O_849,N_18727,N_19712);
xor UO_850 (O_850,N_18883,N_18248);
nand UO_851 (O_851,N_19426,N_17580);
and UO_852 (O_852,N_15958,N_15188);
xor UO_853 (O_853,N_19348,N_15723);
or UO_854 (O_854,N_15632,N_17999);
nand UO_855 (O_855,N_17688,N_15809);
nor UO_856 (O_856,N_17512,N_19783);
nand UO_857 (O_857,N_18331,N_17049);
nand UO_858 (O_858,N_16518,N_19292);
xor UO_859 (O_859,N_17260,N_16919);
nor UO_860 (O_860,N_19894,N_16984);
or UO_861 (O_861,N_18747,N_17011);
nand UO_862 (O_862,N_17825,N_16347);
nor UO_863 (O_863,N_17173,N_19084);
xor UO_864 (O_864,N_15713,N_18219);
and UO_865 (O_865,N_18951,N_15489);
nor UO_866 (O_866,N_15219,N_18348);
nand UO_867 (O_867,N_19026,N_16680);
xor UO_868 (O_868,N_16199,N_16166);
and UO_869 (O_869,N_16621,N_18587);
and UO_870 (O_870,N_15584,N_15739);
xnor UO_871 (O_871,N_17650,N_19787);
and UO_872 (O_872,N_15647,N_18967);
xor UO_873 (O_873,N_19044,N_19284);
nand UO_874 (O_874,N_15770,N_16761);
and UO_875 (O_875,N_19278,N_17029);
nand UO_876 (O_876,N_18088,N_19112);
or UO_877 (O_877,N_17702,N_16585);
or UO_878 (O_878,N_17228,N_18832);
nand UO_879 (O_879,N_18685,N_19685);
or UO_880 (O_880,N_19900,N_17236);
nand UO_881 (O_881,N_17433,N_19591);
nor UO_882 (O_882,N_16565,N_19259);
and UO_883 (O_883,N_18729,N_17942);
xnor UO_884 (O_884,N_15376,N_19539);
xnor UO_885 (O_885,N_15351,N_15000);
and UO_886 (O_886,N_18450,N_19834);
nor UO_887 (O_887,N_17256,N_15628);
xor UO_888 (O_888,N_15333,N_16168);
nand UO_889 (O_889,N_19888,N_15745);
nand UO_890 (O_890,N_16576,N_15701);
nor UO_891 (O_891,N_18660,N_17350);
xnor UO_892 (O_892,N_19746,N_16127);
and UO_893 (O_893,N_15794,N_16294);
xor UO_894 (O_894,N_15300,N_18980);
and UO_895 (O_895,N_15618,N_16951);
or UO_896 (O_896,N_19885,N_18403);
xor UO_897 (O_897,N_15774,N_17613);
xnor UO_898 (O_898,N_18393,N_18766);
or UO_899 (O_899,N_18938,N_15017);
nor UO_900 (O_900,N_15175,N_19854);
xnor UO_901 (O_901,N_19740,N_18870);
xnor UO_902 (O_902,N_16099,N_15796);
or UO_903 (O_903,N_18819,N_16101);
or UO_904 (O_904,N_15334,N_17488);
or UO_905 (O_905,N_16089,N_19987);
nor UO_906 (O_906,N_19884,N_15805);
or UO_907 (O_907,N_16027,N_15759);
or UO_908 (O_908,N_17122,N_19003);
nor UO_909 (O_909,N_18152,N_18645);
or UO_910 (O_910,N_18847,N_15905);
nand UO_911 (O_911,N_18402,N_15848);
and UO_912 (O_912,N_18341,N_19123);
or UO_913 (O_913,N_15429,N_18087);
or UO_914 (O_914,N_18827,N_19132);
or UO_915 (O_915,N_15242,N_17658);
xnor UO_916 (O_916,N_17048,N_19280);
nor UO_917 (O_917,N_15817,N_18100);
or UO_918 (O_918,N_15568,N_18271);
or UO_919 (O_919,N_19260,N_17780);
and UO_920 (O_920,N_17360,N_19677);
nand UO_921 (O_921,N_15612,N_18800);
nor UO_922 (O_922,N_17781,N_16753);
or UO_923 (O_923,N_17098,N_17391);
nor UO_924 (O_924,N_17279,N_15697);
nor UO_925 (O_925,N_15552,N_19237);
nor UO_926 (O_926,N_15786,N_17985);
nand UO_927 (O_927,N_15885,N_15255);
nor UO_928 (O_928,N_16857,N_19395);
nor UO_929 (O_929,N_19492,N_18676);
nand UO_930 (O_930,N_16816,N_17598);
xor UO_931 (O_931,N_15945,N_17696);
xnor UO_932 (O_932,N_15586,N_16953);
nor UO_933 (O_933,N_18817,N_15604);
nor UO_934 (O_934,N_15737,N_15036);
and UO_935 (O_935,N_19128,N_19254);
and UO_936 (O_936,N_15748,N_18187);
and UO_937 (O_937,N_16334,N_19451);
xor UO_938 (O_938,N_15902,N_16429);
xnor UO_939 (O_939,N_17990,N_17139);
or UO_940 (O_940,N_18909,N_17806);
xor UO_941 (O_941,N_18534,N_18853);
or UO_942 (O_942,N_18338,N_17024);
nor UO_943 (O_943,N_17496,N_17454);
and UO_944 (O_944,N_18939,N_15655);
xnor UO_945 (O_945,N_18617,N_19416);
xor UO_946 (O_946,N_19486,N_17271);
or UO_947 (O_947,N_15311,N_16824);
nor UO_948 (O_948,N_15579,N_16679);
or UO_949 (O_949,N_18583,N_15457);
xor UO_950 (O_950,N_18721,N_15797);
nor UO_951 (O_951,N_17602,N_15367);
nand UO_952 (O_952,N_17659,N_17383);
or UO_953 (O_953,N_18910,N_17295);
and UO_954 (O_954,N_15224,N_17171);
and UO_955 (O_955,N_19272,N_15518);
nor UO_956 (O_956,N_15990,N_15955);
nand UO_957 (O_957,N_18785,N_18024);
and UO_958 (O_958,N_17617,N_15908);
nand UO_959 (O_959,N_19307,N_19533);
and UO_960 (O_960,N_17680,N_16105);
xnor UO_961 (O_961,N_15925,N_17241);
nand UO_962 (O_962,N_17288,N_19161);
nor UO_963 (O_963,N_19018,N_19212);
nand UO_964 (O_964,N_19096,N_15422);
and UO_965 (O_965,N_16043,N_16650);
nand UO_966 (O_966,N_15539,N_19773);
nor UO_967 (O_967,N_17935,N_18559);
xnor UO_968 (O_968,N_15929,N_17844);
nand UO_969 (O_969,N_18670,N_15393);
nand UO_970 (O_970,N_15325,N_17717);
or UO_971 (O_971,N_18658,N_18860);
nor UO_972 (O_972,N_19014,N_17929);
or UO_973 (O_973,N_15751,N_19593);
nand UO_974 (O_974,N_19226,N_18960);
nor UO_975 (O_975,N_18564,N_15594);
and UO_976 (O_976,N_15519,N_19954);
and UO_977 (O_977,N_18982,N_18973);
nand UO_978 (O_978,N_15076,N_18449);
nor UO_979 (O_979,N_18900,N_19063);
and UO_980 (O_980,N_18031,N_19389);
or UO_981 (O_981,N_18422,N_17134);
nor UO_982 (O_982,N_16982,N_16792);
nand UO_983 (O_983,N_19016,N_19127);
nor UO_984 (O_984,N_19635,N_16988);
and UO_985 (O_985,N_18149,N_18957);
and UO_986 (O_986,N_19496,N_17627);
xnor UO_987 (O_987,N_18437,N_17697);
nor UO_988 (O_988,N_19962,N_18056);
nand UO_989 (O_989,N_19698,N_18904);
nand UO_990 (O_990,N_16863,N_18770);
or UO_991 (O_991,N_16779,N_18307);
xnor UO_992 (O_992,N_15645,N_16815);
xnor UO_993 (O_993,N_16796,N_17129);
nand UO_994 (O_994,N_16205,N_15515);
xor UO_995 (O_995,N_17206,N_17489);
or UO_996 (O_996,N_18359,N_19428);
or UO_997 (O_997,N_16477,N_17891);
nand UO_998 (O_998,N_17783,N_15854);
or UO_999 (O_999,N_19524,N_18743);
or UO_1000 (O_1000,N_18858,N_18268);
nor UO_1001 (O_1001,N_16916,N_18905);
and UO_1002 (O_1002,N_15792,N_19781);
nor UO_1003 (O_1003,N_16791,N_16024);
or UO_1004 (O_1004,N_16297,N_16235);
xnor UO_1005 (O_1005,N_15606,N_17715);
nand UO_1006 (O_1006,N_16820,N_15487);
xor UO_1007 (O_1007,N_16760,N_18004);
xor UO_1008 (O_1008,N_17681,N_19385);
nand UO_1009 (O_1009,N_15397,N_15762);
xnor UO_1010 (O_1010,N_18186,N_19899);
or UO_1011 (O_1011,N_17147,N_15793);
xnor UO_1012 (O_1012,N_17161,N_15609);
nand UO_1013 (O_1013,N_17778,N_15095);
nand UO_1014 (O_1014,N_17632,N_17815);
xor UO_1015 (O_1015,N_16948,N_19499);
and UO_1016 (O_1016,N_19882,N_18032);
xnor UO_1017 (O_1017,N_16379,N_16363);
xnor UO_1018 (O_1018,N_15296,N_19222);
and UO_1019 (O_1019,N_15093,N_16546);
or UO_1020 (O_1020,N_15850,N_18732);
xnor UO_1021 (O_1021,N_19349,N_16582);
xor UO_1022 (O_1022,N_16055,N_19369);
xor UO_1023 (O_1023,N_15654,N_15784);
nor UO_1024 (O_1024,N_16754,N_17713);
nand UO_1025 (O_1025,N_15517,N_16925);
and UO_1026 (O_1026,N_15545,N_19110);
nor UO_1027 (O_1027,N_16187,N_16748);
or UO_1028 (O_1028,N_19507,N_19043);
nand UO_1029 (O_1029,N_19652,N_16522);
nand UO_1030 (O_1030,N_16635,N_15587);
and UO_1031 (O_1031,N_15749,N_18533);
or UO_1032 (O_1032,N_17964,N_15061);
nand UO_1033 (O_1033,N_18020,N_19046);
nand UO_1034 (O_1034,N_18317,N_16482);
and UO_1035 (O_1035,N_16282,N_18080);
nor UO_1036 (O_1036,N_16269,N_18241);
and UO_1037 (O_1037,N_18481,N_19202);
xnor UO_1038 (O_1038,N_19663,N_19456);
nand UO_1039 (O_1039,N_17652,N_19365);
or UO_1040 (O_1040,N_19856,N_18026);
nand UO_1041 (O_1041,N_18336,N_19434);
nor UO_1042 (O_1042,N_17835,N_19310);
and UO_1043 (O_1043,N_16852,N_18830);
nand UO_1044 (O_1044,N_16960,N_15081);
xnor UO_1045 (O_1045,N_19731,N_17876);
xor UO_1046 (O_1046,N_18593,N_16644);
and UO_1047 (O_1047,N_15810,N_17137);
or UO_1048 (O_1048,N_19177,N_16714);
nand UO_1049 (O_1049,N_16441,N_15754);
nor UO_1050 (O_1050,N_16377,N_19546);
nand UO_1051 (O_1051,N_15374,N_16498);
nand UO_1052 (O_1052,N_15607,N_16751);
or UO_1053 (O_1053,N_15933,N_17819);
and UO_1054 (O_1054,N_19017,N_18826);
xor UO_1055 (O_1055,N_17823,N_18948);
nand UO_1056 (O_1056,N_19891,N_15495);
nor UO_1057 (O_1057,N_15349,N_18539);
xnor UO_1058 (O_1058,N_19317,N_16039);
and UO_1059 (O_1059,N_16689,N_15985);
xor UO_1060 (O_1060,N_18500,N_16410);
and UO_1061 (O_1061,N_18039,N_19775);
nand UO_1062 (O_1062,N_15953,N_18335);
and UO_1063 (O_1063,N_17708,N_16613);
xor UO_1064 (O_1064,N_18406,N_18120);
and UO_1065 (O_1065,N_19109,N_17760);
and UO_1066 (O_1066,N_19425,N_19442);
xor UO_1067 (O_1067,N_19135,N_18546);
nand UO_1068 (O_1068,N_15534,N_17040);
nor UO_1069 (O_1069,N_16308,N_15405);
nor UO_1070 (O_1070,N_19287,N_19431);
and UO_1071 (O_1071,N_17120,N_16221);
nand UO_1072 (O_1072,N_15042,N_15016);
nand UO_1073 (O_1073,N_15879,N_17442);
xnor UO_1074 (O_1074,N_18469,N_16923);
and UO_1075 (O_1075,N_17801,N_19769);
nor UO_1076 (O_1076,N_15970,N_18722);
xor UO_1077 (O_1077,N_15622,N_18176);
nor UO_1078 (O_1078,N_18945,N_18728);
or UO_1079 (O_1079,N_15750,N_19541);
nor UO_1080 (O_1080,N_19378,N_19419);
and UO_1081 (O_1081,N_16059,N_17560);
or UO_1082 (O_1082,N_16271,N_18873);
xnor UO_1083 (O_1083,N_15602,N_16976);
xor UO_1084 (O_1084,N_19203,N_18638);
nand UO_1085 (O_1085,N_15238,N_19662);
or UO_1086 (O_1086,N_18168,N_18291);
or UO_1087 (O_1087,N_16874,N_17537);
xnor UO_1088 (O_1088,N_16317,N_17192);
or UO_1089 (O_1089,N_15881,N_19806);
nor UO_1090 (O_1090,N_16704,N_17977);
and UO_1091 (O_1091,N_18189,N_17053);
or UO_1092 (O_1092,N_19994,N_19588);
nand UO_1093 (O_1093,N_16388,N_18240);
xor UO_1094 (O_1094,N_19965,N_19534);
xor UO_1095 (O_1095,N_18833,N_16797);
nor UO_1096 (O_1096,N_18028,N_17515);
or UO_1097 (O_1097,N_18840,N_18809);
or UO_1098 (O_1098,N_17292,N_16548);
nor UO_1099 (O_1099,N_16686,N_15856);
xnor UO_1100 (O_1100,N_15345,N_16943);
or UO_1101 (O_1101,N_15149,N_19683);
nand UO_1102 (O_1102,N_15234,N_18627);
nand UO_1103 (O_1103,N_15150,N_16611);
or UO_1104 (O_1104,N_18086,N_15567);
nor UO_1105 (O_1105,N_15988,N_19409);
and UO_1106 (O_1106,N_17563,N_17138);
or UO_1107 (O_1107,N_15139,N_19579);
nand UO_1108 (O_1108,N_19895,N_17195);
xnor UO_1109 (O_1109,N_16591,N_16287);
or UO_1110 (O_1110,N_17547,N_15914);
nand UO_1111 (O_1111,N_17199,N_18825);
and UO_1112 (O_1112,N_15913,N_19167);
xnor UO_1113 (O_1113,N_18303,N_15200);
nand UO_1114 (O_1114,N_15276,N_16457);
nand UO_1115 (O_1115,N_16601,N_15965);
nor UO_1116 (O_1116,N_16073,N_18019);
or UO_1117 (O_1117,N_19485,N_18412);
xnor UO_1118 (O_1118,N_17827,N_16872);
and UO_1119 (O_1119,N_18389,N_17103);
and UO_1120 (O_1120,N_17465,N_15098);
or UO_1121 (O_1121,N_18751,N_17499);
and UO_1122 (O_1122,N_19242,N_19622);
or UO_1123 (O_1123,N_16763,N_15162);
xnor UO_1124 (O_1124,N_15273,N_19850);
and UO_1125 (O_1125,N_16231,N_18616);
xor UO_1126 (O_1126,N_16227,N_17843);
and UO_1127 (O_1127,N_18185,N_19001);
or UO_1128 (O_1128,N_15728,N_15551);
and UO_1129 (O_1129,N_17877,N_17859);
xor UO_1130 (O_1130,N_17002,N_19498);
nand UO_1131 (O_1131,N_15235,N_15571);
and UO_1132 (O_1132,N_18744,N_17264);
nand UO_1133 (O_1133,N_19138,N_18509);
nand UO_1134 (O_1134,N_19630,N_18581);
nand UO_1135 (O_1135,N_15174,N_19083);
and UO_1136 (O_1136,N_16146,N_19199);
or UO_1137 (O_1137,N_16563,N_19006);
or UO_1138 (O_1138,N_19355,N_16596);
nand UO_1139 (O_1139,N_16489,N_15605);
and UO_1140 (O_1140,N_19086,N_15502);
nand UO_1141 (O_1141,N_19508,N_15335);
nand UO_1142 (O_1142,N_15639,N_16568);
nand UO_1143 (O_1143,N_19841,N_19282);
nor UO_1144 (O_1144,N_18886,N_16192);
nand UO_1145 (O_1145,N_18669,N_15146);
and UO_1146 (O_1146,N_17518,N_15252);
xor UO_1147 (O_1147,N_17232,N_17663);
xor UO_1148 (O_1148,N_15742,N_19518);
xor UO_1149 (O_1149,N_18109,N_19249);
or UO_1150 (O_1150,N_19009,N_18573);
or UO_1151 (O_1151,N_17072,N_19950);
or UO_1152 (O_1152,N_18175,N_19459);
nor UO_1153 (O_1153,N_16408,N_16466);
nor UO_1154 (O_1154,N_17748,N_16239);
nor UO_1155 (O_1155,N_19505,N_19753);
or UO_1156 (O_1156,N_18764,N_18454);
nand UO_1157 (O_1157,N_17721,N_16065);
and UO_1158 (O_1158,N_15833,N_16964);
or UO_1159 (O_1159,N_16935,N_18464);
and UO_1160 (O_1160,N_18941,N_19610);
xor UO_1161 (O_1161,N_17900,N_15847);
and UO_1162 (O_1162,N_16258,N_15940);
nor UO_1163 (O_1163,N_15695,N_18375);
or UO_1164 (O_1164,N_17003,N_15714);
xor UO_1165 (O_1165,N_17588,N_19129);
xor UO_1166 (O_1166,N_15413,N_19209);
and UO_1167 (O_1167,N_18139,N_15173);
or UO_1168 (O_1168,N_18818,N_16405);
nor UO_1169 (O_1169,N_16774,N_16841);
xor UO_1170 (O_1170,N_19246,N_17432);
nand UO_1171 (O_1171,N_19875,N_15034);
nor UO_1172 (O_1172,N_17111,N_16671);
nand UO_1173 (O_1173,N_16056,N_19966);
nor UO_1174 (O_1174,N_19796,N_15932);
nor UO_1175 (O_1175,N_18405,N_18029);
or UO_1176 (O_1176,N_19980,N_15488);
or UO_1177 (O_1177,N_19056,N_18280);
and UO_1178 (O_1178,N_19062,N_19696);
nand UO_1179 (O_1179,N_16854,N_15195);
xor UO_1180 (O_1180,N_15373,N_19396);
nor UO_1181 (O_1181,N_16058,N_18929);
nand UO_1182 (O_1182,N_16499,N_15250);
nand UO_1183 (O_1183,N_16367,N_17101);
nor UO_1184 (O_1184,N_15055,N_19502);
nand UO_1185 (O_1185,N_18922,N_18778);
and UO_1186 (O_1186,N_19824,N_15049);
nor UO_1187 (O_1187,N_18133,N_18548);
or UO_1188 (O_1188,N_16959,N_17880);
or UO_1189 (O_1189,N_16240,N_19750);
nor UO_1190 (O_1190,N_17678,N_15505);
xnor UO_1191 (O_1191,N_18443,N_17959);
xnor UO_1192 (O_1192,N_16583,N_16569);
or UO_1193 (O_1193,N_18674,N_16454);
nor UO_1194 (O_1194,N_15170,N_16741);
nand UO_1195 (O_1195,N_17051,N_16933);
nor UO_1196 (O_1196,N_17293,N_17621);
or UO_1197 (O_1197,N_18306,N_18410);
and UO_1198 (O_1198,N_19861,N_15918);
or UO_1199 (O_1199,N_16507,N_16314);
or UO_1200 (O_1200,N_15312,N_16031);
and UO_1201 (O_1201,N_15033,N_18578);
nand UO_1202 (O_1202,N_17186,N_16830);
xor UO_1203 (O_1203,N_18748,N_16990);
xnor UO_1204 (O_1204,N_19829,N_19394);
or UO_1205 (O_1205,N_17957,N_17500);
xnor UO_1206 (O_1206,N_16619,N_17692);
xnor UO_1207 (O_1207,N_16757,N_18424);
and UO_1208 (O_1208,N_17626,N_19937);
nand UO_1209 (O_1209,N_17962,N_17540);
or UO_1210 (O_1210,N_15791,N_18299);
or UO_1211 (O_1211,N_16888,N_15143);
and UO_1212 (O_1212,N_17016,N_16706);
xnor UO_1213 (O_1213,N_18527,N_16823);
xor UO_1214 (O_1214,N_18691,N_19047);
and UO_1215 (O_1215,N_17981,N_17854);
or UO_1216 (O_1216,N_15656,N_18992);
nor UO_1217 (O_1217,N_16663,N_19719);
nand UO_1218 (O_1218,N_18786,N_18071);
or UO_1219 (O_1219,N_18673,N_19022);
xor UO_1220 (O_1220,N_18273,N_15436);
and UO_1221 (O_1221,N_19449,N_16444);
or UO_1222 (O_1222,N_17333,N_15826);
and UO_1223 (O_1223,N_17390,N_18597);
or UO_1224 (O_1224,N_16851,N_16337);
and UO_1225 (O_1225,N_16439,N_18214);
nand UO_1226 (O_1226,N_17925,N_17498);
nand UO_1227 (O_1227,N_19333,N_18446);
nand UO_1228 (O_1228,N_16467,N_15920);
xnor UO_1229 (O_1229,N_19300,N_18266);
and UO_1230 (O_1230,N_16900,N_18571);
and UO_1231 (O_1231,N_18699,N_17782);
nor UO_1232 (O_1232,N_16209,N_15285);
and UO_1233 (O_1233,N_19473,N_18695);
and UO_1234 (O_1234,N_17898,N_15657);
xnor UO_1235 (O_1235,N_16398,N_17324);
nand UO_1236 (O_1236,N_19709,N_17229);
nand UO_1237 (O_1237,N_19193,N_18178);
nand UO_1238 (O_1238,N_15818,N_16450);
nor UO_1239 (O_1239,N_18245,N_16324);
xor UO_1240 (O_1240,N_17249,N_16066);
or UO_1241 (O_1241,N_17852,N_18844);
and UO_1242 (O_1242,N_19565,N_19092);
nor UO_1243 (O_1243,N_18385,N_17582);
or UO_1244 (O_1244,N_17378,N_16161);
nand UO_1245 (O_1245,N_17400,N_18547);
or UO_1246 (O_1246,N_15507,N_18887);
nand UO_1247 (O_1247,N_16812,N_16912);
and UO_1248 (O_1248,N_19158,N_15189);
or UO_1249 (O_1249,N_16111,N_18739);
or UO_1250 (O_1250,N_19779,N_16285);
nor UO_1251 (O_1251,N_18612,N_19830);
nand UO_1252 (O_1252,N_16246,N_18151);
nand UO_1253 (O_1253,N_15385,N_16188);
nand UO_1254 (O_1254,N_15096,N_16907);
and UO_1255 (O_1255,N_19705,N_17010);
and UO_1256 (O_1256,N_17797,N_19271);
nor UO_1257 (O_1257,N_17178,N_19522);
and UO_1258 (O_1258,N_15211,N_16834);
nand UO_1259 (O_1259,N_17619,N_18767);
and UO_1260 (O_1260,N_17176,N_16384);
xor UO_1261 (O_1261,N_18114,N_19319);
or UO_1262 (O_1262,N_18407,N_15492);
and UO_1263 (O_1263,N_16033,N_19922);
nand UO_1264 (O_1264,N_15435,N_16358);
or UO_1265 (O_1265,N_16219,N_16773);
and UO_1266 (O_1266,N_18899,N_18343);
nand UO_1267 (O_1267,N_17528,N_18377);
and UO_1268 (O_1268,N_16969,N_17297);
nand UO_1269 (O_1269,N_15780,N_15471);
nor UO_1270 (O_1270,N_15694,N_16343);
xnor UO_1271 (O_1271,N_16291,N_15108);
nor UO_1272 (O_1272,N_17892,N_15185);
nor UO_1273 (O_1273,N_15968,N_17743);
and UO_1274 (O_1274,N_16230,N_18391);
nand UO_1275 (O_1275,N_16312,N_18551);
xnor UO_1276 (O_1276,N_15512,N_15212);
or UO_1277 (O_1277,N_15468,N_18969);
nand UO_1278 (O_1278,N_15105,N_19866);
and UO_1279 (O_1279,N_15331,N_19963);
or UO_1280 (O_1280,N_15693,N_17523);
nor UO_1281 (O_1281,N_19019,N_16875);
or UO_1282 (O_1282,N_18972,N_19100);
nor UO_1283 (O_1283,N_17311,N_19870);
and UO_1284 (O_1284,N_18565,N_17338);
xor UO_1285 (O_1285,N_17824,N_18925);
and UO_1286 (O_1286,N_17376,N_18712);
or UO_1287 (O_1287,N_16799,N_17903);
nor UO_1288 (O_1288,N_16106,N_17266);
nand UO_1289 (O_1289,N_17853,N_18436);
or UO_1290 (O_1290,N_19550,N_18733);
nor UO_1291 (O_1291,N_17726,N_15043);
or UO_1292 (O_1292,N_16817,N_16064);
nor UO_1293 (O_1293,N_15665,N_17032);
nand UO_1294 (O_1294,N_19154,N_15516);
and UO_1295 (O_1295,N_16313,N_19405);
xor UO_1296 (O_1296,N_19747,N_18249);
nor UO_1297 (O_1297,N_16254,N_19924);
nand UO_1298 (O_1298,N_18686,N_18801);
and UO_1299 (O_1299,N_15243,N_17932);
nand UO_1300 (O_1300,N_19211,N_15417);
xor UO_1301 (O_1301,N_15117,N_15677);
nand UO_1302 (O_1302,N_19594,N_15291);
or UO_1303 (O_1303,N_17423,N_18304);
nor UO_1304 (O_1304,N_17533,N_17575);
xnor UO_1305 (O_1305,N_17566,N_15408);
nand UO_1306 (O_1306,N_17549,N_19455);
xor UO_1307 (O_1307,N_15501,N_19816);
and UO_1308 (O_1308,N_16629,N_15862);
nand UO_1309 (O_1309,N_18971,N_17538);
nand UO_1310 (O_1310,N_19981,N_15503);
xnor UO_1311 (O_1311,N_17467,N_16890);
xor UO_1312 (O_1312,N_17340,N_18289);
and UO_1313 (O_1313,N_18618,N_18188);
xnor UO_1314 (O_1314,N_15934,N_19568);
or UO_1315 (O_1315,N_18124,N_17920);
nor UO_1316 (O_1316,N_15129,N_15051);
and UO_1317 (O_1317,N_17766,N_15007);
or UO_1318 (O_1318,N_19767,N_16625);
or UO_1319 (O_1319,N_15763,N_19815);
xnor UO_1320 (O_1320,N_16117,N_16962);
or UO_1321 (O_1321,N_16177,N_15338);
or UO_1322 (O_1322,N_19152,N_18150);
xnor UO_1323 (O_1323,N_15127,N_16290);
nor UO_1324 (O_1324,N_17045,N_18089);
nand UO_1325 (O_1325,N_19552,N_17267);
nand UO_1326 (O_1326,N_17200,N_16627);
nand UO_1327 (O_1327,N_19483,N_15734);
or UO_1328 (O_1328,N_18894,N_17604);
xor UO_1329 (O_1329,N_19744,N_15894);
nand UO_1330 (O_1330,N_19754,N_19908);
and UO_1331 (O_1331,N_17737,N_18269);
nor UO_1332 (O_1332,N_19811,N_18737);
xor UO_1333 (O_1333,N_19340,N_17076);
or UO_1334 (O_1334,N_18353,N_18165);
nand UO_1335 (O_1335,N_15215,N_19437);
xnor UO_1336 (O_1336,N_19356,N_16626);
xor UO_1337 (O_1337,N_16270,N_18195);
xor UO_1338 (O_1338,N_18966,N_18298);
xnor UO_1339 (O_1339,N_16116,N_16190);
and UO_1340 (O_1340,N_15259,N_16197);
or UO_1341 (O_1341,N_19328,N_19184);
nor UO_1342 (O_1342,N_15272,N_15901);
xnor UO_1343 (O_1343,N_15186,N_15718);
nand UO_1344 (O_1344,N_18208,N_17214);
nand UO_1345 (O_1345,N_15052,N_17150);
nand UO_1346 (O_1346,N_17299,N_18856);
and UO_1347 (O_1347,N_15578,N_19749);
nand UO_1348 (O_1348,N_16639,N_17462);
xor UO_1349 (O_1349,N_15470,N_19401);
xor UO_1350 (O_1350,N_15118,N_16204);
xor UO_1351 (O_1351,N_16208,N_17960);
nor UO_1352 (O_1352,N_18639,N_16836);
nor UO_1353 (O_1353,N_15307,N_17036);
nand UO_1354 (O_1354,N_16740,N_16130);
or UO_1355 (O_1355,N_17474,N_18048);
or UO_1356 (O_1356,N_15846,N_19989);
and UO_1357 (O_1357,N_17084,N_19329);
and UO_1358 (O_1358,N_15776,N_19490);
nor UO_1359 (O_1359,N_19388,N_19848);
nor UO_1360 (O_1360,N_18725,N_16705);
nor UO_1361 (O_1361,N_15681,N_16995);
and UO_1362 (O_1362,N_16486,N_19993);
or UO_1363 (O_1363,N_16739,N_18720);
nor UO_1364 (O_1364,N_16272,N_16098);
or UO_1365 (O_1365,N_17606,N_19559);
or UO_1366 (O_1366,N_17479,N_19718);
xnor UO_1367 (O_1367,N_19795,N_16849);
nand UO_1368 (O_1368,N_19845,N_18552);
xnor UO_1369 (O_1369,N_16802,N_16949);
or UO_1370 (O_1370,N_19786,N_19327);
xnor UO_1371 (O_1371,N_15365,N_16495);
and UO_1372 (O_1372,N_17494,N_15368);
xnor UO_1373 (O_1373,N_17329,N_17250);
and UO_1374 (O_1374,N_15330,N_16826);
nor UO_1375 (O_1375,N_19628,N_19036);
nor UO_1376 (O_1376,N_18400,N_19085);
nand UO_1377 (O_1377,N_19896,N_15771);
or UO_1378 (O_1378,N_19241,N_19643);
nand UO_1379 (O_1379,N_15090,N_18180);
nor UO_1380 (O_1380,N_18682,N_17447);
or UO_1381 (O_1381,N_15952,N_16307);
xor UO_1382 (O_1382,N_17439,N_17727);
or UO_1383 (O_1383,N_18814,N_18979);
and UO_1384 (O_1384,N_18810,N_16861);
or UO_1385 (O_1385,N_19743,N_15863);
or UO_1386 (O_1386,N_17611,N_18354);
or UO_1387 (O_1387,N_16897,N_19590);
xnor UO_1388 (O_1388,N_19457,N_15395);
nand UO_1389 (O_1389,N_17809,N_16549);
or UO_1390 (O_1390,N_19470,N_17531);
xor UO_1391 (O_1391,N_17583,N_17939);
xnor UO_1392 (O_1392,N_15220,N_18932);
nor UO_1393 (O_1393,N_19760,N_15210);
nand UO_1394 (O_1394,N_16504,N_17581);
nand UO_1395 (O_1395,N_16138,N_15553);
xnor UO_1396 (O_1396,N_16030,N_15841);
and UO_1397 (O_1397,N_19450,N_18014);
or UO_1398 (O_1398,N_17418,N_19717);
xnor UO_1399 (O_1399,N_17238,N_15249);
nand UO_1400 (O_1400,N_16599,N_16345);
nor UO_1401 (O_1401,N_16217,N_16136);
nand UO_1402 (O_1402,N_17701,N_18494);
nor UO_1403 (O_1403,N_16311,N_17151);
xor UO_1404 (O_1404,N_18099,N_19477);
nand UO_1405 (O_1405,N_15631,N_16260);
nor UO_1406 (O_1406,N_16967,N_19971);
xor UO_1407 (O_1407,N_18831,N_19595);
nand UO_1408 (O_1408,N_16480,N_17483);
and UO_1409 (O_1409,N_19690,N_19218);
nor UO_1410 (O_1410,N_19575,N_15580);
xnor UO_1411 (O_1411,N_16615,N_15142);
and UO_1412 (O_1412,N_18036,N_17594);
and UO_1413 (O_1413,N_16357,N_17974);
nand UO_1414 (O_1414,N_19912,N_16051);
nor UO_1415 (O_1415,N_17955,N_19689);
or UO_1416 (O_1416,N_19617,N_18137);
nor UO_1417 (O_1417,N_17954,N_16289);
and UO_1418 (O_1418,N_18401,N_19646);
nand UO_1419 (O_1419,N_17654,N_17438);
nor UO_1420 (O_1420,N_16034,N_16284);
nand UO_1421 (O_1421,N_17106,N_19136);
xor UO_1422 (O_1422,N_17273,N_19614);
or UO_1423 (O_1423,N_17864,N_18872);
and UO_1424 (O_1424,N_16319,N_16610);
or UO_1425 (O_1425,N_16945,N_16931);
xor UO_1426 (O_1426,N_18874,N_15803);
or UO_1427 (O_1427,N_18921,N_19631);
or UO_1428 (O_1428,N_18919,N_18771);
nor UO_1429 (O_1429,N_16860,N_15823);
and UO_1430 (O_1430,N_16886,N_19808);
or UO_1431 (O_1431,N_15446,N_17289);
or UO_1432 (O_1432,N_16532,N_19506);
or UO_1433 (O_1433,N_15904,N_18763);
or UO_1434 (O_1434,N_19782,N_16137);
nand UO_1435 (O_1435,N_18997,N_15416);
nand UO_1436 (O_1436,N_18940,N_18318);
nand UO_1437 (O_1437,N_15752,N_16255);
and UO_1438 (O_1438,N_17290,N_18495);
and UO_1439 (O_1439,N_18305,N_15884);
nand UO_1440 (O_1440,N_19669,N_16570);
nand UO_1441 (O_1441,N_16709,N_19151);
nand UO_1442 (O_1442,N_15388,N_16885);
nor UO_1443 (O_1443,N_19545,N_17352);
and UO_1444 (O_1444,N_15183,N_18279);
nand UO_1445 (O_1445,N_15213,N_15528);
nand UO_1446 (O_1446,N_17037,N_16020);
nand UO_1447 (O_1447,N_16707,N_17733);
nand UO_1448 (O_1448,N_19448,N_19737);
nor UO_1449 (O_1449,N_15961,N_15806);
xnor UO_1450 (O_1450,N_15947,N_17993);
and UO_1451 (O_1451,N_19105,N_15828);
or UO_1452 (O_1452,N_15406,N_18903);
and UO_1453 (O_1453,N_18749,N_18912);
nand UO_1454 (O_1454,N_19290,N_18452);
or UO_1455 (O_1455,N_16212,N_17882);
and UO_1456 (O_1456,N_16224,N_15022);
xor UO_1457 (O_1457,N_18820,N_17629);
or UO_1458 (O_1458,N_17019,N_17174);
nor UO_1459 (O_1459,N_15744,N_15599);
nor UO_1460 (O_1460,N_16133,N_15343);
nor UO_1461 (O_1461,N_17720,N_18090);
or UO_1462 (O_1462,N_18865,N_16067);
xnor UO_1463 (O_1463,N_18119,N_16047);
nand UO_1464 (O_1464,N_18192,N_18501);
nand UO_1465 (O_1465,N_15822,N_18421);
or UO_1466 (O_1466,N_18650,N_16009);
nor UO_1467 (O_1467,N_18958,N_16768);
nor UO_1468 (O_1468,N_19039,N_16448);
xor UO_1469 (O_1469,N_15124,N_19694);
or UO_1470 (O_1470,N_17804,N_18041);
xnor UO_1471 (O_1471,N_18174,N_19521);
nor UO_1472 (O_1472,N_19607,N_17193);
nand UO_1473 (O_1473,N_19074,N_18380);
xnor UO_1474 (O_1474,N_18395,N_17225);
and UO_1475 (O_1475,N_19131,N_15432);
xnor UO_1476 (O_1476,N_19569,N_17335);
nor UO_1477 (O_1477,N_16465,N_17020);
nor UO_1478 (O_1478,N_16764,N_15638);
nor UO_1479 (O_1479,N_16641,N_15350);
or UO_1480 (O_1480,N_19960,N_19137);
and UO_1481 (O_1481,N_15467,N_16876);
nor UO_1482 (O_1482,N_18529,N_16986);
and UO_1483 (O_1483,N_19666,N_18807);
or UO_1484 (O_1484,N_17115,N_19990);
nand UO_1485 (O_1485,N_16057,N_19700);
and UO_1486 (O_1486,N_16474,N_15050);
or UO_1487 (O_1487,N_15104,N_16540);
nor UO_1488 (O_1488,N_19217,N_15767);
and UO_1489 (O_1489,N_18371,N_16194);
and UO_1490 (O_1490,N_17635,N_16002);
or UO_1491 (O_1491,N_19304,N_19862);
nor UO_1492 (O_1492,N_19418,N_19406);
and UO_1493 (O_1493,N_16008,N_15031);
nand UO_1494 (O_1494,N_15106,N_18160);
nor UO_1495 (O_1495,N_17043,N_15574);
or UO_1496 (O_1496,N_19357,N_17365);
and UO_1497 (O_1497,N_19040,N_19839);
nand UO_1498 (O_1498,N_18381,N_18296);
nand UO_1499 (O_1499,N_19691,N_17387);
and UO_1500 (O_1500,N_17773,N_19113);
nor UO_1501 (O_1501,N_16572,N_19190);
xor UO_1502 (O_1502,N_16643,N_16451);
or UO_1503 (O_1503,N_19339,N_18714);
and UO_1504 (O_1504,N_18861,N_16855);
and UO_1505 (O_1505,N_18780,N_16473);
xnor UO_1506 (O_1506,N_15708,N_16977);
nor UO_1507 (O_1507,N_16120,N_18295);
or UO_1508 (O_1508,N_15161,N_19649);
nor UO_1509 (O_1509,N_17154,N_17109);
or UO_1510 (O_1510,N_17484,N_18540);
nand UO_1511 (O_1511,N_15140,N_15363);
and UO_1512 (O_1512,N_15046,N_16535);
and UO_1513 (O_1513,N_16251,N_18138);
and UO_1514 (O_1514,N_17725,N_16460);
or UO_1515 (O_1515,N_17774,N_18614);
xor UO_1516 (O_1516,N_19076,N_17991);
nand UO_1517 (O_1517,N_19247,N_19858);
xnor UO_1518 (O_1518,N_19672,N_16004);
or UO_1519 (O_1519,N_19438,N_15460);
nor UO_1520 (O_1520,N_15067,N_19536);
nand UO_1521 (O_1521,N_18946,N_16766);
nand UO_1522 (O_1522,N_18937,N_16262);
or UO_1523 (O_1523,N_17291,N_16084);
xnor UO_1524 (O_1524,N_15558,N_16519);
or UO_1525 (O_1525,N_18278,N_19373);
nand UO_1526 (O_1526,N_19991,N_16292);
xor UO_1527 (O_1527,N_19909,N_15159);
nor UO_1528 (O_1528,N_18762,N_15072);
nand UO_1529 (O_1529,N_16309,N_18880);
or UO_1530 (O_1530,N_16373,N_16078);
nand UO_1531 (O_1531,N_19061,N_19637);
and UO_1532 (O_1532,N_16594,N_17021);
and UO_1533 (O_1533,N_17916,N_16090);
or UO_1534 (O_1534,N_16958,N_19102);
xor UO_1535 (O_1535,N_17923,N_19474);
xnor UO_1536 (O_1536,N_17091,N_15054);
nand UO_1537 (O_1537,N_19332,N_19337);
or UO_1538 (O_1538,N_19097,N_17747);
xor UO_1539 (O_1539,N_15404,N_19873);
nand UO_1540 (O_1540,N_19948,N_18205);
and UO_1541 (O_1541,N_15700,N_16382);
or UO_1542 (O_1542,N_16846,N_15875);
and UO_1543 (O_1543,N_17031,N_17092);
and UO_1544 (O_1544,N_15403,N_18859);
and UO_1545 (O_1545,N_17000,N_15197);
or UO_1546 (O_1546,N_15857,N_19111);
or UO_1547 (O_1547,N_16941,N_15614);
xnor UO_1548 (O_1548,N_15937,N_15268);
and UO_1549 (O_1549,N_15724,N_17734);
nand UO_1550 (O_1550,N_16299,N_19510);
nor UO_1551 (O_1551,N_17746,N_18514);
nand UO_1552 (O_1552,N_17127,N_17070);
nor UO_1553 (O_1553,N_16348,N_17937);
xor UO_1554 (O_1554,N_15496,N_18396);
and UO_1555 (O_1555,N_15851,N_15909);
nor UO_1556 (O_1556,N_18239,N_19611);
or UO_1557 (O_1557,N_18891,N_18370);
nand UO_1558 (O_1558,N_18955,N_17140);
nand UO_1559 (O_1559,N_19656,N_15788);
nand UO_1560 (O_1560,N_19336,N_19953);
nor UO_1561 (O_1561,N_19283,N_15425);
nor UO_1562 (O_1562,N_19725,N_18131);
nor UO_1563 (O_1563,N_16685,N_17546);
xnor UO_1564 (O_1564,N_16794,N_19149);
and UO_1565 (O_1565,N_15287,N_17539);
nor UO_1566 (O_1566,N_15463,N_18577);
nand UO_1567 (O_1567,N_17906,N_18838);
nor UO_1568 (O_1568,N_18609,N_15756);
or UO_1569 (O_1569,N_19165,N_17410);
nand UO_1570 (O_1570,N_18311,N_15781);
and UO_1571 (O_1571,N_15696,N_18211);
or UO_1572 (O_1572,N_18703,N_19145);
or UO_1573 (O_1573,N_16171,N_18146);
xnor UO_1574 (O_1574,N_17514,N_15223);
nor UO_1575 (O_1575,N_17464,N_19194);
or UO_1576 (O_1576,N_18824,N_19659);
xnor UO_1577 (O_1577,N_17054,N_19695);
or UO_1578 (O_1578,N_17027,N_16050);
and UO_1579 (O_1579,N_18741,N_18908);
or UO_1580 (O_1580,N_15900,N_19342);
and UO_1581 (O_1581,N_15205,N_16442);
and UO_1582 (O_1582,N_15452,N_15844);
nor UO_1583 (O_1583,N_19126,N_16392);
nor UO_1584 (O_1584,N_18113,N_17450);
xor UO_1585 (O_1585,N_19423,N_16128);
nor UO_1586 (O_1586,N_18507,N_15561);
and UO_1587 (O_1587,N_16882,N_18038);
or UO_1588 (O_1588,N_15420,N_18769);
xnor UO_1589 (O_1589,N_15636,N_19221);
nand UO_1590 (O_1590,N_15595,N_17298);
nor UO_1591 (O_1591,N_18349,N_19465);
nor UO_1592 (O_1592,N_16264,N_18901);
xor UO_1593 (O_1593,N_15549,N_17369);
xnor UO_1594 (O_1594,N_16669,N_17113);
xor UO_1595 (O_1595,N_17230,N_18147);
and UO_1596 (O_1596,N_18652,N_18441);
or UO_1597 (O_1597,N_18602,N_15623);
nand UO_1598 (O_1598,N_15768,N_17949);
or UO_1599 (O_1599,N_17938,N_19887);
or UO_1600 (O_1600,N_15265,N_18390);
and UO_1601 (O_1601,N_17004,N_19956);
or UO_1602 (O_1602,N_17837,N_16266);
nor UO_1603 (O_1603,N_18228,N_15381);
nand UO_1604 (O_1604,N_16462,N_15684);
xnor UO_1605 (O_1605,N_18560,N_16702);
and UO_1606 (O_1606,N_16446,N_17143);
xor UO_1607 (O_1607,N_18878,N_15537);
and UO_1608 (O_1608,N_16306,N_19244);
and UO_1609 (O_1609,N_18066,N_18017);
and UO_1610 (O_1610,N_18300,N_17471);
nand UO_1611 (O_1611,N_19415,N_19347);
and UO_1612 (O_1612,N_17947,N_17946);
xnor UO_1613 (O_1613,N_18238,N_17314);
nor UO_1614 (O_1614,N_19757,N_17668);
xnor UO_1615 (O_1615,N_16045,N_16135);
or UO_1616 (O_1616,N_19711,N_18635);
nor UO_1617 (O_1617,N_19377,N_16152);
xor UO_1618 (O_1618,N_17114,N_15755);
nand UO_1619 (O_1619,N_18888,N_17191);
and UO_1620 (O_1620,N_16673,N_15575);
and UO_1621 (O_1621,N_17840,N_16257);
and UO_1622 (O_1622,N_15437,N_19497);
nor UO_1623 (O_1623,N_16895,N_15669);
xnor UO_1624 (O_1624,N_18218,N_19936);
nor UO_1625 (O_1625,N_17131,N_17554);
nor UO_1626 (O_1626,N_17078,N_17270);
and UO_1627 (O_1627,N_17430,N_19452);
and UO_1628 (O_1628,N_15917,N_17941);
and UO_1629 (O_1629,N_19788,N_15461);
and UO_1630 (O_1630,N_19650,N_18863);
and UO_1631 (O_1631,N_15662,N_16703);
and UO_1632 (O_1632,N_18802,N_17277);
or UO_1633 (O_1633,N_17349,N_15782);
nor UO_1634 (O_1634,N_18949,N_15943);
and UO_1635 (O_1635,N_18496,N_19384);
or UO_1636 (O_1636,N_18125,N_18409);
and UO_1637 (O_1637,N_16214,N_19289);
nand UO_1638 (O_1638,N_17259,N_17788);
xnor UO_1639 (O_1639,N_15318,N_19089);
nor UO_1640 (O_1640,N_18611,N_17063);
nand UO_1641 (O_1641,N_19738,N_16795);
or UO_1642 (O_1642,N_19983,N_19542);
or UO_1643 (O_1643,N_17409,N_18082);
and UO_1644 (O_1644,N_16557,N_15766);
nand UO_1645 (O_1645,N_19270,N_16767);
and UO_1646 (O_1646,N_17272,N_17080);
xnor UO_1647 (O_1647,N_19598,N_19263);
xnor UO_1648 (O_1648,N_16220,N_15184);
xnor UO_1649 (O_1649,N_15194,N_19748);
xnor UO_1650 (O_1650,N_15871,N_16399);
nand UO_1651 (O_1651,N_17339,N_18493);
xnor UO_1652 (O_1652,N_16555,N_15690);
nor UO_1653 (O_1653,N_16769,N_17952);
or UO_1654 (O_1654,N_15747,N_15725);
nor UO_1655 (O_1655,N_18568,N_15133);
and UO_1656 (O_1656,N_16810,N_18526);
nand UO_1657 (O_1657,N_19911,N_17655);
and UO_1658 (O_1658,N_17969,N_17302);
nor UO_1659 (O_1659,N_17351,N_18757);
or UO_1660 (O_1660,N_19058,N_17587);
xor UO_1661 (O_1661,N_16755,N_19045);
nor UO_1662 (O_1662,N_18103,N_17784);
xor UO_1663 (O_1663,N_18231,N_15153);
nand UO_1664 (O_1664,N_15712,N_16690);
nand UO_1665 (O_1665,N_15959,N_15071);
or UO_1666 (O_1666,N_17772,N_15160);
and UO_1667 (O_1667,N_16252,N_15753);
nor UO_1668 (O_1668,N_17077,N_16558);
nor UO_1669 (O_1669,N_15332,N_17135);
xor UO_1670 (O_1670,N_19091,N_19480);
or UO_1671 (O_1671,N_16955,N_15689);
or UO_1672 (O_1672,N_18314,N_18538);
xnor UO_1673 (O_1673,N_16256,N_19366);
or UO_1674 (O_1674,N_16554,N_18626);
nor UO_1675 (O_1675,N_19198,N_16413);
nor UO_1676 (O_1676,N_18525,N_18758);
xor UO_1677 (O_1677,N_18482,N_15443);
nor UO_1678 (O_1678,N_15687,N_18716);
and UO_1679 (O_1679,N_19699,N_19651);
nor UO_1680 (O_1680,N_16400,N_15888);
nor UO_1681 (O_1681,N_15086,N_18631);
nor UO_1682 (O_1682,N_17394,N_15588);
nand UO_1683 (O_1683,N_19821,N_15877);
and UO_1684 (O_1684,N_19759,N_15835);
xnor UO_1685 (O_1685,N_15123,N_15950);
or UO_1686 (O_1686,N_17097,N_17198);
and UO_1687 (O_1687,N_17807,N_15014);
and UO_1688 (O_1688,N_15057,N_19825);
nand UO_1689 (O_1689,N_18653,N_17997);
and UO_1690 (O_1690,N_16310,N_15838);
and UO_1691 (O_1691,N_19049,N_17263);
nor UO_1692 (O_1692,N_17317,N_19890);
nand UO_1693 (O_1693,N_16929,N_19576);
xor UO_1694 (O_1694,N_17636,N_17065);
xnor UO_1695 (O_1695,N_16229,N_19073);
and UO_1696 (O_1696,N_16688,N_17130);
and UO_1697 (O_1697,N_19810,N_18213);
and UO_1698 (O_1698,N_16342,N_17933);
and UO_1699 (O_1699,N_16505,N_18369);
and UO_1700 (O_1700,N_15702,N_15298);
or UO_1701 (O_1701,N_17082,N_16786);
nor UO_1702 (O_1702,N_18753,N_18097);
nor UO_1703 (O_1703,N_18777,N_19797);
nor UO_1704 (O_1704,N_15642,N_17965);
nor UO_1705 (O_1705,N_19864,N_17468);
or UO_1706 (O_1706,N_18292,N_18170);
nor UO_1707 (O_1707,N_16155,N_15180);
nor UO_1708 (O_1708,N_18190,N_15286);
xnor UO_1709 (O_1709,N_17532,N_18022);
nor UO_1710 (O_1710,N_18806,N_17085);
or UO_1711 (O_1711,N_19080,N_17090);
or UO_1712 (O_1712,N_16195,N_18848);
nor UO_1713 (O_1713,N_15674,N_16158);
nor UO_1714 (O_1714,N_15360,N_15814);
nand UO_1715 (O_1715,N_17524,N_18953);
and UO_1716 (O_1716,N_16985,N_18475);
xnor UO_1717 (O_1717,N_17088,N_16427);
xor UO_1718 (O_1718,N_18993,N_18115);
and UO_1719 (O_1719,N_18799,N_18708);
and UO_1720 (O_1720,N_18468,N_18554);
or UO_1721 (O_1721,N_15080,N_17834);
nand UO_1722 (O_1722,N_19021,N_15128);
nor UO_1723 (O_1723,N_19851,N_19944);
xnor UO_1724 (O_1724,N_17278,N_19733);
or UO_1725 (O_1725,N_15313,N_16665);
nand UO_1726 (O_1726,N_15800,N_18896);
nand UO_1727 (O_1727,N_17245,N_19517);
xnor UO_1728 (O_1728,N_19874,N_19667);
and UO_1729 (O_1729,N_15523,N_15898);
xnor UO_1730 (O_1730,N_15038,N_19174);
xor UO_1731 (O_1731,N_19785,N_19592);
or UO_1732 (O_1732,N_19055,N_16273);
nand UO_1733 (O_1733,N_18574,N_18458);
nand UO_1734 (O_1734,N_18122,N_18216);
xor UO_1735 (O_1735,N_19011,N_19255);
and UO_1736 (O_1736,N_19294,N_19420);
or UO_1737 (O_1737,N_19180,N_18425);
nor UO_1738 (O_1738,N_17309,N_17684);
nand UO_1739 (O_1739,N_15309,N_17791);
nor UO_1740 (O_1740,N_19478,N_18541);
nor UO_1741 (O_1741,N_19654,N_19371);
or UO_1742 (O_1742,N_17345,N_15241);
nor UO_1743 (O_1743,N_16086,N_18144);
or UO_1744 (O_1744,N_17849,N_17624);
or UO_1745 (O_1745,N_16023,N_16048);
nor UO_1746 (O_1746,N_15986,N_15415);
nand UO_1747 (O_1747,N_19461,N_15316);
and UO_1748 (O_1748,N_17148,N_18959);
or UO_1749 (O_1749,N_19081,N_17881);
nand UO_1750 (O_1750,N_16695,N_18077);
and UO_1751 (O_1751,N_18346,N_17919);
xor UO_1752 (O_1752,N_15289,N_15283);
nor UO_1753 (O_1753,N_15216,N_18603);
nand UO_1754 (O_1754,N_16428,N_19548);
nor UO_1755 (O_1755,N_16397,N_17520);
xor UO_1756 (O_1756,N_19064,N_19925);
nor UO_1757 (O_1757,N_18917,N_17237);
nor UO_1758 (O_1758,N_16487,N_18008);
or UO_1759 (O_1759,N_16564,N_15956);
xnor UO_1760 (O_1760,N_19906,N_19393);
nor UO_1761 (O_1761,N_18136,N_17152);
or UO_1762 (O_1762,N_17509,N_16747);
or UO_1763 (O_1763,N_17924,N_17665);
nand UO_1764 (O_1764,N_18193,N_19463);
xnor UO_1765 (O_1765,N_19957,N_15699);
or UO_1766 (O_1766,N_17449,N_17517);
or UO_1767 (O_1767,N_15088,N_19671);
xnor UO_1768 (O_1768,N_19007,N_19801);
nor UO_1769 (O_1769,N_15169,N_18776);
or UO_1770 (O_1770,N_15924,N_15164);
or UO_1771 (O_1771,N_15860,N_15993);
and UO_1772 (O_1772,N_19755,N_19883);
nor UO_1773 (O_1773,N_17375,N_15671);
nor UO_1774 (O_1774,N_19404,N_18956);
and UO_1775 (O_1775,N_16640,N_19314);
and UO_1776 (O_1776,N_19379,N_18835);
and UO_1777 (O_1777,N_17392,N_16372);
and UO_1778 (O_1778,N_19535,N_17620);
nor UO_1779 (O_1779,N_19935,N_16459);
nand UO_1780 (O_1780,N_16052,N_19820);
nor UO_1781 (O_1781,N_19107,N_16654);
nand UO_1782 (O_1782,N_15923,N_16721);
and UO_1783 (O_1783,N_16461,N_17347);
nor UO_1784 (O_1784,N_19274,N_15740);
xnor UO_1785 (O_1785,N_17472,N_17079);
or UO_1786 (O_1786,N_18076,N_18018);
and UO_1787 (O_1787,N_16154,N_18293);
nand UO_1788 (O_1788,N_16562,N_15377);
or UO_1789 (O_1789,N_19612,N_16987);
nor UO_1790 (O_1790,N_19118,N_19166);
nor UO_1791 (O_1791,N_18163,N_16516);
xor UO_1792 (O_1792,N_15764,N_16911);
and UO_1793 (O_1793,N_18000,N_19269);
or UO_1794 (O_1794,N_18123,N_16940);
or UO_1795 (O_1795,N_15922,N_16153);
nor UO_1796 (O_1796,N_15021,N_15650);
nor UO_1797 (O_1797,N_15165,N_15641);
nand UO_1798 (O_1798,N_15340,N_16438);
nand UO_1799 (O_1799,N_16662,N_18640);
and UO_1800 (O_1800,N_16828,N_15101);
nand UO_1801 (O_1801,N_18460,N_15967);
or UO_1802 (O_1802,N_16097,N_16075);
nor UO_1803 (O_1803,N_17145,N_19807);
nand UO_1804 (O_1804,N_18127,N_17386);
and UO_1805 (O_1805,N_18052,N_17557);
or UO_1806 (O_1806,N_19012,N_15342);
nor UO_1807 (O_1807,N_15045,N_19636);
nand UO_1808 (O_1808,N_19160,N_17644);
nor UO_1809 (O_1809,N_18754,N_17723);
nand UO_1810 (O_1810,N_16100,N_18308);
nor UO_1811 (O_1811,N_17796,N_19973);
or UO_1812 (O_1812,N_16167,N_15975);
nor UO_1813 (O_1813,N_19351,N_17928);
xor UO_1814 (O_1814,N_18854,N_19984);
nand UO_1815 (O_1815,N_19660,N_16696);
xnor UO_1816 (O_1816,N_17211,N_19706);
nor UO_1817 (O_1817,N_19164,N_18025);
nor UO_1818 (O_1818,N_15887,N_18738);
nor UO_1819 (O_1819,N_17865,N_19286);
and UO_1820 (O_1820,N_19634,N_15819);
or UO_1821 (O_1821,N_15984,N_19352);
nand UO_1822 (O_1822,N_17724,N_17393);
and UO_1823 (O_1823,N_16981,N_17372);
and UO_1824 (O_1824,N_15683,N_15646);
nand UO_1825 (O_1825,N_19124,N_16396);
nor UO_1826 (O_1826,N_19942,N_16354);
nor UO_1827 (O_1827,N_18476,N_17601);
xnor UO_1828 (O_1828,N_16022,N_16018);
or UO_1829 (O_1829,N_17970,N_19500);
or UO_1830 (O_1830,N_17730,N_17758);
or UO_1831 (O_1831,N_15816,N_19316);
and UO_1832 (O_1832,N_19176,N_17089);
and UO_1833 (O_1833,N_19432,N_18788);
xor UO_1834 (O_1834,N_18356,N_17075);
xnor UO_1835 (O_1835,N_15615,N_19185);
nand UO_1836 (O_1836,N_17121,N_19897);
nand UO_1837 (O_1837,N_19661,N_17282);
nand UO_1838 (O_1838,N_18274,N_15527);
xnor UO_1839 (O_1839,N_15983,N_16435);
nand UO_1840 (O_1840,N_19604,N_17475);
or UO_1841 (O_1841,N_16525,N_18821);
or UO_1842 (O_1842,N_16620,N_17281);
and UO_1843 (O_1843,N_18263,N_15400);
nand UO_1844 (O_1844,N_16508,N_17677);
or UO_1845 (O_1845,N_16145,N_16376);
or UO_1846 (O_1846,N_17647,N_16623);
xnor UO_1847 (O_1847,N_17107,N_15214);
nor UO_1848 (O_1848,N_16040,N_15063);
nand UO_1849 (O_1849,N_17197,N_15973);
xor UO_1850 (O_1850,N_15611,N_17868);
xor UO_1851 (O_1851,N_15773,N_17984);
nor UO_1852 (O_1852,N_16877,N_17559);
or UO_1853 (O_1853,N_18790,N_16597);
nand UO_1854 (O_1854,N_17425,N_16660);
or UO_1855 (O_1855,N_17368,N_19235);
xnor UO_1856 (O_1856,N_18183,N_19837);
and UO_1857 (O_1857,N_18237,N_18916);
xor UO_1858 (O_1858,N_18429,N_19077);
nand UO_1859 (O_1859,N_16223,N_16819);
nor UO_1860 (O_1860,N_15832,N_18978);
or UO_1861 (O_1861,N_17218,N_16902);
and UO_1862 (O_1862,N_16316,N_17822);
nand UO_1863 (O_1863,N_17683,N_19629);
nand UO_1864 (O_1864,N_15074,N_15475);
nand UO_1865 (O_1865,N_19736,N_15299);
nor UO_1866 (O_1866,N_17209,N_15262);
or UO_1867 (O_1867,N_15522,N_15469);
xor UO_1868 (O_1868,N_17452,N_17251);
and UO_1869 (O_1869,N_18852,N_19946);
xor UO_1870 (O_1870,N_18664,N_16566);
or UO_1871 (O_1871,N_19487,N_15808);
xor UO_1872 (O_1872,N_19985,N_17800);
and UO_1873 (O_1873,N_18444,N_16658);
xnor UO_1874 (O_1874,N_17172,N_17308);
and UO_1875 (O_1875,N_16862,N_17052);
or UO_1876 (O_1876,N_19201,N_17485);
and UO_1877 (O_1877,N_17123,N_15531);
nand UO_1878 (O_1878,N_16114,N_18851);
nand UO_1879 (O_1879,N_17703,N_18656);
or UO_1880 (O_1880,N_17569,N_15876);
xor UO_1881 (O_1881,N_19844,N_16244);
xnor UO_1882 (O_1882,N_19229,N_16930);
nand UO_1883 (O_1883,N_17897,N_19422);
or UO_1884 (O_1884,N_17275,N_16425);
or UO_1885 (O_1885,N_19157,N_16712);
nor UO_1886 (O_1886,N_19197,N_15362);
xor UO_1887 (O_1887,N_17323,N_19297);
or UO_1888 (O_1888,N_15005,N_18212);
xor UO_1889 (O_1889,N_19537,N_19914);
or UO_1890 (O_1890,N_18742,N_17657);
nand UO_1891 (O_1891,N_18316,N_17762);
nand UO_1892 (O_1892,N_15070,N_17744);
and UO_1893 (O_1893,N_15859,N_16880);
or UO_1894 (O_1894,N_18379,N_17858);
nand UO_1895 (O_1895,N_15769,N_17461);
nor UO_1896 (O_1896,N_19928,N_15089);
and UO_1897 (O_1897,N_15661,N_18414);
or UO_1898 (O_1898,N_18857,N_18517);
and UO_1899 (O_1899,N_19216,N_16156);
and UO_1900 (O_1900,N_17116,N_15479);
nand UO_1901 (O_1901,N_17794,N_18388);
xor UO_1902 (O_1902,N_18585,N_15562);
and UO_1903 (O_1903,N_19071,N_15092);
nand UO_1904 (O_1904,N_18223,N_19715);
and UO_1905 (O_1905,N_16847,N_19910);
or UO_1906 (O_1906,N_16044,N_18615);
or UO_1907 (O_1907,N_18340,N_15598);
nand UO_1908 (O_1908,N_16784,N_16301);
nor UO_1909 (O_1909,N_16651,N_19163);
or UO_1910 (O_1910,N_17141,N_19846);
nand UO_1911 (O_1911,N_15426,N_17316);
xnor UO_1912 (O_1912,N_15542,N_18584);
nand UO_1913 (O_1913,N_17637,N_18357);
or UO_1914 (O_1914,N_17845,N_18084);
xnor UO_1915 (O_1915,N_15401,N_19730);
xor UO_1916 (O_1916,N_15116,N_16853);
and UO_1917 (O_1917,N_15880,N_17966);
nor UO_1918 (O_1918,N_15660,N_17342);
or UO_1919 (O_1919,N_18322,N_16469);
and UO_1920 (O_1920,N_16609,N_17280);
nor UO_1921 (O_1921,N_15978,N_15326);
or UO_1922 (O_1922,N_16200,N_18313);
nor UO_1923 (O_1923,N_15002,N_17319);
and UO_1924 (O_1924,N_18497,N_19134);
nand UO_1925 (O_1925,N_16831,N_16141);
and UO_1926 (O_1926,N_18975,N_15939);
xnor UO_1927 (O_1927,N_16295,N_17244);
nand UO_1928 (O_1928,N_17177,N_17473);
or UO_1929 (O_1929,N_17486,N_16000);
and UO_1930 (O_1930,N_16007,N_16248);
nor UO_1931 (O_1931,N_17202,N_16453);
nor UO_1932 (O_1932,N_16957,N_17963);
nand UO_1933 (O_1933,N_17203,N_16871);
nor UO_1934 (O_1934,N_18591,N_16279);
nor UO_1935 (O_1935,N_18528,N_17526);
and UO_1936 (O_1936,N_16743,N_16980);
nand UO_1937 (O_1937,N_19974,N_18116);
nor UO_1938 (O_1938,N_19027,N_16068);
nand UO_1939 (O_1939,N_19139,N_17348);
nand UO_1940 (O_1940,N_16315,N_19813);
or UO_1941 (O_1941,N_19308,N_16731);
nand UO_1942 (O_1942,N_16151,N_17830);
xnor UO_1943 (O_1943,N_19561,N_18718);
xor UO_1944 (O_1944,N_17609,N_16914);
or UO_1945 (O_1945,N_17789,N_15099);
xor UO_1946 (O_1946,N_19516,N_17871);
or UO_1947 (O_1947,N_18225,N_17331);
and UO_1948 (O_1948,N_18360,N_16165);
xor UO_1949 (O_1949,N_17561,N_15711);
nand UO_1950 (O_1950,N_19079,N_18265);
nor UO_1951 (O_1951,N_16808,N_17870);
nor UO_1952 (O_1952,N_16418,N_16501);
xor UO_1953 (O_1953,N_18143,N_18057);
and UO_1954 (O_1954,N_15546,N_18740);
nor UO_1955 (O_1955,N_16433,N_19609);
nand UO_1956 (O_1956,N_18244,N_15566);
nor UO_1957 (O_1957,N_19597,N_15664);
nand UO_1958 (O_1958,N_17971,N_16693);
or UO_1959 (O_1959,N_17821,N_16211);
nor UO_1960 (O_1960,N_17786,N_17769);
and UO_1961 (O_1961,N_17015,N_16389);
xnor UO_1962 (O_1962,N_17574,N_16122);
nand UO_1963 (O_1963,N_15065,N_19303);
xor UO_1964 (O_1964,N_15845,N_18167);
nor UO_1965 (O_1965,N_17050,N_17994);
xor UO_1966 (O_1966,N_16534,N_18855);
and UO_1967 (O_1967,N_18620,N_15543);
nand UO_1968 (O_1968,N_17086,N_18461);
nor UO_1969 (O_1969,N_15137,N_18310);
or UO_1970 (O_1970,N_15451,N_16464);
or UO_1971 (O_1971,N_16891,N_18569);
and UO_1972 (O_1972,N_15163,N_17006);
xor UO_1973 (O_1973,N_17671,N_17307);
nor UO_1974 (O_1974,N_19390,N_18309);
or UO_1975 (O_1975,N_15179,N_19745);
nor UO_1976 (O_1976,N_17404,N_18523);
nor UO_1977 (O_1977,N_16939,N_17208);
xor UO_1978 (O_1978,N_18049,N_17025);
xnor UO_1979 (O_1979,N_17735,N_17112);
nor UO_1980 (O_1980,N_18065,N_16887);
and UO_1981 (O_1981,N_18382,N_19312);
or UO_1982 (O_1982,N_16809,N_16901);
or UO_1983 (O_1983,N_16868,N_16181);
or UO_1984 (O_1984,N_17039,N_15077);
and UO_1985 (O_1985,N_15853,N_18849);
xnor UO_1986 (O_1986,N_18575,N_15058);
xor UO_1987 (O_1987,N_17948,N_17787);
nand UO_1988 (O_1988,N_18198,N_17046);
and UO_1989 (O_1989,N_19827,N_18672);
or UO_1990 (O_1990,N_16478,N_19817);
and UO_1991 (O_1991,N_19281,N_18981);
nand UO_1992 (O_1992,N_17592,N_15691);
and UO_1993 (O_1993,N_17428,N_15514);
or UO_1994 (O_1994,N_18599,N_18985);
or UO_1995 (O_1995,N_18756,N_18397);
and UO_1996 (O_1996,N_19495,N_17504);
nand UO_1997 (O_1997,N_16850,N_19103);
nor UO_1998 (O_1998,N_16430,N_19665);
xnor UO_1999 (O_1999,N_19639,N_19443);
or UO_2000 (O_2000,N_18544,N_18164);
nor UO_2001 (O_2001,N_19065,N_19571);
or UO_2002 (O_2002,N_19934,N_18045);
nand UO_2003 (O_2003,N_16509,N_18641);
nand UO_2004 (O_2004,N_17364,N_16074);
nand UO_2005 (O_2005,N_15538,N_16353);
and UO_2006 (O_2006,N_15529,N_19070);
or UO_2007 (O_2007,N_16378,N_18836);
or UO_2008 (O_2008,N_18055,N_15132);
or UO_2009 (O_2009,N_19686,N_16913);
or UO_2010 (O_2010,N_17255,N_18191);
nand UO_2011 (O_2011,N_17153,N_15706);
and UO_2012 (O_2012,N_19503,N_16330);
or UO_2013 (O_2013,N_16993,N_19860);
xor UO_2014 (O_2014,N_18508,N_15910);
nor UO_2015 (O_2015,N_17888,N_15499);
nor UO_2016 (O_2016,N_18197,N_16005);
nand UO_2017 (O_2017,N_16750,N_15926);
and UO_2018 (O_2018,N_17165,N_17242);
nand UO_2019 (O_2019,N_19567,N_16541);
or UO_2020 (O_2020,N_17699,N_16017);
nand UO_2021 (O_2021,N_16589,N_17126);
nand UO_2022 (O_2022,N_19335,N_15839);
xnor UO_2023 (O_2023,N_19484,N_17408);
nor UO_2024 (O_2024,N_17493,N_19088);
or UO_2025 (O_2025,N_17332,N_16241);
and UO_2026 (O_2026,N_16054,N_16909);
and UO_2027 (O_2027,N_17478,N_16305);
nand UO_2028 (O_2028,N_15855,N_17221);
nor UO_2029 (O_2029,N_19313,N_15858);
or UO_2030 (O_2030,N_18999,N_15027);
nor UO_2031 (O_2031,N_19243,N_19710);
or UO_2032 (O_2032,N_16443,N_18623);
nor UO_2033 (O_2033,N_16883,N_17525);
nand UO_2034 (O_2034,N_15927,N_19066);
or UO_2035 (O_2035,N_16633,N_15916);
nor UO_2036 (O_2036,N_15012,N_19491);
and UO_2037 (O_2037,N_19192,N_18505);
nand UO_2038 (O_2038,N_18154,N_16602);
nor UO_2039 (O_2039,N_18121,N_19995);
and UO_2040 (O_2040,N_18207,N_15427);
and UO_2041 (O_2041,N_15364,N_17886);
xor UO_2042 (O_2042,N_17305,N_16905);
xor UO_2043 (O_2043,N_19621,N_16403);
xor UO_2044 (O_2044,N_17099,N_19620);
or UO_2045 (O_2045,N_19945,N_16012);
xnor UO_2046 (O_2046,N_16070,N_15441);
xor UO_2047 (O_2047,N_16238,N_15494);
nand UO_2048 (O_2048,N_16734,N_15964);
nor UO_2049 (O_2049,N_18892,N_16077);
nand UO_2050 (O_2050,N_17793,N_18637);
xor UO_2051 (O_2051,N_18235,N_19407);
and UO_2052 (O_2052,N_19424,N_19903);
and UO_2053 (O_2053,N_16657,N_18687);
or UO_2054 (O_2054,N_16735,N_16170);
xnor UO_2055 (O_2055,N_18227,N_15941);
nand UO_2056 (O_2056,N_15613,N_18473);
and UO_2057 (O_2057,N_19121,N_16607);
and UO_2058 (O_2058,N_18576,N_17912);
xnor UO_2059 (O_2059,N_16169,N_16488);
nand UO_2060 (O_2060,N_15524,N_15237);
and UO_2061 (O_2061,N_16038,N_15938);
nor UO_2062 (O_2062,N_19879,N_17189);
or UO_2063 (O_2063,N_17463,N_15447);
or UO_2064 (O_2064,N_19225,N_15825);
nand UO_2065 (O_2065,N_15570,N_18362);
nor UO_2066 (O_2066,N_16544,N_19402);
and UO_2067 (O_2067,N_17108,N_19032);
or UO_2068 (O_2068,N_17687,N_19115);
xor UO_2069 (O_2069,N_17487,N_15430);
or UO_2070 (O_2070,N_17294,N_15023);
xor UO_2071 (O_2071,N_19869,N_15458);
nand UO_2072 (O_2072,N_19931,N_18321);
or UO_2073 (O_2073,N_18659,N_17030);
xor UO_2074 (O_2074,N_17353,N_16801);
or UO_2075 (O_2075,N_17196,N_15873);
nand UO_2076 (O_2076,N_16718,N_17768);
and UO_2077 (O_2077,N_19170,N_15303);
or UO_2078 (O_2078,N_15222,N_15637);
nor UO_2079 (O_2079,N_18589,N_18734);
or UO_2080 (O_2080,N_18692,N_15261);
nor UO_2081 (O_2081,N_15230,N_17710);
nand UO_2082 (O_2082,N_19311,N_16079);
nand UO_2083 (O_2083,N_19898,N_16500);
nand UO_2084 (O_2084,N_15064,N_17674);
nor UO_2085 (O_2085,N_15357,N_16434);
nand UO_2086 (O_2086,N_17382,N_16368);
nand UO_2087 (O_2087,N_19372,N_15732);
and UO_2088 (O_2088,N_15555,N_17745);
and UO_2089 (O_2089,N_18345,N_18206);
xor UO_2090 (O_2090,N_18871,N_18302);
and UO_2091 (O_2091,N_15320,N_19140);
and UO_2092 (O_2092,N_15954,N_17558);
nand UO_2093 (O_2093,N_16758,N_18976);
nand UO_2094 (O_2094,N_18906,N_19082);
or UO_2095 (O_2095,N_16692,N_16697);
or UO_2096 (O_2096,N_17133,N_17756);
xor UO_2097 (O_2097,N_19362,N_19777);
and UO_2098 (O_2098,N_16021,N_18805);
and UO_2099 (O_2099,N_15815,N_15765);
nand UO_2100 (O_2100,N_15930,N_16879);
nand UO_2101 (O_2101,N_16604,N_15682);
or UO_2102 (O_2102,N_15204,N_15048);
xor UO_2103 (O_2103,N_19741,N_15347);
nor UO_2104 (O_2104,N_19302,N_16884);
or UO_2105 (O_2105,N_18162,N_19577);
nor UO_2106 (O_2106,N_16730,N_17595);
or UO_2107 (O_2107,N_18063,N_19104);
xor UO_2108 (O_2108,N_15453,N_15297);
xnor UO_2109 (O_2109,N_19657,N_19051);
nand UO_2110 (O_2110,N_19318,N_17551);
or UO_2111 (O_2111,N_16645,N_15783);
nor UO_2112 (O_2112,N_15576,N_19353);
xor UO_2113 (O_2113,N_16110,N_18928);
nor UO_2114 (O_2114,N_18782,N_17972);
or UO_2115 (O_2115,N_16559,N_15069);
nand UO_2116 (O_2116,N_15231,N_17579);
and UO_2117 (O_2117,N_17565,N_16476);
nand UO_2118 (O_2118,N_17188,N_15245);
and UO_2119 (O_2119,N_17361,N_15951);
or UO_2120 (O_2120,N_17631,N_15176);
xor UO_2121 (O_2121,N_16528,N_16822);
or UO_2122 (O_2122,N_17716,N_19472);
nand UO_2123 (O_2123,N_17180,N_18276);
xor UO_2124 (O_2124,N_17274,N_18415);
nor UO_2125 (O_2125,N_15886,N_17212);
nor UO_2126 (O_2126,N_18030,N_18759);
or UO_2127 (O_2127,N_19792,N_17503);
xnor UO_2128 (O_2128,N_16437,N_18561);
nor UO_2129 (O_2129,N_15980,N_16715);
nor UO_2130 (O_2130,N_17814,N_16076);
and UO_2131 (O_2131,N_15789,N_17396);
or UO_2132 (O_2132,N_16423,N_17087);
or UO_2133 (O_2133,N_16531,N_16041);
or UO_2134 (O_2134,N_18222,N_16366);
nand UO_2135 (O_2135,N_15138,N_19940);
or UO_2136 (O_2136,N_17437,N_15897);
xnor UO_2137 (O_2137,N_19207,N_17641);
or UO_2138 (O_2138,N_18822,N_19949);
and UO_2139 (O_2139,N_16944,N_19391);
and UO_2140 (O_2140,N_17124,N_16577);
xor UO_2141 (O_2141,N_16267,N_16206);
nor UO_2142 (O_2142,N_17738,N_18952);
nand UO_2143 (O_2143,N_17638,N_15418);
and UO_2144 (O_2144,N_17490,N_15899);
and UO_2145 (O_2145,N_15526,N_18104);
nand UO_2146 (O_2146,N_17779,N_19727);
xnor UO_2147 (O_2147,N_19381,N_18499);
nor UO_2148 (O_2148,N_15246,N_18483);
xnor UO_2149 (O_2149,N_17838,N_17698);
nor UO_2150 (O_2150,N_17670,N_18684);
or UO_2151 (O_2151,N_16691,N_15131);
nand UO_2152 (O_2152,N_18093,N_17286);
nor UO_2153 (O_2153,N_19467,N_17995);
xnor UO_2154 (O_2154,N_16811,N_15271);
or UO_2155 (O_2155,N_17905,N_19240);
nor UO_2156 (O_2156,N_16189,N_15673);
xnor UO_2157 (O_2157,N_15056,N_15824);
or UO_2158 (O_2158,N_19978,N_15114);
or UO_2159 (O_2159,N_18463,N_16998);
or UO_2160 (O_2160,N_18157,N_16417);
nor UO_2161 (O_2161,N_18516,N_18816);
and UO_2162 (O_2162,N_17752,N_17119);
xnor UO_2163 (O_2163,N_17615,N_17014);
nand UO_2164 (O_2164,N_19543,N_16274);
and UO_2165 (O_2165,N_17066,N_19684);
or UO_2166 (O_2166,N_16514,N_15911);
nand UO_2167 (O_2167,N_18986,N_15094);
xor UO_2168 (O_2168,N_19002,N_17673);
and UO_2169 (O_2169,N_17445,N_15564);
nand UO_2170 (O_2170,N_19075,N_15239);
nand UO_2171 (O_2171,N_15209,N_16280);
xor UO_2172 (O_2172,N_18671,N_18445);
nor UO_2173 (O_2173,N_19640,N_18655);
or UO_2174 (O_2174,N_19551,N_17071);
and UO_2175 (O_2175,N_18521,N_19220);
and UO_2176 (O_2176,N_17336,N_18411);
and UO_2177 (O_2177,N_17283,N_17513);
nand UO_2178 (O_2178,N_18702,N_15569);
or UO_2179 (O_2179,N_17982,N_16970);
nor UO_2180 (O_2180,N_15181,N_17069);
nor UO_2181 (O_2181,N_18841,N_19236);
or UO_2182 (O_2182,N_16176,N_18563);
and UO_2183 (O_2183,N_15867,N_15821);
and UO_2184 (O_2184,N_18286,N_15167);
xor UO_2185 (O_2185,N_16191,N_17915);
nand UO_2186 (O_2186,N_19676,N_17646);
and UO_2187 (O_2187,N_17005,N_17895);
xor UO_2188 (O_2188,N_16496,N_15337);
nor UO_2189 (O_2189,N_19179,N_16983);
nand UO_2190 (O_2190,N_16785,N_18003);
or UO_2191 (O_2191,N_17334,N_17215);
nor UO_2192 (O_2192,N_18342,N_16148);
nor UO_2193 (O_2193,N_18895,N_17252);
nor UO_2194 (O_2194,N_18804,N_15267);
or UO_2195 (O_2195,N_17081,N_15484);
nor UO_2196 (O_2196,N_17651,N_16719);
xor UO_2197 (O_2197,N_17552,N_15820);
xnor UO_2198 (O_2198,N_17419,N_17455);
nand UO_2199 (O_2199,N_16722,N_18479);
nand UO_2200 (O_2200,N_18270,N_16201);
or UO_2201 (O_2201,N_16080,N_15785);
or UO_2202 (O_2202,N_15278,N_15812);
and UO_2203 (O_2203,N_16699,N_15110);
xnor UO_2204 (O_2204,N_19587,N_15921);
nand UO_2205 (O_2205,N_18376,N_17750);
and UO_2206 (O_2206,N_19688,N_19447);
nor UO_2207 (O_2207,N_19641,N_15208);
nor UO_2208 (O_2208,N_16896,N_17676);
xor UO_2209 (O_2209,N_15040,N_19692);
xnor UO_2210 (O_2210,N_19979,N_16821);
nand UO_2211 (O_2211,N_17441,N_19878);
nor UO_2212 (O_2212,N_18942,N_16670);
xnor UO_2213 (O_2213,N_17867,N_19454);
nor UO_2214 (O_2214,N_18332,N_18142);
or UO_2215 (O_2215,N_19756,N_18839);
xnor UO_2216 (O_2216,N_17623,N_16193);
nand UO_2217 (O_2217,N_17125,N_15382);
nand UO_2218 (O_2218,N_19557,N_16630);
or UO_2219 (O_2219,N_15419,N_19466);
nor UO_2220 (O_2220,N_19865,N_18434);
nand UO_2221 (O_2221,N_18926,N_19572);
nor UO_2222 (O_2222,N_19761,N_19400);
xnor UO_2223 (O_2223,N_19462,N_17184);
nand UO_2224 (O_2224,N_17645,N_17482);
nand UO_2225 (O_2225,N_17802,N_18647);
xnor UO_2226 (O_2226,N_19258,N_19189);
nor UO_2227 (O_2227,N_15593,N_17018);
xor UO_2228 (O_2228,N_15028,N_16800);
nand UO_2229 (O_2229,N_15977,N_16338);
nor UO_2230 (O_2230,N_15802,N_19876);
or UO_2231 (O_2231,N_18012,N_17183);
nand UO_2232 (O_2232,N_16600,N_18485);
xnor UO_2233 (O_2233,N_18259,N_19188);
xnor UO_2234 (O_2234,N_17591,N_19600);
and UO_2235 (O_2235,N_19175,N_18108);
xor UO_2236 (O_2236,N_15601,N_17944);
xnor UO_2237 (O_2237,N_18013,N_16838);
nand UO_2238 (O_2238,N_18072,N_19181);
xor UO_2239 (O_2239,N_18075,N_16492);
nor UO_2240 (O_2240,N_16485,N_17889);
or UO_2241 (O_2241,N_16491,N_15872);
nand UO_2242 (O_2242,N_15152,N_17826);
nand UO_2243 (O_2243,N_19716,N_17732);
and UO_2244 (O_2244,N_17026,N_19268);
nand UO_2245 (O_2245,N_19460,N_16016);
nand UO_2246 (O_2246,N_19682,N_15931);
and UO_2247 (O_2247,N_15462,N_17341);
nand UO_2248 (O_2248,N_16989,N_15260);
or UO_2249 (O_2249,N_19778,N_17975);
nand UO_2250 (O_2250,N_18081,N_17013);
xnor UO_2251 (O_2251,N_17397,N_19392);
nor UO_2252 (O_2252,N_19232,N_17776);
nor UO_2253 (O_2253,N_17501,N_17083);
or UO_2254 (O_2254,N_19213,N_18005);
nor UO_2255 (O_2255,N_16025,N_15581);
xor UO_2256 (O_2256,N_17989,N_19814);
or UO_2257 (O_2257,N_18709,N_16638);
nand UO_2258 (O_2258,N_19248,N_18634);
xor UO_2259 (O_2259,N_16511,N_15688);
and UO_2260 (O_2260,N_15729,N_15135);
xor UO_2261 (O_2261,N_18924,N_17296);
and UO_2262 (O_2262,N_15720,N_17618);
or UO_2263 (O_2263,N_15456,N_17686);
and UO_2264 (O_2264,N_19926,N_18011);
nand UO_2265 (O_2265,N_15472,N_17306);
nor UO_2266 (O_2266,N_15865,N_19417);
xor UO_2267 (O_2267,N_17850,N_19306);
xnor UO_2268 (O_2268,N_15171,N_15987);
nor UO_2269 (O_2269,N_18490,N_15630);
xnor UO_2270 (O_2270,N_17175,N_15585);
nor UO_2271 (O_2271,N_15582,N_19707);
and UO_2272 (O_2272,N_16364,N_17367);
or UO_2273 (O_2273,N_17144,N_18203);
nand UO_2274 (O_2274,N_15322,N_18459);
nand UO_2275 (O_2275,N_18046,N_16825);
or UO_2276 (O_2276,N_16503,N_19321);
nand UO_2277 (O_2277,N_16361,N_15158);
nor UO_2278 (O_2278,N_16587,N_19764);
xor UO_2279 (O_2279,N_18064,N_15716);
nor UO_2280 (O_2280,N_19435,N_17599);
or UO_2281 (O_2281,N_19469,N_19172);
or UO_2282 (O_2282,N_15659,N_16759);
nand UO_2283 (O_2283,N_18793,N_18378);
nor UO_2284 (O_2284,N_18667,N_18153);
nor UO_2285 (O_2285,N_17190,N_15717);
xor UO_2286 (O_2286,N_17940,N_15136);
nor UO_2287 (O_2287,N_17511,N_18557);
and UO_2288 (O_2288,N_17205,N_19364);
nor UO_2289 (O_2289,N_17660,N_15675);
and UO_2290 (O_2290,N_16088,N_19048);
xor UO_2291 (O_2291,N_15026,N_15852);
nor UO_2292 (O_2292,N_19619,N_17568);
xnor UO_2293 (O_2293,N_16581,N_19558);
or UO_2294 (O_2294,N_18043,N_17980);
nand UO_2295 (O_2295,N_16393,N_19200);
or UO_2296 (O_2296,N_18070,N_17570);
or UO_2297 (O_2297,N_19766,N_18226);
or UO_2298 (O_2298,N_19489,N_15843);
and UO_2299 (O_2299,N_18983,N_16724);
or UO_2300 (O_2300,N_19375,N_16481);
nor UO_2301 (O_2301,N_16121,N_15375);
and UO_2302 (O_2302,N_18648,N_18760);
nor UO_2303 (O_2303,N_19130,N_16738);
nor UO_2304 (O_2304,N_16617,N_16906);
nand UO_2305 (O_2305,N_19413,N_19627);
xnor UO_2306 (O_2306,N_18947,N_15509);
or UO_2307 (O_2307,N_19528,N_19880);
or UO_2308 (O_2308,N_17413,N_16391);
or UO_2309 (O_2309,N_17761,N_16628);
xnor UO_2310 (O_2310,N_18061,N_17987);
nand UO_2311 (O_2311,N_16539,N_16898);
or UO_2312 (O_2312,N_18813,N_16839);
and UO_2313 (O_2313,N_18451,N_18646);
and UO_2314 (O_2314,N_18783,N_15721);
nor UO_2315 (O_2315,N_18705,N_15102);
and UO_2316 (O_2316,N_19693,N_17812);
nand UO_2317 (O_2317,N_15270,N_18480);
and UO_2318 (O_2318,N_19616,N_15535);
nor UO_2319 (O_2319,N_18698,N_17586);
xnor UO_2320 (O_2320,N_17210,N_17988);
or UO_2321 (O_2321,N_15635,N_16329);
nand UO_2322 (O_2322,N_18181,N_15125);
and UO_2323 (O_2323,N_16652,N_18051);
or UO_2324 (O_2324,N_16036,N_19840);
nor UO_2325 (O_2325,N_17757,N_19540);
nor UO_2326 (O_2326,N_19867,N_17545);
nor UO_2327 (O_2327,N_19905,N_16326);
and UO_2328 (O_2328,N_15969,N_16395);
or UO_2329 (O_2329,N_19608,N_17803);
nand UO_2330 (O_2330,N_16069,N_18202);
or UO_2331 (O_2331,N_16140,N_15550);
nor UO_2332 (O_2332,N_16458,N_15589);
and UO_2333 (O_2333,N_17639,N_18470);
nor UO_2334 (O_2334,N_16723,N_17477);
or UO_2335 (O_2335,N_16588,N_16526);
and UO_2336 (O_2336,N_17110,N_17855);
nand UO_2337 (O_2337,N_18234,N_16085);
and UO_2338 (O_2338,N_15275,N_17866);
nor UO_2339 (O_2339,N_19723,N_17276);
nand UO_2340 (O_2340,N_17326,N_16350);
and UO_2341 (O_2341,N_18098,N_16798);
or UO_2342 (O_2342,N_16908,N_15292);
and UO_2343 (O_2343,N_18252,N_19214);
nand UO_2344 (O_2344,N_15445,N_16869);
nor UO_2345 (O_2345,N_17320,N_17429);
nand UO_2346 (O_2346,N_18690,N_16543);
and UO_2347 (O_2347,N_15449,N_18095);
and UO_2348 (O_2348,N_15103,N_16668);
and UO_2349 (O_2349,N_18488,N_18392);
or UO_2350 (O_2350,N_16374,N_17795);
nor UO_2351 (O_2351,N_16115,N_19538);
xnor UO_2352 (O_2352,N_17921,N_19904);
xor UO_2353 (O_2353,N_16370,N_18531);
nor UO_2354 (O_2354,N_15610,N_18996);
xor UO_2355 (O_2355,N_18042,N_17008);
and UO_2356 (O_2356,N_16552,N_19780);
xnor UO_2357 (O_2357,N_15709,N_15493);
nor UO_2358 (O_2358,N_15703,N_19028);
nor UO_2359 (O_2359,N_19653,N_16134);
xnor UO_2360 (O_2360,N_18141,N_18486);
xnor UO_2361 (O_2361,N_18666,N_19758);
and UO_2362 (O_2362,N_18294,N_15719);
and UO_2363 (O_2363,N_18594,N_15412);
and UO_2364 (O_2364,N_19068,N_15020);
nand UO_2365 (O_2365,N_16475,N_17068);
xnor UO_2366 (O_2366,N_15621,N_15864);
or UO_2367 (O_2367,N_19265,N_18530);
or UO_2368 (O_2368,N_15221,N_18132);
and UO_2369 (O_2369,N_15644,N_16032);
and UO_2370 (O_2370,N_16856,N_15073);
xor UO_2371 (O_2371,N_15597,N_15685);
nor UO_2372 (O_2372,N_19530,N_18255);
or UO_2373 (O_2373,N_19098,N_17869);
nand UO_2374 (O_2374,N_16632,N_16245);
nand UO_2375 (O_2375,N_18440,N_17911);
nor UO_2376 (O_2376,N_19482,N_15548);
or UO_2377 (O_2377,N_17362,N_17741);
nand UO_2378 (O_2378,N_19298,N_16394);
nor UO_2379 (O_2379,N_19276,N_15433);
nand UO_2380 (O_2380,N_18477,N_18688);
xor UO_2381 (O_2381,N_19586,N_19322);
xnor UO_2382 (O_2382,N_15206,N_18283);
and UO_2383 (O_2383,N_16293,N_16026);
nor UO_2384 (O_2384,N_16493,N_17411);
xnor UO_2385 (O_2385,N_16530,N_15018);
and UO_2386 (O_2386,N_16323,N_17321);
nand UO_2387 (O_2387,N_17731,N_15346);
nand UO_2388 (O_2388,N_15202,N_19742);
xor UO_2389 (O_2389,N_15652,N_16062);
and UO_2390 (O_2390,N_18101,N_18710);
nand UO_2391 (O_2391,N_19204,N_16804);
xnor UO_2392 (O_2392,N_16083,N_19458);
nand UO_2393 (O_2393,N_17510,N_17672);
xnor UO_2394 (O_2394,N_15256,N_16456);
nand UO_2395 (O_2395,N_19430,N_18715);
nand UO_2396 (O_2396,N_17357,N_19998);
xor UO_2397 (O_2397,N_19233,N_19855);
nand UO_2398 (O_2398,N_15648,N_17536);
and UO_2399 (O_2399,N_18351,N_19178);
xor UO_2400 (O_2400,N_19383,N_19182);
or UO_2401 (O_2401,N_15201,N_16726);
nand UO_2402 (O_2402,N_16349,N_18361);
nor UO_2403 (O_2403,N_18264,N_15282);
xnor UO_2404 (O_2404,N_18106,N_16149);
nor UO_2405 (O_2405,N_17578,N_16878);
nand UO_2406 (O_2406,N_19187,N_16131);
xor UO_2407 (O_2407,N_15778,N_19961);
or UO_2408 (O_2408,N_19791,N_16560);
xor UO_2409 (O_2409,N_16728,N_15643);
nor UO_2410 (O_2410,N_15359,N_19849);
nand UO_2411 (O_2411,N_19739,N_18961);
xnor UO_2412 (O_2412,N_19210,N_15120);
nor UO_2413 (O_2413,N_18823,N_16997);
nor UO_2414 (O_2414,N_19227,N_17979);
or UO_2415 (O_2415,N_18970,N_19029);
nor UO_2416 (O_2416,N_15474,N_17007);
nand UO_2417 (O_2417,N_16215,N_18654);
xnor UO_2418 (O_2418,N_16616,N_17953);
xnor UO_2419 (O_2419,N_17223,N_16172);
and UO_2420 (O_2420,N_16218,N_15668);
xnor UO_2421 (O_2421,N_16756,N_15741);
and UO_2422 (O_2422,N_15464,N_16793);
and UO_2423 (O_2423,N_16362,N_16708);
and UO_2424 (O_2424,N_16143,N_15109);
or UO_2425 (O_2425,N_17406,N_18242);
or UO_2426 (O_2426,N_15082,N_17736);
and UO_2427 (O_2427,N_18128,N_18869);
nor UO_2428 (O_2428,N_18837,N_16339);
and UO_2429 (O_2429,N_18118,N_19343);
nor UO_2430 (O_2430,N_19615,N_18233);
xor UO_2431 (O_2431,N_15560,N_16622);
nand UO_2432 (O_2432,N_18489,N_18812);
nand UO_2433 (O_2433,N_18697,N_17918);
or UO_2434 (O_2434,N_15156,N_18931);
and UO_2435 (O_2435,N_19668,N_19309);
and UO_2436 (O_2436,N_19915,N_16996);
nor UO_2437 (O_2437,N_15465,N_17370);
and UO_2438 (O_2438,N_15015,N_16510);
or UO_2439 (O_2439,N_16390,N_17359);
xnor UO_2440 (O_2440,N_18678,N_18668);
nor UO_2441 (O_2441,N_15866,N_15226);
and UO_2442 (O_2442,N_18251,N_16634);
or UO_2443 (O_2443,N_16506,N_15277);
or UO_2444 (O_2444,N_17689,N_15148);
xnor UO_2445 (O_2445,N_17179,N_19315);
and UO_2446 (O_2446,N_16842,N_19030);
or UO_2447 (O_2447,N_16737,N_17022);
nor UO_2448 (O_2448,N_18007,N_16966);
nand UO_2449 (O_2449,N_19005,N_18601);
or UO_2450 (O_2450,N_15746,N_18194);
xnor UO_2451 (O_2451,N_16159,N_17160);
nor UO_2452 (O_2452,N_18875,N_18328);
xnor UO_2453 (O_2453,N_18325,N_19583);
xor UO_2454 (O_2454,N_16965,N_19024);
xnor UO_2455 (O_2455,N_19439,N_15257);
or UO_2456 (O_2456,N_15024,N_17718);
or UO_2457 (O_2457,N_18927,N_19223);
nand UO_2458 (O_2458,N_17664,N_15236);
xnor UO_2459 (O_2459,N_17041,N_17023);
nor UO_2460 (O_2460,N_16186,N_17169);
nor UO_2461 (O_2461,N_15490,N_15378);
and UO_2462 (O_2462,N_16113,N_18323);
or UO_2463 (O_2463,N_15596,N_19638);
and UO_2464 (O_2464,N_16920,N_16687);
nor UO_2465 (O_2465,N_19000,N_15649);
nor UO_2466 (O_2466,N_16561,N_18285);
nand UO_2467 (O_2467,N_18765,N_16336);
nand UO_2468 (O_2468,N_17571,N_16447);
xnor UO_2469 (O_2469,N_15882,N_18413);
and UO_2470 (O_2470,N_17535,N_18134);
or UO_2471 (O_2471,N_17590,N_19464);
or UO_2472 (O_2472,N_16118,N_15147);
and UO_2473 (O_2473,N_16848,N_17322);
nor UO_2474 (O_2474,N_15030,N_17813);
and UO_2475 (O_2475,N_16455,N_15354);
nand UO_2476 (O_2476,N_17446,N_15889);
or UO_2477 (O_2477,N_16932,N_17694);
and UO_2478 (O_2478,N_18272,N_18001);
or UO_2479 (O_2479,N_16470,N_15532);
nand UO_2480 (O_2480,N_17614,N_17100);
nand UO_2481 (O_2481,N_17775,N_18427);
xor UO_2482 (O_2482,N_19835,N_18352);
nor UO_2483 (O_2483,N_19224,N_19288);
xnor UO_2484 (O_2484,N_18253,N_19790);
nand UO_2485 (O_2485,N_16567,N_19722);
or UO_2486 (O_2486,N_19386,N_18267);
nor UO_2487 (O_2487,N_17162,N_16513);
and UO_2488 (O_2488,N_16300,N_17913);
and UO_2489 (O_2489,N_18936,N_17495);
and UO_2490 (O_2490,N_16579,N_15966);
or UO_2491 (O_2491,N_18745,N_15193);
nor UO_2492 (O_2492,N_16666,N_19976);
or UO_2493 (O_2493,N_19501,N_16593);
nor UO_2494 (O_2494,N_15896,N_18761);
and UO_2495 (O_2495,N_18779,N_18914);
or UO_2496 (O_2496,N_18337,N_16452);
nand UO_2497 (O_2497,N_16091,N_18642);
nor UO_2498 (O_2498,N_15995,N_17312);
nand UO_2499 (O_2499,N_15963,N_16333);
endmodule