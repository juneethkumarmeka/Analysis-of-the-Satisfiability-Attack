module basic_500_3000_500_40_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_383,In_144);
nor U1 (N_1,In_117,In_248);
xor U2 (N_2,In_293,In_56);
or U3 (N_3,In_187,In_235);
and U4 (N_4,In_23,In_53);
xor U5 (N_5,In_54,In_331);
nor U6 (N_6,In_20,In_364);
nand U7 (N_7,In_438,In_468);
nor U8 (N_8,In_406,In_34);
xor U9 (N_9,In_116,In_232);
and U10 (N_10,In_487,In_47);
or U11 (N_11,In_340,In_243);
nor U12 (N_12,In_211,In_407);
nand U13 (N_13,In_264,In_239);
and U14 (N_14,In_21,In_404);
nand U15 (N_15,In_63,In_473);
or U16 (N_16,In_50,In_332);
nor U17 (N_17,In_5,In_15);
or U18 (N_18,In_263,In_316);
nor U19 (N_19,In_206,In_95);
nand U20 (N_20,In_469,In_443);
or U21 (N_21,In_265,In_393);
nand U22 (N_22,In_382,In_164);
and U23 (N_23,In_376,In_268);
nor U24 (N_24,In_9,In_387);
or U25 (N_25,In_4,In_452);
and U26 (N_26,In_104,In_30);
nor U27 (N_27,In_202,In_292);
and U28 (N_28,In_167,In_346);
nand U29 (N_29,In_358,In_130);
or U30 (N_30,In_470,In_17);
nor U31 (N_31,In_299,In_223);
nor U32 (N_32,In_445,In_241);
or U33 (N_33,In_166,In_279);
nand U34 (N_34,In_363,In_408);
nand U35 (N_35,In_267,In_476);
or U36 (N_36,In_124,In_96);
nor U37 (N_37,In_188,In_399);
nor U38 (N_38,In_397,In_155);
xnor U39 (N_39,In_296,In_386);
or U40 (N_40,In_466,In_147);
or U41 (N_41,In_249,In_411);
nand U42 (N_42,In_24,In_234);
nor U43 (N_43,In_325,In_361);
and U44 (N_44,In_403,In_431);
nor U45 (N_45,In_495,In_127);
xor U46 (N_46,In_151,In_150);
xor U47 (N_47,In_143,In_118);
nor U48 (N_48,In_488,In_204);
and U49 (N_49,In_308,In_252);
nor U50 (N_50,In_351,In_61);
nor U51 (N_51,In_314,In_230);
nor U52 (N_52,In_297,In_149);
or U53 (N_53,In_245,In_425);
or U54 (N_54,In_214,In_44);
and U55 (N_55,In_240,In_375);
nor U56 (N_56,In_19,In_218);
or U57 (N_57,In_496,In_289);
nand U58 (N_58,In_137,In_13);
or U59 (N_59,In_76,In_79);
and U60 (N_60,In_162,In_210);
nor U61 (N_61,In_339,In_153);
nand U62 (N_62,In_25,In_298);
or U63 (N_63,In_57,In_335);
and U64 (N_64,In_189,In_48);
nor U65 (N_65,In_329,In_80);
nand U66 (N_66,In_420,In_78);
or U67 (N_67,In_8,In_284);
and U68 (N_68,In_379,In_456);
xor U69 (N_69,In_246,In_472);
nor U70 (N_70,In_269,In_108);
nor U71 (N_71,In_374,In_98);
nand U72 (N_72,In_471,In_126);
or U73 (N_73,In_287,In_280);
or U74 (N_74,In_122,In_457);
xnor U75 (N_75,In_312,N_29);
and U76 (N_76,In_353,N_11);
and U77 (N_77,In_109,In_486);
or U78 (N_78,In_40,In_221);
or U79 (N_79,N_9,In_326);
or U80 (N_80,In_302,In_238);
and U81 (N_81,In_177,In_207);
and U82 (N_82,In_318,In_89);
or U83 (N_83,In_391,In_401);
nor U84 (N_84,In_52,N_0);
and U85 (N_85,In_183,In_32);
nand U86 (N_86,In_58,In_338);
and U87 (N_87,In_424,In_36);
nor U88 (N_88,In_110,In_208);
and U89 (N_89,In_205,In_430);
nand U90 (N_90,In_303,In_444);
or U91 (N_91,N_57,In_484);
and U92 (N_92,In_286,In_134);
and U93 (N_93,In_306,In_1);
and U94 (N_94,In_259,In_491);
and U95 (N_95,In_184,N_70);
or U96 (N_96,In_45,In_291);
nor U97 (N_97,In_275,In_366);
and U98 (N_98,In_145,In_442);
xor U99 (N_99,N_59,N_15);
or U100 (N_100,In_454,In_344);
nor U101 (N_101,In_38,In_323);
nand U102 (N_102,In_405,In_136);
or U103 (N_103,In_428,In_451);
nand U104 (N_104,In_490,In_283);
and U105 (N_105,In_141,In_59);
or U106 (N_106,In_389,In_313);
or U107 (N_107,In_181,In_493);
or U108 (N_108,In_474,In_41);
and U109 (N_109,N_35,In_160);
or U110 (N_110,In_278,In_453);
xor U111 (N_111,In_435,In_138);
nor U112 (N_112,In_419,In_485);
or U113 (N_113,In_460,In_200);
nor U114 (N_114,In_394,N_17);
nor U115 (N_115,In_90,In_18);
or U116 (N_116,In_288,In_72);
and U117 (N_117,In_87,In_237);
or U118 (N_118,In_14,N_27);
and U119 (N_119,In_414,N_67);
nand U120 (N_120,In_274,In_311);
or U121 (N_121,In_295,In_43);
nand U122 (N_122,In_370,In_333);
and U123 (N_123,N_61,In_65);
or U124 (N_124,In_436,In_261);
or U125 (N_125,In_185,In_262);
or U126 (N_126,In_481,In_494);
nor U127 (N_127,N_73,In_254);
nand U128 (N_128,In_342,N_8);
or U129 (N_129,In_103,In_349);
and U130 (N_130,In_448,In_3);
and U131 (N_131,In_356,In_154);
nand U132 (N_132,In_133,In_480);
nand U133 (N_133,In_381,In_402);
or U134 (N_134,In_482,In_176);
xnor U135 (N_135,In_434,In_336);
nand U136 (N_136,In_31,In_27);
or U137 (N_137,In_132,In_173);
nand U138 (N_138,In_68,In_463);
and U139 (N_139,In_266,In_228);
nor U140 (N_140,In_368,In_139);
nand U141 (N_141,In_128,In_179);
nand U142 (N_142,In_307,In_146);
or U143 (N_143,In_180,In_123);
and U144 (N_144,N_14,In_37);
and U145 (N_145,In_74,In_92);
or U146 (N_146,In_464,In_22);
or U147 (N_147,In_450,In_385);
nor U148 (N_148,N_18,In_354);
nor U149 (N_149,In_193,In_71);
nand U150 (N_150,In_222,N_62);
nor U151 (N_151,N_146,In_330);
or U152 (N_152,N_130,In_158);
and U153 (N_153,N_2,N_81);
nand U154 (N_154,In_174,In_465);
nor U155 (N_155,N_142,In_119);
nand U156 (N_156,N_87,In_219);
nor U157 (N_157,In_461,In_350);
nor U158 (N_158,N_32,In_82);
xor U159 (N_159,In_301,N_105);
nand U160 (N_160,In_422,N_101);
nor U161 (N_161,In_337,N_91);
xor U162 (N_162,In_321,N_68);
and U163 (N_163,In_91,N_28);
nor U164 (N_164,N_138,In_449);
nand U165 (N_165,In_310,In_194);
and U166 (N_166,N_54,In_328);
and U167 (N_167,In_86,In_462);
nor U168 (N_168,In_26,N_93);
nor U169 (N_169,In_201,In_343);
nor U170 (N_170,In_140,N_79);
nand U171 (N_171,In_62,In_441);
xor U172 (N_172,N_50,In_131);
nor U173 (N_173,In_215,In_7);
or U174 (N_174,In_304,N_133);
nor U175 (N_175,N_124,In_395);
xnor U176 (N_176,N_117,In_384);
and U177 (N_177,In_300,In_69);
and U178 (N_178,N_84,N_136);
and U179 (N_179,N_98,In_172);
and U180 (N_180,In_135,N_49);
or U181 (N_181,N_33,In_429);
and U182 (N_182,In_273,N_149);
nor U183 (N_183,In_341,N_64);
or U184 (N_184,In_28,In_94);
or U185 (N_185,N_39,In_250);
and U186 (N_186,In_369,In_372);
or U187 (N_187,In_225,In_16);
or U188 (N_188,N_21,In_11);
and U189 (N_189,In_322,In_197);
nand U190 (N_190,N_66,In_352);
xnor U191 (N_191,In_73,In_55);
and U192 (N_192,N_114,N_112);
nand U193 (N_193,In_226,In_209);
and U194 (N_194,In_182,In_388);
xor U195 (N_195,In_51,N_147);
and U196 (N_196,N_108,N_16);
nand U197 (N_197,In_113,N_13);
and U198 (N_198,In_359,In_46);
or U199 (N_199,In_497,In_365);
and U200 (N_200,In_426,In_196);
xor U201 (N_201,N_45,In_255);
nand U202 (N_202,In_360,N_126);
nor U203 (N_203,N_24,In_244);
or U204 (N_204,In_270,In_165);
nand U205 (N_205,N_132,In_120);
and U206 (N_206,N_116,In_437);
and U207 (N_207,N_90,In_175);
and U208 (N_208,N_12,In_276);
nor U209 (N_209,In_392,In_492);
or U210 (N_210,N_80,N_74);
nor U211 (N_211,N_46,In_0);
and U212 (N_212,N_58,N_43);
or U213 (N_213,N_139,N_78);
nand U214 (N_214,In_271,In_12);
or U215 (N_215,N_100,In_373);
and U216 (N_216,In_439,N_145);
nor U217 (N_217,N_106,N_26);
nand U218 (N_218,In_75,In_446);
and U219 (N_219,N_53,In_77);
nor U220 (N_220,N_95,N_19);
or U221 (N_221,In_242,In_413);
nand U222 (N_222,In_229,N_115);
nand U223 (N_223,In_129,In_447);
or U224 (N_224,In_418,N_82);
or U225 (N_225,N_222,N_44);
nand U226 (N_226,In_290,N_71);
and U227 (N_227,In_224,N_191);
xnor U228 (N_228,In_67,In_467);
and U229 (N_229,In_217,In_168);
and U230 (N_230,N_144,N_162);
xor U231 (N_231,In_459,In_88);
and U232 (N_232,N_220,N_161);
and U233 (N_233,N_184,N_170);
nor U234 (N_234,N_107,N_76);
nor U235 (N_235,In_33,N_119);
nand U236 (N_236,In_440,In_216);
nand U237 (N_237,In_29,In_281);
xnor U238 (N_238,In_64,In_191);
nor U239 (N_239,In_192,N_206);
xor U240 (N_240,N_180,In_35);
and U241 (N_241,N_160,In_81);
or U242 (N_242,In_148,In_60);
or U243 (N_243,N_164,In_2);
or U244 (N_244,N_171,N_224);
nand U245 (N_245,In_121,In_114);
nand U246 (N_246,In_475,N_195);
nor U247 (N_247,In_417,In_294);
and U248 (N_248,N_199,N_196);
nand U249 (N_249,In_320,N_182);
xor U250 (N_250,N_77,N_131);
and U251 (N_251,In_421,In_49);
and U252 (N_252,N_113,N_159);
and U253 (N_253,N_173,In_499);
or U254 (N_254,In_285,N_75);
or U255 (N_255,In_112,In_236);
nor U256 (N_256,N_22,N_127);
nand U257 (N_257,N_34,In_315);
nand U258 (N_258,In_39,In_427);
or U259 (N_259,In_203,In_93);
and U260 (N_260,N_135,N_52);
or U261 (N_261,N_151,In_347);
and U262 (N_262,N_125,N_211);
xnor U263 (N_263,In_157,N_176);
xnor U264 (N_264,In_66,N_41);
or U265 (N_265,In_345,In_97);
nand U266 (N_266,N_109,In_309);
nand U267 (N_267,In_396,In_100);
or U268 (N_268,N_129,In_319);
and U269 (N_269,In_362,N_186);
nand U270 (N_270,N_85,In_260);
and U271 (N_271,N_157,N_204);
xnor U272 (N_272,In_231,In_101);
nand U273 (N_273,N_200,N_123);
xor U274 (N_274,In_455,N_179);
or U275 (N_275,In_458,N_201);
xor U276 (N_276,N_69,In_105);
and U277 (N_277,N_202,In_478);
nand U278 (N_278,N_166,N_193);
nand U279 (N_279,In_195,N_219);
nand U280 (N_280,In_398,N_187);
nor U281 (N_281,In_377,In_348);
or U282 (N_282,In_498,In_390);
and U283 (N_283,N_3,N_55);
xnor U284 (N_284,In_115,N_118);
and U285 (N_285,N_141,In_152);
nand U286 (N_286,N_192,N_42);
nor U287 (N_287,In_416,N_122);
nand U288 (N_288,N_209,N_23);
nand U289 (N_289,N_178,In_247);
nand U290 (N_290,In_102,N_172);
nand U291 (N_291,In_380,N_40);
and U292 (N_292,In_423,N_152);
and U293 (N_293,In_415,In_324);
or U294 (N_294,In_433,N_47);
or U295 (N_295,In_410,N_218);
or U296 (N_296,N_94,In_483);
nand U297 (N_297,N_104,In_169);
nor U298 (N_298,In_371,In_277);
or U299 (N_299,N_168,N_83);
and U300 (N_300,N_30,N_205);
and U301 (N_301,N_289,N_269);
and U302 (N_302,In_412,N_110);
nor U303 (N_303,N_298,In_357);
nand U304 (N_304,N_274,In_190);
nand U305 (N_305,N_213,N_270);
nor U306 (N_306,N_158,In_355);
or U307 (N_307,N_212,N_299);
and U308 (N_308,In_42,N_278);
nor U309 (N_309,N_245,N_150);
and U310 (N_310,In_272,N_89);
xnor U311 (N_311,In_111,In_233);
nor U312 (N_312,N_185,In_186);
xor U313 (N_313,In_258,In_432);
and U314 (N_314,In_212,N_153);
or U315 (N_315,In_198,N_283);
xor U316 (N_316,N_163,N_143);
and U317 (N_317,N_262,N_72);
xnor U318 (N_318,N_92,N_276);
and U319 (N_319,In_367,N_267);
and U320 (N_320,N_241,N_226);
or U321 (N_321,N_225,N_292);
xor U322 (N_322,N_174,In_477);
or U323 (N_323,In_171,N_148);
nor U324 (N_324,N_266,N_291);
xnor U325 (N_325,N_167,N_120);
nand U326 (N_326,N_154,In_479);
nand U327 (N_327,In_409,N_25);
and U328 (N_328,In_256,N_10);
or U329 (N_329,N_235,N_216);
nand U330 (N_330,In_10,In_327);
and U331 (N_331,N_121,N_254);
nor U332 (N_332,N_242,N_258);
nor U333 (N_333,N_51,N_128);
nand U334 (N_334,In_159,N_155);
or U335 (N_335,In_70,In_142);
xnor U336 (N_336,N_137,N_247);
and U337 (N_337,N_239,N_243);
nand U338 (N_338,N_257,In_257);
nor U339 (N_339,N_233,N_197);
or U340 (N_340,N_240,N_5);
nor U341 (N_341,N_111,In_107);
nor U342 (N_342,N_36,N_256);
and U343 (N_343,N_177,N_96);
and U344 (N_344,N_296,N_37);
or U345 (N_345,N_255,N_103);
or U346 (N_346,N_97,In_378);
xnor U347 (N_347,In_213,N_280);
or U348 (N_348,In_161,N_281);
nor U349 (N_349,N_229,N_4);
nor U350 (N_350,N_230,N_134);
nand U351 (N_351,N_214,In_85);
or U352 (N_352,N_210,N_287);
or U353 (N_353,N_252,In_83);
nand U354 (N_354,N_65,In_6);
xor U355 (N_355,In_106,N_234);
and U356 (N_356,N_286,N_265);
or U357 (N_357,In_227,N_275);
or U358 (N_358,In_334,N_223);
and U359 (N_359,N_190,N_288);
and U360 (N_360,N_237,N_188);
xnor U361 (N_361,N_181,N_246);
or U362 (N_362,N_175,N_273);
or U363 (N_363,In_317,N_249);
or U364 (N_364,N_86,N_284);
nor U365 (N_365,In_178,In_170);
and U366 (N_366,In_84,N_290);
nor U367 (N_367,N_285,In_305);
and U368 (N_368,N_293,N_268);
nand U369 (N_369,In_251,N_6);
or U370 (N_370,N_194,N_261);
nor U371 (N_371,In_220,N_221);
nor U372 (N_372,N_165,N_238);
or U373 (N_373,N_277,In_489);
xnor U374 (N_374,N_156,N_264);
nand U375 (N_375,N_329,N_373);
or U376 (N_376,N_309,N_341);
nand U377 (N_377,N_321,N_362);
and U378 (N_378,N_345,N_336);
and U379 (N_379,N_228,N_320);
or U380 (N_380,N_359,N_342);
nand U381 (N_381,N_232,N_349);
nand U382 (N_382,N_348,N_355);
or U383 (N_383,N_305,N_302);
and U384 (N_384,N_318,N_263);
nor U385 (N_385,N_260,N_323);
and U386 (N_386,N_20,N_282);
and U387 (N_387,N_227,N_358);
nand U388 (N_388,N_183,N_38);
and U389 (N_389,N_295,In_156);
and U390 (N_390,N_271,N_368);
or U391 (N_391,N_315,N_319);
nand U392 (N_392,In_282,N_328);
nor U393 (N_393,N_272,N_99);
xnor U394 (N_394,N_325,N_365);
nor U395 (N_395,N_340,N_364);
and U396 (N_396,N_253,N_331);
nand U397 (N_397,N_279,N_208);
nand U398 (N_398,N_140,N_169);
nor U399 (N_399,N_313,N_335);
xor U400 (N_400,N_250,N_317);
xnor U401 (N_401,N_48,N_346);
nor U402 (N_402,N_1,N_369);
or U403 (N_403,N_198,N_306);
or U404 (N_404,N_327,N_360);
and U405 (N_405,N_352,N_334);
and U406 (N_406,N_344,N_351);
nor U407 (N_407,In_99,N_310);
or U408 (N_408,N_338,N_316);
nand U409 (N_409,N_339,N_297);
nor U410 (N_410,N_372,N_374);
nor U411 (N_411,N_371,N_63);
or U412 (N_412,N_314,In_400);
and U413 (N_413,N_312,N_244);
or U414 (N_414,N_311,In_163);
nor U415 (N_415,N_354,In_253);
xnor U416 (N_416,N_294,In_125);
and U417 (N_417,N_236,N_56);
or U418 (N_418,N_353,N_301);
and U419 (N_419,N_343,In_199);
and U420 (N_420,N_60,N_203);
or U421 (N_421,N_217,N_102);
nor U422 (N_422,N_215,N_307);
nor U423 (N_423,N_300,N_303);
nand U424 (N_424,N_259,N_248);
and U425 (N_425,N_350,N_357);
or U426 (N_426,N_370,N_31);
nor U427 (N_427,N_308,N_330);
or U428 (N_428,N_363,N_347);
nor U429 (N_429,N_324,N_7);
and U430 (N_430,N_251,N_207);
and U431 (N_431,N_322,N_361);
or U432 (N_432,N_332,N_333);
nor U433 (N_433,N_231,N_88);
and U434 (N_434,N_356,N_304);
xnor U435 (N_435,N_326,N_189);
or U436 (N_436,N_366,N_367);
or U437 (N_437,N_337,N_99);
xor U438 (N_438,N_307,N_297);
nor U439 (N_439,N_363,N_362);
nand U440 (N_440,In_163,N_324);
and U441 (N_441,N_311,N_366);
nand U442 (N_442,N_294,N_369);
and U443 (N_443,N_198,N_7);
and U444 (N_444,N_358,N_369);
xor U445 (N_445,N_294,N_259);
nand U446 (N_446,N_208,N_353);
nand U447 (N_447,N_48,N_251);
or U448 (N_448,N_367,N_349);
nand U449 (N_449,N_317,N_351);
nand U450 (N_450,N_420,N_391);
nor U451 (N_451,N_429,N_417);
and U452 (N_452,N_407,N_442);
nand U453 (N_453,N_439,N_428);
and U454 (N_454,N_403,N_376);
and U455 (N_455,N_430,N_432);
and U456 (N_456,N_418,N_382);
nor U457 (N_457,N_427,N_408);
or U458 (N_458,N_434,N_393);
nand U459 (N_459,N_413,N_416);
xor U460 (N_460,N_435,N_443);
xor U461 (N_461,N_402,N_381);
nor U462 (N_462,N_387,N_383);
nand U463 (N_463,N_385,N_409);
nor U464 (N_464,N_410,N_404);
nor U465 (N_465,N_438,N_448);
nor U466 (N_466,N_419,N_394);
xnor U467 (N_467,N_398,N_433);
nand U468 (N_468,N_379,N_378);
nand U469 (N_469,N_380,N_395);
or U470 (N_470,N_406,N_400);
and U471 (N_471,N_377,N_401);
and U472 (N_472,N_446,N_386);
and U473 (N_473,N_424,N_375);
nor U474 (N_474,N_426,N_449);
nor U475 (N_475,N_414,N_445);
or U476 (N_476,N_396,N_384);
nor U477 (N_477,N_405,N_425);
nor U478 (N_478,N_392,N_412);
or U479 (N_479,N_411,N_431);
xnor U480 (N_480,N_390,N_440);
nand U481 (N_481,N_389,N_444);
nand U482 (N_482,N_415,N_399);
and U483 (N_483,N_436,N_422);
and U484 (N_484,N_441,N_421);
and U485 (N_485,N_397,N_388);
nor U486 (N_486,N_423,N_437);
nand U487 (N_487,N_447,N_395);
or U488 (N_488,N_376,N_412);
nor U489 (N_489,N_397,N_442);
nor U490 (N_490,N_436,N_392);
nor U491 (N_491,N_411,N_401);
or U492 (N_492,N_426,N_445);
nor U493 (N_493,N_407,N_417);
nor U494 (N_494,N_424,N_400);
nand U495 (N_495,N_382,N_394);
and U496 (N_496,N_416,N_409);
nor U497 (N_497,N_398,N_385);
nor U498 (N_498,N_380,N_403);
nor U499 (N_499,N_447,N_382);
or U500 (N_500,N_425,N_447);
and U501 (N_501,N_390,N_381);
nand U502 (N_502,N_435,N_431);
xor U503 (N_503,N_382,N_431);
nor U504 (N_504,N_421,N_411);
and U505 (N_505,N_391,N_444);
nor U506 (N_506,N_376,N_432);
or U507 (N_507,N_430,N_421);
nand U508 (N_508,N_397,N_401);
nor U509 (N_509,N_434,N_431);
nand U510 (N_510,N_447,N_448);
and U511 (N_511,N_432,N_390);
nor U512 (N_512,N_440,N_447);
nor U513 (N_513,N_435,N_427);
and U514 (N_514,N_412,N_403);
nand U515 (N_515,N_380,N_416);
nor U516 (N_516,N_393,N_423);
nor U517 (N_517,N_393,N_446);
and U518 (N_518,N_403,N_422);
nand U519 (N_519,N_375,N_414);
nand U520 (N_520,N_416,N_376);
nor U521 (N_521,N_395,N_442);
and U522 (N_522,N_430,N_412);
or U523 (N_523,N_427,N_415);
nand U524 (N_524,N_438,N_443);
and U525 (N_525,N_480,N_451);
xor U526 (N_526,N_500,N_477);
and U527 (N_527,N_514,N_486);
or U528 (N_528,N_518,N_517);
nand U529 (N_529,N_457,N_495);
nor U530 (N_530,N_478,N_505);
or U531 (N_531,N_519,N_515);
and U532 (N_532,N_521,N_453);
xnor U533 (N_533,N_493,N_456);
nor U534 (N_534,N_501,N_504);
and U535 (N_535,N_474,N_462);
nand U536 (N_536,N_455,N_491);
nor U537 (N_537,N_499,N_485);
nor U538 (N_538,N_470,N_475);
or U539 (N_539,N_497,N_516);
nand U540 (N_540,N_492,N_520);
xor U541 (N_541,N_502,N_513);
and U542 (N_542,N_461,N_490);
or U543 (N_543,N_508,N_494);
xor U544 (N_544,N_503,N_496);
nand U545 (N_545,N_481,N_512);
or U546 (N_546,N_522,N_471);
or U547 (N_547,N_507,N_487);
nor U548 (N_548,N_450,N_510);
or U549 (N_549,N_464,N_466);
nand U550 (N_550,N_459,N_473);
or U551 (N_551,N_460,N_498);
nand U552 (N_552,N_511,N_479);
nand U553 (N_553,N_506,N_458);
and U554 (N_554,N_488,N_465);
and U555 (N_555,N_463,N_523);
and U556 (N_556,N_476,N_489);
or U557 (N_557,N_524,N_484);
nand U558 (N_558,N_469,N_454);
or U559 (N_559,N_452,N_467);
xor U560 (N_560,N_468,N_472);
nor U561 (N_561,N_482,N_483);
nand U562 (N_562,N_509,N_486);
or U563 (N_563,N_465,N_460);
xor U564 (N_564,N_473,N_511);
or U565 (N_565,N_462,N_451);
or U566 (N_566,N_503,N_498);
and U567 (N_567,N_497,N_493);
and U568 (N_568,N_468,N_517);
or U569 (N_569,N_490,N_498);
nor U570 (N_570,N_459,N_474);
and U571 (N_571,N_507,N_471);
and U572 (N_572,N_507,N_473);
nor U573 (N_573,N_502,N_520);
or U574 (N_574,N_509,N_466);
xor U575 (N_575,N_505,N_451);
nor U576 (N_576,N_476,N_470);
nor U577 (N_577,N_510,N_480);
nand U578 (N_578,N_455,N_516);
or U579 (N_579,N_483,N_474);
or U580 (N_580,N_515,N_518);
nand U581 (N_581,N_451,N_523);
nor U582 (N_582,N_490,N_460);
nand U583 (N_583,N_510,N_514);
nor U584 (N_584,N_450,N_452);
nor U585 (N_585,N_512,N_496);
or U586 (N_586,N_476,N_493);
nand U587 (N_587,N_466,N_478);
or U588 (N_588,N_483,N_499);
xor U589 (N_589,N_488,N_512);
or U590 (N_590,N_503,N_477);
nand U591 (N_591,N_457,N_517);
nor U592 (N_592,N_500,N_451);
nand U593 (N_593,N_450,N_518);
or U594 (N_594,N_480,N_490);
or U595 (N_595,N_491,N_472);
and U596 (N_596,N_490,N_458);
xor U597 (N_597,N_509,N_517);
or U598 (N_598,N_524,N_466);
nand U599 (N_599,N_454,N_514);
nor U600 (N_600,N_539,N_583);
nor U601 (N_601,N_548,N_532);
and U602 (N_602,N_545,N_558);
nand U603 (N_603,N_550,N_572);
nor U604 (N_604,N_597,N_538);
nand U605 (N_605,N_540,N_593);
and U606 (N_606,N_531,N_595);
nor U607 (N_607,N_575,N_533);
nor U608 (N_608,N_567,N_571);
xor U609 (N_609,N_586,N_525);
and U610 (N_610,N_544,N_546);
nand U611 (N_611,N_592,N_552);
nand U612 (N_612,N_594,N_581);
and U613 (N_613,N_557,N_561);
nand U614 (N_614,N_589,N_537);
and U615 (N_615,N_591,N_536);
nor U616 (N_616,N_562,N_553);
xnor U617 (N_617,N_578,N_590);
or U618 (N_618,N_535,N_574);
nand U619 (N_619,N_543,N_547);
xnor U620 (N_620,N_527,N_570);
nor U621 (N_621,N_573,N_587);
nand U622 (N_622,N_598,N_534);
nand U623 (N_623,N_564,N_599);
nor U624 (N_624,N_588,N_528);
and U625 (N_625,N_529,N_577);
nand U626 (N_626,N_554,N_556);
xor U627 (N_627,N_580,N_555);
nand U628 (N_628,N_551,N_566);
nor U629 (N_629,N_526,N_596);
or U630 (N_630,N_579,N_563);
and U631 (N_631,N_530,N_542);
or U632 (N_632,N_549,N_584);
or U633 (N_633,N_585,N_569);
and U634 (N_634,N_541,N_560);
nor U635 (N_635,N_565,N_582);
or U636 (N_636,N_559,N_576);
and U637 (N_637,N_568,N_591);
and U638 (N_638,N_547,N_562);
nor U639 (N_639,N_558,N_585);
nor U640 (N_640,N_558,N_596);
and U641 (N_641,N_551,N_593);
xor U642 (N_642,N_527,N_556);
nand U643 (N_643,N_525,N_546);
xnor U644 (N_644,N_546,N_587);
and U645 (N_645,N_526,N_533);
nor U646 (N_646,N_530,N_583);
or U647 (N_647,N_557,N_590);
or U648 (N_648,N_591,N_565);
nand U649 (N_649,N_537,N_560);
or U650 (N_650,N_525,N_536);
nor U651 (N_651,N_571,N_542);
nor U652 (N_652,N_554,N_533);
nor U653 (N_653,N_582,N_539);
and U654 (N_654,N_579,N_552);
or U655 (N_655,N_562,N_578);
nor U656 (N_656,N_555,N_576);
nor U657 (N_657,N_581,N_527);
and U658 (N_658,N_586,N_553);
and U659 (N_659,N_528,N_585);
or U660 (N_660,N_537,N_567);
nor U661 (N_661,N_546,N_545);
and U662 (N_662,N_529,N_599);
nand U663 (N_663,N_599,N_583);
nor U664 (N_664,N_541,N_586);
or U665 (N_665,N_534,N_540);
and U666 (N_666,N_544,N_588);
or U667 (N_667,N_555,N_530);
nor U668 (N_668,N_541,N_557);
or U669 (N_669,N_579,N_587);
or U670 (N_670,N_566,N_574);
and U671 (N_671,N_558,N_598);
or U672 (N_672,N_569,N_567);
xnor U673 (N_673,N_543,N_590);
and U674 (N_674,N_581,N_571);
nand U675 (N_675,N_637,N_618);
xnor U676 (N_676,N_662,N_653);
or U677 (N_677,N_639,N_630);
or U678 (N_678,N_612,N_671);
xor U679 (N_679,N_619,N_665);
or U680 (N_680,N_627,N_650);
and U681 (N_681,N_607,N_615);
or U682 (N_682,N_644,N_669);
xor U683 (N_683,N_658,N_666);
or U684 (N_684,N_640,N_614);
nand U685 (N_685,N_624,N_617);
or U686 (N_686,N_655,N_672);
or U687 (N_687,N_636,N_674);
nor U688 (N_688,N_664,N_654);
nor U689 (N_689,N_651,N_620);
and U690 (N_690,N_648,N_652);
nand U691 (N_691,N_668,N_656);
nor U692 (N_692,N_659,N_609);
and U693 (N_693,N_638,N_605);
nand U694 (N_694,N_645,N_642);
or U695 (N_695,N_616,N_673);
nand U696 (N_696,N_600,N_629);
xnor U697 (N_697,N_663,N_626);
nand U698 (N_698,N_660,N_667);
and U699 (N_699,N_631,N_601);
and U700 (N_700,N_625,N_643);
or U701 (N_701,N_610,N_649);
or U702 (N_702,N_622,N_670);
and U703 (N_703,N_635,N_634);
nand U704 (N_704,N_611,N_647);
nor U705 (N_705,N_606,N_602);
nand U706 (N_706,N_633,N_613);
nand U707 (N_707,N_641,N_661);
and U708 (N_708,N_603,N_621);
or U709 (N_709,N_632,N_623);
or U710 (N_710,N_657,N_628);
or U711 (N_711,N_646,N_608);
xnor U712 (N_712,N_604,N_657);
and U713 (N_713,N_636,N_667);
or U714 (N_714,N_672,N_632);
nor U715 (N_715,N_651,N_674);
or U716 (N_716,N_639,N_620);
nand U717 (N_717,N_668,N_653);
xnor U718 (N_718,N_666,N_669);
nor U719 (N_719,N_654,N_606);
nor U720 (N_720,N_614,N_633);
and U721 (N_721,N_635,N_653);
xor U722 (N_722,N_628,N_616);
nand U723 (N_723,N_648,N_630);
nor U724 (N_724,N_642,N_612);
nand U725 (N_725,N_636,N_634);
and U726 (N_726,N_661,N_634);
xnor U727 (N_727,N_649,N_609);
and U728 (N_728,N_648,N_610);
nor U729 (N_729,N_613,N_660);
nor U730 (N_730,N_643,N_658);
or U731 (N_731,N_639,N_606);
xnor U732 (N_732,N_636,N_657);
xor U733 (N_733,N_607,N_642);
nand U734 (N_734,N_629,N_633);
nand U735 (N_735,N_613,N_657);
xor U736 (N_736,N_607,N_638);
xnor U737 (N_737,N_641,N_649);
and U738 (N_738,N_642,N_622);
nor U739 (N_739,N_611,N_609);
or U740 (N_740,N_622,N_617);
or U741 (N_741,N_666,N_605);
or U742 (N_742,N_673,N_652);
and U743 (N_743,N_620,N_662);
nor U744 (N_744,N_674,N_626);
or U745 (N_745,N_630,N_626);
nand U746 (N_746,N_662,N_659);
nor U747 (N_747,N_670,N_630);
and U748 (N_748,N_660,N_615);
and U749 (N_749,N_660,N_662);
or U750 (N_750,N_740,N_702);
and U751 (N_751,N_719,N_744);
nand U752 (N_752,N_696,N_742);
nor U753 (N_753,N_720,N_710);
nor U754 (N_754,N_717,N_686);
nand U755 (N_755,N_681,N_743);
nand U756 (N_756,N_722,N_749);
nand U757 (N_757,N_746,N_676);
or U758 (N_758,N_731,N_690);
nand U759 (N_759,N_689,N_725);
xor U760 (N_760,N_695,N_704);
nand U761 (N_761,N_716,N_739);
and U762 (N_762,N_692,N_687);
nor U763 (N_763,N_693,N_707);
or U764 (N_764,N_698,N_713);
xor U765 (N_765,N_714,N_684);
or U766 (N_766,N_705,N_691);
and U767 (N_767,N_706,N_747);
and U768 (N_768,N_721,N_732);
nand U769 (N_769,N_748,N_745);
nor U770 (N_770,N_735,N_701);
nor U771 (N_771,N_712,N_715);
or U772 (N_772,N_697,N_736);
nor U773 (N_773,N_699,N_730);
nor U774 (N_774,N_679,N_677);
xor U775 (N_775,N_682,N_683);
nor U776 (N_776,N_708,N_685);
nand U777 (N_777,N_738,N_680);
nor U778 (N_778,N_741,N_727);
nand U779 (N_779,N_729,N_737);
nor U780 (N_780,N_723,N_728);
and U781 (N_781,N_694,N_726);
or U782 (N_782,N_703,N_733);
or U783 (N_783,N_724,N_678);
and U784 (N_784,N_718,N_709);
nand U785 (N_785,N_700,N_734);
nor U786 (N_786,N_688,N_675);
xnor U787 (N_787,N_711,N_701);
nand U788 (N_788,N_705,N_683);
or U789 (N_789,N_716,N_717);
nor U790 (N_790,N_734,N_710);
and U791 (N_791,N_701,N_707);
nand U792 (N_792,N_716,N_706);
or U793 (N_793,N_702,N_685);
xnor U794 (N_794,N_684,N_679);
nor U795 (N_795,N_698,N_706);
and U796 (N_796,N_687,N_748);
and U797 (N_797,N_727,N_686);
nand U798 (N_798,N_692,N_749);
or U799 (N_799,N_705,N_724);
nand U800 (N_800,N_731,N_736);
nor U801 (N_801,N_681,N_719);
and U802 (N_802,N_701,N_733);
and U803 (N_803,N_747,N_677);
and U804 (N_804,N_715,N_687);
nor U805 (N_805,N_737,N_716);
or U806 (N_806,N_732,N_675);
nor U807 (N_807,N_722,N_707);
nand U808 (N_808,N_689,N_735);
nor U809 (N_809,N_702,N_707);
nand U810 (N_810,N_717,N_737);
nand U811 (N_811,N_689,N_704);
or U812 (N_812,N_742,N_681);
nand U813 (N_813,N_688,N_710);
nor U814 (N_814,N_696,N_679);
xor U815 (N_815,N_695,N_741);
nand U816 (N_816,N_746,N_694);
nand U817 (N_817,N_684,N_701);
or U818 (N_818,N_675,N_696);
nand U819 (N_819,N_738,N_746);
nand U820 (N_820,N_704,N_694);
nand U821 (N_821,N_738,N_711);
nand U822 (N_822,N_725,N_732);
nor U823 (N_823,N_730,N_696);
xor U824 (N_824,N_683,N_679);
or U825 (N_825,N_809,N_751);
or U826 (N_826,N_770,N_763);
nor U827 (N_827,N_777,N_756);
and U828 (N_828,N_766,N_765);
and U829 (N_829,N_816,N_820);
and U830 (N_830,N_805,N_788);
nand U831 (N_831,N_771,N_782);
and U832 (N_832,N_755,N_772);
and U833 (N_833,N_779,N_787);
nand U834 (N_834,N_790,N_802);
and U835 (N_835,N_759,N_800);
and U836 (N_836,N_821,N_753);
and U837 (N_837,N_808,N_822);
xnor U838 (N_838,N_791,N_781);
xor U839 (N_839,N_794,N_793);
and U840 (N_840,N_769,N_807);
and U841 (N_841,N_798,N_778);
and U842 (N_842,N_811,N_762);
nor U843 (N_843,N_789,N_796);
and U844 (N_844,N_824,N_815);
nor U845 (N_845,N_786,N_774);
nor U846 (N_846,N_799,N_784);
xor U847 (N_847,N_819,N_773);
or U848 (N_848,N_823,N_783);
xnor U849 (N_849,N_785,N_810);
nand U850 (N_850,N_754,N_752);
nor U851 (N_851,N_757,N_814);
nor U852 (N_852,N_801,N_813);
or U853 (N_853,N_812,N_780);
xor U854 (N_854,N_804,N_768);
xnor U855 (N_855,N_795,N_775);
nand U856 (N_856,N_761,N_767);
or U857 (N_857,N_764,N_758);
nor U858 (N_858,N_792,N_760);
nand U859 (N_859,N_803,N_817);
nand U860 (N_860,N_818,N_797);
nand U861 (N_861,N_750,N_776);
xnor U862 (N_862,N_806,N_807);
or U863 (N_863,N_823,N_769);
and U864 (N_864,N_793,N_808);
and U865 (N_865,N_751,N_779);
nor U866 (N_866,N_803,N_751);
and U867 (N_867,N_784,N_786);
and U868 (N_868,N_767,N_772);
or U869 (N_869,N_760,N_772);
nor U870 (N_870,N_802,N_766);
or U871 (N_871,N_754,N_780);
xor U872 (N_872,N_780,N_757);
xnor U873 (N_873,N_780,N_766);
nand U874 (N_874,N_818,N_762);
nor U875 (N_875,N_774,N_821);
or U876 (N_876,N_772,N_759);
nand U877 (N_877,N_813,N_783);
or U878 (N_878,N_807,N_765);
or U879 (N_879,N_776,N_824);
or U880 (N_880,N_753,N_758);
or U881 (N_881,N_799,N_790);
and U882 (N_882,N_759,N_819);
or U883 (N_883,N_778,N_776);
nand U884 (N_884,N_788,N_777);
nor U885 (N_885,N_754,N_804);
and U886 (N_886,N_776,N_765);
nand U887 (N_887,N_779,N_758);
or U888 (N_888,N_784,N_797);
nand U889 (N_889,N_778,N_811);
nand U890 (N_890,N_754,N_770);
and U891 (N_891,N_797,N_778);
or U892 (N_892,N_760,N_750);
xnor U893 (N_893,N_802,N_775);
and U894 (N_894,N_752,N_771);
xor U895 (N_895,N_805,N_777);
or U896 (N_896,N_763,N_807);
or U897 (N_897,N_799,N_802);
and U898 (N_898,N_750,N_790);
or U899 (N_899,N_801,N_817);
xor U900 (N_900,N_864,N_878);
nand U901 (N_901,N_879,N_830);
nand U902 (N_902,N_860,N_854);
nand U903 (N_903,N_861,N_836);
nor U904 (N_904,N_898,N_849);
nor U905 (N_905,N_871,N_850);
nor U906 (N_906,N_856,N_876);
nor U907 (N_907,N_839,N_843);
nand U908 (N_908,N_825,N_887);
and U909 (N_909,N_838,N_847);
xor U910 (N_910,N_828,N_881);
xnor U911 (N_911,N_851,N_870);
nor U912 (N_912,N_873,N_855);
and U913 (N_913,N_895,N_865);
or U914 (N_914,N_833,N_834);
or U915 (N_915,N_837,N_884);
and U916 (N_916,N_882,N_826);
nor U917 (N_917,N_889,N_852);
nand U918 (N_918,N_899,N_892);
nand U919 (N_919,N_875,N_853);
nor U920 (N_920,N_829,N_848);
and U921 (N_921,N_840,N_894);
nor U922 (N_922,N_886,N_883);
nand U923 (N_923,N_832,N_858);
nand U924 (N_924,N_857,N_874);
nor U925 (N_925,N_845,N_859);
nand U926 (N_926,N_897,N_835);
xor U927 (N_927,N_869,N_863);
or U928 (N_928,N_841,N_893);
nor U929 (N_929,N_891,N_844);
xor U930 (N_930,N_827,N_877);
xor U931 (N_931,N_896,N_888);
and U932 (N_932,N_890,N_831);
nor U933 (N_933,N_880,N_846);
and U934 (N_934,N_862,N_866);
or U935 (N_935,N_842,N_872);
xnor U936 (N_936,N_867,N_885);
nor U937 (N_937,N_868,N_844);
or U938 (N_938,N_896,N_863);
and U939 (N_939,N_843,N_834);
or U940 (N_940,N_833,N_860);
nand U941 (N_941,N_873,N_856);
or U942 (N_942,N_883,N_898);
or U943 (N_943,N_831,N_837);
nand U944 (N_944,N_832,N_857);
or U945 (N_945,N_874,N_826);
nand U946 (N_946,N_881,N_893);
or U947 (N_947,N_843,N_871);
nor U948 (N_948,N_897,N_886);
and U949 (N_949,N_852,N_857);
or U950 (N_950,N_851,N_887);
or U951 (N_951,N_832,N_834);
nand U952 (N_952,N_883,N_875);
nor U953 (N_953,N_874,N_839);
nor U954 (N_954,N_854,N_868);
nand U955 (N_955,N_888,N_842);
or U956 (N_956,N_875,N_852);
or U957 (N_957,N_827,N_878);
nor U958 (N_958,N_880,N_871);
and U959 (N_959,N_863,N_866);
xor U960 (N_960,N_837,N_897);
nor U961 (N_961,N_840,N_893);
nand U962 (N_962,N_840,N_827);
or U963 (N_963,N_886,N_825);
nor U964 (N_964,N_833,N_886);
or U965 (N_965,N_850,N_842);
nand U966 (N_966,N_848,N_853);
or U967 (N_967,N_888,N_876);
xor U968 (N_968,N_898,N_885);
xor U969 (N_969,N_852,N_860);
nand U970 (N_970,N_857,N_845);
and U971 (N_971,N_870,N_875);
nor U972 (N_972,N_895,N_859);
and U973 (N_973,N_891,N_861);
or U974 (N_974,N_843,N_830);
nand U975 (N_975,N_966,N_918);
nor U976 (N_976,N_943,N_922);
or U977 (N_977,N_926,N_965);
nand U978 (N_978,N_919,N_913);
and U979 (N_979,N_900,N_954);
nor U980 (N_980,N_931,N_909);
or U981 (N_981,N_935,N_948);
nor U982 (N_982,N_934,N_970);
nand U983 (N_983,N_925,N_944);
or U984 (N_984,N_914,N_920);
or U985 (N_985,N_967,N_937);
and U986 (N_986,N_950,N_928);
nor U987 (N_987,N_947,N_964);
or U988 (N_988,N_930,N_908);
nand U989 (N_989,N_969,N_916);
nor U990 (N_990,N_904,N_924);
or U991 (N_991,N_961,N_907);
or U992 (N_992,N_945,N_973);
or U993 (N_993,N_959,N_915);
and U994 (N_994,N_910,N_941);
nand U995 (N_995,N_956,N_936);
or U996 (N_996,N_952,N_933);
and U997 (N_997,N_911,N_901);
xnor U998 (N_998,N_921,N_957);
nand U999 (N_999,N_939,N_912);
and U1000 (N_1000,N_903,N_932);
and U1001 (N_1001,N_951,N_972);
xor U1002 (N_1002,N_923,N_958);
or U1003 (N_1003,N_906,N_938);
or U1004 (N_1004,N_902,N_962);
nor U1005 (N_1005,N_974,N_917);
xor U1006 (N_1006,N_929,N_971);
nand U1007 (N_1007,N_940,N_949);
and U1008 (N_1008,N_953,N_963);
or U1009 (N_1009,N_968,N_955);
nand U1010 (N_1010,N_960,N_942);
xor U1011 (N_1011,N_946,N_905);
and U1012 (N_1012,N_927,N_947);
and U1013 (N_1013,N_963,N_954);
nand U1014 (N_1014,N_902,N_958);
nor U1015 (N_1015,N_958,N_935);
or U1016 (N_1016,N_929,N_909);
and U1017 (N_1017,N_974,N_951);
and U1018 (N_1018,N_956,N_925);
nor U1019 (N_1019,N_940,N_923);
xor U1020 (N_1020,N_932,N_943);
or U1021 (N_1021,N_914,N_974);
and U1022 (N_1022,N_947,N_944);
nand U1023 (N_1023,N_964,N_944);
nor U1024 (N_1024,N_905,N_900);
and U1025 (N_1025,N_910,N_973);
nand U1026 (N_1026,N_906,N_901);
and U1027 (N_1027,N_926,N_930);
nand U1028 (N_1028,N_907,N_951);
and U1029 (N_1029,N_958,N_915);
and U1030 (N_1030,N_941,N_938);
nand U1031 (N_1031,N_902,N_960);
nor U1032 (N_1032,N_960,N_934);
nand U1033 (N_1033,N_944,N_941);
and U1034 (N_1034,N_944,N_970);
xor U1035 (N_1035,N_968,N_901);
nand U1036 (N_1036,N_906,N_950);
or U1037 (N_1037,N_935,N_923);
xor U1038 (N_1038,N_910,N_907);
nor U1039 (N_1039,N_937,N_972);
nor U1040 (N_1040,N_921,N_930);
nand U1041 (N_1041,N_954,N_971);
nor U1042 (N_1042,N_907,N_903);
nand U1043 (N_1043,N_914,N_910);
and U1044 (N_1044,N_964,N_948);
nand U1045 (N_1045,N_945,N_951);
nor U1046 (N_1046,N_939,N_900);
or U1047 (N_1047,N_916,N_900);
nor U1048 (N_1048,N_908,N_905);
and U1049 (N_1049,N_924,N_950);
nand U1050 (N_1050,N_976,N_1031);
or U1051 (N_1051,N_975,N_1008);
and U1052 (N_1052,N_1036,N_1026);
or U1053 (N_1053,N_987,N_1018);
or U1054 (N_1054,N_978,N_986);
and U1055 (N_1055,N_1046,N_1019);
xor U1056 (N_1056,N_1038,N_1027);
or U1057 (N_1057,N_1045,N_1035);
and U1058 (N_1058,N_1015,N_1042);
and U1059 (N_1059,N_1032,N_1005);
nor U1060 (N_1060,N_1044,N_1020);
and U1061 (N_1061,N_1013,N_995);
nor U1062 (N_1062,N_1010,N_1041);
or U1063 (N_1063,N_1033,N_1011);
nand U1064 (N_1064,N_989,N_1012);
and U1065 (N_1065,N_990,N_1022);
or U1066 (N_1066,N_1034,N_1028);
nor U1067 (N_1067,N_988,N_977);
or U1068 (N_1068,N_1023,N_1049);
nor U1069 (N_1069,N_1039,N_993);
or U1070 (N_1070,N_1014,N_982);
nor U1071 (N_1071,N_984,N_1017);
nor U1072 (N_1072,N_1043,N_1025);
xnor U1073 (N_1073,N_998,N_981);
or U1074 (N_1074,N_1016,N_999);
nor U1075 (N_1075,N_1000,N_1002);
and U1076 (N_1076,N_1040,N_1004);
xnor U1077 (N_1077,N_992,N_1009);
nand U1078 (N_1078,N_1021,N_1001);
nor U1079 (N_1079,N_1007,N_979);
nand U1080 (N_1080,N_994,N_1030);
nor U1081 (N_1081,N_983,N_1024);
or U1082 (N_1082,N_1047,N_996);
and U1083 (N_1083,N_991,N_980);
or U1084 (N_1084,N_1048,N_997);
or U1085 (N_1085,N_985,N_1003);
nand U1086 (N_1086,N_1006,N_1029);
nand U1087 (N_1087,N_1037,N_1010);
nand U1088 (N_1088,N_1008,N_1033);
nand U1089 (N_1089,N_1033,N_996);
and U1090 (N_1090,N_993,N_1009);
or U1091 (N_1091,N_980,N_1004);
nor U1092 (N_1092,N_998,N_1005);
or U1093 (N_1093,N_1011,N_1039);
and U1094 (N_1094,N_1013,N_1046);
or U1095 (N_1095,N_1023,N_981);
or U1096 (N_1096,N_1020,N_1011);
or U1097 (N_1097,N_977,N_1017);
nor U1098 (N_1098,N_1031,N_993);
and U1099 (N_1099,N_1035,N_1013);
and U1100 (N_1100,N_1007,N_1019);
and U1101 (N_1101,N_990,N_1004);
or U1102 (N_1102,N_1015,N_1031);
or U1103 (N_1103,N_1006,N_1035);
or U1104 (N_1104,N_987,N_1034);
and U1105 (N_1105,N_1006,N_1011);
and U1106 (N_1106,N_1028,N_1005);
nor U1107 (N_1107,N_1040,N_1038);
nor U1108 (N_1108,N_1012,N_1034);
or U1109 (N_1109,N_986,N_980);
nor U1110 (N_1110,N_1023,N_1021);
nand U1111 (N_1111,N_1001,N_991);
nor U1112 (N_1112,N_1007,N_990);
or U1113 (N_1113,N_1000,N_1018);
nand U1114 (N_1114,N_1009,N_991);
nor U1115 (N_1115,N_1019,N_1005);
or U1116 (N_1116,N_1049,N_1032);
or U1117 (N_1117,N_1001,N_1007);
and U1118 (N_1118,N_989,N_1032);
or U1119 (N_1119,N_1035,N_1033);
nand U1120 (N_1120,N_1006,N_984);
nor U1121 (N_1121,N_997,N_1035);
and U1122 (N_1122,N_1027,N_1040);
and U1123 (N_1123,N_1008,N_976);
nand U1124 (N_1124,N_984,N_1030);
nor U1125 (N_1125,N_1119,N_1066);
nor U1126 (N_1126,N_1081,N_1121);
nand U1127 (N_1127,N_1059,N_1083);
nor U1128 (N_1128,N_1087,N_1072);
nor U1129 (N_1129,N_1101,N_1055);
xor U1130 (N_1130,N_1063,N_1099);
nand U1131 (N_1131,N_1096,N_1124);
nand U1132 (N_1132,N_1080,N_1118);
and U1133 (N_1133,N_1060,N_1076);
nand U1134 (N_1134,N_1095,N_1104);
nor U1135 (N_1135,N_1106,N_1088);
and U1136 (N_1136,N_1093,N_1057);
xor U1137 (N_1137,N_1082,N_1054);
nand U1138 (N_1138,N_1111,N_1079);
or U1139 (N_1139,N_1123,N_1061);
or U1140 (N_1140,N_1073,N_1103);
xnor U1141 (N_1141,N_1108,N_1091);
nor U1142 (N_1142,N_1089,N_1056);
nor U1143 (N_1143,N_1086,N_1051);
nand U1144 (N_1144,N_1090,N_1058);
and U1145 (N_1145,N_1052,N_1120);
nand U1146 (N_1146,N_1085,N_1065);
nand U1147 (N_1147,N_1114,N_1077);
nand U1148 (N_1148,N_1074,N_1094);
nor U1149 (N_1149,N_1071,N_1062);
or U1150 (N_1150,N_1068,N_1107);
or U1151 (N_1151,N_1067,N_1069);
and U1152 (N_1152,N_1064,N_1092);
nand U1153 (N_1153,N_1050,N_1117);
nor U1154 (N_1154,N_1078,N_1102);
nor U1155 (N_1155,N_1105,N_1053);
and U1156 (N_1156,N_1122,N_1112);
and U1157 (N_1157,N_1110,N_1113);
nand U1158 (N_1158,N_1075,N_1084);
or U1159 (N_1159,N_1097,N_1116);
and U1160 (N_1160,N_1115,N_1098);
nand U1161 (N_1161,N_1070,N_1109);
and U1162 (N_1162,N_1100,N_1079);
xnor U1163 (N_1163,N_1093,N_1100);
and U1164 (N_1164,N_1059,N_1106);
and U1165 (N_1165,N_1097,N_1102);
and U1166 (N_1166,N_1057,N_1080);
or U1167 (N_1167,N_1068,N_1055);
or U1168 (N_1168,N_1069,N_1099);
and U1169 (N_1169,N_1087,N_1092);
or U1170 (N_1170,N_1109,N_1103);
nor U1171 (N_1171,N_1079,N_1103);
nand U1172 (N_1172,N_1075,N_1060);
or U1173 (N_1173,N_1085,N_1086);
nor U1174 (N_1174,N_1073,N_1100);
nor U1175 (N_1175,N_1076,N_1119);
nor U1176 (N_1176,N_1114,N_1067);
and U1177 (N_1177,N_1106,N_1053);
or U1178 (N_1178,N_1080,N_1050);
and U1179 (N_1179,N_1099,N_1052);
nand U1180 (N_1180,N_1053,N_1060);
or U1181 (N_1181,N_1107,N_1093);
xnor U1182 (N_1182,N_1105,N_1113);
or U1183 (N_1183,N_1119,N_1117);
or U1184 (N_1184,N_1100,N_1068);
xnor U1185 (N_1185,N_1086,N_1118);
and U1186 (N_1186,N_1116,N_1122);
and U1187 (N_1187,N_1106,N_1065);
nand U1188 (N_1188,N_1067,N_1099);
xor U1189 (N_1189,N_1116,N_1070);
and U1190 (N_1190,N_1092,N_1108);
xor U1191 (N_1191,N_1119,N_1120);
nor U1192 (N_1192,N_1115,N_1053);
xnor U1193 (N_1193,N_1093,N_1065);
and U1194 (N_1194,N_1077,N_1104);
nand U1195 (N_1195,N_1055,N_1082);
nand U1196 (N_1196,N_1122,N_1123);
and U1197 (N_1197,N_1085,N_1050);
nand U1198 (N_1198,N_1082,N_1101);
nor U1199 (N_1199,N_1064,N_1102);
and U1200 (N_1200,N_1133,N_1147);
or U1201 (N_1201,N_1166,N_1172);
nand U1202 (N_1202,N_1155,N_1179);
nor U1203 (N_1203,N_1132,N_1195);
nor U1204 (N_1204,N_1148,N_1129);
nor U1205 (N_1205,N_1127,N_1189);
nor U1206 (N_1206,N_1178,N_1143);
nand U1207 (N_1207,N_1126,N_1131);
nand U1208 (N_1208,N_1162,N_1142);
nand U1209 (N_1209,N_1137,N_1176);
and U1210 (N_1210,N_1175,N_1146);
nand U1211 (N_1211,N_1144,N_1159);
and U1212 (N_1212,N_1185,N_1141);
or U1213 (N_1213,N_1163,N_1165);
nor U1214 (N_1214,N_1152,N_1198);
or U1215 (N_1215,N_1173,N_1177);
and U1216 (N_1216,N_1157,N_1174);
nand U1217 (N_1217,N_1151,N_1181);
xnor U1218 (N_1218,N_1130,N_1183);
and U1219 (N_1219,N_1186,N_1190);
xor U1220 (N_1220,N_1135,N_1199);
nor U1221 (N_1221,N_1187,N_1188);
or U1222 (N_1222,N_1140,N_1145);
or U1223 (N_1223,N_1158,N_1192);
nand U1224 (N_1224,N_1139,N_1182);
nor U1225 (N_1225,N_1138,N_1136);
nor U1226 (N_1226,N_1191,N_1180);
nand U1227 (N_1227,N_1134,N_1171);
nand U1228 (N_1228,N_1164,N_1194);
xor U1229 (N_1229,N_1160,N_1170);
nor U1230 (N_1230,N_1167,N_1154);
nand U1231 (N_1231,N_1128,N_1169);
nor U1232 (N_1232,N_1168,N_1196);
or U1233 (N_1233,N_1153,N_1150);
and U1234 (N_1234,N_1149,N_1156);
and U1235 (N_1235,N_1184,N_1193);
xor U1236 (N_1236,N_1161,N_1125);
nand U1237 (N_1237,N_1197,N_1173);
xnor U1238 (N_1238,N_1137,N_1181);
or U1239 (N_1239,N_1147,N_1136);
nor U1240 (N_1240,N_1157,N_1173);
nor U1241 (N_1241,N_1167,N_1178);
nor U1242 (N_1242,N_1170,N_1191);
or U1243 (N_1243,N_1197,N_1164);
nor U1244 (N_1244,N_1191,N_1184);
and U1245 (N_1245,N_1190,N_1137);
nand U1246 (N_1246,N_1149,N_1140);
xnor U1247 (N_1247,N_1154,N_1169);
and U1248 (N_1248,N_1182,N_1155);
or U1249 (N_1249,N_1128,N_1139);
nand U1250 (N_1250,N_1138,N_1145);
xnor U1251 (N_1251,N_1156,N_1170);
nand U1252 (N_1252,N_1175,N_1159);
or U1253 (N_1253,N_1193,N_1125);
nor U1254 (N_1254,N_1147,N_1194);
nor U1255 (N_1255,N_1126,N_1135);
or U1256 (N_1256,N_1179,N_1186);
or U1257 (N_1257,N_1186,N_1171);
or U1258 (N_1258,N_1152,N_1185);
nor U1259 (N_1259,N_1134,N_1159);
and U1260 (N_1260,N_1126,N_1138);
nor U1261 (N_1261,N_1131,N_1140);
and U1262 (N_1262,N_1190,N_1132);
nand U1263 (N_1263,N_1163,N_1169);
or U1264 (N_1264,N_1152,N_1169);
and U1265 (N_1265,N_1193,N_1154);
nand U1266 (N_1266,N_1127,N_1144);
nor U1267 (N_1267,N_1172,N_1146);
nand U1268 (N_1268,N_1154,N_1138);
or U1269 (N_1269,N_1173,N_1128);
and U1270 (N_1270,N_1191,N_1171);
and U1271 (N_1271,N_1128,N_1177);
nand U1272 (N_1272,N_1142,N_1165);
nand U1273 (N_1273,N_1179,N_1182);
or U1274 (N_1274,N_1170,N_1178);
or U1275 (N_1275,N_1212,N_1245);
or U1276 (N_1276,N_1253,N_1239);
and U1277 (N_1277,N_1247,N_1240);
and U1278 (N_1278,N_1214,N_1271);
nand U1279 (N_1279,N_1238,N_1224);
and U1280 (N_1280,N_1207,N_1232);
nor U1281 (N_1281,N_1203,N_1251);
xor U1282 (N_1282,N_1249,N_1263);
and U1283 (N_1283,N_1206,N_1274);
and U1284 (N_1284,N_1216,N_1223);
nor U1285 (N_1285,N_1272,N_1273);
and U1286 (N_1286,N_1246,N_1248);
nor U1287 (N_1287,N_1261,N_1234);
and U1288 (N_1288,N_1250,N_1225);
nand U1289 (N_1289,N_1220,N_1211);
xor U1290 (N_1290,N_1201,N_1242);
nand U1291 (N_1291,N_1228,N_1236);
xor U1292 (N_1292,N_1218,N_1265);
and U1293 (N_1293,N_1237,N_1267);
nand U1294 (N_1294,N_1230,N_1256);
and U1295 (N_1295,N_1227,N_1233);
nor U1296 (N_1296,N_1270,N_1217);
or U1297 (N_1297,N_1204,N_1235);
nor U1298 (N_1298,N_1226,N_1257);
and U1299 (N_1299,N_1255,N_1222);
and U1300 (N_1300,N_1252,N_1210);
nor U1301 (N_1301,N_1205,N_1258);
or U1302 (N_1302,N_1244,N_1241);
nand U1303 (N_1303,N_1254,N_1221);
xor U1304 (N_1304,N_1264,N_1266);
nor U1305 (N_1305,N_1215,N_1219);
nor U1306 (N_1306,N_1209,N_1231);
nor U1307 (N_1307,N_1202,N_1262);
or U1308 (N_1308,N_1229,N_1269);
nor U1309 (N_1309,N_1260,N_1243);
nor U1310 (N_1310,N_1200,N_1208);
or U1311 (N_1311,N_1259,N_1213);
nor U1312 (N_1312,N_1268,N_1263);
nor U1313 (N_1313,N_1210,N_1270);
nand U1314 (N_1314,N_1205,N_1252);
or U1315 (N_1315,N_1204,N_1202);
nand U1316 (N_1316,N_1237,N_1251);
nand U1317 (N_1317,N_1202,N_1225);
nand U1318 (N_1318,N_1200,N_1229);
and U1319 (N_1319,N_1204,N_1232);
nand U1320 (N_1320,N_1214,N_1251);
nand U1321 (N_1321,N_1255,N_1267);
nor U1322 (N_1322,N_1248,N_1272);
and U1323 (N_1323,N_1216,N_1254);
and U1324 (N_1324,N_1228,N_1268);
nand U1325 (N_1325,N_1260,N_1208);
and U1326 (N_1326,N_1212,N_1250);
and U1327 (N_1327,N_1249,N_1205);
and U1328 (N_1328,N_1272,N_1218);
nand U1329 (N_1329,N_1224,N_1247);
or U1330 (N_1330,N_1210,N_1232);
or U1331 (N_1331,N_1234,N_1236);
and U1332 (N_1332,N_1262,N_1235);
nor U1333 (N_1333,N_1267,N_1215);
xnor U1334 (N_1334,N_1260,N_1263);
nand U1335 (N_1335,N_1230,N_1236);
and U1336 (N_1336,N_1219,N_1203);
xor U1337 (N_1337,N_1253,N_1213);
and U1338 (N_1338,N_1209,N_1212);
xnor U1339 (N_1339,N_1257,N_1216);
and U1340 (N_1340,N_1200,N_1264);
or U1341 (N_1341,N_1201,N_1221);
or U1342 (N_1342,N_1218,N_1208);
nor U1343 (N_1343,N_1201,N_1232);
and U1344 (N_1344,N_1254,N_1237);
nand U1345 (N_1345,N_1233,N_1250);
nor U1346 (N_1346,N_1253,N_1217);
nand U1347 (N_1347,N_1264,N_1252);
or U1348 (N_1348,N_1229,N_1228);
and U1349 (N_1349,N_1273,N_1212);
and U1350 (N_1350,N_1302,N_1285);
or U1351 (N_1351,N_1309,N_1319);
nor U1352 (N_1352,N_1346,N_1329);
nor U1353 (N_1353,N_1348,N_1284);
nor U1354 (N_1354,N_1303,N_1291);
nor U1355 (N_1355,N_1308,N_1289);
or U1356 (N_1356,N_1340,N_1313);
and U1357 (N_1357,N_1321,N_1338);
nor U1358 (N_1358,N_1283,N_1298);
nand U1359 (N_1359,N_1278,N_1306);
nand U1360 (N_1360,N_1320,N_1318);
xor U1361 (N_1361,N_1330,N_1323);
xor U1362 (N_1362,N_1310,N_1326);
or U1363 (N_1363,N_1279,N_1324);
xnor U1364 (N_1364,N_1281,N_1296);
and U1365 (N_1365,N_1342,N_1295);
and U1366 (N_1366,N_1305,N_1304);
nand U1367 (N_1367,N_1336,N_1314);
nor U1368 (N_1368,N_1300,N_1275);
xnor U1369 (N_1369,N_1286,N_1335);
or U1370 (N_1370,N_1349,N_1293);
xor U1371 (N_1371,N_1277,N_1311);
nor U1372 (N_1372,N_1316,N_1307);
or U1373 (N_1373,N_1315,N_1337);
nor U1374 (N_1374,N_1344,N_1297);
nor U1375 (N_1375,N_1322,N_1339);
nand U1376 (N_1376,N_1282,N_1294);
nor U1377 (N_1377,N_1333,N_1325);
nand U1378 (N_1378,N_1312,N_1288);
nor U1379 (N_1379,N_1327,N_1287);
xnor U1380 (N_1380,N_1343,N_1332);
xnor U1381 (N_1381,N_1317,N_1299);
or U1382 (N_1382,N_1347,N_1280);
nor U1383 (N_1383,N_1331,N_1290);
nor U1384 (N_1384,N_1345,N_1301);
nand U1385 (N_1385,N_1292,N_1334);
nand U1386 (N_1386,N_1341,N_1276);
xor U1387 (N_1387,N_1328,N_1277);
xor U1388 (N_1388,N_1332,N_1338);
nor U1389 (N_1389,N_1283,N_1324);
and U1390 (N_1390,N_1296,N_1292);
nor U1391 (N_1391,N_1315,N_1333);
or U1392 (N_1392,N_1317,N_1339);
nand U1393 (N_1393,N_1323,N_1290);
nand U1394 (N_1394,N_1280,N_1325);
or U1395 (N_1395,N_1341,N_1298);
or U1396 (N_1396,N_1321,N_1332);
nand U1397 (N_1397,N_1344,N_1343);
and U1398 (N_1398,N_1288,N_1308);
or U1399 (N_1399,N_1326,N_1329);
nand U1400 (N_1400,N_1324,N_1282);
and U1401 (N_1401,N_1333,N_1327);
nor U1402 (N_1402,N_1303,N_1282);
or U1403 (N_1403,N_1309,N_1336);
xnor U1404 (N_1404,N_1332,N_1335);
and U1405 (N_1405,N_1333,N_1284);
nand U1406 (N_1406,N_1284,N_1294);
and U1407 (N_1407,N_1343,N_1308);
nor U1408 (N_1408,N_1344,N_1277);
xnor U1409 (N_1409,N_1327,N_1291);
nor U1410 (N_1410,N_1312,N_1335);
nand U1411 (N_1411,N_1322,N_1286);
or U1412 (N_1412,N_1298,N_1312);
nand U1413 (N_1413,N_1304,N_1299);
nand U1414 (N_1414,N_1306,N_1343);
or U1415 (N_1415,N_1297,N_1290);
or U1416 (N_1416,N_1311,N_1335);
nor U1417 (N_1417,N_1280,N_1295);
and U1418 (N_1418,N_1346,N_1296);
nor U1419 (N_1419,N_1321,N_1303);
and U1420 (N_1420,N_1282,N_1296);
nand U1421 (N_1421,N_1308,N_1348);
nand U1422 (N_1422,N_1279,N_1318);
nor U1423 (N_1423,N_1292,N_1304);
nor U1424 (N_1424,N_1315,N_1299);
xor U1425 (N_1425,N_1414,N_1364);
and U1426 (N_1426,N_1407,N_1411);
and U1427 (N_1427,N_1419,N_1369);
and U1428 (N_1428,N_1381,N_1368);
nand U1429 (N_1429,N_1358,N_1387);
xor U1430 (N_1430,N_1354,N_1363);
xnor U1431 (N_1431,N_1402,N_1377);
and U1432 (N_1432,N_1422,N_1362);
and U1433 (N_1433,N_1413,N_1382);
nor U1434 (N_1434,N_1374,N_1391);
nor U1435 (N_1435,N_1393,N_1361);
nor U1436 (N_1436,N_1351,N_1376);
nor U1437 (N_1437,N_1378,N_1416);
or U1438 (N_1438,N_1396,N_1365);
nand U1439 (N_1439,N_1415,N_1409);
nand U1440 (N_1440,N_1408,N_1379);
or U1441 (N_1441,N_1372,N_1367);
nand U1442 (N_1442,N_1398,N_1352);
or U1443 (N_1443,N_1406,N_1385);
nor U1444 (N_1444,N_1366,N_1386);
nand U1445 (N_1445,N_1389,N_1418);
xnor U1446 (N_1446,N_1357,N_1388);
or U1447 (N_1447,N_1380,N_1417);
and U1448 (N_1448,N_1355,N_1395);
or U1449 (N_1449,N_1400,N_1397);
nor U1450 (N_1450,N_1420,N_1371);
and U1451 (N_1451,N_1394,N_1350);
nand U1452 (N_1452,N_1423,N_1405);
xor U1453 (N_1453,N_1384,N_1403);
nor U1454 (N_1454,N_1424,N_1404);
nand U1455 (N_1455,N_1410,N_1401);
nor U1456 (N_1456,N_1390,N_1373);
and U1457 (N_1457,N_1360,N_1359);
or U1458 (N_1458,N_1370,N_1353);
nand U1459 (N_1459,N_1392,N_1421);
nand U1460 (N_1460,N_1412,N_1356);
nand U1461 (N_1461,N_1375,N_1383);
and U1462 (N_1462,N_1399,N_1405);
nand U1463 (N_1463,N_1424,N_1396);
and U1464 (N_1464,N_1377,N_1367);
and U1465 (N_1465,N_1381,N_1387);
and U1466 (N_1466,N_1351,N_1397);
xor U1467 (N_1467,N_1366,N_1421);
nand U1468 (N_1468,N_1378,N_1410);
nand U1469 (N_1469,N_1374,N_1363);
nor U1470 (N_1470,N_1397,N_1355);
xor U1471 (N_1471,N_1395,N_1372);
or U1472 (N_1472,N_1400,N_1358);
xnor U1473 (N_1473,N_1386,N_1421);
or U1474 (N_1474,N_1412,N_1384);
xor U1475 (N_1475,N_1374,N_1415);
or U1476 (N_1476,N_1422,N_1403);
nor U1477 (N_1477,N_1381,N_1397);
nand U1478 (N_1478,N_1353,N_1388);
and U1479 (N_1479,N_1387,N_1386);
nor U1480 (N_1480,N_1398,N_1358);
nand U1481 (N_1481,N_1404,N_1373);
nand U1482 (N_1482,N_1402,N_1405);
xor U1483 (N_1483,N_1397,N_1391);
or U1484 (N_1484,N_1401,N_1423);
or U1485 (N_1485,N_1382,N_1420);
or U1486 (N_1486,N_1362,N_1409);
nor U1487 (N_1487,N_1423,N_1417);
or U1488 (N_1488,N_1359,N_1412);
or U1489 (N_1489,N_1353,N_1412);
and U1490 (N_1490,N_1388,N_1350);
or U1491 (N_1491,N_1366,N_1416);
or U1492 (N_1492,N_1356,N_1369);
or U1493 (N_1493,N_1403,N_1360);
nand U1494 (N_1494,N_1395,N_1370);
or U1495 (N_1495,N_1366,N_1356);
or U1496 (N_1496,N_1362,N_1385);
or U1497 (N_1497,N_1421,N_1375);
nand U1498 (N_1498,N_1389,N_1392);
and U1499 (N_1499,N_1369,N_1359);
and U1500 (N_1500,N_1431,N_1483);
or U1501 (N_1501,N_1474,N_1471);
and U1502 (N_1502,N_1451,N_1485);
and U1503 (N_1503,N_1468,N_1477);
nor U1504 (N_1504,N_1498,N_1489);
nor U1505 (N_1505,N_1467,N_1437);
xnor U1506 (N_1506,N_1458,N_1432);
or U1507 (N_1507,N_1426,N_1425);
or U1508 (N_1508,N_1482,N_1443);
or U1509 (N_1509,N_1488,N_1453);
xnor U1510 (N_1510,N_1463,N_1454);
nor U1511 (N_1511,N_1461,N_1430);
or U1512 (N_1512,N_1492,N_1427);
nand U1513 (N_1513,N_1442,N_1473);
nor U1514 (N_1514,N_1470,N_1434);
and U1515 (N_1515,N_1444,N_1487);
nor U1516 (N_1516,N_1491,N_1490);
nand U1517 (N_1517,N_1476,N_1450);
xor U1518 (N_1518,N_1481,N_1462);
and U1519 (N_1519,N_1475,N_1441);
and U1520 (N_1520,N_1438,N_1464);
nand U1521 (N_1521,N_1447,N_1428);
and U1522 (N_1522,N_1460,N_1440);
and U1523 (N_1523,N_1469,N_1433);
nor U1524 (N_1524,N_1457,N_1499);
nor U1525 (N_1525,N_1484,N_1439);
nand U1526 (N_1526,N_1445,N_1478);
and U1527 (N_1527,N_1455,N_1449);
and U1528 (N_1528,N_1446,N_1495);
and U1529 (N_1529,N_1486,N_1435);
or U1530 (N_1530,N_1494,N_1452);
and U1531 (N_1531,N_1436,N_1479);
nand U1532 (N_1532,N_1429,N_1497);
or U1533 (N_1533,N_1480,N_1466);
and U1534 (N_1534,N_1448,N_1496);
nand U1535 (N_1535,N_1456,N_1472);
nor U1536 (N_1536,N_1459,N_1493);
or U1537 (N_1537,N_1465,N_1457);
xnor U1538 (N_1538,N_1433,N_1478);
or U1539 (N_1539,N_1475,N_1478);
and U1540 (N_1540,N_1444,N_1471);
and U1541 (N_1541,N_1496,N_1483);
xor U1542 (N_1542,N_1452,N_1429);
or U1543 (N_1543,N_1480,N_1454);
xor U1544 (N_1544,N_1449,N_1495);
or U1545 (N_1545,N_1473,N_1452);
nand U1546 (N_1546,N_1440,N_1477);
or U1547 (N_1547,N_1441,N_1436);
nand U1548 (N_1548,N_1495,N_1428);
or U1549 (N_1549,N_1481,N_1476);
and U1550 (N_1550,N_1427,N_1431);
nand U1551 (N_1551,N_1443,N_1442);
and U1552 (N_1552,N_1485,N_1466);
nor U1553 (N_1553,N_1458,N_1466);
nor U1554 (N_1554,N_1481,N_1455);
nor U1555 (N_1555,N_1459,N_1471);
nor U1556 (N_1556,N_1442,N_1446);
nor U1557 (N_1557,N_1469,N_1465);
and U1558 (N_1558,N_1426,N_1427);
and U1559 (N_1559,N_1459,N_1445);
nand U1560 (N_1560,N_1475,N_1433);
and U1561 (N_1561,N_1450,N_1456);
nor U1562 (N_1562,N_1469,N_1436);
and U1563 (N_1563,N_1481,N_1467);
nand U1564 (N_1564,N_1445,N_1484);
nand U1565 (N_1565,N_1464,N_1449);
or U1566 (N_1566,N_1439,N_1445);
nand U1567 (N_1567,N_1449,N_1448);
nor U1568 (N_1568,N_1443,N_1478);
nand U1569 (N_1569,N_1454,N_1434);
or U1570 (N_1570,N_1446,N_1444);
nand U1571 (N_1571,N_1465,N_1444);
nand U1572 (N_1572,N_1464,N_1470);
or U1573 (N_1573,N_1426,N_1467);
and U1574 (N_1574,N_1448,N_1451);
nor U1575 (N_1575,N_1553,N_1541);
xnor U1576 (N_1576,N_1542,N_1517);
nor U1577 (N_1577,N_1556,N_1568);
xnor U1578 (N_1578,N_1512,N_1539);
and U1579 (N_1579,N_1508,N_1558);
or U1580 (N_1580,N_1565,N_1552);
or U1581 (N_1581,N_1528,N_1524);
and U1582 (N_1582,N_1530,N_1500);
nand U1583 (N_1583,N_1506,N_1550);
or U1584 (N_1584,N_1544,N_1567);
nor U1585 (N_1585,N_1520,N_1569);
xnor U1586 (N_1586,N_1536,N_1564);
or U1587 (N_1587,N_1509,N_1514);
and U1588 (N_1588,N_1573,N_1572);
and U1589 (N_1589,N_1526,N_1502);
nand U1590 (N_1590,N_1563,N_1549);
nor U1591 (N_1591,N_1570,N_1515);
nand U1592 (N_1592,N_1534,N_1557);
and U1593 (N_1593,N_1503,N_1537);
and U1594 (N_1594,N_1540,N_1559);
or U1595 (N_1595,N_1571,N_1511);
nand U1596 (N_1596,N_1560,N_1538);
xnor U1597 (N_1597,N_1504,N_1543);
and U1598 (N_1598,N_1513,N_1562);
or U1599 (N_1599,N_1545,N_1554);
or U1600 (N_1600,N_1525,N_1516);
nor U1601 (N_1601,N_1518,N_1561);
nor U1602 (N_1602,N_1547,N_1523);
xor U1603 (N_1603,N_1548,N_1510);
nor U1604 (N_1604,N_1546,N_1527);
nor U1605 (N_1605,N_1521,N_1531);
nand U1606 (N_1606,N_1535,N_1501);
or U1607 (N_1607,N_1551,N_1505);
nand U1608 (N_1608,N_1533,N_1522);
nor U1609 (N_1609,N_1529,N_1532);
nand U1610 (N_1610,N_1555,N_1574);
nand U1611 (N_1611,N_1507,N_1519);
or U1612 (N_1612,N_1566,N_1557);
xnor U1613 (N_1613,N_1549,N_1532);
or U1614 (N_1614,N_1513,N_1567);
xor U1615 (N_1615,N_1573,N_1571);
xnor U1616 (N_1616,N_1510,N_1569);
nor U1617 (N_1617,N_1565,N_1562);
or U1618 (N_1618,N_1522,N_1545);
nor U1619 (N_1619,N_1530,N_1510);
nor U1620 (N_1620,N_1535,N_1524);
or U1621 (N_1621,N_1547,N_1562);
nor U1622 (N_1622,N_1558,N_1568);
nor U1623 (N_1623,N_1510,N_1517);
or U1624 (N_1624,N_1501,N_1564);
xnor U1625 (N_1625,N_1556,N_1539);
xor U1626 (N_1626,N_1528,N_1510);
and U1627 (N_1627,N_1515,N_1543);
or U1628 (N_1628,N_1547,N_1536);
nand U1629 (N_1629,N_1564,N_1574);
nand U1630 (N_1630,N_1553,N_1522);
and U1631 (N_1631,N_1546,N_1512);
nor U1632 (N_1632,N_1520,N_1512);
or U1633 (N_1633,N_1512,N_1540);
nor U1634 (N_1634,N_1544,N_1525);
and U1635 (N_1635,N_1510,N_1539);
and U1636 (N_1636,N_1515,N_1557);
xor U1637 (N_1637,N_1505,N_1502);
nor U1638 (N_1638,N_1529,N_1524);
nor U1639 (N_1639,N_1508,N_1559);
nor U1640 (N_1640,N_1502,N_1501);
or U1641 (N_1641,N_1552,N_1568);
nand U1642 (N_1642,N_1567,N_1530);
nor U1643 (N_1643,N_1501,N_1506);
nor U1644 (N_1644,N_1563,N_1524);
nor U1645 (N_1645,N_1559,N_1572);
nor U1646 (N_1646,N_1557,N_1550);
nand U1647 (N_1647,N_1564,N_1554);
xnor U1648 (N_1648,N_1506,N_1525);
and U1649 (N_1649,N_1559,N_1510);
nor U1650 (N_1650,N_1582,N_1594);
or U1651 (N_1651,N_1621,N_1641);
xnor U1652 (N_1652,N_1595,N_1610);
nand U1653 (N_1653,N_1637,N_1646);
nor U1654 (N_1654,N_1640,N_1596);
nand U1655 (N_1655,N_1630,N_1636);
or U1656 (N_1656,N_1581,N_1587);
nor U1657 (N_1657,N_1644,N_1600);
nor U1658 (N_1658,N_1626,N_1604);
and U1659 (N_1659,N_1588,N_1616);
and U1660 (N_1660,N_1584,N_1638);
xnor U1661 (N_1661,N_1649,N_1645);
nand U1662 (N_1662,N_1635,N_1602);
nand U1663 (N_1663,N_1617,N_1639);
nor U1664 (N_1664,N_1612,N_1642);
nor U1665 (N_1665,N_1627,N_1577);
nand U1666 (N_1666,N_1619,N_1608);
nor U1667 (N_1667,N_1611,N_1605);
and U1668 (N_1668,N_1580,N_1648);
nand U1669 (N_1669,N_1606,N_1632);
nor U1670 (N_1670,N_1603,N_1615);
xor U1671 (N_1671,N_1590,N_1628);
and U1672 (N_1672,N_1601,N_1633);
and U1673 (N_1673,N_1622,N_1631);
or U1674 (N_1674,N_1618,N_1576);
or U1675 (N_1675,N_1575,N_1629);
or U1676 (N_1676,N_1579,N_1586);
xnor U1677 (N_1677,N_1634,N_1591);
nor U1678 (N_1678,N_1609,N_1597);
xor U1679 (N_1679,N_1592,N_1643);
or U1680 (N_1680,N_1599,N_1614);
or U1681 (N_1681,N_1607,N_1624);
and U1682 (N_1682,N_1620,N_1647);
nor U1683 (N_1683,N_1583,N_1625);
or U1684 (N_1684,N_1585,N_1623);
nand U1685 (N_1685,N_1613,N_1593);
nand U1686 (N_1686,N_1589,N_1578);
or U1687 (N_1687,N_1598,N_1577);
nand U1688 (N_1688,N_1614,N_1582);
or U1689 (N_1689,N_1588,N_1587);
xnor U1690 (N_1690,N_1614,N_1646);
and U1691 (N_1691,N_1648,N_1635);
nand U1692 (N_1692,N_1643,N_1616);
and U1693 (N_1693,N_1598,N_1587);
nor U1694 (N_1694,N_1577,N_1634);
xnor U1695 (N_1695,N_1648,N_1610);
nor U1696 (N_1696,N_1612,N_1620);
or U1697 (N_1697,N_1636,N_1611);
and U1698 (N_1698,N_1605,N_1595);
nand U1699 (N_1699,N_1611,N_1603);
or U1700 (N_1700,N_1586,N_1625);
nor U1701 (N_1701,N_1638,N_1641);
nor U1702 (N_1702,N_1600,N_1624);
nand U1703 (N_1703,N_1587,N_1634);
or U1704 (N_1704,N_1605,N_1592);
and U1705 (N_1705,N_1611,N_1626);
nand U1706 (N_1706,N_1616,N_1587);
and U1707 (N_1707,N_1575,N_1592);
nor U1708 (N_1708,N_1582,N_1583);
nand U1709 (N_1709,N_1636,N_1643);
xor U1710 (N_1710,N_1585,N_1632);
or U1711 (N_1711,N_1589,N_1649);
nand U1712 (N_1712,N_1628,N_1599);
nor U1713 (N_1713,N_1582,N_1589);
nor U1714 (N_1714,N_1632,N_1592);
nand U1715 (N_1715,N_1597,N_1595);
nor U1716 (N_1716,N_1583,N_1643);
nand U1717 (N_1717,N_1605,N_1599);
nor U1718 (N_1718,N_1633,N_1622);
nand U1719 (N_1719,N_1628,N_1637);
or U1720 (N_1720,N_1595,N_1614);
and U1721 (N_1721,N_1580,N_1600);
and U1722 (N_1722,N_1640,N_1611);
nor U1723 (N_1723,N_1600,N_1637);
or U1724 (N_1724,N_1600,N_1585);
and U1725 (N_1725,N_1683,N_1686);
nor U1726 (N_1726,N_1650,N_1700);
or U1727 (N_1727,N_1659,N_1713);
and U1728 (N_1728,N_1680,N_1695);
or U1729 (N_1729,N_1687,N_1661);
or U1730 (N_1730,N_1692,N_1662);
and U1731 (N_1731,N_1678,N_1693);
nand U1732 (N_1732,N_1704,N_1706);
nand U1733 (N_1733,N_1685,N_1660);
and U1734 (N_1734,N_1689,N_1719);
nand U1735 (N_1735,N_1657,N_1710);
and U1736 (N_1736,N_1676,N_1653);
nand U1737 (N_1737,N_1663,N_1651);
or U1738 (N_1738,N_1664,N_1668);
nor U1739 (N_1739,N_1715,N_1709);
xnor U1740 (N_1740,N_1690,N_1711);
and U1741 (N_1741,N_1724,N_1669);
or U1742 (N_1742,N_1666,N_1712);
nor U1743 (N_1743,N_1688,N_1702);
nand U1744 (N_1744,N_1696,N_1707);
nand U1745 (N_1745,N_1698,N_1717);
nor U1746 (N_1746,N_1723,N_1652);
and U1747 (N_1747,N_1656,N_1667);
xor U1748 (N_1748,N_1677,N_1671);
nor U1749 (N_1749,N_1722,N_1718);
nand U1750 (N_1750,N_1701,N_1684);
or U1751 (N_1751,N_1714,N_1673);
and U1752 (N_1752,N_1681,N_1675);
nor U1753 (N_1753,N_1716,N_1691);
nor U1754 (N_1754,N_1679,N_1697);
and U1755 (N_1755,N_1703,N_1720);
and U1756 (N_1756,N_1670,N_1682);
nor U1757 (N_1757,N_1655,N_1699);
nor U1758 (N_1758,N_1654,N_1665);
and U1759 (N_1759,N_1705,N_1674);
nand U1760 (N_1760,N_1658,N_1672);
xor U1761 (N_1761,N_1694,N_1708);
xor U1762 (N_1762,N_1721,N_1693);
nor U1763 (N_1763,N_1685,N_1678);
and U1764 (N_1764,N_1665,N_1663);
or U1765 (N_1765,N_1708,N_1693);
xor U1766 (N_1766,N_1718,N_1707);
or U1767 (N_1767,N_1700,N_1723);
nor U1768 (N_1768,N_1664,N_1709);
and U1769 (N_1769,N_1662,N_1722);
nor U1770 (N_1770,N_1672,N_1660);
and U1771 (N_1771,N_1720,N_1719);
nor U1772 (N_1772,N_1711,N_1693);
nor U1773 (N_1773,N_1704,N_1668);
xor U1774 (N_1774,N_1723,N_1716);
nor U1775 (N_1775,N_1706,N_1660);
xnor U1776 (N_1776,N_1662,N_1665);
nor U1777 (N_1777,N_1694,N_1653);
and U1778 (N_1778,N_1696,N_1683);
and U1779 (N_1779,N_1652,N_1691);
and U1780 (N_1780,N_1708,N_1657);
nand U1781 (N_1781,N_1665,N_1702);
nor U1782 (N_1782,N_1693,N_1698);
nor U1783 (N_1783,N_1712,N_1686);
xor U1784 (N_1784,N_1713,N_1693);
nor U1785 (N_1785,N_1692,N_1707);
or U1786 (N_1786,N_1652,N_1689);
nand U1787 (N_1787,N_1692,N_1717);
nand U1788 (N_1788,N_1680,N_1720);
xnor U1789 (N_1789,N_1669,N_1715);
and U1790 (N_1790,N_1682,N_1698);
nand U1791 (N_1791,N_1658,N_1718);
or U1792 (N_1792,N_1677,N_1661);
xnor U1793 (N_1793,N_1660,N_1697);
or U1794 (N_1794,N_1702,N_1677);
or U1795 (N_1795,N_1723,N_1675);
nor U1796 (N_1796,N_1658,N_1724);
or U1797 (N_1797,N_1660,N_1662);
nand U1798 (N_1798,N_1690,N_1669);
nor U1799 (N_1799,N_1666,N_1688);
nor U1800 (N_1800,N_1740,N_1771);
nor U1801 (N_1801,N_1751,N_1732);
nor U1802 (N_1802,N_1797,N_1776);
nand U1803 (N_1803,N_1763,N_1789);
and U1804 (N_1804,N_1768,N_1777);
or U1805 (N_1805,N_1785,N_1745);
nor U1806 (N_1806,N_1727,N_1759);
or U1807 (N_1807,N_1786,N_1750);
nor U1808 (N_1808,N_1766,N_1760);
or U1809 (N_1809,N_1775,N_1791);
nor U1810 (N_1810,N_1737,N_1772);
nor U1811 (N_1811,N_1781,N_1731);
and U1812 (N_1812,N_1755,N_1741);
and U1813 (N_1813,N_1774,N_1780);
and U1814 (N_1814,N_1729,N_1738);
or U1815 (N_1815,N_1794,N_1767);
nand U1816 (N_1816,N_1733,N_1769);
nor U1817 (N_1817,N_1788,N_1725);
nor U1818 (N_1818,N_1761,N_1773);
and U1819 (N_1819,N_1757,N_1736);
and U1820 (N_1820,N_1739,N_1795);
or U1821 (N_1821,N_1730,N_1793);
nand U1822 (N_1822,N_1778,N_1783);
or U1823 (N_1823,N_1756,N_1784);
xnor U1824 (N_1824,N_1726,N_1762);
xor U1825 (N_1825,N_1796,N_1742);
xor U1826 (N_1826,N_1779,N_1747);
nor U1827 (N_1827,N_1765,N_1746);
or U1828 (N_1828,N_1728,N_1743);
and U1829 (N_1829,N_1754,N_1744);
nor U1830 (N_1830,N_1792,N_1753);
nor U1831 (N_1831,N_1790,N_1782);
and U1832 (N_1832,N_1770,N_1758);
and U1833 (N_1833,N_1735,N_1787);
and U1834 (N_1834,N_1798,N_1749);
or U1835 (N_1835,N_1764,N_1799);
nand U1836 (N_1836,N_1734,N_1748);
and U1837 (N_1837,N_1752,N_1748);
nand U1838 (N_1838,N_1783,N_1784);
nor U1839 (N_1839,N_1788,N_1762);
xnor U1840 (N_1840,N_1785,N_1799);
and U1841 (N_1841,N_1760,N_1789);
nor U1842 (N_1842,N_1789,N_1747);
or U1843 (N_1843,N_1795,N_1791);
xor U1844 (N_1844,N_1778,N_1758);
nor U1845 (N_1845,N_1790,N_1794);
or U1846 (N_1846,N_1742,N_1745);
nor U1847 (N_1847,N_1798,N_1792);
or U1848 (N_1848,N_1798,N_1750);
nand U1849 (N_1849,N_1783,N_1769);
nand U1850 (N_1850,N_1728,N_1729);
nor U1851 (N_1851,N_1732,N_1799);
or U1852 (N_1852,N_1752,N_1740);
xnor U1853 (N_1853,N_1765,N_1767);
nor U1854 (N_1854,N_1780,N_1775);
and U1855 (N_1855,N_1792,N_1740);
and U1856 (N_1856,N_1770,N_1738);
and U1857 (N_1857,N_1746,N_1733);
nand U1858 (N_1858,N_1733,N_1764);
and U1859 (N_1859,N_1754,N_1725);
nand U1860 (N_1860,N_1733,N_1761);
and U1861 (N_1861,N_1727,N_1798);
nor U1862 (N_1862,N_1793,N_1791);
or U1863 (N_1863,N_1791,N_1740);
nand U1864 (N_1864,N_1728,N_1790);
xnor U1865 (N_1865,N_1766,N_1777);
nor U1866 (N_1866,N_1742,N_1792);
nand U1867 (N_1867,N_1787,N_1799);
nor U1868 (N_1868,N_1757,N_1739);
and U1869 (N_1869,N_1750,N_1784);
xnor U1870 (N_1870,N_1752,N_1759);
xnor U1871 (N_1871,N_1727,N_1771);
or U1872 (N_1872,N_1778,N_1756);
nand U1873 (N_1873,N_1742,N_1751);
nand U1874 (N_1874,N_1726,N_1774);
xor U1875 (N_1875,N_1860,N_1826);
nand U1876 (N_1876,N_1817,N_1835);
or U1877 (N_1877,N_1842,N_1832);
nand U1878 (N_1878,N_1849,N_1818);
and U1879 (N_1879,N_1831,N_1851);
nor U1880 (N_1880,N_1830,N_1837);
xor U1881 (N_1881,N_1862,N_1812);
nor U1882 (N_1882,N_1845,N_1873);
or U1883 (N_1883,N_1840,N_1811);
or U1884 (N_1884,N_1859,N_1819);
and U1885 (N_1885,N_1872,N_1854);
and U1886 (N_1886,N_1871,N_1814);
nor U1887 (N_1887,N_1857,N_1825);
xor U1888 (N_1888,N_1852,N_1844);
nand U1889 (N_1889,N_1810,N_1846);
and U1890 (N_1890,N_1815,N_1801);
and U1891 (N_1891,N_1848,N_1804);
xor U1892 (N_1892,N_1805,N_1858);
and U1893 (N_1893,N_1866,N_1853);
nor U1894 (N_1894,N_1800,N_1841);
nor U1895 (N_1895,N_1809,N_1864);
or U1896 (N_1896,N_1855,N_1823);
nor U1897 (N_1897,N_1870,N_1867);
or U1898 (N_1898,N_1874,N_1827);
nor U1899 (N_1899,N_1803,N_1863);
and U1900 (N_1900,N_1816,N_1808);
or U1901 (N_1901,N_1828,N_1839);
and U1902 (N_1902,N_1807,N_1856);
or U1903 (N_1903,N_1820,N_1821);
or U1904 (N_1904,N_1834,N_1802);
nor U1905 (N_1905,N_1813,N_1850);
or U1906 (N_1906,N_1824,N_1833);
and U1907 (N_1907,N_1869,N_1829);
and U1908 (N_1908,N_1865,N_1806);
nand U1909 (N_1909,N_1836,N_1847);
nand U1910 (N_1910,N_1838,N_1861);
nand U1911 (N_1911,N_1822,N_1868);
nor U1912 (N_1912,N_1843,N_1804);
xnor U1913 (N_1913,N_1804,N_1862);
and U1914 (N_1914,N_1850,N_1804);
or U1915 (N_1915,N_1874,N_1848);
nand U1916 (N_1916,N_1816,N_1828);
or U1917 (N_1917,N_1824,N_1838);
nor U1918 (N_1918,N_1806,N_1807);
nor U1919 (N_1919,N_1803,N_1858);
or U1920 (N_1920,N_1871,N_1845);
or U1921 (N_1921,N_1814,N_1825);
xor U1922 (N_1922,N_1863,N_1834);
or U1923 (N_1923,N_1804,N_1830);
xor U1924 (N_1924,N_1863,N_1854);
nand U1925 (N_1925,N_1807,N_1839);
nand U1926 (N_1926,N_1820,N_1806);
or U1927 (N_1927,N_1809,N_1820);
or U1928 (N_1928,N_1812,N_1822);
nand U1929 (N_1929,N_1804,N_1855);
nor U1930 (N_1930,N_1810,N_1818);
or U1931 (N_1931,N_1808,N_1827);
and U1932 (N_1932,N_1864,N_1846);
nand U1933 (N_1933,N_1870,N_1849);
nor U1934 (N_1934,N_1839,N_1871);
nand U1935 (N_1935,N_1808,N_1823);
nor U1936 (N_1936,N_1863,N_1827);
nand U1937 (N_1937,N_1866,N_1822);
or U1938 (N_1938,N_1862,N_1849);
nand U1939 (N_1939,N_1821,N_1805);
or U1940 (N_1940,N_1866,N_1865);
nand U1941 (N_1941,N_1863,N_1835);
or U1942 (N_1942,N_1837,N_1841);
and U1943 (N_1943,N_1801,N_1804);
nor U1944 (N_1944,N_1866,N_1821);
nand U1945 (N_1945,N_1813,N_1826);
and U1946 (N_1946,N_1800,N_1823);
nor U1947 (N_1947,N_1871,N_1865);
nand U1948 (N_1948,N_1860,N_1813);
and U1949 (N_1949,N_1803,N_1825);
nand U1950 (N_1950,N_1913,N_1883);
and U1951 (N_1951,N_1942,N_1893);
or U1952 (N_1952,N_1925,N_1929);
and U1953 (N_1953,N_1909,N_1943);
and U1954 (N_1954,N_1896,N_1918);
or U1955 (N_1955,N_1931,N_1911);
or U1956 (N_1956,N_1927,N_1928);
nor U1957 (N_1957,N_1920,N_1908);
and U1958 (N_1958,N_1887,N_1924);
nor U1959 (N_1959,N_1895,N_1898);
and U1960 (N_1960,N_1948,N_1939);
nor U1961 (N_1961,N_1905,N_1876);
nor U1962 (N_1962,N_1888,N_1914);
and U1963 (N_1963,N_1936,N_1880);
and U1964 (N_1964,N_1949,N_1889);
and U1965 (N_1965,N_1884,N_1917);
and U1966 (N_1966,N_1932,N_1879);
or U1967 (N_1967,N_1894,N_1897);
and U1968 (N_1968,N_1875,N_1912);
nand U1969 (N_1969,N_1900,N_1892);
xnor U1970 (N_1970,N_1899,N_1919);
nand U1971 (N_1971,N_1926,N_1885);
nand U1972 (N_1972,N_1933,N_1891);
xnor U1973 (N_1973,N_1930,N_1940);
nor U1974 (N_1974,N_1916,N_1901);
and U1975 (N_1975,N_1882,N_1922);
nor U1976 (N_1976,N_1878,N_1945);
nor U1977 (N_1977,N_1923,N_1946);
nand U1978 (N_1978,N_1881,N_1941);
nor U1979 (N_1979,N_1937,N_1915);
and U1980 (N_1980,N_1935,N_1890);
nand U1981 (N_1981,N_1906,N_1910);
nand U1982 (N_1982,N_1904,N_1877);
nor U1983 (N_1983,N_1907,N_1886);
nor U1984 (N_1984,N_1902,N_1947);
nand U1985 (N_1985,N_1903,N_1944);
and U1986 (N_1986,N_1921,N_1934);
xnor U1987 (N_1987,N_1938,N_1935);
nand U1988 (N_1988,N_1905,N_1903);
xor U1989 (N_1989,N_1877,N_1918);
nand U1990 (N_1990,N_1907,N_1944);
nand U1991 (N_1991,N_1932,N_1905);
and U1992 (N_1992,N_1908,N_1902);
nand U1993 (N_1993,N_1893,N_1918);
nor U1994 (N_1994,N_1939,N_1923);
nand U1995 (N_1995,N_1907,N_1936);
and U1996 (N_1996,N_1924,N_1948);
and U1997 (N_1997,N_1901,N_1946);
nand U1998 (N_1998,N_1877,N_1905);
and U1999 (N_1999,N_1934,N_1920);
nor U2000 (N_2000,N_1910,N_1937);
xor U2001 (N_2001,N_1917,N_1905);
and U2002 (N_2002,N_1893,N_1940);
or U2003 (N_2003,N_1936,N_1886);
nand U2004 (N_2004,N_1949,N_1929);
nand U2005 (N_2005,N_1918,N_1886);
or U2006 (N_2006,N_1880,N_1927);
xor U2007 (N_2007,N_1933,N_1923);
nor U2008 (N_2008,N_1911,N_1923);
and U2009 (N_2009,N_1921,N_1925);
or U2010 (N_2010,N_1876,N_1881);
or U2011 (N_2011,N_1917,N_1939);
or U2012 (N_2012,N_1937,N_1878);
xnor U2013 (N_2013,N_1894,N_1888);
nor U2014 (N_2014,N_1899,N_1892);
nor U2015 (N_2015,N_1921,N_1909);
nor U2016 (N_2016,N_1895,N_1902);
and U2017 (N_2017,N_1894,N_1948);
nor U2018 (N_2018,N_1896,N_1913);
and U2019 (N_2019,N_1943,N_1947);
nand U2020 (N_2020,N_1925,N_1884);
nor U2021 (N_2021,N_1922,N_1938);
or U2022 (N_2022,N_1922,N_1928);
xor U2023 (N_2023,N_1930,N_1944);
and U2024 (N_2024,N_1919,N_1934);
nand U2025 (N_2025,N_1970,N_2014);
or U2026 (N_2026,N_1994,N_2022);
and U2027 (N_2027,N_1960,N_1978);
nor U2028 (N_2028,N_2021,N_1972);
xor U2029 (N_2029,N_1963,N_2016);
nand U2030 (N_2030,N_1977,N_1951);
nand U2031 (N_2031,N_2012,N_2023);
or U2032 (N_2032,N_2020,N_1993);
xnor U2033 (N_2033,N_1991,N_1967);
nor U2034 (N_2034,N_1987,N_1974);
nand U2035 (N_2035,N_1953,N_1965);
nor U2036 (N_2036,N_2004,N_1990);
xnor U2037 (N_2037,N_1961,N_1962);
and U2038 (N_2038,N_1959,N_1996);
or U2039 (N_2039,N_1957,N_1971);
or U2040 (N_2040,N_1968,N_2013);
nor U2041 (N_2041,N_2017,N_2002);
or U2042 (N_2042,N_1985,N_2005);
or U2043 (N_2043,N_1988,N_2006);
nand U2044 (N_2044,N_2015,N_1979);
or U2045 (N_2045,N_1950,N_1969);
and U2046 (N_2046,N_2010,N_1966);
nor U2047 (N_2047,N_1954,N_1984);
nor U2048 (N_2048,N_1995,N_1992);
or U2049 (N_2049,N_2008,N_1952);
xor U2050 (N_2050,N_1976,N_1981);
and U2051 (N_2051,N_1956,N_1997);
nor U2052 (N_2052,N_1980,N_2003);
and U2053 (N_2053,N_1989,N_1982);
nor U2054 (N_2054,N_2007,N_1975);
and U2055 (N_2055,N_2018,N_1983);
nor U2056 (N_2056,N_2019,N_2001);
xor U2057 (N_2057,N_2009,N_2024);
nor U2058 (N_2058,N_1958,N_1964);
or U2059 (N_2059,N_1998,N_1955);
nand U2060 (N_2060,N_1986,N_2011);
xnor U2061 (N_2061,N_1999,N_2000);
or U2062 (N_2062,N_1973,N_2020);
nor U2063 (N_2063,N_2013,N_1960);
or U2064 (N_2064,N_1996,N_1966);
nand U2065 (N_2065,N_1957,N_1972);
nor U2066 (N_2066,N_1957,N_2024);
nand U2067 (N_2067,N_2020,N_2007);
xor U2068 (N_2068,N_1987,N_1991);
nor U2069 (N_2069,N_1971,N_1950);
or U2070 (N_2070,N_1957,N_2015);
and U2071 (N_2071,N_2004,N_1977);
nor U2072 (N_2072,N_1999,N_2017);
or U2073 (N_2073,N_1966,N_1979);
nand U2074 (N_2074,N_1974,N_2017);
and U2075 (N_2075,N_2024,N_1969);
nand U2076 (N_2076,N_1993,N_1956);
xor U2077 (N_2077,N_1954,N_1994);
nand U2078 (N_2078,N_1981,N_1993);
and U2079 (N_2079,N_1981,N_1977);
and U2080 (N_2080,N_2014,N_1958);
nor U2081 (N_2081,N_2007,N_1999);
nand U2082 (N_2082,N_1970,N_1960);
and U2083 (N_2083,N_2022,N_1996);
nor U2084 (N_2084,N_1992,N_1984);
nand U2085 (N_2085,N_1999,N_2021);
nor U2086 (N_2086,N_2009,N_2023);
nand U2087 (N_2087,N_1976,N_2006);
nand U2088 (N_2088,N_1995,N_1982);
or U2089 (N_2089,N_1961,N_1964);
nand U2090 (N_2090,N_2011,N_1955);
or U2091 (N_2091,N_1979,N_2007);
xor U2092 (N_2092,N_1966,N_1964);
and U2093 (N_2093,N_1991,N_1986);
nand U2094 (N_2094,N_2007,N_1950);
nor U2095 (N_2095,N_1975,N_2024);
and U2096 (N_2096,N_1950,N_1951);
and U2097 (N_2097,N_1962,N_1992);
nand U2098 (N_2098,N_1989,N_1977);
or U2099 (N_2099,N_1978,N_1973);
nor U2100 (N_2100,N_2043,N_2026);
or U2101 (N_2101,N_2057,N_2046);
or U2102 (N_2102,N_2098,N_2066);
nor U2103 (N_2103,N_2028,N_2070);
nand U2104 (N_2104,N_2088,N_2081);
nand U2105 (N_2105,N_2051,N_2037);
nand U2106 (N_2106,N_2069,N_2062);
nor U2107 (N_2107,N_2080,N_2092);
xnor U2108 (N_2108,N_2054,N_2064);
nand U2109 (N_2109,N_2091,N_2084);
nand U2110 (N_2110,N_2065,N_2052);
and U2111 (N_2111,N_2039,N_2053);
nand U2112 (N_2112,N_2089,N_2056);
or U2113 (N_2113,N_2082,N_2068);
or U2114 (N_2114,N_2076,N_2058);
nor U2115 (N_2115,N_2049,N_2048);
and U2116 (N_2116,N_2095,N_2079);
nand U2117 (N_2117,N_2072,N_2031);
nand U2118 (N_2118,N_2038,N_2078);
nand U2119 (N_2119,N_2044,N_2029);
and U2120 (N_2120,N_2075,N_2093);
or U2121 (N_2121,N_2097,N_2060);
nor U2122 (N_2122,N_2045,N_2030);
or U2123 (N_2123,N_2042,N_2055);
nand U2124 (N_2124,N_2059,N_2036);
and U2125 (N_2125,N_2086,N_2067);
or U2126 (N_2126,N_2099,N_2047);
nor U2127 (N_2127,N_2035,N_2077);
and U2128 (N_2128,N_2096,N_2041);
and U2129 (N_2129,N_2087,N_2027);
or U2130 (N_2130,N_2090,N_2073);
nand U2131 (N_2131,N_2063,N_2033);
nand U2132 (N_2132,N_2040,N_2083);
nand U2133 (N_2133,N_2025,N_2085);
xnor U2134 (N_2134,N_2071,N_2050);
nor U2135 (N_2135,N_2094,N_2034);
or U2136 (N_2136,N_2032,N_2074);
and U2137 (N_2137,N_2061,N_2096);
nor U2138 (N_2138,N_2042,N_2080);
nand U2139 (N_2139,N_2098,N_2034);
and U2140 (N_2140,N_2098,N_2064);
or U2141 (N_2141,N_2040,N_2035);
nand U2142 (N_2142,N_2092,N_2040);
nor U2143 (N_2143,N_2076,N_2073);
and U2144 (N_2144,N_2046,N_2040);
nor U2145 (N_2145,N_2057,N_2060);
and U2146 (N_2146,N_2077,N_2080);
nand U2147 (N_2147,N_2090,N_2036);
or U2148 (N_2148,N_2064,N_2074);
or U2149 (N_2149,N_2061,N_2042);
or U2150 (N_2150,N_2040,N_2057);
nand U2151 (N_2151,N_2080,N_2026);
and U2152 (N_2152,N_2048,N_2040);
nand U2153 (N_2153,N_2095,N_2061);
nor U2154 (N_2154,N_2079,N_2069);
and U2155 (N_2155,N_2027,N_2081);
xnor U2156 (N_2156,N_2045,N_2084);
nand U2157 (N_2157,N_2097,N_2077);
or U2158 (N_2158,N_2082,N_2034);
or U2159 (N_2159,N_2070,N_2092);
and U2160 (N_2160,N_2095,N_2088);
and U2161 (N_2161,N_2092,N_2025);
nand U2162 (N_2162,N_2054,N_2061);
nor U2163 (N_2163,N_2056,N_2031);
and U2164 (N_2164,N_2032,N_2030);
or U2165 (N_2165,N_2052,N_2054);
or U2166 (N_2166,N_2052,N_2086);
nor U2167 (N_2167,N_2025,N_2094);
or U2168 (N_2168,N_2036,N_2061);
and U2169 (N_2169,N_2052,N_2033);
and U2170 (N_2170,N_2091,N_2070);
nand U2171 (N_2171,N_2051,N_2042);
nand U2172 (N_2172,N_2092,N_2089);
nor U2173 (N_2173,N_2099,N_2083);
xor U2174 (N_2174,N_2062,N_2093);
or U2175 (N_2175,N_2173,N_2142);
or U2176 (N_2176,N_2119,N_2100);
xor U2177 (N_2177,N_2105,N_2170);
nand U2178 (N_2178,N_2148,N_2145);
nand U2179 (N_2179,N_2159,N_2103);
nand U2180 (N_2180,N_2132,N_2127);
or U2181 (N_2181,N_2124,N_2165);
or U2182 (N_2182,N_2123,N_2140);
or U2183 (N_2183,N_2109,N_2115);
nand U2184 (N_2184,N_2152,N_2144);
nor U2185 (N_2185,N_2106,N_2111);
xor U2186 (N_2186,N_2160,N_2156);
or U2187 (N_2187,N_2174,N_2134);
nor U2188 (N_2188,N_2133,N_2162);
or U2189 (N_2189,N_2157,N_2147);
xnor U2190 (N_2190,N_2135,N_2141);
nor U2191 (N_2191,N_2120,N_2117);
xnor U2192 (N_2192,N_2166,N_2139);
nand U2193 (N_2193,N_2129,N_2108);
or U2194 (N_2194,N_2155,N_2154);
nand U2195 (N_2195,N_2168,N_2110);
nor U2196 (N_2196,N_2169,N_2136);
nand U2197 (N_2197,N_2102,N_2172);
nor U2198 (N_2198,N_2153,N_2150);
nand U2199 (N_2199,N_2146,N_2116);
and U2200 (N_2200,N_2161,N_2167);
or U2201 (N_2201,N_2130,N_2113);
and U2202 (N_2202,N_2151,N_2121);
nand U2203 (N_2203,N_2101,N_2137);
or U2204 (N_2204,N_2107,N_2114);
and U2205 (N_2205,N_2104,N_2118);
nand U2206 (N_2206,N_2126,N_2149);
or U2207 (N_2207,N_2128,N_2171);
and U2208 (N_2208,N_2112,N_2164);
or U2209 (N_2209,N_2138,N_2143);
nor U2210 (N_2210,N_2163,N_2131);
or U2211 (N_2211,N_2158,N_2122);
xnor U2212 (N_2212,N_2125,N_2140);
nor U2213 (N_2213,N_2146,N_2162);
and U2214 (N_2214,N_2121,N_2104);
nor U2215 (N_2215,N_2125,N_2122);
nor U2216 (N_2216,N_2127,N_2116);
nor U2217 (N_2217,N_2135,N_2111);
xnor U2218 (N_2218,N_2167,N_2169);
nand U2219 (N_2219,N_2157,N_2159);
nand U2220 (N_2220,N_2168,N_2113);
and U2221 (N_2221,N_2156,N_2105);
xor U2222 (N_2222,N_2140,N_2114);
xor U2223 (N_2223,N_2169,N_2124);
nor U2224 (N_2224,N_2157,N_2151);
xor U2225 (N_2225,N_2131,N_2149);
and U2226 (N_2226,N_2120,N_2108);
and U2227 (N_2227,N_2170,N_2109);
or U2228 (N_2228,N_2128,N_2110);
nor U2229 (N_2229,N_2123,N_2142);
nor U2230 (N_2230,N_2138,N_2121);
xnor U2231 (N_2231,N_2102,N_2152);
nor U2232 (N_2232,N_2172,N_2133);
nor U2233 (N_2233,N_2110,N_2123);
or U2234 (N_2234,N_2162,N_2139);
and U2235 (N_2235,N_2124,N_2101);
and U2236 (N_2236,N_2121,N_2160);
or U2237 (N_2237,N_2122,N_2166);
nor U2238 (N_2238,N_2140,N_2134);
nor U2239 (N_2239,N_2140,N_2115);
xnor U2240 (N_2240,N_2155,N_2147);
xor U2241 (N_2241,N_2152,N_2172);
and U2242 (N_2242,N_2151,N_2101);
nand U2243 (N_2243,N_2133,N_2110);
nand U2244 (N_2244,N_2130,N_2132);
nor U2245 (N_2245,N_2129,N_2163);
and U2246 (N_2246,N_2154,N_2131);
nor U2247 (N_2247,N_2103,N_2115);
and U2248 (N_2248,N_2132,N_2171);
nor U2249 (N_2249,N_2135,N_2160);
nand U2250 (N_2250,N_2215,N_2189);
nor U2251 (N_2251,N_2178,N_2230);
nand U2252 (N_2252,N_2193,N_2222);
or U2253 (N_2253,N_2236,N_2223);
and U2254 (N_2254,N_2188,N_2217);
and U2255 (N_2255,N_2225,N_2247);
nor U2256 (N_2256,N_2210,N_2243);
nand U2257 (N_2257,N_2177,N_2195);
or U2258 (N_2258,N_2226,N_2228);
xnor U2259 (N_2259,N_2199,N_2197);
or U2260 (N_2260,N_2204,N_2227);
xnor U2261 (N_2261,N_2184,N_2182);
nand U2262 (N_2262,N_2190,N_2218);
and U2263 (N_2263,N_2235,N_2185);
nor U2264 (N_2264,N_2209,N_2181);
nand U2265 (N_2265,N_2196,N_2179);
nor U2266 (N_2266,N_2237,N_2187);
and U2267 (N_2267,N_2207,N_2180);
xor U2268 (N_2268,N_2198,N_2221);
nor U2269 (N_2269,N_2213,N_2234);
xnor U2270 (N_2270,N_2231,N_2192);
and U2271 (N_2271,N_2194,N_2244);
nor U2272 (N_2272,N_2245,N_2239);
nor U2273 (N_2273,N_2241,N_2212);
nor U2274 (N_2274,N_2246,N_2175);
nor U2275 (N_2275,N_2248,N_2206);
nand U2276 (N_2276,N_2208,N_2232);
nor U2277 (N_2277,N_2211,N_2202);
and U2278 (N_2278,N_2238,N_2186);
and U2279 (N_2279,N_2242,N_2220);
nand U2280 (N_2280,N_2201,N_2224);
or U2281 (N_2281,N_2240,N_2205);
nand U2282 (N_2282,N_2249,N_2216);
xor U2283 (N_2283,N_2229,N_2191);
nor U2284 (N_2284,N_2219,N_2200);
nor U2285 (N_2285,N_2233,N_2203);
nand U2286 (N_2286,N_2214,N_2183);
nor U2287 (N_2287,N_2176,N_2183);
or U2288 (N_2288,N_2177,N_2230);
and U2289 (N_2289,N_2211,N_2184);
or U2290 (N_2290,N_2226,N_2205);
and U2291 (N_2291,N_2238,N_2216);
xnor U2292 (N_2292,N_2230,N_2219);
or U2293 (N_2293,N_2197,N_2222);
nand U2294 (N_2294,N_2187,N_2197);
and U2295 (N_2295,N_2233,N_2194);
nand U2296 (N_2296,N_2199,N_2185);
nand U2297 (N_2297,N_2203,N_2232);
or U2298 (N_2298,N_2213,N_2200);
or U2299 (N_2299,N_2236,N_2224);
and U2300 (N_2300,N_2200,N_2177);
nor U2301 (N_2301,N_2185,N_2203);
nand U2302 (N_2302,N_2212,N_2192);
nor U2303 (N_2303,N_2225,N_2219);
and U2304 (N_2304,N_2212,N_2188);
xor U2305 (N_2305,N_2232,N_2191);
or U2306 (N_2306,N_2191,N_2222);
nor U2307 (N_2307,N_2229,N_2217);
nor U2308 (N_2308,N_2198,N_2194);
nor U2309 (N_2309,N_2221,N_2188);
or U2310 (N_2310,N_2242,N_2230);
nor U2311 (N_2311,N_2236,N_2191);
nor U2312 (N_2312,N_2189,N_2187);
nor U2313 (N_2313,N_2180,N_2212);
nand U2314 (N_2314,N_2232,N_2231);
nor U2315 (N_2315,N_2190,N_2207);
and U2316 (N_2316,N_2190,N_2247);
nor U2317 (N_2317,N_2226,N_2210);
or U2318 (N_2318,N_2249,N_2226);
nor U2319 (N_2319,N_2230,N_2194);
xor U2320 (N_2320,N_2227,N_2200);
nor U2321 (N_2321,N_2205,N_2200);
nand U2322 (N_2322,N_2239,N_2246);
and U2323 (N_2323,N_2202,N_2219);
xor U2324 (N_2324,N_2176,N_2181);
nand U2325 (N_2325,N_2266,N_2290);
nor U2326 (N_2326,N_2312,N_2308);
xnor U2327 (N_2327,N_2264,N_2269);
and U2328 (N_2328,N_2297,N_2298);
nand U2329 (N_2329,N_2296,N_2280);
or U2330 (N_2330,N_2294,N_2281);
xnor U2331 (N_2331,N_2284,N_2309);
and U2332 (N_2332,N_2282,N_2291);
nand U2333 (N_2333,N_2307,N_2287);
or U2334 (N_2334,N_2299,N_2311);
nand U2335 (N_2335,N_2262,N_2259);
or U2336 (N_2336,N_2320,N_2256);
xnor U2337 (N_2337,N_2319,N_2283);
and U2338 (N_2338,N_2306,N_2302);
or U2339 (N_2339,N_2301,N_2272);
xnor U2340 (N_2340,N_2268,N_2260);
and U2341 (N_2341,N_2321,N_2279);
xor U2342 (N_2342,N_2257,N_2323);
nor U2343 (N_2343,N_2254,N_2276);
or U2344 (N_2344,N_2261,N_2278);
nand U2345 (N_2345,N_2315,N_2316);
nand U2346 (N_2346,N_2253,N_2292);
and U2347 (N_2347,N_2250,N_2317);
or U2348 (N_2348,N_2251,N_2252);
nor U2349 (N_2349,N_2285,N_2313);
nor U2350 (N_2350,N_2324,N_2255);
nand U2351 (N_2351,N_2295,N_2258);
or U2352 (N_2352,N_2286,N_2318);
nand U2353 (N_2353,N_2265,N_2274);
nand U2354 (N_2354,N_2273,N_2303);
nor U2355 (N_2355,N_2322,N_2275);
and U2356 (N_2356,N_2270,N_2304);
or U2357 (N_2357,N_2288,N_2289);
nor U2358 (N_2358,N_2300,N_2293);
nor U2359 (N_2359,N_2271,N_2263);
nand U2360 (N_2360,N_2310,N_2305);
or U2361 (N_2361,N_2277,N_2314);
nand U2362 (N_2362,N_2267,N_2296);
or U2363 (N_2363,N_2277,N_2297);
nor U2364 (N_2364,N_2270,N_2277);
and U2365 (N_2365,N_2264,N_2309);
and U2366 (N_2366,N_2256,N_2304);
nor U2367 (N_2367,N_2316,N_2321);
nand U2368 (N_2368,N_2318,N_2313);
and U2369 (N_2369,N_2262,N_2254);
nor U2370 (N_2370,N_2324,N_2278);
nand U2371 (N_2371,N_2289,N_2307);
nand U2372 (N_2372,N_2273,N_2306);
and U2373 (N_2373,N_2281,N_2251);
nor U2374 (N_2374,N_2254,N_2300);
and U2375 (N_2375,N_2265,N_2318);
nand U2376 (N_2376,N_2288,N_2270);
or U2377 (N_2377,N_2266,N_2265);
or U2378 (N_2378,N_2315,N_2252);
nor U2379 (N_2379,N_2263,N_2269);
and U2380 (N_2380,N_2310,N_2318);
or U2381 (N_2381,N_2316,N_2294);
nor U2382 (N_2382,N_2295,N_2309);
nand U2383 (N_2383,N_2303,N_2296);
xor U2384 (N_2384,N_2313,N_2273);
and U2385 (N_2385,N_2266,N_2287);
nand U2386 (N_2386,N_2286,N_2279);
and U2387 (N_2387,N_2304,N_2267);
nor U2388 (N_2388,N_2285,N_2278);
and U2389 (N_2389,N_2303,N_2265);
xnor U2390 (N_2390,N_2312,N_2262);
and U2391 (N_2391,N_2276,N_2287);
xnor U2392 (N_2392,N_2253,N_2294);
or U2393 (N_2393,N_2268,N_2254);
nand U2394 (N_2394,N_2292,N_2306);
and U2395 (N_2395,N_2265,N_2275);
or U2396 (N_2396,N_2311,N_2258);
or U2397 (N_2397,N_2308,N_2276);
nor U2398 (N_2398,N_2301,N_2255);
xor U2399 (N_2399,N_2278,N_2321);
xor U2400 (N_2400,N_2332,N_2388);
and U2401 (N_2401,N_2345,N_2346);
or U2402 (N_2402,N_2348,N_2357);
or U2403 (N_2403,N_2329,N_2371);
nor U2404 (N_2404,N_2365,N_2368);
and U2405 (N_2405,N_2376,N_2356);
and U2406 (N_2406,N_2331,N_2354);
nor U2407 (N_2407,N_2359,N_2361);
nor U2408 (N_2408,N_2336,N_2363);
nand U2409 (N_2409,N_2369,N_2343);
nor U2410 (N_2410,N_2344,N_2374);
and U2411 (N_2411,N_2338,N_2373);
xnor U2412 (N_2412,N_2347,N_2379);
nand U2413 (N_2413,N_2386,N_2358);
or U2414 (N_2414,N_2362,N_2383);
and U2415 (N_2415,N_2399,N_2335);
and U2416 (N_2416,N_2325,N_2392);
and U2417 (N_2417,N_2398,N_2337);
nand U2418 (N_2418,N_2377,N_2384);
and U2419 (N_2419,N_2326,N_2366);
or U2420 (N_2420,N_2367,N_2393);
nand U2421 (N_2421,N_2378,N_2370);
nor U2422 (N_2422,N_2372,N_2364);
or U2423 (N_2423,N_2328,N_2390);
nor U2424 (N_2424,N_2334,N_2385);
nor U2425 (N_2425,N_2350,N_2341);
nand U2426 (N_2426,N_2382,N_2395);
or U2427 (N_2427,N_2387,N_2360);
nand U2428 (N_2428,N_2380,N_2396);
and U2429 (N_2429,N_2330,N_2340);
nand U2430 (N_2430,N_2349,N_2355);
xnor U2431 (N_2431,N_2352,N_2397);
xnor U2432 (N_2432,N_2327,N_2333);
xnor U2433 (N_2433,N_2342,N_2394);
nor U2434 (N_2434,N_2375,N_2353);
and U2435 (N_2435,N_2351,N_2389);
nand U2436 (N_2436,N_2391,N_2381);
nand U2437 (N_2437,N_2339,N_2334);
nand U2438 (N_2438,N_2364,N_2352);
or U2439 (N_2439,N_2338,N_2374);
nor U2440 (N_2440,N_2381,N_2383);
nand U2441 (N_2441,N_2367,N_2361);
or U2442 (N_2442,N_2334,N_2387);
nor U2443 (N_2443,N_2366,N_2327);
or U2444 (N_2444,N_2336,N_2373);
nand U2445 (N_2445,N_2327,N_2386);
nor U2446 (N_2446,N_2386,N_2339);
and U2447 (N_2447,N_2383,N_2358);
nor U2448 (N_2448,N_2353,N_2342);
nor U2449 (N_2449,N_2335,N_2370);
nand U2450 (N_2450,N_2384,N_2362);
nand U2451 (N_2451,N_2329,N_2388);
nand U2452 (N_2452,N_2330,N_2377);
and U2453 (N_2453,N_2349,N_2325);
nor U2454 (N_2454,N_2337,N_2331);
or U2455 (N_2455,N_2368,N_2388);
nor U2456 (N_2456,N_2387,N_2362);
and U2457 (N_2457,N_2353,N_2349);
nor U2458 (N_2458,N_2369,N_2363);
nor U2459 (N_2459,N_2349,N_2375);
or U2460 (N_2460,N_2365,N_2355);
nand U2461 (N_2461,N_2332,N_2339);
or U2462 (N_2462,N_2380,N_2325);
nor U2463 (N_2463,N_2342,N_2387);
and U2464 (N_2464,N_2372,N_2345);
nor U2465 (N_2465,N_2388,N_2369);
nand U2466 (N_2466,N_2360,N_2376);
nor U2467 (N_2467,N_2358,N_2347);
nand U2468 (N_2468,N_2372,N_2362);
and U2469 (N_2469,N_2393,N_2372);
nand U2470 (N_2470,N_2382,N_2372);
or U2471 (N_2471,N_2341,N_2393);
nor U2472 (N_2472,N_2369,N_2348);
and U2473 (N_2473,N_2329,N_2373);
nand U2474 (N_2474,N_2372,N_2380);
nor U2475 (N_2475,N_2412,N_2466);
nand U2476 (N_2476,N_2401,N_2421);
nand U2477 (N_2477,N_2471,N_2433);
nor U2478 (N_2478,N_2434,N_2430);
xnor U2479 (N_2479,N_2468,N_2442);
nor U2480 (N_2480,N_2447,N_2432);
nand U2481 (N_2481,N_2400,N_2414);
nand U2482 (N_2482,N_2470,N_2436);
nand U2483 (N_2483,N_2406,N_2423);
or U2484 (N_2484,N_2419,N_2457);
nor U2485 (N_2485,N_2458,N_2426);
nand U2486 (N_2486,N_2451,N_2461);
and U2487 (N_2487,N_2445,N_2444);
or U2488 (N_2488,N_2452,N_2415);
nand U2489 (N_2489,N_2463,N_2437);
or U2490 (N_2490,N_2402,N_2455);
nand U2491 (N_2491,N_2448,N_2450);
and U2492 (N_2492,N_2405,N_2418);
or U2493 (N_2493,N_2428,N_2422);
and U2494 (N_2494,N_2439,N_2449);
nand U2495 (N_2495,N_2420,N_2453);
and U2496 (N_2496,N_2464,N_2404);
or U2497 (N_2497,N_2454,N_2467);
xnor U2498 (N_2498,N_2427,N_2409);
nand U2499 (N_2499,N_2424,N_2407);
nand U2500 (N_2500,N_2435,N_2429);
or U2501 (N_2501,N_2456,N_2469);
nor U2502 (N_2502,N_2462,N_2460);
nand U2503 (N_2503,N_2472,N_2431);
xnor U2504 (N_2504,N_2425,N_2441);
and U2505 (N_2505,N_2410,N_2440);
or U2506 (N_2506,N_2411,N_2443);
and U2507 (N_2507,N_2473,N_2438);
and U2508 (N_2508,N_2446,N_2403);
nor U2509 (N_2509,N_2417,N_2465);
nor U2510 (N_2510,N_2474,N_2413);
xnor U2511 (N_2511,N_2459,N_2408);
or U2512 (N_2512,N_2416,N_2469);
or U2513 (N_2513,N_2457,N_2431);
and U2514 (N_2514,N_2444,N_2440);
and U2515 (N_2515,N_2474,N_2435);
nor U2516 (N_2516,N_2457,N_2413);
or U2517 (N_2517,N_2414,N_2465);
or U2518 (N_2518,N_2468,N_2436);
and U2519 (N_2519,N_2427,N_2462);
nand U2520 (N_2520,N_2451,N_2438);
xor U2521 (N_2521,N_2465,N_2405);
or U2522 (N_2522,N_2429,N_2449);
or U2523 (N_2523,N_2434,N_2426);
and U2524 (N_2524,N_2402,N_2429);
or U2525 (N_2525,N_2424,N_2403);
nand U2526 (N_2526,N_2414,N_2416);
or U2527 (N_2527,N_2439,N_2460);
nor U2528 (N_2528,N_2436,N_2460);
or U2529 (N_2529,N_2461,N_2448);
or U2530 (N_2530,N_2433,N_2446);
and U2531 (N_2531,N_2412,N_2461);
nand U2532 (N_2532,N_2453,N_2435);
or U2533 (N_2533,N_2447,N_2463);
and U2534 (N_2534,N_2429,N_2473);
or U2535 (N_2535,N_2466,N_2410);
nor U2536 (N_2536,N_2436,N_2471);
xor U2537 (N_2537,N_2449,N_2446);
nor U2538 (N_2538,N_2422,N_2406);
or U2539 (N_2539,N_2467,N_2425);
and U2540 (N_2540,N_2432,N_2419);
nand U2541 (N_2541,N_2452,N_2434);
or U2542 (N_2542,N_2426,N_2438);
nor U2543 (N_2543,N_2472,N_2449);
xor U2544 (N_2544,N_2448,N_2400);
xor U2545 (N_2545,N_2422,N_2412);
nor U2546 (N_2546,N_2468,N_2472);
nand U2547 (N_2547,N_2473,N_2423);
nand U2548 (N_2548,N_2406,N_2417);
nand U2549 (N_2549,N_2455,N_2419);
or U2550 (N_2550,N_2495,N_2548);
or U2551 (N_2551,N_2537,N_2476);
xnor U2552 (N_2552,N_2542,N_2515);
nand U2553 (N_2553,N_2538,N_2485);
and U2554 (N_2554,N_2481,N_2516);
or U2555 (N_2555,N_2480,N_2475);
or U2556 (N_2556,N_2482,N_2518);
or U2557 (N_2557,N_2510,N_2541);
or U2558 (N_2558,N_2533,N_2501);
nor U2559 (N_2559,N_2490,N_2502);
nand U2560 (N_2560,N_2498,N_2489);
nand U2561 (N_2561,N_2499,N_2539);
and U2562 (N_2562,N_2530,N_2494);
xor U2563 (N_2563,N_2524,N_2503);
nor U2564 (N_2564,N_2488,N_2513);
nor U2565 (N_2565,N_2483,N_2527);
and U2566 (N_2566,N_2500,N_2497);
or U2567 (N_2567,N_2544,N_2523);
nor U2568 (N_2568,N_2519,N_2504);
or U2569 (N_2569,N_2514,N_2491);
or U2570 (N_2570,N_2522,N_2545);
nor U2571 (N_2571,N_2493,N_2478);
and U2572 (N_2572,N_2546,N_2536);
nand U2573 (N_2573,N_2532,N_2484);
or U2574 (N_2574,N_2549,N_2531);
and U2575 (N_2575,N_2526,N_2529);
nor U2576 (N_2576,N_2508,N_2543);
nor U2577 (N_2577,N_2479,N_2511);
or U2578 (N_2578,N_2487,N_2477);
nor U2579 (N_2579,N_2509,N_2534);
xor U2580 (N_2580,N_2535,N_2517);
nand U2581 (N_2581,N_2528,N_2520);
or U2582 (N_2582,N_2496,N_2540);
or U2583 (N_2583,N_2512,N_2492);
nor U2584 (N_2584,N_2507,N_2506);
nor U2585 (N_2585,N_2505,N_2521);
nor U2586 (N_2586,N_2547,N_2525);
or U2587 (N_2587,N_2486,N_2502);
nand U2588 (N_2588,N_2497,N_2524);
and U2589 (N_2589,N_2476,N_2549);
xnor U2590 (N_2590,N_2493,N_2513);
nor U2591 (N_2591,N_2486,N_2524);
and U2592 (N_2592,N_2524,N_2514);
nor U2593 (N_2593,N_2493,N_2506);
nand U2594 (N_2594,N_2503,N_2548);
nand U2595 (N_2595,N_2484,N_2503);
nor U2596 (N_2596,N_2482,N_2504);
nor U2597 (N_2597,N_2539,N_2477);
or U2598 (N_2598,N_2480,N_2515);
and U2599 (N_2599,N_2510,N_2487);
nor U2600 (N_2600,N_2507,N_2505);
or U2601 (N_2601,N_2538,N_2547);
xnor U2602 (N_2602,N_2535,N_2539);
and U2603 (N_2603,N_2533,N_2487);
nand U2604 (N_2604,N_2479,N_2478);
xor U2605 (N_2605,N_2540,N_2536);
nand U2606 (N_2606,N_2533,N_2525);
nor U2607 (N_2607,N_2508,N_2493);
or U2608 (N_2608,N_2499,N_2486);
or U2609 (N_2609,N_2507,N_2544);
nor U2610 (N_2610,N_2477,N_2507);
or U2611 (N_2611,N_2484,N_2505);
nor U2612 (N_2612,N_2477,N_2549);
nand U2613 (N_2613,N_2509,N_2513);
nor U2614 (N_2614,N_2485,N_2546);
and U2615 (N_2615,N_2476,N_2534);
xnor U2616 (N_2616,N_2528,N_2527);
and U2617 (N_2617,N_2538,N_2503);
nor U2618 (N_2618,N_2523,N_2547);
xnor U2619 (N_2619,N_2540,N_2502);
xor U2620 (N_2620,N_2476,N_2548);
xor U2621 (N_2621,N_2489,N_2538);
nor U2622 (N_2622,N_2501,N_2477);
nor U2623 (N_2623,N_2522,N_2508);
and U2624 (N_2624,N_2523,N_2482);
and U2625 (N_2625,N_2622,N_2558);
or U2626 (N_2626,N_2574,N_2572);
nor U2627 (N_2627,N_2623,N_2600);
nor U2628 (N_2628,N_2593,N_2585);
or U2629 (N_2629,N_2596,N_2559);
and U2630 (N_2630,N_2564,N_2556);
or U2631 (N_2631,N_2588,N_2553);
nand U2632 (N_2632,N_2601,N_2618);
nor U2633 (N_2633,N_2598,N_2604);
nor U2634 (N_2634,N_2560,N_2555);
nand U2635 (N_2635,N_2569,N_2614);
nor U2636 (N_2636,N_2602,N_2617);
nor U2637 (N_2637,N_2619,N_2580);
xor U2638 (N_2638,N_2608,N_2551);
nand U2639 (N_2639,N_2550,N_2595);
or U2640 (N_2640,N_2565,N_2568);
and U2641 (N_2641,N_2563,N_2613);
and U2642 (N_2642,N_2599,N_2612);
nand U2643 (N_2643,N_2582,N_2594);
or U2644 (N_2644,N_2557,N_2567);
and U2645 (N_2645,N_2552,N_2571);
or U2646 (N_2646,N_2573,N_2609);
nand U2647 (N_2647,N_2616,N_2581);
or U2648 (N_2648,N_2611,N_2562);
or U2649 (N_2649,N_2603,N_2624);
xor U2650 (N_2650,N_2587,N_2561);
nor U2651 (N_2651,N_2605,N_2610);
and U2652 (N_2652,N_2592,N_2607);
nand U2653 (N_2653,N_2577,N_2606);
and U2654 (N_2654,N_2554,N_2590);
or U2655 (N_2655,N_2578,N_2579);
nand U2656 (N_2656,N_2597,N_2615);
or U2657 (N_2657,N_2575,N_2591);
nand U2658 (N_2658,N_2621,N_2589);
nor U2659 (N_2659,N_2566,N_2583);
nor U2660 (N_2660,N_2576,N_2586);
nor U2661 (N_2661,N_2620,N_2570);
and U2662 (N_2662,N_2584,N_2587);
nor U2663 (N_2663,N_2581,N_2620);
nand U2664 (N_2664,N_2596,N_2562);
nand U2665 (N_2665,N_2572,N_2580);
or U2666 (N_2666,N_2558,N_2567);
and U2667 (N_2667,N_2564,N_2550);
nand U2668 (N_2668,N_2592,N_2583);
nor U2669 (N_2669,N_2570,N_2559);
nand U2670 (N_2670,N_2607,N_2608);
and U2671 (N_2671,N_2593,N_2624);
or U2672 (N_2672,N_2608,N_2616);
and U2673 (N_2673,N_2604,N_2572);
and U2674 (N_2674,N_2593,N_2580);
or U2675 (N_2675,N_2614,N_2558);
nand U2676 (N_2676,N_2575,N_2606);
nand U2677 (N_2677,N_2597,N_2581);
and U2678 (N_2678,N_2616,N_2623);
and U2679 (N_2679,N_2581,N_2563);
xnor U2680 (N_2680,N_2566,N_2564);
nand U2681 (N_2681,N_2554,N_2592);
nand U2682 (N_2682,N_2572,N_2581);
and U2683 (N_2683,N_2613,N_2576);
nand U2684 (N_2684,N_2578,N_2606);
or U2685 (N_2685,N_2580,N_2624);
and U2686 (N_2686,N_2578,N_2586);
nor U2687 (N_2687,N_2584,N_2616);
and U2688 (N_2688,N_2570,N_2564);
or U2689 (N_2689,N_2608,N_2594);
and U2690 (N_2690,N_2599,N_2589);
nand U2691 (N_2691,N_2603,N_2612);
nor U2692 (N_2692,N_2571,N_2562);
nor U2693 (N_2693,N_2615,N_2593);
nor U2694 (N_2694,N_2597,N_2623);
xnor U2695 (N_2695,N_2602,N_2557);
nand U2696 (N_2696,N_2623,N_2601);
and U2697 (N_2697,N_2577,N_2585);
or U2698 (N_2698,N_2602,N_2598);
and U2699 (N_2699,N_2611,N_2559);
and U2700 (N_2700,N_2681,N_2669);
nor U2701 (N_2701,N_2659,N_2666);
and U2702 (N_2702,N_2636,N_2695);
nor U2703 (N_2703,N_2673,N_2632);
nand U2704 (N_2704,N_2641,N_2640);
nor U2705 (N_2705,N_2686,N_2692);
nor U2706 (N_2706,N_2680,N_2690);
nor U2707 (N_2707,N_2644,N_2672);
and U2708 (N_2708,N_2633,N_2675);
or U2709 (N_2709,N_2691,N_2689);
and U2710 (N_2710,N_2626,N_2645);
nand U2711 (N_2711,N_2650,N_2667);
or U2712 (N_2712,N_2671,N_2696);
xnor U2713 (N_2713,N_2656,N_2627);
xnor U2714 (N_2714,N_2654,N_2651);
nor U2715 (N_2715,N_2646,N_2628);
and U2716 (N_2716,N_2648,N_2658);
or U2717 (N_2717,N_2668,N_2643);
and U2718 (N_2718,N_2642,N_2649);
nor U2719 (N_2719,N_2685,N_2655);
nand U2720 (N_2720,N_2661,N_2664);
nand U2721 (N_2721,N_2637,N_2677);
and U2722 (N_2722,N_2674,N_2676);
nor U2723 (N_2723,N_2660,N_2635);
nand U2724 (N_2724,N_2682,N_2687);
nand U2725 (N_2725,N_2693,N_2625);
nand U2726 (N_2726,N_2630,N_2697);
nor U2727 (N_2727,N_2694,N_2678);
nor U2728 (N_2728,N_2665,N_2639);
and U2729 (N_2729,N_2688,N_2631);
nor U2730 (N_2730,N_2657,N_2698);
nand U2731 (N_2731,N_2647,N_2638);
nor U2732 (N_2732,N_2679,N_2634);
nand U2733 (N_2733,N_2683,N_2670);
or U2734 (N_2734,N_2652,N_2663);
xnor U2735 (N_2735,N_2629,N_2653);
xor U2736 (N_2736,N_2662,N_2699);
nand U2737 (N_2737,N_2684,N_2633);
nand U2738 (N_2738,N_2679,N_2683);
or U2739 (N_2739,N_2628,N_2635);
nand U2740 (N_2740,N_2650,N_2687);
xor U2741 (N_2741,N_2675,N_2656);
nor U2742 (N_2742,N_2652,N_2669);
nand U2743 (N_2743,N_2695,N_2659);
nor U2744 (N_2744,N_2677,N_2633);
and U2745 (N_2745,N_2627,N_2680);
nor U2746 (N_2746,N_2687,N_2698);
nand U2747 (N_2747,N_2659,N_2650);
and U2748 (N_2748,N_2651,N_2690);
nor U2749 (N_2749,N_2648,N_2697);
and U2750 (N_2750,N_2685,N_2668);
nor U2751 (N_2751,N_2653,N_2674);
and U2752 (N_2752,N_2637,N_2669);
and U2753 (N_2753,N_2643,N_2684);
and U2754 (N_2754,N_2669,N_2648);
xor U2755 (N_2755,N_2644,N_2638);
nand U2756 (N_2756,N_2679,N_2671);
nor U2757 (N_2757,N_2650,N_2651);
nor U2758 (N_2758,N_2692,N_2632);
and U2759 (N_2759,N_2680,N_2655);
nor U2760 (N_2760,N_2676,N_2682);
and U2761 (N_2761,N_2691,N_2682);
or U2762 (N_2762,N_2694,N_2683);
and U2763 (N_2763,N_2673,N_2634);
nor U2764 (N_2764,N_2683,N_2636);
or U2765 (N_2765,N_2640,N_2678);
or U2766 (N_2766,N_2644,N_2695);
and U2767 (N_2767,N_2674,N_2666);
and U2768 (N_2768,N_2655,N_2638);
or U2769 (N_2769,N_2680,N_2664);
or U2770 (N_2770,N_2671,N_2664);
and U2771 (N_2771,N_2650,N_2632);
nand U2772 (N_2772,N_2673,N_2686);
and U2773 (N_2773,N_2639,N_2648);
or U2774 (N_2774,N_2650,N_2674);
or U2775 (N_2775,N_2710,N_2762);
and U2776 (N_2776,N_2754,N_2752);
and U2777 (N_2777,N_2741,N_2772);
nor U2778 (N_2778,N_2711,N_2749);
and U2779 (N_2779,N_2755,N_2736);
and U2780 (N_2780,N_2757,N_2761);
and U2781 (N_2781,N_2702,N_2759);
or U2782 (N_2782,N_2745,N_2735);
nor U2783 (N_2783,N_2768,N_2773);
or U2784 (N_2784,N_2766,N_2729);
nor U2785 (N_2785,N_2706,N_2743);
nand U2786 (N_2786,N_2756,N_2769);
nand U2787 (N_2787,N_2753,N_2712);
or U2788 (N_2788,N_2765,N_2716);
nor U2789 (N_2789,N_2701,N_2714);
or U2790 (N_2790,N_2732,N_2771);
or U2791 (N_2791,N_2707,N_2767);
and U2792 (N_2792,N_2748,N_2728);
nand U2793 (N_2793,N_2760,N_2740);
nand U2794 (N_2794,N_2705,N_2725);
nor U2795 (N_2795,N_2734,N_2715);
nor U2796 (N_2796,N_2750,N_2703);
nor U2797 (N_2797,N_2739,N_2717);
nand U2798 (N_2798,N_2724,N_2727);
nand U2799 (N_2799,N_2751,N_2742);
and U2800 (N_2800,N_2721,N_2704);
nor U2801 (N_2801,N_2764,N_2774);
nor U2802 (N_2802,N_2730,N_2763);
and U2803 (N_2803,N_2709,N_2700);
nor U2804 (N_2804,N_2708,N_2722);
or U2805 (N_2805,N_2718,N_2713);
or U2806 (N_2806,N_2747,N_2746);
and U2807 (N_2807,N_2719,N_2738);
or U2808 (N_2808,N_2731,N_2720);
or U2809 (N_2809,N_2770,N_2758);
and U2810 (N_2810,N_2726,N_2733);
and U2811 (N_2811,N_2723,N_2744);
and U2812 (N_2812,N_2737,N_2740);
nor U2813 (N_2813,N_2711,N_2754);
or U2814 (N_2814,N_2722,N_2704);
nor U2815 (N_2815,N_2760,N_2756);
nor U2816 (N_2816,N_2753,N_2707);
nor U2817 (N_2817,N_2700,N_2739);
or U2818 (N_2818,N_2700,N_2718);
or U2819 (N_2819,N_2719,N_2706);
nand U2820 (N_2820,N_2734,N_2728);
nand U2821 (N_2821,N_2718,N_2772);
nor U2822 (N_2822,N_2708,N_2729);
and U2823 (N_2823,N_2707,N_2717);
or U2824 (N_2824,N_2755,N_2712);
nor U2825 (N_2825,N_2720,N_2725);
nor U2826 (N_2826,N_2709,N_2738);
nand U2827 (N_2827,N_2715,N_2769);
and U2828 (N_2828,N_2716,N_2771);
and U2829 (N_2829,N_2709,N_2764);
nand U2830 (N_2830,N_2703,N_2731);
and U2831 (N_2831,N_2709,N_2749);
and U2832 (N_2832,N_2729,N_2743);
nor U2833 (N_2833,N_2724,N_2769);
nor U2834 (N_2834,N_2745,N_2756);
nor U2835 (N_2835,N_2766,N_2711);
and U2836 (N_2836,N_2721,N_2764);
nor U2837 (N_2837,N_2716,N_2711);
nor U2838 (N_2838,N_2740,N_2700);
or U2839 (N_2839,N_2753,N_2761);
nor U2840 (N_2840,N_2713,N_2772);
and U2841 (N_2841,N_2755,N_2714);
or U2842 (N_2842,N_2700,N_2707);
nor U2843 (N_2843,N_2761,N_2772);
nor U2844 (N_2844,N_2710,N_2756);
or U2845 (N_2845,N_2717,N_2767);
and U2846 (N_2846,N_2740,N_2748);
nor U2847 (N_2847,N_2773,N_2772);
nand U2848 (N_2848,N_2754,N_2763);
and U2849 (N_2849,N_2755,N_2726);
nor U2850 (N_2850,N_2814,N_2775);
or U2851 (N_2851,N_2836,N_2790);
and U2852 (N_2852,N_2808,N_2820);
xnor U2853 (N_2853,N_2804,N_2816);
or U2854 (N_2854,N_2835,N_2791);
nor U2855 (N_2855,N_2778,N_2789);
nor U2856 (N_2856,N_2831,N_2846);
nor U2857 (N_2857,N_2830,N_2783);
nand U2858 (N_2858,N_2832,N_2822);
and U2859 (N_2859,N_2795,N_2839);
xnor U2860 (N_2860,N_2779,N_2780);
and U2861 (N_2861,N_2802,N_2801);
nor U2862 (N_2862,N_2818,N_2793);
and U2863 (N_2863,N_2826,N_2813);
nand U2864 (N_2864,N_2842,N_2841);
nor U2865 (N_2865,N_2798,N_2845);
or U2866 (N_2866,N_2799,N_2781);
nand U2867 (N_2867,N_2815,N_2838);
and U2868 (N_2868,N_2807,N_2823);
or U2869 (N_2869,N_2787,N_2788);
nor U2870 (N_2870,N_2800,N_2821);
and U2871 (N_2871,N_2805,N_2829);
xor U2872 (N_2872,N_2819,N_2786);
nand U2873 (N_2873,N_2810,N_2784);
nor U2874 (N_2874,N_2824,N_2840);
nand U2875 (N_2875,N_2834,N_2843);
or U2876 (N_2876,N_2811,N_2794);
nand U2877 (N_2877,N_2776,N_2844);
and U2878 (N_2878,N_2833,N_2828);
nor U2879 (N_2879,N_2827,N_2825);
or U2880 (N_2880,N_2785,N_2796);
or U2881 (N_2881,N_2803,N_2777);
nand U2882 (N_2882,N_2806,N_2817);
or U2883 (N_2883,N_2849,N_2848);
nand U2884 (N_2884,N_2809,N_2782);
nor U2885 (N_2885,N_2847,N_2797);
or U2886 (N_2886,N_2792,N_2812);
nor U2887 (N_2887,N_2837,N_2825);
or U2888 (N_2888,N_2814,N_2833);
nor U2889 (N_2889,N_2802,N_2776);
or U2890 (N_2890,N_2818,N_2800);
and U2891 (N_2891,N_2781,N_2828);
and U2892 (N_2892,N_2836,N_2805);
nand U2893 (N_2893,N_2787,N_2775);
nor U2894 (N_2894,N_2790,N_2798);
and U2895 (N_2895,N_2848,N_2835);
nor U2896 (N_2896,N_2786,N_2805);
nand U2897 (N_2897,N_2803,N_2829);
xor U2898 (N_2898,N_2834,N_2797);
nand U2899 (N_2899,N_2806,N_2827);
nor U2900 (N_2900,N_2812,N_2823);
nand U2901 (N_2901,N_2842,N_2832);
or U2902 (N_2902,N_2788,N_2802);
nor U2903 (N_2903,N_2829,N_2826);
nor U2904 (N_2904,N_2787,N_2780);
xnor U2905 (N_2905,N_2821,N_2848);
and U2906 (N_2906,N_2838,N_2780);
nand U2907 (N_2907,N_2815,N_2792);
and U2908 (N_2908,N_2798,N_2775);
nor U2909 (N_2909,N_2779,N_2778);
nor U2910 (N_2910,N_2792,N_2785);
or U2911 (N_2911,N_2775,N_2825);
and U2912 (N_2912,N_2820,N_2825);
or U2913 (N_2913,N_2796,N_2808);
nand U2914 (N_2914,N_2847,N_2788);
nand U2915 (N_2915,N_2780,N_2809);
nor U2916 (N_2916,N_2844,N_2842);
or U2917 (N_2917,N_2814,N_2832);
or U2918 (N_2918,N_2795,N_2832);
nand U2919 (N_2919,N_2807,N_2837);
xor U2920 (N_2920,N_2841,N_2786);
nand U2921 (N_2921,N_2806,N_2820);
nand U2922 (N_2922,N_2787,N_2829);
nand U2923 (N_2923,N_2804,N_2792);
nand U2924 (N_2924,N_2834,N_2802);
or U2925 (N_2925,N_2883,N_2867);
and U2926 (N_2926,N_2894,N_2860);
and U2927 (N_2927,N_2906,N_2902);
nor U2928 (N_2928,N_2919,N_2898);
xnor U2929 (N_2929,N_2921,N_2862);
or U2930 (N_2930,N_2915,N_2923);
nor U2931 (N_2931,N_2904,N_2899);
or U2932 (N_2932,N_2891,N_2878);
and U2933 (N_2933,N_2874,N_2877);
and U2934 (N_2934,N_2893,N_2869);
nor U2935 (N_2935,N_2924,N_2908);
nand U2936 (N_2936,N_2864,N_2901);
nand U2937 (N_2937,N_2900,N_2870);
nand U2938 (N_2938,N_2873,N_2911);
and U2939 (N_2939,N_2855,N_2889);
and U2940 (N_2940,N_2851,N_2909);
and U2941 (N_2941,N_2875,N_2897);
xor U2942 (N_2942,N_2916,N_2922);
nor U2943 (N_2943,N_2881,N_2910);
and U2944 (N_2944,N_2880,N_2856);
nand U2945 (N_2945,N_2896,N_2884);
nand U2946 (N_2946,N_2871,N_2872);
and U2947 (N_2947,N_2885,N_2912);
and U2948 (N_2948,N_2852,N_2850);
nand U2949 (N_2949,N_2895,N_2892);
nor U2950 (N_2950,N_2859,N_2865);
xor U2951 (N_2951,N_2866,N_2913);
xnor U2952 (N_2952,N_2917,N_2886);
xnor U2953 (N_2953,N_2853,N_2890);
xnor U2954 (N_2954,N_2879,N_2918);
or U2955 (N_2955,N_2903,N_2876);
or U2956 (N_2956,N_2920,N_2882);
xor U2957 (N_2957,N_2905,N_2857);
nand U2958 (N_2958,N_2907,N_2888);
nand U2959 (N_2959,N_2858,N_2887);
xor U2960 (N_2960,N_2914,N_2868);
nor U2961 (N_2961,N_2863,N_2854);
or U2962 (N_2962,N_2861,N_2856);
nor U2963 (N_2963,N_2862,N_2850);
and U2964 (N_2964,N_2887,N_2857);
and U2965 (N_2965,N_2910,N_2896);
nand U2966 (N_2966,N_2918,N_2905);
and U2967 (N_2967,N_2884,N_2892);
and U2968 (N_2968,N_2855,N_2883);
and U2969 (N_2969,N_2912,N_2869);
or U2970 (N_2970,N_2878,N_2906);
nand U2971 (N_2971,N_2888,N_2873);
and U2972 (N_2972,N_2868,N_2856);
or U2973 (N_2973,N_2919,N_2866);
and U2974 (N_2974,N_2911,N_2874);
nand U2975 (N_2975,N_2893,N_2918);
nor U2976 (N_2976,N_2891,N_2918);
nor U2977 (N_2977,N_2924,N_2858);
and U2978 (N_2978,N_2878,N_2892);
xor U2979 (N_2979,N_2922,N_2921);
nor U2980 (N_2980,N_2889,N_2896);
nor U2981 (N_2981,N_2903,N_2869);
or U2982 (N_2982,N_2904,N_2902);
nor U2983 (N_2983,N_2882,N_2868);
nor U2984 (N_2984,N_2922,N_2883);
nor U2985 (N_2985,N_2911,N_2920);
nor U2986 (N_2986,N_2899,N_2886);
or U2987 (N_2987,N_2852,N_2904);
and U2988 (N_2988,N_2911,N_2879);
nor U2989 (N_2989,N_2872,N_2911);
or U2990 (N_2990,N_2880,N_2869);
xor U2991 (N_2991,N_2875,N_2898);
nand U2992 (N_2992,N_2860,N_2850);
nor U2993 (N_2993,N_2916,N_2902);
or U2994 (N_2994,N_2898,N_2924);
nand U2995 (N_2995,N_2885,N_2877);
nor U2996 (N_2996,N_2908,N_2919);
nand U2997 (N_2997,N_2914,N_2897);
nor U2998 (N_2998,N_2861,N_2878);
and U2999 (N_2999,N_2879,N_2893);
and UO_0 (O_0,N_2999,N_2961);
nor UO_1 (O_1,N_2980,N_2928);
xnor UO_2 (O_2,N_2992,N_2994);
or UO_3 (O_3,N_2981,N_2952);
and UO_4 (O_4,N_2955,N_2932);
nand UO_5 (O_5,N_2960,N_2974);
or UO_6 (O_6,N_2979,N_2971);
nor UO_7 (O_7,N_2946,N_2951);
xor UO_8 (O_8,N_2964,N_2963);
or UO_9 (O_9,N_2935,N_2941);
and UO_10 (O_10,N_2993,N_2985);
or UO_11 (O_11,N_2953,N_2986);
nand UO_12 (O_12,N_2977,N_2968);
nand UO_13 (O_13,N_2933,N_2959);
nand UO_14 (O_14,N_2996,N_2965);
or UO_15 (O_15,N_2970,N_2930);
and UO_16 (O_16,N_2990,N_2984);
nor UO_17 (O_17,N_2954,N_2972);
nand UO_18 (O_18,N_2945,N_2982);
nor UO_19 (O_19,N_2949,N_2926);
nor UO_20 (O_20,N_2978,N_2934);
nor UO_21 (O_21,N_2997,N_2929);
nor UO_22 (O_22,N_2939,N_2958);
nor UO_23 (O_23,N_2957,N_2938);
nor UO_24 (O_24,N_2950,N_2998);
or UO_25 (O_25,N_2969,N_2962);
nand UO_26 (O_26,N_2942,N_2936);
nor UO_27 (O_27,N_2983,N_2976);
and UO_28 (O_28,N_2943,N_2940);
nor UO_29 (O_29,N_2987,N_2991);
or UO_30 (O_30,N_2988,N_2927);
and UO_31 (O_31,N_2947,N_2973);
or UO_32 (O_32,N_2989,N_2975);
xor UO_33 (O_33,N_2966,N_2948);
or UO_34 (O_34,N_2956,N_2944);
and UO_35 (O_35,N_2967,N_2937);
nor UO_36 (O_36,N_2995,N_2931);
nor UO_37 (O_37,N_2925,N_2958);
or UO_38 (O_38,N_2968,N_2937);
and UO_39 (O_39,N_2956,N_2973);
nor UO_40 (O_40,N_2996,N_2932);
and UO_41 (O_41,N_2947,N_2969);
and UO_42 (O_42,N_2952,N_2966);
nor UO_43 (O_43,N_2956,N_2974);
nor UO_44 (O_44,N_2956,N_2997);
nor UO_45 (O_45,N_2955,N_2946);
or UO_46 (O_46,N_2927,N_2996);
nand UO_47 (O_47,N_2952,N_2971);
and UO_48 (O_48,N_2978,N_2941);
nor UO_49 (O_49,N_2941,N_2959);
nor UO_50 (O_50,N_2941,N_2997);
and UO_51 (O_51,N_2960,N_2942);
nand UO_52 (O_52,N_2991,N_2980);
nand UO_53 (O_53,N_2984,N_2995);
or UO_54 (O_54,N_2987,N_2982);
or UO_55 (O_55,N_2985,N_2937);
or UO_56 (O_56,N_2935,N_2956);
and UO_57 (O_57,N_2995,N_2974);
or UO_58 (O_58,N_2945,N_2961);
nor UO_59 (O_59,N_2946,N_2929);
xnor UO_60 (O_60,N_2949,N_2971);
or UO_61 (O_61,N_2999,N_2926);
nand UO_62 (O_62,N_2992,N_2952);
or UO_63 (O_63,N_2925,N_2967);
nor UO_64 (O_64,N_2985,N_2964);
nor UO_65 (O_65,N_2938,N_2965);
nor UO_66 (O_66,N_2930,N_2936);
nor UO_67 (O_67,N_2995,N_2934);
nor UO_68 (O_68,N_2945,N_2939);
xnor UO_69 (O_69,N_2969,N_2981);
nand UO_70 (O_70,N_2929,N_2960);
nor UO_71 (O_71,N_2959,N_2997);
nand UO_72 (O_72,N_2952,N_2953);
nor UO_73 (O_73,N_2960,N_2937);
nand UO_74 (O_74,N_2930,N_2993);
nand UO_75 (O_75,N_2937,N_2992);
xnor UO_76 (O_76,N_2928,N_2951);
and UO_77 (O_77,N_2960,N_2949);
and UO_78 (O_78,N_2959,N_2944);
nand UO_79 (O_79,N_2965,N_2977);
xor UO_80 (O_80,N_2930,N_2969);
or UO_81 (O_81,N_2970,N_2979);
nor UO_82 (O_82,N_2964,N_2943);
or UO_83 (O_83,N_2983,N_2988);
nand UO_84 (O_84,N_2925,N_2986);
and UO_85 (O_85,N_2976,N_2965);
and UO_86 (O_86,N_2947,N_2976);
nand UO_87 (O_87,N_2972,N_2968);
and UO_88 (O_88,N_2963,N_2939);
or UO_89 (O_89,N_2955,N_2975);
and UO_90 (O_90,N_2969,N_2953);
nor UO_91 (O_91,N_2994,N_2934);
xnor UO_92 (O_92,N_2925,N_2968);
xor UO_93 (O_93,N_2968,N_2956);
and UO_94 (O_94,N_2970,N_2937);
or UO_95 (O_95,N_2994,N_2965);
nor UO_96 (O_96,N_2984,N_2973);
and UO_97 (O_97,N_2983,N_2967);
or UO_98 (O_98,N_2977,N_2997);
nand UO_99 (O_99,N_2938,N_2974);
or UO_100 (O_100,N_2983,N_2929);
or UO_101 (O_101,N_2950,N_2993);
nand UO_102 (O_102,N_2957,N_2959);
nor UO_103 (O_103,N_2950,N_2927);
nand UO_104 (O_104,N_2936,N_2986);
nand UO_105 (O_105,N_2939,N_2933);
xor UO_106 (O_106,N_2960,N_2932);
or UO_107 (O_107,N_2975,N_2998);
nand UO_108 (O_108,N_2984,N_2932);
and UO_109 (O_109,N_2930,N_2979);
nor UO_110 (O_110,N_2948,N_2977);
or UO_111 (O_111,N_2934,N_2935);
xnor UO_112 (O_112,N_2958,N_2929);
nor UO_113 (O_113,N_2944,N_2980);
nand UO_114 (O_114,N_2990,N_2959);
nand UO_115 (O_115,N_2975,N_2973);
or UO_116 (O_116,N_2969,N_2963);
nor UO_117 (O_117,N_2942,N_2986);
or UO_118 (O_118,N_2965,N_2956);
or UO_119 (O_119,N_2944,N_2972);
nor UO_120 (O_120,N_2937,N_2957);
or UO_121 (O_121,N_2955,N_2966);
nor UO_122 (O_122,N_2952,N_2954);
xnor UO_123 (O_123,N_2931,N_2950);
xnor UO_124 (O_124,N_2928,N_2965);
nor UO_125 (O_125,N_2962,N_2978);
nand UO_126 (O_126,N_2954,N_2974);
nor UO_127 (O_127,N_2965,N_2975);
or UO_128 (O_128,N_2948,N_2932);
and UO_129 (O_129,N_2949,N_2935);
or UO_130 (O_130,N_2945,N_2978);
and UO_131 (O_131,N_2991,N_2967);
and UO_132 (O_132,N_2964,N_2987);
or UO_133 (O_133,N_2944,N_2935);
or UO_134 (O_134,N_2930,N_2984);
nand UO_135 (O_135,N_2961,N_2957);
nand UO_136 (O_136,N_2990,N_2975);
or UO_137 (O_137,N_2931,N_2958);
or UO_138 (O_138,N_2957,N_2984);
nor UO_139 (O_139,N_2975,N_2946);
and UO_140 (O_140,N_2978,N_2936);
xor UO_141 (O_141,N_2935,N_2983);
xor UO_142 (O_142,N_2929,N_2944);
and UO_143 (O_143,N_2991,N_2988);
nor UO_144 (O_144,N_2925,N_2931);
and UO_145 (O_145,N_2954,N_2965);
or UO_146 (O_146,N_2991,N_2930);
xor UO_147 (O_147,N_2985,N_2946);
or UO_148 (O_148,N_2983,N_2932);
and UO_149 (O_149,N_2993,N_2962);
nand UO_150 (O_150,N_2970,N_2965);
nand UO_151 (O_151,N_2976,N_2945);
or UO_152 (O_152,N_2995,N_2959);
or UO_153 (O_153,N_2935,N_2987);
and UO_154 (O_154,N_2993,N_2933);
nor UO_155 (O_155,N_2982,N_2927);
nand UO_156 (O_156,N_2939,N_2940);
nor UO_157 (O_157,N_2969,N_2951);
nor UO_158 (O_158,N_2957,N_2949);
nand UO_159 (O_159,N_2980,N_2994);
or UO_160 (O_160,N_2967,N_2953);
and UO_161 (O_161,N_2955,N_2928);
and UO_162 (O_162,N_2935,N_2999);
nor UO_163 (O_163,N_2953,N_2996);
nand UO_164 (O_164,N_2959,N_2976);
nand UO_165 (O_165,N_2963,N_2995);
xor UO_166 (O_166,N_2926,N_2991);
or UO_167 (O_167,N_2929,N_2936);
or UO_168 (O_168,N_2927,N_2953);
xor UO_169 (O_169,N_2996,N_2978);
nand UO_170 (O_170,N_2962,N_2988);
nand UO_171 (O_171,N_2981,N_2999);
and UO_172 (O_172,N_2961,N_2940);
nor UO_173 (O_173,N_2986,N_2981);
or UO_174 (O_174,N_2925,N_2971);
or UO_175 (O_175,N_2925,N_2954);
nand UO_176 (O_176,N_2945,N_2925);
or UO_177 (O_177,N_2930,N_2932);
or UO_178 (O_178,N_2968,N_2992);
nor UO_179 (O_179,N_2990,N_2967);
nand UO_180 (O_180,N_2949,N_2996);
nand UO_181 (O_181,N_2995,N_2996);
or UO_182 (O_182,N_2977,N_2971);
or UO_183 (O_183,N_2983,N_2996);
and UO_184 (O_184,N_2962,N_2949);
and UO_185 (O_185,N_2965,N_2931);
nor UO_186 (O_186,N_2937,N_2934);
or UO_187 (O_187,N_2941,N_2982);
xor UO_188 (O_188,N_2981,N_2994);
and UO_189 (O_189,N_2959,N_2974);
and UO_190 (O_190,N_2988,N_2979);
nor UO_191 (O_191,N_2937,N_2962);
and UO_192 (O_192,N_2931,N_2996);
nor UO_193 (O_193,N_2969,N_2948);
nor UO_194 (O_194,N_2953,N_2934);
nor UO_195 (O_195,N_2926,N_2964);
or UO_196 (O_196,N_2972,N_2982);
and UO_197 (O_197,N_2942,N_2966);
nor UO_198 (O_198,N_2995,N_2977);
or UO_199 (O_199,N_2963,N_2935);
xor UO_200 (O_200,N_2986,N_2959);
or UO_201 (O_201,N_2964,N_2950);
or UO_202 (O_202,N_2936,N_2958);
xnor UO_203 (O_203,N_2949,N_2952);
or UO_204 (O_204,N_2936,N_2949);
or UO_205 (O_205,N_2956,N_2945);
nand UO_206 (O_206,N_2950,N_2968);
and UO_207 (O_207,N_2930,N_2925);
nand UO_208 (O_208,N_2971,N_2942);
and UO_209 (O_209,N_2956,N_2954);
nand UO_210 (O_210,N_2973,N_2953);
nor UO_211 (O_211,N_2936,N_2972);
nand UO_212 (O_212,N_2985,N_2957);
or UO_213 (O_213,N_2925,N_2952);
or UO_214 (O_214,N_2930,N_2998);
nand UO_215 (O_215,N_2953,N_2943);
and UO_216 (O_216,N_2939,N_2968);
nand UO_217 (O_217,N_2983,N_2948);
xnor UO_218 (O_218,N_2995,N_2955);
and UO_219 (O_219,N_2978,N_2939);
or UO_220 (O_220,N_2947,N_2990);
nand UO_221 (O_221,N_2980,N_2951);
and UO_222 (O_222,N_2938,N_2945);
or UO_223 (O_223,N_2956,N_2958);
nand UO_224 (O_224,N_2958,N_2932);
nand UO_225 (O_225,N_2995,N_2956);
or UO_226 (O_226,N_2994,N_2938);
nand UO_227 (O_227,N_2927,N_2994);
nand UO_228 (O_228,N_2925,N_2950);
nor UO_229 (O_229,N_2985,N_2979);
and UO_230 (O_230,N_2959,N_2948);
and UO_231 (O_231,N_2929,N_2966);
nand UO_232 (O_232,N_2941,N_2930);
nand UO_233 (O_233,N_2992,N_2925);
nor UO_234 (O_234,N_2936,N_2957);
xor UO_235 (O_235,N_2954,N_2999);
and UO_236 (O_236,N_2986,N_2990);
or UO_237 (O_237,N_2986,N_2967);
and UO_238 (O_238,N_2960,N_2963);
nor UO_239 (O_239,N_2946,N_2931);
xor UO_240 (O_240,N_2932,N_2965);
nand UO_241 (O_241,N_2980,N_2943);
nand UO_242 (O_242,N_2975,N_2940);
nand UO_243 (O_243,N_2980,N_2959);
nor UO_244 (O_244,N_2966,N_2981);
nor UO_245 (O_245,N_2943,N_2966);
nand UO_246 (O_246,N_2991,N_2982);
nor UO_247 (O_247,N_2974,N_2975);
and UO_248 (O_248,N_2936,N_2959);
and UO_249 (O_249,N_2949,N_2942);
or UO_250 (O_250,N_2997,N_2967);
nand UO_251 (O_251,N_2979,N_2994);
nor UO_252 (O_252,N_2999,N_2978);
and UO_253 (O_253,N_2939,N_2947);
xor UO_254 (O_254,N_2944,N_2933);
and UO_255 (O_255,N_2969,N_2944);
nor UO_256 (O_256,N_2969,N_2985);
nor UO_257 (O_257,N_2943,N_2989);
nor UO_258 (O_258,N_2966,N_2957);
nand UO_259 (O_259,N_2942,N_2972);
xnor UO_260 (O_260,N_2943,N_2928);
or UO_261 (O_261,N_2933,N_2952);
or UO_262 (O_262,N_2933,N_2985);
or UO_263 (O_263,N_2977,N_2962);
nand UO_264 (O_264,N_2940,N_2998);
or UO_265 (O_265,N_2978,N_2998);
and UO_266 (O_266,N_2997,N_2947);
nand UO_267 (O_267,N_2963,N_2992);
nand UO_268 (O_268,N_2979,N_2992);
nor UO_269 (O_269,N_2939,N_2942);
nor UO_270 (O_270,N_2964,N_2978);
nand UO_271 (O_271,N_2963,N_2989);
or UO_272 (O_272,N_2957,N_2991);
xnor UO_273 (O_273,N_2964,N_2938);
or UO_274 (O_274,N_2986,N_2965);
or UO_275 (O_275,N_2932,N_2946);
or UO_276 (O_276,N_2952,N_2951);
and UO_277 (O_277,N_2999,N_2931);
and UO_278 (O_278,N_2961,N_2938);
and UO_279 (O_279,N_2927,N_2938);
and UO_280 (O_280,N_2952,N_2939);
nand UO_281 (O_281,N_2930,N_2992);
nand UO_282 (O_282,N_2925,N_2947);
nand UO_283 (O_283,N_2959,N_2940);
and UO_284 (O_284,N_2959,N_2950);
nand UO_285 (O_285,N_2964,N_2956);
nand UO_286 (O_286,N_2977,N_2991);
nand UO_287 (O_287,N_2937,N_2979);
nor UO_288 (O_288,N_2947,N_2995);
and UO_289 (O_289,N_2966,N_2984);
and UO_290 (O_290,N_2984,N_2933);
and UO_291 (O_291,N_2938,N_2991);
or UO_292 (O_292,N_2954,N_2981);
or UO_293 (O_293,N_2949,N_2937);
or UO_294 (O_294,N_2995,N_2969);
or UO_295 (O_295,N_2938,N_2985);
or UO_296 (O_296,N_2927,N_2941);
or UO_297 (O_297,N_2989,N_2955);
and UO_298 (O_298,N_2989,N_2936);
or UO_299 (O_299,N_2976,N_2925);
nand UO_300 (O_300,N_2966,N_2934);
and UO_301 (O_301,N_2931,N_2926);
or UO_302 (O_302,N_2929,N_2980);
xor UO_303 (O_303,N_2951,N_2931);
xnor UO_304 (O_304,N_2977,N_2951);
or UO_305 (O_305,N_2995,N_2950);
or UO_306 (O_306,N_2957,N_2965);
or UO_307 (O_307,N_2975,N_2985);
and UO_308 (O_308,N_2950,N_2992);
or UO_309 (O_309,N_2934,N_2976);
xor UO_310 (O_310,N_2954,N_2969);
nand UO_311 (O_311,N_2980,N_2988);
xnor UO_312 (O_312,N_2940,N_2944);
or UO_313 (O_313,N_2983,N_2991);
and UO_314 (O_314,N_2952,N_2998);
and UO_315 (O_315,N_2932,N_2951);
nor UO_316 (O_316,N_2949,N_2994);
and UO_317 (O_317,N_2966,N_2931);
nand UO_318 (O_318,N_2964,N_2990);
and UO_319 (O_319,N_2965,N_2933);
and UO_320 (O_320,N_2939,N_2980);
nor UO_321 (O_321,N_2952,N_2968);
xnor UO_322 (O_322,N_2930,N_2937);
and UO_323 (O_323,N_2967,N_2964);
or UO_324 (O_324,N_2946,N_2978);
nor UO_325 (O_325,N_2999,N_2998);
nor UO_326 (O_326,N_2960,N_2979);
or UO_327 (O_327,N_2932,N_2935);
and UO_328 (O_328,N_2977,N_2932);
xor UO_329 (O_329,N_2936,N_2988);
nand UO_330 (O_330,N_2991,N_2997);
and UO_331 (O_331,N_2976,N_2930);
nor UO_332 (O_332,N_2975,N_2937);
and UO_333 (O_333,N_2981,N_2928);
or UO_334 (O_334,N_2946,N_2988);
nand UO_335 (O_335,N_2987,N_2976);
nor UO_336 (O_336,N_2984,N_2955);
and UO_337 (O_337,N_2996,N_2952);
nand UO_338 (O_338,N_2954,N_2957);
xor UO_339 (O_339,N_2997,N_2961);
or UO_340 (O_340,N_2984,N_2999);
xnor UO_341 (O_341,N_2948,N_2944);
nor UO_342 (O_342,N_2993,N_2988);
nor UO_343 (O_343,N_2926,N_2948);
xnor UO_344 (O_344,N_2994,N_2955);
and UO_345 (O_345,N_2949,N_2969);
nor UO_346 (O_346,N_2946,N_2933);
or UO_347 (O_347,N_2968,N_2929);
nand UO_348 (O_348,N_2954,N_2960);
nor UO_349 (O_349,N_2988,N_2933);
nand UO_350 (O_350,N_2929,N_2926);
xnor UO_351 (O_351,N_2952,N_2989);
nor UO_352 (O_352,N_2961,N_2967);
or UO_353 (O_353,N_2958,N_2950);
and UO_354 (O_354,N_2943,N_2965);
and UO_355 (O_355,N_2954,N_2967);
or UO_356 (O_356,N_2990,N_2974);
and UO_357 (O_357,N_2957,N_2976);
or UO_358 (O_358,N_2957,N_2973);
nand UO_359 (O_359,N_2990,N_2971);
and UO_360 (O_360,N_2927,N_2956);
or UO_361 (O_361,N_2994,N_2926);
and UO_362 (O_362,N_2994,N_2941);
and UO_363 (O_363,N_2968,N_2978);
xor UO_364 (O_364,N_2945,N_2970);
xnor UO_365 (O_365,N_2991,N_2942);
nand UO_366 (O_366,N_2958,N_2962);
xnor UO_367 (O_367,N_2999,N_2972);
nand UO_368 (O_368,N_2925,N_2929);
nor UO_369 (O_369,N_2974,N_2932);
nor UO_370 (O_370,N_2983,N_2986);
or UO_371 (O_371,N_2990,N_2985);
nor UO_372 (O_372,N_2936,N_2939);
nand UO_373 (O_373,N_2947,N_2994);
nor UO_374 (O_374,N_2987,N_2929);
or UO_375 (O_375,N_2985,N_2968);
xor UO_376 (O_376,N_2957,N_2927);
and UO_377 (O_377,N_2962,N_2929);
xnor UO_378 (O_378,N_2984,N_2979);
and UO_379 (O_379,N_2994,N_2982);
or UO_380 (O_380,N_2963,N_2974);
or UO_381 (O_381,N_2971,N_2933);
or UO_382 (O_382,N_2928,N_2986);
xnor UO_383 (O_383,N_2951,N_2939);
or UO_384 (O_384,N_2967,N_2979);
and UO_385 (O_385,N_2997,N_2979);
nand UO_386 (O_386,N_2970,N_2934);
xnor UO_387 (O_387,N_2998,N_2936);
or UO_388 (O_388,N_2993,N_2984);
and UO_389 (O_389,N_2993,N_2953);
nor UO_390 (O_390,N_2941,N_2999);
nor UO_391 (O_391,N_2993,N_2964);
and UO_392 (O_392,N_2927,N_2986);
nand UO_393 (O_393,N_2959,N_2987);
xnor UO_394 (O_394,N_2962,N_2989);
or UO_395 (O_395,N_2964,N_2954);
and UO_396 (O_396,N_2961,N_2953);
nand UO_397 (O_397,N_2951,N_2927);
or UO_398 (O_398,N_2979,N_2957);
nor UO_399 (O_399,N_2967,N_2975);
nand UO_400 (O_400,N_2987,N_2974);
nand UO_401 (O_401,N_2958,N_2953);
and UO_402 (O_402,N_2946,N_2950);
nor UO_403 (O_403,N_2933,N_2937);
and UO_404 (O_404,N_2962,N_2983);
xnor UO_405 (O_405,N_2965,N_2972);
xnor UO_406 (O_406,N_2967,N_2936);
nand UO_407 (O_407,N_2994,N_2951);
and UO_408 (O_408,N_2970,N_2986);
nand UO_409 (O_409,N_2986,N_2998);
and UO_410 (O_410,N_2986,N_2954);
xor UO_411 (O_411,N_2943,N_2990);
and UO_412 (O_412,N_2953,N_2944);
and UO_413 (O_413,N_2934,N_2977);
nand UO_414 (O_414,N_2945,N_2944);
nor UO_415 (O_415,N_2999,N_2976);
and UO_416 (O_416,N_2988,N_2986);
nand UO_417 (O_417,N_2949,N_2968);
nand UO_418 (O_418,N_2982,N_2973);
and UO_419 (O_419,N_2953,N_2978);
and UO_420 (O_420,N_2925,N_2965);
or UO_421 (O_421,N_2927,N_2985);
and UO_422 (O_422,N_2956,N_2979);
nor UO_423 (O_423,N_2955,N_2957);
and UO_424 (O_424,N_2995,N_2983);
and UO_425 (O_425,N_2957,N_2956);
nand UO_426 (O_426,N_2943,N_2982);
or UO_427 (O_427,N_2992,N_2997);
or UO_428 (O_428,N_2943,N_2927);
nand UO_429 (O_429,N_2945,N_2968);
and UO_430 (O_430,N_2946,N_2949);
xnor UO_431 (O_431,N_2956,N_2982);
nor UO_432 (O_432,N_2978,N_2935);
nor UO_433 (O_433,N_2964,N_2953);
or UO_434 (O_434,N_2966,N_2939);
or UO_435 (O_435,N_2983,N_2993);
nand UO_436 (O_436,N_2982,N_2937);
and UO_437 (O_437,N_2957,N_2972);
xnor UO_438 (O_438,N_2945,N_2980);
nand UO_439 (O_439,N_2983,N_2969);
nor UO_440 (O_440,N_2962,N_2991);
and UO_441 (O_441,N_2950,N_2957);
and UO_442 (O_442,N_2994,N_2990);
and UO_443 (O_443,N_2977,N_2953);
or UO_444 (O_444,N_2979,N_2995);
and UO_445 (O_445,N_2999,N_2944);
nand UO_446 (O_446,N_2957,N_2925);
nand UO_447 (O_447,N_2950,N_2997);
and UO_448 (O_448,N_2990,N_2998);
or UO_449 (O_449,N_2953,N_2998);
and UO_450 (O_450,N_2947,N_2966);
and UO_451 (O_451,N_2985,N_2959);
xnor UO_452 (O_452,N_2972,N_2996);
nor UO_453 (O_453,N_2955,N_2976);
or UO_454 (O_454,N_2998,N_2970);
or UO_455 (O_455,N_2995,N_2930);
and UO_456 (O_456,N_2985,N_2956);
nand UO_457 (O_457,N_2937,N_2929);
xnor UO_458 (O_458,N_2946,N_2971);
or UO_459 (O_459,N_2940,N_2932);
or UO_460 (O_460,N_2965,N_2959);
nand UO_461 (O_461,N_2944,N_2951);
and UO_462 (O_462,N_2951,N_2945);
nor UO_463 (O_463,N_2964,N_2983);
or UO_464 (O_464,N_2956,N_2984);
nor UO_465 (O_465,N_2991,N_2965);
or UO_466 (O_466,N_2990,N_2948);
and UO_467 (O_467,N_2969,N_2946);
or UO_468 (O_468,N_2979,N_2973);
and UO_469 (O_469,N_2940,N_2929);
or UO_470 (O_470,N_2931,N_2980);
or UO_471 (O_471,N_2941,N_2960);
nand UO_472 (O_472,N_2996,N_2964);
xor UO_473 (O_473,N_2960,N_2938);
or UO_474 (O_474,N_2948,N_2960);
nor UO_475 (O_475,N_2961,N_2943);
and UO_476 (O_476,N_2994,N_2991);
nor UO_477 (O_477,N_2942,N_2933);
and UO_478 (O_478,N_2931,N_2972);
or UO_479 (O_479,N_2928,N_2944);
and UO_480 (O_480,N_2964,N_2942);
and UO_481 (O_481,N_2983,N_2951);
xor UO_482 (O_482,N_2944,N_2986);
and UO_483 (O_483,N_2992,N_2990);
nand UO_484 (O_484,N_2977,N_2978);
and UO_485 (O_485,N_2982,N_2979);
nand UO_486 (O_486,N_2940,N_2987);
nor UO_487 (O_487,N_2925,N_2940);
nor UO_488 (O_488,N_2987,N_2928);
and UO_489 (O_489,N_2971,N_2986);
nor UO_490 (O_490,N_2947,N_2983);
and UO_491 (O_491,N_2989,N_2950);
and UO_492 (O_492,N_2935,N_2979);
nand UO_493 (O_493,N_2936,N_2971);
nor UO_494 (O_494,N_2954,N_2989);
nor UO_495 (O_495,N_2965,N_2936);
and UO_496 (O_496,N_2941,N_2977);
xor UO_497 (O_497,N_2979,N_2974);
or UO_498 (O_498,N_2960,N_2925);
or UO_499 (O_499,N_2984,N_2925);
endmodule