module basic_750_5000_1000_5_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_314,In_561);
nor U1 (N_1,In_742,In_463);
or U2 (N_2,In_665,In_533);
and U3 (N_3,In_103,In_380);
nor U4 (N_4,In_303,In_136);
or U5 (N_5,In_372,In_143);
nand U6 (N_6,In_526,In_87);
nor U7 (N_7,In_546,In_114);
or U8 (N_8,In_277,In_569);
and U9 (N_9,In_185,In_284);
nor U10 (N_10,In_333,In_106);
nor U11 (N_11,In_265,In_699);
xor U12 (N_12,In_565,In_743);
xnor U13 (N_13,In_370,In_134);
and U14 (N_14,In_127,In_153);
nor U15 (N_15,In_667,In_334);
nand U16 (N_16,In_191,In_724);
xor U17 (N_17,In_392,In_749);
and U18 (N_18,In_394,In_340);
xor U19 (N_19,In_27,In_4);
or U20 (N_20,In_92,In_607);
or U21 (N_21,In_734,In_249);
nor U22 (N_22,In_43,In_503);
xor U23 (N_23,In_579,In_436);
or U24 (N_24,In_157,In_105);
or U25 (N_25,In_696,In_327);
nor U26 (N_26,In_304,In_337);
and U27 (N_27,In_728,In_470);
nor U28 (N_28,In_266,In_414);
and U29 (N_29,In_345,In_140);
or U30 (N_30,In_94,In_735);
or U31 (N_31,In_8,In_244);
nor U32 (N_32,In_443,In_286);
xor U33 (N_33,In_212,In_60);
and U34 (N_34,In_705,In_586);
and U35 (N_35,In_637,In_694);
or U36 (N_36,In_176,In_13);
nor U37 (N_37,In_226,In_72);
xor U38 (N_38,In_150,In_505);
or U39 (N_39,In_604,In_90);
nand U40 (N_40,In_440,In_307);
and U41 (N_41,In_231,In_241);
and U42 (N_42,In_74,In_164);
and U43 (N_43,In_585,In_373);
or U44 (N_44,In_525,In_224);
nor U45 (N_45,In_182,In_410);
xnor U46 (N_46,In_454,In_678);
or U47 (N_47,In_99,In_687);
nand U48 (N_48,In_568,In_530);
and U49 (N_49,In_52,In_395);
nand U50 (N_50,In_118,In_207);
or U51 (N_51,In_278,In_268);
xor U52 (N_52,In_700,In_196);
nor U53 (N_53,In_315,In_670);
nand U54 (N_54,In_747,In_712);
or U55 (N_55,In_643,In_89);
xnor U56 (N_56,In_706,In_381);
xor U57 (N_57,In_56,In_205);
nor U58 (N_58,In_177,In_431);
nand U59 (N_59,In_623,In_635);
nor U60 (N_60,In_343,In_350);
nor U61 (N_61,In_233,In_326);
xor U62 (N_62,In_459,In_632);
and U63 (N_63,In_650,In_547);
nor U64 (N_64,In_296,In_225);
and U65 (N_65,In_281,In_512);
nor U66 (N_66,In_285,In_276);
xnor U67 (N_67,In_722,In_3);
nor U68 (N_68,In_252,In_647);
and U69 (N_69,In_692,In_393);
and U70 (N_70,In_214,In_336);
xor U71 (N_71,In_596,In_360);
nor U72 (N_72,In_36,In_29);
nand U73 (N_73,In_654,In_536);
or U74 (N_74,In_234,In_527);
nand U75 (N_75,In_96,In_709);
nand U76 (N_76,In_169,In_313);
nand U77 (N_77,In_550,In_270);
nand U78 (N_78,In_489,In_368);
and U79 (N_79,In_476,In_497);
nand U80 (N_80,In_7,In_203);
and U81 (N_81,In_494,In_739);
or U82 (N_82,In_475,In_479);
xor U83 (N_83,In_59,In_119);
or U84 (N_84,In_61,In_523);
xor U85 (N_85,In_197,In_58);
nor U86 (N_86,In_675,In_112);
xnor U87 (N_87,In_450,In_642);
xnor U88 (N_88,In_673,In_445);
nor U89 (N_89,In_657,In_655);
nand U90 (N_90,In_40,In_358);
nor U91 (N_91,In_236,In_206);
nor U92 (N_92,In_415,In_543);
and U93 (N_93,In_35,In_291);
nand U94 (N_94,In_218,In_256);
nand U95 (N_95,In_733,In_575);
nor U96 (N_96,In_9,In_247);
or U97 (N_97,In_329,In_80);
or U98 (N_98,In_748,In_455);
xnor U99 (N_99,In_316,In_560);
or U100 (N_100,In_110,In_534);
nor U101 (N_101,In_298,In_466);
nor U102 (N_102,In_482,In_698);
or U103 (N_103,In_625,In_230);
nand U104 (N_104,In_194,In_605);
nand U105 (N_105,In_332,In_460);
or U106 (N_106,In_498,In_366);
xor U107 (N_107,In_640,In_383);
nand U108 (N_108,In_702,In_406);
nor U109 (N_109,In_155,In_583);
nor U110 (N_110,In_135,In_578);
nand U111 (N_111,In_402,In_184);
and U112 (N_112,In_597,In_146);
or U113 (N_113,In_438,In_81);
nand U114 (N_114,In_587,In_15);
xor U115 (N_115,In_279,In_591);
xor U116 (N_116,In_188,In_297);
nand U117 (N_117,In_319,In_282);
or U118 (N_118,In_172,In_636);
nor U119 (N_119,In_129,In_506);
nand U120 (N_120,In_631,In_317);
and U121 (N_121,In_500,In_502);
and U122 (N_122,In_581,In_420);
or U123 (N_123,In_183,In_166);
xnor U124 (N_124,In_697,In_412);
and U125 (N_125,In_684,In_311);
nand U126 (N_126,In_38,In_111);
and U127 (N_127,In_202,In_49);
nor U128 (N_128,In_362,In_131);
nor U129 (N_129,In_156,In_309);
xor U130 (N_130,In_483,In_389);
and U131 (N_131,In_490,In_144);
and U132 (N_132,In_645,In_659);
or U133 (N_133,In_613,In_25);
xnor U134 (N_134,In_713,In_626);
nand U135 (N_135,In_727,In_537);
xor U136 (N_136,In_151,In_710);
xor U137 (N_137,In_610,In_357);
or U138 (N_138,In_528,In_539);
xnor U139 (N_139,In_181,In_18);
nand U140 (N_140,In_718,In_294);
nor U141 (N_141,In_208,In_227);
or U142 (N_142,In_142,In_573);
nand U143 (N_143,In_464,In_744);
or U144 (N_144,In_385,In_159);
nor U145 (N_145,In_299,In_620);
and U146 (N_146,In_167,In_514);
nor U147 (N_147,In_63,In_215);
xnor U148 (N_148,In_474,In_308);
nor U149 (N_149,In_520,In_64);
nor U150 (N_150,In_186,In_86);
xnor U151 (N_151,In_149,In_283);
xor U152 (N_152,In_486,In_574);
or U153 (N_153,In_369,In_648);
or U154 (N_154,In_419,In_651);
and U155 (N_155,In_467,In_342);
or U156 (N_156,In_658,In_264);
xnor U157 (N_157,In_522,In_446);
and U158 (N_158,In_639,In_617);
nor U159 (N_159,In_109,In_367);
nor U160 (N_160,In_740,In_187);
xnor U161 (N_161,In_353,In_564);
and U162 (N_162,In_418,In_97);
xnor U163 (N_163,In_469,In_243);
nor U164 (N_164,In_571,In_535);
nor U165 (N_165,In_201,In_34);
and U166 (N_166,In_671,In_708);
nor U167 (N_167,In_551,In_220);
and U168 (N_168,In_508,In_375);
and U169 (N_169,In_171,In_179);
nand U170 (N_170,In_354,In_683);
or U171 (N_171,In_1,In_161);
or U172 (N_172,In_745,In_677);
nor U173 (N_173,In_458,In_524);
nand U174 (N_174,In_462,In_257);
xnor U175 (N_175,In_359,In_158);
xor U176 (N_176,In_473,In_273);
and U177 (N_177,In_595,In_554);
or U178 (N_178,In_618,In_387);
or U179 (N_179,In_53,In_444);
and U180 (N_180,In_646,In_468);
nand U181 (N_181,In_2,In_556);
nor U182 (N_182,In_344,In_19);
xor U183 (N_183,In_199,In_269);
or U184 (N_184,In_104,In_17);
or U185 (N_185,In_292,In_472);
or U186 (N_186,In_725,In_261);
nand U187 (N_187,In_666,In_178);
nand U188 (N_188,In_662,In_634);
xor U189 (N_189,In_251,In_132);
nor U190 (N_190,In_555,In_192);
or U191 (N_191,In_71,In_588);
and U192 (N_192,In_240,In_679);
nor U193 (N_193,In_130,In_390);
or U194 (N_194,In_141,In_685);
or U195 (N_195,In_211,In_552);
or U196 (N_196,In_20,In_47);
nor U197 (N_197,In_511,In_624);
nand U198 (N_198,In_95,In_532);
and U199 (N_199,In_544,In_424);
nor U200 (N_200,In_545,In_125);
nand U201 (N_201,In_324,In_300);
nor U202 (N_202,In_113,In_165);
and U203 (N_203,In_352,In_638);
or U204 (N_204,In_39,In_229);
nor U205 (N_205,In_374,In_235);
xor U206 (N_206,In_190,In_57);
xor U207 (N_207,In_173,In_77);
or U208 (N_208,In_69,In_693);
nor U209 (N_209,In_616,In_719);
nand U210 (N_210,In_433,In_541);
nand U211 (N_211,In_396,In_656);
xor U212 (N_212,In_409,In_14);
or U213 (N_213,In_200,In_477);
and U214 (N_214,In_355,In_653);
nand U215 (N_215,In_107,In_121);
and U216 (N_216,In_364,In_253);
nand U217 (N_217,In_495,In_398);
nor U218 (N_218,In_301,In_453);
and U219 (N_219,In_622,In_447);
or U220 (N_220,In_519,In_714);
and U221 (N_221,In_515,In_239);
or U222 (N_222,In_471,In_397);
and U223 (N_223,In_538,In_377);
nand U224 (N_224,In_633,In_37);
nor U225 (N_225,In_717,In_137);
and U226 (N_226,In_295,In_703);
xor U227 (N_227,In_488,In_701);
xor U228 (N_228,In_189,In_576);
nor U229 (N_229,In_430,In_160);
or U230 (N_230,In_128,In_644);
xor U231 (N_231,In_65,In_404);
or U232 (N_232,In_451,In_46);
xor U233 (N_233,In_28,In_549);
nand U234 (N_234,In_401,In_41);
and U235 (N_235,In_271,In_5);
xor U236 (N_236,In_246,In_391);
or U237 (N_237,In_501,In_163);
nand U238 (N_238,In_24,In_288);
and U239 (N_239,In_154,In_711);
xnor U240 (N_240,In_162,In_628);
nor U241 (N_241,In_738,In_82);
and U242 (N_242,In_630,In_351);
nor U243 (N_243,In_91,In_382);
xor U244 (N_244,In_741,In_54);
nand U245 (N_245,In_139,In_223);
nor U246 (N_246,In_310,In_553);
nand U247 (N_247,In_590,In_210);
nand U248 (N_248,In_50,In_723);
or U249 (N_249,In_598,In_649);
xnor U250 (N_250,In_384,In_682);
nand U251 (N_251,In_260,In_540);
nor U252 (N_252,In_388,In_238);
nor U253 (N_253,In_250,In_518);
or U254 (N_254,In_102,In_108);
and U255 (N_255,In_79,In_306);
and U256 (N_256,In_558,In_611);
or U257 (N_257,In_70,In_66);
or U258 (N_258,In_413,In_690);
nand U259 (N_259,In_660,In_716);
xor U260 (N_260,In_510,In_441);
nor U261 (N_261,In_221,In_98);
and U262 (N_262,In_562,In_122);
nand U263 (N_263,In_715,In_688);
and U264 (N_264,In_290,In_361);
nand U265 (N_265,In_442,In_195);
nor U266 (N_266,In_330,In_485);
or U267 (N_267,In_487,In_606);
and U268 (N_268,In_517,In_504);
nand U269 (N_269,In_493,In_216);
and U270 (N_270,In_593,In_531);
xnor U271 (N_271,In_434,In_602);
xnor U272 (N_272,In_492,In_346);
and U273 (N_273,In_435,In_85);
nor U274 (N_274,In_707,In_465);
and U275 (N_275,In_736,In_376);
and U276 (N_276,In_117,In_423);
xnor U277 (N_277,In_147,In_305);
nand U278 (N_278,In_612,In_730);
xnor U279 (N_279,In_426,In_21);
xor U280 (N_280,In_228,In_509);
nor U281 (N_281,In_363,In_180);
nor U282 (N_282,In_542,In_417);
or U283 (N_283,In_582,In_674);
and U284 (N_284,In_681,In_323);
xnor U285 (N_285,In_600,In_204);
nor U286 (N_286,In_746,In_428);
or U287 (N_287,In_403,In_16);
and U288 (N_288,In_341,In_322);
nand U289 (N_289,In_209,In_672);
or U290 (N_290,In_62,In_6);
xnor U291 (N_291,In_348,In_601);
nor U292 (N_292,In_100,In_347);
xnor U293 (N_293,In_680,In_289);
and U294 (N_294,In_83,In_513);
and U295 (N_295,In_45,In_386);
nand U296 (N_296,In_263,In_664);
nor U297 (N_297,In_302,In_272);
or U298 (N_298,In_33,In_621);
or U299 (N_299,In_349,In_557);
xor U300 (N_300,In_242,In_55);
or U301 (N_301,In_76,In_175);
xnor U302 (N_302,In_484,In_720);
or U303 (N_303,In_321,In_356);
nand U304 (N_304,In_429,In_481);
nand U305 (N_305,In_267,In_48);
nand U306 (N_306,In_44,In_439);
nor U307 (N_307,In_101,In_255);
xnor U308 (N_308,In_115,In_668);
nor U309 (N_309,In_721,In_732);
or U310 (N_310,In_254,In_609);
and U311 (N_311,In_152,In_193);
nor U312 (N_312,In_30,In_331);
and U313 (N_313,In_10,In_23);
xnor U314 (N_314,In_174,In_259);
xnor U315 (N_315,In_478,In_335);
xnor U316 (N_316,In_262,In_275);
xnor U317 (N_317,In_168,In_400);
and U318 (N_318,In_365,In_449);
nor U319 (N_319,In_287,In_695);
or U320 (N_320,In_42,In_516);
or U321 (N_321,In_661,In_222);
xor U322 (N_322,In_437,In_75);
or U323 (N_323,In_427,In_22);
and U324 (N_324,In_32,In_480);
or U325 (N_325,In_258,In_126);
xor U326 (N_326,In_123,In_457);
and U327 (N_327,In_170,In_217);
nand U328 (N_328,In_245,In_198);
xor U329 (N_329,In_641,In_456);
nand U330 (N_330,In_78,In_88);
and U331 (N_331,In_448,In_563);
nand U332 (N_332,In_84,In_577);
nand U333 (N_333,In_31,In_599);
nand U334 (N_334,In_237,In_669);
nand U335 (N_335,In_379,In_726);
xnor U336 (N_336,In_138,In_603);
nand U337 (N_337,In_452,In_691);
or U338 (N_338,In_507,In_594);
or U339 (N_339,In_320,In_312);
xnor U340 (N_340,In_422,In_248);
nor U341 (N_341,In_405,In_572);
nor U342 (N_342,In_592,In_145);
or U343 (N_343,In_68,In_608);
and U344 (N_344,In_213,In_339);
nor U345 (N_345,In_499,In_116);
and U346 (N_346,In_73,In_521);
xnor U347 (N_347,In_432,In_425);
nor U348 (N_348,In_580,In_619);
nor U349 (N_349,In_51,In_663);
nor U350 (N_350,In_731,In_614);
nor U351 (N_351,In_318,In_737);
nand U352 (N_352,In_11,In_559);
and U353 (N_353,In_399,In_421);
nand U354 (N_354,In_529,In_496);
or U355 (N_355,In_567,In_93);
xnor U356 (N_356,In_408,In_548);
xnor U357 (N_357,In_12,In_491);
nand U358 (N_358,In_676,In_371);
xnor U359 (N_359,In_378,In_274);
or U360 (N_360,In_629,In_148);
nand U361 (N_361,In_26,In_461);
or U362 (N_362,In_338,In_120);
and U363 (N_363,In_729,In_584);
or U364 (N_364,In_0,In_133);
nor U365 (N_365,In_686,In_67);
nor U366 (N_366,In_570,In_293);
nor U367 (N_367,In_411,In_566);
or U368 (N_368,In_219,In_416);
or U369 (N_369,In_704,In_280);
nand U370 (N_370,In_328,In_689);
xnor U371 (N_371,In_589,In_407);
nor U372 (N_372,In_627,In_232);
nor U373 (N_373,In_615,In_652);
xor U374 (N_374,In_124,In_325);
xor U375 (N_375,In_131,In_301);
and U376 (N_376,In_200,In_182);
and U377 (N_377,In_387,In_9);
nand U378 (N_378,In_107,In_504);
and U379 (N_379,In_347,In_127);
nand U380 (N_380,In_605,In_224);
or U381 (N_381,In_190,In_556);
xor U382 (N_382,In_83,In_406);
xor U383 (N_383,In_745,In_587);
nand U384 (N_384,In_269,In_44);
nand U385 (N_385,In_537,In_621);
xnor U386 (N_386,In_725,In_309);
and U387 (N_387,In_6,In_628);
nor U388 (N_388,In_293,In_729);
nor U389 (N_389,In_450,In_494);
xor U390 (N_390,In_479,In_178);
and U391 (N_391,In_8,In_509);
xor U392 (N_392,In_477,In_241);
xnor U393 (N_393,In_154,In_224);
or U394 (N_394,In_704,In_442);
nand U395 (N_395,In_362,In_574);
xor U396 (N_396,In_495,In_163);
or U397 (N_397,In_363,In_60);
nand U398 (N_398,In_590,In_250);
nor U399 (N_399,In_684,In_421);
nor U400 (N_400,In_108,In_31);
or U401 (N_401,In_67,In_312);
and U402 (N_402,In_84,In_590);
xnor U403 (N_403,In_43,In_323);
and U404 (N_404,In_548,In_27);
nor U405 (N_405,In_54,In_406);
xnor U406 (N_406,In_512,In_655);
nor U407 (N_407,In_430,In_150);
nor U408 (N_408,In_556,In_181);
xnor U409 (N_409,In_619,In_482);
nor U410 (N_410,In_393,In_154);
xnor U411 (N_411,In_336,In_408);
xor U412 (N_412,In_132,In_268);
or U413 (N_413,In_180,In_564);
nand U414 (N_414,In_61,In_697);
or U415 (N_415,In_384,In_735);
or U416 (N_416,In_39,In_648);
xor U417 (N_417,In_322,In_585);
nand U418 (N_418,In_672,In_457);
and U419 (N_419,In_497,In_477);
xnor U420 (N_420,In_576,In_373);
nor U421 (N_421,In_414,In_31);
nand U422 (N_422,In_141,In_536);
or U423 (N_423,In_519,In_326);
and U424 (N_424,In_123,In_67);
or U425 (N_425,In_717,In_393);
or U426 (N_426,In_323,In_115);
and U427 (N_427,In_224,In_11);
nor U428 (N_428,In_252,In_490);
nor U429 (N_429,In_352,In_119);
nor U430 (N_430,In_237,In_605);
or U431 (N_431,In_579,In_196);
xnor U432 (N_432,In_721,In_230);
xnor U433 (N_433,In_670,In_46);
and U434 (N_434,In_440,In_436);
nand U435 (N_435,In_147,In_650);
xnor U436 (N_436,In_139,In_126);
and U437 (N_437,In_672,In_379);
and U438 (N_438,In_538,In_732);
xnor U439 (N_439,In_161,In_190);
xnor U440 (N_440,In_9,In_374);
and U441 (N_441,In_153,In_372);
xnor U442 (N_442,In_695,In_586);
nor U443 (N_443,In_67,In_23);
nand U444 (N_444,In_671,In_365);
xor U445 (N_445,In_533,In_364);
xnor U446 (N_446,In_35,In_231);
nand U447 (N_447,In_478,In_253);
nor U448 (N_448,In_14,In_514);
xor U449 (N_449,In_115,In_81);
nand U450 (N_450,In_611,In_226);
nor U451 (N_451,In_419,In_254);
xor U452 (N_452,In_430,In_193);
and U453 (N_453,In_213,In_593);
nand U454 (N_454,In_74,In_154);
and U455 (N_455,In_697,In_420);
nand U456 (N_456,In_357,In_343);
nand U457 (N_457,In_12,In_289);
xnor U458 (N_458,In_490,In_42);
and U459 (N_459,In_398,In_4);
nand U460 (N_460,In_426,In_69);
nand U461 (N_461,In_286,In_41);
xor U462 (N_462,In_68,In_682);
nand U463 (N_463,In_158,In_673);
xnor U464 (N_464,In_187,In_252);
and U465 (N_465,In_252,In_662);
and U466 (N_466,In_303,In_682);
nand U467 (N_467,In_471,In_254);
or U468 (N_468,In_392,In_659);
nor U469 (N_469,In_77,In_13);
and U470 (N_470,In_123,In_196);
xor U471 (N_471,In_702,In_678);
nor U472 (N_472,In_402,In_152);
nand U473 (N_473,In_71,In_256);
nor U474 (N_474,In_594,In_601);
nor U475 (N_475,In_130,In_179);
nor U476 (N_476,In_451,In_65);
or U477 (N_477,In_549,In_713);
nor U478 (N_478,In_648,In_663);
nand U479 (N_479,In_175,In_571);
or U480 (N_480,In_162,In_308);
and U481 (N_481,In_443,In_617);
xnor U482 (N_482,In_568,In_224);
nor U483 (N_483,In_446,In_675);
or U484 (N_484,In_481,In_492);
xor U485 (N_485,In_213,In_518);
and U486 (N_486,In_351,In_566);
and U487 (N_487,In_185,In_549);
nand U488 (N_488,In_331,In_691);
and U489 (N_489,In_595,In_489);
nand U490 (N_490,In_711,In_352);
nor U491 (N_491,In_690,In_261);
or U492 (N_492,In_595,In_342);
nor U493 (N_493,In_514,In_3);
and U494 (N_494,In_7,In_297);
or U495 (N_495,In_549,In_25);
nand U496 (N_496,In_92,In_22);
xnor U497 (N_497,In_94,In_318);
or U498 (N_498,In_368,In_444);
xor U499 (N_499,In_254,In_162);
and U500 (N_500,In_154,In_115);
xor U501 (N_501,In_546,In_723);
nor U502 (N_502,In_618,In_344);
nor U503 (N_503,In_728,In_386);
nand U504 (N_504,In_180,In_549);
and U505 (N_505,In_341,In_238);
nor U506 (N_506,In_157,In_257);
nor U507 (N_507,In_374,In_97);
and U508 (N_508,In_521,In_663);
xor U509 (N_509,In_494,In_435);
or U510 (N_510,In_176,In_235);
nand U511 (N_511,In_26,In_170);
nand U512 (N_512,In_698,In_744);
xnor U513 (N_513,In_714,In_627);
xnor U514 (N_514,In_321,In_404);
nor U515 (N_515,In_152,In_468);
xor U516 (N_516,In_24,In_258);
or U517 (N_517,In_457,In_508);
nand U518 (N_518,In_595,In_441);
or U519 (N_519,In_426,In_7);
nand U520 (N_520,In_523,In_247);
xor U521 (N_521,In_224,In_433);
xnor U522 (N_522,In_132,In_9);
nand U523 (N_523,In_206,In_305);
xor U524 (N_524,In_359,In_165);
nand U525 (N_525,In_744,In_524);
or U526 (N_526,In_667,In_618);
xnor U527 (N_527,In_596,In_443);
xnor U528 (N_528,In_345,In_276);
or U529 (N_529,In_281,In_735);
or U530 (N_530,In_746,In_103);
xor U531 (N_531,In_389,In_3);
nand U532 (N_532,In_610,In_103);
and U533 (N_533,In_744,In_293);
nor U534 (N_534,In_231,In_196);
and U535 (N_535,In_727,In_578);
nor U536 (N_536,In_653,In_628);
nand U537 (N_537,In_111,In_22);
and U538 (N_538,In_356,In_384);
and U539 (N_539,In_229,In_321);
and U540 (N_540,In_154,In_305);
and U541 (N_541,In_69,In_647);
and U542 (N_542,In_26,In_382);
nor U543 (N_543,In_565,In_338);
nor U544 (N_544,In_77,In_593);
nor U545 (N_545,In_592,In_181);
or U546 (N_546,In_717,In_734);
xor U547 (N_547,In_681,In_108);
or U548 (N_548,In_662,In_251);
nor U549 (N_549,In_265,In_48);
and U550 (N_550,In_151,In_430);
xor U551 (N_551,In_329,In_436);
xnor U552 (N_552,In_79,In_562);
and U553 (N_553,In_641,In_110);
or U554 (N_554,In_442,In_517);
nand U555 (N_555,In_628,In_357);
nor U556 (N_556,In_741,In_695);
or U557 (N_557,In_738,In_54);
nor U558 (N_558,In_417,In_585);
nor U559 (N_559,In_274,In_355);
xor U560 (N_560,In_265,In_324);
nand U561 (N_561,In_1,In_685);
or U562 (N_562,In_95,In_411);
nand U563 (N_563,In_702,In_258);
and U564 (N_564,In_360,In_113);
xor U565 (N_565,In_654,In_423);
nor U566 (N_566,In_231,In_361);
xnor U567 (N_567,In_579,In_477);
and U568 (N_568,In_478,In_115);
or U569 (N_569,In_505,In_377);
xor U570 (N_570,In_612,In_697);
nand U571 (N_571,In_743,In_379);
nor U572 (N_572,In_251,In_468);
nand U573 (N_573,In_332,In_49);
xor U574 (N_574,In_452,In_743);
xor U575 (N_575,In_395,In_35);
or U576 (N_576,In_634,In_297);
nand U577 (N_577,In_442,In_191);
or U578 (N_578,In_665,In_35);
or U579 (N_579,In_436,In_141);
xnor U580 (N_580,In_636,In_200);
nand U581 (N_581,In_309,In_666);
nor U582 (N_582,In_407,In_177);
xor U583 (N_583,In_155,In_356);
or U584 (N_584,In_452,In_386);
nand U585 (N_585,In_586,In_673);
and U586 (N_586,In_297,In_561);
and U587 (N_587,In_547,In_408);
nor U588 (N_588,In_638,In_139);
nor U589 (N_589,In_324,In_450);
or U590 (N_590,In_297,In_264);
and U591 (N_591,In_239,In_363);
xnor U592 (N_592,In_407,In_169);
and U593 (N_593,In_15,In_69);
and U594 (N_594,In_539,In_52);
nor U595 (N_595,In_525,In_740);
nor U596 (N_596,In_185,In_237);
or U597 (N_597,In_265,In_635);
or U598 (N_598,In_658,In_715);
nand U599 (N_599,In_221,In_330);
nand U600 (N_600,In_581,In_171);
or U601 (N_601,In_126,In_647);
xnor U602 (N_602,In_315,In_299);
and U603 (N_603,In_179,In_60);
xnor U604 (N_604,In_601,In_488);
nand U605 (N_605,In_497,In_395);
and U606 (N_606,In_444,In_694);
nor U607 (N_607,In_682,In_247);
xor U608 (N_608,In_612,In_619);
and U609 (N_609,In_721,In_270);
and U610 (N_610,In_384,In_558);
nor U611 (N_611,In_729,In_244);
and U612 (N_612,In_283,In_195);
nand U613 (N_613,In_86,In_152);
xnor U614 (N_614,In_62,In_536);
nand U615 (N_615,In_684,In_594);
nand U616 (N_616,In_114,In_93);
or U617 (N_617,In_511,In_166);
nand U618 (N_618,In_212,In_19);
xor U619 (N_619,In_390,In_354);
and U620 (N_620,In_103,In_554);
and U621 (N_621,In_173,In_466);
or U622 (N_622,In_550,In_194);
or U623 (N_623,In_40,In_303);
nor U624 (N_624,In_480,In_412);
or U625 (N_625,In_94,In_486);
nor U626 (N_626,In_652,In_59);
nor U627 (N_627,In_264,In_534);
xor U628 (N_628,In_673,In_606);
nor U629 (N_629,In_427,In_566);
xor U630 (N_630,In_211,In_195);
and U631 (N_631,In_663,In_575);
xnor U632 (N_632,In_481,In_524);
or U633 (N_633,In_119,In_82);
xor U634 (N_634,In_33,In_441);
nand U635 (N_635,In_591,In_19);
nand U636 (N_636,In_254,In_524);
xor U637 (N_637,In_454,In_36);
nor U638 (N_638,In_91,In_208);
nor U639 (N_639,In_92,In_317);
or U640 (N_640,In_206,In_230);
nand U641 (N_641,In_450,In_679);
nand U642 (N_642,In_171,In_562);
nand U643 (N_643,In_464,In_127);
and U644 (N_644,In_408,In_660);
nand U645 (N_645,In_192,In_510);
or U646 (N_646,In_264,In_684);
nor U647 (N_647,In_42,In_519);
nand U648 (N_648,In_2,In_706);
and U649 (N_649,In_59,In_744);
and U650 (N_650,In_155,In_57);
or U651 (N_651,In_604,In_132);
xor U652 (N_652,In_4,In_596);
or U653 (N_653,In_169,In_653);
nand U654 (N_654,In_159,In_67);
or U655 (N_655,In_475,In_236);
or U656 (N_656,In_581,In_460);
or U657 (N_657,In_213,In_144);
or U658 (N_658,In_17,In_289);
nand U659 (N_659,In_174,In_139);
nand U660 (N_660,In_394,In_414);
and U661 (N_661,In_270,In_97);
or U662 (N_662,In_254,In_477);
nand U663 (N_663,In_516,In_609);
nand U664 (N_664,In_722,In_129);
nor U665 (N_665,In_217,In_563);
nor U666 (N_666,In_231,In_697);
nand U667 (N_667,In_683,In_285);
and U668 (N_668,In_380,In_263);
nor U669 (N_669,In_69,In_613);
nor U670 (N_670,In_417,In_494);
and U671 (N_671,In_118,In_67);
nand U672 (N_672,In_629,In_69);
nor U673 (N_673,In_152,In_503);
nand U674 (N_674,In_624,In_227);
nand U675 (N_675,In_68,In_131);
nor U676 (N_676,In_219,In_451);
and U677 (N_677,In_728,In_426);
nor U678 (N_678,In_542,In_21);
nor U679 (N_679,In_577,In_117);
nor U680 (N_680,In_663,In_606);
nor U681 (N_681,In_319,In_258);
nand U682 (N_682,In_744,In_418);
nand U683 (N_683,In_194,In_191);
nand U684 (N_684,In_146,In_612);
nor U685 (N_685,In_382,In_355);
nand U686 (N_686,In_641,In_100);
and U687 (N_687,In_241,In_303);
xnor U688 (N_688,In_535,In_179);
xnor U689 (N_689,In_155,In_386);
nor U690 (N_690,In_32,In_285);
nand U691 (N_691,In_179,In_10);
or U692 (N_692,In_615,In_518);
xor U693 (N_693,In_555,In_738);
and U694 (N_694,In_53,In_192);
or U695 (N_695,In_345,In_163);
xor U696 (N_696,In_109,In_288);
nand U697 (N_697,In_154,In_438);
nor U698 (N_698,In_312,In_378);
or U699 (N_699,In_371,In_700);
or U700 (N_700,In_260,In_168);
xnor U701 (N_701,In_196,In_731);
xor U702 (N_702,In_320,In_567);
xor U703 (N_703,In_660,In_1);
nor U704 (N_704,In_202,In_3);
nand U705 (N_705,In_462,In_164);
nand U706 (N_706,In_322,In_169);
nor U707 (N_707,In_635,In_606);
nor U708 (N_708,In_269,In_130);
or U709 (N_709,In_700,In_104);
or U710 (N_710,In_558,In_570);
nand U711 (N_711,In_663,In_483);
nor U712 (N_712,In_503,In_561);
or U713 (N_713,In_294,In_497);
nor U714 (N_714,In_536,In_454);
xor U715 (N_715,In_330,In_476);
xor U716 (N_716,In_575,In_146);
nand U717 (N_717,In_43,In_7);
and U718 (N_718,In_550,In_35);
nor U719 (N_719,In_227,In_325);
nand U720 (N_720,In_396,In_368);
nor U721 (N_721,In_308,In_383);
nor U722 (N_722,In_64,In_444);
xor U723 (N_723,In_329,In_235);
or U724 (N_724,In_135,In_261);
nor U725 (N_725,In_53,In_705);
or U726 (N_726,In_579,In_458);
and U727 (N_727,In_330,In_462);
nor U728 (N_728,In_357,In_640);
or U729 (N_729,In_239,In_155);
or U730 (N_730,In_248,In_63);
xor U731 (N_731,In_686,In_525);
and U732 (N_732,In_80,In_459);
nand U733 (N_733,In_740,In_364);
nand U734 (N_734,In_504,In_560);
or U735 (N_735,In_478,In_63);
nand U736 (N_736,In_207,In_443);
nor U737 (N_737,In_135,In_122);
or U738 (N_738,In_500,In_342);
nand U739 (N_739,In_245,In_217);
or U740 (N_740,In_400,In_677);
and U741 (N_741,In_116,In_399);
xnor U742 (N_742,In_10,In_589);
nor U743 (N_743,In_99,In_601);
xor U744 (N_744,In_179,In_45);
xnor U745 (N_745,In_108,In_373);
or U746 (N_746,In_262,In_466);
nor U747 (N_747,In_583,In_316);
xnor U748 (N_748,In_648,In_220);
xor U749 (N_749,In_437,In_514);
and U750 (N_750,In_98,In_451);
and U751 (N_751,In_282,In_515);
nor U752 (N_752,In_145,In_305);
or U753 (N_753,In_293,In_550);
nand U754 (N_754,In_652,In_74);
nor U755 (N_755,In_544,In_648);
nor U756 (N_756,In_442,In_362);
and U757 (N_757,In_542,In_190);
nor U758 (N_758,In_357,In_212);
or U759 (N_759,In_336,In_696);
nor U760 (N_760,In_576,In_453);
and U761 (N_761,In_144,In_97);
and U762 (N_762,In_33,In_706);
nand U763 (N_763,In_586,In_682);
nor U764 (N_764,In_557,In_392);
nand U765 (N_765,In_356,In_150);
nand U766 (N_766,In_290,In_642);
or U767 (N_767,In_155,In_568);
or U768 (N_768,In_730,In_335);
or U769 (N_769,In_175,In_734);
nand U770 (N_770,In_215,In_136);
nor U771 (N_771,In_661,In_415);
nand U772 (N_772,In_708,In_741);
nand U773 (N_773,In_76,In_662);
nand U774 (N_774,In_497,In_660);
nor U775 (N_775,In_447,In_20);
xnor U776 (N_776,In_665,In_29);
xnor U777 (N_777,In_677,In_373);
nand U778 (N_778,In_197,In_66);
xor U779 (N_779,In_436,In_694);
nor U780 (N_780,In_281,In_712);
and U781 (N_781,In_550,In_425);
nor U782 (N_782,In_480,In_309);
nor U783 (N_783,In_706,In_389);
nand U784 (N_784,In_90,In_722);
nand U785 (N_785,In_429,In_113);
xnor U786 (N_786,In_662,In_278);
nand U787 (N_787,In_701,In_367);
and U788 (N_788,In_145,In_714);
xor U789 (N_789,In_588,In_4);
or U790 (N_790,In_316,In_105);
nand U791 (N_791,In_515,In_214);
or U792 (N_792,In_734,In_452);
nor U793 (N_793,In_501,In_243);
or U794 (N_794,In_505,In_445);
nand U795 (N_795,In_645,In_535);
or U796 (N_796,In_258,In_356);
or U797 (N_797,In_227,In_9);
nor U798 (N_798,In_387,In_571);
or U799 (N_799,In_436,In_549);
xor U800 (N_800,In_138,In_206);
nor U801 (N_801,In_715,In_274);
and U802 (N_802,In_4,In_104);
xor U803 (N_803,In_451,In_169);
nand U804 (N_804,In_721,In_464);
xnor U805 (N_805,In_33,In_742);
and U806 (N_806,In_597,In_257);
or U807 (N_807,In_64,In_476);
nand U808 (N_808,In_148,In_48);
nor U809 (N_809,In_434,In_233);
and U810 (N_810,In_711,In_6);
nor U811 (N_811,In_13,In_21);
nor U812 (N_812,In_274,In_181);
or U813 (N_813,In_232,In_31);
and U814 (N_814,In_167,In_66);
nor U815 (N_815,In_35,In_348);
nand U816 (N_816,In_264,In_529);
xor U817 (N_817,In_564,In_411);
xnor U818 (N_818,In_563,In_520);
nor U819 (N_819,In_590,In_720);
or U820 (N_820,In_372,In_690);
xnor U821 (N_821,In_248,In_263);
and U822 (N_822,In_82,In_376);
xnor U823 (N_823,In_727,In_269);
and U824 (N_824,In_565,In_179);
or U825 (N_825,In_709,In_695);
xnor U826 (N_826,In_63,In_428);
xor U827 (N_827,In_344,In_552);
and U828 (N_828,In_708,In_174);
nor U829 (N_829,In_593,In_587);
xnor U830 (N_830,In_200,In_301);
xor U831 (N_831,In_192,In_617);
nor U832 (N_832,In_128,In_522);
nor U833 (N_833,In_304,In_163);
xnor U834 (N_834,In_343,In_503);
or U835 (N_835,In_174,In_706);
or U836 (N_836,In_725,In_83);
or U837 (N_837,In_715,In_697);
xor U838 (N_838,In_342,In_545);
xnor U839 (N_839,In_128,In_403);
xor U840 (N_840,In_265,In_612);
xnor U841 (N_841,In_101,In_712);
nor U842 (N_842,In_539,In_662);
or U843 (N_843,In_69,In_440);
nand U844 (N_844,In_344,In_367);
nand U845 (N_845,In_626,In_171);
xor U846 (N_846,In_341,In_454);
and U847 (N_847,In_110,In_523);
xnor U848 (N_848,In_275,In_719);
nor U849 (N_849,In_179,In_541);
nor U850 (N_850,In_246,In_206);
nand U851 (N_851,In_320,In_586);
xnor U852 (N_852,In_691,In_635);
nand U853 (N_853,In_281,In_114);
xor U854 (N_854,In_697,In_602);
or U855 (N_855,In_159,In_427);
xnor U856 (N_856,In_684,In_695);
xor U857 (N_857,In_314,In_518);
nor U858 (N_858,In_558,In_222);
and U859 (N_859,In_385,In_408);
xnor U860 (N_860,In_385,In_431);
or U861 (N_861,In_614,In_112);
nor U862 (N_862,In_277,In_727);
or U863 (N_863,In_654,In_292);
nand U864 (N_864,In_597,In_270);
nor U865 (N_865,In_339,In_24);
and U866 (N_866,In_368,In_480);
nor U867 (N_867,In_504,In_187);
nand U868 (N_868,In_414,In_492);
xor U869 (N_869,In_107,In_219);
xnor U870 (N_870,In_450,In_48);
xor U871 (N_871,In_117,In_480);
nor U872 (N_872,In_641,In_734);
xnor U873 (N_873,In_22,In_64);
nand U874 (N_874,In_3,In_670);
nor U875 (N_875,In_360,In_438);
or U876 (N_876,In_689,In_358);
nor U877 (N_877,In_128,In_88);
nor U878 (N_878,In_305,In_658);
and U879 (N_879,In_410,In_364);
and U880 (N_880,In_447,In_465);
xnor U881 (N_881,In_162,In_285);
xor U882 (N_882,In_504,In_674);
and U883 (N_883,In_614,In_333);
nor U884 (N_884,In_518,In_514);
and U885 (N_885,In_299,In_708);
nor U886 (N_886,In_483,In_183);
and U887 (N_887,In_183,In_278);
or U888 (N_888,In_474,In_735);
or U889 (N_889,In_46,In_254);
and U890 (N_890,In_624,In_169);
xnor U891 (N_891,In_607,In_275);
nand U892 (N_892,In_431,In_278);
nand U893 (N_893,In_550,In_377);
nor U894 (N_894,In_536,In_671);
and U895 (N_895,In_427,In_656);
nand U896 (N_896,In_373,In_460);
nand U897 (N_897,In_553,In_256);
nand U898 (N_898,In_54,In_294);
xor U899 (N_899,In_562,In_738);
or U900 (N_900,In_332,In_410);
nor U901 (N_901,In_553,In_133);
and U902 (N_902,In_92,In_499);
and U903 (N_903,In_192,In_388);
nand U904 (N_904,In_547,In_554);
nand U905 (N_905,In_120,In_593);
nor U906 (N_906,In_123,In_526);
or U907 (N_907,In_44,In_105);
nor U908 (N_908,In_108,In_606);
and U909 (N_909,In_568,In_320);
nand U910 (N_910,In_258,In_582);
nor U911 (N_911,In_534,In_214);
and U912 (N_912,In_641,In_716);
xor U913 (N_913,In_604,In_160);
and U914 (N_914,In_54,In_393);
nor U915 (N_915,In_598,In_39);
xnor U916 (N_916,In_269,In_283);
nand U917 (N_917,In_552,In_663);
or U918 (N_918,In_293,In_144);
nand U919 (N_919,In_483,In_252);
xnor U920 (N_920,In_655,In_98);
nor U921 (N_921,In_299,In_377);
and U922 (N_922,In_458,In_373);
and U923 (N_923,In_218,In_699);
or U924 (N_924,In_160,In_248);
nand U925 (N_925,In_19,In_115);
xor U926 (N_926,In_201,In_630);
or U927 (N_927,In_653,In_363);
xnor U928 (N_928,In_27,In_644);
or U929 (N_929,In_98,In_270);
nand U930 (N_930,In_402,In_274);
nor U931 (N_931,In_88,In_596);
nor U932 (N_932,In_251,In_486);
xnor U933 (N_933,In_426,In_107);
xor U934 (N_934,In_424,In_2);
or U935 (N_935,In_477,In_717);
or U936 (N_936,In_699,In_691);
nor U937 (N_937,In_103,In_422);
nand U938 (N_938,In_211,In_649);
and U939 (N_939,In_713,In_451);
xnor U940 (N_940,In_512,In_321);
nor U941 (N_941,In_166,In_100);
and U942 (N_942,In_598,In_233);
nor U943 (N_943,In_554,In_114);
xnor U944 (N_944,In_607,In_479);
xor U945 (N_945,In_377,In_362);
nand U946 (N_946,In_240,In_715);
xnor U947 (N_947,In_581,In_310);
or U948 (N_948,In_729,In_144);
or U949 (N_949,In_378,In_636);
nor U950 (N_950,In_384,In_686);
nor U951 (N_951,In_506,In_279);
and U952 (N_952,In_491,In_327);
nor U953 (N_953,In_693,In_714);
nor U954 (N_954,In_467,In_193);
xor U955 (N_955,In_390,In_618);
xor U956 (N_956,In_68,In_725);
and U957 (N_957,In_44,In_556);
nor U958 (N_958,In_92,In_329);
and U959 (N_959,In_123,In_462);
xnor U960 (N_960,In_145,In_671);
or U961 (N_961,In_208,In_738);
or U962 (N_962,In_370,In_445);
xnor U963 (N_963,In_292,In_188);
nand U964 (N_964,In_743,In_187);
or U965 (N_965,In_454,In_261);
or U966 (N_966,In_457,In_495);
xnor U967 (N_967,In_58,In_510);
xnor U968 (N_968,In_495,In_272);
nor U969 (N_969,In_633,In_296);
nor U970 (N_970,In_81,In_455);
nor U971 (N_971,In_489,In_370);
nand U972 (N_972,In_504,In_425);
xnor U973 (N_973,In_250,In_2);
nor U974 (N_974,In_623,In_487);
nor U975 (N_975,In_38,In_179);
nand U976 (N_976,In_216,In_311);
xnor U977 (N_977,In_506,In_423);
and U978 (N_978,In_188,In_692);
xor U979 (N_979,In_2,In_115);
and U980 (N_980,In_21,In_554);
and U981 (N_981,In_40,In_131);
or U982 (N_982,In_19,In_327);
nand U983 (N_983,In_394,In_284);
or U984 (N_984,In_546,In_745);
and U985 (N_985,In_377,In_144);
nor U986 (N_986,In_214,In_432);
nand U987 (N_987,In_534,In_221);
xor U988 (N_988,In_221,In_178);
xor U989 (N_989,In_444,In_19);
or U990 (N_990,In_510,In_718);
or U991 (N_991,In_681,In_407);
or U992 (N_992,In_98,In_646);
nand U993 (N_993,In_106,In_75);
and U994 (N_994,In_698,In_590);
xnor U995 (N_995,In_164,In_725);
nor U996 (N_996,In_548,In_517);
nand U997 (N_997,In_730,In_76);
or U998 (N_998,In_246,In_3);
nor U999 (N_999,In_298,In_672);
and U1000 (N_1000,N_769,N_388);
nand U1001 (N_1001,N_620,N_339);
xnor U1002 (N_1002,N_170,N_162);
xor U1003 (N_1003,N_423,N_666);
xnor U1004 (N_1004,N_457,N_483);
or U1005 (N_1005,N_587,N_466);
xnor U1006 (N_1006,N_186,N_880);
xor U1007 (N_1007,N_503,N_919);
and U1008 (N_1008,N_567,N_878);
or U1009 (N_1009,N_836,N_366);
nor U1010 (N_1010,N_692,N_204);
nor U1011 (N_1011,N_991,N_763);
xor U1012 (N_1012,N_363,N_813);
or U1013 (N_1013,N_888,N_87);
and U1014 (N_1014,N_273,N_944);
nand U1015 (N_1015,N_771,N_632);
nor U1016 (N_1016,N_461,N_234);
or U1017 (N_1017,N_743,N_459);
xnor U1018 (N_1018,N_84,N_702);
or U1019 (N_1019,N_392,N_464);
and U1020 (N_1020,N_798,N_19);
nor U1021 (N_1021,N_724,N_241);
and U1022 (N_1022,N_785,N_201);
nand U1023 (N_1023,N_165,N_476);
or U1024 (N_1024,N_866,N_868);
or U1025 (N_1025,N_473,N_191);
nand U1026 (N_1026,N_312,N_727);
nor U1027 (N_1027,N_558,N_905);
nand U1028 (N_1028,N_540,N_542);
or U1029 (N_1029,N_906,N_681);
nand U1030 (N_1030,N_313,N_50);
nor U1031 (N_1031,N_62,N_573);
and U1032 (N_1032,N_135,N_437);
nor U1033 (N_1033,N_380,N_74);
xnor U1034 (N_1034,N_990,N_235);
or U1035 (N_1035,N_5,N_83);
nand U1036 (N_1036,N_401,N_912);
nor U1037 (N_1037,N_284,N_54);
and U1038 (N_1038,N_570,N_285);
and U1039 (N_1039,N_141,N_148);
and U1040 (N_1040,N_161,N_139);
nor U1041 (N_1041,N_99,N_978);
or U1042 (N_1042,N_296,N_143);
xnor U1043 (N_1043,N_242,N_908);
or U1044 (N_1044,N_815,N_864);
xor U1045 (N_1045,N_755,N_623);
nand U1046 (N_1046,N_968,N_300);
xnor U1047 (N_1047,N_480,N_914);
xor U1048 (N_1048,N_26,N_262);
nand U1049 (N_1049,N_215,N_647);
or U1050 (N_1050,N_520,N_48);
and U1051 (N_1051,N_848,N_71);
or U1052 (N_1052,N_106,N_895);
nand U1053 (N_1053,N_90,N_598);
or U1054 (N_1054,N_206,N_89);
or U1055 (N_1055,N_147,N_605);
nor U1056 (N_1056,N_629,N_420);
and U1057 (N_1057,N_155,N_863);
xor U1058 (N_1058,N_935,N_431);
xnor U1059 (N_1059,N_472,N_178);
nand U1060 (N_1060,N_543,N_131);
or U1061 (N_1061,N_784,N_993);
nand U1062 (N_1062,N_512,N_827);
xnor U1063 (N_1063,N_208,N_387);
or U1064 (N_1064,N_280,N_331);
nand U1065 (N_1065,N_283,N_153);
and U1066 (N_1066,N_744,N_151);
xnor U1067 (N_1067,N_706,N_341);
nand U1068 (N_1068,N_6,N_602);
xor U1069 (N_1069,N_484,N_889);
nand U1070 (N_1070,N_219,N_997);
nor U1071 (N_1071,N_574,N_482);
nand U1072 (N_1072,N_586,N_557);
or U1073 (N_1073,N_876,N_212);
nand U1074 (N_1074,N_651,N_531);
nor U1075 (N_1075,N_528,N_500);
nor U1076 (N_1076,N_224,N_918);
and U1077 (N_1077,N_290,N_677);
nor U1078 (N_1078,N_199,N_60);
nor U1079 (N_1079,N_794,N_317);
nor U1080 (N_1080,N_514,N_103);
nand U1081 (N_1081,N_266,N_843);
and U1082 (N_1082,N_240,N_228);
nand U1083 (N_1083,N_220,N_109);
or U1084 (N_1084,N_672,N_221);
nor U1085 (N_1085,N_776,N_370);
and U1086 (N_1086,N_497,N_728);
nand U1087 (N_1087,N_805,N_988);
nor U1088 (N_1088,N_149,N_941);
nand U1089 (N_1089,N_320,N_675);
and U1090 (N_1090,N_205,N_845);
or U1091 (N_1091,N_806,N_683);
nand U1092 (N_1092,N_882,N_577);
nor U1093 (N_1093,N_898,N_433);
nand U1094 (N_1094,N_717,N_377);
or U1095 (N_1095,N_166,N_674);
and U1096 (N_1096,N_569,N_307);
nand U1097 (N_1097,N_347,N_597);
and U1098 (N_1098,N_957,N_646);
and U1099 (N_1099,N_571,N_269);
xnor U1100 (N_1100,N_64,N_849);
or U1101 (N_1101,N_892,N_731);
or U1102 (N_1102,N_323,N_438);
or U1103 (N_1103,N_841,N_216);
xor U1104 (N_1104,N_682,N_819);
xor U1105 (N_1105,N_72,N_174);
xor U1106 (N_1106,N_625,N_777);
or U1107 (N_1107,N_455,N_17);
nor U1108 (N_1108,N_182,N_98);
and U1109 (N_1109,N_578,N_126);
xnor U1110 (N_1110,N_720,N_939);
or U1111 (N_1111,N_385,N_874);
and U1112 (N_1112,N_328,N_984);
nor U1113 (N_1113,N_18,N_448);
or U1114 (N_1114,N_555,N_343);
nor U1115 (N_1115,N_523,N_788);
and U1116 (N_1116,N_900,N_817);
nor U1117 (N_1117,N_1,N_705);
nor U1118 (N_1118,N_263,N_913);
nor U1119 (N_1119,N_907,N_248);
nand U1120 (N_1120,N_286,N_245);
nand U1121 (N_1121,N_21,N_383);
xor U1122 (N_1122,N_257,N_207);
and U1123 (N_1123,N_45,N_773);
or U1124 (N_1124,N_443,N_405);
xnor U1125 (N_1125,N_894,N_113);
nand U1126 (N_1126,N_757,N_65);
nor U1127 (N_1127,N_156,N_14);
xnor U1128 (N_1128,N_872,N_904);
and U1129 (N_1129,N_942,N_856);
and U1130 (N_1130,N_222,N_188);
or U1131 (N_1131,N_886,N_999);
nor U1132 (N_1132,N_859,N_739);
nor U1133 (N_1133,N_229,N_590);
nor U1134 (N_1134,N_548,N_460);
or U1135 (N_1135,N_979,N_440);
nand U1136 (N_1136,N_662,N_432);
nor U1137 (N_1137,N_795,N_3);
xor U1138 (N_1138,N_452,N_218);
and U1139 (N_1139,N_709,N_334);
xnor U1140 (N_1140,N_688,N_227);
nand U1141 (N_1141,N_852,N_871);
or U1142 (N_1142,N_760,N_934);
or U1143 (N_1143,N_168,N_835);
and U1144 (N_1144,N_25,N_726);
nor U1145 (N_1145,N_697,N_112);
nor U1146 (N_1146,N_346,N_172);
nand U1147 (N_1147,N_575,N_349);
and U1148 (N_1148,N_986,N_853);
nand U1149 (N_1149,N_611,N_115);
nor U1150 (N_1150,N_509,N_716);
or U1151 (N_1151,N_654,N_561);
and U1152 (N_1152,N_943,N_449);
nand U1153 (N_1153,N_247,N_501);
xor U1154 (N_1154,N_899,N_820);
xor U1155 (N_1155,N_649,N_552);
or U1156 (N_1156,N_821,N_873);
or U1157 (N_1157,N_374,N_976);
nand U1158 (N_1158,N_759,N_278);
or U1159 (N_1159,N_336,N_108);
nand U1160 (N_1160,N_487,N_485);
nand U1161 (N_1161,N_936,N_830);
nand U1162 (N_1162,N_801,N_802);
or U1163 (N_1163,N_150,N_354);
and U1164 (N_1164,N_643,N_146);
nand U1165 (N_1165,N_288,N_427);
nand U1166 (N_1166,N_406,N_10);
and U1167 (N_1167,N_152,N_59);
nand U1168 (N_1168,N_468,N_924);
or U1169 (N_1169,N_911,N_787);
nor U1170 (N_1170,N_832,N_2);
and U1171 (N_1171,N_238,N_436);
or U1172 (N_1172,N_816,N_434);
nor U1173 (N_1173,N_511,N_289);
nor U1174 (N_1174,N_992,N_505);
nor U1175 (N_1175,N_127,N_721);
or U1176 (N_1176,N_335,N_167);
and U1177 (N_1177,N_607,N_57);
and U1178 (N_1178,N_606,N_589);
nand U1179 (N_1179,N_9,N_922);
or U1180 (N_1180,N_559,N_446);
nand U1181 (N_1181,N_0,N_198);
nand U1182 (N_1182,N_637,N_946);
or U1183 (N_1183,N_133,N_117);
or U1184 (N_1184,N_489,N_160);
and U1185 (N_1185,N_412,N_545);
or U1186 (N_1186,N_490,N_361);
or U1187 (N_1187,N_407,N_534);
and U1188 (N_1188,N_765,N_745);
nor U1189 (N_1189,N_826,N_439);
or U1190 (N_1190,N_956,N_442);
and U1191 (N_1191,N_85,N_350);
nand U1192 (N_1192,N_197,N_808);
and U1193 (N_1193,N_809,N_416);
xor U1194 (N_1194,N_850,N_768);
nor U1195 (N_1195,N_653,N_703);
xnor U1196 (N_1196,N_16,N_250);
and U1197 (N_1197,N_471,N_121);
or U1198 (N_1198,N_333,N_526);
nand U1199 (N_1199,N_272,N_395);
nand U1200 (N_1200,N_411,N_144);
xnor U1201 (N_1201,N_828,N_137);
nor U1202 (N_1202,N_424,N_28);
nand U1203 (N_1203,N_319,N_226);
and U1204 (N_1204,N_264,N_539);
and U1205 (N_1205,N_404,N_345);
and U1206 (N_1206,N_733,N_231);
or U1207 (N_1207,N_29,N_758);
xor U1208 (N_1208,N_551,N_965);
nor U1209 (N_1209,N_52,N_522);
and U1210 (N_1210,N_642,N_342);
and U1211 (N_1211,N_948,N_546);
xnor U1212 (N_1212,N_428,N_474);
xnor U1213 (N_1213,N_299,N_297);
nand U1214 (N_1214,N_650,N_775);
and U1215 (N_1215,N_734,N_100);
xnor U1216 (N_1216,N_582,N_276);
nor U1217 (N_1217,N_120,N_634);
xnor U1218 (N_1218,N_563,N_790);
and U1219 (N_1219,N_837,N_129);
nor U1220 (N_1220,N_690,N_981);
or U1221 (N_1221,N_196,N_529);
xnor U1222 (N_1222,N_910,N_389);
nor U1223 (N_1223,N_842,N_663);
xor U1224 (N_1224,N_960,N_877);
nand U1225 (N_1225,N_762,N_710);
xnor U1226 (N_1226,N_989,N_124);
nand U1227 (N_1227,N_310,N_736);
or U1228 (N_1228,N_961,N_450);
and U1229 (N_1229,N_419,N_695);
nand U1230 (N_1230,N_295,N_475);
and U1231 (N_1231,N_764,N_527);
and U1232 (N_1232,N_538,N_998);
or U1233 (N_1233,N_536,N_645);
xor U1234 (N_1234,N_977,N_390);
and U1235 (N_1235,N_34,N_256);
nand U1236 (N_1236,N_513,N_12);
xnor U1237 (N_1237,N_870,N_823);
nor U1238 (N_1238,N_967,N_951);
nand U1239 (N_1239,N_963,N_752);
or U1240 (N_1240,N_630,N_732);
nor U1241 (N_1241,N_301,N_970);
and U1242 (N_1242,N_556,N_51);
nor U1243 (N_1243,N_735,N_860);
xnor U1244 (N_1244,N_41,N_565);
and U1245 (N_1245,N_233,N_723);
xor U1246 (N_1246,N_949,N_418);
or U1247 (N_1247,N_581,N_782);
and U1248 (N_1248,N_603,N_619);
and U1249 (N_1249,N_594,N_158);
nor U1250 (N_1250,N_481,N_867);
and U1251 (N_1251,N_495,N_37);
xor U1252 (N_1252,N_772,N_282);
and U1253 (N_1253,N_164,N_40);
or U1254 (N_1254,N_318,N_641);
or U1255 (N_1255,N_959,N_766);
nand U1256 (N_1256,N_644,N_43);
nand U1257 (N_1257,N_524,N_737);
or U1258 (N_1258,N_825,N_122);
xor U1259 (N_1259,N_358,N_314);
nor U1260 (N_1260,N_504,N_394);
and U1261 (N_1261,N_232,N_382);
xnor U1262 (N_1262,N_595,N_969);
nor U1263 (N_1263,N_964,N_4);
and U1264 (N_1264,N_621,N_627);
nand U1265 (N_1265,N_670,N_786);
nand U1266 (N_1266,N_491,N_811);
and U1267 (N_1267,N_796,N_875);
nand U1268 (N_1268,N_415,N_699);
nor U1269 (N_1269,N_937,N_715);
nand U1270 (N_1270,N_770,N_799);
or U1271 (N_1271,N_549,N_375);
or U1272 (N_1272,N_748,N_79);
xnor U1273 (N_1273,N_767,N_492);
and U1274 (N_1274,N_75,N_132);
and U1275 (N_1275,N_96,N_42);
nand U1276 (N_1276,N_324,N_305);
or U1277 (N_1277,N_704,N_869);
nand U1278 (N_1278,N_30,N_180);
nand U1279 (N_1279,N_950,N_923);
nor U1280 (N_1280,N_353,N_142);
nor U1281 (N_1281,N_519,N_95);
and U1282 (N_1282,N_600,N_138);
nand U1283 (N_1283,N_838,N_624);
or U1284 (N_1284,N_508,N_327);
nand U1285 (N_1285,N_69,N_306);
and U1286 (N_1286,N_897,N_680);
or U1287 (N_1287,N_694,N_294);
or U1288 (N_1288,N_277,N_685);
nor U1289 (N_1289,N_67,N_210);
and U1290 (N_1290,N_157,N_309);
nor U1291 (N_1291,N_435,N_616);
nor U1292 (N_1292,N_890,N_93);
nand U1293 (N_1293,N_237,N_154);
nand U1294 (N_1294,N_930,N_348);
xor U1295 (N_1295,N_145,N_244);
or U1296 (N_1296,N_386,N_378);
nand U1297 (N_1297,N_316,N_714);
nor U1298 (N_1298,N_713,N_803);
or U1299 (N_1299,N_271,N_953);
nor U1300 (N_1300,N_917,N_901);
or U1301 (N_1301,N_657,N_639);
or U1302 (N_1302,N_58,N_810);
nor U1303 (N_1303,N_136,N_13);
nand U1304 (N_1304,N_24,N_592);
nor U1305 (N_1305,N_265,N_591);
nand U1306 (N_1306,N_252,N_507);
and U1307 (N_1307,N_622,N_402);
xnor U1308 (N_1308,N_239,N_818);
xor U1309 (N_1309,N_396,N_725);
xnor U1310 (N_1310,N_792,N_615);
xnor U1311 (N_1311,N_477,N_847);
or U1312 (N_1312,N_425,N_995);
and U1313 (N_1313,N_541,N_15);
nand U1314 (N_1314,N_338,N_746);
nand U1315 (N_1315,N_332,N_414);
nor U1316 (N_1316,N_368,N_189);
nand U1317 (N_1317,N_608,N_104);
and U1318 (N_1318,N_330,N_46);
xor U1319 (N_1319,N_669,N_855);
or U1320 (N_1320,N_781,N_833);
or U1321 (N_1321,N_926,N_243);
xor U1322 (N_1322,N_660,N_612);
xnor U1323 (N_1323,N_287,N_369);
or U1324 (N_1324,N_834,N_134);
xnor U1325 (N_1325,N_909,N_8);
or U1326 (N_1326,N_996,N_114);
nor U1327 (N_1327,N_844,N_47);
xor U1328 (N_1328,N_275,N_915);
nand U1329 (N_1329,N_932,N_91);
nor U1330 (N_1330,N_400,N_456);
and U1331 (N_1331,N_214,N_854);
and U1332 (N_1332,N_80,N_499);
and U1333 (N_1333,N_63,N_486);
and U1334 (N_1334,N_696,N_453);
or U1335 (N_1335,N_340,N_711);
nand U1336 (N_1336,N_364,N_693);
or U1337 (N_1337,N_465,N_192);
nor U1338 (N_1338,N_903,N_659);
xnor U1339 (N_1339,N_931,N_195);
xor U1340 (N_1340,N_308,N_70);
and U1341 (N_1341,N_171,N_55);
nor U1342 (N_1342,N_700,N_478);
xnor U1343 (N_1343,N_530,N_268);
xnor U1344 (N_1344,N_209,N_202);
nor U1345 (N_1345,N_322,N_925);
nor U1346 (N_1346,N_974,N_217);
or U1347 (N_1347,N_355,N_367);
or U1348 (N_1348,N_179,N_658);
or U1349 (N_1349,N_691,N_665);
nor U1350 (N_1350,N_173,N_927);
nor U1351 (N_1351,N_566,N_807);
nor U1352 (N_1352,N_94,N_793);
and U1353 (N_1353,N_82,N_140);
nor U1354 (N_1354,N_780,N_896);
and U1355 (N_1355,N_23,N_22);
xor U1356 (N_1356,N_884,N_463);
and U1357 (N_1357,N_78,N_885);
or U1358 (N_1358,N_861,N_640);
nor U1359 (N_1359,N_701,N_223);
and U1360 (N_1360,N_604,N_678);
nor U1361 (N_1361,N_822,N_397);
xor U1362 (N_1362,N_236,N_610);
and U1363 (N_1363,N_86,N_664);
nand U1364 (N_1364,N_130,N_971);
nand U1365 (N_1365,N_159,N_66);
nor U1366 (N_1366,N_97,N_77);
nand U1367 (N_1367,N_311,N_553);
xnor U1368 (N_1368,N_982,N_588);
and U1369 (N_1369,N_506,N_887);
nor U1370 (N_1370,N_261,N_929);
or U1371 (N_1371,N_730,N_116);
xnor U1372 (N_1372,N_200,N_119);
xnor U1373 (N_1373,N_351,N_76);
xnor U1374 (N_1374,N_53,N_426);
nor U1375 (N_1375,N_469,N_413);
nand U1376 (N_1376,N_462,N_61);
xor U1377 (N_1377,N_994,N_980);
and U1378 (N_1378,N_631,N_857);
and U1379 (N_1379,N_56,N_879);
nand U1380 (N_1380,N_410,N_858);
and U1381 (N_1381,N_626,N_648);
nor U1382 (N_1382,N_357,N_955);
nand U1383 (N_1383,N_123,N_814);
or U1384 (N_1384,N_399,N_7);
or U1385 (N_1385,N_128,N_656);
nor U1386 (N_1386,N_454,N_791);
or U1387 (N_1387,N_525,N_441);
or U1388 (N_1388,N_184,N_515);
xor U1389 (N_1389,N_707,N_749);
nand U1390 (N_1390,N_920,N_429);
nand U1391 (N_1391,N_517,N_38);
nor U1392 (N_1392,N_88,N_356);
xor U1393 (N_1393,N_572,N_27);
nand U1394 (N_1394,N_851,N_761);
nand U1395 (N_1395,N_194,N_101);
nand U1396 (N_1396,N_203,N_893);
nand U1397 (N_1397,N_181,N_789);
and U1398 (N_1398,N_32,N_973);
and U1399 (N_1399,N_225,N_190);
or U1400 (N_1400,N_584,N_655);
and U1401 (N_1401,N_176,N_254);
xnor U1402 (N_1402,N_840,N_185);
or U1403 (N_1403,N_628,N_304);
and U1404 (N_1404,N_92,N_279);
and U1405 (N_1405,N_326,N_183);
or U1406 (N_1406,N_741,N_329);
nor U1407 (N_1407,N_676,N_365);
or U1408 (N_1408,N_687,N_337);
nor U1409 (N_1409,N_583,N_494);
nand U1410 (N_1410,N_940,N_444);
and U1411 (N_1411,N_451,N_398);
or U1412 (N_1412,N_881,N_576);
and U1413 (N_1413,N_325,N_747);
nand U1414 (N_1414,N_211,N_20);
nor U1415 (N_1415,N_518,N_712);
xnor U1416 (N_1416,N_972,N_783);
nand U1417 (N_1417,N_599,N_379);
xnor U1418 (N_1418,N_865,N_302);
and U1419 (N_1419,N_298,N_891);
and U1420 (N_1420,N_163,N_636);
or U1421 (N_1421,N_193,N_488);
nor U1422 (N_1422,N_564,N_35);
nand U1423 (N_1423,N_403,N_376);
nor U1424 (N_1424,N_593,N_493);
and U1425 (N_1425,N_479,N_668);
and U1426 (N_1426,N_947,N_824);
nor U1427 (N_1427,N_862,N_422);
and U1428 (N_1428,N_797,N_537);
and U1429 (N_1429,N_118,N_568);
nor U1430 (N_1430,N_609,N_111);
nor U1431 (N_1431,N_708,N_73);
or U1432 (N_1432,N_921,N_105);
xnor U1433 (N_1433,N_804,N_321);
and U1434 (N_1434,N_928,N_177);
and U1435 (N_1435,N_430,N_698);
nand U1436 (N_1436,N_987,N_259);
nor U1437 (N_1437,N_580,N_839);
or U1438 (N_1438,N_303,N_689);
nor U1439 (N_1439,N_585,N_774);
or U1440 (N_1440,N_933,N_958);
or U1441 (N_1441,N_251,N_447);
nand U1442 (N_1442,N_391,N_902);
nand U1443 (N_1443,N_81,N_260);
nand U1444 (N_1444,N_754,N_187);
nand U1445 (N_1445,N_635,N_535);
xnor U1446 (N_1446,N_667,N_722);
or U1447 (N_1447,N_344,N_966);
or U1448 (N_1448,N_255,N_373);
or U1449 (N_1449,N_751,N_230);
and U1450 (N_1450,N_829,N_954);
xor U1451 (N_1451,N_36,N_679);
nand U1452 (N_1452,N_521,N_496);
xor U1453 (N_1453,N_125,N_467);
xor U1454 (N_1454,N_617,N_11);
nor U1455 (N_1455,N_618,N_502);
and U1456 (N_1456,N_938,N_652);
xnor U1457 (N_1457,N_281,N_445);
nand U1458 (N_1458,N_916,N_249);
nand U1459 (N_1459,N_33,N_39);
nand U1460 (N_1460,N_267,N_107);
nand U1461 (N_1461,N_729,N_883);
and U1462 (N_1462,N_384,N_516);
nor U1463 (N_1463,N_246,N_359);
nand U1464 (N_1464,N_719,N_360);
and U1465 (N_1465,N_554,N_169);
or U1466 (N_1466,N_68,N_372);
nand U1467 (N_1467,N_562,N_579);
and U1468 (N_1468,N_983,N_31);
and U1469 (N_1469,N_381,N_750);
xnor U1470 (N_1470,N_532,N_408);
nor U1471 (N_1471,N_470,N_49);
nand U1472 (N_1472,N_684,N_952);
or U1473 (N_1473,N_800,N_945);
or U1474 (N_1474,N_975,N_740);
or U1475 (N_1475,N_421,N_510);
or U1476 (N_1476,N_742,N_44);
and U1477 (N_1477,N_778,N_270);
nor U1478 (N_1478,N_985,N_613);
or U1479 (N_1479,N_550,N_544);
and U1480 (N_1480,N_110,N_962);
xnor U1481 (N_1481,N_671,N_409);
nor U1482 (N_1482,N_547,N_846);
nand U1483 (N_1483,N_291,N_498);
nor U1484 (N_1484,N_661,N_738);
or U1485 (N_1485,N_638,N_458);
xnor U1486 (N_1486,N_601,N_686);
nor U1487 (N_1487,N_293,N_292);
or U1488 (N_1488,N_175,N_831);
and U1489 (N_1489,N_596,N_102);
nand U1490 (N_1490,N_718,N_352);
or U1491 (N_1491,N_213,N_258);
nand U1492 (N_1492,N_362,N_417);
and U1493 (N_1493,N_633,N_812);
nand U1494 (N_1494,N_753,N_533);
xnor U1495 (N_1495,N_253,N_779);
nand U1496 (N_1496,N_371,N_673);
or U1497 (N_1497,N_614,N_393);
xnor U1498 (N_1498,N_756,N_274);
or U1499 (N_1499,N_315,N_560);
nand U1500 (N_1500,N_735,N_293);
nand U1501 (N_1501,N_442,N_566);
and U1502 (N_1502,N_1,N_849);
xnor U1503 (N_1503,N_196,N_325);
and U1504 (N_1504,N_427,N_541);
xnor U1505 (N_1505,N_743,N_437);
nor U1506 (N_1506,N_698,N_584);
nor U1507 (N_1507,N_111,N_448);
nor U1508 (N_1508,N_207,N_810);
xor U1509 (N_1509,N_660,N_513);
or U1510 (N_1510,N_769,N_74);
nand U1511 (N_1511,N_148,N_420);
nand U1512 (N_1512,N_588,N_14);
nand U1513 (N_1513,N_492,N_661);
nor U1514 (N_1514,N_509,N_114);
xor U1515 (N_1515,N_209,N_465);
or U1516 (N_1516,N_211,N_280);
or U1517 (N_1517,N_495,N_975);
or U1518 (N_1518,N_826,N_143);
xnor U1519 (N_1519,N_29,N_419);
nor U1520 (N_1520,N_540,N_59);
xnor U1521 (N_1521,N_437,N_87);
nand U1522 (N_1522,N_574,N_16);
or U1523 (N_1523,N_705,N_345);
xnor U1524 (N_1524,N_201,N_70);
nor U1525 (N_1525,N_411,N_953);
and U1526 (N_1526,N_403,N_333);
nor U1527 (N_1527,N_20,N_413);
or U1528 (N_1528,N_880,N_868);
or U1529 (N_1529,N_387,N_174);
nor U1530 (N_1530,N_916,N_700);
nor U1531 (N_1531,N_313,N_885);
nor U1532 (N_1532,N_272,N_604);
nand U1533 (N_1533,N_238,N_631);
xnor U1534 (N_1534,N_300,N_356);
nor U1535 (N_1535,N_545,N_115);
nor U1536 (N_1536,N_171,N_215);
and U1537 (N_1537,N_830,N_556);
and U1538 (N_1538,N_450,N_407);
and U1539 (N_1539,N_340,N_519);
nand U1540 (N_1540,N_340,N_980);
nand U1541 (N_1541,N_527,N_955);
xnor U1542 (N_1542,N_560,N_40);
xor U1543 (N_1543,N_702,N_627);
nand U1544 (N_1544,N_253,N_54);
or U1545 (N_1545,N_716,N_84);
nor U1546 (N_1546,N_704,N_455);
nand U1547 (N_1547,N_202,N_893);
and U1548 (N_1548,N_357,N_808);
and U1549 (N_1549,N_955,N_286);
and U1550 (N_1550,N_693,N_753);
nand U1551 (N_1551,N_594,N_8);
xnor U1552 (N_1552,N_737,N_877);
nor U1553 (N_1553,N_43,N_671);
or U1554 (N_1554,N_544,N_49);
or U1555 (N_1555,N_159,N_703);
and U1556 (N_1556,N_445,N_211);
xor U1557 (N_1557,N_342,N_772);
and U1558 (N_1558,N_997,N_922);
nand U1559 (N_1559,N_912,N_931);
nor U1560 (N_1560,N_238,N_512);
nand U1561 (N_1561,N_68,N_712);
nand U1562 (N_1562,N_479,N_718);
nor U1563 (N_1563,N_397,N_448);
xor U1564 (N_1564,N_266,N_228);
xnor U1565 (N_1565,N_373,N_765);
and U1566 (N_1566,N_136,N_819);
nor U1567 (N_1567,N_855,N_520);
and U1568 (N_1568,N_857,N_601);
or U1569 (N_1569,N_730,N_775);
nand U1570 (N_1570,N_594,N_527);
nand U1571 (N_1571,N_838,N_772);
nor U1572 (N_1572,N_233,N_48);
nor U1573 (N_1573,N_246,N_691);
xnor U1574 (N_1574,N_887,N_920);
or U1575 (N_1575,N_690,N_908);
xor U1576 (N_1576,N_220,N_103);
or U1577 (N_1577,N_114,N_582);
and U1578 (N_1578,N_184,N_343);
nand U1579 (N_1579,N_590,N_318);
or U1580 (N_1580,N_465,N_244);
or U1581 (N_1581,N_202,N_3);
nand U1582 (N_1582,N_988,N_325);
nor U1583 (N_1583,N_910,N_291);
nor U1584 (N_1584,N_307,N_174);
xor U1585 (N_1585,N_984,N_939);
nand U1586 (N_1586,N_483,N_168);
nand U1587 (N_1587,N_542,N_327);
nand U1588 (N_1588,N_646,N_736);
xor U1589 (N_1589,N_664,N_569);
xnor U1590 (N_1590,N_584,N_624);
nand U1591 (N_1591,N_662,N_126);
and U1592 (N_1592,N_282,N_942);
xor U1593 (N_1593,N_411,N_716);
xor U1594 (N_1594,N_975,N_531);
nand U1595 (N_1595,N_205,N_799);
nor U1596 (N_1596,N_172,N_360);
or U1597 (N_1597,N_719,N_747);
nor U1598 (N_1598,N_608,N_746);
and U1599 (N_1599,N_368,N_211);
or U1600 (N_1600,N_825,N_865);
or U1601 (N_1601,N_430,N_123);
nand U1602 (N_1602,N_391,N_318);
xor U1603 (N_1603,N_478,N_885);
xor U1604 (N_1604,N_350,N_563);
nand U1605 (N_1605,N_879,N_79);
or U1606 (N_1606,N_677,N_343);
or U1607 (N_1607,N_542,N_417);
xnor U1608 (N_1608,N_427,N_118);
xor U1609 (N_1609,N_824,N_79);
xor U1610 (N_1610,N_263,N_717);
and U1611 (N_1611,N_534,N_47);
nand U1612 (N_1612,N_93,N_828);
xor U1613 (N_1613,N_727,N_817);
nor U1614 (N_1614,N_868,N_224);
xnor U1615 (N_1615,N_66,N_247);
and U1616 (N_1616,N_50,N_44);
nand U1617 (N_1617,N_147,N_255);
nor U1618 (N_1618,N_774,N_52);
or U1619 (N_1619,N_297,N_848);
xor U1620 (N_1620,N_557,N_259);
nor U1621 (N_1621,N_741,N_569);
and U1622 (N_1622,N_604,N_223);
nand U1623 (N_1623,N_574,N_713);
or U1624 (N_1624,N_629,N_800);
nor U1625 (N_1625,N_841,N_210);
nand U1626 (N_1626,N_336,N_452);
xor U1627 (N_1627,N_704,N_783);
nand U1628 (N_1628,N_639,N_280);
nor U1629 (N_1629,N_274,N_826);
nor U1630 (N_1630,N_12,N_90);
nand U1631 (N_1631,N_609,N_894);
and U1632 (N_1632,N_601,N_291);
nand U1633 (N_1633,N_877,N_414);
nor U1634 (N_1634,N_809,N_134);
or U1635 (N_1635,N_431,N_499);
or U1636 (N_1636,N_836,N_947);
nor U1637 (N_1637,N_213,N_185);
xor U1638 (N_1638,N_9,N_95);
xnor U1639 (N_1639,N_862,N_883);
and U1640 (N_1640,N_235,N_457);
and U1641 (N_1641,N_540,N_456);
and U1642 (N_1642,N_54,N_928);
nand U1643 (N_1643,N_883,N_585);
nor U1644 (N_1644,N_883,N_955);
and U1645 (N_1645,N_350,N_222);
nand U1646 (N_1646,N_86,N_39);
or U1647 (N_1647,N_657,N_507);
and U1648 (N_1648,N_591,N_385);
xnor U1649 (N_1649,N_773,N_233);
xor U1650 (N_1650,N_459,N_235);
or U1651 (N_1651,N_81,N_995);
and U1652 (N_1652,N_601,N_207);
or U1653 (N_1653,N_140,N_767);
xor U1654 (N_1654,N_761,N_588);
nand U1655 (N_1655,N_308,N_541);
or U1656 (N_1656,N_824,N_559);
nand U1657 (N_1657,N_985,N_303);
nand U1658 (N_1658,N_797,N_425);
or U1659 (N_1659,N_883,N_513);
nand U1660 (N_1660,N_760,N_653);
nand U1661 (N_1661,N_2,N_925);
xnor U1662 (N_1662,N_754,N_148);
xnor U1663 (N_1663,N_957,N_201);
or U1664 (N_1664,N_459,N_828);
nand U1665 (N_1665,N_995,N_653);
or U1666 (N_1666,N_816,N_358);
or U1667 (N_1667,N_372,N_764);
nand U1668 (N_1668,N_170,N_831);
or U1669 (N_1669,N_702,N_810);
or U1670 (N_1670,N_796,N_160);
or U1671 (N_1671,N_567,N_743);
and U1672 (N_1672,N_959,N_5);
xnor U1673 (N_1673,N_817,N_224);
or U1674 (N_1674,N_31,N_368);
nand U1675 (N_1675,N_100,N_488);
xor U1676 (N_1676,N_40,N_669);
nand U1677 (N_1677,N_846,N_850);
nor U1678 (N_1678,N_394,N_862);
and U1679 (N_1679,N_169,N_343);
nand U1680 (N_1680,N_4,N_353);
and U1681 (N_1681,N_361,N_750);
xnor U1682 (N_1682,N_527,N_931);
nor U1683 (N_1683,N_243,N_302);
nand U1684 (N_1684,N_88,N_0);
or U1685 (N_1685,N_62,N_732);
and U1686 (N_1686,N_622,N_768);
nor U1687 (N_1687,N_512,N_557);
or U1688 (N_1688,N_934,N_74);
or U1689 (N_1689,N_910,N_491);
or U1690 (N_1690,N_169,N_170);
nand U1691 (N_1691,N_149,N_899);
nand U1692 (N_1692,N_819,N_75);
nor U1693 (N_1693,N_173,N_126);
nor U1694 (N_1694,N_383,N_24);
nor U1695 (N_1695,N_774,N_532);
nor U1696 (N_1696,N_725,N_935);
or U1697 (N_1697,N_617,N_22);
and U1698 (N_1698,N_870,N_374);
nand U1699 (N_1699,N_361,N_147);
and U1700 (N_1700,N_819,N_889);
and U1701 (N_1701,N_959,N_497);
xor U1702 (N_1702,N_735,N_244);
or U1703 (N_1703,N_947,N_130);
nand U1704 (N_1704,N_830,N_31);
and U1705 (N_1705,N_48,N_567);
and U1706 (N_1706,N_406,N_843);
nand U1707 (N_1707,N_137,N_173);
nand U1708 (N_1708,N_928,N_676);
and U1709 (N_1709,N_609,N_64);
xor U1710 (N_1710,N_90,N_162);
and U1711 (N_1711,N_895,N_475);
nor U1712 (N_1712,N_854,N_402);
nor U1713 (N_1713,N_717,N_174);
nor U1714 (N_1714,N_657,N_904);
nor U1715 (N_1715,N_55,N_801);
xor U1716 (N_1716,N_68,N_617);
and U1717 (N_1717,N_267,N_615);
nor U1718 (N_1718,N_727,N_189);
xor U1719 (N_1719,N_879,N_736);
or U1720 (N_1720,N_667,N_313);
nor U1721 (N_1721,N_762,N_844);
xor U1722 (N_1722,N_976,N_900);
nand U1723 (N_1723,N_731,N_945);
nor U1724 (N_1724,N_394,N_262);
or U1725 (N_1725,N_205,N_258);
and U1726 (N_1726,N_361,N_446);
xor U1727 (N_1727,N_638,N_658);
nor U1728 (N_1728,N_391,N_390);
nand U1729 (N_1729,N_905,N_111);
nor U1730 (N_1730,N_244,N_859);
and U1731 (N_1731,N_184,N_713);
xnor U1732 (N_1732,N_970,N_921);
nor U1733 (N_1733,N_952,N_907);
xor U1734 (N_1734,N_860,N_596);
nor U1735 (N_1735,N_776,N_391);
nor U1736 (N_1736,N_939,N_216);
and U1737 (N_1737,N_166,N_97);
xnor U1738 (N_1738,N_321,N_265);
nand U1739 (N_1739,N_234,N_546);
nand U1740 (N_1740,N_965,N_353);
xnor U1741 (N_1741,N_658,N_117);
nand U1742 (N_1742,N_817,N_281);
nand U1743 (N_1743,N_713,N_643);
or U1744 (N_1744,N_773,N_776);
or U1745 (N_1745,N_931,N_980);
xor U1746 (N_1746,N_353,N_235);
nand U1747 (N_1747,N_957,N_64);
xor U1748 (N_1748,N_91,N_597);
or U1749 (N_1749,N_575,N_66);
or U1750 (N_1750,N_697,N_72);
or U1751 (N_1751,N_61,N_600);
xor U1752 (N_1752,N_246,N_582);
nor U1753 (N_1753,N_137,N_746);
and U1754 (N_1754,N_766,N_272);
and U1755 (N_1755,N_755,N_33);
nand U1756 (N_1756,N_687,N_501);
and U1757 (N_1757,N_707,N_509);
and U1758 (N_1758,N_809,N_822);
and U1759 (N_1759,N_333,N_269);
or U1760 (N_1760,N_716,N_274);
nor U1761 (N_1761,N_790,N_506);
or U1762 (N_1762,N_993,N_131);
xor U1763 (N_1763,N_765,N_659);
nand U1764 (N_1764,N_600,N_918);
nand U1765 (N_1765,N_862,N_667);
xor U1766 (N_1766,N_841,N_576);
and U1767 (N_1767,N_120,N_248);
or U1768 (N_1768,N_873,N_830);
xor U1769 (N_1769,N_588,N_896);
xor U1770 (N_1770,N_971,N_292);
or U1771 (N_1771,N_718,N_292);
nor U1772 (N_1772,N_947,N_715);
or U1773 (N_1773,N_727,N_433);
xnor U1774 (N_1774,N_537,N_75);
and U1775 (N_1775,N_126,N_85);
xor U1776 (N_1776,N_491,N_891);
and U1777 (N_1777,N_67,N_381);
and U1778 (N_1778,N_549,N_162);
nor U1779 (N_1779,N_276,N_837);
nor U1780 (N_1780,N_668,N_804);
or U1781 (N_1781,N_830,N_774);
nor U1782 (N_1782,N_411,N_149);
nand U1783 (N_1783,N_147,N_870);
or U1784 (N_1784,N_865,N_647);
and U1785 (N_1785,N_280,N_162);
xor U1786 (N_1786,N_986,N_344);
nand U1787 (N_1787,N_273,N_579);
or U1788 (N_1788,N_914,N_176);
nand U1789 (N_1789,N_763,N_394);
nor U1790 (N_1790,N_886,N_293);
nor U1791 (N_1791,N_548,N_133);
and U1792 (N_1792,N_118,N_634);
or U1793 (N_1793,N_443,N_49);
nor U1794 (N_1794,N_392,N_650);
nor U1795 (N_1795,N_411,N_699);
nor U1796 (N_1796,N_195,N_694);
nand U1797 (N_1797,N_419,N_626);
or U1798 (N_1798,N_389,N_33);
nor U1799 (N_1799,N_798,N_440);
nand U1800 (N_1800,N_69,N_759);
nand U1801 (N_1801,N_980,N_457);
xnor U1802 (N_1802,N_919,N_572);
xnor U1803 (N_1803,N_523,N_263);
nor U1804 (N_1804,N_650,N_317);
and U1805 (N_1805,N_227,N_205);
and U1806 (N_1806,N_606,N_84);
and U1807 (N_1807,N_985,N_779);
xnor U1808 (N_1808,N_761,N_285);
xnor U1809 (N_1809,N_682,N_927);
xnor U1810 (N_1810,N_85,N_166);
xnor U1811 (N_1811,N_39,N_879);
nor U1812 (N_1812,N_456,N_571);
and U1813 (N_1813,N_572,N_4);
nor U1814 (N_1814,N_693,N_106);
nand U1815 (N_1815,N_886,N_170);
xor U1816 (N_1816,N_351,N_857);
xor U1817 (N_1817,N_51,N_377);
nor U1818 (N_1818,N_915,N_651);
nand U1819 (N_1819,N_693,N_74);
xnor U1820 (N_1820,N_468,N_474);
nand U1821 (N_1821,N_726,N_312);
xor U1822 (N_1822,N_808,N_97);
nand U1823 (N_1823,N_289,N_300);
nand U1824 (N_1824,N_588,N_212);
and U1825 (N_1825,N_460,N_944);
xor U1826 (N_1826,N_261,N_242);
xnor U1827 (N_1827,N_112,N_948);
nand U1828 (N_1828,N_996,N_947);
nor U1829 (N_1829,N_848,N_179);
xnor U1830 (N_1830,N_319,N_628);
nand U1831 (N_1831,N_465,N_676);
nand U1832 (N_1832,N_113,N_465);
and U1833 (N_1833,N_391,N_304);
nand U1834 (N_1834,N_641,N_410);
or U1835 (N_1835,N_675,N_137);
xnor U1836 (N_1836,N_938,N_734);
or U1837 (N_1837,N_392,N_979);
nor U1838 (N_1838,N_819,N_7);
nor U1839 (N_1839,N_488,N_569);
xnor U1840 (N_1840,N_315,N_816);
and U1841 (N_1841,N_57,N_278);
and U1842 (N_1842,N_591,N_296);
and U1843 (N_1843,N_627,N_699);
or U1844 (N_1844,N_524,N_252);
nor U1845 (N_1845,N_835,N_935);
nand U1846 (N_1846,N_435,N_477);
nand U1847 (N_1847,N_257,N_420);
and U1848 (N_1848,N_202,N_884);
nor U1849 (N_1849,N_604,N_521);
nor U1850 (N_1850,N_103,N_8);
or U1851 (N_1851,N_851,N_245);
or U1852 (N_1852,N_492,N_537);
xor U1853 (N_1853,N_651,N_419);
and U1854 (N_1854,N_602,N_25);
nor U1855 (N_1855,N_388,N_69);
and U1856 (N_1856,N_633,N_204);
or U1857 (N_1857,N_812,N_630);
or U1858 (N_1858,N_852,N_786);
nor U1859 (N_1859,N_843,N_367);
nand U1860 (N_1860,N_354,N_604);
xor U1861 (N_1861,N_415,N_603);
nor U1862 (N_1862,N_260,N_937);
and U1863 (N_1863,N_58,N_754);
nor U1864 (N_1864,N_76,N_2);
nor U1865 (N_1865,N_909,N_570);
nand U1866 (N_1866,N_260,N_833);
nor U1867 (N_1867,N_658,N_505);
nor U1868 (N_1868,N_247,N_525);
nand U1869 (N_1869,N_46,N_761);
nand U1870 (N_1870,N_358,N_798);
or U1871 (N_1871,N_189,N_115);
xnor U1872 (N_1872,N_333,N_987);
xor U1873 (N_1873,N_245,N_834);
and U1874 (N_1874,N_283,N_140);
and U1875 (N_1875,N_899,N_421);
or U1876 (N_1876,N_57,N_938);
and U1877 (N_1877,N_564,N_194);
xor U1878 (N_1878,N_285,N_114);
or U1879 (N_1879,N_842,N_196);
nor U1880 (N_1880,N_331,N_177);
or U1881 (N_1881,N_715,N_468);
or U1882 (N_1882,N_997,N_226);
xnor U1883 (N_1883,N_374,N_129);
nor U1884 (N_1884,N_383,N_947);
nand U1885 (N_1885,N_875,N_372);
xor U1886 (N_1886,N_602,N_646);
xor U1887 (N_1887,N_749,N_317);
and U1888 (N_1888,N_209,N_868);
or U1889 (N_1889,N_323,N_439);
xor U1890 (N_1890,N_512,N_418);
xor U1891 (N_1891,N_441,N_145);
and U1892 (N_1892,N_919,N_935);
nand U1893 (N_1893,N_940,N_574);
nand U1894 (N_1894,N_738,N_14);
or U1895 (N_1895,N_847,N_239);
xnor U1896 (N_1896,N_973,N_509);
or U1897 (N_1897,N_765,N_42);
or U1898 (N_1898,N_169,N_740);
nand U1899 (N_1899,N_537,N_650);
nand U1900 (N_1900,N_392,N_447);
and U1901 (N_1901,N_247,N_311);
xnor U1902 (N_1902,N_56,N_948);
nand U1903 (N_1903,N_727,N_934);
nor U1904 (N_1904,N_606,N_116);
nand U1905 (N_1905,N_713,N_121);
nand U1906 (N_1906,N_154,N_25);
nand U1907 (N_1907,N_656,N_788);
or U1908 (N_1908,N_301,N_162);
or U1909 (N_1909,N_979,N_117);
xor U1910 (N_1910,N_912,N_983);
or U1911 (N_1911,N_716,N_674);
or U1912 (N_1912,N_309,N_75);
nor U1913 (N_1913,N_928,N_163);
nand U1914 (N_1914,N_425,N_326);
nor U1915 (N_1915,N_598,N_336);
or U1916 (N_1916,N_153,N_449);
xor U1917 (N_1917,N_392,N_197);
nor U1918 (N_1918,N_741,N_73);
and U1919 (N_1919,N_637,N_764);
xnor U1920 (N_1920,N_54,N_916);
or U1921 (N_1921,N_959,N_842);
or U1922 (N_1922,N_426,N_408);
xnor U1923 (N_1923,N_862,N_923);
and U1924 (N_1924,N_505,N_936);
nor U1925 (N_1925,N_153,N_584);
nand U1926 (N_1926,N_443,N_172);
nor U1927 (N_1927,N_895,N_235);
nand U1928 (N_1928,N_312,N_513);
nor U1929 (N_1929,N_370,N_424);
nor U1930 (N_1930,N_473,N_509);
nor U1931 (N_1931,N_526,N_978);
or U1932 (N_1932,N_826,N_669);
or U1933 (N_1933,N_824,N_613);
nand U1934 (N_1934,N_929,N_285);
and U1935 (N_1935,N_374,N_597);
or U1936 (N_1936,N_653,N_83);
xor U1937 (N_1937,N_277,N_180);
nand U1938 (N_1938,N_894,N_215);
and U1939 (N_1939,N_864,N_134);
or U1940 (N_1940,N_95,N_843);
and U1941 (N_1941,N_296,N_528);
nor U1942 (N_1942,N_817,N_815);
nand U1943 (N_1943,N_625,N_994);
nand U1944 (N_1944,N_418,N_962);
nor U1945 (N_1945,N_543,N_388);
nor U1946 (N_1946,N_784,N_576);
nand U1947 (N_1947,N_970,N_992);
and U1948 (N_1948,N_922,N_926);
or U1949 (N_1949,N_275,N_585);
nand U1950 (N_1950,N_953,N_269);
nor U1951 (N_1951,N_822,N_418);
nor U1952 (N_1952,N_157,N_193);
nand U1953 (N_1953,N_833,N_963);
xor U1954 (N_1954,N_554,N_255);
or U1955 (N_1955,N_922,N_363);
xnor U1956 (N_1956,N_353,N_715);
nand U1957 (N_1957,N_466,N_91);
or U1958 (N_1958,N_832,N_701);
or U1959 (N_1959,N_867,N_619);
nor U1960 (N_1960,N_428,N_89);
nor U1961 (N_1961,N_614,N_331);
nand U1962 (N_1962,N_666,N_706);
xnor U1963 (N_1963,N_556,N_588);
nor U1964 (N_1964,N_827,N_464);
and U1965 (N_1965,N_682,N_811);
nand U1966 (N_1966,N_158,N_187);
nand U1967 (N_1967,N_666,N_429);
nor U1968 (N_1968,N_77,N_700);
or U1969 (N_1969,N_654,N_346);
or U1970 (N_1970,N_692,N_884);
xor U1971 (N_1971,N_252,N_977);
nand U1972 (N_1972,N_901,N_674);
xor U1973 (N_1973,N_549,N_45);
nand U1974 (N_1974,N_676,N_702);
and U1975 (N_1975,N_273,N_567);
or U1976 (N_1976,N_79,N_320);
xor U1977 (N_1977,N_590,N_687);
and U1978 (N_1978,N_862,N_223);
nor U1979 (N_1979,N_132,N_653);
nor U1980 (N_1980,N_296,N_382);
nor U1981 (N_1981,N_869,N_708);
nand U1982 (N_1982,N_213,N_265);
xnor U1983 (N_1983,N_488,N_663);
or U1984 (N_1984,N_503,N_407);
xnor U1985 (N_1985,N_582,N_55);
nor U1986 (N_1986,N_566,N_946);
and U1987 (N_1987,N_714,N_241);
nor U1988 (N_1988,N_989,N_972);
and U1989 (N_1989,N_262,N_794);
nand U1990 (N_1990,N_556,N_103);
xor U1991 (N_1991,N_585,N_53);
nand U1992 (N_1992,N_689,N_202);
and U1993 (N_1993,N_658,N_720);
nor U1994 (N_1994,N_257,N_539);
and U1995 (N_1995,N_884,N_713);
or U1996 (N_1996,N_339,N_125);
and U1997 (N_1997,N_28,N_593);
and U1998 (N_1998,N_992,N_629);
nand U1999 (N_1999,N_475,N_928);
or U2000 (N_2000,N_1451,N_1529);
nor U2001 (N_2001,N_1728,N_1426);
or U2002 (N_2002,N_1951,N_1011);
nand U2003 (N_2003,N_1394,N_1143);
nand U2004 (N_2004,N_1806,N_1329);
and U2005 (N_2005,N_1816,N_1095);
nand U2006 (N_2006,N_1714,N_1796);
or U2007 (N_2007,N_1646,N_1495);
nand U2008 (N_2008,N_1212,N_1820);
nand U2009 (N_2009,N_1175,N_1739);
or U2010 (N_2010,N_1323,N_1282);
xor U2011 (N_2011,N_1410,N_1837);
xnor U2012 (N_2012,N_1545,N_1150);
xnor U2013 (N_2013,N_1956,N_1051);
xor U2014 (N_2014,N_1761,N_1690);
nand U2015 (N_2015,N_1784,N_1035);
and U2016 (N_2016,N_1993,N_1102);
nor U2017 (N_2017,N_1340,N_1424);
nand U2018 (N_2018,N_1698,N_1662);
nor U2019 (N_2019,N_1841,N_1613);
or U2020 (N_2020,N_1116,N_1774);
nor U2021 (N_2021,N_1776,N_1049);
nor U2022 (N_2022,N_1239,N_1970);
nor U2023 (N_2023,N_1629,N_1139);
nand U2024 (N_2024,N_1429,N_1787);
xnor U2025 (N_2025,N_1607,N_1103);
and U2026 (N_2026,N_1555,N_1532);
or U2027 (N_2027,N_1125,N_1111);
and U2028 (N_2028,N_1798,N_1325);
nand U2029 (N_2029,N_1098,N_1355);
and U2030 (N_2030,N_1542,N_1588);
and U2031 (N_2031,N_1659,N_1528);
xnor U2032 (N_2032,N_1099,N_1127);
or U2033 (N_2033,N_1348,N_1884);
nand U2034 (N_2034,N_1168,N_1013);
nand U2035 (N_2035,N_1262,N_1014);
xor U2036 (N_2036,N_1151,N_1192);
xor U2037 (N_2037,N_1656,N_1414);
nor U2038 (N_2038,N_1474,N_1802);
nor U2039 (N_2039,N_1950,N_1668);
nor U2040 (N_2040,N_1893,N_1564);
and U2041 (N_2041,N_1493,N_1381);
and U2042 (N_2042,N_1135,N_1601);
nor U2043 (N_2043,N_1123,N_1670);
nand U2044 (N_2044,N_1031,N_1923);
xor U2045 (N_2045,N_1015,N_1310);
or U2046 (N_2046,N_1917,N_1374);
or U2047 (N_2047,N_1856,N_1744);
and U2048 (N_2048,N_1070,N_1830);
or U2049 (N_2049,N_1693,N_1485);
or U2050 (N_2050,N_1423,N_1634);
or U2051 (N_2051,N_1505,N_1782);
nand U2052 (N_2052,N_1315,N_1676);
or U2053 (N_2053,N_1199,N_1063);
nor U2054 (N_2054,N_1964,N_1751);
and U2055 (N_2055,N_1387,N_1560);
nand U2056 (N_2056,N_1688,N_1266);
nand U2057 (N_2057,N_1498,N_1600);
nor U2058 (N_2058,N_1045,N_1370);
or U2059 (N_2059,N_1009,N_1391);
and U2060 (N_2060,N_1172,N_1777);
or U2061 (N_2061,N_1454,N_1548);
and U2062 (N_2062,N_1664,N_1781);
xnor U2063 (N_2063,N_1213,N_1048);
nor U2064 (N_2064,N_1180,N_1492);
xnor U2065 (N_2065,N_1296,N_1399);
or U2066 (N_2066,N_1522,N_1385);
and U2067 (N_2067,N_1733,N_1930);
xor U2068 (N_2068,N_1022,N_1082);
or U2069 (N_2069,N_1582,N_1220);
xor U2070 (N_2070,N_1184,N_1138);
or U2071 (N_2071,N_1487,N_1539);
xor U2072 (N_2072,N_1718,N_1390);
and U2073 (N_2073,N_1276,N_1368);
nor U2074 (N_2074,N_1652,N_1680);
xnor U2075 (N_2075,N_1700,N_1566);
nand U2076 (N_2076,N_1218,N_1076);
nand U2077 (N_2077,N_1261,N_1617);
nand U2078 (N_2078,N_1913,N_1156);
nand U2079 (N_2079,N_1105,N_1915);
nor U2080 (N_2080,N_1996,N_1540);
and U2081 (N_2081,N_1640,N_1967);
and U2082 (N_2082,N_1779,N_1214);
or U2083 (N_2083,N_1023,N_1840);
xor U2084 (N_2084,N_1790,N_1242);
nor U2085 (N_2085,N_1585,N_1369);
nand U2086 (N_2086,N_1789,N_1421);
nand U2087 (N_2087,N_1875,N_1223);
nand U2088 (N_2088,N_1148,N_1435);
and U2089 (N_2089,N_1926,N_1365);
nand U2090 (N_2090,N_1230,N_1976);
nand U2091 (N_2091,N_1551,N_1635);
nand U2092 (N_2092,N_1822,N_1019);
nor U2093 (N_2093,N_1624,N_1060);
nor U2094 (N_2094,N_1232,N_1459);
nor U2095 (N_2095,N_1517,N_1354);
nor U2096 (N_2096,N_1734,N_1080);
nand U2097 (N_2097,N_1270,N_1701);
nand U2098 (N_2098,N_1267,N_1537);
nor U2099 (N_2099,N_1484,N_1050);
and U2100 (N_2100,N_1215,N_1389);
nor U2101 (N_2101,N_1181,N_1397);
and U2102 (N_2102,N_1715,N_1709);
or U2103 (N_2103,N_1762,N_1705);
and U2104 (N_2104,N_1749,N_1987);
nand U2105 (N_2105,N_1843,N_1895);
nor U2106 (N_2106,N_1256,N_1641);
or U2107 (N_2107,N_1874,N_1431);
and U2108 (N_2108,N_1592,N_1834);
and U2109 (N_2109,N_1274,N_1176);
or U2110 (N_2110,N_1977,N_1570);
nand U2111 (N_2111,N_1581,N_1314);
nor U2112 (N_2112,N_1727,N_1032);
nor U2113 (N_2113,N_1058,N_1773);
nand U2114 (N_2114,N_1377,N_1378);
xnor U2115 (N_2115,N_1625,N_1322);
xnor U2116 (N_2116,N_1189,N_1870);
and U2117 (N_2117,N_1170,N_1809);
and U2118 (N_2118,N_1633,N_1651);
nand U2119 (N_2119,N_1444,N_1699);
nor U2120 (N_2120,N_1083,N_1178);
xor U2121 (N_2121,N_1952,N_1141);
nand U2122 (N_2122,N_1469,N_1490);
or U2123 (N_2123,N_1210,N_1117);
xnor U2124 (N_2124,N_1330,N_1692);
and U2125 (N_2125,N_1860,N_1363);
xnor U2126 (N_2126,N_1631,N_1114);
nor U2127 (N_2127,N_1938,N_1188);
xnor U2128 (N_2128,N_1879,N_1754);
or U2129 (N_2129,N_1053,N_1963);
xor U2130 (N_2130,N_1826,N_1571);
nand U2131 (N_2131,N_1406,N_1654);
or U2132 (N_2132,N_1351,N_1061);
xnor U2133 (N_2133,N_1932,N_1765);
or U2134 (N_2134,N_1726,N_1954);
or U2135 (N_2135,N_1085,N_1136);
xnor U2136 (N_2136,N_1752,N_1708);
xor U2137 (N_2137,N_1758,N_1088);
nor U2138 (N_2138,N_1590,N_1476);
nand U2139 (N_2139,N_1200,N_1778);
nor U2140 (N_2140,N_1515,N_1272);
nand U2141 (N_2141,N_1612,N_1979);
xor U2142 (N_2142,N_1059,N_1033);
xnor U2143 (N_2143,N_1079,N_1383);
xnor U2144 (N_2144,N_1258,N_1093);
and U2145 (N_2145,N_1679,N_1801);
and U2146 (N_2146,N_1810,N_1823);
xor U2147 (N_2147,N_1149,N_1650);
or U2148 (N_2148,N_1717,N_1681);
or U2149 (N_2149,N_1824,N_1862);
nand U2150 (N_2150,N_1658,N_1040);
xor U2151 (N_2151,N_1850,N_1042);
or U2152 (N_2152,N_1614,N_1283);
nand U2153 (N_2153,N_1968,N_1236);
nand U2154 (N_2154,N_1317,N_1247);
nand U2155 (N_2155,N_1273,N_1328);
and U2156 (N_2156,N_1320,N_1575);
nor U2157 (N_2157,N_1392,N_1871);
and U2158 (N_2158,N_1027,N_1831);
or U2159 (N_2159,N_1024,N_1911);
xor U2160 (N_2160,N_1246,N_1417);
xnor U2161 (N_2161,N_1838,N_1825);
or U2162 (N_2162,N_1747,N_1685);
and U2163 (N_2163,N_1936,N_1939);
nor U2164 (N_2164,N_1249,N_1073);
nand U2165 (N_2165,N_1089,N_1846);
xnor U2166 (N_2166,N_1442,N_1710);
xor U2167 (N_2167,N_1240,N_1005);
nand U2168 (N_2168,N_1395,N_1942);
or U2169 (N_2169,N_1037,N_1064);
or U2170 (N_2170,N_1056,N_1286);
and U2171 (N_2171,N_1769,N_1881);
nor U2172 (N_2172,N_1300,N_1890);
nand U2173 (N_2173,N_1373,N_1508);
xnor U2174 (N_2174,N_1120,N_1554);
nor U2175 (N_2175,N_1853,N_1722);
or U2176 (N_2176,N_1947,N_1356);
or U2177 (N_2177,N_1546,N_1263);
and U2178 (N_2178,N_1524,N_1388);
xnor U2179 (N_2179,N_1494,N_1807);
nand U2180 (N_2180,N_1367,N_1422);
nand U2181 (N_2181,N_1233,N_1234);
nand U2182 (N_2182,N_1477,N_1396);
nor U2183 (N_2183,N_1922,N_1346);
xor U2184 (N_2184,N_1489,N_1580);
and U2185 (N_2185,N_1814,N_1780);
nand U2186 (N_2186,N_1413,N_1596);
xor U2187 (N_2187,N_1924,N_1731);
nand U2188 (N_2188,N_1157,N_1131);
nor U2189 (N_2189,N_1128,N_1497);
nor U2190 (N_2190,N_1159,N_1756);
or U2191 (N_2191,N_1799,N_1339);
and U2192 (N_2192,N_1966,N_1108);
and U2193 (N_2193,N_1092,N_1001);
nor U2194 (N_2194,N_1857,N_1880);
xor U2195 (N_2195,N_1632,N_1643);
nand U2196 (N_2196,N_1434,N_1158);
nor U2197 (N_2197,N_1649,N_1411);
xor U2198 (N_2198,N_1458,N_1671);
xnor U2199 (N_2199,N_1074,N_1735);
or U2200 (N_2200,N_1081,N_1347);
nor U2201 (N_2201,N_1353,N_1763);
xnor U2202 (N_2202,N_1195,N_1177);
and U2203 (N_2203,N_1994,N_1301);
nor U2204 (N_2204,N_1238,N_1479);
and U2205 (N_2205,N_1989,N_1606);
and U2206 (N_2206,N_1943,N_1109);
nor U2207 (N_2207,N_1309,N_1648);
xor U2208 (N_2208,N_1808,N_1729);
and U2209 (N_2209,N_1376,N_1420);
xnor U2210 (N_2210,N_1096,N_1738);
or U2211 (N_2211,N_1842,N_1360);
and U2212 (N_2212,N_1684,N_1137);
and U2213 (N_2213,N_1227,N_1750);
nand U2214 (N_2214,N_1552,N_1711);
and U2215 (N_2215,N_1400,N_1427);
and U2216 (N_2216,N_1721,N_1813);
nand U2217 (N_2217,N_1441,N_1990);
or U2218 (N_2218,N_1980,N_1271);
and U2219 (N_2219,N_1401,N_1338);
or U2220 (N_2220,N_1541,N_1304);
and U2221 (N_2221,N_1334,N_1983);
xnor U2222 (N_2222,N_1029,N_1337);
and U2223 (N_2223,N_1277,N_1350);
and U2224 (N_2224,N_1839,N_1386);
nand U2225 (N_2225,N_1669,N_1453);
nand U2226 (N_2226,N_1677,N_1844);
xnor U2227 (N_2227,N_1436,N_1878);
xnor U2228 (N_2228,N_1285,N_1847);
nor U2229 (N_2229,N_1342,N_1598);
nor U2230 (N_2230,N_1660,N_1294);
and U2231 (N_2231,N_1362,N_1891);
and U2232 (N_2232,N_1835,N_1785);
nor U2233 (N_2233,N_1297,N_1130);
and U2234 (N_2234,N_1534,N_1461);
or U2235 (N_2235,N_1740,N_1343);
xnor U2236 (N_2236,N_1892,N_1572);
nor U2237 (N_2237,N_1478,N_1775);
nand U2238 (N_2238,N_1403,N_1169);
or U2239 (N_2239,N_1129,N_1229);
nor U2240 (N_2240,N_1443,N_1584);
or U2241 (N_2241,N_1278,N_1628);
or U2242 (N_2242,N_1741,N_1591);
nor U2243 (N_2243,N_1961,N_1384);
and U2244 (N_2244,N_1193,N_1179);
and U2245 (N_2245,N_1565,N_1518);
or U2246 (N_2246,N_1510,N_1766);
and U2247 (N_2247,N_1861,N_1488);
nand U2248 (N_2248,N_1284,N_1483);
nand U2249 (N_2249,N_1521,N_1456);
and U2250 (N_2250,N_1764,N_1683);
and U2251 (N_2251,N_1302,N_1480);
nand U2252 (N_2252,N_1800,N_1203);
xor U2253 (N_2253,N_1167,N_1174);
and U2254 (N_2254,N_1595,N_1324);
or U2255 (N_2255,N_1797,N_1228);
or U2256 (N_2256,N_1470,N_1771);
xor U2257 (N_2257,N_1182,N_1568);
xor U2258 (N_2258,N_1768,N_1665);
and U2259 (N_2259,N_1269,N_1561);
or U2260 (N_2260,N_1969,N_1438);
and U2261 (N_2261,N_1010,N_1481);
and U2262 (N_2262,N_1204,N_1516);
xnor U2263 (N_2263,N_1465,N_1620);
or U2264 (N_2264,N_1039,N_1231);
nor U2265 (N_2265,N_1133,N_1254);
nor U2266 (N_2266,N_1927,N_1319);
xor U2267 (N_2267,N_1087,N_1557);
nor U2268 (N_2268,N_1290,N_1982);
or U2269 (N_2269,N_1712,N_1412);
and U2270 (N_2270,N_1851,N_1110);
or U2271 (N_2271,N_1241,N_1473);
nor U2272 (N_2272,N_1985,N_1567);
nand U2273 (N_2273,N_1618,N_1602);
xor U2274 (N_2274,N_1859,N_1308);
and U2275 (N_2275,N_1526,N_1866);
xnor U2276 (N_2276,N_1068,N_1770);
nor U2277 (N_2277,N_1720,N_1146);
or U2278 (N_2278,N_1046,N_1445);
and U2279 (N_2279,N_1667,N_1101);
or U2280 (N_2280,N_1358,N_1268);
or U2281 (N_2281,N_1817,N_1933);
xnor U2282 (N_2282,N_1094,N_1535);
or U2283 (N_2283,N_1736,N_1243);
nor U2284 (N_2284,N_1957,N_1171);
or U2285 (N_2285,N_1183,N_1615);
nand U2286 (N_2286,N_1682,N_1275);
and U2287 (N_2287,N_1124,N_1637);
xor U2288 (N_2288,N_1995,N_1065);
nor U2289 (N_2289,N_1702,N_1678);
nand U2290 (N_2290,N_1724,N_1198);
or U2291 (N_2291,N_1292,N_1075);
and U2292 (N_2292,N_1439,N_1812);
or U2293 (N_2293,N_1432,N_1916);
or U2294 (N_2294,N_1446,N_1788);
nand U2295 (N_2295,N_1716,N_1921);
and U2296 (N_2296,N_1937,N_1706);
nand U2297 (N_2297,N_1886,N_1673);
and U2298 (N_2298,N_1084,N_1639);
and U2299 (N_2299,N_1527,N_1636);
nor U2300 (N_2300,N_1556,N_1972);
and U2301 (N_2301,N_1865,N_1071);
nand U2302 (N_2302,N_1196,N_1577);
nand U2303 (N_2303,N_1044,N_1463);
nand U2304 (N_2304,N_1608,N_1644);
nand U2305 (N_2305,N_1472,N_1553);
xnor U2306 (N_2306,N_1448,N_1255);
and U2307 (N_2307,N_1760,N_1929);
and U2308 (N_2308,N_1536,N_1610);
xor U2309 (N_2309,N_1455,N_1904);
nand U2310 (N_2310,N_1311,N_1407);
nor U2311 (N_2311,N_1344,N_1202);
and U2312 (N_2312,N_1858,N_1988);
or U2313 (N_2313,N_1173,N_1819);
or U2314 (N_2314,N_1437,N_1327);
or U2315 (N_2315,N_1657,N_1783);
nor U2316 (N_2316,N_1949,N_1619);
and U2317 (N_2317,N_1888,N_1898);
nor U2318 (N_2318,N_1579,N_1899);
xor U2319 (N_2319,N_1440,N_1306);
xnor U2320 (N_2320,N_1547,N_1666);
and U2321 (N_2321,N_1333,N_1025);
nand U2322 (N_2322,N_1845,N_1482);
xor U2323 (N_2323,N_1538,N_1121);
xnor U2324 (N_2324,N_1550,N_1511);
or U2325 (N_2325,N_1047,N_1486);
or U2326 (N_2326,N_1250,N_1998);
nand U2327 (N_2327,N_1772,N_1134);
or U2328 (N_2328,N_1205,N_1549);
or U2329 (N_2329,N_1832,N_1279);
and U2330 (N_2330,N_1876,N_1902);
and U2331 (N_2331,N_1583,N_1316);
nor U2332 (N_2332,N_1638,N_1020);
nand U2333 (N_2333,N_1222,N_1259);
nand U2334 (N_2334,N_1107,N_1520);
or U2335 (N_2335,N_1901,N_1000);
and U2336 (N_2336,N_1464,N_1460);
nor U2337 (N_2337,N_1689,N_1992);
or U2338 (N_2338,N_1237,N_1499);
or U2339 (N_2339,N_1593,N_1409);
nand U2340 (N_2340,N_1017,N_1719);
nor U2341 (N_2341,N_1466,N_1119);
nand U2342 (N_2342,N_1375,N_1090);
or U2343 (N_2343,N_1616,N_1543);
nor U2344 (N_2344,N_1405,N_1674);
nor U2345 (N_2345,N_1594,N_1757);
xor U2346 (N_2346,N_1208,N_1863);
or U2347 (N_2347,N_1450,N_1743);
xor U2348 (N_2348,N_1162,N_1906);
nand U2349 (N_2349,N_1126,N_1836);
or U2350 (N_2350,N_1882,N_1069);
nand U2351 (N_2351,N_1611,N_1475);
xnor U2352 (N_2352,N_1038,N_1257);
or U2353 (N_2353,N_1006,N_1811);
nor U2354 (N_2354,N_1251,N_1221);
and U2355 (N_2355,N_1372,N_1398);
nand U2356 (N_2356,N_1896,N_1603);
or U2357 (N_2357,N_1855,N_1004);
and U2358 (N_2358,N_1621,N_1305);
nor U2359 (N_2359,N_1948,N_1026);
nand U2360 (N_2360,N_1960,N_1113);
or U2361 (N_2361,N_1604,N_1883);
nor U2362 (N_2362,N_1295,N_1867);
nand U2363 (N_2363,N_1007,N_1626);
or U2364 (N_2364,N_1872,N_1514);
nand U2365 (N_2365,N_1746,N_1359);
xor U2366 (N_2366,N_1946,N_1054);
and U2367 (N_2367,N_1122,N_1622);
xnor U2368 (N_2368,N_1792,N_1852);
xor U2369 (N_2369,N_1958,N_1163);
or U2370 (N_2370,N_1818,N_1264);
or U2371 (N_2371,N_1647,N_1512);
and U2372 (N_2372,N_1209,N_1245);
xnor U2373 (N_2373,N_1036,N_1118);
xor U2374 (N_2374,N_1513,N_1185);
nor U2375 (N_2375,N_1288,N_1828);
nor U2376 (N_2376,N_1753,N_1380);
and U2377 (N_2377,N_1574,N_1144);
and U2378 (N_2378,N_1166,N_1132);
xnor U2379 (N_2379,N_1165,N_1018);
nand U2380 (N_2380,N_1462,N_1945);
nor U2381 (N_2381,N_1544,N_1804);
and U2382 (N_2382,N_1326,N_1978);
and U2383 (N_2383,N_1897,N_1578);
nor U2384 (N_2384,N_1419,N_1312);
or U2385 (N_2385,N_1889,N_1145);
or U2386 (N_2386,N_1894,N_1815);
xor U2387 (N_2387,N_1931,N_1253);
nand U2388 (N_2388,N_1500,N_1885);
or U2389 (N_2389,N_1759,N_1062);
xnor U2390 (N_2390,N_1280,N_1364);
and U2391 (N_2391,N_1224,N_1941);
or U2392 (N_2392,N_1928,N_1737);
nand U2393 (N_2393,N_1791,N_1919);
nand U2394 (N_2394,N_1335,N_1627);
nand U2395 (N_2395,N_1106,N_1697);
and U2396 (N_2396,N_1704,N_1336);
nand U2397 (N_2397,N_1864,N_1955);
xnor U2398 (N_2398,N_1057,N_1519);
and U2399 (N_2399,N_1732,N_1501);
and U2400 (N_2400,N_1293,N_1586);
nand U2401 (N_2401,N_1379,N_1194);
and U2402 (N_2402,N_1905,N_1869);
nand U2403 (N_2403,N_1873,N_1154);
xor U2404 (N_2404,N_1086,N_1587);
or U2405 (N_2405,N_1216,N_1408);
or U2406 (N_2406,N_1503,N_1211);
nand U2407 (N_2407,N_1558,N_1341);
nand U2408 (N_2408,N_1981,N_1723);
and U2409 (N_2409,N_1908,N_1016);
or U2410 (N_2410,N_1959,N_1912);
or U2411 (N_2411,N_1447,N_1371);
nand U2412 (N_2412,N_1509,N_1973);
xnor U2413 (N_2413,N_1352,N_1331);
nand U2414 (N_2414,N_1307,N_1248);
and U2415 (N_2415,N_1217,N_1206);
xnor U2416 (N_2416,N_1191,N_1393);
and U2417 (N_2417,N_1907,N_1900);
and U2418 (N_2418,N_1531,N_1313);
nand U2419 (N_2419,N_1115,N_1416);
or U2420 (N_2420,N_1597,N_1748);
xor U2421 (N_2421,N_1833,N_1940);
or U2422 (N_2422,N_1999,N_1506);
nand U2423 (N_2423,N_1965,N_1997);
and U2424 (N_2424,N_1298,N_1918);
nand U2425 (N_2425,N_1696,N_1091);
nand U2426 (N_2426,N_1755,N_1260);
nor U2427 (N_2427,N_1795,N_1072);
or U2428 (N_2428,N_1944,N_1100);
nand U2429 (N_2429,N_1425,N_1415);
and U2430 (N_2430,N_1028,N_1829);
or U2431 (N_2431,N_1471,N_1827);
or U2432 (N_2432,N_1645,N_1112);
xnor U2433 (N_2433,N_1226,N_1920);
xnor U2434 (N_2434,N_1569,N_1642);
or U2435 (N_2435,N_1030,N_1767);
or U2436 (N_2436,N_1848,N_1868);
or U2437 (N_2437,N_1219,N_1910);
xnor U2438 (N_2438,N_1887,N_1877);
or U2439 (N_2439,N_1041,N_1694);
xnor U2440 (N_2440,N_1034,N_1077);
nor U2441 (N_2441,N_1468,N_1713);
nor U2442 (N_2442,N_1687,N_1067);
xor U2443 (N_2443,N_1052,N_1366);
and U2444 (N_2444,N_1573,N_1742);
or U2445 (N_2445,N_1730,N_1186);
xnor U2446 (N_2446,N_1332,N_1623);
and U2447 (N_2447,N_1078,N_1055);
nor U2448 (N_2448,N_1299,N_1021);
nor U2449 (N_2449,N_1686,N_1097);
nor U2450 (N_2450,N_1382,N_1975);
or U2451 (N_2451,N_1703,N_1428);
or U2452 (N_2452,N_1653,N_1452);
and U2453 (N_2453,N_1805,N_1925);
nor U2454 (N_2454,N_1794,N_1161);
and U2455 (N_2455,N_1589,N_1559);
xnor U2456 (N_2456,N_1287,N_1562);
and U2457 (N_2457,N_1207,N_1457);
or U2458 (N_2458,N_1008,N_1402);
nand U2459 (N_2459,N_1190,N_1530);
nand U2460 (N_2460,N_1563,N_1854);
nand U2461 (N_2461,N_1914,N_1909);
and U2462 (N_2462,N_1821,N_1630);
nand U2463 (N_2463,N_1793,N_1962);
or U2464 (N_2464,N_1433,N_1576);
and U2465 (N_2465,N_1707,N_1675);
or U2466 (N_2466,N_1786,N_1849);
nor U2467 (N_2467,N_1935,N_1012);
xor U2468 (N_2468,N_1745,N_1655);
or U2469 (N_2469,N_1695,N_1953);
nand U2470 (N_2470,N_1318,N_1974);
or U2471 (N_2471,N_1523,N_1349);
nand U2472 (N_2472,N_1252,N_1691);
and U2473 (N_2473,N_1533,N_1043);
nand U2474 (N_2474,N_1599,N_1984);
or U2475 (N_2475,N_1986,N_1345);
nand U2476 (N_2476,N_1225,N_1507);
xnor U2477 (N_2477,N_1449,N_1164);
xnor U2478 (N_2478,N_1160,N_1066);
and U2479 (N_2479,N_1903,N_1663);
or U2480 (N_2480,N_1725,N_1152);
nand U2481 (N_2481,N_1991,N_1244);
xor U2482 (N_2482,N_1525,N_1971);
or U2483 (N_2483,N_1605,N_1404);
nor U2484 (N_2484,N_1321,N_1672);
nor U2485 (N_2485,N_1155,N_1142);
nand U2486 (N_2486,N_1418,N_1661);
and U2487 (N_2487,N_1289,N_1361);
and U2488 (N_2488,N_1291,N_1303);
nor U2489 (N_2489,N_1430,N_1147);
and U2490 (N_2490,N_1201,N_1491);
or U2491 (N_2491,N_1104,N_1609);
nand U2492 (N_2492,N_1934,N_1187);
or U2493 (N_2493,N_1504,N_1502);
nand U2494 (N_2494,N_1467,N_1803);
and U2495 (N_2495,N_1357,N_1197);
nor U2496 (N_2496,N_1002,N_1153);
and U2497 (N_2497,N_1496,N_1265);
or U2498 (N_2498,N_1140,N_1235);
xor U2499 (N_2499,N_1003,N_1281);
nor U2500 (N_2500,N_1520,N_1983);
nor U2501 (N_2501,N_1413,N_1392);
nor U2502 (N_2502,N_1625,N_1639);
xnor U2503 (N_2503,N_1233,N_1821);
or U2504 (N_2504,N_1701,N_1666);
or U2505 (N_2505,N_1020,N_1045);
and U2506 (N_2506,N_1593,N_1115);
and U2507 (N_2507,N_1909,N_1898);
or U2508 (N_2508,N_1773,N_1474);
or U2509 (N_2509,N_1159,N_1158);
and U2510 (N_2510,N_1409,N_1089);
and U2511 (N_2511,N_1086,N_1453);
nor U2512 (N_2512,N_1016,N_1441);
and U2513 (N_2513,N_1270,N_1617);
nand U2514 (N_2514,N_1286,N_1960);
and U2515 (N_2515,N_1207,N_1833);
and U2516 (N_2516,N_1804,N_1032);
and U2517 (N_2517,N_1973,N_1978);
nor U2518 (N_2518,N_1065,N_1034);
xnor U2519 (N_2519,N_1930,N_1800);
or U2520 (N_2520,N_1881,N_1846);
and U2521 (N_2521,N_1759,N_1050);
nor U2522 (N_2522,N_1356,N_1438);
nor U2523 (N_2523,N_1542,N_1225);
and U2524 (N_2524,N_1205,N_1391);
nand U2525 (N_2525,N_1255,N_1534);
xnor U2526 (N_2526,N_1868,N_1242);
and U2527 (N_2527,N_1313,N_1912);
nand U2528 (N_2528,N_1059,N_1276);
xnor U2529 (N_2529,N_1635,N_1678);
xor U2530 (N_2530,N_1399,N_1422);
or U2531 (N_2531,N_1863,N_1801);
and U2532 (N_2532,N_1382,N_1220);
nor U2533 (N_2533,N_1325,N_1627);
nor U2534 (N_2534,N_1859,N_1884);
xnor U2535 (N_2535,N_1610,N_1185);
xnor U2536 (N_2536,N_1532,N_1886);
or U2537 (N_2537,N_1819,N_1304);
xor U2538 (N_2538,N_1564,N_1873);
xnor U2539 (N_2539,N_1375,N_1264);
nand U2540 (N_2540,N_1670,N_1586);
nand U2541 (N_2541,N_1815,N_1434);
and U2542 (N_2542,N_1309,N_1972);
xor U2543 (N_2543,N_1498,N_1581);
and U2544 (N_2544,N_1936,N_1086);
nand U2545 (N_2545,N_1939,N_1126);
and U2546 (N_2546,N_1354,N_1522);
nand U2547 (N_2547,N_1593,N_1073);
or U2548 (N_2548,N_1565,N_1696);
nor U2549 (N_2549,N_1112,N_1044);
nand U2550 (N_2550,N_1045,N_1493);
nor U2551 (N_2551,N_1460,N_1722);
xor U2552 (N_2552,N_1259,N_1568);
or U2553 (N_2553,N_1433,N_1232);
or U2554 (N_2554,N_1616,N_1887);
xor U2555 (N_2555,N_1058,N_1126);
nor U2556 (N_2556,N_1187,N_1108);
nand U2557 (N_2557,N_1807,N_1405);
nand U2558 (N_2558,N_1000,N_1146);
and U2559 (N_2559,N_1885,N_1575);
xor U2560 (N_2560,N_1538,N_1920);
nand U2561 (N_2561,N_1912,N_1906);
nor U2562 (N_2562,N_1560,N_1020);
nand U2563 (N_2563,N_1726,N_1011);
nand U2564 (N_2564,N_1345,N_1475);
or U2565 (N_2565,N_1136,N_1753);
nor U2566 (N_2566,N_1240,N_1524);
nor U2567 (N_2567,N_1896,N_1147);
nor U2568 (N_2568,N_1042,N_1317);
nand U2569 (N_2569,N_1611,N_1074);
nor U2570 (N_2570,N_1079,N_1548);
nand U2571 (N_2571,N_1053,N_1096);
xor U2572 (N_2572,N_1779,N_1591);
or U2573 (N_2573,N_1596,N_1923);
or U2574 (N_2574,N_1530,N_1000);
and U2575 (N_2575,N_1644,N_1351);
or U2576 (N_2576,N_1069,N_1745);
xnor U2577 (N_2577,N_1214,N_1218);
and U2578 (N_2578,N_1040,N_1773);
or U2579 (N_2579,N_1631,N_1953);
and U2580 (N_2580,N_1059,N_1111);
and U2581 (N_2581,N_1575,N_1529);
and U2582 (N_2582,N_1535,N_1796);
xor U2583 (N_2583,N_1078,N_1777);
or U2584 (N_2584,N_1812,N_1925);
nor U2585 (N_2585,N_1653,N_1677);
nor U2586 (N_2586,N_1553,N_1559);
nor U2587 (N_2587,N_1228,N_1350);
or U2588 (N_2588,N_1595,N_1006);
nand U2589 (N_2589,N_1877,N_1424);
nand U2590 (N_2590,N_1011,N_1779);
or U2591 (N_2591,N_1078,N_1386);
xor U2592 (N_2592,N_1526,N_1814);
nand U2593 (N_2593,N_1817,N_1382);
xnor U2594 (N_2594,N_1561,N_1348);
nand U2595 (N_2595,N_1013,N_1192);
and U2596 (N_2596,N_1899,N_1606);
and U2597 (N_2597,N_1126,N_1652);
or U2598 (N_2598,N_1094,N_1755);
nand U2599 (N_2599,N_1743,N_1988);
or U2600 (N_2600,N_1245,N_1098);
or U2601 (N_2601,N_1939,N_1893);
xor U2602 (N_2602,N_1977,N_1461);
or U2603 (N_2603,N_1731,N_1061);
and U2604 (N_2604,N_1366,N_1814);
xor U2605 (N_2605,N_1364,N_1179);
nand U2606 (N_2606,N_1472,N_1424);
nor U2607 (N_2607,N_1418,N_1451);
and U2608 (N_2608,N_1658,N_1848);
nand U2609 (N_2609,N_1620,N_1028);
nand U2610 (N_2610,N_1082,N_1984);
nor U2611 (N_2611,N_1694,N_1467);
or U2612 (N_2612,N_1869,N_1406);
nand U2613 (N_2613,N_1973,N_1724);
nand U2614 (N_2614,N_1802,N_1725);
or U2615 (N_2615,N_1667,N_1451);
and U2616 (N_2616,N_1425,N_1103);
xnor U2617 (N_2617,N_1023,N_1119);
nor U2618 (N_2618,N_1714,N_1481);
nor U2619 (N_2619,N_1893,N_1847);
or U2620 (N_2620,N_1001,N_1033);
and U2621 (N_2621,N_1747,N_1511);
nand U2622 (N_2622,N_1918,N_1052);
and U2623 (N_2623,N_1721,N_1427);
and U2624 (N_2624,N_1601,N_1716);
nor U2625 (N_2625,N_1674,N_1491);
and U2626 (N_2626,N_1483,N_1091);
or U2627 (N_2627,N_1697,N_1223);
nand U2628 (N_2628,N_1713,N_1539);
or U2629 (N_2629,N_1327,N_1816);
or U2630 (N_2630,N_1357,N_1437);
xnor U2631 (N_2631,N_1805,N_1286);
nor U2632 (N_2632,N_1015,N_1844);
nor U2633 (N_2633,N_1866,N_1666);
xnor U2634 (N_2634,N_1048,N_1868);
nor U2635 (N_2635,N_1878,N_1388);
or U2636 (N_2636,N_1697,N_1896);
xnor U2637 (N_2637,N_1784,N_1293);
nor U2638 (N_2638,N_1288,N_1462);
nand U2639 (N_2639,N_1689,N_1714);
and U2640 (N_2640,N_1215,N_1250);
nand U2641 (N_2641,N_1608,N_1231);
nor U2642 (N_2642,N_1908,N_1192);
or U2643 (N_2643,N_1207,N_1943);
nor U2644 (N_2644,N_1094,N_1104);
xor U2645 (N_2645,N_1813,N_1261);
and U2646 (N_2646,N_1576,N_1922);
nand U2647 (N_2647,N_1793,N_1728);
nor U2648 (N_2648,N_1139,N_1768);
and U2649 (N_2649,N_1318,N_1054);
and U2650 (N_2650,N_1143,N_1505);
nor U2651 (N_2651,N_1337,N_1326);
nor U2652 (N_2652,N_1599,N_1516);
and U2653 (N_2653,N_1050,N_1564);
xor U2654 (N_2654,N_1023,N_1033);
xor U2655 (N_2655,N_1296,N_1837);
nor U2656 (N_2656,N_1694,N_1676);
or U2657 (N_2657,N_1141,N_1960);
xor U2658 (N_2658,N_1143,N_1868);
xnor U2659 (N_2659,N_1173,N_1969);
or U2660 (N_2660,N_1632,N_1865);
and U2661 (N_2661,N_1136,N_1795);
nand U2662 (N_2662,N_1046,N_1045);
and U2663 (N_2663,N_1377,N_1793);
nor U2664 (N_2664,N_1074,N_1885);
and U2665 (N_2665,N_1553,N_1988);
nor U2666 (N_2666,N_1862,N_1635);
xnor U2667 (N_2667,N_1041,N_1584);
xnor U2668 (N_2668,N_1085,N_1451);
xnor U2669 (N_2669,N_1560,N_1732);
or U2670 (N_2670,N_1475,N_1389);
xor U2671 (N_2671,N_1620,N_1656);
xor U2672 (N_2672,N_1327,N_1649);
and U2673 (N_2673,N_1805,N_1547);
nor U2674 (N_2674,N_1375,N_1910);
nand U2675 (N_2675,N_1107,N_1657);
and U2676 (N_2676,N_1575,N_1071);
xnor U2677 (N_2677,N_1982,N_1713);
nand U2678 (N_2678,N_1795,N_1459);
xnor U2679 (N_2679,N_1987,N_1996);
or U2680 (N_2680,N_1324,N_1691);
and U2681 (N_2681,N_1400,N_1157);
nand U2682 (N_2682,N_1687,N_1953);
or U2683 (N_2683,N_1836,N_1020);
and U2684 (N_2684,N_1047,N_1503);
nand U2685 (N_2685,N_1568,N_1056);
xor U2686 (N_2686,N_1435,N_1518);
xnor U2687 (N_2687,N_1650,N_1922);
and U2688 (N_2688,N_1479,N_1003);
nand U2689 (N_2689,N_1923,N_1543);
and U2690 (N_2690,N_1574,N_1165);
nand U2691 (N_2691,N_1551,N_1458);
and U2692 (N_2692,N_1942,N_1254);
or U2693 (N_2693,N_1141,N_1925);
xnor U2694 (N_2694,N_1098,N_1271);
and U2695 (N_2695,N_1214,N_1706);
xnor U2696 (N_2696,N_1925,N_1789);
nor U2697 (N_2697,N_1782,N_1139);
nand U2698 (N_2698,N_1915,N_1462);
nor U2699 (N_2699,N_1654,N_1374);
and U2700 (N_2700,N_1206,N_1761);
and U2701 (N_2701,N_1578,N_1196);
or U2702 (N_2702,N_1555,N_1029);
and U2703 (N_2703,N_1587,N_1844);
xnor U2704 (N_2704,N_1585,N_1914);
and U2705 (N_2705,N_1953,N_1343);
or U2706 (N_2706,N_1596,N_1709);
or U2707 (N_2707,N_1376,N_1129);
and U2708 (N_2708,N_1182,N_1051);
xnor U2709 (N_2709,N_1111,N_1854);
xor U2710 (N_2710,N_1812,N_1289);
or U2711 (N_2711,N_1920,N_1430);
or U2712 (N_2712,N_1619,N_1136);
or U2713 (N_2713,N_1869,N_1795);
or U2714 (N_2714,N_1336,N_1082);
or U2715 (N_2715,N_1045,N_1812);
nand U2716 (N_2716,N_1794,N_1590);
and U2717 (N_2717,N_1162,N_1585);
xnor U2718 (N_2718,N_1510,N_1516);
nor U2719 (N_2719,N_1509,N_1395);
and U2720 (N_2720,N_1065,N_1352);
xnor U2721 (N_2721,N_1961,N_1666);
and U2722 (N_2722,N_1961,N_1673);
and U2723 (N_2723,N_1842,N_1188);
or U2724 (N_2724,N_1287,N_1714);
nand U2725 (N_2725,N_1772,N_1356);
or U2726 (N_2726,N_1234,N_1428);
xor U2727 (N_2727,N_1147,N_1159);
or U2728 (N_2728,N_1666,N_1587);
or U2729 (N_2729,N_1335,N_1254);
nand U2730 (N_2730,N_1308,N_1814);
nand U2731 (N_2731,N_1490,N_1289);
nand U2732 (N_2732,N_1508,N_1110);
nor U2733 (N_2733,N_1862,N_1633);
and U2734 (N_2734,N_1624,N_1728);
xor U2735 (N_2735,N_1514,N_1196);
or U2736 (N_2736,N_1337,N_1440);
or U2737 (N_2737,N_1905,N_1233);
nor U2738 (N_2738,N_1404,N_1984);
xnor U2739 (N_2739,N_1945,N_1864);
xnor U2740 (N_2740,N_1111,N_1771);
and U2741 (N_2741,N_1667,N_1481);
and U2742 (N_2742,N_1585,N_1408);
nor U2743 (N_2743,N_1339,N_1487);
nor U2744 (N_2744,N_1343,N_1742);
or U2745 (N_2745,N_1542,N_1555);
and U2746 (N_2746,N_1219,N_1101);
and U2747 (N_2747,N_1990,N_1229);
nor U2748 (N_2748,N_1735,N_1056);
xor U2749 (N_2749,N_1385,N_1474);
nand U2750 (N_2750,N_1565,N_1759);
xor U2751 (N_2751,N_1110,N_1895);
and U2752 (N_2752,N_1126,N_1805);
and U2753 (N_2753,N_1147,N_1764);
nor U2754 (N_2754,N_1320,N_1324);
or U2755 (N_2755,N_1956,N_1928);
xnor U2756 (N_2756,N_1137,N_1773);
nor U2757 (N_2757,N_1494,N_1055);
xor U2758 (N_2758,N_1721,N_1886);
nand U2759 (N_2759,N_1134,N_1826);
xor U2760 (N_2760,N_1586,N_1537);
or U2761 (N_2761,N_1181,N_1893);
or U2762 (N_2762,N_1350,N_1998);
nor U2763 (N_2763,N_1619,N_1142);
nor U2764 (N_2764,N_1872,N_1866);
or U2765 (N_2765,N_1152,N_1761);
or U2766 (N_2766,N_1847,N_1989);
or U2767 (N_2767,N_1637,N_1075);
xnor U2768 (N_2768,N_1424,N_1997);
xnor U2769 (N_2769,N_1860,N_1244);
nand U2770 (N_2770,N_1763,N_1775);
nand U2771 (N_2771,N_1197,N_1119);
or U2772 (N_2772,N_1448,N_1784);
nand U2773 (N_2773,N_1790,N_1156);
nand U2774 (N_2774,N_1501,N_1664);
or U2775 (N_2775,N_1815,N_1431);
nand U2776 (N_2776,N_1400,N_1803);
xnor U2777 (N_2777,N_1669,N_1633);
nor U2778 (N_2778,N_1645,N_1840);
xor U2779 (N_2779,N_1162,N_1243);
nand U2780 (N_2780,N_1950,N_1952);
and U2781 (N_2781,N_1489,N_1199);
nor U2782 (N_2782,N_1643,N_1927);
or U2783 (N_2783,N_1006,N_1745);
nor U2784 (N_2784,N_1593,N_1424);
and U2785 (N_2785,N_1872,N_1850);
or U2786 (N_2786,N_1619,N_1751);
nand U2787 (N_2787,N_1891,N_1472);
or U2788 (N_2788,N_1836,N_1622);
or U2789 (N_2789,N_1886,N_1473);
xnor U2790 (N_2790,N_1825,N_1612);
or U2791 (N_2791,N_1828,N_1661);
or U2792 (N_2792,N_1530,N_1261);
xor U2793 (N_2793,N_1357,N_1251);
and U2794 (N_2794,N_1046,N_1814);
nor U2795 (N_2795,N_1903,N_1747);
and U2796 (N_2796,N_1301,N_1560);
and U2797 (N_2797,N_1867,N_1948);
xor U2798 (N_2798,N_1461,N_1729);
nand U2799 (N_2799,N_1242,N_1018);
and U2800 (N_2800,N_1654,N_1746);
and U2801 (N_2801,N_1664,N_1884);
nand U2802 (N_2802,N_1986,N_1135);
and U2803 (N_2803,N_1974,N_1600);
xor U2804 (N_2804,N_1742,N_1494);
nand U2805 (N_2805,N_1729,N_1051);
xnor U2806 (N_2806,N_1389,N_1983);
nand U2807 (N_2807,N_1945,N_1333);
xor U2808 (N_2808,N_1367,N_1018);
and U2809 (N_2809,N_1273,N_1890);
nor U2810 (N_2810,N_1400,N_1196);
nor U2811 (N_2811,N_1082,N_1949);
and U2812 (N_2812,N_1768,N_1391);
xor U2813 (N_2813,N_1591,N_1023);
or U2814 (N_2814,N_1392,N_1925);
and U2815 (N_2815,N_1981,N_1835);
nand U2816 (N_2816,N_1713,N_1347);
nor U2817 (N_2817,N_1090,N_1570);
xnor U2818 (N_2818,N_1038,N_1503);
xnor U2819 (N_2819,N_1187,N_1295);
and U2820 (N_2820,N_1321,N_1647);
and U2821 (N_2821,N_1988,N_1944);
or U2822 (N_2822,N_1969,N_1792);
and U2823 (N_2823,N_1385,N_1037);
and U2824 (N_2824,N_1880,N_1396);
nand U2825 (N_2825,N_1143,N_1817);
or U2826 (N_2826,N_1519,N_1701);
or U2827 (N_2827,N_1522,N_1693);
xnor U2828 (N_2828,N_1626,N_1106);
and U2829 (N_2829,N_1490,N_1458);
and U2830 (N_2830,N_1331,N_1743);
and U2831 (N_2831,N_1669,N_1603);
or U2832 (N_2832,N_1890,N_1656);
and U2833 (N_2833,N_1682,N_1906);
and U2834 (N_2834,N_1126,N_1286);
and U2835 (N_2835,N_1560,N_1627);
xor U2836 (N_2836,N_1835,N_1342);
nand U2837 (N_2837,N_1433,N_1208);
or U2838 (N_2838,N_1722,N_1173);
and U2839 (N_2839,N_1063,N_1478);
xor U2840 (N_2840,N_1987,N_1242);
nor U2841 (N_2841,N_1554,N_1807);
nor U2842 (N_2842,N_1737,N_1673);
and U2843 (N_2843,N_1202,N_1164);
nor U2844 (N_2844,N_1703,N_1344);
xnor U2845 (N_2845,N_1512,N_1490);
and U2846 (N_2846,N_1308,N_1377);
or U2847 (N_2847,N_1154,N_1217);
or U2848 (N_2848,N_1148,N_1214);
or U2849 (N_2849,N_1795,N_1309);
nor U2850 (N_2850,N_1512,N_1768);
or U2851 (N_2851,N_1988,N_1855);
xnor U2852 (N_2852,N_1485,N_1573);
nor U2853 (N_2853,N_1870,N_1143);
or U2854 (N_2854,N_1881,N_1629);
or U2855 (N_2855,N_1008,N_1795);
xnor U2856 (N_2856,N_1678,N_1624);
and U2857 (N_2857,N_1264,N_1056);
xnor U2858 (N_2858,N_1493,N_1236);
xnor U2859 (N_2859,N_1959,N_1257);
xor U2860 (N_2860,N_1758,N_1781);
and U2861 (N_2861,N_1285,N_1262);
nand U2862 (N_2862,N_1203,N_1378);
xnor U2863 (N_2863,N_1930,N_1688);
or U2864 (N_2864,N_1971,N_1020);
nand U2865 (N_2865,N_1695,N_1298);
or U2866 (N_2866,N_1112,N_1439);
or U2867 (N_2867,N_1318,N_1891);
or U2868 (N_2868,N_1476,N_1226);
and U2869 (N_2869,N_1282,N_1892);
nand U2870 (N_2870,N_1878,N_1835);
nand U2871 (N_2871,N_1679,N_1991);
or U2872 (N_2872,N_1040,N_1841);
or U2873 (N_2873,N_1053,N_1846);
and U2874 (N_2874,N_1436,N_1238);
nand U2875 (N_2875,N_1647,N_1690);
nand U2876 (N_2876,N_1482,N_1598);
nor U2877 (N_2877,N_1151,N_1486);
and U2878 (N_2878,N_1822,N_1493);
xnor U2879 (N_2879,N_1357,N_1393);
nand U2880 (N_2880,N_1657,N_1558);
and U2881 (N_2881,N_1969,N_1362);
nor U2882 (N_2882,N_1174,N_1289);
nor U2883 (N_2883,N_1474,N_1188);
xnor U2884 (N_2884,N_1093,N_1819);
xor U2885 (N_2885,N_1417,N_1248);
xor U2886 (N_2886,N_1611,N_1604);
and U2887 (N_2887,N_1001,N_1160);
nand U2888 (N_2888,N_1269,N_1746);
and U2889 (N_2889,N_1762,N_1898);
or U2890 (N_2890,N_1424,N_1731);
nand U2891 (N_2891,N_1797,N_1278);
nand U2892 (N_2892,N_1210,N_1660);
xnor U2893 (N_2893,N_1279,N_1083);
nor U2894 (N_2894,N_1751,N_1758);
xor U2895 (N_2895,N_1653,N_1740);
nor U2896 (N_2896,N_1449,N_1452);
nor U2897 (N_2897,N_1855,N_1920);
or U2898 (N_2898,N_1109,N_1879);
or U2899 (N_2899,N_1677,N_1042);
xor U2900 (N_2900,N_1324,N_1803);
and U2901 (N_2901,N_1713,N_1205);
and U2902 (N_2902,N_1962,N_1602);
xor U2903 (N_2903,N_1165,N_1281);
nor U2904 (N_2904,N_1788,N_1932);
nand U2905 (N_2905,N_1869,N_1193);
nor U2906 (N_2906,N_1330,N_1608);
and U2907 (N_2907,N_1530,N_1046);
xnor U2908 (N_2908,N_1002,N_1068);
or U2909 (N_2909,N_1545,N_1634);
xor U2910 (N_2910,N_1345,N_1224);
nand U2911 (N_2911,N_1185,N_1337);
nor U2912 (N_2912,N_1281,N_1592);
and U2913 (N_2913,N_1279,N_1922);
xnor U2914 (N_2914,N_1578,N_1321);
or U2915 (N_2915,N_1082,N_1773);
or U2916 (N_2916,N_1143,N_1880);
and U2917 (N_2917,N_1543,N_1200);
nand U2918 (N_2918,N_1005,N_1406);
xnor U2919 (N_2919,N_1648,N_1233);
xnor U2920 (N_2920,N_1600,N_1063);
nand U2921 (N_2921,N_1023,N_1711);
or U2922 (N_2922,N_1532,N_1029);
and U2923 (N_2923,N_1979,N_1673);
xnor U2924 (N_2924,N_1712,N_1341);
xnor U2925 (N_2925,N_1577,N_1687);
or U2926 (N_2926,N_1571,N_1225);
nor U2927 (N_2927,N_1817,N_1061);
or U2928 (N_2928,N_1802,N_1654);
and U2929 (N_2929,N_1522,N_1077);
nand U2930 (N_2930,N_1026,N_1598);
or U2931 (N_2931,N_1052,N_1299);
nand U2932 (N_2932,N_1159,N_1374);
nor U2933 (N_2933,N_1551,N_1397);
and U2934 (N_2934,N_1572,N_1725);
and U2935 (N_2935,N_1238,N_1513);
and U2936 (N_2936,N_1377,N_1695);
nor U2937 (N_2937,N_1386,N_1340);
and U2938 (N_2938,N_1137,N_1558);
and U2939 (N_2939,N_1085,N_1179);
nand U2940 (N_2940,N_1285,N_1573);
and U2941 (N_2941,N_1027,N_1026);
xnor U2942 (N_2942,N_1483,N_1395);
or U2943 (N_2943,N_1388,N_1271);
and U2944 (N_2944,N_1956,N_1677);
and U2945 (N_2945,N_1602,N_1719);
and U2946 (N_2946,N_1147,N_1585);
or U2947 (N_2947,N_1158,N_1333);
xor U2948 (N_2948,N_1182,N_1716);
and U2949 (N_2949,N_1558,N_1874);
nand U2950 (N_2950,N_1394,N_1733);
xor U2951 (N_2951,N_1368,N_1035);
and U2952 (N_2952,N_1823,N_1970);
nor U2953 (N_2953,N_1052,N_1587);
xnor U2954 (N_2954,N_1094,N_1462);
nor U2955 (N_2955,N_1586,N_1591);
or U2956 (N_2956,N_1203,N_1380);
and U2957 (N_2957,N_1968,N_1494);
xor U2958 (N_2958,N_1349,N_1632);
nand U2959 (N_2959,N_1146,N_1426);
xor U2960 (N_2960,N_1827,N_1243);
nor U2961 (N_2961,N_1691,N_1479);
nor U2962 (N_2962,N_1877,N_1063);
nor U2963 (N_2963,N_1036,N_1555);
or U2964 (N_2964,N_1446,N_1128);
or U2965 (N_2965,N_1026,N_1513);
or U2966 (N_2966,N_1131,N_1895);
or U2967 (N_2967,N_1358,N_1742);
nand U2968 (N_2968,N_1026,N_1190);
nand U2969 (N_2969,N_1583,N_1417);
nor U2970 (N_2970,N_1930,N_1837);
nand U2971 (N_2971,N_1028,N_1294);
or U2972 (N_2972,N_1039,N_1467);
or U2973 (N_2973,N_1720,N_1361);
nor U2974 (N_2974,N_1124,N_1270);
or U2975 (N_2975,N_1758,N_1952);
nand U2976 (N_2976,N_1402,N_1637);
nand U2977 (N_2977,N_1827,N_1874);
xor U2978 (N_2978,N_1015,N_1948);
xor U2979 (N_2979,N_1374,N_1635);
xor U2980 (N_2980,N_1172,N_1540);
nand U2981 (N_2981,N_1866,N_1685);
xnor U2982 (N_2982,N_1149,N_1615);
and U2983 (N_2983,N_1494,N_1045);
and U2984 (N_2984,N_1629,N_1826);
xnor U2985 (N_2985,N_1291,N_1212);
nand U2986 (N_2986,N_1719,N_1775);
or U2987 (N_2987,N_1648,N_1490);
or U2988 (N_2988,N_1120,N_1237);
or U2989 (N_2989,N_1927,N_1380);
and U2990 (N_2990,N_1142,N_1267);
nand U2991 (N_2991,N_1605,N_1333);
xnor U2992 (N_2992,N_1295,N_1950);
nand U2993 (N_2993,N_1486,N_1301);
xnor U2994 (N_2994,N_1562,N_1768);
xor U2995 (N_2995,N_1437,N_1288);
and U2996 (N_2996,N_1111,N_1775);
nand U2997 (N_2997,N_1236,N_1270);
and U2998 (N_2998,N_1458,N_1806);
or U2999 (N_2999,N_1664,N_1892);
xor U3000 (N_3000,N_2640,N_2677);
nand U3001 (N_3001,N_2723,N_2029);
nor U3002 (N_3002,N_2061,N_2241);
nor U3003 (N_3003,N_2831,N_2216);
xnor U3004 (N_3004,N_2433,N_2016);
nor U3005 (N_3005,N_2945,N_2778);
and U3006 (N_3006,N_2467,N_2396);
and U3007 (N_3007,N_2857,N_2953);
and U3008 (N_3008,N_2874,N_2887);
nand U3009 (N_3009,N_2878,N_2611);
xor U3010 (N_3010,N_2872,N_2641);
nor U3011 (N_3011,N_2686,N_2163);
or U3012 (N_3012,N_2576,N_2375);
xor U3013 (N_3013,N_2646,N_2757);
xor U3014 (N_3014,N_2080,N_2420);
nand U3015 (N_3015,N_2924,N_2739);
or U3016 (N_3016,N_2367,N_2803);
nor U3017 (N_3017,N_2028,N_2973);
nand U3018 (N_3018,N_2620,N_2910);
nand U3019 (N_3019,N_2208,N_2868);
and U3020 (N_3020,N_2115,N_2227);
and U3021 (N_3021,N_2372,N_2344);
or U3022 (N_3022,N_2161,N_2599);
nor U3023 (N_3023,N_2993,N_2896);
nand U3024 (N_3024,N_2350,N_2383);
nand U3025 (N_3025,N_2410,N_2880);
xor U3026 (N_3026,N_2533,N_2962);
and U3027 (N_3027,N_2624,N_2477);
nand U3028 (N_3028,N_2837,N_2829);
nor U3029 (N_3029,N_2863,N_2370);
or U3030 (N_3030,N_2499,N_2283);
or U3031 (N_3031,N_2230,N_2716);
xnor U3032 (N_3032,N_2675,N_2135);
xor U3033 (N_3033,N_2510,N_2722);
xor U3034 (N_3034,N_2751,N_2264);
xor U3035 (N_3035,N_2813,N_2101);
nor U3036 (N_3036,N_2219,N_2622);
or U3037 (N_3037,N_2472,N_2178);
nor U3038 (N_3038,N_2685,N_2545);
nand U3039 (N_3039,N_2743,N_2421);
nor U3040 (N_3040,N_2681,N_2475);
and U3041 (N_3041,N_2205,N_2489);
nand U3042 (N_3042,N_2218,N_2112);
xor U3043 (N_3043,N_2428,N_2939);
nor U3044 (N_3044,N_2592,N_2495);
xnor U3045 (N_3045,N_2690,N_2667);
nor U3046 (N_3046,N_2921,N_2360);
nand U3047 (N_3047,N_2144,N_2278);
xnor U3048 (N_3048,N_2182,N_2940);
xor U3049 (N_3049,N_2904,N_2736);
nand U3050 (N_3050,N_2177,N_2676);
nand U3051 (N_3051,N_2267,N_2563);
and U3052 (N_3052,N_2152,N_2326);
and U3053 (N_3053,N_2578,N_2132);
nor U3054 (N_3054,N_2379,N_2341);
or U3055 (N_3055,N_2330,N_2537);
nor U3056 (N_3056,N_2765,N_2565);
nor U3057 (N_3057,N_2167,N_2405);
or U3058 (N_3058,N_2170,N_2842);
or U3059 (N_3059,N_2562,N_2998);
or U3060 (N_3060,N_2841,N_2927);
xnor U3061 (N_3061,N_2884,N_2965);
xnor U3062 (N_3062,N_2391,N_2388);
and U3063 (N_3063,N_2631,N_2932);
nand U3064 (N_3064,N_2046,N_2791);
nor U3065 (N_3065,N_2120,N_2859);
xor U3066 (N_3066,N_2542,N_2465);
nand U3067 (N_3067,N_2134,N_2756);
or U3068 (N_3068,N_2990,N_2610);
or U3069 (N_3069,N_2256,N_2529);
xor U3070 (N_3070,N_2777,N_2853);
xor U3071 (N_3071,N_2892,N_2009);
or U3072 (N_3072,N_2678,N_2030);
or U3073 (N_3073,N_2301,N_2649);
nand U3074 (N_3074,N_2509,N_2710);
nand U3075 (N_3075,N_2065,N_2325);
and U3076 (N_3076,N_2987,N_2110);
or U3077 (N_3077,N_2508,N_2732);
nor U3078 (N_3078,N_2642,N_2556);
nor U3079 (N_3079,N_2770,N_2655);
and U3080 (N_3080,N_2126,N_2031);
nand U3081 (N_3081,N_2225,N_2012);
and U3082 (N_3082,N_2005,N_2176);
or U3083 (N_3083,N_2385,N_2106);
xor U3084 (N_3084,N_2458,N_2724);
and U3085 (N_3085,N_2543,N_2483);
or U3086 (N_3086,N_2520,N_2203);
nor U3087 (N_3087,N_2395,N_2362);
or U3088 (N_3088,N_2586,N_2306);
and U3089 (N_3089,N_2334,N_2290);
xnor U3090 (N_3090,N_2077,N_2915);
nand U3091 (N_3091,N_2625,N_2279);
and U3092 (N_3092,N_2527,N_2574);
nand U3093 (N_3093,N_2022,N_2053);
and U3094 (N_3094,N_2984,N_2960);
nor U3095 (N_3095,N_2528,N_2389);
and U3096 (N_3096,N_2930,N_2036);
xnor U3097 (N_3097,N_2839,N_2346);
nand U3098 (N_3098,N_2522,N_2222);
nand U3099 (N_3099,N_2013,N_2840);
or U3100 (N_3100,N_2011,N_2081);
or U3101 (N_3101,N_2503,N_2616);
nor U3102 (N_3102,N_2828,N_2551);
nand U3103 (N_3103,N_2913,N_2179);
or U3104 (N_3104,N_2619,N_2038);
or U3105 (N_3105,N_2213,N_2003);
or U3106 (N_3106,N_2986,N_2727);
nor U3107 (N_3107,N_2902,N_2974);
or U3108 (N_3108,N_2844,N_2284);
or U3109 (N_3109,N_2571,N_2714);
and U3110 (N_3110,N_2443,N_2800);
nand U3111 (N_3111,N_2014,N_2358);
nand U3112 (N_3112,N_2249,N_2246);
xor U3113 (N_3113,N_2444,N_2183);
or U3114 (N_3114,N_2487,N_2501);
nor U3115 (N_3115,N_2607,N_2122);
nor U3116 (N_3116,N_2833,N_2351);
xor U3117 (N_3117,N_2459,N_2972);
xnor U3118 (N_3118,N_2700,N_2816);
nor U3119 (N_3119,N_2398,N_2426);
nand U3120 (N_3120,N_2039,N_2174);
nor U3121 (N_3121,N_2266,N_2790);
xor U3122 (N_3122,N_2253,N_2883);
nor U3123 (N_3123,N_2867,N_2804);
nand U3124 (N_3124,N_2713,N_2779);
xor U3125 (N_3125,N_2149,N_2357);
nor U3126 (N_3126,N_2125,N_2672);
nand U3127 (N_3127,N_2289,N_2068);
nor U3128 (N_3128,N_2796,N_2273);
nor U3129 (N_3129,N_2479,N_2514);
nor U3130 (N_3130,N_2659,N_2295);
and U3131 (N_3131,N_2873,N_2876);
nor U3132 (N_3132,N_2905,N_2063);
xnor U3133 (N_3133,N_2964,N_2783);
nor U3134 (N_3134,N_2270,N_2834);
nand U3135 (N_3135,N_2078,N_2526);
and U3136 (N_3136,N_2536,N_2604);
nand U3137 (N_3137,N_2890,N_2166);
nand U3138 (N_3138,N_2133,N_2687);
nor U3139 (N_3139,N_2084,N_2623);
nand U3140 (N_3140,N_2762,N_2436);
nand U3141 (N_3141,N_2440,N_2425);
xor U3142 (N_3142,N_2768,N_2188);
xor U3143 (N_3143,N_2159,N_2140);
xor U3144 (N_3144,N_2200,N_2382);
or U3145 (N_3145,N_2582,N_2606);
xor U3146 (N_3146,N_2347,N_2075);
xor U3147 (N_3147,N_2434,N_2708);
nand U3148 (N_3148,N_2861,N_2747);
xnor U3149 (N_3149,N_2956,N_2474);
or U3150 (N_3150,N_2697,N_2558);
and U3151 (N_3151,N_2401,N_2507);
nor U3152 (N_3152,N_2229,N_2052);
xor U3153 (N_3153,N_2911,N_2715);
nand U3154 (N_3154,N_2925,N_2946);
xor U3155 (N_3155,N_2460,N_2966);
and U3156 (N_3156,N_2314,N_2299);
or U3157 (N_3157,N_2608,N_2516);
xnor U3158 (N_3158,N_2320,N_2919);
or U3159 (N_3159,N_2407,N_2801);
nand U3160 (N_3160,N_2390,N_2086);
nor U3161 (N_3161,N_2845,N_2798);
xnor U3162 (N_3162,N_2532,N_2894);
and U3163 (N_3163,N_2119,N_2171);
nor U3164 (N_3164,N_2585,N_2186);
nand U3165 (N_3165,N_2486,N_2949);
nor U3166 (N_3166,N_2473,N_2775);
xor U3167 (N_3167,N_2044,N_2024);
nand U3168 (N_3168,N_2809,N_2753);
xor U3169 (N_3169,N_2652,N_2212);
nor U3170 (N_3170,N_2497,N_2846);
or U3171 (N_3171,N_2750,N_2157);
and U3172 (N_3172,N_2999,N_2830);
nor U3173 (N_3173,N_2037,N_2976);
nor U3174 (N_3174,N_2234,N_2089);
or U3175 (N_3175,N_2312,N_2018);
xnor U3176 (N_3176,N_2605,N_2573);
nand U3177 (N_3177,N_2445,N_2780);
and U3178 (N_3178,N_2466,N_2478);
nor U3179 (N_3179,N_2746,N_2788);
nor U3180 (N_3180,N_2142,N_2096);
nand U3181 (N_3181,N_2546,N_2258);
xnor U3182 (N_3182,N_2615,N_2431);
or U3183 (N_3183,N_2963,N_2327);
xnor U3184 (N_3184,N_2450,N_2799);
or U3185 (N_3185,N_2198,N_2280);
or U3186 (N_3186,N_2088,N_2943);
nand U3187 (N_3187,N_2627,N_2498);
or U3188 (N_3188,N_2238,N_2090);
and U3189 (N_3189,N_2260,N_2257);
nand U3190 (N_3190,N_2189,N_2297);
xnor U3191 (N_3191,N_2855,N_2394);
xor U3192 (N_3192,N_2359,N_2087);
xnor U3193 (N_3193,N_2158,N_2162);
nand U3194 (N_3194,N_2482,N_2912);
or U3195 (N_3195,N_2983,N_2718);
and U3196 (N_3196,N_2534,N_2849);
nor U3197 (N_3197,N_2506,N_2632);
or U3198 (N_3198,N_2083,N_2742);
and U3199 (N_3199,N_2108,N_2923);
and U3200 (N_3200,N_2082,N_2215);
or U3201 (N_3201,N_2393,N_2704);
and U3202 (N_3202,N_2042,N_2626);
nand U3203 (N_3203,N_2356,N_2552);
xnor U3204 (N_3204,N_2244,N_2680);
or U3205 (N_3205,N_2588,N_2684);
nor U3206 (N_3206,N_2457,N_2559);
xor U3207 (N_3207,N_2151,N_2899);
nor U3208 (N_3208,N_2755,N_2261);
nor U3209 (N_3209,N_2291,N_2569);
nor U3210 (N_3210,N_2865,N_2852);
or U3211 (N_3211,N_2647,N_2381);
xnor U3212 (N_3212,N_2802,N_2432);
nand U3213 (N_3213,N_2936,N_2363);
nor U3214 (N_3214,N_2102,N_2259);
nand U3215 (N_3215,N_2977,N_2373);
and U3216 (N_3216,N_2468,N_2958);
nand U3217 (N_3217,N_2763,N_2638);
nor U3218 (N_3218,N_2232,N_2748);
or U3219 (N_3219,N_2579,N_2926);
nor U3220 (N_3220,N_2826,N_2601);
and U3221 (N_3221,N_2719,N_2717);
or U3222 (N_3222,N_2760,N_2709);
xnor U3223 (N_3223,N_2099,N_2664);
nand U3224 (N_3224,N_2069,N_2199);
nand U3225 (N_3225,N_2231,N_2792);
and U3226 (N_3226,N_2376,N_2095);
nor U3227 (N_3227,N_2143,N_2113);
nor U3228 (N_3228,N_2494,N_2181);
or U3229 (N_3229,N_2172,N_2961);
or U3230 (N_3230,N_2348,N_2034);
xor U3231 (N_3231,N_2427,N_2412);
nor U3232 (N_3232,N_2860,N_2617);
nand U3233 (N_3233,N_2774,N_2980);
xor U3234 (N_3234,N_2773,N_2352);
nand U3235 (N_3235,N_2302,N_2703);
or U3236 (N_3236,N_2057,N_2059);
and U3237 (N_3237,N_2251,N_2692);
and U3238 (N_3238,N_2707,N_2272);
nand U3239 (N_3239,N_2173,N_2952);
or U3240 (N_3240,N_2187,N_2738);
or U3241 (N_3241,N_2531,N_2305);
xnor U3242 (N_3242,N_2490,N_2265);
or U3243 (N_3243,N_2093,N_2404);
nand U3244 (N_3244,N_2207,N_2918);
nand U3245 (N_3245,N_2150,N_2463);
nand U3246 (N_3246,N_2164,N_2544);
xnor U3247 (N_3247,N_2233,N_2369);
or U3248 (N_3248,N_2553,N_2787);
xnor U3249 (N_3249,N_2997,N_2076);
nand U3250 (N_3250,N_2055,N_2643);
nor U3251 (N_3251,N_2674,N_2070);
nor U3252 (N_3252,N_2567,N_2098);
xor U3253 (N_3253,N_2848,N_2668);
xnor U3254 (N_3254,N_2262,N_2535);
nor U3255 (N_3255,N_2824,N_2835);
xor U3256 (N_3256,N_2094,N_2679);
xnor U3257 (N_3257,N_2492,N_2733);
xor U3258 (N_3258,N_2741,N_2731);
and U3259 (N_3259,N_2758,N_2555);
nand U3260 (N_3260,N_2851,N_2593);
or U3261 (N_3261,N_2575,N_2339);
and U3262 (N_3262,N_2671,N_2959);
and U3263 (N_3263,N_2496,N_2017);
nor U3264 (N_3264,N_2197,N_2196);
xor U3265 (N_3265,N_2767,N_2612);
and U3266 (N_3266,N_2764,N_2456);
or U3267 (N_3267,N_2694,N_2843);
xor U3268 (N_3268,N_2072,N_2885);
nand U3269 (N_3269,N_2554,N_2942);
nand U3270 (N_3270,N_2309,N_2202);
nand U3271 (N_3271,N_2332,N_2480);
nor U3272 (N_3272,N_2191,N_2361);
and U3273 (N_3273,N_2399,N_2331);
and U3274 (N_3274,N_2111,N_2900);
or U3275 (N_3275,N_2613,N_2138);
nor U3276 (N_3276,N_2937,N_2277);
nor U3277 (N_3277,N_2064,N_2602);
and U3278 (N_3278,N_2006,N_2705);
nand U3279 (N_3279,N_2248,N_2985);
xnor U3280 (N_3280,N_2008,N_2201);
or U3281 (N_3281,N_2644,N_2665);
xor U3282 (N_3282,N_2629,N_2317);
and U3283 (N_3283,N_2002,N_2311);
nor U3284 (N_3284,N_2618,N_2524);
nor U3285 (N_3285,N_2598,N_2307);
or U3286 (N_3286,N_2462,N_2169);
or U3287 (N_3287,N_2673,N_2403);
nand U3288 (N_3288,N_2822,N_2085);
nand U3289 (N_3289,N_2470,N_2645);
or U3290 (N_3290,N_2109,N_2239);
nand U3291 (N_3291,N_2744,N_2806);
nand U3292 (N_3292,N_2712,N_2603);
xnor U3293 (N_3293,N_2782,N_2862);
or U3294 (N_3294,N_2888,N_2435);
xor U3295 (N_3295,N_2663,N_2971);
xnor U3296 (N_3296,N_2145,N_2377);
xnor U3297 (N_3297,N_2660,N_2365);
nor U3298 (N_3298,N_2988,N_2335);
nor U3299 (N_3299,N_2541,N_2041);
xnor U3300 (N_3300,N_2931,N_2349);
or U3301 (N_3301,N_2446,N_2570);
and U3302 (N_3302,N_2204,N_2228);
nor U3303 (N_3303,N_2877,N_2650);
and U3304 (N_3304,N_2130,N_2293);
or U3305 (N_3305,N_2304,N_2185);
or U3306 (N_3306,N_2286,N_2243);
or U3307 (N_3307,N_2116,N_2015);
xnor U3308 (N_3308,N_2066,N_2975);
nor U3309 (N_3309,N_2235,N_2236);
nand U3310 (N_3310,N_2836,N_2411);
xnor U3311 (N_3311,N_2048,N_2454);
and U3312 (N_3312,N_2338,N_2354);
and U3313 (N_3313,N_2019,N_2417);
or U3314 (N_3314,N_2693,N_2969);
xor U3315 (N_3315,N_2045,N_2097);
and U3316 (N_3316,N_2916,N_2515);
xor U3317 (N_3317,N_2004,N_2165);
nor U3318 (N_3318,N_2384,N_2139);
xnor U3319 (N_3319,N_2720,N_2269);
or U3320 (N_3320,N_2451,N_2124);
xnor U3321 (N_3321,N_2691,N_2319);
nor U3322 (N_3322,N_2895,N_2734);
xnor U3323 (N_3323,N_2387,N_2922);
xnor U3324 (N_3324,N_2807,N_2415);
nand U3325 (N_3325,N_2485,N_2091);
and U3326 (N_3326,N_2117,N_2190);
xor U3327 (N_3327,N_2493,N_2060);
nand U3328 (N_3328,N_2073,N_2092);
xor U3329 (N_3329,N_2192,N_2023);
and U3330 (N_3330,N_2662,N_2898);
or U3331 (N_3331,N_2100,N_2504);
or U3332 (N_3332,N_2147,N_2408);
and U3333 (N_3333,N_2580,N_2512);
xnor U3334 (N_3334,N_2220,N_2146);
and U3335 (N_3335,N_2523,N_2226);
and U3336 (N_3336,N_2530,N_2423);
and U3337 (N_3337,N_2875,N_2772);
nor U3338 (N_3338,N_2298,N_2995);
nor U3339 (N_3339,N_2505,N_2525);
and U3340 (N_3340,N_2056,N_2950);
nor U3341 (N_3341,N_2893,N_2242);
or U3342 (N_3342,N_2818,N_2769);
and U3343 (N_3343,N_2886,N_2609);
nand U3344 (N_3344,N_2929,N_2104);
nand U3345 (N_3345,N_2706,N_2035);
and U3346 (N_3346,N_2500,N_2429);
nor U3347 (N_3347,N_2838,N_2808);
or U3348 (N_3348,N_2827,N_2817);
xor U3349 (N_3349,N_2564,N_2321);
or U3350 (N_3350,N_2441,N_2118);
nand U3351 (N_3351,N_2587,N_2521);
nor U3352 (N_3352,N_2914,N_2903);
nor U3353 (N_3353,N_2548,N_2547);
or U3354 (N_3354,N_2658,N_2378);
and U3355 (N_3355,N_2418,N_2539);
nand U3356 (N_3356,N_2549,N_2870);
xnor U3357 (N_3357,N_2637,N_2577);
nor U3358 (N_3358,N_2067,N_2250);
nor U3359 (N_3359,N_2566,N_2823);
xor U3360 (N_3360,N_2968,N_2560);
xor U3361 (N_3361,N_2364,N_2310);
or U3362 (N_3362,N_2979,N_2255);
nor U3363 (N_3363,N_2288,N_2957);
nand U3364 (N_3364,N_2944,N_2424);
nand U3365 (N_3365,N_2449,N_2648);
nand U3366 (N_3366,N_2336,N_2287);
and U3367 (N_3367,N_2448,N_2337);
xor U3368 (N_3368,N_2954,N_2864);
nand U3369 (N_3369,N_2211,N_2333);
nor U3370 (N_3370,N_2811,N_2810);
and U3371 (N_3371,N_2471,N_2657);
nor U3372 (N_3372,N_2633,N_2745);
or U3373 (N_3373,N_2702,N_2907);
or U3374 (N_3374,N_2184,N_2353);
nor U3375 (N_3375,N_2933,N_2634);
or U3376 (N_3376,N_2308,N_2656);
nand U3377 (N_3377,N_2917,N_2355);
nor U3378 (N_3378,N_2889,N_2481);
and U3379 (N_3379,N_2047,N_2442);
and U3380 (N_3380,N_2324,N_2785);
or U3381 (N_3381,N_2160,N_2721);
nand U3382 (N_3382,N_2461,N_2561);
nand U3383 (N_3383,N_2300,N_2274);
nand U3384 (N_3384,N_2318,N_2982);
nand U3385 (N_3385,N_2402,N_2316);
and U3386 (N_3386,N_2107,N_2654);
xor U3387 (N_3387,N_2303,N_2121);
nand U3388 (N_3388,N_2906,N_2292);
nand U3389 (N_3389,N_2214,N_2600);
nor U3390 (N_3390,N_2621,N_2469);
or U3391 (N_3391,N_2127,N_2635);
and U3392 (N_3392,N_2881,N_2007);
nor U3393 (N_3393,N_2858,N_2491);
nor U3394 (N_3394,N_2815,N_2814);
and U3395 (N_3395,N_2245,N_2550);
xnor U3396 (N_3396,N_2832,N_2026);
nor U3397 (N_3397,N_2313,N_2711);
or U3398 (N_3398,N_2455,N_2821);
xnor U3399 (N_3399,N_2572,N_2540);
xor U3400 (N_3400,N_2025,N_2033);
and U3401 (N_3401,N_2597,N_2994);
and U3402 (N_3402,N_2947,N_2049);
and U3403 (N_3403,N_2074,N_2051);
nor U3404 (N_3404,N_2345,N_2032);
xnor U3405 (N_3405,N_2934,N_2271);
nand U3406 (N_3406,N_2992,N_2368);
nand U3407 (N_3407,N_2058,N_2175);
and U3408 (N_3408,N_2502,N_2343);
nor U3409 (N_3409,N_2413,N_2276);
and U3410 (N_3410,N_2754,N_2464);
xnor U3411 (N_3411,N_2438,N_2154);
and U3412 (N_3412,N_2776,N_2978);
nor U3413 (N_3413,N_2043,N_2630);
and U3414 (N_3414,N_2866,N_2027);
xor U3415 (N_3415,N_2825,N_2847);
nand U3416 (N_3416,N_2136,N_2414);
nand U3417 (N_3417,N_2437,N_2000);
nor U3418 (N_3418,N_2488,N_2392);
nor U3419 (N_3419,N_2210,N_2050);
or U3420 (N_3420,N_2315,N_2137);
and U3421 (N_3421,N_2797,N_2682);
nand U3422 (N_3422,N_2584,N_2380);
and U3423 (N_3423,N_2409,N_2856);
and U3424 (N_3424,N_2614,N_2581);
nand U3425 (N_3425,N_2282,N_2871);
and U3426 (N_3426,N_2020,N_2168);
and U3427 (N_3427,N_2590,N_2735);
xnor U3428 (N_3428,N_2400,N_2247);
xnor U3429 (N_3429,N_2850,N_2951);
or U3430 (N_3430,N_2209,N_2596);
xnor U3431 (N_3431,N_2941,N_2696);
nand U3432 (N_3432,N_2557,N_2153);
nand U3433 (N_3433,N_2237,N_2021);
or U3434 (N_3434,N_2766,N_2195);
xor U3435 (N_3435,N_2698,N_2156);
or U3436 (N_3436,N_2517,N_2967);
nor U3437 (N_3437,N_2430,N_2955);
nor U3438 (N_3438,N_2194,N_2938);
nand U3439 (N_3439,N_2761,N_2920);
xor U3440 (N_3440,N_2795,N_2131);
xor U3441 (N_3441,N_2141,N_2476);
nand U3442 (N_3442,N_2285,N_2416);
or U3443 (N_3443,N_2908,N_2819);
xor U3444 (N_3444,N_2366,N_2948);
or U3445 (N_3445,N_2224,N_2386);
nand U3446 (N_3446,N_2740,N_2786);
nor U3447 (N_3447,N_2591,N_2897);
nand U3448 (N_3448,N_2294,N_2729);
xor U3449 (N_3449,N_2538,N_2820);
xnor U3450 (N_3450,N_2079,N_2519);
or U3451 (N_3451,N_2728,N_2726);
xor U3452 (N_3452,N_2651,N_2103);
or U3453 (N_3453,N_2771,N_2759);
xor U3454 (N_3454,N_2989,N_2981);
and U3455 (N_3455,N_2328,N_2275);
nand U3456 (N_3456,N_2594,N_2781);
and U3457 (N_3457,N_2737,N_2221);
or U3458 (N_3458,N_2901,N_2661);
and U3459 (N_3459,N_2447,N_2374);
nand U3460 (N_3460,N_2653,N_2263);
nand U3461 (N_3461,N_2909,N_2636);
xnor U3462 (N_3462,N_2928,N_2595);
and U3463 (N_3463,N_2040,N_2683);
nand U3464 (N_3464,N_2406,N_2439);
and U3465 (N_3465,N_2254,N_2518);
xor U3466 (N_3466,N_2062,N_2484);
or U3467 (N_3467,N_2155,N_2670);
nand U3468 (N_3468,N_2180,N_2114);
and U3469 (N_3469,N_2419,N_2730);
xor U3470 (N_3470,N_2340,N_2010);
or U3471 (N_3471,N_2991,N_2752);
nand U3472 (N_3472,N_2701,N_2879);
nand U3473 (N_3473,N_2789,N_2193);
xor U3474 (N_3474,N_2322,N_2001);
xor U3475 (N_3475,N_2996,N_2217);
nand U3476 (N_3476,N_2794,N_2869);
or U3477 (N_3477,N_2628,N_2281);
nor U3478 (N_3478,N_2129,N_2639);
and U3479 (N_3479,N_2296,N_2128);
or U3480 (N_3480,N_2511,N_2123);
xnor U3481 (N_3481,N_2513,N_2784);
and U3482 (N_3482,N_2240,N_2689);
or U3483 (N_3483,N_2329,N_2323);
nand U3484 (N_3484,N_2422,N_2568);
or U3485 (N_3485,N_2970,N_2725);
nor U3486 (N_3486,N_2453,N_2695);
and U3487 (N_3487,N_2054,N_2583);
nand U3488 (N_3488,N_2749,N_2699);
xor U3489 (N_3489,N_2589,N_2371);
and U3490 (N_3490,N_2206,N_2688);
xor U3491 (N_3491,N_2105,N_2452);
xor U3492 (N_3492,N_2891,N_2397);
nor U3493 (N_3493,N_2268,N_2223);
xor U3494 (N_3494,N_2854,N_2882);
nor U3495 (N_3495,N_2812,N_2071);
or U3496 (N_3496,N_2935,N_2669);
nand U3497 (N_3497,N_2252,N_2805);
xnor U3498 (N_3498,N_2148,N_2793);
xnor U3499 (N_3499,N_2342,N_2666);
nand U3500 (N_3500,N_2195,N_2841);
and U3501 (N_3501,N_2710,N_2473);
and U3502 (N_3502,N_2737,N_2473);
and U3503 (N_3503,N_2514,N_2320);
nor U3504 (N_3504,N_2643,N_2843);
or U3505 (N_3505,N_2834,N_2477);
and U3506 (N_3506,N_2186,N_2371);
xor U3507 (N_3507,N_2251,N_2905);
or U3508 (N_3508,N_2065,N_2949);
or U3509 (N_3509,N_2836,N_2597);
or U3510 (N_3510,N_2079,N_2690);
nor U3511 (N_3511,N_2669,N_2924);
nand U3512 (N_3512,N_2224,N_2903);
or U3513 (N_3513,N_2425,N_2653);
or U3514 (N_3514,N_2859,N_2604);
and U3515 (N_3515,N_2178,N_2675);
nand U3516 (N_3516,N_2406,N_2836);
xor U3517 (N_3517,N_2074,N_2715);
or U3518 (N_3518,N_2502,N_2151);
nor U3519 (N_3519,N_2523,N_2868);
and U3520 (N_3520,N_2574,N_2577);
or U3521 (N_3521,N_2731,N_2653);
nor U3522 (N_3522,N_2961,N_2372);
or U3523 (N_3523,N_2277,N_2515);
nand U3524 (N_3524,N_2678,N_2955);
nand U3525 (N_3525,N_2770,N_2960);
xor U3526 (N_3526,N_2151,N_2988);
nand U3527 (N_3527,N_2030,N_2950);
nor U3528 (N_3528,N_2652,N_2883);
nor U3529 (N_3529,N_2026,N_2483);
or U3530 (N_3530,N_2574,N_2309);
and U3531 (N_3531,N_2202,N_2469);
nand U3532 (N_3532,N_2701,N_2125);
xnor U3533 (N_3533,N_2455,N_2475);
and U3534 (N_3534,N_2163,N_2503);
or U3535 (N_3535,N_2789,N_2523);
nand U3536 (N_3536,N_2141,N_2130);
nor U3537 (N_3537,N_2930,N_2798);
or U3538 (N_3538,N_2889,N_2090);
nand U3539 (N_3539,N_2753,N_2194);
or U3540 (N_3540,N_2556,N_2647);
nand U3541 (N_3541,N_2720,N_2365);
nor U3542 (N_3542,N_2918,N_2616);
xor U3543 (N_3543,N_2021,N_2191);
and U3544 (N_3544,N_2445,N_2242);
xor U3545 (N_3545,N_2447,N_2937);
nor U3546 (N_3546,N_2835,N_2103);
xnor U3547 (N_3547,N_2890,N_2504);
and U3548 (N_3548,N_2107,N_2775);
nand U3549 (N_3549,N_2939,N_2157);
or U3550 (N_3550,N_2162,N_2310);
or U3551 (N_3551,N_2964,N_2588);
and U3552 (N_3552,N_2474,N_2733);
nor U3553 (N_3553,N_2393,N_2447);
and U3554 (N_3554,N_2348,N_2406);
and U3555 (N_3555,N_2145,N_2436);
xor U3556 (N_3556,N_2539,N_2930);
nand U3557 (N_3557,N_2602,N_2507);
or U3558 (N_3558,N_2563,N_2289);
and U3559 (N_3559,N_2826,N_2736);
nand U3560 (N_3560,N_2399,N_2232);
or U3561 (N_3561,N_2908,N_2853);
xnor U3562 (N_3562,N_2911,N_2328);
nand U3563 (N_3563,N_2440,N_2178);
or U3564 (N_3564,N_2386,N_2700);
nor U3565 (N_3565,N_2607,N_2452);
xnor U3566 (N_3566,N_2298,N_2880);
or U3567 (N_3567,N_2110,N_2674);
or U3568 (N_3568,N_2285,N_2533);
xor U3569 (N_3569,N_2790,N_2290);
and U3570 (N_3570,N_2120,N_2804);
nor U3571 (N_3571,N_2830,N_2566);
and U3572 (N_3572,N_2960,N_2437);
and U3573 (N_3573,N_2215,N_2886);
xnor U3574 (N_3574,N_2853,N_2708);
xor U3575 (N_3575,N_2118,N_2168);
nor U3576 (N_3576,N_2506,N_2533);
or U3577 (N_3577,N_2260,N_2661);
or U3578 (N_3578,N_2657,N_2907);
and U3579 (N_3579,N_2873,N_2494);
nor U3580 (N_3580,N_2125,N_2891);
and U3581 (N_3581,N_2031,N_2401);
nand U3582 (N_3582,N_2261,N_2146);
xor U3583 (N_3583,N_2556,N_2921);
nor U3584 (N_3584,N_2706,N_2955);
or U3585 (N_3585,N_2058,N_2331);
or U3586 (N_3586,N_2082,N_2464);
nor U3587 (N_3587,N_2993,N_2555);
nor U3588 (N_3588,N_2985,N_2265);
or U3589 (N_3589,N_2152,N_2752);
and U3590 (N_3590,N_2333,N_2574);
or U3591 (N_3591,N_2142,N_2419);
xnor U3592 (N_3592,N_2635,N_2492);
nand U3593 (N_3593,N_2191,N_2161);
xor U3594 (N_3594,N_2788,N_2632);
and U3595 (N_3595,N_2395,N_2223);
and U3596 (N_3596,N_2073,N_2868);
or U3597 (N_3597,N_2866,N_2286);
or U3598 (N_3598,N_2873,N_2857);
and U3599 (N_3599,N_2030,N_2366);
nor U3600 (N_3600,N_2227,N_2688);
xnor U3601 (N_3601,N_2858,N_2733);
or U3602 (N_3602,N_2780,N_2512);
or U3603 (N_3603,N_2066,N_2262);
nand U3604 (N_3604,N_2516,N_2740);
nor U3605 (N_3605,N_2230,N_2183);
nand U3606 (N_3606,N_2350,N_2467);
nor U3607 (N_3607,N_2468,N_2980);
and U3608 (N_3608,N_2216,N_2586);
and U3609 (N_3609,N_2877,N_2380);
or U3610 (N_3610,N_2539,N_2064);
and U3611 (N_3611,N_2638,N_2803);
nor U3612 (N_3612,N_2287,N_2649);
or U3613 (N_3613,N_2125,N_2801);
nand U3614 (N_3614,N_2904,N_2767);
or U3615 (N_3615,N_2674,N_2137);
nor U3616 (N_3616,N_2951,N_2295);
nand U3617 (N_3617,N_2019,N_2758);
xor U3618 (N_3618,N_2450,N_2271);
nand U3619 (N_3619,N_2403,N_2234);
and U3620 (N_3620,N_2916,N_2067);
xor U3621 (N_3621,N_2417,N_2316);
and U3622 (N_3622,N_2485,N_2149);
or U3623 (N_3623,N_2183,N_2835);
xor U3624 (N_3624,N_2438,N_2186);
and U3625 (N_3625,N_2319,N_2157);
or U3626 (N_3626,N_2085,N_2363);
xor U3627 (N_3627,N_2581,N_2303);
xor U3628 (N_3628,N_2351,N_2535);
or U3629 (N_3629,N_2864,N_2066);
and U3630 (N_3630,N_2503,N_2338);
and U3631 (N_3631,N_2458,N_2212);
xor U3632 (N_3632,N_2573,N_2458);
or U3633 (N_3633,N_2094,N_2148);
and U3634 (N_3634,N_2489,N_2427);
or U3635 (N_3635,N_2485,N_2279);
or U3636 (N_3636,N_2188,N_2786);
and U3637 (N_3637,N_2544,N_2651);
nand U3638 (N_3638,N_2340,N_2088);
and U3639 (N_3639,N_2889,N_2829);
or U3640 (N_3640,N_2047,N_2190);
or U3641 (N_3641,N_2406,N_2640);
xor U3642 (N_3642,N_2624,N_2729);
xnor U3643 (N_3643,N_2274,N_2674);
or U3644 (N_3644,N_2906,N_2341);
xnor U3645 (N_3645,N_2506,N_2279);
and U3646 (N_3646,N_2264,N_2824);
nand U3647 (N_3647,N_2103,N_2694);
nand U3648 (N_3648,N_2192,N_2850);
and U3649 (N_3649,N_2313,N_2224);
and U3650 (N_3650,N_2637,N_2496);
or U3651 (N_3651,N_2040,N_2505);
nor U3652 (N_3652,N_2783,N_2298);
nand U3653 (N_3653,N_2655,N_2416);
nand U3654 (N_3654,N_2699,N_2444);
xnor U3655 (N_3655,N_2950,N_2084);
xor U3656 (N_3656,N_2414,N_2533);
xnor U3657 (N_3657,N_2892,N_2820);
nor U3658 (N_3658,N_2554,N_2829);
nor U3659 (N_3659,N_2374,N_2353);
or U3660 (N_3660,N_2839,N_2932);
xor U3661 (N_3661,N_2254,N_2335);
nand U3662 (N_3662,N_2898,N_2187);
and U3663 (N_3663,N_2180,N_2395);
and U3664 (N_3664,N_2940,N_2654);
nor U3665 (N_3665,N_2975,N_2929);
or U3666 (N_3666,N_2565,N_2119);
nand U3667 (N_3667,N_2653,N_2433);
and U3668 (N_3668,N_2669,N_2056);
or U3669 (N_3669,N_2843,N_2540);
nand U3670 (N_3670,N_2514,N_2591);
and U3671 (N_3671,N_2439,N_2247);
or U3672 (N_3672,N_2888,N_2920);
nor U3673 (N_3673,N_2462,N_2546);
or U3674 (N_3674,N_2756,N_2102);
nor U3675 (N_3675,N_2133,N_2846);
and U3676 (N_3676,N_2147,N_2366);
nor U3677 (N_3677,N_2383,N_2578);
nand U3678 (N_3678,N_2127,N_2752);
xor U3679 (N_3679,N_2655,N_2229);
nand U3680 (N_3680,N_2885,N_2991);
or U3681 (N_3681,N_2674,N_2552);
xor U3682 (N_3682,N_2368,N_2302);
and U3683 (N_3683,N_2500,N_2961);
nor U3684 (N_3684,N_2001,N_2636);
xnor U3685 (N_3685,N_2432,N_2185);
and U3686 (N_3686,N_2647,N_2289);
nand U3687 (N_3687,N_2166,N_2792);
xnor U3688 (N_3688,N_2616,N_2953);
or U3689 (N_3689,N_2942,N_2322);
and U3690 (N_3690,N_2656,N_2694);
nand U3691 (N_3691,N_2967,N_2738);
xor U3692 (N_3692,N_2756,N_2844);
nor U3693 (N_3693,N_2012,N_2296);
nor U3694 (N_3694,N_2332,N_2734);
or U3695 (N_3695,N_2813,N_2941);
or U3696 (N_3696,N_2696,N_2577);
nand U3697 (N_3697,N_2024,N_2520);
xor U3698 (N_3698,N_2661,N_2553);
or U3699 (N_3699,N_2759,N_2809);
xnor U3700 (N_3700,N_2620,N_2089);
and U3701 (N_3701,N_2566,N_2225);
nand U3702 (N_3702,N_2470,N_2111);
nor U3703 (N_3703,N_2667,N_2473);
nand U3704 (N_3704,N_2991,N_2235);
or U3705 (N_3705,N_2970,N_2153);
nand U3706 (N_3706,N_2410,N_2196);
nor U3707 (N_3707,N_2451,N_2231);
or U3708 (N_3708,N_2425,N_2311);
or U3709 (N_3709,N_2822,N_2509);
nand U3710 (N_3710,N_2773,N_2636);
nand U3711 (N_3711,N_2494,N_2965);
and U3712 (N_3712,N_2574,N_2717);
or U3713 (N_3713,N_2944,N_2933);
nand U3714 (N_3714,N_2464,N_2547);
nor U3715 (N_3715,N_2353,N_2997);
or U3716 (N_3716,N_2489,N_2936);
nand U3717 (N_3717,N_2773,N_2724);
and U3718 (N_3718,N_2774,N_2694);
or U3719 (N_3719,N_2366,N_2924);
nand U3720 (N_3720,N_2108,N_2380);
and U3721 (N_3721,N_2098,N_2409);
nor U3722 (N_3722,N_2677,N_2955);
or U3723 (N_3723,N_2494,N_2936);
or U3724 (N_3724,N_2104,N_2699);
or U3725 (N_3725,N_2457,N_2464);
and U3726 (N_3726,N_2532,N_2861);
nand U3727 (N_3727,N_2435,N_2297);
and U3728 (N_3728,N_2221,N_2309);
nand U3729 (N_3729,N_2146,N_2518);
nor U3730 (N_3730,N_2584,N_2731);
xnor U3731 (N_3731,N_2101,N_2567);
nor U3732 (N_3732,N_2845,N_2828);
or U3733 (N_3733,N_2171,N_2174);
nor U3734 (N_3734,N_2006,N_2517);
and U3735 (N_3735,N_2719,N_2508);
xnor U3736 (N_3736,N_2380,N_2405);
nand U3737 (N_3737,N_2063,N_2047);
nor U3738 (N_3738,N_2570,N_2341);
nor U3739 (N_3739,N_2124,N_2291);
and U3740 (N_3740,N_2835,N_2278);
xnor U3741 (N_3741,N_2253,N_2737);
nor U3742 (N_3742,N_2269,N_2809);
nor U3743 (N_3743,N_2882,N_2913);
nor U3744 (N_3744,N_2657,N_2215);
or U3745 (N_3745,N_2165,N_2217);
nand U3746 (N_3746,N_2423,N_2697);
xor U3747 (N_3747,N_2370,N_2593);
nand U3748 (N_3748,N_2297,N_2607);
xor U3749 (N_3749,N_2759,N_2651);
nand U3750 (N_3750,N_2644,N_2479);
xnor U3751 (N_3751,N_2246,N_2708);
and U3752 (N_3752,N_2263,N_2124);
nor U3753 (N_3753,N_2967,N_2444);
or U3754 (N_3754,N_2132,N_2669);
nand U3755 (N_3755,N_2664,N_2690);
nor U3756 (N_3756,N_2977,N_2141);
nand U3757 (N_3757,N_2136,N_2623);
nand U3758 (N_3758,N_2192,N_2870);
or U3759 (N_3759,N_2242,N_2488);
or U3760 (N_3760,N_2213,N_2623);
and U3761 (N_3761,N_2943,N_2965);
nand U3762 (N_3762,N_2084,N_2299);
nor U3763 (N_3763,N_2288,N_2943);
xor U3764 (N_3764,N_2285,N_2747);
and U3765 (N_3765,N_2537,N_2889);
xnor U3766 (N_3766,N_2275,N_2921);
and U3767 (N_3767,N_2916,N_2870);
nor U3768 (N_3768,N_2945,N_2313);
xnor U3769 (N_3769,N_2426,N_2747);
or U3770 (N_3770,N_2999,N_2417);
xnor U3771 (N_3771,N_2213,N_2986);
nand U3772 (N_3772,N_2265,N_2479);
nand U3773 (N_3773,N_2568,N_2034);
nor U3774 (N_3774,N_2385,N_2492);
or U3775 (N_3775,N_2419,N_2384);
nand U3776 (N_3776,N_2584,N_2271);
nor U3777 (N_3777,N_2531,N_2735);
nand U3778 (N_3778,N_2235,N_2537);
nor U3779 (N_3779,N_2691,N_2448);
or U3780 (N_3780,N_2209,N_2351);
xnor U3781 (N_3781,N_2714,N_2306);
nand U3782 (N_3782,N_2582,N_2701);
nor U3783 (N_3783,N_2864,N_2206);
nor U3784 (N_3784,N_2632,N_2657);
nand U3785 (N_3785,N_2280,N_2595);
and U3786 (N_3786,N_2859,N_2671);
or U3787 (N_3787,N_2331,N_2072);
and U3788 (N_3788,N_2567,N_2341);
or U3789 (N_3789,N_2261,N_2421);
xnor U3790 (N_3790,N_2399,N_2641);
xor U3791 (N_3791,N_2408,N_2988);
and U3792 (N_3792,N_2204,N_2273);
and U3793 (N_3793,N_2263,N_2036);
or U3794 (N_3794,N_2180,N_2279);
and U3795 (N_3795,N_2129,N_2903);
and U3796 (N_3796,N_2423,N_2365);
xor U3797 (N_3797,N_2069,N_2176);
or U3798 (N_3798,N_2700,N_2420);
nand U3799 (N_3799,N_2853,N_2369);
nor U3800 (N_3800,N_2869,N_2799);
xor U3801 (N_3801,N_2953,N_2918);
xor U3802 (N_3802,N_2840,N_2573);
nor U3803 (N_3803,N_2430,N_2908);
xor U3804 (N_3804,N_2543,N_2401);
nor U3805 (N_3805,N_2199,N_2829);
and U3806 (N_3806,N_2661,N_2494);
nor U3807 (N_3807,N_2932,N_2573);
nand U3808 (N_3808,N_2718,N_2636);
nand U3809 (N_3809,N_2390,N_2948);
nand U3810 (N_3810,N_2874,N_2675);
nand U3811 (N_3811,N_2514,N_2654);
nand U3812 (N_3812,N_2558,N_2840);
nor U3813 (N_3813,N_2401,N_2519);
nor U3814 (N_3814,N_2132,N_2453);
or U3815 (N_3815,N_2862,N_2030);
and U3816 (N_3816,N_2379,N_2948);
nand U3817 (N_3817,N_2996,N_2468);
nand U3818 (N_3818,N_2482,N_2694);
and U3819 (N_3819,N_2140,N_2839);
and U3820 (N_3820,N_2879,N_2688);
and U3821 (N_3821,N_2624,N_2419);
and U3822 (N_3822,N_2024,N_2034);
and U3823 (N_3823,N_2591,N_2026);
nand U3824 (N_3824,N_2363,N_2105);
nor U3825 (N_3825,N_2477,N_2494);
nand U3826 (N_3826,N_2423,N_2775);
xnor U3827 (N_3827,N_2582,N_2906);
nor U3828 (N_3828,N_2676,N_2523);
or U3829 (N_3829,N_2661,N_2679);
and U3830 (N_3830,N_2951,N_2033);
and U3831 (N_3831,N_2148,N_2166);
nand U3832 (N_3832,N_2852,N_2497);
xor U3833 (N_3833,N_2020,N_2904);
nand U3834 (N_3834,N_2596,N_2123);
xnor U3835 (N_3835,N_2570,N_2620);
nand U3836 (N_3836,N_2031,N_2768);
nor U3837 (N_3837,N_2478,N_2462);
xnor U3838 (N_3838,N_2822,N_2343);
nor U3839 (N_3839,N_2712,N_2111);
nor U3840 (N_3840,N_2281,N_2877);
xnor U3841 (N_3841,N_2160,N_2506);
and U3842 (N_3842,N_2671,N_2205);
nand U3843 (N_3843,N_2135,N_2462);
nor U3844 (N_3844,N_2070,N_2062);
or U3845 (N_3845,N_2104,N_2752);
xor U3846 (N_3846,N_2172,N_2971);
nand U3847 (N_3847,N_2827,N_2989);
or U3848 (N_3848,N_2559,N_2383);
xnor U3849 (N_3849,N_2324,N_2580);
or U3850 (N_3850,N_2637,N_2752);
or U3851 (N_3851,N_2368,N_2770);
and U3852 (N_3852,N_2826,N_2283);
nand U3853 (N_3853,N_2947,N_2210);
or U3854 (N_3854,N_2552,N_2225);
nand U3855 (N_3855,N_2603,N_2022);
xor U3856 (N_3856,N_2112,N_2144);
or U3857 (N_3857,N_2550,N_2679);
xnor U3858 (N_3858,N_2005,N_2660);
nand U3859 (N_3859,N_2497,N_2261);
nand U3860 (N_3860,N_2596,N_2155);
nor U3861 (N_3861,N_2841,N_2474);
nand U3862 (N_3862,N_2795,N_2840);
or U3863 (N_3863,N_2352,N_2040);
and U3864 (N_3864,N_2658,N_2113);
or U3865 (N_3865,N_2844,N_2011);
and U3866 (N_3866,N_2413,N_2634);
nor U3867 (N_3867,N_2790,N_2746);
and U3868 (N_3868,N_2864,N_2458);
and U3869 (N_3869,N_2912,N_2512);
xor U3870 (N_3870,N_2576,N_2095);
nor U3871 (N_3871,N_2301,N_2829);
xor U3872 (N_3872,N_2403,N_2685);
and U3873 (N_3873,N_2860,N_2477);
nand U3874 (N_3874,N_2490,N_2507);
nand U3875 (N_3875,N_2133,N_2205);
and U3876 (N_3876,N_2621,N_2537);
nand U3877 (N_3877,N_2447,N_2193);
nand U3878 (N_3878,N_2716,N_2200);
nand U3879 (N_3879,N_2064,N_2924);
nand U3880 (N_3880,N_2928,N_2543);
nand U3881 (N_3881,N_2100,N_2684);
or U3882 (N_3882,N_2850,N_2629);
or U3883 (N_3883,N_2587,N_2135);
xor U3884 (N_3884,N_2739,N_2643);
nand U3885 (N_3885,N_2251,N_2935);
xor U3886 (N_3886,N_2417,N_2233);
nor U3887 (N_3887,N_2753,N_2125);
nand U3888 (N_3888,N_2700,N_2087);
nor U3889 (N_3889,N_2866,N_2395);
or U3890 (N_3890,N_2703,N_2847);
or U3891 (N_3891,N_2741,N_2875);
xnor U3892 (N_3892,N_2734,N_2252);
nor U3893 (N_3893,N_2602,N_2925);
or U3894 (N_3894,N_2732,N_2268);
nand U3895 (N_3895,N_2920,N_2007);
or U3896 (N_3896,N_2312,N_2815);
and U3897 (N_3897,N_2946,N_2280);
or U3898 (N_3898,N_2927,N_2805);
and U3899 (N_3899,N_2727,N_2671);
or U3900 (N_3900,N_2353,N_2144);
xor U3901 (N_3901,N_2882,N_2368);
xnor U3902 (N_3902,N_2400,N_2617);
or U3903 (N_3903,N_2605,N_2765);
nor U3904 (N_3904,N_2514,N_2162);
and U3905 (N_3905,N_2058,N_2002);
or U3906 (N_3906,N_2176,N_2100);
xor U3907 (N_3907,N_2806,N_2596);
nand U3908 (N_3908,N_2972,N_2630);
or U3909 (N_3909,N_2762,N_2264);
nor U3910 (N_3910,N_2623,N_2546);
or U3911 (N_3911,N_2038,N_2575);
xnor U3912 (N_3912,N_2439,N_2622);
nand U3913 (N_3913,N_2584,N_2683);
nand U3914 (N_3914,N_2433,N_2440);
nor U3915 (N_3915,N_2575,N_2462);
nand U3916 (N_3916,N_2699,N_2600);
nand U3917 (N_3917,N_2137,N_2234);
and U3918 (N_3918,N_2344,N_2521);
xnor U3919 (N_3919,N_2834,N_2735);
xnor U3920 (N_3920,N_2512,N_2168);
xnor U3921 (N_3921,N_2969,N_2601);
nand U3922 (N_3922,N_2627,N_2713);
nor U3923 (N_3923,N_2930,N_2744);
and U3924 (N_3924,N_2853,N_2175);
nor U3925 (N_3925,N_2218,N_2995);
nand U3926 (N_3926,N_2223,N_2539);
or U3927 (N_3927,N_2720,N_2004);
nor U3928 (N_3928,N_2124,N_2563);
xor U3929 (N_3929,N_2027,N_2600);
and U3930 (N_3930,N_2886,N_2639);
or U3931 (N_3931,N_2539,N_2344);
and U3932 (N_3932,N_2483,N_2204);
nand U3933 (N_3933,N_2389,N_2394);
xor U3934 (N_3934,N_2036,N_2807);
xnor U3935 (N_3935,N_2668,N_2015);
or U3936 (N_3936,N_2925,N_2148);
xnor U3937 (N_3937,N_2356,N_2633);
or U3938 (N_3938,N_2422,N_2267);
and U3939 (N_3939,N_2565,N_2778);
and U3940 (N_3940,N_2879,N_2679);
nor U3941 (N_3941,N_2928,N_2426);
nor U3942 (N_3942,N_2092,N_2268);
nor U3943 (N_3943,N_2122,N_2180);
and U3944 (N_3944,N_2725,N_2714);
xnor U3945 (N_3945,N_2195,N_2762);
nand U3946 (N_3946,N_2209,N_2326);
xnor U3947 (N_3947,N_2705,N_2480);
nand U3948 (N_3948,N_2935,N_2083);
nand U3949 (N_3949,N_2164,N_2677);
and U3950 (N_3950,N_2350,N_2576);
xor U3951 (N_3951,N_2702,N_2348);
xnor U3952 (N_3952,N_2367,N_2475);
xor U3953 (N_3953,N_2608,N_2340);
nand U3954 (N_3954,N_2646,N_2119);
nor U3955 (N_3955,N_2416,N_2048);
or U3956 (N_3956,N_2604,N_2568);
or U3957 (N_3957,N_2586,N_2339);
or U3958 (N_3958,N_2534,N_2144);
or U3959 (N_3959,N_2392,N_2372);
nand U3960 (N_3960,N_2513,N_2411);
xor U3961 (N_3961,N_2985,N_2043);
and U3962 (N_3962,N_2613,N_2176);
nand U3963 (N_3963,N_2251,N_2589);
or U3964 (N_3964,N_2445,N_2116);
nand U3965 (N_3965,N_2763,N_2550);
nor U3966 (N_3966,N_2769,N_2480);
xor U3967 (N_3967,N_2081,N_2919);
xor U3968 (N_3968,N_2599,N_2777);
nand U3969 (N_3969,N_2703,N_2676);
nor U3970 (N_3970,N_2352,N_2672);
and U3971 (N_3971,N_2392,N_2892);
or U3972 (N_3972,N_2114,N_2932);
nor U3973 (N_3973,N_2716,N_2185);
and U3974 (N_3974,N_2509,N_2939);
or U3975 (N_3975,N_2578,N_2727);
nor U3976 (N_3976,N_2353,N_2099);
nor U3977 (N_3977,N_2468,N_2811);
and U3978 (N_3978,N_2395,N_2171);
nand U3979 (N_3979,N_2305,N_2100);
nor U3980 (N_3980,N_2250,N_2096);
nand U3981 (N_3981,N_2895,N_2766);
and U3982 (N_3982,N_2331,N_2349);
nor U3983 (N_3983,N_2784,N_2369);
nand U3984 (N_3984,N_2997,N_2472);
or U3985 (N_3985,N_2919,N_2467);
nand U3986 (N_3986,N_2013,N_2385);
or U3987 (N_3987,N_2591,N_2106);
xnor U3988 (N_3988,N_2572,N_2483);
nand U3989 (N_3989,N_2372,N_2057);
nor U3990 (N_3990,N_2212,N_2010);
nor U3991 (N_3991,N_2360,N_2285);
or U3992 (N_3992,N_2407,N_2952);
nand U3993 (N_3993,N_2335,N_2293);
nor U3994 (N_3994,N_2797,N_2266);
nand U3995 (N_3995,N_2995,N_2447);
and U3996 (N_3996,N_2137,N_2421);
xor U3997 (N_3997,N_2352,N_2200);
nor U3998 (N_3998,N_2951,N_2679);
nand U3999 (N_3999,N_2246,N_2083);
or U4000 (N_4000,N_3399,N_3401);
xor U4001 (N_4001,N_3215,N_3291);
xnor U4002 (N_4002,N_3369,N_3659);
nor U4003 (N_4003,N_3122,N_3031);
and U4004 (N_4004,N_3212,N_3879);
xnor U4005 (N_4005,N_3042,N_3715);
xnor U4006 (N_4006,N_3668,N_3863);
or U4007 (N_4007,N_3253,N_3465);
nand U4008 (N_4008,N_3374,N_3266);
nand U4009 (N_4009,N_3514,N_3023);
and U4010 (N_4010,N_3492,N_3595);
nor U4011 (N_4011,N_3414,N_3798);
xnor U4012 (N_4012,N_3724,N_3098);
nor U4013 (N_4013,N_3976,N_3300);
xor U4014 (N_4014,N_3845,N_3411);
xor U4015 (N_4015,N_3982,N_3282);
nand U4016 (N_4016,N_3048,N_3925);
xnor U4017 (N_4017,N_3051,N_3679);
and U4018 (N_4018,N_3788,N_3706);
and U4019 (N_4019,N_3174,N_3487);
and U4020 (N_4020,N_3755,N_3373);
or U4021 (N_4021,N_3442,N_3546);
and U4022 (N_4022,N_3379,N_3025);
or U4023 (N_4023,N_3992,N_3571);
and U4024 (N_4024,N_3349,N_3314);
or U4025 (N_4025,N_3406,N_3702);
or U4026 (N_4026,N_3592,N_3240);
nand U4027 (N_4027,N_3527,N_3566);
nand U4028 (N_4028,N_3880,N_3631);
and U4029 (N_4029,N_3780,N_3607);
nor U4030 (N_4030,N_3513,N_3856);
and U4031 (N_4031,N_3508,N_3108);
nand U4032 (N_4032,N_3929,N_3172);
or U4033 (N_4033,N_3959,N_3061);
xnor U4034 (N_4034,N_3783,N_3146);
nor U4035 (N_4035,N_3320,N_3611);
nor U4036 (N_4036,N_3425,N_3207);
nand U4037 (N_4037,N_3481,N_3342);
nor U4038 (N_4038,N_3228,N_3101);
nand U4039 (N_4039,N_3325,N_3745);
or U4040 (N_4040,N_3111,N_3383);
nor U4041 (N_4041,N_3941,N_3472);
or U4042 (N_4042,N_3700,N_3616);
or U4043 (N_4043,N_3524,N_3348);
or U4044 (N_4044,N_3775,N_3115);
and U4045 (N_4045,N_3877,N_3157);
xnor U4046 (N_4046,N_3405,N_3971);
nor U4047 (N_4047,N_3210,N_3004);
xnor U4048 (N_4048,N_3366,N_3757);
nor U4049 (N_4049,N_3244,N_3462);
nand U4050 (N_4050,N_3554,N_3063);
or U4051 (N_4051,N_3445,N_3623);
or U4052 (N_4052,N_3365,N_3562);
nand U4053 (N_4053,N_3091,N_3183);
xor U4054 (N_4054,N_3728,N_3867);
nand U4055 (N_4055,N_3648,N_3036);
xnor U4056 (N_4056,N_3764,N_3092);
nor U4057 (N_4057,N_3910,N_3854);
or U4058 (N_4058,N_3693,N_3579);
and U4059 (N_4059,N_3694,N_3956);
xor U4060 (N_4060,N_3301,N_3541);
or U4061 (N_4061,N_3243,N_3664);
nand U4062 (N_4062,N_3802,N_3915);
and U4063 (N_4063,N_3681,N_3621);
or U4064 (N_4064,N_3958,N_3433);
nand U4065 (N_4065,N_3520,N_3467);
nor U4066 (N_4066,N_3797,N_3066);
nor U4067 (N_4067,N_3476,N_3273);
or U4068 (N_4068,N_3874,N_3153);
nand U4069 (N_4069,N_3135,N_3474);
or U4070 (N_4070,N_3489,N_3670);
or U4071 (N_4071,N_3404,N_3924);
and U4072 (N_4072,N_3417,N_3974);
nor U4073 (N_4073,N_3175,N_3677);
or U4074 (N_4074,N_3627,N_3857);
and U4075 (N_4075,N_3418,N_3713);
nor U4076 (N_4076,N_3493,N_3263);
or U4077 (N_4077,N_3899,N_3671);
nand U4078 (N_4078,N_3011,N_3707);
xnor U4079 (N_4079,N_3573,N_3550);
nand U4080 (N_4080,N_3129,N_3130);
xnor U4081 (N_4081,N_3390,N_3722);
and U4082 (N_4082,N_3475,N_3164);
and U4083 (N_4083,N_3261,N_3416);
nand U4084 (N_4084,N_3464,N_3766);
nor U4085 (N_4085,N_3620,N_3890);
or U4086 (N_4086,N_3944,N_3269);
nor U4087 (N_4087,N_3270,N_3154);
or U4088 (N_4088,N_3962,N_3860);
xnor U4089 (N_4089,N_3807,N_3099);
xor U4090 (N_4090,N_3653,N_3605);
xor U4091 (N_4091,N_3217,N_3556);
xor U4092 (N_4092,N_3892,N_3703);
or U4093 (N_4093,N_3463,N_3704);
and U4094 (N_4094,N_3371,N_3306);
nor U4095 (N_4095,N_3771,N_3555);
nand U4096 (N_4096,N_3444,N_3260);
and U4097 (N_4097,N_3937,N_3778);
and U4098 (N_4098,N_3523,N_3312);
nand U4099 (N_4099,N_3906,N_3237);
or U4100 (N_4100,N_3491,N_3165);
xor U4101 (N_4101,N_3361,N_3341);
or U4102 (N_4102,N_3537,N_3821);
nand U4103 (N_4103,N_3255,N_3156);
xnor U4104 (N_4104,N_3787,N_3859);
or U4105 (N_4105,N_3034,N_3120);
nor U4106 (N_4106,N_3948,N_3458);
nand U4107 (N_4107,N_3311,N_3285);
nor U4108 (N_4108,N_3055,N_3482);
or U4109 (N_4109,N_3988,N_3678);
nand U4110 (N_4110,N_3152,N_3330);
xor U4111 (N_4111,N_3104,N_3299);
nor U4112 (N_4112,N_3049,N_3375);
xnor U4113 (N_4113,N_3795,N_3690);
and U4114 (N_4114,N_3904,N_3675);
xor U4115 (N_4115,N_3391,N_3252);
xor U4116 (N_4116,N_3498,N_3117);
xor U4117 (N_4117,N_3598,N_3995);
or U4118 (N_4118,N_3264,N_3274);
or U4119 (N_4119,N_3786,N_3714);
or U4120 (N_4120,N_3202,N_3769);
nor U4121 (N_4121,N_3984,N_3068);
nor U4122 (N_4122,N_3112,N_3913);
nand U4123 (N_4123,N_3497,N_3238);
and U4124 (N_4124,N_3485,N_3058);
nor U4125 (N_4125,N_3125,N_3869);
or U4126 (N_4126,N_3222,N_3056);
xor U4127 (N_4127,N_3624,N_3750);
or U4128 (N_4128,N_3754,N_3993);
nand U4129 (N_4129,N_3567,N_3332);
or U4130 (N_4130,N_3533,N_3712);
or U4131 (N_4131,N_3582,N_3136);
nor U4132 (N_4132,N_3114,N_3897);
xnor U4133 (N_4133,N_3116,N_3473);
xnor U4134 (N_4134,N_3727,N_3310);
nor U4135 (N_4135,N_3149,N_3811);
or U4136 (N_4136,N_3448,N_3538);
nor U4137 (N_4137,N_3643,N_3697);
and U4138 (N_4138,N_3708,N_3219);
and U4139 (N_4139,N_3640,N_3022);
nor U4140 (N_4140,N_3759,N_3224);
xnor U4141 (N_4141,N_3593,N_3415);
nand U4142 (N_4142,N_3437,N_3740);
nor U4143 (N_4143,N_3326,N_3572);
xnor U4144 (N_4144,N_3903,N_3526);
xor U4145 (N_4145,N_3124,N_3355);
xor U4146 (N_4146,N_3638,N_3357);
xor U4147 (N_4147,N_3020,N_3543);
nand U4148 (N_4148,N_3635,N_3050);
and U4149 (N_4149,N_3466,N_3198);
nand U4150 (N_4150,N_3468,N_3015);
xnor U4151 (N_4151,N_3730,N_3356);
or U4152 (N_4152,N_3434,N_3074);
and U4153 (N_4153,N_3059,N_3280);
nor U4154 (N_4154,N_3109,N_3604);
and U4155 (N_4155,N_3189,N_3214);
nor U4156 (N_4156,N_3762,N_3600);
nor U4157 (N_4157,N_3557,N_3096);
and U4158 (N_4158,N_3873,N_3179);
or U4159 (N_4159,N_3585,N_3477);
and U4160 (N_4160,N_3725,N_3580);
xor U4161 (N_4161,N_3118,N_3594);
xor U4162 (N_4162,N_3753,N_3053);
xor U4163 (N_4163,N_3826,N_3323);
or U4164 (N_4164,N_3934,N_3281);
nand U4165 (N_4165,N_3551,N_3632);
nand U4166 (N_4166,N_3946,N_3652);
nand U4167 (N_4167,N_3177,N_3601);
nand U4168 (N_4168,N_3184,N_3749);
or U4169 (N_4169,N_3824,N_3794);
nor U4170 (N_4170,N_3721,N_3163);
and U4171 (N_4171,N_3254,N_3071);
and U4172 (N_4172,N_3303,N_3279);
and U4173 (N_4173,N_3268,N_3609);
xor U4174 (N_4174,N_3459,N_3338);
nand U4175 (N_4175,N_3241,N_3045);
xnor U4176 (N_4176,N_3235,N_3901);
or U4177 (N_4177,N_3486,N_3139);
xnor U4178 (N_4178,N_3287,N_3980);
xor U4179 (N_4179,N_3446,N_3319);
nor U4180 (N_4180,N_3169,N_3449);
nand U4181 (N_4181,N_3460,N_3699);
and U4182 (N_4182,N_3077,N_3686);
or U4183 (N_4183,N_3825,N_3996);
xor U4184 (N_4184,N_3171,N_3606);
xor U4185 (N_4185,N_3997,N_3711);
nand U4186 (N_4186,N_3443,N_3256);
nor U4187 (N_4187,N_3176,N_3005);
nor U4188 (N_4188,N_3168,N_3999);
xnor U4189 (N_4189,N_3024,N_3830);
nor U4190 (N_4190,N_3160,N_3367);
and U4191 (N_4191,N_3204,N_3297);
and U4192 (N_4192,N_3480,N_3608);
nand U4193 (N_4193,N_3181,N_3196);
xor U4194 (N_4194,N_3003,N_3190);
xnor U4195 (N_4195,N_3781,N_3471);
and U4196 (N_4196,N_3872,N_3292);
and U4197 (N_4197,N_3351,N_3855);
or U4198 (N_4198,N_3536,N_3695);
or U4199 (N_4199,N_3803,N_3547);
nor U4200 (N_4200,N_3575,N_3747);
xor U4201 (N_4201,N_3046,N_3994);
nand U4202 (N_4202,N_3683,N_3666);
and U4203 (N_4203,N_3088,N_3603);
or U4204 (N_4204,N_3075,N_3065);
nor U4205 (N_4205,N_3896,N_3954);
or U4206 (N_4206,N_3134,N_3614);
or U4207 (N_4207,N_3871,N_3990);
or U4208 (N_4208,N_3552,N_3322);
nand U4209 (N_4209,N_3876,N_3333);
or U4210 (N_4210,N_3398,N_3983);
nor U4211 (N_4211,N_3245,N_3938);
nor U4212 (N_4212,N_3021,N_3942);
nor U4213 (N_4213,N_3558,N_3344);
nor U4214 (N_4214,N_3284,N_3751);
nand U4215 (N_4215,N_3343,N_3364);
or U4216 (N_4216,N_3085,N_3395);
nor U4217 (N_4217,N_3569,N_3836);
nor U4218 (N_4218,N_3862,N_3738);
and U4219 (N_4219,N_3353,N_3810);
and U4220 (N_4220,N_3288,N_3622);
nand U4221 (N_4221,N_3935,N_3090);
or U4222 (N_4222,N_3731,N_3597);
nand U4223 (N_4223,N_3345,N_3528);
xor U4224 (N_4224,N_3461,N_3150);
and U4225 (N_4225,N_3438,N_3436);
xnor U4226 (N_4226,N_3248,N_3969);
nand U4227 (N_4227,N_3973,N_3972);
nor U4228 (N_4228,N_3510,N_3895);
or U4229 (N_4229,N_3372,N_3362);
or U4230 (N_4230,N_3073,N_3133);
or U4231 (N_4231,N_3363,N_3483);
or U4232 (N_4232,N_3806,N_3271);
or U4233 (N_4233,N_3232,N_3885);
or U4234 (N_4234,N_3216,N_3397);
and U4235 (N_4235,N_3809,N_3815);
or U4236 (N_4236,N_3734,N_3672);
or U4237 (N_4237,N_3853,N_3574);
xnor U4238 (N_4238,N_3739,N_3911);
and U4239 (N_4239,N_3535,N_3080);
nand U4240 (N_4240,N_3705,N_3441);
and U4241 (N_4241,N_3435,N_3752);
or U4242 (N_4242,N_3408,N_3262);
xnor U4243 (N_4243,N_3503,N_3384);
nand U4244 (N_4244,N_3777,N_3522);
nand U4245 (N_4245,N_3186,N_3298);
or U4246 (N_4246,N_3852,N_3131);
nor U4247 (N_4247,N_3170,N_3865);
nand U4248 (N_4248,N_3278,N_3737);
xnor U4249 (N_4249,N_3199,N_3121);
and U4250 (N_4250,N_3456,N_3804);
or U4251 (N_4251,N_3576,N_3007);
nor U4252 (N_4252,N_3043,N_3933);
and U4253 (N_4253,N_3293,N_3336);
nand U4254 (N_4254,N_3661,N_3975);
or U4255 (N_4255,N_3894,N_3741);
and U4256 (N_4256,N_3054,N_3642);
or U4257 (N_4257,N_3392,N_3064);
nand U4258 (N_4258,N_3633,N_3113);
nor U4259 (N_4259,N_3354,N_3626);
nor U4260 (N_4260,N_3192,N_3589);
xor U4261 (N_4261,N_3187,N_3422);
nor U4262 (N_4262,N_3878,N_3968);
nand U4263 (N_4263,N_3818,N_3094);
xnor U4264 (N_4264,N_3917,N_3035);
nor U4265 (N_4265,N_3805,N_3837);
and U4266 (N_4266,N_3955,N_3506);
nand U4267 (N_4267,N_3615,N_3507);
nand U4268 (N_4268,N_3394,N_3010);
nand U4269 (N_4269,N_3258,N_3978);
xor U4270 (N_4270,N_3765,N_3516);
xnor U4271 (N_4271,N_3613,N_3540);
nor U4272 (N_4272,N_3410,N_3823);
xnor U4273 (N_4273,N_3950,N_3820);
xor U4274 (N_4274,N_3286,N_3329);
or U4275 (N_4275,N_3610,N_3421);
nand U4276 (N_4276,N_3315,N_3313);
or U4277 (N_4277,N_3309,N_3561);
xor U4278 (N_4278,N_3719,N_3733);
nor U4279 (N_4279,N_3389,N_3432);
nor U4280 (N_4280,N_3521,N_3839);
nand U4281 (N_4281,N_3221,N_3742);
or U4282 (N_4282,N_3070,N_3039);
xor U4283 (N_4283,N_3017,N_3834);
or U4284 (N_4284,N_3902,N_3939);
nor U4285 (N_4285,N_3454,N_3674);
xor U4286 (N_4286,N_3455,N_3819);
xor U4287 (N_4287,N_3000,N_3205);
nand U4288 (N_4288,N_3927,N_3531);
and U4289 (N_4289,N_3137,N_3801);
nor U4290 (N_4290,N_3145,N_3223);
or U4291 (N_4291,N_3583,N_3584);
xnor U4292 (N_4292,N_3866,N_3518);
and U4293 (N_4293,N_3760,N_3726);
nor U4294 (N_4294,N_3026,N_3928);
or U4295 (N_4295,N_3380,N_3612);
or U4296 (N_4296,N_3930,N_3542);
and U4297 (N_4297,N_3662,N_3440);
nor U4298 (N_4298,N_3967,N_3308);
xnor U4299 (N_4299,N_3086,N_3785);
xnor U4300 (N_4300,N_3041,N_3986);
and U4301 (N_4301,N_3529,N_3140);
nor U4302 (N_4302,N_3530,N_3985);
and U4303 (N_4303,N_3525,N_3509);
nand U4304 (N_4304,N_3790,N_3875);
or U4305 (N_4305,N_3359,N_3057);
nor U4306 (N_4306,N_3987,N_3779);
and U4307 (N_4307,N_3965,N_3393);
or U4308 (N_4308,N_3549,N_3898);
nand U4309 (N_4309,N_3470,N_3206);
nand U4310 (N_4310,N_3701,N_3409);
nor U4311 (N_4311,N_3716,N_3267);
nor U4312 (N_4312,N_3961,N_3013);
xnor U4313 (N_4313,N_3447,N_3833);
or U4314 (N_4314,N_3776,N_3484);
or U4315 (N_4315,N_3816,N_3912);
xor U4316 (N_4316,N_3377,N_3062);
xnor U4317 (N_4317,N_3123,N_3012);
nand U4318 (N_4318,N_3100,N_3193);
nand U4319 (N_4319,N_3658,N_3352);
xor U4320 (N_4320,N_3296,N_3209);
or U4321 (N_4321,N_3155,N_3981);
xnor U4322 (N_4322,N_3226,N_3439);
xor U4323 (N_4323,N_3893,N_3709);
and U4324 (N_4324,N_3923,N_3849);
nor U4325 (N_4325,N_3891,N_3103);
and U4326 (N_4326,N_3568,N_3494);
and U4327 (N_4327,N_3989,N_3814);
xnor U4328 (N_4328,N_3289,N_3864);
xnor U4329 (N_4329,N_3040,N_3774);
xor U4330 (N_4330,N_3147,N_3951);
xnor U4331 (N_4331,N_3964,N_3502);
or U4332 (N_4332,N_3478,N_3387);
nor U4333 (N_4333,N_3106,N_3431);
nand U4334 (N_4334,N_3386,N_3072);
xor U4335 (N_4335,N_3213,N_3499);
nor U4336 (N_4336,N_3316,N_3014);
or U4337 (N_4337,N_3501,N_3963);
or U4338 (N_4338,N_3843,N_3334);
nor U4339 (N_4339,N_3423,N_3835);
and U4340 (N_4340,N_3926,N_3947);
xor U4341 (N_4341,N_3838,N_3655);
nor U4342 (N_4342,N_3799,N_3909);
nor U4343 (N_4343,N_3469,N_3553);
xor U4344 (N_4344,N_3259,N_3102);
nor U4345 (N_4345,N_3692,N_3630);
and U4346 (N_4346,N_3305,N_3644);
nor U4347 (N_4347,N_3784,N_3490);
and U4348 (N_4348,N_3360,N_3126);
nand U4349 (N_4349,N_3685,N_3647);
and U4350 (N_4350,N_3908,N_3680);
and U4351 (N_4351,N_3560,N_3078);
and U4352 (N_4352,N_3868,N_3002);
and U4353 (N_4353,N_3654,N_3141);
xor U4354 (N_4354,N_3639,N_3596);
xnor U4355 (N_4355,N_3663,N_3105);
and U4356 (N_4356,N_3687,N_3208);
nand U4357 (N_4357,N_3318,N_3945);
nor U4358 (N_4358,N_3087,N_3698);
nand U4359 (N_4359,N_3496,N_3628);
nor U4360 (N_4360,N_3773,N_3173);
or U4361 (N_4361,N_3918,N_3511);
nand U4362 (N_4362,N_3304,N_3257);
nor U4363 (N_4363,N_3038,N_3230);
xor U4364 (N_4364,N_3500,N_3841);
or U4365 (N_4365,N_3166,N_3646);
xor U4366 (N_4366,N_3559,N_3870);
or U4367 (N_4367,N_3931,N_3563);
nand U4368 (N_4368,N_3220,N_3182);
xor U4369 (N_4369,N_3729,N_3167);
and U4370 (N_4370,N_3744,N_3669);
xor U4371 (N_4371,N_3407,N_3132);
nor U4372 (N_4372,N_3382,N_3327);
nand U4373 (N_4373,N_3162,N_3717);
or U4374 (N_4374,N_3019,N_3539);
nand U4375 (N_4375,N_3665,N_3159);
xor U4376 (N_4376,N_3651,N_3921);
nand U4377 (N_4377,N_3907,N_3889);
or U4378 (N_4378,N_3932,N_3916);
and U4379 (N_4379,N_3185,N_3376);
xor U4380 (N_4380,N_3335,N_3515);
nor U4381 (N_4381,N_3427,N_3089);
and U4382 (N_4382,N_3684,N_3791);
nor U4383 (N_4383,N_3812,N_3277);
xnor U4384 (N_4384,N_3519,N_3808);
nand U4385 (N_4385,N_3718,N_3337);
and U4386 (N_4386,N_3998,N_3792);
xor U4387 (N_4387,N_3018,N_3689);
xor U4388 (N_4388,N_3505,N_3844);
nand U4389 (N_4389,N_3504,N_3370);
nand U4390 (N_4390,N_3676,N_3246);
nand U4391 (N_4391,N_3142,N_3957);
nor U4392 (N_4392,N_3800,N_3251);
xor U4393 (N_4393,N_3381,N_3625);
xor U4394 (N_4394,N_3636,N_3829);
and U4395 (N_4395,N_3746,N_3424);
nand U4396 (N_4396,N_3067,N_3302);
xnor U4397 (N_4397,N_3832,N_3158);
or U4398 (N_4398,N_3645,N_3107);
and U4399 (N_4399,N_3250,N_3940);
nand U4400 (N_4400,N_3403,N_3242);
nor U4401 (N_4401,N_3758,N_3883);
and U4402 (N_4402,N_3548,N_3861);
xor U4403 (N_4403,N_3236,N_3884);
xor U4404 (N_4404,N_3720,N_3736);
xor U4405 (N_4405,N_3060,N_3001);
nor U4406 (N_4406,N_3688,N_3827);
nand U4407 (N_4407,N_3634,N_3570);
nor U4408 (N_4408,N_3346,N_3770);
xnor U4409 (N_4409,N_3368,N_3590);
nor U4410 (N_4410,N_3195,N_3905);
nand U4411 (N_4411,N_3822,N_3828);
and U4412 (N_4412,N_3008,N_3188);
nor U4413 (N_4413,N_3032,N_3201);
nor U4414 (N_4414,N_3307,N_3385);
xnor U4415 (N_4415,N_3637,N_3846);
nor U4416 (N_4416,N_3479,N_3656);
and U4417 (N_4417,N_3030,N_3900);
nor U4418 (N_4418,N_3339,N_3850);
nor U4419 (N_4419,N_3991,N_3817);
nand U4420 (N_4420,N_3457,N_3881);
or U4421 (N_4421,N_3922,N_3710);
xor U4422 (N_4422,N_3272,N_3952);
nand U4423 (N_4423,N_3813,N_3691);
nor U4424 (N_4424,N_3276,N_3265);
or U4425 (N_4425,N_3960,N_3290);
xor U4426 (N_4426,N_3450,N_3488);
and U4427 (N_4427,N_3082,N_3180);
or U4428 (N_4428,N_3097,N_3970);
and U4429 (N_4429,N_3378,N_3295);
nand U4430 (N_4430,N_3657,N_3979);
nor U4431 (N_4431,N_3936,N_3197);
xor U4432 (N_4432,N_3200,N_3402);
and U4433 (N_4433,N_3682,N_3888);
nand U4434 (N_4434,N_3761,N_3842);
xnor U4435 (N_4435,N_3079,N_3234);
xnor U4436 (N_4436,N_3793,N_3429);
nand U4437 (N_4437,N_3565,N_3696);
nand U4438 (N_4438,N_3083,N_3044);
xnor U4439 (N_4439,N_3851,N_3178);
nor U4440 (N_4440,N_3452,N_3577);
nand U4441 (N_4441,N_3191,N_3420);
nor U4442 (N_4442,N_3649,N_3789);
nand U4443 (N_4443,N_3396,N_3069);
or U4444 (N_4444,N_3599,N_3831);
xor U4445 (N_4445,N_3016,N_3581);
or U4446 (N_4446,N_3028,N_3110);
nand U4447 (N_4447,N_3275,N_3629);
xnor U4448 (N_4448,N_3358,N_3564);
and U4449 (N_4449,N_3587,N_3194);
or U4450 (N_4450,N_3009,N_3148);
nor U4451 (N_4451,N_3430,N_3578);
nand U4452 (N_4452,N_3037,N_3027);
or U4453 (N_4453,N_3588,N_3847);
nor U4454 (N_4454,N_3047,N_3426);
nand U4455 (N_4455,N_3419,N_3328);
nand U4456 (N_4456,N_3227,N_3667);
xor U4457 (N_4457,N_3211,N_3350);
nor U4458 (N_4458,N_3660,N_3138);
or U4459 (N_4459,N_3914,N_3886);
or U4460 (N_4460,N_3324,N_3650);
nand U4461 (N_4461,N_3767,N_3919);
or U4462 (N_4462,N_3081,N_3119);
or U4463 (N_4463,N_3768,N_3735);
or U4464 (N_4464,N_3495,N_3532);
or U4465 (N_4465,N_3413,N_3756);
nor U4466 (N_4466,N_3029,N_3591);
or U4467 (N_4467,N_3517,N_3249);
nand U4468 (N_4468,N_3545,N_3340);
xor U4469 (N_4469,N_3128,N_3641);
xnor U4470 (N_4470,N_3006,N_3151);
nand U4471 (N_4471,N_3161,N_3239);
or U4472 (N_4472,N_3943,N_3076);
nor U4473 (N_4473,N_3321,N_3748);
nor U4474 (N_4474,N_3618,N_3127);
and U4475 (N_4475,N_3203,N_3084);
or U4476 (N_4476,N_3772,N_3882);
nor U4477 (N_4477,N_3052,N_3143);
nor U4478 (N_4478,N_3966,N_3586);
xnor U4479 (N_4479,N_3920,N_3796);
or U4480 (N_4480,N_3451,N_3231);
nor U4481 (N_4481,N_3723,N_3317);
xnor U4482 (N_4482,N_3887,N_3294);
nor U4483 (N_4483,N_3544,N_3453);
and U4484 (N_4484,N_3233,N_3673);
or U4485 (N_4485,N_3225,N_3953);
or U4486 (N_4486,N_3412,N_3617);
or U4487 (N_4487,N_3512,N_3229);
and U4488 (N_4488,N_3602,N_3840);
nand U4489 (N_4489,N_3033,N_3858);
and U4490 (N_4490,N_3095,N_3848);
and U4491 (N_4491,N_3347,N_3400);
and U4492 (N_4492,N_3093,N_3782);
nor U4493 (N_4493,N_3247,N_3283);
and U4494 (N_4494,N_3388,N_3763);
nor U4495 (N_4495,N_3619,N_3977);
and U4496 (N_4496,N_3732,N_3428);
or U4497 (N_4497,N_3534,N_3144);
or U4498 (N_4498,N_3949,N_3218);
xor U4499 (N_4499,N_3331,N_3743);
or U4500 (N_4500,N_3431,N_3379);
nand U4501 (N_4501,N_3847,N_3192);
or U4502 (N_4502,N_3343,N_3450);
nand U4503 (N_4503,N_3987,N_3946);
nor U4504 (N_4504,N_3514,N_3618);
nand U4505 (N_4505,N_3710,N_3508);
and U4506 (N_4506,N_3529,N_3692);
xor U4507 (N_4507,N_3023,N_3268);
nand U4508 (N_4508,N_3523,N_3170);
nor U4509 (N_4509,N_3085,N_3624);
or U4510 (N_4510,N_3705,N_3987);
or U4511 (N_4511,N_3714,N_3434);
nor U4512 (N_4512,N_3991,N_3519);
xor U4513 (N_4513,N_3753,N_3982);
or U4514 (N_4514,N_3948,N_3346);
xor U4515 (N_4515,N_3001,N_3090);
nor U4516 (N_4516,N_3620,N_3975);
nor U4517 (N_4517,N_3017,N_3805);
and U4518 (N_4518,N_3251,N_3385);
or U4519 (N_4519,N_3030,N_3707);
nor U4520 (N_4520,N_3087,N_3532);
and U4521 (N_4521,N_3852,N_3809);
and U4522 (N_4522,N_3613,N_3700);
nand U4523 (N_4523,N_3853,N_3373);
nand U4524 (N_4524,N_3897,N_3825);
nor U4525 (N_4525,N_3124,N_3806);
xor U4526 (N_4526,N_3296,N_3781);
or U4527 (N_4527,N_3489,N_3346);
xor U4528 (N_4528,N_3775,N_3323);
or U4529 (N_4529,N_3082,N_3370);
or U4530 (N_4530,N_3989,N_3738);
xor U4531 (N_4531,N_3360,N_3701);
xor U4532 (N_4532,N_3566,N_3409);
nand U4533 (N_4533,N_3511,N_3857);
nand U4534 (N_4534,N_3661,N_3617);
xnor U4535 (N_4535,N_3639,N_3461);
nand U4536 (N_4536,N_3635,N_3149);
xnor U4537 (N_4537,N_3374,N_3874);
nor U4538 (N_4538,N_3973,N_3930);
nor U4539 (N_4539,N_3740,N_3625);
nand U4540 (N_4540,N_3213,N_3765);
nor U4541 (N_4541,N_3287,N_3208);
xor U4542 (N_4542,N_3271,N_3876);
and U4543 (N_4543,N_3884,N_3585);
xor U4544 (N_4544,N_3737,N_3476);
or U4545 (N_4545,N_3791,N_3797);
and U4546 (N_4546,N_3909,N_3668);
and U4547 (N_4547,N_3672,N_3376);
nor U4548 (N_4548,N_3051,N_3542);
and U4549 (N_4549,N_3277,N_3477);
nor U4550 (N_4550,N_3382,N_3766);
or U4551 (N_4551,N_3273,N_3992);
nor U4552 (N_4552,N_3544,N_3411);
xor U4553 (N_4553,N_3120,N_3278);
xnor U4554 (N_4554,N_3792,N_3753);
nand U4555 (N_4555,N_3186,N_3473);
or U4556 (N_4556,N_3482,N_3295);
or U4557 (N_4557,N_3966,N_3885);
xnor U4558 (N_4558,N_3664,N_3840);
nor U4559 (N_4559,N_3573,N_3906);
and U4560 (N_4560,N_3946,N_3003);
and U4561 (N_4561,N_3844,N_3319);
xor U4562 (N_4562,N_3377,N_3542);
xor U4563 (N_4563,N_3931,N_3642);
nor U4564 (N_4564,N_3355,N_3037);
or U4565 (N_4565,N_3731,N_3769);
and U4566 (N_4566,N_3307,N_3700);
xor U4567 (N_4567,N_3431,N_3430);
or U4568 (N_4568,N_3712,N_3896);
nand U4569 (N_4569,N_3304,N_3969);
or U4570 (N_4570,N_3057,N_3143);
nand U4571 (N_4571,N_3571,N_3456);
nand U4572 (N_4572,N_3226,N_3262);
and U4573 (N_4573,N_3375,N_3884);
xor U4574 (N_4574,N_3490,N_3294);
xnor U4575 (N_4575,N_3901,N_3341);
or U4576 (N_4576,N_3699,N_3356);
and U4577 (N_4577,N_3476,N_3956);
nor U4578 (N_4578,N_3420,N_3816);
and U4579 (N_4579,N_3319,N_3296);
or U4580 (N_4580,N_3358,N_3592);
nand U4581 (N_4581,N_3002,N_3416);
nor U4582 (N_4582,N_3270,N_3315);
nand U4583 (N_4583,N_3616,N_3081);
or U4584 (N_4584,N_3227,N_3664);
nor U4585 (N_4585,N_3232,N_3114);
or U4586 (N_4586,N_3097,N_3122);
nor U4587 (N_4587,N_3588,N_3995);
nand U4588 (N_4588,N_3524,N_3761);
nor U4589 (N_4589,N_3553,N_3883);
and U4590 (N_4590,N_3639,N_3097);
or U4591 (N_4591,N_3980,N_3894);
xor U4592 (N_4592,N_3074,N_3424);
or U4593 (N_4593,N_3123,N_3637);
nor U4594 (N_4594,N_3574,N_3703);
and U4595 (N_4595,N_3092,N_3105);
nand U4596 (N_4596,N_3367,N_3273);
xnor U4597 (N_4597,N_3311,N_3762);
or U4598 (N_4598,N_3478,N_3721);
nor U4599 (N_4599,N_3921,N_3976);
nor U4600 (N_4600,N_3430,N_3956);
and U4601 (N_4601,N_3166,N_3700);
or U4602 (N_4602,N_3450,N_3387);
or U4603 (N_4603,N_3119,N_3442);
and U4604 (N_4604,N_3957,N_3550);
nand U4605 (N_4605,N_3504,N_3820);
nor U4606 (N_4606,N_3845,N_3804);
or U4607 (N_4607,N_3334,N_3027);
xor U4608 (N_4608,N_3559,N_3384);
nor U4609 (N_4609,N_3675,N_3396);
xor U4610 (N_4610,N_3989,N_3907);
nor U4611 (N_4611,N_3255,N_3034);
nand U4612 (N_4612,N_3539,N_3117);
or U4613 (N_4613,N_3429,N_3768);
xnor U4614 (N_4614,N_3058,N_3167);
or U4615 (N_4615,N_3706,N_3074);
nor U4616 (N_4616,N_3658,N_3588);
or U4617 (N_4617,N_3354,N_3620);
xor U4618 (N_4618,N_3842,N_3705);
nand U4619 (N_4619,N_3037,N_3426);
nand U4620 (N_4620,N_3412,N_3875);
or U4621 (N_4621,N_3390,N_3580);
nor U4622 (N_4622,N_3108,N_3134);
xnor U4623 (N_4623,N_3155,N_3129);
xor U4624 (N_4624,N_3272,N_3825);
nor U4625 (N_4625,N_3429,N_3704);
nor U4626 (N_4626,N_3522,N_3144);
and U4627 (N_4627,N_3695,N_3568);
or U4628 (N_4628,N_3711,N_3691);
and U4629 (N_4629,N_3036,N_3841);
xor U4630 (N_4630,N_3498,N_3097);
nand U4631 (N_4631,N_3196,N_3931);
and U4632 (N_4632,N_3494,N_3689);
nand U4633 (N_4633,N_3107,N_3113);
nand U4634 (N_4634,N_3609,N_3933);
nor U4635 (N_4635,N_3508,N_3532);
or U4636 (N_4636,N_3715,N_3858);
and U4637 (N_4637,N_3797,N_3926);
nor U4638 (N_4638,N_3929,N_3482);
nand U4639 (N_4639,N_3092,N_3032);
nand U4640 (N_4640,N_3951,N_3158);
nor U4641 (N_4641,N_3526,N_3618);
or U4642 (N_4642,N_3491,N_3703);
or U4643 (N_4643,N_3189,N_3862);
nand U4644 (N_4644,N_3949,N_3272);
and U4645 (N_4645,N_3440,N_3953);
nand U4646 (N_4646,N_3058,N_3341);
xnor U4647 (N_4647,N_3244,N_3417);
nor U4648 (N_4648,N_3722,N_3313);
nand U4649 (N_4649,N_3619,N_3214);
nand U4650 (N_4650,N_3063,N_3183);
or U4651 (N_4651,N_3388,N_3755);
xor U4652 (N_4652,N_3549,N_3590);
xnor U4653 (N_4653,N_3959,N_3312);
or U4654 (N_4654,N_3206,N_3753);
or U4655 (N_4655,N_3429,N_3010);
nor U4656 (N_4656,N_3499,N_3249);
nor U4657 (N_4657,N_3894,N_3912);
nand U4658 (N_4658,N_3032,N_3845);
xnor U4659 (N_4659,N_3285,N_3740);
and U4660 (N_4660,N_3457,N_3961);
nand U4661 (N_4661,N_3578,N_3600);
xnor U4662 (N_4662,N_3449,N_3122);
nand U4663 (N_4663,N_3571,N_3077);
nand U4664 (N_4664,N_3819,N_3563);
or U4665 (N_4665,N_3431,N_3159);
or U4666 (N_4666,N_3890,N_3719);
xor U4667 (N_4667,N_3536,N_3581);
and U4668 (N_4668,N_3986,N_3908);
or U4669 (N_4669,N_3333,N_3298);
xor U4670 (N_4670,N_3611,N_3848);
nor U4671 (N_4671,N_3198,N_3488);
or U4672 (N_4672,N_3479,N_3162);
or U4673 (N_4673,N_3964,N_3646);
or U4674 (N_4674,N_3060,N_3393);
and U4675 (N_4675,N_3912,N_3090);
nor U4676 (N_4676,N_3625,N_3680);
nor U4677 (N_4677,N_3378,N_3446);
and U4678 (N_4678,N_3292,N_3570);
xor U4679 (N_4679,N_3046,N_3922);
nand U4680 (N_4680,N_3501,N_3217);
or U4681 (N_4681,N_3525,N_3501);
or U4682 (N_4682,N_3156,N_3489);
nand U4683 (N_4683,N_3982,N_3739);
or U4684 (N_4684,N_3041,N_3012);
and U4685 (N_4685,N_3168,N_3254);
and U4686 (N_4686,N_3261,N_3844);
or U4687 (N_4687,N_3771,N_3321);
and U4688 (N_4688,N_3170,N_3155);
nor U4689 (N_4689,N_3628,N_3258);
xor U4690 (N_4690,N_3478,N_3555);
and U4691 (N_4691,N_3313,N_3387);
nor U4692 (N_4692,N_3867,N_3908);
nor U4693 (N_4693,N_3142,N_3983);
or U4694 (N_4694,N_3058,N_3132);
or U4695 (N_4695,N_3149,N_3052);
xnor U4696 (N_4696,N_3828,N_3030);
nand U4697 (N_4697,N_3601,N_3940);
xor U4698 (N_4698,N_3177,N_3095);
nand U4699 (N_4699,N_3295,N_3647);
nor U4700 (N_4700,N_3388,N_3516);
or U4701 (N_4701,N_3190,N_3029);
and U4702 (N_4702,N_3019,N_3351);
or U4703 (N_4703,N_3306,N_3777);
nor U4704 (N_4704,N_3635,N_3485);
and U4705 (N_4705,N_3356,N_3719);
and U4706 (N_4706,N_3699,N_3672);
nand U4707 (N_4707,N_3236,N_3071);
nor U4708 (N_4708,N_3869,N_3882);
nand U4709 (N_4709,N_3370,N_3176);
nor U4710 (N_4710,N_3008,N_3659);
nand U4711 (N_4711,N_3154,N_3012);
nand U4712 (N_4712,N_3010,N_3446);
xnor U4713 (N_4713,N_3030,N_3260);
or U4714 (N_4714,N_3754,N_3853);
xnor U4715 (N_4715,N_3240,N_3013);
xor U4716 (N_4716,N_3011,N_3766);
or U4717 (N_4717,N_3239,N_3520);
xor U4718 (N_4718,N_3001,N_3155);
or U4719 (N_4719,N_3416,N_3936);
nand U4720 (N_4720,N_3884,N_3862);
nand U4721 (N_4721,N_3845,N_3861);
nor U4722 (N_4722,N_3150,N_3122);
nor U4723 (N_4723,N_3478,N_3380);
and U4724 (N_4724,N_3581,N_3059);
xor U4725 (N_4725,N_3670,N_3987);
and U4726 (N_4726,N_3098,N_3478);
or U4727 (N_4727,N_3295,N_3629);
or U4728 (N_4728,N_3738,N_3618);
and U4729 (N_4729,N_3841,N_3521);
xor U4730 (N_4730,N_3889,N_3307);
nor U4731 (N_4731,N_3749,N_3143);
nor U4732 (N_4732,N_3931,N_3312);
nor U4733 (N_4733,N_3936,N_3113);
xnor U4734 (N_4734,N_3771,N_3710);
xor U4735 (N_4735,N_3567,N_3687);
nor U4736 (N_4736,N_3290,N_3694);
nand U4737 (N_4737,N_3373,N_3055);
xnor U4738 (N_4738,N_3461,N_3736);
or U4739 (N_4739,N_3008,N_3126);
and U4740 (N_4740,N_3141,N_3558);
or U4741 (N_4741,N_3464,N_3722);
or U4742 (N_4742,N_3465,N_3153);
and U4743 (N_4743,N_3021,N_3780);
nand U4744 (N_4744,N_3716,N_3417);
nor U4745 (N_4745,N_3989,N_3342);
nor U4746 (N_4746,N_3881,N_3183);
and U4747 (N_4747,N_3890,N_3391);
nor U4748 (N_4748,N_3419,N_3180);
nand U4749 (N_4749,N_3333,N_3581);
or U4750 (N_4750,N_3390,N_3205);
nor U4751 (N_4751,N_3902,N_3265);
nand U4752 (N_4752,N_3239,N_3839);
nor U4753 (N_4753,N_3287,N_3678);
and U4754 (N_4754,N_3452,N_3326);
nand U4755 (N_4755,N_3837,N_3713);
xor U4756 (N_4756,N_3481,N_3600);
nor U4757 (N_4757,N_3795,N_3954);
or U4758 (N_4758,N_3536,N_3086);
or U4759 (N_4759,N_3150,N_3179);
nor U4760 (N_4760,N_3467,N_3683);
nand U4761 (N_4761,N_3445,N_3826);
nand U4762 (N_4762,N_3992,N_3711);
nor U4763 (N_4763,N_3416,N_3909);
xnor U4764 (N_4764,N_3200,N_3912);
nand U4765 (N_4765,N_3179,N_3965);
and U4766 (N_4766,N_3543,N_3107);
nand U4767 (N_4767,N_3789,N_3479);
and U4768 (N_4768,N_3770,N_3307);
and U4769 (N_4769,N_3662,N_3852);
nor U4770 (N_4770,N_3193,N_3946);
or U4771 (N_4771,N_3838,N_3682);
nor U4772 (N_4772,N_3315,N_3089);
and U4773 (N_4773,N_3201,N_3604);
and U4774 (N_4774,N_3652,N_3035);
xor U4775 (N_4775,N_3411,N_3781);
or U4776 (N_4776,N_3705,N_3467);
nor U4777 (N_4777,N_3651,N_3478);
xnor U4778 (N_4778,N_3736,N_3126);
and U4779 (N_4779,N_3058,N_3085);
or U4780 (N_4780,N_3330,N_3225);
nand U4781 (N_4781,N_3865,N_3813);
and U4782 (N_4782,N_3475,N_3544);
and U4783 (N_4783,N_3992,N_3725);
xor U4784 (N_4784,N_3141,N_3698);
xnor U4785 (N_4785,N_3220,N_3162);
nor U4786 (N_4786,N_3366,N_3981);
and U4787 (N_4787,N_3544,N_3220);
xnor U4788 (N_4788,N_3474,N_3611);
nand U4789 (N_4789,N_3463,N_3284);
nand U4790 (N_4790,N_3850,N_3080);
nand U4791 (N_4791,N_3124,N_3451);
xor U4792 (N_4792,N_3356,N_3403);
nor U4793 (N_4793,N_3856,N_3535);
nor U4794 (N_4794,N_3042,N_3794);
and U4795 (N_4795,N_3562,N_3042);
nor U4796 (N_4796,N_3577,N_3701);
or U4797 (N_4797,N_3912,N_3495);
nand U4798 (N_4798,N_3074,N_3865);
or U4799 (N_4799,N_3193,N_3341);
nor U4800 (N_4800,N_3004,N_3659);
nor U4801 (N_4801,N_3617,N_3249);
nor U4802 (N_4802,N_3795,N_3558);
xor U4803 (N_4803,N_3892,N_3752);
and U4804 (N_4804,N_3363,N_3780);
xnor U4805 (N_4805,N_3980,N_3160);
nor U4806 (N_4806,N_3967,N_3842);
nand U4807 (N_4807,N_3096,N_3111);
nand U4808 (N_4808,N_3664,N_3690);
and U4809 (N_4809,N_3369,N_3661);
nand U4810 (N_4810,N_3500,N_3435);
or U4811 (N_4811,N_3117,N_3052);
or U4812 (N_4812,N_3862,N_3580);
xnor U4813 (N_4813,N_3186,N_3352);
and U4814 (N_4814,N_3028,N_3281);
nand U4815 (N_4815,N_3983,N_3110);
nor U4816 (N_4816,N_3484,N_3265);
nor U4817 (N_4817,N_3198,N_3272);
or U4818 (N_4818,N_3318,N_3590);
nor U4819 (N_4819,N_3701,N_3645);
nand U4820 (N_4820,N_3470,N_3504);
or U4821 (N_4821,N_3507,N_3174);
nand U4822 (N_4822,N_3480,N_3078);
xor U4823 (N_4823,N_3599,N_3483);
or U4824 (N_4824,N_3492,N_3440);
nor U4825 (N_4825,N_3518,N_3347);
nand U4826 (N_4826,N_3906,N_3115);
xor U4827 (N_4827,N_3805,N_3116);
xor U4828 (N_4828,N_3069,N_3726);
xnor U4829 (N_4829,N_3451,N_3994);
xor U4830 (N_4830,N_3400,N_3677);
nor U4831 (N_4831,N_3921,N_3597);
xor U4832 (N_4832,N_3971,N_3361);
nand U4833 (N_4833,N_3630,N_3668);
nand U4834 (N_4834,N_3776,N_3243);
and U4835 (N_4835,N_3248,N_3851);
or U4836 (N_4836,N_3889,N_3176);
and U4837 (N_4837,N_3286,N_3620);
xnor U4838 (N_4838,N_3066,N_3734);
nand U4839 (N_4839,N_3907,N_3590);
nand U4840 (N_4840,N_3648,N_3682);
nor U4841 (N_4841,N_3142,N_3716);
and U4842 (N_4842,N_3918,N_3686);
nor U4843 (N_4843,N_3212,N_3848);
and U4844 (N_4844,N_3769,N_3654);
and U4845 (N_4845,N_3830,N_3850);
and U4846 (N_4846,N_3902,N_3428);
nand U4847 (N_4847,N_3443,N_3099);
nand U4848 (N_4848,N_3642,N_3623);
xnor U4849 (N_4849,N_3631,N_3901);
or U4850 (N_4850,N_3656,N_3768);
and U4851 (N_4851,N_3688,N_3737);
or U4852 (N_4852,N_3889,N_3489);
nand U4853 (N_4853,N_3179,N_3998);
and U4854 (N_4854,N_3024,N_3378);
xnor U4855 (N_4855,N_3872,N_3002);
xor U4856 (N_4856,N_3667,N_3672);
and U4857 (N_4857,N_3554,N_3105);
and U4858 (N_4858,N_3111,N_3058);
and U4859 (N_4859,N_3568,N_3778);
xnor U4860 (N_4860,N_3629,N_3473);
nor U4861 (N_4861,N_3960,N_3377);
nand U4862 (N_4862,N_3906,N_3938);
xor U4863 (N_4863,N_3423,N_3099);
and U4864 (N_4864,N_3900,N_3175);
and U4865 (N_4865,N_3575,N_3573);
xnor U4866 (N_4866,N_3629,N_3766);
and U4867 (N_4867,N_3418,N_3779);
nor U4868 (N_4868,N_3671,N_3368);
nand U4869 (N_4869,N_3788,N_3385);
nor U4870 (N_4870,N_3611,N_3952);
nor U4871 (N_4871,N_3896,N_3316);
or U4872 (N_4872,N_3010,N_3116);
and U4873 (N_4873,N_3157,N_3087);
xnor U4874 (N_4874,N_3289,N_3517);
xor U4875 (N_4875,N_3072,N_3646);
nand U4876 (N_4876,N_3185,N_3909);
nand U4877 (N_4877,N_3497,N_3893);
xor U4878 (N_4878,N_3735,N_3430);
nor U4879 (N_4879,N_3995,N_3275);
xor U4880 (N_4880,N_3316,N_3194);
and U4881 (N_4881,N_3863,N_3639);
or U4882 (N_4882,N_3760,N_3054);
or U4883 (N_4883,N_3193,N_3979);
or U4884 (N_4884,N_3920,N_3558);
xor U4885 (N_4885,N_3170,N_3826);
and U4886 (N_4886,N_3371,N_3481);
xnor U4887 (N_4887,N_3765,N_3580);
and U4888 (N_4888,N_3961,N_3481);
xor U4889 (N_4889,N_3752,N_3438);
xnor U4890 (N_4890,N_3195,N_3126);
nand U4891 (N_4891,N_3374,N_3699);
or U4892 (N_4892,N_3185,N_3327);
xnor U4893 (N_4893,N_3041,N_3226);
or U4894 (N_4894,N_3437,N_3162);
or U4895 (N_4895,N_3739,N_3534);
and U4896 (N_4896,N_3397,N_3819);
nand U4897 (N_4897,N_3639,N_3860);
and U4898 (N_4898,N_3750,N_3848);
nor U4899 (N_4899,N_3208,N_3624);
xor U4900 (N_4900,N_3124,N_3345);
and U4901 (N_4901,N_3530,N_3979);
nand U4902 (N_4902,N_3862,N_3677);
and U4903 (N_4903,N_3119,N_3301);
or U4904 (N_4904,N_3325,N_3424);
nand U4905 (N_4905,N_3329,N_3361);
nand U4906 (N_4906,N_3151,N_3611);
and U4907 (N_4907,N_3808,N_3866);
and U4908 (N_4908,N_3091,N_3803);
xnor U4909 (N_4909,N_3633,N_3229);
xor U4910 (N_4910,N_3445,N_3018);
nor U4911 (N_4911,N_3556,N_3315);
nor U4912 (N_4912,N_3185,N_3579);
and U4913 (N_4913,N_3452,N_3351);
or U4914 (N_4914,N_3269,N_3718);
xor U4915 (N_4915,N_3096,N_3266);
xor U4916 (N_4916,N_3996,N_3951);
nor U4917 (N_4917,N_3510,N_3749);
nor U4918 (N_4918,N_3654,N_3454);
or U4919 (N_4919,N_3677,N_3110);
or U4920 (N_4920,N_3942,N_3647);
xor U4921 (N_4921,N_3442,N_3312);
nand U4922 (N_4922,N_3141,N_3560);
nor U4923 (N_4923,N_3981,N_3307);
or U4924 (N_4924,N_3646,N_3983);
nor U4925 (N_4925,N_3682,N_3936);
nor U4926 (N_4926,N_3580,N_3874);
and U4927 (N_4927,N_3287,N_3311);
nand U4928 (N_4928,N_3369,N_3811);
and U4929 (N_4929,N_3902,N_3412);
xnor U4930 (N_4930,N_3143,N_3740);
and U4931 (N_4931,N_3743,N_3523);
and U4932 (N_4932,N_3687,N_3377);
or U4933 (N_4933,N_3174,N_3445);
nand U4934 (N_4934,N_3494,N_3920);
and U4935 (N_4935,N_3949,N_3036);
and U4936 (N_4936,N_3895,N_3180);
nand U4937 (N_4937,N_3986,N_3332);
nor U4938 (N_4938,N_3158,N_3250);
or U4939 (N_4939,N_3266,N_3824);
or U4940 (N_4940,N_3188,N_3989);
and U4941 (N_4941,N_3002,N_3988);
xnor U4942 (N_4942,N_3333,N_3172);
or U4943 (N_4943,N_3541,N_3072);
xor U4944 (N_4944,N_3622,N_3090);
and U4945 (N_4945,N_3196,N_3872);
nor U4946 (N_4946,N_3403,N_3489);
or U4947 (N_4947,N_3705,N_3494);
nand U4948 (N_4948,N_3549,N_3787);
or U4949 (N_4949,N_3609,N_3697);
or U4950 (N_4950,N_3081,N_3169);
xor U4951 (N_4951,N_3570,N_3510);
nor U4952 (N_4952,N_3487,N_3772);
and U4953 (N_4953,N_3386,N_3326);
nor U4954 (N_4954,N_3882,N_3633);
and U4955 (N_4955,N_3637,N_3208);
or U4956 (N_4956,N_3638,N_3857);
and U4957 (N_4957,N_3779,N_3562);
xor U4958 (N_4958,N_3585,N_3074);
nand U4959 (N_4959,N_3529,N_3736);
xor U4960 (N_4960,N_3409,N_3810);
xnor U4961 (N_4961,N_3606,N_3149);
or U4962 (N_4962,N_3725,N_3253);
xnor U4963 (N_4963,N_3635,N_3156);
xor U4964 (N_4964,N_3525,N_3056);
or U4965 (N_4965,N_3140,N_3217);
nand U4966 (N_4966,N_3031,N_3526);
or U4967 (N_4967,N_3541,N_3807);
xnor U4968 (N_4968,N_3521,N_3262);
nor U4969 (N_4969,N_3000,N_3272);
nor U4970 (N_4970,N_3335,N_3648);
xor U4971 (N_4971,N_3739,N_3694);
and U4972 (N_4972,N_3309,N_3480);
xor U4973 (N_4973,N_3551,N_3014);
nor U4974 (N_4974,N_3497,N_3464);
or U4975 (N_4975,N_3010,N_3047);
nor U4976 (N_4976,N_3126,N_3408);
nand U4977 (N_4977,N_3028,N_3855);
nand U4978 (N_4978,N_3881,N_3532);
and U4979 (N_4979,N_3455,N_3660);
nor U4980 (N_4980,N_3043,N_3692);
xnor U4981 (N_4981,N_3995,N_3700);
or U4982 (N_4982,N_3960,N_3932);
nand U4983 (N_4983,N_3554,N_3180);
nand U4984 (N_4984,N_3080,N_3408);
nor U4985 (N_4985,N_3207,N_3735);
nor U4986 (N_4986,N_3954,N_3544);
nor U4987 (N_4987,N_3558,N_3465);
nand U4988 (N_4988,N_3077,N_3988);
nor U4989 (N_4989,N_3175,N_3903);
nor U4990 (N_4990,N_3741,N_3985);
xnor U4991 (N_4991,N_3904,N_3488);
nand U4992 (N_4992,N_3953,N_3452);
or U4993 (N_4993,N_3969,N_3980);
nand U4994 (N_4994,N_3513,N_3723);
xor U4995 (N_4995,N_3896,N_3110);
xor U4996 (N_4996,N_3967,N_3981);
nor U4997 (N_4997,N_3358,N_3309);
xnor U4998 (N_4998,N_3185,N_3736);
xnor U4999 (N_4999,N_3012,N_3540);
and UO_0 (O_0,N_4496,N_4046);
or UO_1 (O_1,N_4919,N_4832);
xnor UO_2 (O_2,N_4209,N_4129);
xor UO_3 (O_3,N_4284,N_4847);
and UO_4 (O_4,N_4225,N_4518);
nor UO_5 (O_5,N_4632,N_4493);
and UO_6 (O_6,N_4054,N_4727);
nor UO_7 (O_7,N_4611,N_4325);
or UO_8 (O_8,N_4636,N_4554);
xor UO_9 (O_9,N_4059,N_4675);
or UO_10 (O_10,N_4703,N_4365);
nor UO_11 (O_11,N_4689,N_4717);
nand UO_12 (O_12,N_4011,N_4126);
nand UO_13 (O_13,N_4634,N_4159);
and UO_14 (O_14,N_4378,N_4375);
or UO_15 (O_15,N_4094,N_4362);
or UO_16 (O_16,N_4440,N_4409);
nor UO_17 (O_17,N_4055,N_4733);
nor UO_18 (O_18,N_4737,N_4827);
nand UO_19 (O_19,N_4572,N_4565);
or UO_20 (O_20,N_4039,N_4594);
nand UO_21 (O_21,N_4937,N_4718);
and UO_22 (O_22,N_4665,N_4296);
nand UO_23 (O_23,N_4807,N_4122);
or UO_24 (O_24,N_4528,N_4691);
nand UO_25 (O_25,N_4941,N_4147);
and UO_26 (O_26,N_4647,N_4025);
xor UO_27 (O_27,N_4419,N_4512);
nand UO_28 (O_28,N_4970,N_4204);
xnor UO_29 (O_29,N_4006,N_4854);
xnor UO_30 (O_30,N_4692,N_4433);
nor UO_31 (O_31,N_4959,N_4875);
or UO_32 (O_32,N_4395,N_4598);
xnor UO_33 (O_33,N_4307,N_4868);
or UO_34 (O_34,N_4569,N_4196);
nor UO_35 (O_35,N_4627,N_4568);
or UO_36 (O_36,N_4228,N_4274);
xnor UO_37 (O_37,N_4774,N_4741);
nor UO_38 (O_38,N_4795,N_4547);
nand UO_39 (O_39,N_4803,N_4575);
xnor UO_40 (O_40,N_4898,N_4946);
nor UO_41 (O_41,N_4430,N_4294);
or UO_42 (O_42,N_4455,N_4157);
nor UO_43 (O_43,N_4182,N_4206);
nor UO_44 (O_44,N_4422,N_4109);
nand UO_45 (O_45,N_4155,N_4889);
and UO_46 (O_46,N_4527,N_4673);
nor UO_47 (O_47,N_4826,N_4071);
xnor UO_48 (O_48,N_4251,N_4498);
or UO_49 (O_49,N_4186,N_4887);
or UO_50 (O_50,N_4077,N_4616);
and UO_51 (O_51,N_4661,N_4404);
or UO_52 (O_52,N_4530,N_4885);
xor UO_53 (O_53,N_4957,N_4886);
nor UO_54 (O_54,N_4060,N_4269);
nand UO_55 (O_55,N_4825,N_4953);
and UO_56 (O_56,N_4470,N_4442);
xnor UO_57 (O_57,N_4163,N_4371);
nand UO_58 (O_58,N_4856,N_4949);
xnor UO_59 (O_59,N_4605,N_4858);
and UO_60 (O_60,N_4379,N_4050);
nor UO_61 (O_61,N_4845,N_4564);
nor UO_62 (O_62,N_4263,N_4456);
or UO_63 (O_63,N_4922,N_4870);
xor UO_64 (O_64,N_4292,N_4576);
or UO_65 (O_65,N_4821,N_4846);
or UO_66 (O_66,N_4863,N_4045);
and UO_67 (O_67,N_4747,N_4871);
or UO_68 (O_68,N_4955,N_4231);
nor UO_69 (O_69,N_4696,N_4043);
or UO_70 (O_70,N_4932,N_4893);
xor UO_71 (O_71,N_4763,N_4326);
nor UO_72 (O_72,N_4383,N_4694);
or UO_73 (O_73,N_4287,N_4698);
or UO_74 (O_74,N_4744,N_4766);
and UO_75 (O_75,N_4911,N_4002);
nor UO_76 (O_76,N_4264,N_4724);
or UO_77 (O_77,N_4116,N_4139);
xor UO_78 (O_78,N_4562,N_4024);
or UO_79 (O_79,N_4065,N_4981);
xor UO_80 (O_80,N_4161,N_4780);
nor UO_81 (O_81,N_4468,N_4393);
xnor UO_82 (O_82,N_4867,N_4786);
xor UO_83 (O_83,N_4872,N_4255);
and UO_84 (O_84,N_4464,N_4657);
or UO_85 (O_85,N_4349,N_4162);
nand UO_86 (O_86,N_4436,N_4978);
or UO_87 (O_87,N_4506,N_4303);
or UO_88 (O_88,N_4909,N_4034);
and UO_89 (O_89,N_4544,N_4708);
nand UO_90 (O_90,N_4093,N_4447);
or UO_91 (O_91,N_4335,N_4275);
or UO_92 (O_92,N_4824,N_4452);
nor UO_93 (O_93,N_4180,N_4902);
xnor UO_94 (O_94,N_4642,N_4352);
xnor UO_95 (O_95,N_4101,N_4535);
xor UO_96 (O_96,N_4646,N_4697);
nor UO_97 (O_97,N_4439,N_4449);
or UO_98 (O_98,N_4347,N_4167);
and UO_99 (O_99,N_4224,N_4521);
or UO_100 (O_100,N_4441,N_4991);
nor UO_101 (O_101,N_4629,N_4551);
xor UO_102 (O_102,N_4876,N_4009);
or UO_103 (O_103,N_4604,N_4019);
nor UO_104 (O_104,N_4390,N_4380);
nand UO_105 (O_105,N_4382,N_4731);
nand UO_106 (O_106,N_4138,N_4150);
nand UO_107 (O_107,N_4654,N_4202);
xnor UO_108 (O_108,N_4467,N_4730);
or UO_109 (O_109,N_4450,N_4534);
or UO_110 (O_110,N_4295,N_4492);
nor UO_111 (O_111,N_4877,N_4631);
xor UO_112 (O_112,N_4980,N_4189);
and UO_113 (O_113,N_4427,N_4280);
xnor UO_114 (O_114,N_4338,N_4341);
nand UO_115 (O_115,N_4505,N_4324);
xnor UO_116 (O_116,N_4644,N_4448);
or UO_117 (O_117,N_4557,N_4223);
and UO_118 (O_118,N_4394,N_4205);
xnor UO_119 (O_119,N_4706,N_4148);
and UO_120 (O_120,N_4879,N_4884);
nand UO_121 (O_121,N_4805,N_4705);
or UO_122 (O_122,N_4235,N_4811);
and UO_123 (O_123,N_4855,N_4250);
nor UO_124 (O_124,N_4735,N_4729);
nor UO_125 (O_125,N_4415,N_4773);
nand UO_126 (O_126,N_4023,N_4587);
nor UO_127 (O_127,N_4517,N_4291);
and UO_128 (O_128,N_4089,N_4012);
xor UO_129 (O_129,N_4286,N_4169);
xnor UO_130 (O_130,N_4712,N_4482);
xor UO_131 (O_131,N_4110,N_4866);
nor UO_132 (O_132,N_4972,N_4686);
xor UO_133 (O_133,N_4154,N_4016);
and UO_134 (O_134,N_4796,N_4750);
nand UO_135 (O_135,N_4105,N_4925);
nor UO_136 (O_136,N_4305,N_4072);
nand UO_137 (O_137,N_4031,N_4038);
or UO_138 (O_138,N_4745,N_4004);
nand UO_139 (O_139,N_4342,N_4860);
nand UO_140 (O_140,N_4074,N_4090);
xnor UO_141 (O_141,N_4082,N_4222);
and UO_142 (O_142,N_4999,N_4923);
nand UO_143 (O_143,N_4620,N_4471);
nand UO_144 (O_144,N_4797,N_4302);
and UO_145 (O_145,N_4571,N_4080);
nor UO_146 (O_146,N_4670,N_4556);
or UO_147 (O_147,N_4668,N_4314);
or UO_148 (O_148,N_4865,N_4309);
and UO_149 (O_149,N_4172,N_4483);
and UO_150 (O_150,N_4903,N_4906);
nand UO_151 (O_151,N_4160,N_4293);
xor UO_152 (O_152,N_4348,N_4794);
or UO_153 (O_153,N_4707,N_4974);
and UO_154 (O_154,N_4332,N_4713);
nand UO_155 (O_155,N_4850,N_4883);
xnor UO_156 (O_156,N_4133,N_4244);
or UO_157 (O_157,N_4986,N_4954);
or UO_158 (O_158,N_4823,N_4297);
or UO_159 (O_159,N_4299,N_4306);
nor UO_160 (O_160,N_4641,N_4520);
and UO_161 (O_161,N_4486,N_4005);
and UO_162 (O_162,N_4915,N_4835);
nand UO_163 (O_163,N_4234,N_4951);
or UO_164 (O_164,N_4385,N_4767);
xnor UO_165 (O_165,N_4056,N_4036);
or UO_166 (O_166,N_4519,N_4555);
nor UO_167 (O_167,N_4366,N_4892);
and UO_168 (O_168,N_4330,N_4920);
and UO_169 (O_169,N_4831,N_4201);
or UO_170 (O_170,N_4621,N_4400);
or UO_171 (O_171,N_4660,N_4114);
xor UO_172 (O_172,N_4873,N_4128);
nor UO_173 (O_173,N_4630,N_4804);
xor UO_174 (O_174,N_4355,N_4061);
or UO_175 (O_175,N_4663,N_4104);
nor UO_176 (O_176,N_4316,N_4064);
or UO_177 (O_177,N_4282,N_4417);
or UO_178 (O_178,N_4788,N_4523);
or UO_179 (O_179,N_4402,N_4364);
or UO_180 (O_180,N_4754,N_4221);
or UO_181 (O_181,N_4240,N_4232);
nand UO_182 (O_182,N_4115,N_4158);
nand UO_183 (O_183,N_4762,N_4494);
nand UO_184 (O_184,N_4757,N_4559);
xor UO_185 (O_185,N_4723,N_4117);
nand UO_186 (O_186,N_4934,N_4929);
nor UO_187 (O_187,N_4136,N_4853);
xor UO_188 (O_188,N_4022,N_4177);
and UO_189 (O_189,N_4431,N_4103);
nor UO_190 (O_190,N_4210,N_4288);
xnor UO_191 (O_191,N_4833,N_4687);
or UO_192 (O_192,N_4709,N_4588);
xor UO_193 (O_193,N_4398,N_4843);
or UO_194 (O_194,N_4121,N_4361);
or UO_195 (O_195,N_4191,N_4168);
nor UO_196 (O_196,N_4253,N_4720);
nand UO_197 (O_197,N_4507,N_4830);
nor UO_198 (O_198,N_4049,N_4198);
xnor UO_199 (O_199,N_4127,N_4514);
xnor UO_200 (O_200,N_4683,N_4944);
and UO_201 (O_201,N_4451,N_4770);
nor UO_202 (O_202,N_4042,N_4053);
nand UO_203 (O_203,N_4239,N_4216);
and UO_204 (O_204,N_4227,N_4533);
or UO_205 (O_205,N_4051,N_4541);
nor UO_206 (O_206,N_4472,N_4891);
nor UO_207 (O_207,N_4271,N_4617);
or UO_208 (O_208,N_4078,N_4693);
nand UO_209 (O_209,N_4539,N_4372);
or UO_210 (O_210,N_4553,N_4597);
and UO_211 (O_211,N_4118,N_4401);
xnor UO_212 (O_212,N_4685,N_4552);
xnor UO_213 (O_213,N_4261,N_4279);
nand UO_214 (O_214,N_4041,N_4258);
and UO_215 (O_215,N_4021,N_4376);
or UO_216 (O_216,N_4392,N_4268);
xnor UO_217 (O_217,N_4503,N_4443);
nand UO_218 (O_218,N_4246,N_4752);
or UO_219 (O_219,N_4580,N_4839);
or UO_220 (O_220,N_4236,N_4195);
xnor UO_221 (O_221,N_4008,N_4312);
nand UO_222 (O_222,N_4680,N_4298);
xnor UO_223 (O_223,N_4396,N_4940);
and UO_224 (O_224,N_4537,N_4146);
or UO_225 (O_225,N_4912,N_4622);
and UO_226 (O_226,N_4397,N_4732);
and UO_227 (O_227,N_4655,N_4548);
xor UO_228 (O_228,N_4311,N_4181);
nand UO_229 (O_229,N_4200,N_4781);
and UO_230 (O_230,N_4098,N_4124);
nand UO_231 (O_231,N_4817,N_4600);
nor UO_232 (O_232,N_4852,N_4926);
nand UO_233 (O_233,N_4910,N_4350);
nand UO_234 (O_234,N_4070,N_4319);
xor UO_235 (O_235,N_4207,N_4377);
xnor UO_236 (O_236,N_4682,N_4131);
nand UO_237 (O_237,N_4414,N_4585);
or UO_238 (O_238,N_4984,N_4097);
and UO_239 (O_239,N_4017,N_4841);
or UO_240 (O_240,N_4895,N_4462);
xor UO_241 (O_241,N_4990,N_4194);
or UO_242 (O_242,N_4864,N_4029);
xnor UO_243 (O_243,N_4649,N_4982);
nor UO_244 (O_244,N_4849,N_4466);
or UO_245 (O_245,N_4413,N_4609);
or UO_246 (O_246,N_4501,N_4272);
or UO_247 (O_247,N_4453,N_4339);
nor UO_248 (O_248,N_4119,N_4679);
or UO_249 (O_249,N_4259,N_4578);
xor UO_250 (O_250,N_4775,N_4187);
and UO_251 (O_251,N_4882,N_4476);
or UO_252 (O_252,N_4896,N_4595);
or UO_253 (O_253,N_4549,N_4862);
xor UO_254 (O_254,N_4593,N_4715);
xnor UO_255 (O_255,N_4120,N_4701);
nor UO_256 (O_256,N_4488,N_4928);
nor UO_257 (O_257,N_4360,N_4894);
xor UO_258 (O_258,N_4151,N_4249);
nand UO_259 (O_259,N_4418,N_4123);
nand UO_260 (O_260,N_4966,N_4844);
xnor UO_261 (O_261,N_4596,N_4048);
xnor UO_262 (O_262,N_4057,N_4145);
nor UO_263 (O_263,N_4897,N_4459);
or UO_264 (O_264,N_4226,N_4818);
or UO_265 (O_265,N_4522,N_4574);
xnor UO_266 (O_266,N_4545,N_4810);
nor UO_267 (O_267,N_4676,N_4822);
and UO_268 (O_268,N_4538,N_4516);
nand UO_269 (O_269,N_4407,N_4277);
and UO_270 (O_270,N_4344,N_4434);
and UO_271 (O_271,N_4058,N_4076);
nor UO_272 (O_272,N_4607,N_4997);
nand UO_273 (O_273,N_4267,N_4370);
or UO_274 (O_274,N_4323,N_4003);
and UO_275 (O_275,N_4814,N_4812);
nand UO_276 (O_276,N_4586,N_4658);
xnor UO_277 (O_277,N_4589,N_4423);
or UO_278 (O_278,N_4710,N_4608);
and UO_279 (O_279,N_4285,N_4721);
nand UO_280 (O_280,N_4343,N_4113);
nor UO_281 (O_281,N_4432,N_4052);
or UO_282 (O_282,N_4753,N_4142);
and UO_283 (O_283,N_4230,N_4792);
or UO_284 (O_284,N_4170,N_4075);
nand UO_285 (O_285,N_4478,N_4315);
or UO_286 (O_286,N_4577,N_4363);
or UO_287 (O_287,N_4933,N_4211);
nor UO_288 (O_288,N_4640,N_4469);
nand UO_289 (O_289,N_4973,N_4664);
or UO_290 (O_290,N_4977,N_4130);
and UO_291 (O_291,N_4878,N_4612);
or UO_292 (O_292,N_4386,N_4270);
and UO_293 (O_293,N_4066,N_4965);
xor UO_294 (O_294,N_4426,N_4531);
xor UO_295 (O_295,N_4579,N_4681);
xnor UO_296 (O_296,N_4489,N_4214);
or UO_297 (O_297,N_4874,N_4975);
or UO_298 (O_298,N_4958,N_4667);
and UO_299 (O_299,N_4633,N_4678);
and UO_300 (O_300,N_4152,N_4495);
xnor UO_301 (O_301,N_4725,N_4190);
xor UO_302 (O_302,N_4592,N_4337);
nand UO_303 (O_303,N_4801,N_4704);
or UO_304 (O_304,N_4789,N_4816);
or UO_305 (O_305,N_4582,N_4083);
and UO_306 (O_306,N_4790,N_4178);
and UO_307 (O_307,N_4281,N_4081);
or UO_308 (O_308,N_4857,N_4917);
or UO_309 (O_309,N_4477,N_4027);
and UO_310 (O_310,N_4765,N_4618);
nand UO_311 (O_311,N_4111,N_4444);
xor UO_312 (O_312,N_4635,N_4387);
nand UO_313 (O_313,N_4748,N_4106);
nor UO_314 (O_314,N_4719,N_4174);
and UO_315 (O_315,N_4650,N_4963);
nand UO_316 (O_316,N_4907,N_4914);
and UO_317 (O_317,N_4425,N_4799);
or UO_318 (O_318,N_4809,N_4626);
xor UO_319 (O_319,N_4782,N_4173);
nor UO_320 (O_320,N_4695,N_4329);
nand UO_321 (O_321,N_4784,N_4610);
nand UO_322 (O_322,N_4688,N_4952);
nand UO_323 (O_323,N_4840,N_4546);
and UO_324 (O_324,N_4384,N_4904);
and UO_325 (O_325,N_4930,N_4219);
nor UO_326 (O_326,N_4563,N_4987);
and UO_327 (O_327,N_4671,N_4308);
nand UO_328 (O_328,N_4497,N_4445);
or UO_329 (O_329,N_4761,N_4751);
xnor UO_330 (O_330,N_4156,N_4073);
and UO_331 (O_331,N_4192,N_4399);
and UO_332 (O_332,N_4838,N_4095);
nor UO_333 (O_333,N_4345,N_4842);
nand UO_334 (O_334,N_4229,N_4581);
nand UO_335 (O_335,N_4273,N_4561);
nand UO_336 (O_336,N_4651,N_4573);
nor UO_337 (O_337,N_4599,N_4096);
nor UO_338 (O_338,N_4143,N_4331);
nand UO_339 (O_339,N_4026,N_4550);
and UO_340 (O_340,N_4254,N_4916);
or UO_341 (O_341,N_4032,N_4743);
and UO_342 (O_342,N_4102,N_4989);
nor UO_343 (O_343,N_4524,N_4726);
and UO_344 (O_344,N_4995,N_4346);
nor UO_345 (O_345,N_4416,N_4092);
nand UO_346 (O_346,N_4403,N_4764);
nand UO_347 (O_347,N_4834,N_4067);
nand UO_348 (O_348,N_4357,N_4480);
nand UO_349 (O_349,N_4746,N_4890);
and UO_350 (O_350,N_4458,N_4457);
xnor UO_351 (O_351,N_4526,N_4310);
nand UO_352 (O_352,N_4406,N_4939);
or UO_353 (O_353,N_4241,N_4491);
xnor UO_354 (O_354,N_4962,N_4590);
nor UO_355 (O_355,N_4772,N_4233);
xor UO_356 (O_356,N_4736,N_4454);
nand UO_357 (O_357,N_4313,N_4243);
nand UO_358 (O_358,N_4791,N_4602);
and UO_359 (O_359,N_4567,N_4193);
xnor UO_360 (O_360,N_4669,N_4945);
or UO_361 (O_361,N_4013,N_4601);
nand UO_362 (O_362,N_4769,N_4125);
nand UO_363 (O_363,N_4742,N_4921);
nand UO_364 (O_364,N_4188,N_4529);
and UO_365 (O_365,N_4513,N_4508);
xnor UO_366 (O_366,N_4583,N_4321);
or UO_367 (O_367,N_4829,N_4499);
and UO_368 (O_368,N_4322,N_4040);
and UO_369 (O_369,N_4475,N_4820);
or UO_370 (O_370,N_4802,N_4135);
nand UO_371 (O_371,N_4936,N_4359);
or UO_372 (O_372,N_4779,N_4994);
xnor UO_373 (O_373,N_4619,N_4532);
or UO_374 (O_374,N_4652,N_4428);
nand UO_375 (O_375,N_4044,N_4461);
xor UO_376 (O_376,N_4213,N_4639);
and UO_377 (O_377,N_4108,N_4134);
and UO_378 (O_378,N_4484,N_4301);
nand UO_379 (O_379,N_4711,N_4373);
and UO_380 (O_380,N_4446,N_4938);
nor UO_381 (O_381,N_4935,N_4140);
or UO_382 (O_382,N_4179,N_4672);
or UO_383 (O_383,N_4030,N_4424);
nand UO_384 (O_384,N_4199,N_4100);
nand UO_385 (O_385,N_4327,N_4502);
nor UO_386 (O_386,N_4785,N_4351);
and UO_387 (O_387,N_4768,N_4252);
and UO_388 (O_388,N_4317,N_4215);
xnor UO_389 (O_389,N_4086,N_4778);
xor UO_390 (O_390,N_4175,N_4388);
and UO_391 (O_391,N_4353,N_4808);
xnor UO_392 (O_392,N_4988,N_4540);
and UO_393 (O_393,N_4410,N_4624);
nor UO_394 (O_394,N_4653,N_4197);
nand UO_395 (O_395,N_4389,N_4684);
nor UO_396 (O_396,N_4289,N_4956);
nor UO_397 (O_397,N_4776,N_4141);
nand UO_398 (O_398,N_4437,N_4460);
nand UO_399 (O_399,N_4405,N_4656);
or UO_400 (O_400,N_4218,N_4212);
and UO_401 (O_401,N_4381,N_4047);
xor UO_402 (O_402,N_4429,N_4908);
or UO_403 (O_403,N_4993,N_4001);
nor UO_404 (O_404,N_4165,N_4515);
nor UO_405 (O_405,N_4543,N_4290);
nand UO_406 (O_406,N_4511,N_4968);
nand UO_407 (O_407,N_4421,N_4144);
and UO_408 (O_408,N_4828,N_4690);
nand UO_409 (O_409,N_4777,N_4967);
nand UO_410 (O_410,N_4237,N_4248);
or UO_411 (O_411,N_4334,N_4570);
nand UO_412 (O_412,N_4560,N_4033);
nor UO_413 (O_413,N_4755,N_4037);
or UO_414 (O_414,N_4203,N_4340);
nand UO_415 (O_415,N_4463,N_4943);
nand UO_416 (O_416,N_4411,N_4806);
nor UO_417 (O_417,N_4132,N_4913);
and UO_418 (O_418,N_4931,N_4606);
nand UO_419 (O_419,N_4948,N_4759);
or UO_420 (O_420,N_4185,N_4176);
xor UO_421 (O_421,N_4510,N_4961);
and UO_422 (O_422,N_4015,N_4674);
and UO_423 (O_423,N_4623,N_4659);
xnor UO_424 (O_424,N_4412,N_4500);
or UO_425 (O_425,N_4566,N_4479);
or UO_426 (O_426,N_4542,N_4473);
or UO_427 (O_427,N_4000,N_4740);
nand UO_428 (O_428,N_4088,N_4739);
or UO_429 (O_429,N_4063,N_4242);
and UO_430 (O_430,N_4408,N_4615);
and UO_431 (O_431,N_4899,N_4525);
and UO_432 (O_432,N_4354,N_4262);
nor UO_433 (O_433,N_4699,N_4591);
and UO_434 (O_434,N_4278,N_4010);
and UO_435 (O_435,N_4260,N_4584);
or UO_436 (O_436,N_4628,N_4485);
xnor UO_437 (O_437,N_4558,N_4998);
nor UO_438 (O_438,N_4771,N_4979);
or UO_439 (O_439,N_4734,N_4256);
nand UO_440 (O_440,N_4880,N_4356);
and UO_441 (O_441,N_4783,N_4099);
and UO_442 (O_442,N_4300,N_4819);
or UO_443 (O_443,N_4662,N_4881);
nor UO_444 (O_444,N_4836,N_4068);
nand UO_445 (O_445,N_4018,N_4069);
or UO_446 (O_446,N_4062,N_4677);
nor UO_447 (O_447,N_4374,N_4815);
and UO_448 (O_448,N_4798,N_4166);
nor UO_449 (O_449,N_4787,N_4112);
xor UO_450 (O_450,N_4079,N_4369);
nand UO_451 (O_451,N_4217,N_4666);
or UO_452 (O_452,N_4333,N_4265);
or UO_453 (O_453,N_4487,N_4869);
and UO_454 (O_454,N_4481,N_4391);
xor UO_455 (O_455,N_4020,N_4028);
or UO_456 (O_456,N_4851,N_4367);
nand UO_457 (O_457,N_4368,N_4184);
or UO_458 (O_458,N_4942,N_4304);
xor UO_459 (O_459,N_4220,N_4861);
and UO_460 (O_460,N_4318,N_4465);
xor UO_461 (O_461,N_4714,N_4245);
nor UO_462 (O_462,N_4837,N_4107);
and UO_463 (O_463,N_4964,N_4971);
nand UO_464 (O_464,N_4438,N_4085);
or UO_465 (O_465,N_4960,N_4625);
nor UO_466 (O_466,N_4700,N_4336);
or UO_467 (O_467,N_4183,N_4283);
xor UO_468 (O_468,N_4613,N_4638);
xnor UO_469 (O_469,N_4760,N_4490);
xnor UO_470 (O_470,N_4257,N_4950);
nor UO_471 (O_471,N_4996,N_4084);
xor UO_472 (O_472,N_4648,N_4149);
and UO_473 (O_473,N_4645,N_4976);
or UO_474 (O_474,N_4164,N_4983);
and UO_475 (O_475,N_4992,N_4536);
nor UO_476 (O_476,N_4509,N_4171);
and UO_477 (O_477,N_4924,N_4927);
xnor UO_478 (O_478,N_4153,N_4137);
xor UO_479 (O_479,N_4756,N_4728);
xor UO_480 (O_480,N_4328,N_4320);
or UO_481 (O_481,N_4643,N_4800);
nand UO_482 (O_482,N_4900,N_4266);
or UO_483 (O_483,N_4888,N_4007);
xor UO_484 (O_484,N_4358,N_4969);
nor UO_485 (O_485,N_4603,N_4985);
xor UO_486 (O_486,N_4014,N_4813);
and UO_487 (O_487,N_4208,N_4702);
xnor UO_488 (O_488,N_4238,N_4087);
nor UO_489 (O_489,N_4637,N_4716);
or UO_490 (O_490,N_4474,N_4947);
nand UO_491 (O_491,N_4504,N_4905);
xor UO_492 (O_492,N_4722,N_4793);
and UO_493 (O_493,N_4614,N_4859);
nor UO_494 (O_494,N_4901,N_4091);
and UO_495 (O_495,N_4420,N_4035);
or UO_496 (O_496,N_4758,N_4247);
or UO_497 (O_497,N_4918,N_4276);
or UO_498 (O_498,N_4435,N_4738);
nand UO_499 (O_499,N_4848,N_4749);
xnor UO_500 (O_500,N_4927,N_4739);
and UO_501 (O_501,N_4804,N_4050);
xor UO_502 (O_502,N_4227,N_4911);
and UO_503 (O_503,N_4616,N_4355);
and UO_504 (O_504,N_4747,N_4335);
nand UO_505 (O_505,N_4686,N_4802);
nand UO_506 (O_506,N_4401,N_4177);
nand UO_507 (O_507,N_4376,N_4285);
nor UO_508 (O_508,N_4575,N_4925);
nand UO_509 (O_509,N_4887,N_4294);
nor UO_510 (O_510,N_4500,N_4526);
nor UO_511 (O_511,N_4633,N_4088);
nor UO_512 (O_512,N_4596,N_4210);
xnor UO_513 (O_513,N_4783,N_4628);
or UO_514 (O_514,N_4614,N_4513);
nor UO_515 (O_515,N_4315,N_4611);
nor UO_516 (O_516,N_4676,N_4671);
nor UO_517 (O_517,N_4444,N_4665);
xor UO_518 (O_518,N_4649,N_4363);
nor UO_519 (O_519,N_4548,N_4714);
nor UO_520 (O_520,N_4029,N_4673);
xnor UO_521 (O_521,N_4398,N_4538);
and UO_522 (O_522,N_4057,N_4859);
xor UO_523 (O_523,N_4893,N_4650);
nor UO_524 (O_524,N_4326,N_4058);
nor UO_525 (O_525,N_4511,N_4338);
nand UO_526 (O_526,N_4192,N_4311);
or UO_527 (O_527,N_4052,N_4428);
xor UO_528 (O_528,N_4563,N_4568);
or UO_529 (O_529,N_4625,N_4544);
nand UO_530 (O_530,N_4402,N_4791);
xor UO_531 (O_531,N_4464,N_4196);
xor UO_532 (O_532,N_4072,N_4999);
xor UO_533 (O_533,N_4419,N_4881);
nor UO_534 (O_534,N_4468,N_4615);
or UO_535 (O_535,N_4249,N_4714);
nor UO_536 (O_536,N_4909,N_4378);
nor UO_537 (O_537,N_4786,N_4861);
nand UO_538 (O_538,N_4878,N_4643);
xnor UO_539 (O_539,N_4737,N_4002);
xnor UO_540 (O_540,N_4375,N_4847);
nand UO_541 (O_541,N_4913,N_4210);
and UO_542 (O_542,N_4693,N_4122);
and UO_543 (O_543,N_4624,N_4760);
and UO_544 (O_544,N_4220,N_4885);
and UO_545 (O_545,N_4733,N_4215);
nand UO_546 (O_546,N_4678,N_4884);
xnor UO_547 (O_547,N_4949,N_4052);
nor UO_548 (O_548,N_4537,N_4143);
xnor UO_549 (O_549,N_4432,N_4985);
and UO_550 (O_550,N_4426,N_4081);
or UO_551 (O_551,N_4224,N_4096);
and UO_552 (O_552,N_4779,N_4910);
nand UO_553 (O_553,N_4296,N_4904);
nand UO_554 (O_554,N_4485,N_4220);
and UO_555 (O_555,N_4298,N_4217);
nor UO_556 (O_556,N_4511,N_4655);
or UO_557 (O_557,N_4660,N_4596);
xor UO_558 (O_558,N_4397,N_4660);
or UO_559 (O_559,N_4624,N_4843);
xor UO_560 (O_560,N_4841,N_4218);
and UO_561 (O_561,N_4263,N_4634);
xor UO_562 (O_562,N_4038,N_4101);
xor UO_563 (O_563,N_4105,N_4170);
nor UO_564 (O_564,N_4860,N_4865);
nor UO_565 (O_565,N_4327,N_4249);
xor UO_566 (O_566,N_4877,N_4257);
xnor UO_567 (O_567,N_4718,N_4807);
and UO_568 (O_568,N_4084,N_4628);
xor UO_569 (O_569,N_4891,N_4671);
or UO_570 (O_570,N_4314,N_4790);
xnor UO_571 (O_571,N_4800,N_4935);
and UO_572 (O_572,N_4594,N_4396);
nor UO_573 (O_573,N_4823,N_4339);
or UO_574 (O_574,N_4668,N_4604);
nor UO_575 (O_575,N_4464,N_4702);
xor UO_576 (O_576,N_4606,N_4018);
xnor UO_577 (O_577,N_4606,N_4141);
or UO_578 (O_578,N_4522,N_4620);
xor UO_579 (O_579,N_4447,N_4995);
or UO_580 (O_580,N_4045,N_4980);
xnor UO_581 (O_581,N_4090,N_4660);
or UO_582 (O_582,N_4289,N_4227);
xor UO_583 (O_583,N_4320,N_4225);
and UO_584 (O_584,N_4291,N_4759);
or UO_585 (O_585,N_4933,N_4579);
nor UO_586 (O_586,N_4510,N_4281);
and UO_587 (O_587,N_4776,N_4372);
and UO_588 (O_588,N_4847,N_4894);
or UO_589 (O_589,N_4472,N_4162);
xnor UO_590 (O_590,N_4620,N_4598);
and UO_591 (O_591,N_4505,N_4922);
xor UO_592 (O_592,N_4105,N_4751);
nor UO_593 (O_593,N_4836,N_4175);
nor UO_594 (O_594,N_4078,N_4931);
or UO_595 (O_595,N_4014,N_4791);
and UO_596 (O_596,N_4467,N_4343);
and UO_597 (O_597,N_4414,N_4566);
nor UO_598 (O_598,N_4963,N_4291);
nor UO_599 (O_599,N_4961,N_4043);
and UO_600 (O_600,N_4218,N_4743);
nand UO_601 (O_601,N_4723,N_4440);
nand UO_602 (O_602,N_4370,N_4385);
nor UO_603 (O_603,N_4179,N_4226);
nand UO_604 (O_604,N_4582,N_4173);
nor UO_605 (O_605,N_4531,N_4109);
nand UO_606 (O_606,N_4234,N_4286);
xor UO_607 (O_607,N_4145,N_4883);
nand UO_608 (O_608,N_4104,N_4410);
xnor UO_609 (O_609,N_4870,N_4343);
or UO_610 (O_610,N_4585,N_4451);
nor UO_611 (O_611,N_4551,N_4976);
nor UO_612 (O_612,N_4119,N_4144);
or UO_613 (O_613,N_4986,N_4304);
nand UO_614 (O_614,N_4226,N_4488);
and UO_615 (O_615,N_4716,N_4001);
and UO_616 (O_616,N_4960,N_4449);
nand UO_617 (O_617,N_4100,N_4069);
xor UO_618 (O_618,N_4478,N_4328);
or UO_619 (O_619,N_4397,N_4867);
and UO_620 (O_620,N_4610,N_4783);
nor UO_621 (O_621,N_4668,N_4560);
or UO_622 (O_622,N_4735,N_4962);
nand UO_623 (O_623,N_4009,N_4726);
nor UO_624 (O_624,N_4218,N_4162);
and UO_625 (O_625,N_4352,N_4132);
nand UO_626 (O_626,N_4817,N_4011);
nand UO_627 (O_627,N_4478,N_4452);
xnor UO_628 (O_628,N_4282,N_4574);
nor UO_629 (O_629,N_4039,N_4969);
or UO_630 (O_630,N_4489,N_4947);
or UO_631 (O_631,N_4434,N_4072);
xor UO_632 (O_632,N_4404,N_4054);
or UO_633 (O_633,N_4238,N_4275);
xor UO_634 (O_634,N_4918,N_4755);
and UO_635 (O_635,N_4783,N_4933);
nand UO_636 (O_636,N_4409,N_4979);
xnor UO_637 (O_637,N_4954,N_4575);
or UO_638 (O_638,N_4827,N_4235);
or UO_639 (O_639,N_4187,N_4252);
or UO_640 (O_640,N_4410,N_4323);
nand UO_641 (O_641,N_4255,N_4710);
nand UO_642 (O_642,N_4059,N_4131);
or UO_643 (O_643,N_4107,N_4931);
nand UO_644 (O_644,N_4458,N_4073);
nor UO_645 (O_645,N_4012,N_4336);
and UO_646 (O_646,N_4912,N_4676);
or UO_647 (O_647,N_4365,N_4976);
nand UO_648 (O_648,N_4616,N_4499);
and UO_649 (O_649,N_4607,N_4147);
nor UO_650 (O_650,N_4952,N_4747);
or UO_651 (O_651,N_4862,N_4411);
xnor UO_652 (O_652,N_4308,N_4266);
nor UO_653 (O_653,N_4188,N_4577);
xnor UO_654 (O_654,N_4872,N_4573);
xnor UO_655 (O_655,N_4626,N_4305);
or UO_656 (O_656,N_4504,N_4521);
xor UO_657 (O_657,N_4389,N_4896);
nor UO_658 (O_658,N_4363,N_4179);
xnor UO_659 (O_659,N_4089,N_4119);
nand UO_660 (O_660,N_4132,N_4259);
xnor UO_661 (O_661,N_4406,N_4194);
or UO_662 (O_662,N_4293,N_4987);
xor UO_663 (O_663,N_4059,N_4301);
xnor UO_664 (O_664,N_4575,N_4812);
xor UO_665 (O_665,N_4086,N_4606);
xor UO_666 (O_666,N_4580,N_4467);
xnor UO_667 (O_667,N_4981,N_4150);
or UO_668 (O_668,N_4068,N_4350);
xor UO_669 (O_669,N_4076,N_4825);
xor UO_670 (O_670,N_4526,N_4449);
nor UO_671 (O_671,N_4876,N_4566);
nor UO_672 (O_672,N_4755,N_4097);
and UO_673 (O_673,N_4832,N_4950);
or UO_674 (O_674,N_4671,N_4539);
nand UO_675 (O_675,N_4020,N_4119);
and UO_676 (O_676,N_4178,N_4317);
nor UO_677 (O_677,N_4756,N_4008);
or UO_678 (O_678,N_4020,N_4888);
xor UO_679 (O_679,N_4515,N_4915);
nand UO_680 (O_680,N_4063,N_4610);
or UO_681 (O_681,N_4799,N_4007);
nand UO_682 (O_682,N_4516,N_4062);
and UO_683 (O_683,N_4441,N_4174);
nor UO_684 (O_684,N_4086,N_4928);
and UO_685 (O_685,N_4864,N_4186);
xnor UO_686 (O_686,N_4866,N_4947);
nor UO_687 (O_687,N_4539,N_4177);
or UO_688 (O_688,N_4113,N_4012);
xnor UO_689 (O_689,N_4625,N_4630);
xor UO_690 (O_690,N_4096,N_4745);
and UO_691 (O_691,N_4589,N_4309);
nand UO_692 (O_692,N_4621,N_4443);
and UO_693 (O_693,N_4732,N_4110);
xor UO_694 (O_694,N_4571,N_4932);
xor UO_695 (O_695,N_4515,N_4577);
xor UO_696 (O_696,N_4736,N_4552);
and UO_697 (O_697,N_4083,N_4700);
xnor UO_698 (O_698,N_4847,N_4102);
nor UO_699 (O_699,N_4113,N_4065);
nand UO_700 (O_700,N_4076,N_4293);
nand UO_701 (O_701,N_4849,N_4391);
and UO_702 (O_702,N_4253,N_4482);
or UO_703 (O_703,N_4408,N_4519);
or UO_704 (O_704,N_4776,N_4120);
or UO_705 (O_705,N_4486,N_4019);
xnor UO_706 (O_706,N_4323,N_4919);
xor UO_707 (O_707,N_4112,N_4577);
and UO_708 (O_708,N_4861,N_4606);
and UO_709 (O_709,N_4304,N_4130);
nand UO_710 (O_710,N_4866,N_4612);
nand UO_711 (O_711,N_4117,N_4419);
xor UO_712 (O_712,N_4057,N_4628);
and UO_713 (O_713,N_4825,N_4744);
nor UO_714 (O_714,N_4517,N_4452);
xnor UO_715 (O_715,N_4847,N_4546);
and UO_716 (O_716,N_4141,N_4901);
or UO_717 (O_717,N_4457,N_4043);
nor UO_718 (O_718,N_4769,N_4176);
nor UO_719 (O_719,N_4314,N_4311);
nor UO_720 (O_720,N_4989,N_4719);
nor UO_721 (O_721,N_4555,N_4640);
and UO_722 (O_722,N_4527,N_4489);
nor UO_723 (O_723,N_4331,N_4879);
or UO_724 (O_724,N_4992,N_4358);
and UO_725 (O_725,N_4567,N_4810);
xnor UO_726 (O_726,N_4156,N_4400);
or UO_727 (O_727,N_4656,N_4014);
or UO_728 (O_728,N_4662,N_4161);
nand UO_729 (O_729,N_4052,N_4009);
xnor UO_730 (O_730,N_4869,N_4884);
nand UO_731 (O_731,N_4510,N_4652);
nand UO_732 (O_732,N_4924,N_4408);
nand UO_733 (O_733,N_4053,N_4480);
nor UO_734 (O_734,N_4694,N_4427);
nor UO_735 (O_735,N_4400,N_4106);
and UO_736 (O_736,N_4905,N_4922);
xor UO_737 (O_737,N_4782,N_4701);
nor UO_738 (O_738,N_4818,N_4328);
xnor UO_739 (O_739,N_4985,N_4103);
nand UO_740 (O_740,N_4276,N_4702);
and UO_741 (O_741,N_4308,N_4658);
nor UO_742 (O_742,N_4795,N_4596);
nor UO_743 (O_743,N_4469,N_4583);
and UO_744 (O_744,N_4142,N_4127);
nand UO_745 (O_745,N_4481,N_4697);
nand UO_746 (O_746,N_4669,N_4705);
xnor UO_747 (O_747,N_4268,N_4349);
and UO_748 (O_748,N_4036,N_4518);
nand UO_749 (O_749,N_4999,N_4860);
nand UO_750 (O_750,N_4755,N_4153);
xnor UO_751 (O_751,N_4403,N_4397);
xnor UO_752 (O_752,N_4323,N_4490);
and UO_753 (O_753,N_4159,N_4374);
and UO_754 (O_754,N_4245,N_4283);
nor UO_755 (O_755,N_4753,N_4466);
nor UO_756 (O_756,N_4246,N_4794);
nand UO_757 (O_757,N_4812,N_4918);
and UO_758 (O_758,N_4282,N_4498);
or UO_759 (O_759,N_4245,N_4040);
or UO_760 (O_760,N_4681,N_4813);
nor UO_761 (O_761,N_4555,N_4887);
or UO_762 (O_762,N_4603,N_4466);
nor UO_763 (O_763,N_4403,N_4195);
xnor UO_764 (O_764,N_4600,N_4449);
xnor UO_765 (O_765,N_4058,N_4859);
xnor UO_766 (O_766,N_4702,N_4674);
or UO_767 (O_767,N_4443,N_4499);
nand UO_768 (O_768,N_4826,N_4852);
nor UO_769 (O_769,N_4184,N_4162);
xor UO_770 (O_770,N_4974,N_4929);
nand UO_771 (O_771,N_4106,N_4253);
xnor UO_772 (O_772,N_4094,N_4743);
nand UO_773 (O_773,N_4087,N_4255);
nor UO_774 (O_774,N_4879,N_4866);
nor UO_775 (O_775,N_4168,N_4894);
and UO_776 (O_776,N_4091,N_4163);
nand UO_777 (O_777,N_4989,N_4059);
nand UO_778 (O_778,N_4775,N_4549);
xnor UO_779 (O_779,N_4218,N_4977);
xor UO_780 (O_780,N_4626,N_4736);
and UO_781 (O_781,N_4152,N_4553);
nor UO_782 (O_782,N_4496,N_4984);
nand UO_783 (O_783,N_4528,N_4699);
or UO_784 (O_784,N_4323,N_4096);
nand UO_785 (O_785,N_4283,N_4678);
nand UO_786 (O_786,N_4377,N_4264);
xor UO_787 (O_787,N_4921,N_4270);
nand UO_788 (O_788,N_4083,N_4208);
xor UO_789 (O_789,N_4187,N_4877);
nor UO_790 (O_790,N_4552,N_4154);
or UO_791 (O_791,N_4488,N_4263);
nor UO_792 (O_792,N_4761,N_4703);
nand UO_793 (O_793,N_4657,N_4441);
xor UO_794 (O_794,N_4363,N_4540);
nor UO_795 (O_795,N_4807,N_4603);
nor UO_796 (O_796,N_4377,N_4987);
or UO_797 (O_797,N_4259,N_4472);
xnor UO_798 (O_798,N_4991,N_4537);
or UO_799 (O_799,N_4553,N_4338);
nor UO_800 (O_800,N_4944,N_4746);
nor UO_801 (O_801,N_4964,N_4696);
xor UO_802 (O_802,N_4829,N_4718);
xnor UO_803 (O_803,N_4795,N_4119);
xnor UO_804 (O_804,N_4906,N_4643);
and UO_805 (O_805,N_4480,N_4419);
nand UO_806 (O_806,N_4164,N_4939);
nor UO_807 (O_807,N_4147,N_4458);
and UO_808 (O_808,N_4126,N_4274);
and UO_809 (O_809,N_4086,N_4323);
and UO_810 (O_810,N_4488,N_4185);
xnor UO_811 (O_811,N_4755,N_4520);
xnor UO_812 (O_812,N_4669,N_4055);
and UO_813 (O_813,N_4908,N_4602);
nor UO_814 (O_814,N_4344,N_4035);
and UO_815 (O_815,N_4640,N_4139);
nand UO_816 (O_816,N_4364,N_4393);
nor UO_817 (O_817,N_4928,N_4607);
nand UO_818 (O_818,N_4214,N_4375);
nor UO_819 (O_819,N_4318,N_4754);
and UO_820 (O_820,N_4926,N_4098);
xnor UO_821 (O_821,N_4043,N_4708);
or UO_822 (O_822,N_4371,N_4823);
nor UO_823 (O_823,N_4034,N_4434);
and UO_824 (O_824,N_4403,N_4272);
or UO_825 (O_825,N_4610,N_4027);
nor UO_826 (O_826,N_4402,N_4957);
xor UO_827 (O_827,N_4758,N_4378);
nor UO_828 (O_828,N_4918,N_4582);
xnor UO_829 (O_829,N_4080,N_4165);
nor UO_830 (O_830,N_4475,N_4982);
xor UO_831 (O_831,N_4826,N_4650);
nor UO_832 (O_832,N_4479,N_4896);
nand UO_833 (O_833,N_4657,N_4002);
nor UO_834 (O_834,N_4413,N_4829);
nor UO_835 (O_835,N_4608,N_4408);
xnor UO_836 (O_836,N_4720,N_4119);
or UO_837 (O_837,N_4357,N_4708);
xor UO_838 (O_838,N_4600,N_4940);
and UO_839 (O_839,N_4394,N_4118);
and UO_840 (O_840,N_4794,N_4873);
or UO_841 (O_841,N_4813,N_4883);
and UO_842 (O_842,N_4336,N_4793);
or UO_843 (O_843,N_4051,N_4324);
xor UO_844 (O_844,N_4120,N_4818);
nand UO_845 (O_845,N_4312,N_4686);
nand UO_846 (O_846,N_4441,N_4391);
nand UO_847 (O_847,N_4272,N_4004);
and UO_848 (O_848,N_4443,N_4279);
xnor UO_849 (O_849,N_4481,N_4766);
nor UO_850 (O_850,N_4276,N_4379);
nor UO_851 (O_851,N_4325,N_4271);
and UO_852 (O_852,N_4686,N_4364);
nand UO_853 (O_853,N_4925,N_4336);
nor UO_854 (O_854,N_4692,N_4119);
nor UO_855 (O_855,N_4938,N_4176);
and UO_856 (O_856,N_4226,N_4157);
xnor UO_857 (O_857,N_4694,N_4808);
nor UO_858 (O_858,N_4531,N_4662);
xor UO_859 (O_859,N_4645,N_4992);
or UO_860 (O_860,N_4838,N_4111);
xor UO_861 (O_861,N_4122,N_4817);
and UO_862 (O_862,N_4883,N_4617);
or UO_863 (O_863,N_4530,N_4097);
xnor UO_864 (O_864,N_4401,N_4617);
nand UO_865 (O_865,N_4462,N_4541);
nor UO_866 (O_866,N_4863,N_4091);
or UO_867 (O_867,N_4329,N_4598);
nor UO_868 (O_868,N_4269,N_4088);
or UO_869 (O_869,N_4467,N_4885);
and UO_870 (O_870,N_4295,N_4147);
nor UO_871 (O_871,N_4918,N_4246);
nand UO_872 (O_872,N_4687,N_4711);
and UO_873 (O_873,N_4872,N_4350);
and UO_874 (O_874,N_4928,N_4157);
or UO_875 (O_875,N_4892,N_4069);
xor UO_876 (O_876,N_4614,N_4133);
nor UO_877 (O_877,N_4966,N_4032);
nor UO_878 (O_878,N_4670,N_4203);
nand UO_879 (O_879,N_4141,N_4919);
nor UO_880 (O_880,N_4624,N_4041);
nand UO_881 (O_881,N_4192,N_4135);
or UO_882 (O_882,N_4217,N_4539);
or UO_883 (O_883,N_4542,N_4434);
and UO_884 (O_884,N_4255,N_4362);
nor UO_885 (O_885,N_4758,N_4143);
and UO_886 (O_886,N_4069,N_4173);
nand UO_887 (O_887,N_4654,N_4671);
and UO_888 (O_888,N_4694,N_4581);
or UO_889 (O_889,N_4491,N_4828);
nor UO_890 (O_890,N_4283,N_4392);
or UO_891 (O_891,N_4317,N_4474);
nand UO_892 (O_892,N_4168,N_4971);
and UO_893 (O_893,N_4196,N_4486);
xor UO_894 (O_894,N_4682,N_4187);
nand UO_895 (O_895,N_4921,N_4511);
nand UO_896 (O_896,N_4580,N_4256);
xor UO_897 (O_897,N_4168,N_4928);
xor UO_898 (O_898,N_4580,N_4847);
xor UO_899 (O_899,N_4963,N_4981);
nor UO_900 (O_900,N_4937,N_4406);
or UO_901 (O_901,N_4511,N_4927);
nand UO_902 (O_902,N_4745,N_4719);
nor UO_903 (O_903,N_4658,N_4791);
nor UO_904 (O_904,N_4856,N_4773);
nor UO_905 (O_905,N_4515,N_4426);
nand UO_906 (O_906,N_4123,N_4315);
and UO_907 (O_907,N_4593,N_4582);
nor UO_908 (O_908,N_4252,N_4361);
nand UO_909 (O_909,N_4615,N_4875);
nor UO_910 (O_910,N_4673,N_4582);
nor UO_911 (O_911,N_4526,N_4636);
nand UO_912 (O_912,N_4907,N_4198);
nand UO_913 (O_913,N_4769,N_4615);
nor UO_914 (O_914,N_4266,N_4713);
or UO_915 (O_915,N_4623,N_4131);
or UO_916 (O_916,N_4243,N_4262);
nand UO_917 (O_917,N_4351,N_4774);
nand UO_918 (O_918,N_4598,N_4545);
or UO_919 (O_919,N_4376,N_4074);
nand UO_920 (O_920,N_4125,N_4120);
xnor UO_921 (O_921,N_4464,N_4547);
or UO_922 (O_922,N_4948,N_4110);
nor UO_923 (O_923,N_4254,N_4171);
and UO_924 (O_924,N_4673,N_4930);
nand UO_925 (O_925,N_4115,N_4368);
xnor UO_926 (O_926,N_4456,N_4346);
nor UO_927 (O_927,N_4293,N_4099);
or UO_928 (O_928,N_4731,N_4171);
or UO_929 (O_929,N_4282,N_4324);
nor UO_930 (O_930,N_4512,N_4092);
and UO_931 (O_931,N_4105,N_4267);
and UO_932 (O_932,N_4982,N_4774);
and UO_933 (O_933,N_4998,N_4095);
and UO_934 (O_934,N_4681,N_4737);
xnor UO_935 (O_935,N_4920,N_4269);
and UO_936 (O_936,N_4829,N_4167);
nor UO_937 (O_937,N_4175,N_4516);
and UO_938 (O_938,N_4450,N_4809);
or UO_939 (O_939,N_4804,N_4715);
nor UO_940 (O_940,N_4897,N_4601);
or UO_941 (O_941,N_4912,N_4944);
nor UO_942 (O_942,N_4180,N_4574);
nor UO_943 (O_943,N_4762,N_4061);
nand UO_944 (O_944,N_4545,N_4517);
xor UO_945 (O_945,N_4936,N_4668);
nand UO_946 (O_946,N_4336,N_4316);
or UO_947 (O_947,N_4060,N_4540);
xor UO_948 (O_948,N_4045,N_4638);
xnor UO_949 (O_949,N_4301,N_4151);
nor UO_950 (O_950,N_4372,N_4211);
and UO_951 (O_951,N_4039,N_4331);
nor UO_952 (O_952,N_4506,N_4624);
nand UO_953 (O_953,N_4720,N_4293);
or UO_954 (O_954,N_4840,N_4770);
or UO_955 (O_955,N_4417,N_4302);
nor UO_956 (O_956,N_4475,N_4208);
nand UO_957 (O_957,N_4773,N_4907);
or UO_958 (O_958,N_4574,N_4791);
or UO_959 (O_959,N_4911,N_4877);
and UO_960 (O_960,N_4692,N_4586);
or UO_961 (O_961,N_4376,N_4487);
xnor UO_962 (O_962,N_4625,N_4444);
nor UO_963 (O_963,N_4586,N_4718);
or UO_964 (O_964,N_4245,N_4833);
nor UO_965 (O_965,N_4430,N_4371);
and UO_966 (O_966,N_4266,N_4821);
and UO_967 (O_967,N_4184,N_4633);
and UO_968 (O_968,N_4144,N_4673);
or UO_969 (O_969,N_4723,N_4997);
nor UO_970 (O_970,N_4275,N_4369);
nor UO_971 (O_971,N_4477,N_4563);
and UO_972 (O_972,N_4685,N_4622);
nand UO_973 (O_973,N_4943,N_4535);
or UO_974 (O_974,N_4361,N_4198);
nand UO_975 (O_975,N_4264,N_4826);
and UO_976 (O_976,N_4196,N_4245);
and UO_977 (O_977,N_4407,N_4284);
or UO_978 (O_978,N_4214,N_4528);
and UO_979 (O_979,N_4151,N_4455);
nor UO_980 (O_980,N_4696,N_4810);
xnor UO_981 (O_981,N_4327,N_4414);
or UO_982 (O_982,N_4159,N_4636);
nand UO_983 (O_983,N_4059,N_4278);
nor UO_984 (O_984,N_4440,N_4030);
nor UO_985 (O_985,N_4238,N_4033);
xnor UO_986 (O_986,N_4885,N_4757);
nor UO_987 (O_987,N_4159,N_4084);
or UO_988 (O_988,N_4404,N_4166);
or UO_989 (O_989,N_4799,N_4286);
or UO_990 (O_990,N_4316,N_4509);
nand UO_991 (O_991,N_4241,N_4931);
xnor UO_992 (O_992,N_4859,N_4225);
nor UO_993 (O_993,N_4328,N_4027);
nand UO_994 (O_994,N_4160,N_4654);
nand UO_995 (O_995,N_4096,N_4259);
nor UO_996 (O_996,N_4911,N_4919);
and UO_997 (O_997,N_4554,N_4090);
or UO_998 (O_998,N_4399,N_4083);
or UO_999 (O_999,N_4582,N_4311);
endmodule