module basic_3000_30000_3500_10_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_1065,In_1258);
nand U1 (N_1,In_303,In_1598);
xor U2 (N_2,In_124,In_1834);
or U3 (N_3,In_2250,In_2534);
nand U4 (N_4,In_2057,In_2527);
nor U5 (N_5,In_1767,In_1497);
nand U6 (N_6,In_2221,In_1285);
nand U7 (N_7,In_2547,In_2574);
nor U8 (N_8,In_2260,In_2202);
and U9 (N_9,In_982,In_943);
or U10 (N_10,In_2207,In_1018);
or U11 (N_11,In_2892,In_2881);
nor U12 (N_12,In_222,In_740);
and U13 (N_13,In_1079,In_2418);
or U14 (N_14,In_438,In_692);
and U15 (N_15,In_728,In_2432);
nor U16 (N_16,In_2307,In_1352);
xnor U17 (N_17,In_1701,In_1003);
xor U18 (N_18,In_2135,In_1212);
and U19 (N_19,In_2867,In_1215);
nand U20 (N_20,In_1973,In_1957);
or U21 (N_21,In_1382,In_1988);
and U22 (N_22,In_2518,In_1318);
and U23 (N_23,In_635,In_2817);
nor U24 (N_24,In_1297,In_1322);
nor U25 (N_25,In_915,In_2709);
nor U26 (N_26,In_1929,In_2297);
and U27 (N_27,In_622,In_1177);
nand U28 (N_28,In_2106,In_150);
or U29 (N_29,In_318,In_2830);
nor U30 (N_30,In_923,In_989);
and U31 (N_31,In_2062,In_731);
nand U32 (N_32,In_2801,In_236);
nor U33 (N_33,In_440,In_2998);
xor U34 (N_34,In_2684,In_146);
xnor U35 (N_35,In_426,In_257);
xnor U36 (N_36,In_1566,In_1151);
xnor U37 (N_37,In_1800,In_1797);
nand U38 (N_38,In_2490,In_925);
nor U39 (N_39,In_1176,In_118);
and U40 (N_40,In_2988,In_2002);
xnor U41 (N_41,In_909,In_1931);
xor U42 (N_42,In_2852,In_745);
and U43 (N_43,In_194,In_2918);
nand U44 (N_44,In_1491,In_1062);
xnor U45 (N_45,In_2103,In_1189);
nand U46 (N_46,In_2741,In_2276);
or U47 (N_47,In_1265,In_1156);
and U48 (N_48,In_1299,In_2083);
nand U49 (N_49,In_722,In_1480);
xor U50 (N_50,In_1599,In_956);
or U51 (N_51,In_2258,In_1493);
nand U52 (N_52,In_511,In_2790);
and U53 (N_53,In_2400,In_1969);
nor U54 (N_54,In_2020,In_1096);
xor U55 (N_55,In_2049,In_1788);
xnor U56 (N_56,In_1585,In_1120);
or U57 (N_57,In_1292,In_206);
or U58 (N_58,In_1467,In_788);
and U59 (N_59,In_2621,In_1708);
nor U60 (N_60,In_1905,In_2027);
or U61 (N_61,In_872,In_1015);
xor U62 (N_62,In_1434,In_1635);
nand U63 (N_63,In_2774,In_623);
nand U64 (N_64,In_2039,In_980);
nand U65 (N_65,In_2491,In_499);
nor U66 (N_66,In_1354,In_3);
and U67 (N_67,In_1745,In_2249);
or U68 (N_68,In_397,In_315);
xor U69 (N_69,In_239,In_476);
or U70 (N_70,In_2128,In_1192);
nor U71 (N_71,In_2509,In_83);
xnor U72 (N_72,In_940,In_2657);
and U73 (N_73,In_1774,In_2174);
xnor U74 (N_74,In_409,In_2540);
xor U75 (N_75,In_1684,In_541);
or U76 (N_76,In_81,In_2559);
and U77 (N_77,In_2392,In_2612);
nand U78 (N_78,In_2653,In_132);
and U79 (N_79,In_1455,In_2126);
and U80 (N_80,In_1183,In_733);
nand U81 (N_81,In_952,In_2452);
and U82 (N_82,In_805,In_1019);
nor U83 (N_83,In_212,In_108);
xnor U84 (N_84,In_2633,In_2665);
nand U85 (N_85,In_1617,In_404);
and U86 (N_86,In_1794,In_475);
and U87 (N_87,In_162,In_1966);
and U88 (N_88,In_2847,In_1216);
xor U89 (N_89,In_2829,In_636);
xor U90 (N_90,In_505,In_981);
and U91 (N_91,In_596,In_2733);
nand U92 (N_92,In_447,In_2778);
nor U93 (N_93,In_710,In_1396);
nor U94 (N_94,In_1013,In_695);
and U95 (N_95,In_2632,In_2893);
xor U96 (N_96,In_2934,In_2552);
or U97 (N_97,In_977,In_2691);
nand U98 (N_98,In_1228,In_429);
and U99 (N_99,In_1512,In_2754);
and U100 (N_100,In_2254,In_2320);
nand U101 (N_101,In_2065,In_608);
xnor U102 (N_102,In_539,In_2155);
and U103 (N_103,In_2642,In_1364);
xor U104 (N_104,In_361,In_2375);
and U105 (N_105,In_1024,In_815);
xor U106 (N_106,In_804,In_899);
nand U107 (N_107,In_2596,In_2915);
nor U108 (N_108,In_2047,In_610);
nand U109 (N_109,In_347,In_1443);
nand U110 (N_110,In_2343,In_2603);
xor U111 (N_111,In_929,In_2854);
or U112 (N_112,In_882,In_504);
xor U113 (N_113,In_2616,In_219);
nand U114 (N_114,In_282,In_2129);
nor U115 (N_115,In_1017,In_1411);
xor U116 (N_116,In_2462,In_2654);
nand U117 (N_117,In_2206,In_1476);
xor U118 (N_118,In_170,In_2025);
nor U119 (N_119,In_91,In_1914);
or U120 (N_120,In_2506,In_1539);
and U121 (N_121,In_1325,In_297);
nand U122 (N_122,In_799,In_864);
nor U123 (N_123,In_2765,In_1716);
xor U124 (N_124,In_163,In_2874);
xor U125 (N_125,In_1501,In_1742);
and U126 (N_126,In_164,In_574);
and U127 (N_127,In_421,In_2210);
nor U128 (N_128,In_2600,In_1779);
xor U129 (N_129,In_384,In_1038);
or U130 (N_130,In_1317,In_2233);
and U131 (N_131,In_2676,In_2976);
nand U132 (N_132,In_1239,In_594);
nor U133 (N_133,In_2118,In_1372);
nand U134 (N_134,In_1217,In_2700);
nor U135 (N_135,In_552,In_79);
nand U136 (N_136,In_1913,In_1181);
or U137 (N_137,In_2377,In_1843);
and U138 (N_138,In_1655,In_904);
and U139 (N_139,In_1141,In_2245);
and U140 (N_140,In_1266,In_1826);
nor U141 (N_141,In_2869,In_2929);
and U142 (N_142,In_46,In_2115);
xor U143 (N_143,In_1390,In_2521);
xor U144 (N_144,In_152,In_1238);
and U145 (N_145,In_143,In_427);
or U146 (N_146,In_2463,In_202);
nor U147 (N_147,In_2932,In_410);
and U148 (N_148,In_2764,In_2394);
nor U149 (N_149,In_372,In_2017);
nor U150 (N_150,In_756,In_2641);
xor U151 (N_151,In_1223,In_1681);
and U152 (N_152,In_2219,In_1268);
or U153 (N_153,In_1053,In_1306);
nand U154 (N_154,In_1996,In_1486);
xor U155 (N_155,In_311,In_588);
and U156 (N_156,In_828,In_822);
nand U157 (N_157,In_924,In_198);
nand U158 (N_158,In_618,In_839);
nor U159 (N_159,In_530,In_825);
nand U160 (N_160,In_2190,In_2409);
xnor U161 (N_161,In_184,In_750);
nor U162 (N_162,In_1994,In_2987);
nor U163 (N_163,In_1336,In_605);
or U164 (N_164,In_2040,In_1169);
xnor U165 (N_165,In_1144,In_1232);
nand U166 (N_166,In_2051,In_918);
nor U167 (N_167,In_1457,In_320);
nor U168 (N_168,In_2385,In_1555);
nor U169 (N_169,In_387,In_378);
or U170 (N_170,In_2136,In_1004);
nand U171 (N_171,In_2413,In_415);
and U172 (N_172,In_1546,In_2211);
xor U173 (N_173,In_935,In_2763);
or U174 (N_174,In_2557,In_2434);
nor U175 (N_175,In_734,In_1508);
xor U176 (N_176,In_1876,In_1646);
xor U177 (N_177,In_1472,In_246);
nor U178 (N_178,In_2648,In_992);
nand U179 (N_179,In_893,In_2422);
xor U180 (N_180,In_1631,In_2526);
xor U181 (N_181,In_2080,In_2026);
and U182 (N_182,In_1234,In_1267);
xor U183 (N_183,In_1262,In_418);
nand U184 (N_184,In_11,In_2531);
nor U185 (N_185,In_2538,In_1888);
nand U186 (N_186,In_2322,In_966);
or U187 (N_187,In_2873,In_1245);
and U188 (N_188,In_1959,In_1670);
nor U189 (N_189,In_2991,In_531);
or U190 (N_190,In_506,In_1880);
nand U191 (N_191,In_241,In_1580);
nand U192 (N_192,In_1178,In_2139);
nand U193 (N_193,In_189,In_324);
xnor U194 (N_194,In_2837,In_265);
nand U195 (N_195,In_856,In_1344);
or U196 (N_196,In_806,In_881);
nor U197 (N_197,In_2092,In_1901);
nand U198 (N_198,In_1606,In_1121);
nand U199 (N_199,In_2662,In_99);
nand U200 (N_200,In_2104,In_730);
and U201 (N_201,In_349,In_2528);
nor U202 (N_202,In_483,In_1224);
and U203 (N_203,In_52,In_2146);
and U204 (N_204,In_1662,In_2124);
nand U205 (N_205,In_225,In_609);
or U206 (N_206,In_2220,In_1253);
and U207 (N_207,In_1822,In_2154);
or U208 (N_208,In_2485,In_326);
and U209 (N_209,In_2795,In_2113);
nor U210 (N_210,In_457,In_1068);
xnor U211 (N_211,In_1470,In_2328);
nor U212 (N_212,In_721,In_270);
nand U213 (N_213,In_14,In_2339);
nand U214 (N_214,In_912,In_777);
and U215 (N_215,In_773,In_28);
nor U216 (N_216,In_2548,In_816);
and U217 (N_217,In_876,In_66);
and U218 (N_218,In_2515,In_253);
nand U219 (N_219,In_634,In_2205);
xnor U220 (N_220,In_2985,In_2169);
nand U221 (N_221,In_2454,In_2724);
nand U222 (N_222,In_897,In_602);
nor U223 (N_223,In_50,In_2259);
xor U224 (N_224,In_611,In_1586);
xor U225 (N_225,In_1851,In_2832);
nand U226 (N_226,In_857,In_1984);
xor U227 (N_227,In_2969,In_808);
and U228 (N_228,In_2925,In_727);
or U229 (N_229,In_1620,In_1621);
and U230 (N_230,In_1423,In_1401);
and U231 (N_231,In_1678,In_2660);
and U232 (N_232,In_479,In_1874);
nand U233 (N_233,In_1628,In_1793);
nor U234 (N_234,In_1375,In_2467);
xor U235 (N_235,In_153,In_1837);
nand U236 (N_236,In_354,In_1029);
or U237 (N_237,In_2979,In_294);
xor U238 (N_238,In_1408,In_2672);
nand U239 (N_239,In_1052,In_2348);
nand U240 (N_240,In_2806,In_1664);
xnor U241 (N_241,In_2488,In_1772);
and U242 (N_242,In_2808,In_2279);
nor U243 (N_243,In_1526,In_2038);
nand U244 (N_244,In_420,In_1857);
nor U245 (N_245,In_1836,In_2738);
and U246 (N_246,In_2313,In_895);
nand U247 (N_247,In_1552,In_889);
or U248 (N_248,In_2086,In_358);
nor U249 (N_249,In_2519,In_954);
and U250 (N_250,In_1712,In_2530);
and U251 (N_251,In_879,In_380);
nand U252 (N_252,In_2912,In_2833);
nor U253 (N_253,In_1485,In_550);
xnor U254 (N_254,In_2785,In_2889);
and U255 (N_255,In_2666,In_412);
nor U256 (N_256,In_2029,In_1484);
and U257 (N_257,In_2698,In_2678);
and U258 (N_258,In_1468,In_1391);
nand U259 (N_259,In_1722,In_1859);
xor U260 (N_260,In_2284,In_2142);
or U261 (N_261,In_1203,In_215);
xnor U262 (N_262,In_1867,In_1140);
nor U263 (N_263,In_428,In_686);
xnor U264 (N_264,In_1264,In_1393);
xor U265 (N_265,In_1944,In_1179);
and U266 (N_266,In_843,In_1608);
and U267 (N_267,In_2402,In_2081);
or U268 (N_268,In_310,In_2586);
and U269 (N_269,In_1247,In_2296);
nor U270 (N_270,In_2865,In_2478);
nor U271 (N_271,In_2070,In_1110);
nand U272 (N_272,In_1761,In_2508);
xnor U273 (N_273,In_156,In_2165);
xnor U274 (N_274,In_1051,In_997);
xnor U275 (N_275,In_698,In_2560);
xnor U276 (N_276,In_1440,In_1927);
or U277 (N_277,In_2597,In_2366);
nor U278 (N_278,In_2371,In_2228);
and U279 (N_279,In_17,In_110);
or U280 (N_280,In_1269,In_1616);
nor U281 (N_281,In_709,In_2683);
nand U282 (N_282,In_580,In_2697);
xor U283 (N_283,In_942,In_2333);
nand U284 (N_284,In_1031,In_2201);
nor U285 (N_285,In_293,In_54);
or U286 (N_286,In_639,In_154);
xnor U287 (N_287,In_1803,In_724);
nand U288 (N_288,In_300,In_308);
xor U289 (N_289,In_1645,In_2293);
nand U290 (N_290,In_1782,In_1474);
xor U291 (N_291,In_2318,In_1168);
and U292 (N_292,In_1809,In_795);
or U293 (N_293,In_2706,In_810);
xnor U294 (N_294,In_1385,In_1962);
nand U295 (N_295,In_339,In_1473);
xor U296 (N_296,In_2567,In_762);
nor U297 (N_297,In_1271,In_2855);
nor U298 (N_298,In_1928,In_2747);
nand U299 (N_299,In_175,In_1078);
nor U300 (N_300,In_841,In_1821);
nand U301 (N_301,In_2156,In_624);
or U302 (N_302,In_1074,In_829);
and U303 (N_303,In_811,In_1918);
and U304 (N_304,In_48,In_1101);
and U305 (N_305,In_467,In_2068);
nor U306 (N_306,In_2649,In_1106);
or U307 (N_307,In_934,In_669);
xnor U308 (N_308,In_2093,In_325);
and U309 (N_309,In_963,In_675);
nor U310 (N_310,In_544,In_1230);
xnor U311 (N_311,In_430,In_482);
or U312 (N_312,In_478,In_1376);
xnor U313 (N_313,In_2175,In_2448);
nor U314 (N_314,In_2390,In_1981);
or U315 (N_315,In_459,In_1193);
and U316 (N_316,In_2,In_2084);
nor U317 (N_317,In_97,In_2480);
nor U318 (N_318,In_1668,In_2010);
xor U319 (N_319,In_2794,In_1482);
and U320 (N_320,In_565,In_1725);
nand U321 (N_321,In_2652,In_2003);
and U322 (N_322,In_706,In_1991);
and U323 (N_323,In_1533,In_1743);
nor U324 (N_324,In_654,In_2168);
nor U325 (N_325,In_1827,In_456);
nand U326 (N_326,In_149,In_2464);
or U327 (N_327,In_2252,In_115);
xnor U328 (N_328,In_1477,In_76);
nand U329 (N_329,In_350,In_2071);
and U330 (N_330,In_2606,In_321);
xnor U331 (N_331,In_619,In_1281);
or U332 (N_332,In_2525,In_2466);
nor U333 (N_333,In_1817,In_411);
and U334 (N_334,In_986,In_1511);
or U335 (N_335,In_535,In_359);
or U336 (N_336,In_355,In_1567);
nand U337 (N_337,In_922,In_148);
xnor U338 (N_338,In_174,In_2564);
nor U339 (N_339,In_2565,In_95);
and U340 (N_340,In_1414,In_489);
and U341 (N_341,In_2674,In_2317);
nand U342 (N_342,In_1498,In_262);
or U343 (N_343,In_2631,In_363);
xor U344 (N_344,In_51,In_130);
or U345 (N_345,In_250,In_2048);
nor U346 (N_346,In_2311,In_582);
and U347 (N_347,In_1211,In_1956);
and U348 (N_348,In_1590,In_1202);
xor U349 (N_349,In_106,In_168);
xor U350 (N_350,In_662,In_1321);
and U351 (N_351,In_2599,In_1201);
or U352 (N_352,In_2791,In_1448);
xnor U353 (N_353,In_2090,In_2831);
and U354 (N_354,In_1802,In_2489);
and U355 (N_355,In_560,In_2849);
and U356 (N_356,In_754,In_1075);
or U357 (N_357,In_1064,In_13);
and U358 (N_358,In_1296,In_525);
nand U359 (N_359,In_524,In_465);
nand U360 (N_360,In_94,In_2421);
xor U361 (N_361,In_2766,In_1399);
or U362 (N_362,In_158,In_1431);
or U363 (N_363,In_1190,In_1444);
and U364 (N_364,In_2581,In_371);
nor U365 (N_365,In_2486,In_1707);
nor U366 (N_366,In_2590,In_2520);
and U367 (N_367,In_823,In_254);
and U368 (N_368,In_119,In_2938);
nand U369 (N_369,In_1738,In_453);
or U370 (N_370,In_2809,In_1618);
nand U371 (N_371,In_2571,In_758);
nor U372 (N_372,In_2983,In_68);
nor U373 (N_373,In_2445,In_1593);
xor U374 (N_374,In_668,In_2189);
nor U375 (N_375,In_2037,In_1895);
and U376 (N_376,In_911,In_1600);
and U377 (N_377,In_1965,In_1244);
xnor U378 (N_378,In_323,In_538);
nor U379 (N_379,In_1,In_587);
and U380 (N_380,In_1324,In_906);
xor U381 (N_381,In_77,In_2378);
and U382 (N_382,In_2812,In_655);
nor U383 (N_383,In_1311,In_2088);
and U384 (N_384,In_1881,In_2417);
xor U385 (N_385,In_2423,In_2303);
nand U386 (N_386,In_1977,In_1624);
nand U387 (N_387,In_1879,In_2588);
or U388 (N_388,In_187,In_1556);
or U389 (N_389,In_2426,In_2050);
or U390 (N_390,In_2412,In_492);
nand U391 (N_391,In_1020,In_542);
or U392 (N_392,In_1161,In_2277);
nor U393 (N_393,In_2441,In_1577);
xor U394 (N_394,In_931,In_1206);
or U395 (N_395,In_836,In_945);
nand U396 (N_396,In_1419,In_1221);
and U397 (N_397,In_2000,In_1919);
or U398 (N_398,In_480,In_1661);
and U399 (N_399,In_2793,In_2714);
nand U400 (N_400,In_1775,In_2141);
nand U401 (N_401,In_1058,In_1528);
nand U402 (N_402,In_1846,In_2671);
xnor U403 (N_403,In_78,In_786);
nand U404 (N_404,In_201,In_2550);
nand U405 (N_405,In_2900,In_2109);
nor U406 (N_406,In_995,In_1786);
and U407 (N_407,In_2059,In_2238);
and U408 (N_408,In_632,In_2194);
or U409 (N_409,In_2294,In_1912);
and U410 (N_410,In_2213,In_1500);
or U411 (N_411,In_2924,In_2171);
nand U412 (N_412,In_1502,In_548);
or U413 (N_413,In_264,In_2326);
nand U414 (N_414,In_833,In_1773);
nand U415 (N_415,In_1524,In_140);
and U416 (N_416,In_1307,In_1014);
nor U417 (N_417,In_1792,In_135);
or U418 (N_418,In_2404,In_2816);
nor U419 (N_419,In_1514,In_2431);
or U420 (N_420,In_1993,In_2046);
nand U421 (N_421,In_183,In_63);
and U422 (N_422,In_769,In_2569);
nand U423 (N_423,In_1925,In_1790);
or U424 (N_424,In_2759,In_1093);
nor U425 (N_425,In_1142,In_543);
nor U426 (N_426,In_689,In_919);
and U427 (N_427,In_2879,In_1255);
or U428 (N_428,In_1111,In_2060);
and U429 (N_429,In_1808,In_2860);
nor U430 (N_430,In_1873,In_2330);
or U431 (N_431,In_528,In_968);
xnor U432 (N_432,In_2089,In_1717);
xor U433 (N_433,In_330,In_557);
nor U434 (N_434,In_2393,In_1025);
nand U435 (N_435,In_327,In_1237);
xor U436 (N_436,In_8,In_288);
xor U437 (N_437,In_1407,In_933);
or U438 (N_438,In_2353,In_2681);
nor U439 (N_439,In_2907,In_2278);
or U440 (N_440,In_988,In_1081);
or U441 (N_441,In_1172,In_2300);
nor U442 (N_442,In_1804,In_653);
or U443 (N_443,In_1103,In_369);
xnor U444 (N_444,In_2713,In_1222);
and U445 (N_445,In_2044,In_920);
nand U446 (N_446,In_2111,In_2425);
nand U447 (N_447,In_2166,In_2601);
or U448 (N_448,In_1679,In_80);
xor U449 (N_449,In_1291,In_491);
nor U450 (N_450,In_1739,In_693);
nor U451 (N_451,In_2123,In_2471);
nor U452 (N_452,In_1591,In_2614);
and U453 (N_453,In_290,In_1341);
nor U454 (N_454,In_285,In_739);
xnor U455 (N_455,In_1955,In_337);
nor U456 (N_456,In_416,In_2777);
and U457 (N_457,In_2043,In_1254);
nand U458 (N_458,In_658,In_367);
nand U459 (N_459,In_737,In_680);
or U460 (N_460,In_2744,In_335);
or U461 (N_461,In_1884,In_1711);
xor U462 (N_462,In_2209,In_913);
and U463 (N_463,In_213,In_555);
or U464 (N_464,In_1397,In_1510);
xor U465 (N_465,In_809,In_2750);
nor U466 (N_466,In_2449,In_29);
nor U467 (N_467,In_2056,In_136);
and U468 (N_468,In_2585,In_2164);
and U469 (N_469,In_651,In_2041);
and U470 (N_470,In_2256,In_2511);
and U471 (N_471,In_1687,In_1350);
and U472 (N_472,In_1116,In_2708);
xnor U473 (N_473,In_278,In_2913);
or U474 (N_474,In_1858,In_2183);
nor U475 (N_475,In_551,In_533);
and U476 (N_476,In_2381,In_1882);
nor U477 (N_477,In_1752,In_233);
nor U478 (N_478,In_850,In_987);
or U479 (N_479,In_2298,In_2236);
and U480 (N_480,In_1349,In_2610);
xnor U481 (N_481,In_2703,In_2916);
xor U482 (N_482,In_855,In_2069);
or U483 (N_483,In_1820,In_334);
xnor U484 (N_484,In_2216,In_1578);
xor U485 (N_485,In_672,In_584);
nor U486 (N_486,In_1762,In_699);
and U487 (N_487,In_396,In_1138);
and U488 (N_488,In_2470,In_1850);
or U489 (N_489,In_1398,In_7);
nand U490 (N_490,In_2736,In_2973);
nor U491 (N_491,In_785,In_33);
or U492 (N_492,In_144,In_1034);
and U493 (N_493,In_819,In_1449);
nor U494 (N_494,In_1421,In_697);
nand U495 (N_495,In_374,In_2710);
or U496 (N_496,In_1780,In_1011);
xor U497 (N_497,In_1134,In_2577);
and U498 (N_498,In_1844,In_592);
nand U499 (N_499,In_1367,In_1806);
and U500 (N_500,In_2570,In_2208);
xnor U501 (N_501,In_2920,In_2563);
xnor U502 (N_502,In_1191,In_1728);
nand U503 (N_503,In_1359,In_892);
or U504 (N_504,In_306,In_783);
xnor U505 (N_505,In_2994,In_1758);
and U506 (N_506,In_1220,In_1921);
nand U507 (N_507,In_2292,In_2715);
nand U508 (N_508,In_1922,In_442);
or U509 (N_509,In_2628,In_2487);
and U510 (N_510,In_534,In_26);
or U511 (N_511,In_2620,In_2325);
nand U512 (N_512,In_263,In_790);
nor U513 (N_513,In_1086,In_600);
nor U514 (N_514,In_2203,In_238);
or U515 (N_515,In_96,In_1887);
xor U516 (N_516,In_1562,In_826);
xnor U517 (N_517,In_1633,In_1750);
xor U518 (N_518,In_1136,In_793);
or U519 (N_519,In_1710,In_2953);
nor U520 (N_520,In_1769,In_1233);
or U521 (N_521,In_688,In_2196);
or U522 (N_522,In_513,In_678);
xor U523 (N_523,In_272,In_1579);
nand U524 (N_524,In_2321,In_142);
nor U525 (N_525,In_615,In_2134);
nor U526 (N_526,In_1316,In_366);
nor U527 (N_527,In_2416,In_1404);
xnor U528 (N_528,In_1824,In_2504);
nand U529 (N_529,In_1564,In_392);
and U530 (N_530,In_1418,In_936);
xor U531 (N_531,In_2618,In_1863);
or U532 (N_532,In_853,In_2419);
xor U533 (N_533,In_2182,In_1274);
or U534 (N_534,In_2549,In_2611);
and U535 (N_535,In_1466,In_2382);
and U536 (N_536,In_2078,In_2992);
nor U537 (N_537,In_502,In_439);
or U538 (N_538,In_1329,In_1847);
nor U539 (N_539,In_2021,In_1160);
and U540 (N_540,In_1632,In_1864);
xor U541 (N_541,In_2836,In_817);
nor U542 (N_542,In_2323,In_2359);
nand U543 (N_543,In_1719,In_569);
nand U544 (N_544,In_2268,In_23);
xnor U545 (N_545,In_501,In_2158);
nor U546 (N_546,In_1518,In_962);
xor U547 (N_547,In_1595,In_2484);
and U548 (N_548,In_2099,In_1164);
or U549 (N_549,In_2064,In_2450);
or U550 (N_550,In_2898,In_620);
and U551 (N_551,In_322,In_908);
and U552 (N_552,In_838,In_357);
or U553 (N_553,In_2316,In_1060);
or U554 (N_554,In_648,In_226);
xnor U555 (N_555,In_1968,In_1734);
nor U556 (N_556,In_1532,In_2908);
nand U557 (N_557,In_1417,In_946);
nor U558 (N_558,In_998,In_1866);
or U559 (N_559,In_760,In_2602);
or U560 (N_560,In_1009,In_2122);
nand U561 (N_561,In_2232,In_362);
nand U562 (N_562,In_1277,In_88);
or U563 (N_563,In_1900,In_953);
or U564 (N_564,In_1787,In_2595);
or U565 (N_565,In_990,In_666);
nor U566 (N_566,In_1601,In_1105);
and U567 (N_567,In_2167,In_333);
xor U568 (N_568,In_1205,In_652);
nand U569 (N_569,In_1462,In_2712);
nand U570 (N_570,In_407,In_317);
nor U571 (N_571,In_2161,In_526);
and U572 (N_572,In_631,In_1509);
nor U573 (N_573,In_1522,In_2192);
xor U574 (N_574,In_2825,In_529);
xnor U575 (N_575,In_180,In_56);
nand U576 (N_576,In_736,In_218);
and U577 (N_577,In_1200,In_782);
nand U578 (N_578,In_1494,In_1607);
or U579 (N_579,In_970,In_247);
nand U580 (N_580,In_1924,In_304);
nor U581 (N_581,In_865,In_1043);
and U582 (N_582,In_2857,In_2076);
xor U583 (N_583,In_1173,In_967);
nor U584 (N_584,In_167,In_2362);
nor U585 (N_585,In_495,In_1461);
and U586 (N_586,In_2755,In_959);
and U587 (N_587,In_1938,In_67);
and U588 (N_588,In_1990,In_877);
nand U589 (N_589,In_2481,In_1446);
nor U590 (N_590,In_1805,In_852);
xor U591 (N_591,In_390,In_196);
or U592 (N_592,In_313,In_606);
xnor U593 (N_593,In_1940,In_207);
and U594 (N_594,In_789,In_685);
nand U595 (N_595,In_1478,In_1471);
xnor U596 (N_596,In_472,In_72);
or U597 (N_597,In_832,In_868);
or U598 (N_598,In_1764,In_2877);
or U599 (N_599,In_991,In_1706);
and U600 (N_600,In_794,In_1293);
or U601 (N_601,In_599,In_2922);
nor U602 (N_602,In_2177,In_2798);
xor U603 (N_603,In_2927,In_2771);
or U604 (N_604,In_1463,In_1823);
xnor U605 (N_605,In_2958,In_1044);
nand U606 (N_606,In_1961,In_419);
and U607 (N_607,In_1543,In_1958);
nand U608 (N_608,In_650,In_1073);
nor U609 (N_609,In_477,In_2435);
and U610 (N_610,In_2499,In_468);
or U611 (N_611,In_711,In_1852);
xor U612 (N_612,In_20,In_831);
nand U613 (N_613,In_1312,In_1123);
nor U614 (N_614,In_2589,In_2661);
or U615 (N_615,In_1436,In_2286);
xor U616 (N_616,In_2533,In_296);
or U617 (N_617,In_2054,In_1226);
and U618 (N_618,In_649,In_2797);
nor U619 (N_619,In_295,In_422);
or U620 (N_620,In_2289,In_2336);
nand U621 (N_621,In_604,In_2690);
nand U622 (N_622,In_1865,In_1174);
and U623 (N_623,In_2880,In_2227);
or U624 (N_624,In_176,In_1795);
xor U625 (N_625,In_572,In_2592);
nor U626 (N_626,In_2888,In_2758);
nand U627 (N_627,In_352,In_111);
xor U628 (N_628,In_1856,In_1897);
nand U629 (N_629,In_19,In_2420);
and U630 (N_630,In_2143,In_948);
nand U631 (N_631,In_1736,In_1377);
nand U632 (N_632,In_1974,In_1481);
xor U633 (N_633,In_2670,In_2947);
and U634 (N_634,In_2989,In_960);
nor U635 (N_635,In_1149,In_1548);
nand U636 (N_636,In_1571,In_2761);
or U637 (N_637,In_2305,In_1666);
xor U638 (N_638,In_2077,In_1871);
or U639 (N_639,In_1235,In_2162);
or U640 (N_640,In_503,In_1680);
xnor U641 (N_641,In_2770,In_1315);
xor U642 (N_642,In_702,In_1295);
or U643 (N_643,In_1057,In_1853);
nand U644 (N_644,In_2680,In_732);
or U645 (N_645,In_2767,In_1090);
nor U646 (N_646,In_1339,In_1849);
nand U647 (N_647,In_1980,In_1989);
nor U648 (N_648,In_2748,In_1935);
and U649 (N_649,In_21,In_1531);
or U650 (N_650,In_2875,In_570);
xnor U651 (N_651,In_2545,In_2848);
nor U652 (N_652,In_1159,In_1771);
nor U653 (N_653,In_2095,In_1107);
xor U654 (N_654,In_1405,In_1675);
nor U655 (N_655,In_863,In_2910);
nor U656 (N_656,In_2802,In_2803);
and U657 (N_657,In_1252,In_1198);
xnor U658 (N_658,In_2186,In_230);
nor U659 (N_659,In_2501,In_1162);
or U660 (N_660,In_1288,In_166);
and U661 (N_661,In_340,In_114);
nand U662 (N_662,In_220,In_244);
xnor U663 (N_663,In_1721,In_1796);
nor U664 (N_664,In_329,In_1970);
xnor U665 (N_665,In_866,In_116);
and U666 (N_666,In_1126,In_2087);
or U667 (N_667,In_1129,In_49);
nand U668 (N_668,In_2082,In_1042);
nand U669 (N_669,In_2970,In_667);
or U670 (N_670,In_1442,In_2447);
nor U671 (N_671,In_1576,In_771);
nand U672 (N_672,In_1054,In_1939);
nand U673 (N_673,In_1976,In_1100);
and U674 (N_674,In_353,In_1569);
nand U675 (N_675,In_2152,In_1056);
xnor U676 (N_676,In_1006,In_1634);
nand U677 (N_677,In_2822,In_1902);
xor U678 (N_678,In_2891,In_1972);
nor U679 (N_679,In_2160,In_537);
nand U680 (N_680,In_645,In_1830);
nor U681 (N_681,In_802,In_1095);
or U682 (N_682,In_1860,In_319);
or U683 (N_683,In_848,In_209);
or U684 (N_684,In_926,In_586);
or U685 (N_685,In_1702,In_2255);
xor U686 (N_686,In_1848,In_1669);
xor U687 (N_687,In_1798,In_1819);
or U688 (N_688,In_2862,In_1032);
or U689 (N_689,In_1813,In_2309);
and U690 (N_690,In_2742,In_509);
and U691 (N_691,In_1059,In_2212);
nor U692 (N_692,In_2372,In_1839);
or U693 (N_693,In_9,In_1582);
or U694 (N_694,In_1303,In_1158);
and U695 (N_695,In_1642,In_1656);
nor U696 (N_696,In_849,In_2475);
or U697 (N_697,In_1219,In_93);
nand U698 (N_698,In_2625,In_894);
nor U699 (N_699,In_275,In_2923);
and U700 (N_700,In_338,In_979);
nor U701 (N_701,In_2477,In_2796);
xnor U702 (N_702,In_385,In_55);
nand U703 (N_703,In_1611,In_2959);
xor U704 (N_704,In_2248,In_707);
nor U705 (N_705,In_1196,In_1425);
nand U706 (N_706,In_2948,In_417);
and U707 (N_707,In_1186,In_2360);
and U708 (N_708,In_1026,In_446);
xor U709 (N_709,In_2728,In_1394);
nand U710 (N_710,In_2695,In_549);
nand U711 (N_711,In_603,In_1535);
nor U712 (N_712,In_2919,In_84);
xor U713 (N_713,In_1868,In_2542);
and U714 (N_714,In_2694,In_2304);
or U715 (N_715,In_445,In_1542);
or U716 (N_716,In_719,In_1197);
nand U717 (N_717,In_2473,In_1084);
nand U718 (N_718,In_1596,In_1333);
nor U719 (N_719,In_1454,In_2647);
and U720 (N_720,In_1686,In_1132);
nor U721 (N_721,In_1609,In_1378);
nor U722 (N_722,In_563,In_835);
and U723 (N_723,In_2935,In_1908);
or U724 (N_724,In_2532,In_1521);
nor U725 (N_725,In_2365,In_1182);
or U726 (N_726,In_1135,In_614);
or U727 (N_727,In_2474,In_2566);
or U728 (N_728,In_1886,In_1125);
nand U729 (N_729,In_1683,In_2737);
xnor U730 (N_730,In_1952,In_554);
or U731 (N_731,In_748,In_883);
and U732 (N_732,In_1108,In_2349);
and U733 (N_733,In_1650,In_1870);
or U734 (N_734,In_999,In_186);
and U735 (N_735,In_2894,In_558);
nor U736 (N_736,In_527,In_1010);
nor U737 (N_737,In_723,In_2823);
or U738 (N_738,In_399,In_2960);
nand U739 (N_739,In_2997,In_2483);
xor U740 (N_740,In_481,In_1433);
nand U741 (N_741,In_128,In_2458);
xor U742 (N_742,In_712,In_2096);
or U743 (N_743,In_2114,In_1713);
or U744 (N_744,In_1995,In_1022);
nand U745 (N_745,In_1838,In_867);
nor U746 (N_746,In_1428,In_1112);
xnor U747 (N_747,In_121,In_2615);
and U748 (N_748,In_2977,In_2962);
or U749 (N_749,In_1515,In_2931);
or U750 (N_750,In_2288,In_641);
nor U751 (N_751,In_2792,In_2373);
nor U752 (N_752,In_1381,In_356);
or U753 (N_753,In_647,In_102);
xnor U754 (N_754,In_444,In_2398);
xnor U755 (N_755,In_2553,In_776);
nor U756 (N_756,In_2121,In_1049);
and U757 (N_757,In_1409,In_1978);
nand U758 (N_758,In_488,In_2344);
nor U759 (N_759,In_2826,In_2905);
and U760 (N_760,In_101,In_484);
or U761 (N_761,In_2885,In_1979);
xnor U762 (N_762,In_2800,In_573);
nor U763 (N_763,In_2153,In_65);
nor U764 (N_764,In_778,In_1050);
nand U765 (N_765,In_1236,In_2200);
xor U766 (N_766,In_1208,In_2178);
xnor U767 (N_767,In_2950,In_2045);
nand U768 (N_768,In_1282,In_2329);
and U769 (N_769,In_2376,In_2579);
nor U770 (N_770,In_1122,In_1915);
xor U771 (N_771,In_449,In_2004);
or U772 (N_772,In_2768,In_854);
or U773 (N_773,In_2215,In_1594);
xnor U774 (N_774,In_1213,In_2815);
nor U775 (N_775,In_2858,In_1347);
xnor U776 (N_776,In_1504,In_1674);
or U777 (N_777,In_1963,In_2537);
nor U778 (N_778,In_944,In_302);
nor U779 (N_779,In_1592,In_1726);
xnor U780 (N_780,In_2942,In_227);
and U781 (N_781,In_90,In_1360);
and U782 (N_782,In_681,In_1276);
xnor U783 (N_783,In_1891,In_1127);
or U784 (N_784,In_2952,In_1241);
and U785 (N_785,In_1613,In_178);
nor U786 (N_786,In_2841,In_2696);
nand U787 (N_787,In_2144,In_1356);
xnor U788 (N_788,In_2561,In_2267);
and U789 (N_789,In_965,In_1027);
nand U790 (N_790,In_1623,In_898);
xnor U791 (N_791,In_345,In_2246);
and U792 (N_792,In_2351,In_2584);
xnor U793 (N_793,In_1246,In_696);
nand U794 (N_794,In_461,In_2338);
and U795 (N_795,In_2157,In_2895);
nor U796 (N_796,In_978,In_328);
xnor U797 (N_797,In_2149,In_452);
or U798 (N_798,In_2145,In_601);
or U799 (N_799,In_532,In_30);
or U800 (N_800,In_2810,In_1384);
xor U801 (N_801,In_1640,In_1584);
xor U802 (N_802,In_2845,In_2756);
nor U803 (N_803,In_284,In_661);
xor U804 (N_804,In_1072,In_774);
nand U805 (N_805,In_2007,In_1167);
xor U806 (N_806,In_1537,In_2677);
nand U807 (N_807,In_2414,In_910);
or U808 (N_808,In_767,In_2568);
and U809 (N_809,In_2995,In_298);
or U810 (N_810,In_204,In_2269);
or U811 (N_811,In_1348,In_1115);
nand U812 (N_812,In_1342,In_765);
nand U813 (N_813,In_1340,In_1549);
nand U814 (N_814,In_2990,In_2405);
and U815 (N_815,In_798,In_1305);
nand U816 (N_816,In_1696,In_2536);
nand U817 (N_817,In_331,In_2578);
or U818 (N_818,In_1740,In_376);
or U819 (N_819,In_133,In_2052);
xnor U820 (N_820,In_928,In_1561);
and U821 (N_821,In_2368,In_342);
xnor U822 (N_822,In_2493,In_2819);
and U823 (N_823,In_75,In_947);
and U824 (N_824,In_2955,In_2265);
or U825 (N_825,In_1904,In_432);
nor U826 (N_826,In_1899,In_2928);
xnor U827 (N_827,In_2851,In_905);
nand U828 (N_828,In_1503,In_2639);
nor U829 (N_829,In_2406,In_1697);
or U830 (N_830,In_880,In_2844);
and U831 (N_831,In_2996,In_2685);
nand U832 (N_832,In_801,In_1002);
nor U833 (N_833,In_1730,In_621);
nand U834 (N_834,In_1544,In_2859);
xor U835 (N_835,In_1691,In_414);
or U836 (N_836,In_1063,In_2780);
and U837 (N_837,In_2386,In_307);
nor U838 (N_838,In_1997,In_1704);
or U839 (N_839,In_896,In_1094);
nor U840 (N_840,In_2085,In_58);
or U841 (N_841,In_2302,In_2576);
or U842 (N_842,In_2753,In_964);
and U843 (N_843,In_508,In_2909);
xor U844 (N_844,In_791,In_2433);
nand U845 (N_845,In_2866,In_597);
and U846 (N_846,In_394,In_1597);
nand U847 (N_847,In_665,In_1080);
and U848 (N_848,In_2439,In_2966);
nand U849 (N_849,In_2762,In_2273);
nor U850 (N_850,In_299,In_1259);
and U851 (N_851,In_1923,In_2074);
and U852 (N_852,In_1671,In_1104);
or U853 (N_853,In_1210,In_60);
or U854 (N_854,In_2619,In_1644);
nand U855 (N_855,In_1840,In_1709);
nand U856 (N_856,In_1568,In_1157);
and U857 (N_857,In_1861,In_2876);
nor U858 (N_858,In_131,In_784);
nor U859 (N_859,In_775,In_1983);
nand U860 (N_860,In_1165,In_448);
xor U861 (N_861,In_1439,In_344);
or U862 (N_862,In_454,In_1610);
nand U863 (N_863,In_22,In_1626);
xnor U864 (N_864,In_2783,In_844);
nor U865 (N_865,In_2840,In_571);
nor U866 (N_866,In_471,In_120);
nor U867 (N_867,In_455,In_1415);
xnor U868 (N_868,In_2341,In_1765);
nor U869 (N_869,In_2554,In_2315);
xor U870 (N_870,In_2035,In_424);
and U871 (N_871,In_2001,In_229);
nor U872 (N_872,In_2786,In_729);
or U873 (N_873,In_1748,In_37);
xnor U874 (N_874,In_1479,In_402);
or U875 (N_875,In_145,In_1048);
nand U876 (N_876,In_930,In_2751);
nand U877 (N_877,In_2902,In_123);
xor U878 (N_878,In_2172,In_1658);
and U879 (N_879,In_738,In_2726);
nand U880 (N_880,In_1812,In_2197);
nand U881 (N_881,In_743,In_2395);
or U882 (N_882,In_2008,In_2494);
and U883 (N_883,In_2842,In_1128);
or U884 (N_884,In_2355,In_112);
and U885 (N_885,In_2608,In_2340);
or U886 (N_886,In_1374,In_1061);
nand U887 (N_887,In_2701,In_1652);
and U888 (N_888,In_1170,In_2498);
nand U889 (N_889,In_16,In_796);
nor U890 (N_890,In_1791,In_2239);
or U891 (N_891,In_1445,In_1801);
xor U892 (N_892,In_1099,In_486);
nor U893 (N_893,In_1368,In_2374);
xnor U894 (N_894,In_1967,In_1131);
nand U895 (N_895,In_2675,In_1999);
xor U896 (N_896,In_1087,In_1343);
and U897 (N_897,In_2669,In_955);
nand U898 (N_898,In_1227,In_1930);
nor U899 (N_899,In_2954,In_42);
nor U900 (N_900,In_441,In_2229);
xor U901 (N_901,In_2667,In_2933);
and U902 (N_902,In_1363,In_958);
xor U903 (N_903,In_562,In_2367);
nand U904 (N_904,In_957,In_71);
xnor U905 (N_905,In_1685,In_2032);
xnor U906 (N_906,In_1714,In_637);
xnor U907 (N_907,In_2410,In_1829);
nor U908 (N_908,In_85,In_2673);
or U909 (N_909,In_1814,In_2878);
and U910 (N_910,In_1451,In_368);
xnor U911 (N_911,In_2735,In_1314);
nand U912 (N_912,In_1872,In_405);
nor U913 (N_913,In_1163,In_1047);
and U914 (N_914,In_1615,In_173);
xor U915 (N_915,In_951,In_1355);
nand U916 (N_916,In_851,In_2776);
nand U917 (N_917,In_684,In_1300);
xor U918 (N_918,In_377,In_2028);
or U919 (N_919,In_2187,In_1893);
and U920 (N_920,In_2218,In_2732);
nor U921 (N_921,In_1587,In_2941);
and U922 (N_922,In_763,In_1889);
nor U923 (N_923,In_1799,In_682);
or U924 (N_924,In_1387,In_268);
xor U925 (N_925,In_2274,In_1744);
xor U926 (N_926,In_314,In_1450);
and U927 (N_927,In_31,In_1229);
nand U928 (N_928,In_2835,In_82);
nand U929 (N_929,In_2147,In_2937);
xor U930 (N_930,In_2306,In_364);
xnor U931 (N_931,In_2799,In_521);
xnor U932 (N_932,In_1937,In_2644);
and U933 (N_933,In_283,In_1133);
and U934 (N_934,In_1496,In_2723);
xnor U935 (N_935,In_564,In_961);
xor U936 (N_936,In_39,In_1332);
or U937 (N_937,In_1572,In_193);
nand U938 (N_938,In_443,In_1781);
and U939 (N_939,In_579,In_2856);
or U940 (N_940,In_228,In_858);
or U941 (N_941,In_772,In_1067);
or U942 (N_942,In_1351,In_182);
and U943 (N_943,In_2193,In_887);
xor U944 (N_944,In_1070,In_2112);
xor U945 (N_945,In_2965,In_2573);
and U946 (N_946,In_820,In_379);
and U947 (N_947,In_1926,In_2789);
and U948 (N_948,In_1747,In_2752);
xnor U949 (N_949,In_1209,In_2347);
and U950 (N_950,In_1789,In_2609);
and U951 (N_951,In_498,In_2903);
nor U952 (N_952,In_1638,In_2853);
and U953 (N_953,In_2191,In_500);
or U954 (N_954,In_1388,In_2383);
nand U955 (N_955,In_607,In_199);
and U956 (N_956,In_1092,In_2163);
xnor U957 (N_957,In_2717,In_98);
nand U958 (N_958,In_2813,In_141);
or U959 (N_959,In_464,In_1371);
and U960 (N_960,In_2230,In_1153);
nand U961 (N_961,In_2012,In_914);
nand U962 (N_962,In_2073,In_2495);
nor U963 (N_963,In_1637,In_2058);
nand U964 (N_964,In_2716,In_972);
nor U965 (N_965,In_470,In_1688);
nor U966 (N_966,In_1328,In_1218);
nand U967 (N_967,In_2999,In_2686);
nor U968 (N_968,In_2524,In_561);
and U969 (N_969,In_208,In_1960);
nand U970 (N_970,In_861,In_2199);
nor U971 (N_971,In_1892,In_1166);
or U972 (N_972,In_1530,In_1651);
and U973 (N_973,In_2514,In_2984);
nor U974 (N_974,In_2350,In_240);
and U975 (N_975,In_2870,In_2897);
or U976 (N_976,In_2529,In_493);
nand U977 (N_977,In_1828,In_1759);
nor U978 (N_978,In_434,In_566);
nand U979 (N_979,In_2424,In_1214);
nor U980 (N_980,In_1604,In_2023);
nor U981 (N_981,In_749,In_2290);
xnor U982 (N_982,In_1818,In_2787);
or U983 (N_983,In_2460,In_1554);
and U984 (N_984,In_463,In_2871);
nand U985 (N_985,In_59,In_2334);
or U986 (N_986,In_205,In_44);
xnor U987 (N_987,In_40,In_1732);
nor U988 (N_988,In_2818,In_1558);
nor U989 (N_989,In_1951,In_2282);
or U990 (N_990,In_2492,In_1429);
nor U991 (N_991,In_2411,In_814);
nor U992 (N_992,In_2517,In_403);
or U993 (N_993,In_834,In_759);
nor U994 (N_994,In_2692,In_2469);
xnor U995 (N_995,In_1559,In_1447);
or U996 (N_996,In_45,In_109);
xnor U997 (N_997,In_683,In_2668);
xor U998 (N_998,In_269,In_1520);
xor U999 (N_999,In_633,In_2266);
or U1000 (N_1000,In_1689,In_1066);
xor U1001 (N_1001,In_2415,In_1947);
nand U1002 (N_1002,In_2176,In_1435);
xnor U1003 (N_1003,In_2119,In_2456);
nor U1004 (N_1004,In_1249,In_1036);
xor U1005 (N_1005,In_1589,In_2281);
or U1006 (N_1006,In_1353,In_1365);
xor U1007 (N_1007,In_1643,In_211);
xnor U1008 (N_1008,In_1304,In_2993);
and U1009 (N_1009,In_2868,In_237);
nor U1010 (N_1010,In_891,In_984);
nand U1011 (N_1011,In_2624,In_1456);
and U1012 (N_1012,In_126,In_391);
and U1013 (N_1013,In_1379,In_2555);
nand U1014 (N_1014,In_1320,In_32);
and U1015 (N_1015,In_2882,In_2185);
and U1016 (N_1016,In_1290,In_2428);
nand U1017 (N_1017,In_1735,In_994);
and U1018 (N_1018,In_2222,In_1119);
xnor U1019 (N_1019,In_224,In_1426);
xnor U1020 (N_1020,In_2271,In_1831);
nor U1021 (N_1021,In_553,In_630);
nor U1022 (N_1022,In_1877,In_613);
and U1023 (N_1023,In_2828,In_1124);
nand U1024 (N_1024,In_871,In_2730);
xnor U1025 (N_1025,In_885,In_1420);
xor U1026 (N_1026,In_1037,In_1541);
xor U1027 (N_1027,In_1323,In_628);
nor U1028 (N_1028,In_2500,In_53);
and U1029 (N_1029,In_1603,In_1091);
and U1030 (N_1030,In_2914,In_276);
nor U1031 (N_1031,In_2594,In_1835);
nand U1032 (N_1032,In_2689,In_100);
or U1033 (N_1033,In_974,In_1807);
or U1034 (N_1034,In_1630,In_292);
nand U1035 (N_1035,In_2587,In_617);
nor U1036 (N_1036,In_2358,In_2283);
xnor U1037 (N_1037,In_2324,In_2436);
and U1038 (N_1038,In_2505,In_523);
nand U1039 (N_1039,In_281,In_181);
nand U1040 (N_1040,In_1677,In_2663);
nand U1041 (N_1041,In_1289,In_2226);
or U1042 (N_1042,In_547,In_2319);
or U1043 (N_1043,In_1145,In_2834);
nand U1044 (N_1044,In_1021,In_134);
and U1045 (N_1045,In_1180,In_2138);
nand U1046 (N_1046,In_2688,In_1553);
nor U1047 (N_1047,In_1097,In_138);
nand U1048 (N_1048,In_266,In_1184);
and U1049 (N_1049,In_846,In_2188);
and U1050 (N_1050,In_2539,In_937);
and U1051 (N_1051,In_1001,In_2890);
and U1052 (N_1052,In_382,In_2015);
xnor U1053 (N_1053,In_1517,In_18);
and U1054 (N_1054,In_2440,In_1760);
nand U1055 (N_1055,In_2370,In_2640);
nor U1056 (N_1056,In_1910,In_221);
xor U1057 (N_1057,In_2479,In_2443);
xnor U1058 (N_1058,In_291,In_1647);
xor U1059 (N_1059,In_2627,In_2811);
nand U1060 (N_1060,In_191,In_274);
nand U1061 (N_1061,In_1076,In_2613);
xnor U1062 (N_1062,In_1971,In_2593);
nand U1063 (N_1063,In_2014,In_2263);
xor U1064 (N_1064,In_2575,In_1437);
xor U1065 (N_1065,In_638,In_973);
nand U1066 (N_1066,In_2132,In_705);
and U1067 (N_1067,In_1648,In_1248);
and U1068 (N_1068,In_589,In_216);
and U1069 (N_1069,In_1155,In_125);
and U1070 (N_1070,In_859,In_676);
or U1071 (N_1071,In_1143,In_581);
nand U1072 (N_1072,In_1361,In_1413);
nor U1073 (N_1073,In_1943,In_1260);
nor U1074 (N_1074,In_2749,In_2658);
nor U1075 (N_1075,In_386,In_1298);
nand U1076 (N_1076,In_1041,In_1672);
and U1077 (N_1077,In_2814,In_567);
nor U1078 (N_1078,In_1402,In_1251);
or U1079 (N_1079,In_2846,In_890);
and U1080 (N_1080,In_670,In_625);
or U1081 (N_1081,In_255,In_1302);
and U1082 (N_1082,In_1495,In_73);
nand U1083 (N_1083,In_2861,In_1023);
and U1084 (N_1084,In_57,In_1040);
and U1085 (N_1085,In_2917,In_277);
and U1086 (N_1086,In_2127,In_2150);
or U1087 (N_1087,In_1287,In_336);
nand U1088 (N_1088,In_2510,In_2332);
nor U1089 (N_1089,In_593,In_2335);
or U1090 (N_1090,In_1529,In_1069);
and U1091 (N_1091,In_1894,In_2497);
nor U1092 (N_1092,In_406,In_2261);
and U1093 (N_1093,In_2978,In_2729);
or U1094 (N_1094,In_400,In_2108);
nor U1095 (N_1095,In_169,In_536);
nand U1096 (N_1096,In_1649,In_2327);
nor U1097 (N_1097,In_886,In_2389);
nor U1098 (N_1098,In_2971,In_2380);
xnor U1099 (N_1099,In_1715,In_900);
or U1100 (N_1100,In_2872,In_1194);
and U1101 (N_1101,In_2107,In_1146);
xor U1102 (N_1102,In_1581,In_642);
nand U1103 (N_1103,In_2522,In_436);
nand U1104 (N_1104,In_2719,In_907);
or U1105 (N_1105,In_1389,In_1560);
or U1106 (N_1106,In_2705,In_1492);
xor U1107 (N_1107,In_720,In_781);
or U1108 (N_1108,In_2407,In_117);
xnor U1109 (N_1109,In_1906,In_2638);
and U1110 (N_1110,In_1896,In_1016);
nand U1111 (N_1111,In_1563,In_1854);
xnor U1112 (N_1112,In_1286,In_627);
xnor U1113 (N_1113,In_1653,In_1438);
and U1114 (N_1114,In_917,In_2257);
xor U1115 (N_1115,In_1148,In_787);
nor U1116 (N_1116,In_375,In_260);
or U1117 (N_1117,In_474,In_1953);
and U1118 (N_1118,In_2067,In_2939);
nand U1119 (N_1119,In_1945,In_2217);
xnor U1120 (N_1120,In_1622,In_161);
xor U1121 (N_1121,In_1845,In_2446);
nand U1122 (N_1122,In_1383,In_1083);
xor U1123 (N_1123,In_1331,In_2682);
nor U1124 (N_1124,In_746,In_383);
or U1125 (N_1125,In_1139,In_2745);
nand U1126 (N_1126,In_1987,In_1513);
nor U1127 (N_1127,In_1207,In_1724);
nand U1128 (N_1128,In_2921,In_1109);
and U1129 (N_1129,In_985,In_1948);
nor U1130 (N_1130,In_1283,In_1629);
nor U1131 (N_1131,In_190,In_2125);
or U1132 (N_1132,In_1030,In_171);
and U1133 (N_1133,In_1416,In_862);
nand U1134 (N_1134,In_2551,In_346);
and U1135 (N_1135,In_2739,In_1986);
or U1136 (N_1136,In_1012,In_5);
or U1137 (N_1137,In_1700,In_1841);
or U1138 (N_1138,In_2399,In_1452);
or U1139 (N_1139,In_1369,In_1313);
nor U1140 (N_1140,In_2946,In_1692);
xor U1141 (N_1141,In_1427,In_1733);
or U1142 (N_1142,In_713,In_522);
nor U1143 (N_1143,In_1263,In_2721);
and U1144 (N_1144,In_1204,In_1516);
xor U1145 (N_1145,In_1309,In_1345);
nor U1146 (N_1146,In_425,In_870);
nor U1147 (N_1147,In_1605,In_1694);
and U1148 (N_1148,In_129,In_2451);
nor U1149 (N_1149,In_2472,In_691);
xor U1150 (N_1150,In_2943,In_747);
or U1151 (N_1151,In_2896,In_1187);
and U1152 (N_1152,In_1506,In_1627);
xor U1153 (N_1153,In_559,In_1756);
or U1154 (N_1154,In_214,In_1551);
and U1155 (N_1155,In_1272,In_1256);
nor U1156 (N_1156,In_1464,In_2204);
nor U1157 (N_1157,In_1660,In_159);
xnor U1158 (N_1158,In_2179,In_797);
and U1159 (N_1159,In_2331,In_2173);
nand U1160 (N_1160,In_1741,In_515);
or U1161 (N_1161,In_373,In_1770);
and U1162 (N_1162,In_2270,In_381);
nor U1163 (N_1163,In_520,In_2617);
and U1164 (N_1164,In_941,In_1550);
nor U1165 (N_1165,In_2033,In_873);
and U1166 (N_1166,In_1982,In_487);
or U1167 (N_1167,In_842,In_1855);
and U1168 (N_1168,In_1039,In_1885);
or U1169 (N_1169,In_1294,In_2225);
xnor U1170 (N_1170,In_1907,In_27);
nor U1171 (N_1171,In_287,In_2784);
or U1172 (N_1172,In_1946,In_245);
nor U1173 (N_1173,In_1534,In_1777);
xor U1174 (N_1174,In_2637,In_1614);
xor U1175 (N_1175,In_1718,In_770);
nor U1176 (N_1176,In_2357,In_2731);
or U1177 (N_1177,In_435,In_1920);
xnor U1178 (N_1178,In_370,In_2591);
nand U1179 (N_1179,In_812,In_1519);
nand U1180 (N_1180,In_2131,In_518);
xor U1181 (N_1181,In_761,In_2117);
and U1182 (N_1182,In_1195,In_2251);
nor U1183 (N_1183,In_1422,In_360);
nor U1184 (N_1184,In_687,In_971);
and U1185 (N_1185,In_2727,In_1507);
or U1186 (N_1186,In_1357,In_1583);
or U1187 (N_1187,In_2444,In_1319);
xor U1188 (N_1188,In_2235,In_1330);
nand U1189 (N_1189,In_309,In_701);
nor U1190 (N_1190,In_1334,In_2906);
and U1191 (N_1191,In_2746,In_2116);
xor U1192 (N_1192,In_2013,In_751);
or U1193 (N_1193,In_494,In_388);
nand U1194 (N_1194,In_755,In_1089);
nor U1195 (N_1195,In_735,In_195);
or U1196 (N_1196,In_35,In_903);
xnor U1197 (N_1197,In_1729,In_1008);
xnor U1198 (N_1198,In_1639,In_2097);
nor U1199 (N_1199,In_92,In_1406);
and U1200 (N_1200,In_807,In_185);
and U1201 (N_1201,In_2582,In_2031);
nor U1202 (N_1202,In_2711,In_2718);
xor U1203 (N_1203,In_1720,In_1250);
xnor U1204 (N_1204,In_1475,In_725);
nor U1205 (N_1205,In_2769,In_1954);
nor U1206 (N_1206,In_2936,In_2388);
xnor U1207 (N_1207,In_2636,In_1778);
and U1208 (N_1208,In_2234,In_203);
xor U1209 (N_1209,In_1273,In_2133);
and U1210 (N_1210,In_1005,In_1625);
and U1211 (N_1211,In_2280,In_1395);
and U1212 (N_1212,In_1284,In_813);
and U1213 (N_1213,In_2883,In_1088);
nor U1214 (N_1214,In_2098,In_2646);
xnor U1215 (N_1215,In_2244,In_1751);
nand U1216 (N_1216,In_663,In_2195);
and U1217 (N_1217,In_192,In_2105);
xnor U1218 (N_1218,In_177,In_726);
xor U1219 (N_1219,In_2036,In_1000);
nand U1220 (N_1220,In_1883,In_949);
nor U1221 (N_1221,In_2101,In_2275);
xnor U1222 (N_1222,In_217,In_578);
xor U1223 (N_1223,In_151,In_1574);
nor U1224 (N_1224,In_590,In_1147);
xnor U1225 (N_1225,In_800,In_1705);
and U1226 (N_1226,In_2899,In_1667);
or U1227 (N_1227,In_1171,In_715);
xnor U1228 (N_1228,In_2693,In_2720);
nor U1229 (N_1229,In_1753,In_1573);
and U1230 (N_1230,In_1055,In_433);
xnor U1231 (N_1231,In_305,In_473);
nor U1232 (N_1232,In_2805,In_1113);
xor U1233 (N_1233,In_516,In_1035);
or U1234 (N_1234,In_393,In_916);
nand U1235 (N_1235,In_1460,In_1727);
xor U1236 (N_1236,In_1370,In_519);
or U1237 (N_1237,In_2053,In_744);
and U1238 (N_1238,In_2363,In_679);
nor U1239 (N_1239,In_2310,In_1188);
xor U1240 (N_1240,In_6,In_2253);
xnor U1241 (N_1241,In_2430,In_2626);
and U1242 (N_1242,In_671,In_2760);
nor U1243 (N_1243,In_395,In_1832);
and U1244 (N_1244,In_2772,In_2352);
xnor U1245 (N_1245,In_2272,In_2198);
and U1246 (N_1246,In_824,In_2384);
nor U1247 (N_1247,In_577,In_2151);
and U1248 (N_1248,In_2986,In_1746);
xnor U1249 (N_1249,In_1301,In_1137);
xnor U1250 (N_1250,In_512,In_462);
xor U1251 (N_1251,In_252,In_1665);
nand U1252 (N_1252,In_677,In_401);
or U1253 (N_1253,In_2982,In_2964);
xnor U1254 (N_1254,In_2159,In_316);
and U1255 (N_1255,In_43,In_2623);
and U1256 (N_1256,In_752,In_2572);
and U1257 (N_1257,In_2804,In_450);
or U1258 (N_1258,In_708,In_2102);
nor U1259 (N_1259,In_1175,In_764);
or U1260 (N_1260,In_2775,In_38);
nand U1261 (N_1261,In_2887,In_612);
nor U1262 (N_1262,In_2629,In_753);
xor U1263 (N_1263,In_2401,In_1310);
xor U1264 (N_1264,In_137,In_490);
or U1265 (N_1265,In_64,In_2643);
nor U1266 (N_1266,In_1045,In_2180);
and U1267 (N_1267,In_932,In_2782);
nor U1268 (N_1268,In_2788,In_1279);
or U1269 (N_1269,In_598,In_2607);
nor U1270 (N_1270,In_279,In_2006);
xnor U1271 (N_1271,In_2072,In_107);
or U1272 (N_1272,In_1757,In_1934);
or U1273 (N_1273,In_2516,In_2512);
and U1274 (N_1274,In_1949,In_837);
nor U1275 (N_1275,In_2655,In_717);
xnor U1276 (N_1276,In_591,In_2757);
xnor U1277 (N_1277,In_803,In_1862);
nand U1278 (N_1278,In_779,In_1505);
xnor U1279 (N_1279,In_89,In_1380);
nor U1280 (N_1280,In_1588,In_2827);
and U1281 (N_1281,In_1890,In_2061);
xnor U1282 (N_1282,In_1150,In_1489);
nor U1283 (N_1283,In_1703,In_860);
nor U1284 (N_1284,In_1575,In_1565);
nor U1285 (N_1285,In_1082,In_2285);
or U1286 (N_1286,In_2886,In_1257);
xor U1287 (N_1287,In_1154,In_1878);
or U1288 (N_1288,In_2901,In_2562);
and U1289 (N_1289,In_1085,In_2295);
and U1290 (N_1290,In_2438,In_2009);
xnor U1291 (N_1291,In_2140,In_2503);
and U1292 (N_1292,In_2461,In_1825);
and U1293 (N_1293,In_2634,In_2264);
xor U1294 (N_1294,In_1499,In_2957);
nor U1295 (N_1295,In_975,In_1749);
nor U1296 (N_1296,In_2476,In_460);
nor U1297 (N_1297,In_1185,In_657);
or U1298 (N_1298,In_1737,In_1964);
xnor U1299 (N_1299,In_1636,In_2240);
and U1300 (N_1300,In_1545,In_1326);
nand U1301 (N_1301,In_1917,In_1071);
xnor U1302 (N_1302,In_2016,In_2821);
nor U1303 (N_1303,In_673,In_1430);
or U1304 (N_1304,In_1483,In_1366);
or U1305 (N_1305,In_2342,In_1942);
and U1306 (N_1306,In_289,In_103);
or U1307 (N_1307,In_2968,In_510);
nor U1308 (N_1308,In_2598,In_792);
xnor U1309 (N_1309,In_232,In_1776);
xor U1310 (N_1310,In_249,In_1676);
and U1311 (N_1311,In_575,In_1308);
or U1312 (N_1312,In_1373,In_234);
and U1313 (N_1313,In_2231,In_2635);
nand U1314 (N_1314,In_1199,In_2949);
nand U1315 (N_1315,In_1916,In_1488);
xnor U1316 (N_1316,In_408,In_902);
and U1317 (N_1317,In_200,In_2005);
nor U1318 (N_1318,In_766,In_2387);
nand U1319 (N_1319,In_343,In_2940);
nand U1320 (N_1320,In_273,In_1424);
or U1321 (N_1321,In_2308,In_2030);
or U1322 (N_1322,In_1641,In_1875);
xor U1323 (N_1323,In_223,In_1540);
nor U1324 (N_1324,In_1682,In_248);
or U1325 (N_1325,In_437,In_2651);
or U1326 (N_1326,In_1130,In_2650);
xnor U1327 (N_1327,In_1114,In_1243);
nand U1328 (N_1328,In_139,In_2022);
or U1329 (N_1329,In_2850,In_1410);
or U1330 (N_1330,In_1763,In_2314);
nor U1331 (N_1331,In_1240,In_1403);
or U1332 (N_1332,In_1538,In_127);
nor U1333 (N_1333,In_2465,In_2679);
nor U1334 (N_1334,In_2224,In_2482);
nor U1335 (N_1335,In_2556,In_1261);
or U1336 (N_1336,In_1975,In_0);
or U1337 (N_1337,In_1412,In_398);
nand U1338 (N_1338,In_1998,In_939);
nor U1339 (N_1339,In_458,In_2427);
and U1340 (N_1340,In_10,In_2018);
nand U1341 (N_1341,In_271,In_2312);
and U1342 (N_1342,In_1392,In_1950);
and U1343 (N_1343,In_2247,In_1102);
and U1344 (N_1344,In_583,In_179);
xor U1345 (N_1345,In_845,In_2956);
or U1346 (N_1346,In_1337,In_2243);
xnor U1347 (N_1347,In_2702,In_546);
or U1348 (N_1348,In_847,In_2019);
nor U1349 (N_1349,In_1225,In_1327);
or U1350 (N_1350,In_884,In_2214);
nor U1351 (N_1351,In_466,In_61);
nor U1352 (N_1352,In_87,In_2241);
or U1353 (N_1353,In_496,In_25);
nor U1354 (N_1354,In_1270,In_1547);
and U1355 (N_1355,In_2725,In_280);
or U1356 (N_1356,In_258,In_104);
nand U1357 (N_1357,In_2094,In_1698);
or U1358 (N_1358,In_2262,In_2963);
and U1359 (N_1359,In_1231,In_2961);
nand U1360 (N_1360,In_2100,In_1941);
and U1361 (N_1361,In_1673,In_2541);
or U1362 (N_1362,In_996,In_165);
or U1363 (N_1363,In_2967,In_1490);
xnor U1364 (N_1364,In_2063,In_595);
and U1365 (N_1365,In_768,In_2291);
and U1366 (N_1366,In_113,In_242);
or U1367 (N_1367,In_24,In_351);
nor U1368 (N_1368,In_251,In_568);
xnor U1369 (N_1369,In_15,In_2839);
or U1370 (N_1370,In_1400,In_2722);
nand U1371 (N_1371,In_2137,In_2945);
nor U1372 (N_1372,In_874,In_1386);
and U1373 (N_1373,In_1766,In_2622);
xor U1374 (N_1374,In_869,In_2075);
nor U1375 (N_1375,In_1985,In_629);
or U1376 (N_1376,In_2699,In_1046);
nand U1377 (N_1377,In_1936,In_1458);
or U1378 (N_1378,In_1842,In_2301);
or U1379 (N_1379,In_2743,In_172);
nor U1380 (N_1380,In_1118,In_2926);
nand U1381 (N_1381,In_155,In_2605);
and U1382 (N_1382,In_514,In_2974);
and U1383 (N_1383,In_1695,In_431);
and U1384 (N_1384,In_1242,In_2843);
xnor U1385 (N_1385,In_827,In_2944);
xor U1386 (N_1386,In_62,In_664);
nand U1387 (N_1387,In_703,In_780);
nand U1388 (N_1388,In_2904,In_1432);
and U1389 (N_1389,In_1525,In_901);
nand U1390 (N_1390,In_1487,In_2630);
nand U1391 (N_1391,In_517,In_576);
and U1392 (N_1392,In_714,In_1933);
xor U1393 (N_1393,In_1911,In_1536);
or U1394 (N_1394,In_1783,In_2011);
xnor U1395 (N_1395,In_921,In_1028);
nor U1396 (N_1396,In_2523,In_2513);
and U1397 (N_1397,In_34,In_616);
xnor U1398 (N_1398,In_210,In_1659);
nor U1399 (N_1399,In_12,In_1335);
and U1400 (N_1400,In_2287,In_2740);
nor U1401 (N_1401,In_700,In_1903);
nand U1402 (N_1402,In_423,In_2459);
or U1403 (N_1403,In_2535,In_1815);
and U1404 (N_1404,In_1346,In_41);
nand U1405 (N_1405,In_1619,In_2496);
and U1406 (N_1406,In_2981,In_188);
and U1407 (N_1407,In_1077,In_389);
nand U1408 (N_1408,In_2659,In_1358);
xor U1409 (N_1409,In_2507,In_2863);
or U1410 (N_1410,In_1654,In_2437);
or U1411 (N_1411,In_950,In_2397);
nand U1412 (N_1412,In_1152,In_2664);
xor U1413 (N_1413,In_2704,In_976);
nor U1414 (N_1414,In_1098,In_261);
nor U1415 (N_1415,In_2237,In_2369);
nand U1416 (N_1416,In_830,In_1816);
or U1417 (N_1417,In_2379,In_938);
nand U1418 (N_1418,In_742,In_1898);
nand U1419 (N_1419,In_2807,In_1570);
nand U1420 (N_1420,In_875,In_1657);
xor U1421 (N_1421,In_659,In_741);
xnor U1422 (N_1422,In_1527,In_2110);
nor U1423 (N_1423,In_231,In_507);
xnor U1424 (N_1424,In_2170,In_2656);
and U1425 (N_1425,In_1602,In_1465);
nor U1426 (N_1426,In_2468,In_718);
or U1427 (N_1427,In_2502,In_643);
xor U1428 (N_1428,In_2838,In_757);
and U1429 (N_1429,In_2034,In_2864);
or U1430 (N_1430,In_105,In_2911);
nor U1431 (N_1431,In_1810,In_1557);
or U1432 (N_1432,In_451,In_2066);
and U1433 (N_1433,In_2354,In_2687);
xnor U1434 (N_1434,In_2148,In_243);
nand U1435 (N_1435,In_147,In_1690);
nor U1436 (N_1436,In_1278,In_993);
and U1437 (N_1437,In_1909,In_2396);
xor U1438 (N_1438,In_2181,In_157);
xnor U1439 (N_1439,In_256,In_2364);
nor U1440 (N_1440,In_1338,In_840);
and U1441 (N_1441,In_69,In_2356);
nor U1442 (N_1442,In_1754,In_1785);
nand U1443 (N_1443,In_1768,In_160);
or U1444 (N_1444,In_2024,In_2543);
or U1445 (N_1445,In_74,In_2773);
nand U1446 (N_1446,In_626,In_47);
and U1447 (N_1447,In_1992,In_1932);
nor U1448 (N_1448,In_2346,In_704);
xnor U1449 (N_1449,In_197,In_2980);
xnor U1450 (N_1450,In_2223,In_122);
xor U1451 (N_1451,In_2604,In_1033);
nor U1452 (N_1452,In_2824,In_2429);
xor U1453 (N_1453,In_2975,In_1441);
xnor U1454 (N_1454,In_2734,In_674);
nor U1455 (N_1455,In_2130,In_694);
nor U1456 (N_1456,In_2408,In_2544);
nand U1457 (N_1457,In_1869,In_2455);
nor U1458 (N_1458,In_348,In_2120);
and U1459 (N_1459,In_1811,In_2820);
nor U1460 (N_1460,In_2345,In_2055);
or U1461 (N_1461,In_2184,In_2299);
nor U1462 (N_1462,In_1453,In_888);
or U1463 (N_1463,In_690,In_2558);
xor U1464 (N_1464,In_267,In_1117);
xor U1465 (N_1465,In_2583,In_2042);
and U1466 (N_1466,In_2337,In_1784);
nor U1467 (N_1467,In_2091,In_2930);
nor U1468 (N_1468,In_1280,In_983);
nand U1469 (N_1469,In_556,In_1523);
nor U1470 (N_1470,In_1755,In_585);
and U1471 (N_1471,In_1459,In_545);
xnor U1472 (N_1472,In_1663,In_235);
xnor U1473 (N_1473,In_469,In_2781);
and U1474 (N_1474,In_2391,In_927);
nand U1475 (N_1475,In_1731,In_312);
or U1476 (N_1476,In_4,In_86);
xor U1477 (N_1477,In_1612,In_2403);
and U1478 (N_1478,In_1699,In_497);
or U1479 (N_1479,In_2442,In_2779);
or U1480 (N_1480,In_656,In_2645);
nand U1481 (N_1481,In_1362,In_70);
nand U1482 (N_1482,In_259,In_485);
nand U1483 (N_1483,In_2884,In_2242);
and U1484 (N_1484,In_1693,In_716);
and U1485 (N_1485,In_540,In_2453);
xnor U1486 (N_1486,In_2546,In_2457);
xor U1487 (N_1487,In_1833,In_2079);
and U1488 (N_1488,In_36,In_878);
and U1489 (N_1489,In_644,In_2707);
xor U1490 (N_1490,In_332,In_969);
nor U1491 (N_1491,In_365,In_640);
nand U1492 (N_1492,In_1723,In_1469);
or U1493 (N_1493,In_660,In_301);
nand U1494 (N_1494,In_413,In_2361);
nor U1495 (N_1495,In_646,In_2580);
or U1496 (N_1496,In_286,In_1275);
and U1497 (N_1497,In_2972,In_818);
nand U1498 (N_1498,In_821,In_1007);
nand U1499 (N_1499,In_341,In_2951);
or U1500 (N_1500,In_1675,In_2042);
or U1501 (N_1501,In_2662,In_1479);
nor U1502 (N_1502,In_151,In_1806);
or U1503 (N_1503,In_1501,In_1688);
nor U1504 (N_1504,In_2565,In_398);
and U1505 (N_1505,In_2061,In_2416);
xnor U1506 (N_1506,In_1734,In_795);
or U1507 (N_1507,In_2329,In_1009);
nor U1508 (N_1508,In_1195,In_1149);
nand U1509 (N_1509,In_1277,In_741);
nor U1510 (N_1510,In_634,In_371);
nor U1511 (N_1511,In_2398,In_1744);
or U1512 (N_1512,In_2921,In_2416);
nor U1513 (N_1513,In_1355,In_1391);
xor U1514 (N_1514,In_1919,In_1964);
and U1515 (N_1515,In_1992,In_1522);
or U1516 (N_1516,In_2533,In_582);
or U1517 (N_1517,In_624,In_825);
nand U1518 (N_1518,In_344,In_929);
xor U1519 (N_1519,In_1771,In_2147);
or U1520 (N_1520,In_1887,In_420);
nand U1521 (N_1521,In_2699,In_2312);
nand U1522 (N_1522,In_2443,In_776);
nor U1523 (N_1523,In_721,In_2583);
nand U1524 (N_1524,In_62,In_1667);
nor U1525 (N_1525,In_2436,In_6);
nor U1526 (N_1526,In_2530,In_65);
nor U1527 (N_1527,In_813,In_2427);
nand U1528 (N_1528,In_353,In_1241);
and U1529 (N_1529,In_1670,In_19);
nor U1530 (N_1530,In_2106,In_2051);
and U1531 (N_1531,In_1966,In_1036);
nand U1532 (N_1532,In_2036,In_773);
and U1533 (N_1533,In_2553,In_2486);
nand U1534 (N_1534,In_1243,In_2207);
nand U1535 (N_1535,In_1266,In_1837);
nor U1536 (N_1536,In_878,In_2588);
xor U1537 (N_1537,In_1345,In_2122);
nand U1538 (N_1538,In_199,In_1314);
nor U1539 (N_1539,In_751,In_2938);
and U1540 (N_1540,In_1681,In_1289);
nor U1541 (N_1541,In_2617,In_1251);
or U1542 (N_1542,In_2718,In_1858);
nand U1543 (N_1543,In_184,In_595);
nor U1544 (N_1544,In_1782,In_2943);
or U1545 (N_1545,In_1112,In_1082);
or U1546 (N_1546,In_1705,In_2473);
and U1547 (N_1547,In_1378,In_2536);
nor U1548 (N_1548,In_2957,In_561);
nand U1549 (N_1549,In_311,In_1010);
or U1550 (N_1550,In_759,In_1644);
or U1551 (N_1551,In_2860,In_36);
or U1552 (N_1552,In_1047,In_2906);
nand U1553 (N_1553,In_1847,In_735);
and U1554 (N_1554,In_11,In_1940);
xor U1555 (N_1555,In_834,In_2722);
or U1556 (N_1556,In_1846,In_2875);
nor U1557 (N_1557,In_2385,In_1574);
and U1558 (N_1558,In_2293,In_1226);
or U1559 (N_1559,In_1132,In_2770);
nand U1560 (N_1560,In_409,In_418);
nor U1561 (N_1561,In_1492,In_982);
and U1562 (N_1562,In_1388,In_2854);
xnor U1563 (N_1563,In_772,In_2153);
and U1564 (N_1564,In_1649,In_532);
nand U1565 (N_1565,In_887,In_1892);
or U1566 (N_1566,In_2590,In_2223);
nand U1567 (N_1567,In_101,In_31);
nor U1568 (N_1568,In_2675,In_2091);
nand U1569 (N_1569,In_30,In_1689);
nand U1570 (N_1570,In_2190,In_2383);
xor U1571 (N_1571,In_2188,In_461);
and U1572 (N_1572,In_1831,In_964);
nand U1573 (N_1573,In_1788,In_11);
nand U1574 (N_1574,In_2971,In_2297);
nor U1575 (N_1575,In_2041,In_227);
xnor U1576 (N_1576,In_1285,In_2446);
nand U1577 (N_1577,In_2934,In_2649);
or U1578 (N_1578,In_284,In_747);
nor U1579 (N_1579,In_879,In_1737);
xor U1580 (N_1580,In_425,In_198);
and U1581 (N_1581,In_2112,In_2643);
nand U1582 (N_1582,In_2604,In_1192);
and U1583 (N_1583,In_1805,In_1082);
and U1584 (N_1584,In_1592,In_892);
xnor U1585 (N_1585,In_2612,In_1578);
or U1586 (N_1586,In_1864,In_1377);
or U1587 (N_1587,In_1146,In_998);
nand U1588 (N_1588,In_229,In_257);
and U1589 (N_1589,In_2215,In_2477);
and U1590 (N_1590,In_2877,In_1340);
and U1591 (N_1591,In_265,In_2418);
and U1592 (N_1592,In_2921,In_2783);
nor U1593 (N_1593,In_334,In_2050);
or U1594 (N_1594,In_2936,In_1041);
xor U1595 (N_1595,In_933,In_2689);
nor U1596 (N_1596,In_1126,In_2267);
and U1597 (N_1597,In_2756,In_839);
nor U1598 (N_1598,In_2883,In_360);
xnor U1599 (N_1599,In_27,In_317);
nor U1600 (N_1600,In_2599,In_1194);
or U1601 (N_1601,In_2197,In_1272);
or U1602 (N_1602,In_1496,In_1120);
xor U1603 (N_1603,In_1148,In_2245);
nor U1604 (N_1604,In_754,In_205);
nor U1605 (N_1605,In_2588,In_2493);
or U1606 (N_1606,In_2746,In_975);
nor U1607 (N_1607,In_1231,In_945);
xnor U1608 (N_1608,In_2368,In_1649);
nand U1609 (N_1609,In_2419,In_1472);
nand U1610 (N_1610,In_1312,In_1090);
and U1611 (N_1611,In_2516,In_702);
or U1612 (N_1612,In_431,In_271);
xnor U1613 (N_1613,In_1342,In_1948);
or U1614 (N_1614,In_2853,In_874);
nand U1615 (N_1615,In_2198,In_2933);
or U1616 (N_1616,In_1992,In_1830);
or U1617 (N_1617,In_1339,In_91);
nand U1618 (N_1618,In_2735,In_2693);
nor U1619 (N_1619,In_781,In_2064);
or U1620 (N_1620,In_1020,In_2368);
xnor U1621 (N_1621,In_805,In_2133);
or U1622 (N_1622,In_2950,In_1950);
nor U1623 (N_1623,In_1691,In_288);
nand U1624 (N_1624,In_381,In_748);
nor U1625 (N_1625,In_1971,In_192);
nor U1626 (N_1626,In_1059,In_1945);
and U1627 (N_1627,In_2173,In_215);
nand U1628 (N_1628,In_1187,In_1532);
nor U1629 (N_1629,In_291,In_1626);
and U1630 (N_1630,In_1388,In_1057);
nand U1631 (N_1631,In_2825,In_1674);
or U1632 (N_1632,In_2156,In_2559);
and U1633 (N_1633,In_633,In_1830);
and U1634 (N_1634,In_2659,In_877);
and U1635 (N_1635,In_79,In_1908);
and U1636 (N_1636,In_778,In_1655);
nand U1637 (N_1637,In_166,In_162);
or U1638 (N_1638,In_0,In_1898);
nand U1639 (N_1639,In_1220,In_311);
xor U1640 (N_1640,In_1594,In_2454);
xnor U1641 (N_1641,In_1099,In_567);
xnor U1642 (N_1642,In_1409,In_1442);
nor U1643 (N_1643,In_1268,In_1737);
xor U1644 (N_1644,In_1285,In_2440);
or U1645 (N_1645,In_852,In_2274);
or U1646 (N_1646,In_611,In_797);
nand U1647 (N_1647,In_80,In_1346);
nand U1648 (N_1648,In_1231,In_1797);
nor U1649 (N_1649,In_2157,In_2897);
xnor U1650 (N_1650,In_101,In_1417);
and U1651 (N_1651,In_1166,In_919);
or U1652 (N_1652,In_2049,In_2475);
xor U1653 (N_1653,In_1977,In_912);
or U1654 (N_1654,In_219,In_2786);
and U1655 (N_1655,In_685,In_2463);
and U1656 (N_1656,In_770,In_2707);
or U1657 (N_1657,In_2973,In_1610);
nor U1658 (N_1658,In_1424,In_819);
and U1659 (N_1659,In_70,In_1419);
or U1660 (N_1660,In_2361,In_1865);
xor U1661 (N_1661,In_1595,In_2866);
nand U1662 (N_1662,In_1977,In_914);
xor U1663 (N_1663,In_2957,In_2565);
nand U1664 (N_1664,In_2943,In_721);
nor U1665 (N_1665,In_1191,In_569);
nand U1666 (N_1666,In_2694,In_70);
nand U1667 (N_1667,In_25,In_1772);
xnor U1668 (N_1668,In_51,In_1215);
and U1669 (N_1669,In_523,In_2253);
nand U1670 (N_1670,In_1234,In_2177);
or U1671 (N_1671,In_1817,In_227);
or U1672 (N_1672,In_2567,In_1238);
nand U1673 (N_1673,In_2830,In_368);
or U1674 (N_1674,In_2719,In_1997);
or U1675 (N_1675,In_1359,In_1926);
nand U1676 (N_1676,In_1199,In_2818);
and U1677 (N_1677,In_2750,In_2783);
and U1678 (N_1678,In_2048,In_481);
xor U1679 (N_1679,In_2577,In_309);
nor U1680 (N_1680,In_1023,In_2949);
nand U1681 (N_1681,In_926,In_1961);
nand U1682 (N_1682,In_902,In_2069);
nand U1683 (N_1683,In_2665,In_471);
nand U1684 (N_1684,In_2987,In_74);
and U1685 (N_1685,In_2300,In_1469);
nand U1686 (N_1686,In_485,In_213);
nor U1687 (N_1687,In_2315,In_2705);
nor U1688 (N_1688,In_2632,In_2291);
and U1689 (N_1689,In_297,In_2485);
xnor U1690 (N_1690,In_1749,In_1955);
nand U1691 (N_1691,In_2409,In_258);
nor U1692 (N_1692,In_266,In_1869);
xnor U1693 (N_1693,In_1899,In_2052);
or U1694 (N_1694,In_509,In_2102);
and U1695 (N_1695,In_2700,In_992);
or U1696 (N_1696,In_1905,In_354);
xor U1697 (N_1697,In_1154,In_2915);
or U1698 (N_1698,In_2823,In_1140);
or U1699 (N_1699,In_1936,In_480);
or U1700 (N_1700,In_2800,In_2713);
nor U1701 (N_1701,In_2687,In_2413);
xor U1702 (N_1702,In_215,In_470);
nand U1703 (N_1703,In_2456,In_1583);
or U1704 (N_1704,In_2140,In_1956);
or U1705 (N_1705,In_2590,In_2152);
nor U1706 (N_1706,In_1651,In_880);
and U1707 (N_1707,In_2372,In_1001);
or U1708 (N_1708,In_2075,In_2602);
and U1709 (N_1709,In_957,In_476);
or U1710 (N_1710,In_1150,In_516);
or U1711 (N_1711,In_1320,In_2802);
xnor U1712 (N_1712,In_315,In_2658);
nor U1713 (N_1713,In_1508,In_484);
nand U1714 (N_1714,In_1846,In_330);
and U1715 (N_1715,In_1154,In_2183);
nand U1716 (N_1716,In_2105,In_951);
xor U1717 (N_1717,In_2756,In_516);
xnor U1718 (N_1718,In_2752,In_944);
nor U1719 (N_1719,In_1205,In_2386);
xnor U1720 (N_1720,In_1218,In_2810);
xor U1721 (N_1721,In_2960,In_2929);
and U1722 (N_1722,In_1062,In_996);
nor U1723 (N_1723,In_1164,In_352);
nor U1724 (N_1724,In_1993,In_2108);
nor U1725 (N_1725,In_2224,In_2372);
xnor U1726 (N_1726,In_1759,In_1888);
or U1727 (N_1727,In_2915,In_1920);
or U1728 (N_1728,In_494,In_1266);
xnor U1729 (N_1729,In_2838,In_2062);
nor U1730 (N_1730,In_911,In_39);
and U1731 (N_1731,In_2884,In_2586);
xor U1732 (N_1732,In_1256,In_1050);
xor U1733 (N_1733,In_1257,In_1886);
and U1734 (N_1734,In_105,In_5);
xnor U1735 (N_1735,In_1439,In_558);
nand U1736 (N_1736,In_878,In_2417);
or U1737 (N_1737,In_273,In_1934);
or U1738 (N_1738,In_1023,In_1010);
or U1739 (N_1739,In_678,In_2124);
xnor U1740 (N_1740,In_420,In_779);
or U1741 (N_1741,In_2615,In_2888);
or U1742 (N_1742,In_2308,In_2078);
or U1743 (N_1743,In_2456,In_1202);
nand U1744 (N_1744,In_562,In_402);
nand U1745 (N_1745,In_25,In_808);
xnor U1746 (N_1746,In_2406,In_1802);
or U1747 (N_1747,In_423,In_2266);
xnor U1748 (N_1748,In_918,In_2701);
xnor U1749 (N_1749,In_1655,In_862);
and U1750 (N_1750,In_2298,In_1552);
xor U1751 (N_1751,In_1008,In_273);
or U1752 (N_1752,In_523,In_382);
or U1753 (N_1753,In_1374,In_1342);
or U1754 (N_1754,In_465,In_2485);
or U1755 (N_1755,In_471,In_1432);
and U1756 (N_1756,In_1890,In_657);
nand U1757 (N_1757,In_1311,In_2191);
nand U1758 (N_1758,In_2934,In_903);
nand U1759 (N_1759,In_1622,In_293);
or U1760 (N_1760,In_438,In_2792);
or U1761 (N_1761,In_257,In_702);
nor U1762 (N_1762,In_1403,In_1306);
and U1763 (N_1763,In_1815,In_2709);
and U1764 (N_1764,In_1057,In_884);
nand U1765 (N_1765,In_588,In_2306);
or U1766 (N_1766,In_2063,In_859);
nand U1767 (N_1767,In_1183,In_1573);
and U1768 (N_1768,In_1562,In_2828);
and U1769 (N_1769,In_224,In_6);
and U1770 (N_1770,In_998,In_1901);
xor U1771 (N_1771,In_418,In_395);
and U1772 (N_1772,In_1388,In_1975);
and U1773 (N_1773,In_1607,In_1351);
or U1774 (N_1774,In_377,In_497);
nor U1775 (N_1775,In_1107,In_2198);
nand U1776 (N_1776,In_2796,In_2011);
xor U1777 (N_1777,In_2506,In_1941);
nor U1778 (N_1778,In_494,In_2484);
and U1779 (N_1779,In_335,In_2391);
nor U1780 (N_1780,In_1396,In_436);
nand U1781 (N_1781,In_2825,In_2466);
nand U1782 (N_1782,In_1874,In_2037);
or U1783 (N_1783,In_2057,In_2547);
and U1784 (N_1784,In_2679,In_577);
xnor U1785 (N_1785,In_530,In_855);
nand U1786 (N_1786,In_1229,In_437);
nand U1787 (N_1787,In_15,In_2648);
nor U1788 (N_1788,In_1621,In_2949);
nand U1789 (N_1789,In_1822,In_1734);
nand U1790 (N_1790,In_1226,In_1713);
and U1791 (N_1791,In_1685,In_748);
and U1792 (N_1792,In_1909,In_2062);
nand U1793 (N_1793,In_2532,In_1153);
or U1794 (N_1794,In_1157,In_2844);
nor U1795 (N_1795,In_2573,In_849);
nor U1796 (N_1796,In_2809,In_2377);
nand U1797 (N_1797,In_672,In_1927);
and U1798 (N_1798,In_1043,In_253);
or U1799 (N_1799,In_2198,In_2795);
nor U1800 (N_1800,In_1343,In_1278);
and U1801 (N_1801,In_192,In_2407);
nor U1802 (N_1802,In_43,In_2219);
nand U1803 (N_1803,In_1292,In_2445);
or U1804 (N_1804,In_1162,In_2520);
and U1805 (N_1805,In_116,In_2128);
and U1806 (N_1806,In_2782,In_1986);
nand U1807 (N_1807,In_1044,In_1579);
nor U1808 (N_1808,In_360,In_2349);
xnor U1809 (N_1809,In_823,In_1216);
xnor U1810 (N_1810,In_2545,In_972);
and U1811 (N_1811,In_1260,In_1137);
xnor U1812 (N_1812,In_2383,In_609);
or U1813 (N_1813,In_2694,In_1706);
or U1814 (N_1814,In_2523,In_2644);
nand U1815 (N_1815,In_1851,In_1250);
or U1816 (N_1816,In_644,In_1852);
xnor U1817 (N_1817,In_292,In_1602);
and U1818 (N_1818,In_1777,In_2636);
or U1819 (N_1819,In_1138,In_2034);
or U1820 (N_1820,In_1788,In_596);
and U1821 (N_1821,In_1641,In_1260);
xnor U1822 (N_1822,In_484,In_1231);
xor U1823 (N_1823,In_357,In_1622);
nor U1824 (N_1824,In_1767,In_2586);
nand U1825 (N_1825,In_1811,In_2670);
or U1826 (N_1826,In_2915,In_343);
xor U1827 (N_1827,In_2770,In_1008);
nor U1828 (N_1828,In_1365,In_2464);
nand U1829 (N_1829,In_849,In_1968);
nand U1830 (N_1830,In_1352,In_136);
nand U1831 (N_1831,In_2614,In_1321);
and U1832 (N_1832,In_471,In_1893);
xnor U1833 (N_1833,In_1659,In_2417);
and U1834 (N_1834,In_275,In_1567);
or U1835 (N_1835,In_540,In_1263);
and U1836 (N_1836,In_2031,In_1874);
xnor U1837 (N_1837,In_5,In_2305);
and U1838 (N_1838,In_2955,In_1793);
or U1839 (N_1839,In_1465,In_1997);
nor U1840 (N_1840,In_1565,In_1112);
xor U1841 (N_1841,In_485,In_776);
xor U1842 (N_1842,In_2342,In_208);
xor U1843 (N_1843,In_1753,In_661);
nand U1844 (N_1844,In_1289,In_544);
and U1845 (N_1845,In_2824,In_398);
nor U1846 (N_1846,In_1344,In_2583);
or U1847 (N_1847,In_87,In_1321);
nand U1848 (N_1848,In_1063,In_2259);
nor U1849 (N_1849,In_300,In_1429);
nand U1850 (N_1850,In_2296,In_572);
xnor U1851 (N_1851,In_1050,In_2956);
and U1852 (N_1852,In_1504,In_2625);
and U1853 (N_1853,In_1145,In_2498);
and U1854 (N_1854,In_1104,In_1109);
xor U1855 (N_1855,In_141,In_1755);
xnor U1856 (N_1856,In_361,In_2797);
nand U1857 (N_1857,In_859,In_1339);
or U1858 (N_1858,In_983,In_428);
and U1859 (N_1859,In_1191,In_2023);
nand U1860 (N_1860,In_2101,In_2554);
or U1861 (N_1861,In_1646,In_2889);
and U1862 (N_1862,In_2573,In_730);
xnor U1863 (N_1863,In_2132,In_2041);
or U1864 (N_1864,In_2659,In_1238);
nor U1865 (N_1865,In_2724,In_2290);
xnor U1866 (N_1866,In_1635,In_1916);
nand U1867 (N_1867,In_1621,In_2942);
and U1868 (N_1868,In_2582,In_1685);
or U1869 (N_1869,In_1197,In_731);
or U1870 (N_1870,In_612,In_147);
nand U1871 (N_1871,In_1939,In_2871);
nand U1872 (N_1872,In_2078,In_1560);
and U1873 (N_1873,In_2173,In_419);
nand U1874 (N_1874,In_1980,In_1902);
or U1875 (N_1875,In_1474,In_2238);
xor U1876 (N_1876,In_2885,In_433);
and U1877 (N_1877,In_2404,In_1576);
xnor U1878 (N_1878,In_2269,In_2332);
nand U1879 (N_1879,In_1365,In_2148);
xnor U1880 (N_1880,In_1831,In_2055);
xnor U1881 (N_1881,In_2617,In_317);
nand U1882 (N_1882,In_2388,In_1400);
and U1883 (N_1883,In_874,In_219);
xnor U1884 (N_1884,In_2707,In_681);
and U1885 (N_1885,In_1232,In_1687);
and U1886 (N_1886,In_1932,In_637);
or U1887 (N_1887,In_2337,In_2726);
nand U1888 (N_1888,In_462,In_1158);
xnor U1889 (N_1889,In_1989,In_1912);
or U1890 (N_1890,In_863,In_2670);
nor U1891 (N_1891,In_2519,In_467);
nor U1892 (N_1892,In_1820,In_2605);
nand U1893 (N_1893,In_1866,In_753);
nor U1894 (N_1894,In_2184,In_1376);
nor U1895 (N_1895,In_1613,In_31);
or U1896 (N_1896,In_2119,In_445);
or U1897 (N_1897,In_2182,In_48);
and U1898 (N_1898,In_1745,In_2439);
or U1899 (N_1899,In_2895,In_2406);
nand U1900 (N_1900,In_2436,In_2723);
or U1901 (N_1901,In_1838,In_2931);
or U1902 (N_1902,In_884,In_1432);
nand U1903 (N_1903,In_698,In_1402);
nor U1904 (N_1904,In_563,In_278);
nand U1905 (N_1905,In_555,In_2116);
or U1906 (N_1906,In_1963,In_223);
nor U1907 (N_1907,In_1694,In_1216);
or U1908 (N_1908,In_2258,In_1617);
nor U1909 (N_1909,In_2544,In_2536);
nand U1910 (N_1910,In_2373,In_1513);
xnor U1911 (N_1911,In_1949,In_2206);
nand U1912 (N_1912,In_2109,In_97);
and U1913 (N_1913,In_1033,In_908);
nor U1914 (N_1914,In_645,In_712);
or U1915 (N_1915,In_2486,In_610);
or U1916 (N_1916,In_970,In_1402);
xor U1917 (N_1917,In_2686,In_1288);
or U1918 (N_1918,In_296,In_1898);
nor U1919 (N_1919,In_2397,In_2315);
and U1920 (N_1920,In_1264,In_2714);
and U1921 (N_1921,In_1255,In_333);
xor U1922 (N_1922,In_2636,In_320);
nand U1923 (N_1923,In_47,In_935);
or U1924 (N_1924,In_1488,In_509);
xor U1925 (N_1925,In_2521,In_1651);
nand U1926 (N_1926,In_2445,In_505);
or U1927 (N_1927,In_1747,In_492);
nor U1928 (N_1928,In_2404,In_2746);
xnor U1929 (N_1929,In_948,In_2342);
xor U1930 (N_1930,In_2338,In_1184);
or U1931 (N_1931,In_1604,In_1226);
or U1932 (N_1932,In_303,In_2998);
nor U1933 (N_1933,In_2465,In_1236);
and U1934 (N_1934,In_2926,In_422);
nand U1935 (N_1935,In_514,In_2860);
or U1936 (N_1936,In_72,In_742);
nor U1937 (N_1937,In_475,In_2193);
nor U1938 (N_1938,In_1606,In_938);
nand U1939 (N_1939,In_220,In_1302);
xor U1940 (N_1940,In_2740,In_2030);
or U1941 (N_1941,In_2399,In_1021);
or U1942 (N_1942,In_2742,In_1619);
and U1943 (N_1943,In_2051,In_1686);
xnor U1944 (N_1944,In_1109,In_2917);
xnor U1945 (N_1945,In_275,In_1562);
xor U1946 (N_1946,In_1043,In_2388);
and U1947 (N_1947,In_976,In_9);
nor U1948 (N_1948,In_245,In_2692);
nand U1949 (N_1949,In_218,In_2464);
or U1950 (N_1950,In_1800,In_2613);
and U1951 (N_1951,In_2145,In_1211);
and U1952 (N_1952,In_1202,In_1994);
and U1953 (N_1953,In_1348,In_2093);
or U1954 (N_1954,In_2394,In_1904);
nor U1955 (N_1955,In_2918,In_2364);
xor U1956 (N_1956,In_1520,In_1078);
nand U1957 (N_1957,In_2946,In_2755);
or U1958 (N_1958,In_1665,In_2639);
or U1959 (N_1959,In_641,In_158);
xnor U1960 (N_1960,In_1532,In_2409);
nor U1961 (N_1961,In_2502,In_156);
xnor U1962 (N_1962,In_6,In_1394);
nor U1963 (N_1963,In_1777,In_2045);
xnor U1964 (N_1964,In_1025,In_528);
or U1965 (N_1965,In_557,In_1145);
or U1966 (N_1966,In_2357,In_1398);
nor U1967 (N_1967,In_990,In_2813);
and U1968 (N_1968,In_1699,In_2094);
or U1969 (N_1969,In_522,In_702);
or U1970 (N_1970,In_698,In_913);
and U1971 (N_1971,In_156,In_2765);
or U1972 (N_1972,In_2876,In_2824);
and U1973 (N_1973,In_420,In_2770);
or U1974 (N_1974,In_1654,In_2466);
nand U1975 (N_1975,In_2923,In_2351);
or U1976 (N_1976,In_1467,In_1881);
and U1977 (N_1977,In_462,In_146);
nand U1978 (N_1978,In_419,In_774);
or U1979 (N_1979,In_1859,In_2338);
and U1980 (N_1980,In_346,In_462);
nor U1981 (N_1981,In_1437,In_300);
nor U1982 (N_1982,In_411,In_1258);
nand U1983 (N_1983,In_1079,In_649);
nor U1984 (N_1984,In_1991,In_775);
or U1985 (N_1985,In_2910,In_1083);
xor U1986 (N_1986,In_2950,In_2656);
and U1987 (N_1987,In_1690,In_1103);
or U1988 (N_1988,In_1368,In_898);
xnor U1989 (N_1989,In_2112,In_701);
or U1990 (N_1990,In_88,In_2659);
xnor U1991 (N_1991,In_2300,In_2926);
and U1992 (N_1992,In_494,In_2128);
or U1993 (N_1993,In_696,In_583);
xor U1994 (N_1994,In_372,In_1574);
xor U1995 (N_1995,In_430,In_2024);
nand U1996 (N_1996,In_2924,In_1673);
nor U1997 (N_1997,In_2407,In_709);
or U1998 (N_1998,In_2518,In_1739);
or U1999 (N_1999,In_2408,In_1184);
nor U2000 (N_2000,In_1438,In_1427);
or U2001 (N_2001,In_2378,In_1231);
or U2002 (N_2002,In_2496,In_1902);
and U2003 (N_2003,In_2814,In_1712);
nor U2004 (N_2004,In_762,In_2343);
nor U2005 (N_2005,In_156,In_375);
nand U2006 (N_2006,In_769,In_2060);
or U2007 (N_2007,In_1914,In_1294);
xor U2008 (N_2008,In_2809,In_2430);
and U2009 (N_2009,In_1781,In_1519);
or U2010 (N_2010,In_1712,In_1458);
nor U2011 (N_2011,In_2527,In_2369);
and U2012 (N_2012,In_2226,In_1300);
or U2013 (N_2013,In_210,In_1062);
xor U2014 (N_2014,In_942,In_482);
nand U2015 (N_2015,In_2226,In_1492);
xor U2016 (N_2016,In_1528,In_2867);
nor U2017 (N_2017,In_1778,In_2723);
and U2018 (N_2018,In_1966,In_2768);
and U2019 (N_2019,In_2768,In_2302);
or U2020 (N_2020,In_997,In_1961);
xor U2021 (N_2021,In_1245,In_2911);
and U2022 (N_2022,In_1777,In_654);
and U2023 (N_2023,In_2936,In_731);
and U2024 (N_2024,In_1413,In_2158);
nor U2025 (N_2025,In_2556,In_58);
xnor U2026 (N_2026,In_4,In_1357);
and U2027 (N_2027,In_1473,In_1146);
and U2028 (N_2028,In_1907,In_2429);
xnor U2029 (N_2029,In_1847,In_58);
xnor U2030 (N_2030,In_1512,In_997);
and U2031 (N_2031,In_56,In_2424);
nor U2032 (N_2032,In_349,In_2070);
nand U2033 (N_2033,In_16,In_362);
xor U2034 (N_2034,In_1965,In_1737);
nand U2035 (N_2035,In_2408,In_1323);
or U2036 (N_2036,In_1735,In_1251);
nor U2037 (N_2037,In_11,In_1476);
and U2038 (N_2038,In_43,In_1462);
or U2039 (N_2039,In_253,In_1082);
nand U2040 (N_2040,In_208,In_2876);
and U2041 (N_2041,In_2969,In_1174);
and U2042 (N_2042,In_542,In_1222);
xor U2043 (N_2043,In_524,In_2181);
xor U2044 (N_2044,In_1519,In_1684);
nand U2045 (N_2045,In_1592,In_2555);
and U2046 (N_2046,In_1861,In_2674);
and U2047 (N_2047,In_788,In_605);
nand U2048 (N_2048,In_2262,In_1860);
xnor U2049 (N_2049,In_1594,In_834);
nor U2050 (N_2050,In_1684,In_83);
xor U2051 (N_2051,In_2552,In_1677);
and U2052 (N_2052,In_430,In_663);
nand U2053 (N_2053,In_1846,In_1032);
xor U2054 (N_2054,In_1439,In_1736);
nand U2055 (N_2055,In_1477,In_2791);
nor U2056 (N_2056,In_1426,In_1198);
nand U2057 (N_2057,In_593,In_1703);
xnor U2058 (N_2058,In_2757,In_709);
nand U2059 (N_2059,In_1975,In_19);
nand U2060 (N_2060,In_1249,In_931);
and U2061 (N_2061,In_137,In_2140);
or U2062 (N_2062,In_1098,In_1832);
nand U2063 (N_2063,In_207,In_2413);
nand U2064 (N_2064,In_2994,In_1231);
or U2065 (N_2065,In_395,In_603);
and U2066 (N_2066,In_481,In_2287);
nand U2067 (N_2067,In_2392,In_786);
and U2068 (N_2068,In_1936,In_392);
or U2069 (N_2069,In_2384,In_810);
and U2070 (N_2070,In_2108,In_2309);
xor U2071 (N_2071,In_2494,In_1218);
nand U2072 (N_2072,In_185,In_651);
nand U2073 (N_2073,In_516,In_1308);
and U2074 (N_2074,In_434,In_439);
nand U2075 (N_2075,In_994,In_2331);
xnor U2076 (N_2076,In_75,In_192);
and U2077 (N_2077,In_680,In_268);
xor U2078 (N_2078,In_1087,In_360);
nor U2079 (N_2079,In_989,In_1072);
and U2080 (N_2080,In_2143,In_481);
nand U2081 (N_2081,In_2847,In_1945);
nand U2082 (N_2082,In_1202,In_491);
nand U2083 (N_2083,In_2968,In_1975);
and U2084 (N_2084,In_392,In_1837);
and U2085 (N_2085,In_1059,In_2470);
or U2086 (N_2086,In_552,In_2045);
xnor U2087 (N_2087,In_693,In_2205);
and U2088 (N_2088,In_115,In_95);
or U2089 (N_2089,In_375,In_2760);
and U2090 (N_2090,In_1862,In_1706);
xor U2091 (N_2091,In_2391,In_237);
and U2092 (N_2092,In_2132,In_1765);
and U2093 (N_2093,In_2460,In_2832);
or U2094 (N_2094,In_2082,In_577);
or U2095 (N_2095,In_106,In_6);
nor U2096 (N_2096,In_1170,In_1852);
nor U2097 (N_2097,In_2449,In_2788);
or U2098 (N_2098,In_1816,In_210);
nor U2099 (N_2099,In_1687,In_564);
nand U2100 (N_2100,In_2203,In_997);
or U2101 (N_2101,In_298,In_2904);
nor U2102 (N_2102,In_1452,In_2994);
nor U2103 (N_2103,In_1778,In_2710);
and U2104 (N_2104,In_2994,In_841);
or U2105 (N_2105,In_9,In_782);
or U2106 (N_2106,In_847,In_365);
nor U2107 (N_2107,In_2628,In_552);
nand U2108 (N_2108,In_2941,In_559);
and U2109 (N_2109,In_444,In_341);
and U2110 (N_2110,In_2663,In_2158);
and U2111 (N_2111,In_194,In_1698);
or U2112 (N_2112,In_1453,In_903);
nand U2113 (N_2113,In_1207,In_1475);
xor U2114 (N_2114,In_2938,In_2332);
and U2115 (N_2115,In_625,In_2937);
nand U2116 (N_2116,In_2339,In_2792);
xnor U2117 (N_2117,In_2361,In_1693);
and U2118 (N_2118,In_639,In_2369);
or U2119 (N_2119,In_1510,In_1260);
and U2120 (N_2120,In_2085,In_2258);
or U2121 (N_2121,In_2917,In_2289);
xnor U2122 (N_2122,In_355,In_713);
or U2123 (N_2123,In_1524,In_822);
xor U2124 (N_2124,In_1616,In_345);
nor U2125 (N_2125,In_531,In_2208);
and U2126 (N_2126,In_121,In_2133);
or U2127 (N_2127,In_1307,In_79);
or U2128 (N_2128,In_1165,In_313);
or U2129 (N_2129,In_226,In_1535);
xor U2130 (N_2130,In_2804,In_2098);
or U2131 (N_2131,In_1946,In_952);
nor U2132 (N_2132,In_1898,In_2133);
or U2133 (N_2133,In_984,In_2445);
nand U2134 (N_2134,In_80,In_1786);
or U2135 (N_2135,In_2710,In_1068);
nor U2136 (N_2136,In_2895,In_1957);
nor U2137 (N_2137,In_1968,In_2196);
nand U2138 (N_2138,In_333,In_2700);
and U2139 (N_2139,In_763,In_1891);
and U2140 (N_2140,In_2735,In_1608);
and U2141 (N_2141,In_2837,In_2083);
nor U2142 (N_2142,In_575,In_868);
nor U2143 (N_2143,In_25,In_2407);
nand U2144 (N_2144,In_356,In_2631);
nand U2145 (N_2145,In_218,In_2302);
xnor U2146 (N_2146,In_1063,In_818);
nand U2147 (N_2147,In_1864,In_2404);
xnor U2148 (N_2148,In_2810,In_1660);
xnor U2149 (N_2149,In_2822,In_1586);
xor U2150 (N_2150,In_2058,In_2030);
and U2151 (N_2151,In_2593,In_2857);
xnor U2152 (N_2152,In_845,In_8);
nor U2153 (N_2153,In_869,In_399);
and U2154 (N_2154,In_2442,In_1482);
nor U2155 (N_2155,In_801,In_89);
xnor U2156 (N_2156,In_125,In_28);
and U2157 (N_2157,In_909,In_2879);
nand U2158 (N_2158,In_2239,In_1405);
and U2159 (N_2159,In_1685,In_1895);
and U2160 (N_2160,In_417,In_2013);
and U2161 (N_2161,In_1004,In_444);
nand U2162 (N_2162,In_2810,In_206);
xor U2163 (N_2163,In_1136,In_2986);
xor U2164 (N_2164,In_2988,In_337);
or U2165 (N_2165,In_2327,In_2762);
and U2166 (N_2166,In_1666,In_1137);
or U2167 (N_2167,In_2462,In_2617);
xnor U2168 (N_2168,In_288,In_1682);
or U2169 (N_2169,In_351,In_2362);
nand U2170 (N_2170,In_83,In_29);
xnor U2171 (N_2171,In_1622,In_842);
xnor U2172 (N_2172,In_2618,In_806);
nand U2173 (N_2173,In_489,In_269);
xnor U2174 (N_2174,In_1329,In_1788);
xnor U2175 (N_2175,In_2519,In_2240);
and U2176 (N_2176,In_2529,In_444);
or U2177 (N_2177,In_229,In_2509);
and U2178 (N_2178,In_2129,In_782);
nor U2179 (N_2179,In_2424,In_1863);
nand U2180 (N_2180,In_178,In_1991);
or U2181 (N_2181,In_2345,In_2242);
nand U2182 (N_2182,In_715,In_405);
nand U2183 (N_2183,In_2704,In_1914);
nor U2184 (N_2184,In_1832,In_1143);
or U2185 (N_2185,In_1718,In_569);
xor U2186 (N_2186,In_909,In_453);
nand U2187 (N_2187,In_993,In_825);
xor U2188 (N_2188,In_668,In_1895);
or U2189 (N_2189,In_1691,In_2643);
xor U2190 (N_2190,In_2853,In_820);
or U2191 (N_2191,In_1574,In_2341);
and U2192 (N_2192,In_457,In_2976);
or U2193 (N_2193,In_2862,In_2551);
or U2194 (N_2194,In_2785,In_1863);
nor U2195 (N_2195,In_1796,In_2909);
xnor U2196 (N_2196,In_1188,In_2686);
nand U2197 (N_2197,In_1155,In_1793);
or U2198 (N_2198,In_507,In_1483);
nand U2199 (N_2199,In_1536,In_2263);
or U2200 (N_2200,In_2002,In_1839);
nand U2201 (N_2201,In_1747,In_2459);
nand U2202 (N_2202,In_1498,In_1647);
or U2203 (N_2203,In_1940,In_2192);
nor U2204 (N_2204,In_2040,In_900);
xor U2205 (N_2205,In_1812,In_919);
nor U2206 (N_2206,In_183,In_2467);
nor U2207 (N_2207,In_2181,In_1981);
xnor U2208 (N_2208,In_1867,In_1307);
xnor U2209 (N_2209,In_2869,In_1146);
xnor U2210 (N_2210,In_376,In_1359);
or U2211 (N_2211,In_1789,In_141);
or U2212 (N_2212,In_82,In_984);
or U2213 (N_2213,In_631,In_2899);
nand U2214 (N_2214,In_826,In_1042);
and U2215 (N_2215,In_1690,In_389);
xor U2216 (N_2216,In_1075,In_1583);
and U2217 (N_2217,In_169,In_549);
nor U2218 (N_2218,In_1738,In_2886);
nor U2219 (N_2219,In_400,In_1156);
nor U2220 (N_2220,In_2321,In_33);
nor U2221 (N_2221,In_1403,In_1739);
nand U2222 (N_2222,In_400,In_728);
or U2223 (N_2223,In_128,In_814);
nand U2224 (N_2224,In_2374,In_1818);
nor U2225 (N_2225,In_255,In_1628);
nand U2226 (N_2226,In_345,In_255);
xor U2227 (N_2227,In_2379,In_2475);
or U2228 (N_2228,In_1835,In_1043);
nor U2229 (N_2229,In_1426,In_1992);
nor U2230 (N_2230,In_2668,In_2535);
nand U2231 (N_2231,In_1210,In_457);
and U2232 (N_2232,In_1812,In_2581);
xnor U2233 (N_2233,In_1834,In_1758);
xor U2234 (N_2234,In_868,In_1508);
nor U2235 (N_2235,In_1119,In_491);
nand U2236 (N_2236,In_713,In_2199);
and U2237 (N_2237,In_799,In_2228);
or U2238 (N_2238,In_456,In_2136);
nand U2239 (N_2239,In_2298,In_1513);
xor U2240 (N_2240,In_1011,In_1708);
and U2241 (N_2241,In_2630,In_1134);
or U2242 (N_2242,In_1325,In_474);
nand U2243 (N_2243,In_337,In_1115);
nor U2244 (N_2244,In_904,In_2138);
and U2245 (N_2245,In_1919,In_857);
nand U2246 (N_2246,In_320,In_1204);
or U2247 (N_2247,In_1119,In_2881);
nor U2248 (N_2248,In_2758,In_2325);
nor U2249 (N_2249,In_943,In_576);
and U2250 (N_2250,In_2949,In_1163);
and U2251 (N_2251,In_1465,In_1791);
nand U2252 (N_2252,In_66,In_2159);
nor U2253 (N_2253,In_1018,In_549);
nand U2254 (N_2254,In_2963,In_452);
nor U2255 (N_2255,In_613,In_380);
xor U2256 (N_2256,In_156,In_1039);
nand U2257 (N_2257,In_1779,In_497);
xor U2258 (N_2258,In_1024,In_326);
nor U2259 (N_2259,In_2227,In_2233);
and U2260 (N_2260,In_498,In_2432);
and U2261 (N_2261,In_943,In_1446);
or U2262 (N_2262,In_809,In_2645);
nor U2263 (N_2263,In_654,In_1368);
and U2264 (N_2264,In_2945,In_986);
xor U2265 (N_2265,In_2675,In_2403);
nor U2266 (N_2266,In_415,In_309);
nor U2267 (N_2267,In_2035,In_2262);
nand U2268 (N_2268,In_1382,In_2911);
or U2269 (N_2269,In_437,In_490);
nand U2270 (N_2270,In_2475,In_233);
and U2271 (N_2271,In_1114,In_2136);
xnor U2272 (N_2272,In_780,In_2993);
nand U2273 (N_2273,In_1345,In_1727);
nand U2274 (N_2274,In_2975,In_1136);
nor U2275 (N_2275,In_254,In_1806);
and U2276 (N_2276,In_1227,In_2627);
nor U2277 (N_2277,In_1459,In_1371);
nor U2278 (N_2278,In_2242,In_1553);
nor U2279 (N_2279,In_207,In_247);
nor U2280 (N_2280,In_1288,In_1686);
nand U2281 (N_2281,In_2761,In_2733);
nor U2282 (N_2282,In_1438,In_2379);
nor U2283 (N_2283,In_1265,In_1749);
and U2284 (N_2284,In_190,In_719);
xor U2285 (N_2285,In_2613,In_59);
nand U2286 (N_2286,In_1169,In_2628);
xor U2287 (N_2287,In_2864,In_2541);
or U2288 (N_2288,In_770,In_1758);
nand U2289 (N_2289,In_2066,In_1681);
xnor U2290 (N_2290,In_2386,In_2723);
xor U2291 (N_2291,In_490,In_245);
and U2292 (N_2292,In_456,In_1270);
nand U2293 (N_2293,In_1543,In_2012);
nand U2294 (N_2294,In_1561,In_2165);
xor U2295 (N_2295,In_837,In_1229);
nor U2296 (N_2296,In_2481,In_457);
xor U2297 (N_2297,In_2472,In_248);
nand U2298 (N_2298,In_1017,In_2509);
and U2299 (N_2299,In_1258,In_1779);
or U2300 (N_2300,In_2410,In_1053);
or U2301 (N_2301,In_281,In_1884);
xnor U2302 (N_2302,In_1110,In_988);
xor U2303 (N_2303,In_383,In_853);
or U2304 (N_2304,In_1460,In_596);
nor U2305 (N_2305,In_2563,In_1509);
nor U2306 (N_2306,In_1963,In_591);
xor U2307 (N_2307,In_1578,In_2826);
and U2308 (N_2308,In_1127,In_309);
nand U2309 (N_2309,In_1543,In_2295);
and U2310 (N_2310,In_2715,In_317);
nor U2311 (N_2311,In_456,In_1710);
xor U2312 (N_2312,In_284,In_582);
or U2313 (N_2313,In_2117,In_1069);
nand U2314 (N_2314,In_228,In_80);
nand U2315 (N_2315,In_1495,In_1950);
or U2316 (N_2316,In_975,In_2262);
nor U2317 (N_2317,In_1710,In_2181);
or U2318 (N_2318,In_1933,In_2891);
xnor U2319 (N_2319,In_2505,In_2319);
and U2320 (N_2320,In_41,In_1441);
and U2321 (N_2321,In_58,In_1617);
or U2322 (N_2322,In_670,In_189);
or U2323 (N_2323,In_307,In_1170);
nor U2324 (N_2324,In_431,In_2278);
nand U2325 (N_2325,In_1121,In_2128);
xnor U2326 (N_2326,In_2761,In_746);
or U2327 (N_2327,In_2764,In_1196);
xnor U2328 (N_2328,In_47,In_736);
nand U2329 (N_2329,In_2244,In_1370);
nand U2330 (N_2330,In_2710,In_2008);
xnor U2331 (N_2331,In_156,In_2579);
nor U2332 (N_2332,In_2515,In_2853);
nand U2333 (N_2333,In_2662,In_334);
nand U2334 (N_2334,In_898,In_2750);
nor U2335 (N_2335,In_2448,In_2159);
nand U2336 (N_2336,In_2602,In_465);
xor U2337 (N_2337,In_488,In_2517);
nand U2338 (N_2338,In_300,In_623);
nand U2339 (N_2339,In_2089,In_2248);
or U2340 (N_2340,In_1188,In_98);
nand U2341 (N_2341,In_294,In_1304);
and U2342 (N_2342,In_1366,In_2971);
nand U2343 (N_2343,In_1752,In_2423);
nor U2344 (N_2344,In_2033,In_2164);
xor U2345 (N_2345,In_1056,In_448);
and U2346 (N_2346,In_2042,In_96);
and U2347 (N_2347,In_2370,In_488);
or U2348 (N_2348,In_1074,In_1220);
nand U2349 (N_2349,In_42,In_369);
xor U2350 (N_2350,In_1726,In_2567);
nand U2351 (N_2351,In_1345,In_272);
xor U2352 (N_2352,In_1355,In_2410);
nor U2353 (N_2353,In_2048,In_859);
nor U2354 (N_2354,In_379,In_2697);
xnor U2355 (N_2355,In_1214,In_0);
or U2356 (N_2356,In_1914,In_1217);
nor U2357 (N_2357,In_2965,In_623);
nor U2358 (N_2358,In_11,In_2612);
nor U2359 (N_2359,In_2509,In_2370);
nand U2360 (N_2360,In_820,In_2673);
or U2361 (N_2361,In_614,In_1011);
or U2362 (N_2362,In_2923,In_1928);
xor U2363 (N_2363,In_2425,In_1627);
nand U2364 (N_2364,In_1284,In_1128);
nor U2365 (N_2365,In_1163,In_2259);
or U2366 (N_2366,In_1576,In_80);
nand U2367 (N_2367,In_2127,In_2207);
nor U2368 (N_2368,In_2979,In_2329);
xor U2369 (N_2369,In_140,In_1437);
nand U2370 (N_2370,In_716,In_2807);
and U2371 (N_2371,In_1420,In_2952);
and U2372 (N_2372,In_1733,In_1800);
nor U2373 (N_2373,In_2703,In_543);
nor U2374 (N_2374,In_824,In_2002);
nor U2375 (N_2375,In_77,In_1385);
xnor U2376 (N_2376,In_1167,In_983);
and U2377 (N_2377,In_1785,In_1152);
and U2378 (N_2378,In_978,In_4);
xnor U2379 (N_2379,In_481,In_2800);
nor U2380 (N_2380,In_1222,In_2318);
nor U2381 (N_2381,In_2234,In_2152);
nand U2382 (N_2382,In_1483,In_667);
or U2383 (N_2383,In_1084,In_488);
and U2384 (N_2384,In_186,In_2293);
nor U2385 (N_2385,In_113,In_260);
nand U2386 (N_2386,In_2370,In_1450);
or U2387 (N_2387,In_2304,In_2114);
xor U2388 (N_2388,In_2943,In_2509);
nand U2389 (N_2389,In_601,In_184);
nand U2390 (N_2390,In_2966,In_2049);
nand U2391 (N_2391,In_95,In_23);
nand U2392 (N_2392,In_1601,In_2461);
nand U2393 (N_2393,In_664,In_1995);
nand U2394 (N_2394,In_839,In_2188);
nand U2395 (N_2395,In_2884,In_2460);
nand U2396 (N_2396,In_1963,In_2790);
nand U2397 (N_2397,In_2353,In_2500);
nand U2398 (N_2398,In_955,In_2624);
nand U2399 (N_2399,In_1423,In_635);
xnor U2400 (N_2400,In_2435,In_534);
nand U2401 (N_2401,In_717,In_2970);
xor U2402 (N_2402,In_1001,In_600);
or U2403 (N_2403,In_2181,In_1630);
or U2404 (N_2404,In_2060,In_1813);
or U2405 (N_2405,In_232,In_1040);
xnor U2406 (N_2406,In_2056,In_2846);
or U2407 (N_2407,In_1086,In_1696);
or U2408 (N_2408,In_2957,In_675);
xor U2409 (N_2409,In_1699,In_2241);
nand U2410 (N_2410,In_2072,In_1684);
xor U2411 (N_2411,In_388,In_667);
xnor U2412 (N_2412,In_1993,In_2838);
and U2413 (N_2413,In_1046,In_483);
xor U2414 (N_2414,In_2747,In_2427);
or U2415 (N_2415,In_527,In_1723);
or U2416 (N_2416,In_1301,In_2838);
xor U2417 (N_2417,In_543,In_1326);
or U2418 (N_2418,In_1860,In_1808);
xnor U2419 (N_2419,In_1216,In_2759);
or U2420 (N_2420,In_2748,In_2403);
nor U2421 (N_2421,In_1593,In_1687);
or U2422 (N_2422,In_2805,In_340);
xnor U2423 (N_2423,In_524,In_1487);
and U2424 (N_2424,In_2777,In_1766);
xor U2425 (N_2425,In_2591,In_1489);
nor U2426 (N_2426,In_2032,In_121);
and U2427 (N_2427,In_2892,In_1858);
nand U2428 (N_2428,In_1246,In_2541);
xnor U2429 (N_2429,In_820,In_216);
nor U2430 (N_2430,In_2482,In_269);
nand U2431 (N_2431,In_1196,In_1872);
or U2432 (N_2432,In_548,In_80);
xnor U2433 (N_2433,In_476,In_798);
nor U2434 (N_2434,In_1610,In_1104);
nand U2435 (N_2435,In_1046,In_1930);
or U2436 (N_2436,In_2437,In_187);
and U2437 (N_2437,In_2931,In_2893);
nand U2438 (N_2438,In_172,In_544);
nand U2439 (N_2439,In_1541,In_2983);
xor U2440 (N_2440,In_2237,In_2428);
nand U2441 (N_2441,In_323,In_197);
xnor U2442 (N_2442,In_2447,In_358);
nand U2443 (N_2443,In_584,In_2484);
or U2444 (N_2444,In_958,In_1854);
nand U2445 (N_2445,In_72,In_2135);
nor U2446 (N_2446,In_1065,In_275);
nand U2447 (N_2447,In_1912,In_1455);
nor U2448 (N_2448,In_2896,In_79);
or U2449 (N_2449,In_1234,In_2577);
and U2450 (N_2450,In_1008,In_1161);
xnor U2451 (N_2451,In_133,In_1321);
nor U2452 (N_2452,In_2430,In_1556);
or U2453 (N_2453,In_2061,In_2955);
nor U2454 (N_2454,In_249,In_1261);
nor U2455 (N_2455,In_1119,In_2208);
xnor U2456 (N_2456,In_24,In_1250);
or U2457 (N_2457,In_560,In_112);
and U2458 (N_2458,In_876,In_421);
and U2459 (N_2459,In_1986,In_1949);
xor U2460 (N_2460,In_1478,In_223);
or U2461 (N_2461,In_627,In_2374);
nor U2462 (N_2462,In_2492,In_497);
nand U2463 (N_2463,In_2841,In_545);
and U2464 (N_2464,In_2804,In_2111);
nor U2465 (N_2465,In_2338,In_1628);
nor U2466 (N_2466,In_1755,In_2387);
and U2467 (N_2467,In_441,In_1898);
or U2468 (N_2468,In_2617,In_114);
and U2469 (N_2469,In_1815,In_2287);
and U2470 (N_2470,In_2736,In_2236);
and U2471 (N_2471,In_1013,In_1615);
xor U2472 (N_2472,In_458,In_2743);
nand U2473 (N_2473,In_2695,In_1237);
nor U2474 (N_2474,In_2431,In_1735);
nand U2475 (N_2475,In_1018,In_2785);
xor U2476 (N_2476,In_195,In_1225);
nand U2477 (N_2477,In_1271,In_1703);
nand U2478 (N_2478,In_2488,In_2004);
xor U2479 (N_2479,In_139,In_1256);
or U2480 (N_2480,In_2797,In_2263);
xnor U2481 (N_2481,In_2558,In_1392);
nor U2482 (N_2482,In_2234,In_2400);
or U2483 (N_2483,In_1623,In_479);
nand U2484 (N_2484,In_2199,In_172);
xor U2485 (N_2485,In_932,In_601);
nor U2486 (N_2486,In_603,In_2229);
nand U2487 (N_2487,In_833,In_2839);
nand U2488 (N_2488,In_852,In_666);
and U2489 (N_2489,In_475,In_239);
xor U2490 (N_2490,In_1229,In_178);
xnor U2491 (N_2491,In_2837,In_2705);
xnor U2492 (N_2492,In_953,In_918);
or U2493 (N_2493,In_2470,In_2617);
nor U2494 (N_2494,In_477,In_61);
and U2495 (N_2495,In_962,In_2586);
and U2496 (N_2496,In_2228,In_699);
or U2497 (N_2497,In_1412,In_2948);
xor U2498 (N_2498,In_591,In_1802);
and U2499 (N_2499,In_28,In_2274);
xor U2500 (N_2500,In_2863,In_2708);
or U2501 (N_2501,In_1417,In_1443);
nor U2502 (N_2502,In_12,In_2704);
nor U2503 (N_2503,In_791,In_1470);
nor U2504 (N_2504,In_473,In_2262);
xor U2505 (N_2505,In_1009,In_911);
nand U2506 (N_2506,In_1949,In_1348);
nand U2507 (N_2507,In_677,In_855);
xnor U2508 (N_2508,In_1025,In_2960);
nand U2509 (N_2509,In_175,In_2230);
and U2510 (N_2510,In_1997,In_238);
and U2511 (N_2511,In_1984,In_868);
xor U2512 (N_2512,In_45,In_296);
xnor U2513 (N_2513,In_2185,In_593);
or U2514 (N_2514,In_1783,In_2569);
nor U2515 (N_2515,In_1556,In_739);
nor U2516 (N_2516,In_1599,In_2770);
xor U2517 (N_2517,In_575,In_900);
or U2518 (N_2518,In_2197,In_1620);
nand U2519 (N_2519,In_1846,In_2169);
or U2520 (N_2520,In_2325,In_2692);
nor U2521 (N_2521,In_1467,In_968);
xor U2522 (N_2522,In_2947,In_2901);
or U2523 (N_2523,In_1293,In_1556);
and U2524 (N_2524,In_1340,In_2667);
or U2525 (N_2525,In_1169,In_949);
and U2526 (N_2526,In_2646,In_2689);
nor U2527 (N_2527,In_2687,In_332);
and U2528 (N_2528,In_2439,In_1143);
nor U2529 (N_2529,In_13,In_2949);
nor U2530 (N_2530,In_2322,In_2450);
and U2531 (N_2531,In_1807,In_2903);
and U2532 (N_2532,In_990,In_1111);
nor U2533 (N_2533,In_728,In_1395);
xor U2534 (N_2534,In_2270,In_2506);
nor U2535 (N_2535,In_2260,In_1729);
xnor U2536 (N_2536,In_1561,In_683);
and U2537 (N_2537,In_2599,In_959);
or U2538 (N_2538,In_838,In_2338);
and U2539 (N_2539,In_2910,In_2525);
and U2540 (N_2540,In_2282,In_770);
and U2541 (N_2541,In_1978,In_2272);
nor U2542 (N_2542,In_2914,In_2101);
nand U2543 (N_2543,In_2836,In_2821);
and U2544 (N_2544,In_710,In_1426);
nor U2545 (N_2545,In_2772,In_2609);
nand U2546 (N_2546,In_592,In_2166);
nor U2547 (N_2547,In_117,In_537);
xnor U2548 (N_2548,In_753,In_1881);
and U2549 (N_2549,In_2382,In_2360);
and U2550 (N_2550,In_2587,In_333);
nor U2551 (N_2551,In_848,In_933);
and U2552 (N_2552,In_1883,In_2056);
and U2553 (N_2553,In_141,In_624);
and U2554 (N_2554,In_1354,In_20);
nand U2555 (N_2555,In_2475,In_2397);
xor U2556 (N_2556,In_461,In_1531);
and U2557 (N_2557,In_1914,In_295);
xor U2558 (N_2558,In_1168,In_291);
xor U2559 (N_2559,In_1619,In_2502);
and U2560 (N_2560,In_713,In_1427);
nand U2561 (N_2561,In_2089,In_2324);
and U2562 (N_2562,In_2591,In_2545);
or U2563 (N_2563,In_136,In_2172);
or U2564 (N_2564,In_2084,In_2911);
and U2565 (N_2565,In_410,In_1459);
and U2566 (N_2566,In_1855,In_473);
nor U2567 (N_2567,In_1869,In_2493);
or U2568 (N_2568,In_1715,In_27);
xnor U2569 (N_2569,In_177,In_883);
nand U2570 (N_2570,In_824,In_979);
and U2571 (N_2571,In_1966,In_171);
nand U2572 (N_2572,In_2478,In_2043);
xnor U2573 (N_2573,In_2458,In_1948);
nand U2574 (N_2574,In_1958,In_37);
and U2575 (N_2575,In_542,In_697);
or U2576 (N_2576,In_1203,In_1170);
nand U2577 (N_2577,In_2616,In_2199);
nor U2578 (N_2578,In_2083,In_896);
xnor U2579 (N_2579,In_1827,In_1444);
nand U2580 (N_2580,In_1249,In_2996);
or U2581 (N_2581,In_560,In_952);
nor U2582 (N_2582,In_767,In_1148);
and U2583 (N_2583,In_951,In_344);
xnor U2584 (N_2584,In_795,In_0);
xor U2585 (N_2585,In_1466,In_2298);
or U2586 (N_2586,In_1485,In_2194);
and U2587 (N_2587,In_2943,In_2854);
xnor U2588 (N_2588,In_2049,In_604);
and U2589 (N_2589,In_871,In_2778);
and U2590 (N_2590,In_2020,In_14);
or U2591 (N_2591,In_621,In_2554);
or U2592 (N_2592,In_1911,In_1043);
xor U2593 (N_2593,In_208,In_1631);
nor U2594 (N_2594,In_2967,In_2525);
nor U2595 (N_2595,In_1249,In_1658);
nand U2596 (N_2596,In_315,In_2656);
and U2597 (N_2597,In_1778,In_1097);
nor U2598 (N_2598,In_1331,In_2471);
xor U2599 (N_2599,In_1471,In_220);
nand U2600 (N_2600,In_1330,In_879);
or U2601 (N_2601,In_2314,In_1224);
xnor U2602 (N_2602,In_236,In_617);
or U2603 (N_2603,In_2449,In_2463);
nand U2604 (N_2604,In_2149,In_2182);
and U2605 (N_2605,In_390,In_591);
and U2606 (N_2606,In_2648,In_137);
nor U2607 (N_2607,In_1870,In_453);
nand U2608 (N_2608,In_583,In_999);
and U2609 (N_2609,In_1613,In_497);
xor U2610 (N_2610,In_1050,In_1815);
nand U2611 (N_2611,In_1048,In_2027);
and U2612 (N_2612,In_1265,In_352);
nor U2613 (N_2613,In_166,In_1701);
xnor U2614 (N_2614,In_2299,In_1926);
xnor U2615 (N_2615,In_198,In_74);
and U2616 (N_2616,In_259,In_2446);
nor U2617 (N_2617,In_1337,In_511);
or U2618 (N_2618,In_201,In_1463);
nor U2619 (N_2619,In_1206,In_1772);
or U2620 (N_2620,In_997,In_699);
and U2621 (N_2621,In_1599,In_1632);
or U2622 (N_2622,In_718,In_679);
or U2623 (N_2623,In_1389,In_2388);
or U2624 (N_2624,In_1003,In_2274);
and U2625 (N_2625,In_1420,In_1034);
xnor U2626 (N_2626,In_1629,In_2930);
nand U2627 (N_2627,In_1400,In_2315);
nor U2628 (N_2628,In_2944,In_1932);
and U2629 (N_2629,In_2105,In_787);
nor U2630 (N_2630,In_386,In_1477);
xnor U2631 (N_2631,In_1402,In_2067);
nor U2632 (N_2632,In_1583,In_1040);
nand U2633 (N_2633,In_1827,In_2129);
xor U2634 (N_2634,In_2083,In_827);
nand U2635 (N_2635,In_1815,In_1556);
xor U2636 (N_2636,In_2470,In_1431);
nand U2637 (N_2637,In_2878,In_20);
xor U2638 (N_2638,In_88,In_1251);
nor U2639 (N_2639,In_2840,In_2013);
or U2640 (N_2640,In_1330,In_253);
nor U2641 (N_2641,In_2875,In_2021);
and U2642 (N_2642,In_880,In_2521);
nor U2643 (N_2643,In_1065,In_677);
nand U2644 (N_2644,In_1785,In_2991);
nand U2645 (N_2645,In_540,In_1845);
and U2646 (N_2646,In_2106,In_287);
nand U2647 (N_2647,In_449,In_1243);
or U2648 (N_2648,In_2712,In_709);
and U2649 (N_2649,In_2818,In_1721);
nand U2650 (N_2650,In_1364,In_1237);
or U2651 (N_2651,In_1675,In_605);
and U2652 (N_2652,In_1609,In_561);
and U2653 (N_2653,In_1096,In_1337);
xor U2654 (N_2654,In_803,In_873);
or U2655 (N_2655,In_2003,In_2808);
xnor U2656 (N_2656,In_1684,In_46);
or U2657 (N_2657,In_205,In_2227);
or U2658 (N_2658,In_1886,In_1625);
nor U2659 (N_2659,In_1867,In_2719);
xnor U2660 (N_2660,In_113,In_2325);
nand U2661 (N_2661,In_2840,In_2299);
and U2662 (N_2662,In_2348,In_951);
nand U2663 (N_2663,In_2503,In_1049);
xnor U2664 (N_2664,In_1123,In_2166);
xor U2665 (N_2665,In_1084,In_2589);
xor U2666 (N_2666,In_1383,In_1932);
nor U2667 (N_2667,In_78,In_82);
and U2668 (N_2668,In_56,In_857);
xor U2669 (N_2669,In_43,In_2200);
or U2670 (N_2670,In_2307,In_2820);
nand U2671 (N_2671,In_418,In_1537);
or U2672 (N_2672,In_813,In_2495);
and U2673 (N_2673,In_1134,In_763);
xnor U2674 (N_2674,In_1814,In_2206);
nor U2675 (N_2675,In_1629,In_87);
nor U2676 (N_2676,In_1905,In_635);
and U2677 (N_2677,In_2111,In_182);
nor U2678 (N_2678,In_1171,In_1756);
nand U2679 (N_2679,In_563,In_1615);
nand U2680 (N_2680,In_660,In_2399);
and U2681 (N_2681,In_7,In_200);
xnor U2682 (N_2682,In_1496,In_2595);
nand U2683 (N_2683,In_1430,In_1311);
xnor U2684 (N_2684,In_543,In_2424);
xor U2685 (N_2685,In_2721,In_1376);
nor U2686 (N_2686,In_2577,In_490);
and U2687 (N_2687,In_455,In_1824);
and U2688 (N_2688,In_1470,In_1104);
nor U2689 (N_2689,In_2656,In_375);
nand U2690 (N_2690,In_1621,In_939);
nand U2691 (N_2691,In_1369,In_1913);
xor U2692 (N_2692,In_1384,In_458);
or U2693 (N_2693,In_1420,In_1919);
and U2694 (N_2694,In_1973,In_1964);
and U2695 (N_2695,In_2706,In_230);
nor U2696 (N_2696,In_2037,In_21);
xor U2697 (N_2697,In_2470,In_907);
xor U2698 (N_2698,In_1099,In_630);
nand U2699 (N_2699,In_2305,In_1437);
and U2700 (N_2700,In_2104,In_2282);
or U2701 (N_2701,In_2411,In_549);
or U2702 (N_2702,In_2687,In_914);
or U2703 (N_2703,In_1958,In_935);
and U2704 (N_2704,In_1684,In_1951);
and U2705 (N_2705,In_656,In_1581);
nand U2706 (N_2706,In_615,In_1410);
or U2707 (N_2707,In_1074,In_1971);
or U2708 (N_2708,In_1447,In_154);
or U2709 (N_2709,In_1630,In_1945);
or U2710 (N_2710,In_2364,In_1254);
xor U2711 (N_2711,In_1358,In_2696);
or U2712 (N_2712,In_81,In_1726);
nor U2713 (N_2713,In_159,In_1761);
xnor U2714 (N_2714,In_2444,In_2557);
or U2715 (N_2715,In_2450,In_1643);
and U2716 (N_2716,In_2220,In_378);
xnor U2717 (N_2717,In_2335,In_556);
nand U2718 (N_2718,In_2834,In_2755);
and U2719 (N_2719,In_2717,In_549);
or U2720 (N_2720,In_1543,In_574);
nand U2721 (N_2721,In_2527,In_2351);
and U2722 (N_2722,In_1658,In_896);
and U2723 (N_2723,In_580,In_784);
or U2724 (N_2724,In_111,In_2108);
nor U2725 (N_2725,In_273,In_1073);
nor U2726 (N_2726,In_143,In_2857);
xor U2727 (N_2727,In_2246,In_2865);
and U2728 (N_2728,In_1259,In_2154);
xor U2729 (N_2729,In_2581,In_2941);
or U2730 (N_2730,In_2680,In_2518);
nor U2731 (N_2731,In_2273,In_1170);
and U2732 (N_2732,In_957,In_990);
or U2733 (N_2733,In_419,In_2570);
and U2734 (N_2734,In_2064,In_2668);
nand U2735 (N_2735,In_2613,In_2112);
nand U2736 (N_2736,In_303,In_1396);
or U2737 (N_2737,In_1737,In_2083);
or U2738 (N_2738,In_2121,In_2673);
nor U2739 (N_2739,In_1303,In_1352);
nor U2740 (N_2740,In_2766,In_2889);
nor U2741 (N_2741,In_2277,In_1551);
xor U2742 (N_2742,In_1005,In_2711);
xnor U2743 (N_2743,In_1256,In_1784);
nor U2744 (N_2744,In_929,In_2451);
xnor U2745 (N_2745,In_422,In_1966);
and U2746 (N_2746,In_148,In_1370);
xnor U2747 (N_2747,In_2748,In_42);
nand U2748 (N_2748,In_1874,In_2199);
xnor U2749 (N_2749,In_2215,In_2332);
or U2750 (N_2750,In_2992,In_1566);
and U2751 (N_2751,In_2130,In_2295);
or U2752 (N_2752,In_1439,In_2164);
nand U2753 (N_2753,In_1886,In_2177);
nand U2754 (N_2754,In_1262,In_224);
or U2755 (N_2755,In_2432,In_1520);
and U2756 (N_2756,In_2575,In_1304);
and U2757 (N_2757,In_2995,In_1468);
xnor U2758 (N_2758,In_2790,In_829);
xnor U2759 (N_2759,In_1575,In_2986);
or U2760 (N_2760,In_2603,In_2318);
xnor U2761 (N_2761,In_507,In_2345);
and U2762 (N_2762,In_204,In_1987);
nor U2763 (N_2763,In_745,In_813);
or U2764 (N_2764,In_1306,In_2734);
or U2765 (N_2765,In_114,In_1640);
nor U2766 (N_2766,In_1974,In_1813);
and U2767 (N_2767,In_629,In_146);
xnor U2768 (N_2768,In_252,In_2721);
nor U2769 (N_2769,In_346,In_717);
nor U2770 (N_2770,In_1241,In_1158);
nor U2771 (N_2771,In_753,In_1153);
xnor U2772 (N_2772,In_638,In_41);
or U2773 (N_2773,In_1898,In_1691);
nor U2774 (N_2774,In_1423,In_2130);
xnor U2775 (N_2775,In_696,In_2650);
nand U2776 (N_2776,In_2118,In_2391);
nand U2777 (N_2777,In_1013,In_2810);
nand U2778 (N_2778,In_414,In_2037);
and U2779 (N_2779,In_669,In_713);
or U2780 (N_2780,In_1992,In_834);
nand U2781 (N_2781,In_2609,In_960);
nand U2782 (N_2782,In_83,In_2143);
and U2783 (N_2783,In_1123,In_979);
nand U2784 (N_2784,In_2287,In_1905);
nor U2785 (N_2785,In_789,In_2428);
and U2786 (N_2786,In_1029,In_1109);
nor U2787 (N_2787,In_1034,In_1531);
and U2788 (N_2788,In_1938,In_1376);
nand U2789 (N_2789,In_2502,In_1166);
nand U2790 (N_2790,In_615,In_351);
or U2791 (N_2791,In_683,In_343);
or U2792 (N_2792,In_1740,In_1047);
xor U2793 (N_2793,In_2771,In_494);
and U2794 (N_2794,In_1746,In_1486);
or U2795 (N_2795,In_2527,In_1486);
or U2796 (N_2796,In_1541,In_289);
nand U2797 (N_2797,In_2820,In_393);
xnor U2798 (N_2798,In_2808,In_1795);
nand U2799 (N_2799,In_2093,In_2362);
and U2800 (N_2800,In_601,In_2830);
nor U2801 (N_2801,In_165,In_2560);
xor U2802 (N_2802,In_363,In_2301);
xnor U2803 (N_2803,In_2089,In_2718);
and U2804 (N_2804,In_2564,In_704);
nor U2805 (N_2805,In_2996,In_1274);
and U2806 (N_2806,In_668,In_789);
and U2807 (N_2807,In_2395,In_2209);
xnor U2808 (N_2808,In_2928,In_1658);
and U2809 (N_2809,In_1171,In_1845);
and U2810 (N_2810,In_1217,In_1065);
nor U2811 (N_2811,In_2016,In_2487);
nand U2812 (N_2812,In_318,In_2728);
xor U2813 (N_2813,In_2903,In_1830);
nand U2814 (N_2814,In_1004,In_1583);
or U2815 (N_2815,In_2597,In_63);
and U2816 (N_2816,In_1997,In_1683);
nor U2817 (N_2817,In_2946,In_1188);
nor U2818 (N_2818,In_1872,In_2642);
or U2819 (N_2819,In_2978,In_1105);
nand U2820 (N_2820,In_1575,In_1852);
nor U2821 (N_2821,In_954,In_2131);
xor U2822 (N_2822,In_2771,In_710);
and U2823 (N_2823,In_1448,In_2826);
nor U2824 (N_2824,In_490,In_1859);
or U2825 (N_2825,In_915,In_1394);
nor U2826 (N_2826,In_1838,In_1143);
nor U2827 (N_2827,In_1187,In_12);
or U2828 (N_2828,In_655,In_952);
nand U2829 (N_2829,In_2039,In_2290);
or U2830 (N_2830,In_979,In_759);
or U2831 (N_2831,In_2872,In_2269);
nand U2832 (N_2832,In_981,In_1825);
nor U2833 (N_2833,In_1713,In_1380);
or U2834 (N_2834,In_1462,In_354);
nand U2835 (N_2835,In_2577,In_606);
nand U2836 (N_2836,In_628,In_785);
or U2837 (N_2837,In_2051,In_74);
and U2838 (N_2838,In_2979,In_551);
nand U2839 (N_2839,In_2050,In_1969);
or U2840 (N_2840,In_2723,In_463);
nand U2841 (N_2841,In_2006,In_138);
and U2842 (N_2842,In_915,In_335);
nor U2843 (N_2843,In_2564,In_2235);
and U2844 (N_2844,In_931,In_778);
xor U2845 (N_2845,In_2477,In_2249);
xnor U2846 (N_2846,In_2619,In_1557);
nand U2847 (N_2847,In_2645,In_344);
xor U2848 (N_2848,In_1468,In_2130);
nand U2849 (N_2849,In_483,In_2844);
or U2850 (N_2850,In_1689,In_966);
or U2851 (N_2851,In_1844,In_1305);
and U2852 (N_2852,In_1366,In_2976);
xnor U2853 (N_2853,In_124,In_2143);
nand U2854 (N_2854,In_2366,In_2496);
xor U2855 (N_2855,In_1826,In_26);
and U2856 (N_2856,In_2636,In_2313);
xor U2857 (N_2857,In_2532,In_440);
nand U2858 (N_2858,In_2468,In_2062);
and U2859 (N_2859,In_1964,In_1856);
nor U2860 (N_2860,In_2548,In_1289);
nand U2861 (N_2861,In_579,In_541);
xnor U2862 (N_2862,In_1435,In_1572);
nor U2863 (N_2863,In_642,In_790);
xnor U2864 (N_2864,In_2615,In_1736);
or U2865 (N_2865,In_2008,In_1467);
xor U2866 (N_2866,In_377,In_614);
nand U2867 (N_2867,In_1526,In_354);
nand U2868 (N_2868,In_1851,In_2498);
nand U2869 (N_2869,In_1800,In_180);
and U2870 (N_2870,In_2908,In_601);
or U2871 (N_2871,In_2939,In_2317);
nor U2872 (N_2872,In_2279,In_2736);
and U2873 (N_2873,In_1567,In_2269);
or U2874 (N_2874,In_2572,In_1630);
nor U2875 (N_2875,In_1055,In_685);
nand U2876 (N_2876,In_417,In_832);
nor U2877 (N_2877,In_305,In_1848);
nand U2878 (N_2878,In_2719,In_1253);
nand U2879 (N_2879,In_2523,In_2900);
and U2880 (N_2880,In_546,In_1293);
xnor U2881 (N_2881,In_1666,In_555);
xnor U2882 (N_2882,In_2607,In_1040);
xor U2883 (N_2883,In_2362,In_1881);
or U2884 (N_2884,In_1664,In_1013);
nor U2885 (N_2885,In_1253,In_2928);
nor U2886 (N_2886,In_2420,In_1738);
and U2887 (N_2887,In_600,In_1229);
or U2888 (N_2888,In_2313,In_1013);
or U2889 (N_2889,In_283,In_2025);
and U2890 (N_2890,In_2908,In_1548);
xnor U2891 (N_2891,In_2321,In_2296);
xnor U2892 (N_2892,In_438,In_1895);
or U2893 (N_2893,In_2658,In_2970);
xor U2894 (N_2894,In_1682,In_1401);
nor U2895 (N_2895,In_2621,In_2714);
nor U2896 (N_2896,In_1482,In_867);
or U2897 (N_2897,In_2976,In_1047);
or U2898 (N_2898,In_1499,In_2071);
nand U2899 (N_2899,In_31,In_2412);
xnor U2900 (N_2900,In_2798,In_187);
nor U2901 (N_2901,In_1608,In_1158);
and U2902 (N_2902,In_2376,In_2352);
xnor U2903 (N_2903,In_364,In_2416);
or U2904 (N_2904,In_1355,In_740);
nor U2905 (N_2905,In_1353,In_2086);
nand U2906 (N_2906,In_386,In_1648);
and U2907 (N_2907,In_548,In_353);
xnor U2908 (N_2908,In_1444,In_1479);
nor U2909 (N_2909,In_1738,In_94);
or U2910 (N_2910,In_2233,In_1122);
or U2911 (N_2911,In_1389,In_1817);
nand U2912 (N_2912,In_2188,In_1874);
nor U2913 (N_2913,In_1588,In_1129);
or U2914 (N_2914,In_2391,In_520);
nor U2915 (N_2915,In_2563,In_263);
xnor U2916 (N_2916,In_2962,In_604);
or U2917 (N_2917,In_2775,In_43);
xor U2918 (N_2918,In_659,In_2171);
nand U2919 (N_2919,In_1469,In_1356);
nand U2920 (N_2920,In_44,In_585);
xnor U2921 (N_2921,In_1842,In_2010);
nor U2922 (N_2922,In_2001,In_2009);
xnor U2923 (N_2923,In_243,In_2270);
nor U2924 (N_2924,In_2357,In_8);
nand U2925 (N_2925,In_2945,In_271);
or U2926 (N_2926,In_2160,In_2527);
or U2927 (N_2927,In_2893,In_1787);
and U2928 (N_2928,In_1406,In_1913);
xor U2929 (N_2929,In_2691,In_1720);
nor U2930 (N_2930,In_2414,In_1627);
or U2931 (N_2931,In_1699,In_320);
xnor U2932 (N_2932,In_2970,In_1407);
nor U2933 (N_2933,In_1732,In_1233);
nand U2934 (N_2934,In_65,In_2552);
xnor U2935 (N_2935,In_1212,In_1551);
nor U2936 (N_2936,In_1465,In_1332);
nor U2937 (N_2937,In_2323,In_605);
and U2938 (N_2938,In_586,In_2648);
and U2939 (N_2939,In_1518,In_282);
xor U2940 (N_2940,In_1454,In_1215);
xnor U2941 (N_2941,In_1418,In_1425);
nor U2942 (N_2942,In_878,In_2671);
nand U2943 (N_2943,In_1002,In_1534);
or U2944 (N_2944,In_1786,In_372);
nand U2945 (N_2945,In_1369,In_807);
xor U2946 (N_2946,In_2064,In_1806);
xnor U2947 (N_2947,In_656,In_1019);
or U2948 (N_2948,In_1230,In_2446);
nand U2949 (N_2949,In_1380,In_1341);
nor U2950 (N_2950,In_2898,In_2551);
nor U2951 (N_2951,In_2276,In_673);
nor U2952 (N_2952,In_2028,In_2932);
and U2953 (N_2953,In_1373,In_1091);
or U2954 (N_2954,In_943,In_2349);
or U2955 (N_2955,In_1732,In_1725);
and U2956 (N_2956,In_1696,In_553);
or U2957 (N_2957,In_1638,In_1364);
or U2958 (N_2958,In_1378,In_242);
and U2959 (N_2959,In_2276,In_1137);
and U2960 (N_2960,In_1948,In_428);
xnor U2961 (N_2961,In_2251,In_882);
xor U2962 (N_2962,In_1976,In_2418);
nand U2963 (N_2963,In_1289,In_2784);
nor U2964 (N_2964,In_1768,In_579);
xor U2965 (N_2965,In_573,In_2623);
xor U2966 (N_2966,In_515,In_2258);
nand U2967 (N_2967,In_1990,In_931);
nor U2968 (N_2968,In_462,In_2972);
nor U2969 (N_2969,In_1241,In_2903);
nand U2970 (N_2970,In_1013,In_2699);
xnor U2971 (N_2971,In_1913,In_294);
and U2972 (N_2972,In_1456,In_2713);
nand U2973 (N_2973,In_505,In_1247);
nor U2974 (N_2974,In_2520,In_1539);
nor U2975 (N_2975,In_522,In_1622);
nor U2976 (N_2976,In_1955,In_2848);
nor U2977 (N_2977,In_1341,In_1757);
xnor U2978 (N_2978,In_564,In_1699);
nand U2979 (N_2979,In_2644,In_55);
nor U2980 (N_2980,In_1038,In_434);
and U2981 (N_2981,In_2632,In_305);
nor U2982 (N_2982,In_444,In_928);
and U2983 (N_2983,In_2893,In_2136);
and U2984 (N_2984,In_2288,In_917);
xnor U2985 (N_2985,In_2613,In_2997);
and U2986 (N_2986,In_2845,In_1677);
or U2987 (N_2987,In_2253,In_2593);
or U2988 (N_2988,In_1257,In_2566);
nand U2989 (N_2989,In_279,In_1598);
xnor U2990 (N_2990,In_2127,In_1908);
xor U2991 (N_2991,In_1342,In_2371);
xor U2992 (N_2992,In_1481,In_2985);
nor U2993 (N_2993,In_858,In_1635);
nand U2994 (N_2994,In_294,In_1436);
and U2995 (N_2995,In_2424,In_2641);
nor U2996 (N_2996,In_2318,In_1502);
nor U2997 (N_2997,In_2571,In_1339);
or U2998 (N_2998,In_562,In_1794);
nand U2999 (N_2999,In_1075,In_2442);
or U3000 (N_3000,N_1653,N_2013);
xor U3001 (N_3001,N_96,N_2584);
and U3002 (N_3002,N_1666,N_2076);
xnor U3003 (N_3003,N_883,N_271);
and U3004 (N_3004,N_371,N_1596);
nor U3005 (N_3005,N_1227,N_2394);
and U3006 (N_3006,N_1965,N_1082);
xor U3007 (N_3007,N_576,N_695);
nor U3008 (N_3008,N_1345,N_2288);
nand U3009 (N_3009,N_2844,N_4);
and U3010 (N_3010,N_1687,N_2964);
xnor U3011 (N_3011,N_355,N_1179);
nor U3012 (N_3012,N_2215,N_599);
and U3013 (N_3013,N_23,N_1769);
xnor U3014 (N_3014,N_1205,N_2905);
xnor U3015 (N_3015,N_2906,N_2669);
and U3016 (N_3016,N_1754,N_927);
or U3017 (N_3017,N_113,N_59);
and U3018 (N_3018,N_437,N_1838);
and U3019 (N_3019,N_656,N_517);
or U3020 (N_3020,N_2274,N_2008);
nor U3021 (N_3021,N_122,N_317);
or U3022 (N_3022,N_2522,N_1820);
nand U3023 (N_3023,N_1988,N_1591);
xor U3024 (N_3024,N_1540,N_1924);
and U3025 (N_3025,N_1490,N_1245);
or U3026 (N_3026,N_1688,N_752);
nor U3027 (N_3027,N_1684,N_444);
and U3028 (N_3028,N_1894,N_2942);
or U3029 (N_3029,N_2953,N_2428);
xor U3030 (N_3030,N_2852,N_2272);
or U3031 (N_3031,N_786,N_2755);
or U3032 (N_3032,N_873,N_877);
xor U3033 (N_3033,N_1468,N_1292);
or U3034 (N_3034,N_1115,N_1506);
nor U3035 (N_3035,N_2992,N_28);
and U3036 (N_3036,N_2351,N_1430);
nand U3037 (N_3037,N_545,N_2015);
xor U3038 (N_3038,N_109,N_703);
xor U3039 (N_3039,N_1221,N_1146);
xnor U3040 (N_3040,N_2338,N_247);
xor U3041 (N_3041,N_209,N_1404);
nand U3042 (N_3042,N_1600,N_1352);
xor U3043 (N_3043,N_2848,N_1746);
nor U3044 (N_3044,N_2149,N_2750);
nor U3045 (N_3045,N_473,N_1332);
nor U3046 (N_3046,N_742,N_2245);
xnor U3047 (N_3047,N_1952,N_1732);
nand U3048 (N_3048,N_567,N_138);
and U3049 (N_3049,N_2668,N_563);
nor U3050 (N_3050,N_1400,N_453);
or U3051 (N_3051,N_376,N_35);
nand U3052 (N_3052,N_2787,N_52);
nand U3053 (N_3053,N_1062,N_2781);
nand U3054 (N_3054,N_2534,N_2330);
xor U3055 (N_3055,N_1503,N_377);
and U3056 (N_3056,N_1381,N_1390);
nor U3057 (N_3057,N_572,N_442);
nand U3058 (N_3058,N_2975,N_140);
nand U3059 (N_3059,N_2449,N_1071);
and U3060 (N_3060,N_2179,N_1234);
or U3061 (N_3061,N_741,N_1192);
xor U3062 (N_3062,N_2052,N_1464);
nor U3063 (N_3063,N_1862,N_1690);
or U3064 (N_3064,N_1996,N_2025);
xnor U3065 (N_3065,N_756,N_1885);
nor U3066 (N_3066,N_2464,N_1198);
nand U3067 (N_3067,N_68,N_2372);
or U3068 (N_3068,N_869,N_2653);
nor U3069 (N_3069,N_2559,N_1589);
and U3070 (N_3070,N_2317,N_174);
xnor U3071 (N_3071,N_2273,N_78);
and U3072 (N_3072,N_1346,N_1941);
nor U3073 (N_3073,N_1518,N_211);
and U3074 (N_3074,N_2281,N_2078);
nor U3075 (N_3075,N_155,N_801);
or U3076 (N_3076,N_1419,N_2329);
xor U3077 (N_3077,N_1881,N_2827);
and U3078 (N_3078,N_2788,N_2171);
or U3079 (N_3079,N_858,N_2609);
xnor U3080 (N_3080,N_2914,N_487);
or U3081 (N_3081,N_1399,N_540);
xnor U3082 (N_3082,N_507,N_85);
and U3083 (N_3083,N_726,N_445);
and U3084 (N_3084,N_2421,N_2366);
or U3085 (N_3085,N_862,N_2821);
and U3086 (N_3086,N_782,N_2563);
xor U3087 (N_3087,N_2734,N_2298);
and U3088 (N_3088,N_933,N_547);
nor U3089 (N_3089,N_2315,N_1195);
nor U3090 (N_3090,N_1701,N_1066);
nor U3091 (N_3091,N_1855,N_880);
and U3092 (N_3092,N_1489,N_1005);
nor U3093 (N_3093,N_58,N_1465);
xor U3094 (N_3094,N_1868,N_1233);
or U3095 (N_3095,N_776,N_2945);
or U3096 (N_3096,N_210,N_956);
or U3097 (N_3097,N_2102,N_2955);
xor U3098 (N_3098,N_522,N_2976);
nor U3099 (N_3099,N_2003,N_1280);
xnor U3100 (N_3100,N_1241,N_535);
and U3101 (N_3101,N_2334,N_2304);
or U3102 (N_3102,N_215,N_2977);
nor U3103 (N_3103,N_711,N_2856);
or U3104 (N_3104,N_1922,N_2451);
xnor U3105 (N_3105,N_678,N_2937);
nor U3106 (N_3106,N_2615,N_470);
nor U3107 (N_3107,N_1532,N_1129);
or U3108 (N_3108,N_233,N_1957);
nor U3109 (N_3109,N_2608,N_974);
xnor U3110 (N_3110,N_2410,N_870);
and U3111 (N_3111,N_2084,N_2482);
xor U3112 (N_3112,N_2349,N_1015);
xor U3113 (N_3113,N_2499,N_937);
nor U3114 (N_3114,N_1019,N_1869);
and U3115 (N_3115,N_1959,N_1189);
nor U3116 (N_3116,N_2770,N_1255);
nor U3117 (N_3117,N_1874,N_1328);
or U3118 (N_3118,N_2308,N_2158);
and U3119 (N_3119,N_721,N_1824);
and U3120 (N_3120,N_1153,N_1942);
or U3121 (N_3121,N_2047,N_1572);
nand U3122 (N_3122,N_2257,N_464);
nor U3123 (N_3123,N_556,N_1707);
nand U3124 (N_3124,N_2752,N_2037);
xor U3125 (N_3125,N_2347,N_1662);
and U3126 (N_3126,N_244,N_1347);
and U3127 (N_3127,N_2181,N_2425);
nand U3128 (N_3128,N_2870,N_700);
and U3129 (N_3129,N_2424,N_1800);
xor U3130 (N_3130,N_2907,N_1508);
nand U3131 (N_3131,N_762,N_1373);
and U3132 (N_3132,N_2884,N_868);
and U3133 (N_3133,N_2353,N_1987);
and U3134 (N_3134,N_1182,N_45);
nor U3135 (N_3135,N_180,N_821);
nand U3136 (N_3136,N_1393,N_2936);
and U3137 (N_3137,N_1331,N_1394);
nand U3138 (N_3138,N_2164,N_2356);
nand U3139 (N_3139,N_914,N_767);
nand U3140 (N_3140,N_354,N_2323);
xor U3141 (N_3141,N_2939,N_2773);
or U3142 (N_3142,N_1867,N_950);
or U3143 (N_3143,N_739,N_2355);
or U3144 (N_3144,N_475,N_236);
or U3145 (N_3145,N_339,N_1871);
or U3146 (N_3146,N_1156,N_37);
and U3147 (N_3147,N_1112,N_532);
nor U3148 (N_3148,N_2618,N_98);
or U3149 (N_3149,N_2407,N_2784);
nor U3150 (N_3150,N_1674,N_1479);
nand U3151 (N_3151,N_299,N_154);
or U3152 (N_3152,N_986,N_2243);
nand U3153 (N_3153,N_706,N_282);
or U3154 (N_3154,N_1724,N_1206);
xnor U3155 (N_3155,N_2420,N_2761);
or U3156 (N_3156,N_1717,N_2115);
and U3157 (N_3157,N_1744,N_1416);
nor U3158 (N_3158,N_2834,N_2999);
and U3159 (N_3159,N_2006,N_190);
and U3160 (N_3160,N_2389,N_743);
or U3161 (N_3161,N_2333,N_2081);
or U3162 (N_3162,N_2523,N_130);
xor U3163 (N_3163,N_2064,N_2721);
nor U3164 (N_3164,N_660,N_2322);
and U3165 (N_3165,N_2599,N_1178);
and U3166 (N_3166,N_2796,N_1314);
nand U3167 (N_3167,N_474,N_2292);
or U3168 (N_3168,N_922,N_2111);
and U3169 (N_3169,N_2690,N_963);
nor U3170 (N_3170,N_1938,N_1055);
nand U3171 (N_3171,N_395,N_1607);
nand U3172 (N_3172,N_1649,N_367);
and U3173 (N_3173,N_1384,N_1533);
nor U3174 (N_3174,N_1185,N_2726);
nand U3175 (N_3175,N_2984,N_88);
nand U3176 (N_3176,N_2045,N_2851);
xor U3177 (N_3177,N_2344,N_2483);
or U3178 (N_3178,N_1415,N_1782);
xnor U3179 (N_3179,N_2792,N_358);
or U3180 (N_3180,N_2732,N_2168);
nor U3181 (N_3181,N_512,N_398);
nor U3182 (N_3182,N_1307,N_917);
nor U3183 (N_3183,N_796,N_2136);
nor U3184 (N_3184,N_2675,N_1748);
nand U3185 (N_3185,N_218,N_1843);
nand U3186 (N_3186,N_1720,N_2004);
and U3187 (N_3187,N_1380,N_646);
nand U3188 (N_3188,N_2199,N_527);
or U3189 (N_3189,N_222,N_620);
nor U3190 (N_3190,N_2027,N_2881);
nand U3191 (N_3191,N_882,N_1710);
nand U3192 (N_3192,N_1558,N_1485);
nand U3193 (N_3193,N_709,N_2766);
nand U3194 (N_3194,N_593,N_39);
and U3195 (N_3195,N_369,N_1372);
xnor U3196 (N_3196,N_697,N_1186);
or U3197 (N_3197,N_1794,N_318);
and U3198 (N_3198,N_1694,N_2627);
xnor U3199 (N_3199,N_2812,N_894);
and U3200 (N_3200,N_1910,N_1611);
or U3201 (N_3201,N_1190,N_1437);
xnor U3202 (N_3202,N_1308,N_1539);
and U3203 (N_3203,N_2414,N_2090);
or U3204 (N_3204,N_558,N_2221);
nor U3205 (N_3205,N_2177,N_2515);
or U3206 (N_3206,N_1125,N_202);
nor U3207 (N_3207,N_1382,N_2646);
nand U3208 (N_3208,N_2854,N_670);
and U3209 (N_3209,N_328,N_789);
and U3210 (N_3210,N_510,N_2205);
nand U3211 (N_3211,N_2538,N_2652);
or U3212 (N_3212,N_2838,N_2764);
nor U3213 (N_3213,N_1675,N_2579);
xor U3214 (N_3214,N_1525,N_2929);
or U3215 (N_3215,N_261,N_720);
nor U3216 (N_3216,N_2481,N_1946);
nand U3217 (N_3217,N_2542,N_2550);
or U3218 (N_3218,N_362,N_2613);
nor U3219 (N_3219,N_228,N_2461);
or U3220 (N_3220,N_2035,N_1225);
and U3221 (N_3221,N_2456,N_404);
nor U3222 (N_3222,N_1749,N_2485);
nor U3223 (N_3223,N_1529,N_2662);
nor U3224 (N_3224,N_590,N_167);
and U3225 (N_3225,N_1226,N_177);
xor U3226 (N_3226,N_842,N_115);
xnor U3227 (N_3227,N_1063,N_1278);
or U3228 (N_3228,N_1365,N_1698);
or U3229 (N_3229,N_1925,N_133);
nand U3230 (N_3230,N_570,N_588);
or U3231 (N_3231,N_323,N_609);
nand U3232 (N_3232,N_2904,N_1979);
and U3233 (N_3233,N_1072,N_1822);
nor U3234 (N_3234,N_855,N_2930);
nand U3235 (N_3235,N_1745,N_1472);
xor U3236 (N_3236,N_2216,N_2659);
nand U3237 (N_3237,N_2467,N_2445);
xnor U3238 (N_3238,N_2197,N_1099);
xnor U3239 (N_3239,N_1064,N_1269);
xor U3240 (N_3240,N_1994,N_274);
nor U3241 (N_3241,N_685,N_957);
nor U3242 (N_3242,N_669,N_1279);
or U3243 (N_3243,N_509,N_144);
and U3244 (N_3244,N_1931,N_2283);
nand U3245 (N_3245,N_2144,N_2371);
nand U3246 (N_3246,N_1648,N_1126);
nor U3247 (N_3247,N_2561,N_1374);
xor U3248 (N_3248,N_2070,N_2023);
nor U3249 (N_3249,N_1570,N_16);
or U3250 (N_3250,N_2386,N_1050);
nor U3251 (N_3251,N_2002,N_2140);
and U3252 (N_3252,N_1375,N_2790);
nand U3253 (N_3253,N_790,N_116);
xor U3254 (N_3254,N_2074,N_1833);
or U3255 (N_3255,N_1997,N_1344);
xor U3256 (N_3256,N_1722,N_1715);
xor U3257 (N_3257,N_1035,N_771);
and U3258 (N_3258,N_1008,N_2998);
or U3259 (N_3259,N_492,N_2263);
or U3260 (N_3260,N_3,N_1421);
and U3261 (N_3261,N_674,N_2890);
nor U3262 (N_3262,N_2525,N_73);
xor U3263 (N_3263,N_2236,N_2810);
xor U3264 (N_3264,N_958,N_2778);
xor U3265 (N_3265,N_757,N_1049);
or U3266 (N_3266,N_1719,N_2239);
nor U3267 (N_3267,N_1581,N_1013);
nor U3268 (N_3268,N_2963,N_1170);
xor U3269 (N_3269,N_978,N_1056);
and U3270 (N_3270,N_1811,N_2829);
nor U3271 (N_3271,N_1211,N_723);
nor U3272 (N_3272,N_1557,N_575);
and U3273 (N_3273,N_46,N_2670);
nor U3274 (N_3274,N_627,N_1200);
and U3275 (N_3275,N_1368,N_55);
xnor U3276 (N_3276,N_401,N_2435);
nor U3277 (N_3277,N_1040,N_2367);
or U3278 (N_3278,N_2397,N_2224);
nand U3279 (N_3279,N_1247,N_977);
or U3280 (N_3280,N_2970,N_2629);
nand U3281 (N_3281,N_1645,N_225);
nand U3282 (N_3282,N_2649,N_2402);
xor U3283 (N_3283,N_1670,N_1913);
or U3284 (N_3284,N_1058,N_2949);
or U3285 (N_3285,N_319,N_1095);
and U3286 (N_3286,N_886,N_1093);
nor U3287 (N_3287,N_1875,N_179);
xnor U3288 (N_3288,N_1123,N_467);
nand U3289 (N_3289,N_2733,N_2110);
xor U3290 (N_3290,N_2198,N_2092);
nor U3291 (N_3291,N_1903,N_1426);
and U3292 (N_3292,N_132,N_1886);
or U3293 (N_3293,N_2343,N_2417);
and U3294 (N_3294,N_529,N_2153);
nand U3295 (N_3295,N_1174,N_397);
nand U3296 (N_3296,N_272,N_778);
xor U3297 (N_3297,N_2577,N_2665);
xor U3298 (N_3298,N_146,N_1);
xor U3299 (N_3299,N_524,N_949);
nor U3300 (N_3300,N_2959,N_2843);
nor U3301 (N_3301,N_871,N_2352);
nand U3302 (N_3302,N_1943,N_707);
nand U3303 (N_3303,N_1915,N_861);
and U3304 (N_3304,N_1961,N_1628);
nor U3305 (N_3305,N_1378,N_335);
nand U3306 (N_3306,N_1669,N_2728);
nor U3307 (N_3307,N_1309,N_2840);
xor U3308 (N_3308,N_248,N_1220);
xnor U3309 (N_3309,N_1595,N_53);
nor U3310 (N_3310,N_243,N_324);
nor U3311 (N_3311,N_51,N_1691);
xnor U3312 (N_3312,N_2370,N_128);
xor U3313 (N_3313,N_427,N_1459);
xor U3314 (N_3314,N_1851,N_2921);
and U3315 (N_3315,N_773,N_1517);
xnor U3316 (N_3316,N_826,N_447);
xor U3317 (N_3317,N_994,N_1882);
or U3318 (N_3318,N_2383,N_1147);
and U3319 (N_3319,N_1281,N_1379);
or U3320 (N_3320,N_797,N_2173);
nor U3321 (N_3321,N_476,N_2831);
nand U3322 (N_3322,N_734,N_1795);
nor U3323 (N_3323,N_2235,N_1664);
and U3324 (N_3324,N_141,N_284);
xnor U3325 (N_3325,N_391,N_2249);
nand U3326 (N_3326,N_2434,N_1501);
nor U3327 (N_3327,N_1654,N_1919);
nand U3328 (N_3328,N_1983,N_1944);
nor U3329 (N_3329,N_896,N_135);
nand U3330 (N_3330,N_934,N_1340);
nor U3331 (N_3331,N_1999,N_835);
xnor U3332 (N_3332,N_554,N_14);
or U3333 (N_3333,N_1258,N_231);
nand U3334 (N_3334,N_569,N_701);
nand U3335 (N_3335,N_2896,N_2830);
nand U3336 (N_3336,N_1516,N_975);
or U3337 (N_3337,N_1083,N_70);
and U3338 (N_3338,N_1162,N_263);
nor U3339 (N_3339,N_2968,N_746);
or U3340 (N_3340,N_1028,N_2527);
nand U3341 (N_3341,N_2678,N_900);
nand U3342 (N_3342,N_1409,N_2291);
and U3343 (N_3343,N_2611,N_1656);
and U3344 (N_3344,N_2219,N_2278);
nor U3345 (N_3345,N_208,N_1145);
nand U3346 (N_3346,N_938,N_1176);
and U3347 (N_3347,N_148,N_412);
and U3348 (N_3348,N_1445,N_1405);
nand U3349 (N_3349,N_562,N_1462);
nor U3350 (N_3350,N_2794,N_1844);
nand U3351 (N_3351,N_349,N_961);
and U3352 (N_3352,N_1825,N_2429);
nand U3353 (N_3353,N_1630,N_2302);
or U3354 (N_3354,N_1089,N_531);
xnor U3355 (N_3355,N_2807,N_2922);
or U3356 (N_3356,N_2569,N_2030);
xnor U3357 (N_3357,N_1397,N_1197);
or U3358 (N_3358,N_2493,N_2865);
nor U3359 (N_3359,N_705,N_126);
or U3360 (N_3360,N_1482,N_808);
and U3361 (N_3361,N_980,N_1718);
nor U3362 (N_3362,N_2034,N_1545);
and U3363 (N_3363,N_1061,N_1834);
nand U3364 (N_3364,N_2165,N_1584);
and U3365 (N_3365,N_281,N_1889);
nand U3366 (N_3366,N_2676,N_2188);
xor U3367 (N_3367,N_518,N_170);
nand U3368 (N_3368,N_889,N_2935);
nand U3369 (N_3369,N_253,N_1301);
or U3370 (N_3370,N_1579,N_1427);
xor U3371 (N_3371,N_2672,N_1078);
nor U3372 (N_3372,N_1067,N_2319);
nand U3373 (N_3373,N_2062,N_2242);
nand U3374 (N_3374,N_833,N_993);
nor U3375 (N_3375,N_1821,N_2471);
nand U3376 (N_3376,N_366,N_2699);
or U3377 (N_3377,N_268,N_1367);
or U3378 (N_3378,N_1383,N_719);
nor U3379 (N_3379,N_930,N_410);
nor U3380 (N_3380,N_732,N_288);
nor U3381 (N_3381,N_44,N_1904);
or U3382 (N_3382,N_1859,N_1135);
and U3383 (N_3383,N_1695,N_145);
xor U3384 (N_3384,N_10,N_1683);
nand U3385 (N_3385,N_2822,N_2251);
and U3386 (N_3386,N_970,N_2122);
or U3387 (N_3387,N_2825,N_112);
xor U3388 (N_3388,N_1453,N_1187);
nand U3389 (N_3389,N_2007,N_2450);
xor U3390 (N_3390,N_2539,N_805);
or U3391 (N_3391,N_1325,N_1303);
nor U3392 (N_3392,N_2176,N_1703);
and U3393 (N_3393,N_336,N_1998);
and U3394 (N_3394,N_2422,N_1294);
and U3395 (N_3395,N_615,N_1515);
or U3396 (N_3396,N_1288,N_1127);
or U3397 (N_3397,N_331,N_153);
nand U3398 (N_3398,N_1088,N_64);
and U3399 (N_3399,N_2947,N_72);
nand U3400 (N_3400,N_2507,N_2677);
or U3401 (N_3401,N_2400,N_7);
xor U3402 (N_3402,N_1934,N_2031);
nand U3403 (N_3403,N_2850,N_214);
nor U3404 (N_3404,N_1643,N_361);
xnor U3405 (N_3405,N_1918,N_740);
nand U3406 (N_3406,N_1018,N_650);
nand U3407 (N_3407,N_1512,N_2501);
nand U3408 (N_3408,N_1275,N_1796);
xor U3409 (N_3409,N_812,N_2311);
nor U3410 (N_3410,N_2314,N_766);
and U3411 (N_3411,N_2514,N_389);
nor U3412 (N_3412,N_32,N_887);
or U3413 (N_3413,N_1131,N_1150);
and U3414 (N_3414,N_2411,N_1417);
nand U3415 (N_3415,N_2385,N_1299);
and U3416 (N_3416,N_380,N_751);
and U3417 (N_3417,N_1431,N_2944);
and U3418 (N_3418,N_651,N_240);
nor U3419 (N_3419,N_2404,N_1265);
nor U3420 (N_3420,N_2516,N_183);
and U3421 (N_3421,N_2339,N_2119);
or U3422 (N_3422,N_193,N_731);
nand U3423 (N_3423,N_1561,N_530);
nor U3424 (N_3424,N_1553,N_2193);
xor U3425 (N_3425,N_2737,N_1814);
nand U3426 (N_3426,N_2478,N_2020);
nor U3427 (N_3427,N_1457,N_1693);
nor U3428 (N_3428,N_1068,N_69);
nand U3429 (N_3429,N_579,N_1494);
or U3430 (N_3430,N_1230,N_2786);
and U3431 (N_3431,N_2874,N_1967);
or U3432 (N_3432,N_1460,N_1168);
xor U3433 (N_3433,N_850,N_2991);
nand U3434 (N_3434,N_907,N_879);
nor U3435 (N_3435,N_1551,N_2813);
or U3436 (N_3436,N_2066,N_1202);
or U3437 (N_3437,N_2771,N_1335);
nor U3438 (N_3438,N_2496,N_1714);
and U3439 (N_3439,N_691,N_1429);
nor U3440 (N_3440,N_1790,N_560);
nor U3441 (N_3441,N_951,N_124);
nand U3442 (N_3442,N_503,N_121);
nor U3443 (N_3443,N_1535,N_428);
xnor U3444 (N_3444,N_1026,N_1830);
or U3445 (N_3445,N_1636,N_1070);
nand U3446 (N_3446,N_2697,N_769);
or U3447 (N_3447,N_1239,N_733);
or U3448 (N_3448,N_1141,N_2363);
or U3449 (N_3449,N_526,N_2056);
or U3450 (N_3450,N_1916,N_574);
and U3451 (N_3451,N_2475,N_2987);
and U3452 (N_3452,N_981,N_62);
and U3453 (N_3453,N_2634,N_2806);
nand U3454 (N_3454,N_901,N_2);
and U3455 (N_3455,N_1610,N_2377);
nand U3456 (N_3456,N_1935,N_1092);
and U3457 (N_3457,N_1434,N_2857);
xor U3458 (N_3458,N_105,N_1757);
and U3459 (N_3459,N_626,N_2962);
or U3460 (N_3460,N_224,N_2698);
and U3461 (N_3461,N_834,N_1486);
nor U3462 (N_3462,N_1016,N_2526);
or U3463 (N_3463,N_2580,N_1799);
xnor U3464 (N_3464,N_1679,N_2873);
nor U3465 (N_3465,N_1677,N_2715);
or U3466 (N_3466,N_1312,N_2412);
nand U3467 (N_3467,N_2610,N_340);
xnor U3468 (N_3468,N_1094,N_1742);
and U3469 (N_3469,N_2789,N_2446);
or U3470 (N_3470,N_2934,N_928);
xnor U3471 (N_3471,N_2375,N_1229);
nand U3472 (N_3472,N_2918,N_725);
xnor U3473 (N_3473,N_636,N_2549);
and U3474 (N_3474,N_221,N_2100);
nand U3475 (N_3475,N_160,N_264);
nand U3476 (N_3476,N_1210,N_1734);
and U3477 (N_3477,N_1436,N_1163);
nand U3478 (N_3478,N_119,N_286);
and U3479 (N_3479,N_436,N_189);
or U3480 (N_3480,N_992,N_1342);
nand U3481 (N_3481,N_2952,N_2201);
or U3482 (N_3482,N_1333,N_1428);
or U3483 (N_3483,N_143,N_814);
or U3484 (N_3484,N_2529,N_2206);
or U3485 (N_3485,N_2230,N_1559);
or U3486 (N_3486,N_817,N_551);
and U3487 (N_3487,N_2712,N_2300);
and U3488 (N_3488,N_2913,N_1177);
nand U3489 (N_3489,N_1446,N_2418);
nand U3490 (N_3490,N_277,N_591);
nor U3491 (N_3491,N_1706,N_987);
and U3492 (N_3492,N_1025,N_289);
nand U3493 (N_3493,N_832,N_1930);
xor U3494 (N_3494,N_342,N_2423);
or U3495 (N_3495,N_2701,N_448);
and U3496 (N_3496,N_1392,N_2871);
or U3497 (N_3497,N_848,N_2191);
or U3498 (N_3498,N_2231,N_2705);
nand U3499 (N_3499,N_2082,N_1113);
or U3500 (N_3500,N_1117,N_1102);
or U3501 (N_3501,N_2178,N_548);
or U3502 (N_3502,N_1759,N_671);
nor U3503 (N_3503,N_2863,N_954);
nor U3504 (N_3504,N_1296,N_1556);
nor U3505 (N_3505,N_1010,N_2808);
nor U3506 (N_3506,N_1774,N_2837);
and U3507 (N_3507,N_2880,N_1526);
nor U3508 (N_3508,N_24,N_84);
or U3509 (N_3509,N_1403,N_2917);
and U3510 (N_3510,N_2624,N_2448);
or U3511 (N_3511,N_679,N_1080);
nor U3512 (N_3512,N_2911,N_2924);
or U3513 (N_3513,N_2753,N_2462);
nand U3514 (N_3514,N_2544,N_514);
xor U3515 (N_3515,N_27,N_641);
nand U3516 (N_3516,N_1599,N_537);
nor U3517 (N_3517,N_1914,N_2255);
xnor U3518 (N_3518,N_595,N_2065);
nor U3519 (N_3519,N_71,N_586);
or U3520 (N_3520,N_320,N_13);
xor U3521 (N_3521,N_2954,N_2679);
nand U3522 (N_3522,N_2763,N_2557);
nand U3523 (N_3523,N_1511,N_1339);
xor U3524 (N_3524,N_2551,N_1306);
xor U3525 (N_3525,N_754,N_830);
or U3526 (N_3526,N_1563,N_1065);
xnor U3527 (N_3527,N_117,N_2497);
xnor U3528 (N_3528,N_449,N_2271);
or U3529 (N_3529,N_1074,N_405);
and U3530 (N_3530,N_131,N_2050);
or U3531 (N_3531,N_158,N_884);
and U3532 (N_3532,N_800,N_1022);
xnor U3533 (N_3533,N_1672,N_539);
or U3534 (N_3534,N_1667,N_2537);
nand U3535 (N_3535,N_799,N_654);
nand U3536 (N_3536,N_295,N_1921);
or U3537 (N_3537,N_2900,N_2680);
nand U3538 (N_3538,N_387,N_979);
nand U3539 (N_3539,N_676,N_638);
nor U3540 (N_3540,N_321,N_2958);
or U3541 (N_3541,N_785,N_1369);
or U3542 (N_3542,N_673,N_1945);
and U3543 (N_3543,N_684,N_1736);
and U3544 (N_3544,N_1652,N_953);
nor U3545 (N_3545,N_2700,N_1837);
xnor U3546 (N_3546,N_2696,N_2393);
xnor U3547 (N_3547,N_635,N_450);
or U3548 (N_3548,N_238,N_164);
or U3549 (N_3549,N_1826,N_1962);
nor U3550 (N_3550,N_2583,N_2072);
and U3551 (N_3551,N_2345,N_1632);
or U3552 (N_3552,N_2384,N_203);
nor U3553 (N_3553,N_1173,N_852);
xnor U3554 (N_3554,N_892,N_1574);
or U3555 (N_3555,N_2564,N_1450);
xor U3556 (N_3556,N_2574,N_161);
or U3557 (N_3557,N_2284,N_2495);
or U3558 (N_3558,N_2388,N_1951);
nand U3559 (N_3559,N_440,N_2814);
nand U3560 (N_3560,N_2868,N_519);
xnor U3561 (N_3561,N_2555,N_291);
nand U3562 (N_3562,N_1463,N_229);
xnor U3563 (N_3563,N_129,N_2915);
nor U3564 (N_3564,N_81,N_2337);
xnor U3565 (N_3565,N_2093,N_1893);
nand U3566 (N_3566,N_2277,N_1520);
and U3567 (N_3567,N_1326,N_577);
nand U3568 (N_3568,N_2469,N_2196);
xnor U3569 (N_3569,N_201,N_1947);
xor U3570 (N_3570,N_2836,N_1566);
or U3571 (N_3571,N_2455,N_1029);
or U3572 (N_3572,N_469,N_2452);
and U3573 (N_3573,N_486,N_2683);
nand U3574 (N_3574,N_388,N_2572);
and U3575 (N_3575,N_2431,N_1359);
xor U3576 (N_3576,N_2103,N_184);
nand U3577 (N_3577,N_1054,N_881);
nor U3578 (N_3578,N_1633,N_2256);
and U3579 (N_3579,N_1475,N_1223);
nand U3580 (N_3580,N_1524,N_1700);
xnor U3581 (N_3581,N_1454,N_2130);
nand U3582 (N_3582,N_2264,N_710);
nand U3583 (N_3583,N_2085,N_2685);
or U3584 (N_3584,N_418,N_2993);
xor U3585 (N_3585,N_488,N_468);
or U3586 (N_3586,N_456,N_451);
nor U3587 (N_3587,N_1912,N_847);
or U3588 (N_3588,N_2920,N_947);
and U3589 (N_3589,N_2141,N_1194);
or U3590 (N_3590,N_2474,N_911);
or U3591 (N_3591,N_553,N_2494);
nand U3592 (N_3592,N_2211,N_2973);
nand U3593 (N_3593,N_1100,N_254);
nor U3594 (N_3594,N_1160,N_1548);
xnor U3595 (N_3595,N_666,N_316);
xor U3596 (N_3596,N_1217,N_2741);
or U3597 (N_3597,N_2666,N_2369);
or U3598 (N_3598,N_1097,N_1678);
nor U3599 (N_3599,N_2368,N_2287);
xor U3600 (N_3600,N_1978,N_549);
nand U3601 (N_3601,N_2458,N_199);
or U3602 (N_3602,N_1320,N_1528);
and U3603 (N_3603,N_1180,N_192);
nor U3604 (N_3604,N_2687,N_79);
nor U3605 (N_3605,N_1237,N_1057);
nand U3606 (N_3606,N_1905,N_2518);
nand U3607 (N_3607,N_2419,N_2862);
nand U3608 (N_3608,N_631,N_1854);
nand U3609 (N_3609,N_2160,N_1597);
or U3610 (N_3610,N_936,N_2839);
xnor U3611 (N_3611,N_820,N_1646);
nand U3612 (N_3612,N_1906,N_866);
xor U3613 (N_3613,N_2562,N_2466);
or U3614 (N_3614,N_2727,N_944);
and U3615 (N_3615,N_1723,N_1527);
xnor U3616 (N_3616,N_2596,N_1354);
or U3617 (N_3617,N_1817,N_2350);
nand U3618 (N_3618,N_1252,N_843);
or U3619 (N_3619,N_1316,N_2587);
nand U3620 (N_3620,N_1860,N_2606);
xor U3621 (N_3621,N_1804,N_690);
or U3622 (N_3622,N_909,N_2234);
or U3623 (N_3623,N_2380,N_186);
xnor U3624 (N_3624,N_495,N_1165);
and U3625 (N_3625,N_2899,N_465);
or U3626 (N_3626,N_2878,N_809);
nor U3627 (N_3627,N_1603,N_462);
nand U3628 (N_3628,N_828,N_403);
nor U3629 (N_3629,N_1498,N_1992);
and U3630 (N_3630,N_534,N_1612);
nand U3631 (N_3631,N_2782,N_38);
nand U3632 (N_3632,N_182,N_1231);
nor U3633 (N_3633,N_1364,N_602);
or U3634 (N_3634,N_1973,N_1318);
or U3635 (N_3635,N_2460,N_2486);
or U3636 (N_3636,N_2631,N_2745);
nand U3637 (N_3637,N_2437,N_2946);
nor U3638 (N_3638,N_2248,N_1809);
and U3639 (N_3639,N_1411,N_1139);
nand U3640 (N_3640,N_1295,N_1627);
nand U3641 (N_3641,N_1425,N_89);
or U3642 (N_3642,N_689,N_2869);
nor U3643 (N_3643,N_2465,N_1387);
nand U3644 (N_3644,N_2769,N_2046);
nand U3645 (N_3645,N_1521,N_885);
and U3646 (N_3646,N_82,N_2133);
xor U3647 (N_3647,N_582,N_2817);
or U3648 (N_3648,N_33,N_1897);
nand U3649 (N_3649,N_919,N_1161);
or U3650 (N_3650,N_1075,N_941);
xor U3651 (N_3651,N_1266,N_2882);
nand U3652 (N_3652,N_343,N_1249);
and U3653 (N_3653,N_2378,N_1034);
nor U3654 (N_3654,N_1120,N_618);
and U3655 (N_3655,N_2707,N_1353);
or U3656 (N_3656,N_356,N_370);
xor U3657 (N_3657,N_494,N_2226);
nand U3658 (N_3658,N_1504,N_2265);
or U3659 (N_3659,N_303,N_658);
nor U3660 (N_3660,N_472,N_2432);
nor U3661 (N_3661,N_2735,N_2731);
xnor U3662 (N_3662,N_1792,N_1578);
nand U3663 (N_3663,N_730,N_1264);
nor U3664 (N_3664,N_93,N_640);
and U3665 (N_3665,N_2571,N_255);
and U3666 (N_3666,N_1334,N_653);
nand U3667 (N_3667,N_2042,N_838);
nor U3668 (N_3668,N_443,N_2488);
nor U3669 (N_3669,N_2655,N_2044);
xor U3670 (N_3670,N_2585,N_1027);
nor U3671 (N_3671,N_1772,N_597);
or U3672 (N_3672,N_1219,N_2328);
nand U3673 (N_3673,N_95,N_1692);
nor U3674 (N_3674,N_2797,N_500);
nand U3675 (N_3675,N_1196,N_217);
nand U3676 (N_3676,N_598,N_755);
nand U3677 (N_3677,N_1841,N_2359);
nand U3678 (N_3678,N_1474,N_1761);
nand U3679 (N_3679,N_256,N_2553);
or U3680 (N_3680,N_1461,N_1780);
nor U3681 (N_3681,N_2017,N_2398);
nor U3682 (N_3682,N_1891,N_1571);
or U3683 (N_3683,N_2000,N_1507);
or U3684 (N_3684,N_297,N_2641);
nand U3685 (N_3685,N_991,N_2706);
and U3686 (N_3686,N_2433,N_692);
nand U3687 (N_3687,N_1214,N_998);
or U3688 (N_3688,N_523,N_2391);
xor U3689 (N_3689,N_1267,N_2266);
and U3690 (N_3690,N_1676,N_2858);
or U3691 (N_3691,N_80,N_1592);
xor U3692 (N_3692,N_1467,N_829);
and U3693 (N_3693,N_1023,N_600);
nand U3694 (N_3694,N_2187,N_2099);
nor U3695 (N_3695,N_750,N_648);
nand U3696 (N_3696,N_2162,N_219);
nor U3697 (N_3697,N_283,N_2957);
and U3698 (N_3698,N_2594,N_2280);
xnor U3699 (N_3699,N_1297,N_1414);
nand U3700 (N_3700,N_390,N_2041);
or U3701 (N_3701,N_300,N_249);
and U3702 (N_3702,N_330,N_1873);
nand U3703 (N_3703,N_1585,N_378);
xnor U3704 (N_3704,N_840,N_1084);
nor U3705 (N_3705,N_2578,N_2940);
or U3706 (N_3706,N_1251,N_2026);
nand U3707 (N_3707,N_2213,N_2014);
and U3708 (N_3708,N_619,N_423);
nand U3709 (N_3709,N_2269,N_555);
or U3710 (N_3710,N_929,N_1726);
xnor U3711 (N_3711,N_2990,N_2575);
and U3712 (N_3712,N_1836,N_1502);
and U3713 (N_3713,N_2022,N_2320);
nor U3714 (N_3714,N_623,N_365);
xnor U3715 (N_3715,N_2194,N_194);
xnor U3716 (N_3716,N_1522,N_2673);
nor U3717 (N_3717,N_1560,N_637);
nor U3718 (N_3718,N_557,N_2175);
or U3719 (N_3719,N_2276,N_2576);
nor U3720 (N_3720,N_1104,N_1777);
nor U3721 (N_3721,N_2803,N_313);
and U3722 (N_3722,N_1937,N_1847);
or U3723 (N_3723,N_1111,N_2931);
or U3724 (N_3724,N_996,N_2101);
or U3725 (N_3725,N_774,N_1376);
xnor U3726 (N_3726,N_1567,N_333);
and U3727 (N_3727,N_2143,N_1839);
and U3728 (N_3728,N_1940,N_2744);
nand U3729 (N_3729,N_1614,N_2660);
nor U3730 (N_3730,N_508,N_2325);
or U3731 (N_3731,N_411,N_76);
nor U3732 (N_3732,N_538,N_29);
nand U3733 (N_3733,N_1739,N_106);
nor U3734 (N_3734,N_2919,N_426);
or U3735 (N_3735,N_2075,N_2926);
nor U3736 (N_3736,N_2979,N_1444);
or U3737 (N_3737,N_2573,N_2548);
and U3738 (N_3738,N_2617,N_1552);
nor U3739 (N_3739,N_156,N_874);
nor U3740 (N_3740,N_406,N_760);
xor U3741 (N_3741,N_2285,N_2974);
nor U3742 (N_3742,N_1493,N_1663);
xor U3743 (N_3743,N_897,N_1538);
nand U3744 (N_3744,N_2872,N_2702);
and U3745 (N_3745,N_2923,N_2671);
nand U3746 (N_3746,N_213,N_1408);
nor U3747 (N_3747,N_2011,N_2223);
xor U3748 (N_3748,N_1283,N_1069);
xor U3749 (N_3749,N_1420,N_2894);
xor U3750 (N_3750,N_2746,N_1096);
nand U3751 (N_3751,N_48,N_2588);
nand U3752 (N_3752,N_2307,N_2131);
xnor U3753 (N_3753,N_2477,N_347);
nand U3754 (N_3754,N_196,N_1148);
or U3755 (N_3755,N_1171,N_568);
or U3756 (N_3756,N_1256,N_1157);
xor U3757 (N_3757,N_41,N_149);
xor U3758 (N_3758,N_844,N_1151);
or U3759 (N_3759,N_77,N_1808);
xnor U3760 (N_3760,N_75,N_2633);
and U3761 (N_3761,N_1977,N_311);
or U3762 (N_3762,N_1433,N_1576);
or U3763 (N_3763,N_310,N_2847);
nand U3764 (N_3764,N_816,N_1455);
nand U3765 (N_3765,N_1709,N_1133);
or U3766 (N_3766,N_1601,N_795);
and U3767 (N_3767,N_1499,N_825);
or U3768 (N_3768,N_2531,N_1248);
and U3769 (N_3769,N_2748,N_1588);
nand U3770 (N_3770,N_1658,N_2088);
nor U3771 (N_3771,N_2941,N_611);
xor U3772 (N_3772,N_2282,N_227);
nor U3773 (N_3773,N_694,N_417);
nor U3774 (N_3774,N_841,N_2104);
xnor U3775 (N_3775,N_454,N_2714);
and U3776 (N_3776,N_2552,N_2912);
xnor U3777 (N_3777,N_216,N_2346);
nand U3778 (N_3778,N_2048,N_1435);
and U3779 (N_3779,N_1920,N_1032);
or U3780 (N_3780,N_2492,N_120);
nand U3781 (N_3781,N_1398,N_2186);
and U3782 (N_3782,N_1929,N_2730);
and U3783 (N_3783,N_1810,N_2096);
and U3784 (N_3784,N_1228,N_2306);
xor U3785 (N_3785,N_2740,N_614);
or U3786 (N_3786,N_2182,N_1311);
and U3787 (N_3787,N_1106,N_110);
xor U3788 (N_3788,N_2736,N_804);
or U3789 (N_3789,N_2749,N_1043);
and U3790 (N_3790,N_2484,N_2220);
nand U3791 (N_3791,N_2301,N_2005);
nand U3792 (N_3792,N_2094,N_393);
nor U3793 (N_3793,N_578,N_1167);
and U3794 (N_3794,N_972,N_127);
nor U3795 (N_3795,N_764,N_2793);
or U3796 (N_3796,N_2738,N_1835);
nand U3797 (N_3797,N_2866,N_175);
or U3798 (N_3798,N_1031,N_2049);
nor U3799 (N_3799,N_2106,N_737);
or U3800 (N_3800,N_1755,N_668);
and U3801 (N_3801,N_5,N_686);
nor U3802 (N_3802,N_1424,N_2716);
or U3803 (N_3803,N_1037,N_2043);
nor U3804 (N_3804,N_2879,N_47);
xor U3805 (N_3805,N_783,N_455);
nand U3806 (N_3806,N_1386,N_2846);
xnor U3807 (N_3807,N_2358,N_1355);
and U3808 (N_3808,N_2903,N_157);
and U3809 (N_3809,N_2151,N_463);
nor U3810 (N_3810,N_831,N_276);
and U3811 (N_3811,N_384,N_2117);
or U3812 (N_3812,N_1928,N_1659);
nand U3813 (N_3813,N_2693,N_493);
nor U3814 (N_3814,N_2374,N_942);
xor U3815 (N_3815,N_36,N_735);
xor U3816 (N_3816,N_2951,N_2689);
and U3817 (N_3817,N_1621,N_794);
nor U3818 (N_3818,N_2508,N_513);
or U3819 (N_3819,N_853,N_573);
xnor U3820 (N_3820,N_1606,N_1024);
nor U3821 (N_3821,N_2760,N_307);
nand U3822 (N_3822,N_875,N_770);
xnor U3823 (N_3823,N_374,N_1699);
or U3824 (N_3824,N_2779,N_2172);
and U3825 (N_3825,N_287,N_2113);
or U3826 (N_3826,N_2237,N_1682);
xnor U3827 (N_3827,N_1276,N_2505);
xor U3828 (N_3828,N_925,N_2405);
xnor U3829 (N_3829,N_2528,N_441);
xor U3830 (N_3830,N_103,N_608);
and U3831 (N_3831,N_872,N_1547);
and U3832 (N_3832,N_2628,N_2718);
or U3833 (N_3833,N_2381,N_1626);
or U3834 (N_3834,N_1542,N_2443);
nor U3835 (N_3835,N_479,N_2426);
xnor U3836 (N_3836,N_1356,N_478);
nor U3837 (N_3837,N_1480,N_2876);
nor U3838 (N_3838,N_1319,N_34);
nand U3839 (N_3839,N_432,N_893);
xnor U3840 (N_3840,N_559,N_2600);
nor U3841 (N_3841,N_344,N_2073);
and U3842 (N_3842,N_1286,N_696);
or U3843 (N_3843,N_2415,N_863);
and U3844 (N_3844,N_2218,N_856);
xnor U3845 (N_3845,N_2203,N_2650);
and U3846 (N_3846,N_2063,N_293);
and U3847 (N_3847,N_1879,N_2532);
nand U3848 (N_3848,N_1954,N_943);
or U3849 (N_3849,N_2439,N_1496);
xnor U3850 (N_3850,N_1085,N_101);
or U3851 (N_3851,N_2799,N_198);
and U3852 (N_3852,N_2720,N_2901);
nand U3853 (N_3853,N_1725,N_1315);
nor U3854 (N_3854,N_1216,N_854);
nor U3855 (N_3855,N_250,N_102);
and U3856 (N_3856,N_1491,N_1878);
or U3857 (N_3857,N_505,N_332);
or U3858 (N_3858,N_2902,N_687);
and U3859 (N_3859,N_2240,N_2632);
nor U3860 (N_3860,N_2640,N_839);
and U3861 (N_3861,N_2597,N_1616);
and U3862 (N_3862,N_1238,N_2694);
or U3863 (N_3863,N_1550,N_516);
or U3864 (N_3864,N_702,N_1939);
nor U3865 (N_3865,N_2586,N_565);
and U3866 (N_3866,N_946,N_2399);
xor U3867 (N_3867,N_2126,N_891);
nand U3868 (N_3868,N_2742,N_2071);
or U3869 (N_3869,N_2509,N_429);
xnor U3870 (N_3870,N_246,N_2303);
or U3871 (N_3871,N_2392,N_40);
nand U3872 (N_3872,N_1207,N_1721);
or U3873 (N_3873,N_2459,N_1456);
xor U3874 (N_3874,N_1864,N_1696);
and U3875 (N_3875,N_1006,N_2747);
nor U3876 (N_3876,N_837,N_1604);
xnor U3877 (N_3877,N_2595,N_2791);
or U3878 (N_3878,N_2316,N_1149);
xnor U3879 (N_3879,N_1704,N_2086);
xnor U3880 (N_3880,N_2664,N_2853);
and U3881 (N_3881,N_438,N_168);
nor U3882 (N_3882,N_90,N_1003);
xnor U3883 (N_3883,N_1038,N_948);
xor U3884 (N_3884,N_1812,N_2709);
or U3885 (N_3885,N_2118,N_296);
nand U3886 (N_3886,N_1807,N_1017);
xnor U3887 (N_3887,N_2743,N_1770);
xor U3888 (N_3888,N_724,N_1974);
and U3889 (N_3889,N_107,N_2069);
and U3890 (N_3890,N_1500,N_1208);
xnor U3891 (N_3891,N_2212,N_2318);
and U3892 (N_3892,N_2364,N_56);
nor U3893 (N_3893,N_2010,N_2639);
nand U3894 (N_3894,N_1077,N_501);
xor U3895 (N_3895,N_1244,N_66);
xor U3896 (N_3896,N_1853,N_926);
and U3897 (N_3897,N_1963,N_2137);
nor U3898 (N_3898,N_768,N_1785);
and U3899 (N_3899,N_139,N_338);
or U3900 (N_3900,N_2589,N_1737);
and U3901 (N_3901,N_585,N_269);
xnor U3902 (N_3902,N_1981,N_83);
or U3903 (N_3903,N_1213,N_100);
xor U3904 (N_3904,N_2986,N_2895);
and U3905 (N_3905,N_792,N_680);
nor U3906 (N_3906,N_1260,N_2252);
nand U3907 (N_3907,N_604,N_2061);
and U3908 (N_3908,N_2630,N_2174);
and U3909 (N_3909,N_1788,N_1001);
nor U3910 (N_3910,N_2142,N_904);
nand U3911 (N_3911,N_952,N_2202);
nand U3912 (N_3912,N_1901,N_698);
nand U3913 (N_3913,N_2259,N_2120);
xnor U3914 (N_3914,N_908,N_1124);
nand U3915 (N_3915,N_1098,N_2362);
xor U3916 (N_3916,N_2217,N_2965);
or U3917 (N_3917,N_2348,N_1543);
and U3918 (N_3918,N_2607,N_533);
nand U3919 (N_3919,N_306,N_1647);
xnor U3920 (N_3920,N_1519,N_1052);
xnor U3921 (N_3921,N_966,N_632);
nand U3922 (N_3922,N_114,N_1009);
and U3923 (N_3923,N_2826,N_1740);
nand U3924 (N_3924,N_2512,N_1012);
nor U3925 (N_3925,N_571,N_260);
xnor U3926 (N_3926,N_2332,N_1609);
and U3927 (N_3927,N_504,N_744);
or U3928 (N_3928,N_1608,N_584);
or U3929 (N_3929,N_1787,N_1620);
nand U3930 (N_3930,N_1448,N_902);
nand U3931 (N_3931,N_722,N_1483);
nand U3932 (N_3932,N_2795,N_1175);
nand U3933 (N_3933,N_675,N_2554);
nor U3934 (N_3934,N_1731,N_2511);
or U3935 (N_3935,N_2250,N_915);
nor U3936 (N_3936,N_430,N_1768);
xor U3937 (N_3937,N_1564,N_2091);
nand U3938 (N_3938,N_359,N_1051);
xnor U3939 (N_3939,N_1304,N_806);
or U3940 (N_3940,N_212,N_1402);
and U3941 (N_3941,N_2543,N_2816);
nor U3942 (N_3942,N_999,N_396);
and U3943 (N_3943,N_326,N_1366);
nand U3944 (N_3944,N_207,N_1246);
xnor U3945 (N_3945,N_2390,N_1622);
xnor U3946 (N_3946,N_1349,N_895);
and U3947 (N_3947,N_2184,N_727);
nor U3948 (N_3948,N_667,N_2832);
nor U3949 (N_3949,N_341,N_1716);
nand U3950 (N_3950,N_605,N_30);
nor U3951 (N_3951,N_1909,N_625);
xor U3952 (N_3952,N_2185,N_2570);
nor U3953 (N_3953,N_864,N_262);
nand U3954 (N_3954,N_1293,N_541);
nand U3955 (N_3955,N_1285,N_2711);
nand U3956 (N_3956,N_1469,N_2454);
and U3957 (N_3957,N_2222,N_2932);
xor U3958 (N_3958,N_2757,N_2772);
nor U3959 (N_3959,N_1907,N_2297);
nand U3960 (N_3960,N_1466,N_232);
nand U3961 (N_3961,N_960,N_2336);
and U3962 (N_3962,N_1702,N_589);
and U3963 (N_3963,N_350,N_1007);
and U3964 (N_3964,N_924,N_1128);
or U3965 (N_3965,N_497,N_305);
nand U3966 (N_3966,N_748,N_962);
xor U3967 (N_3967,N_1164,N_1243);
nand U3968 (N_3968,N_1534,N_693);
or U3969 (N_3969,N_181,N_1530);
nor U3970 (N_3970,N_2039,N_1932);
nor U3971 (N_3971,N_2710,N_188);
or U3972 (N_3972,N_2506,N_1634);
and U3973 (N_3973,N_1908,N_2107);
and U3974 (N_3974,N_2603,N_2286);
or U3975 (N_3975,N_983,N_251);
nor U3976 (N_3976,N_496,N_1033);
nand U3977 (N_3977,N_273,N_965);
and U3978 (N_3978,N_2510,N_1831);
or U3979 (N_3979,N_2214,N_2756);
xor U3980 (N_3980,N_2621,N_2408);
xnor U3981 (N_3981,N_1727,N_2886);
or U3982 (N_3982,N_2520,N_1641);
or U3983 (N_3983,N_43,N_1509);
nand U3984 (N_3984,N_1555,N_1407);
nand U3985 (N_3985,N_1756,N_729);
or U3986 (N_3986,N_471,N_381);
nand U3987 (N_3987,N_245,N_1593);
nand U3988 (N_3988,N_1590,N_1137);
nor U3989 (N_3989,N_2883,N_1573);
nand U3990 (N_3990,N_543,N_1371);
nor U3991 (N_3991,N_1711,N_1327);
or U3992 (N_3992,N_1781,N_2897);
xor U3993 (N_3993,N_1650,N_811);
xor U3994 (N_3994,N_2635,N_2725);
nand U3995 (N_3995,N_2800,N_2739);
and U3996 (N_3996,N_1505,N_1212);
xor U3997 (N_3997,N_1422,N_940);
nor U3998 (N_3998,N_2309,N_1199);
and U3999 (N_3999,N_2480,N_2801);
nor U4000 (N_4000,N_2247,N_2145);
nand U4001 (N_4001,N_601,N_434);
or U4002 (N_4002,N_2590,N_1014);
nor U4003 (N_4003,N_1458,N_1865);
and U4004 (N_4004,N_1101,N_681);
nand U4005 (N_4005,N_92,N_1546);
xor U4006 (N_4006,N_1958,N_1655);
nor U4007 (N_4007,N_1823,N_2195);
and U4008 (N_4008,N_566,N_2279);
xor U4009 (N_4009,N_191,N_984);
nand U4010 (N_4010,N_431,N_665);
nand U4011 (N_4011,N_781,N_1410);
nand U4012 (N_4012,N_2125,N_6);
nor U4013 (N_4013,N_2530,N_2233);
and U4014 (N_4014,N_2517,N_1786);
xor U4015 (N_4015,N_309,N_360);
nor U4016 (N_4016,N_1852,N_713);
xnor U4017 (N_4017,N_2877,N_2642);
or U4018 (N_4018,N_50,N_2754);
or U4019 (N_4019,N_1298,N_2908);
xor U4020 (N_4020,N_2667,N_2365);
or U4021 (N_4021,N_502,N_1193);
nand U4022 (N_4022,N_2751,N_2124);
nor U4023 (N_4023,N_1091,N_716);
nor U4024 (N_4024,N_91,N_1619);
xor U4025 (N_4025,N_2152,N_2059);
nor U4026 (N_4026,N_621,N_2463);
xnor U4027 (N_4027,N_712,N_2204);
nand U4028 (N_4028,N_2656,N_1569);
and U4029 (N_4029,N_1750,N_1888);
or U4030 (N_4030,N_1268,N_2207);
nor U4031 (N_4031,N_715,N_1577);
nand U4032 (N_4032,N_2139,N_433);
nor U4033 (N_4033,N_1514,N_1531);
nor U4034 (N_4034,N_661,N_1513);
and U4035 (N_4035,N_1263,N_2382);
xor U4036 (N_4036,N_163,N_2688);
and U4037 (N_4037,N_738,N_616);
nor U4038 (N_4038,N_2864,N_1184);
nand U4039 (N_4039,N_592,N_278);
nor U4040 (N_4040,N_482,N_1090);
nor U4041 (N_4041,N_385,N_312);
xnor U4042 (N_4042,N_137,N_1872);
or U4043 (N_4043,N_2258,N_1324);
nand U4044 (N_4044,N_2427,N_1362);
xor U4045 (N_4045,N_1789,N_1130);
nand U4046 (N_4046,N_2995,N_2658);
or U4047 (N_4047,N_1289,N_1159);
xor U4048 (N_4048,N_2909,N_1218);
nand U4049 (N_4049,N_2893,N_2961);
xor U4050 (N_4050,N_939,N_2604);
or U4051 (N_4051,N_49,N_2147);
xnor U4052 (N_4052,N_521,N_910);
xnor U4053 (N_4053,N_2189,N_1041);
xor U4054 (N_4054,N_408,N_2108);
and U4055 (N_4055,N_633,N_759);
or U4056 (N_4056,N_1562,N_2097);
and U4057 (N_4057,N_2326,N_1793);
or U4058 (N_4058,N_1870,N_2053);
xnor U4059 (N_4059,N_2156,N_2982);
nor U4060 (N_4060,N_818,N_2989);
nand U4061 (N_4061,N_134,N_1586);
xor U4062 (N_4062,N_1819,N_301);
nand U4063 (N_4063,N_1240,N_2444);
or U4064 (N_4064,N_2546,N_1565);
nand U4065 (N_4065,N_2009,N_1441);
and U4066 (N_4066,N_2138,N_1203);
and U4067 (N_4067,N_973,N_2373);
or U4068 (N_4068,N_386,N_2060);
nand U4069 (N_4069,N_325,N_1956);
nand U4070 (N_4070,N_1079,N_1510);
nor U4071 (N_4071,N_9,N_2513);
and U4072 (N_4072,N_8,N_1073);
and U4073 (N_4073,N_346,N_416);
xnor U4074 (N_4074,N_2361,N_1271);
nor U4075 (N_4075,N_1661,N_2246);
nor U4076 (N_4076,N_1766,N_2442);
nand U4077 (N_4077,N_736,N_2708);
and U4078 (N_4078,N_968,N_2605);
nand U4079 (N_4079,N_489,N_1284);
xor U4080 (N_4080,N_2722,N_1848);
nor U4081 (N_4081,N_2933,N_1172);
or U4082 (N_4082,N_2971,N_1413);
xnor U4083 (N_4083,N_1358,N_461);
nor U4084 (N_4084,N_2312,N_399);
and U4085 (N_4085,N_292,N_2704);
nor U4086 (N_4086,N_97,N_1389);
xnor U4087 (N_4087,N_1488,N_2341);
nand U4088 (N_4088,N_1116,N_728);
and U4089 (N_4089,N_1477,N_997);
or U4090 (N_4090,N_2227,N_2956);
nand U4091 (N_4091,N_1582,N_617);
nor U4092 (N_4092,N_275,N_777);
nor U4093 (N_4093,N_2244,N_677);
xnor U4094 (N_4094,N_1618,N_1805);
xor U4095 (N_4095,N_31,N_2593);
nand U4096 (N_4096,N_2114,N_682);
xnor U4097 (N_4097,N_878,N_2032);
xor U4098 (N_4098,N_1036,N_466);
xor U4099 (N_4099,N_1338,N_2805);
xor U4100 (N_4100,N_2910,N_1972);
xor U4101 (N_4101,N_2055,N_104);
xnor U4102 (N_4102,N_1273,N_2335);
xnor U4103 (N_4103,N_2016,N_923);
nor U4104 (N_4104,N_1985,N_2568);
or U4105 (N_4105,N_662,N_2406);
and U4106 (N_4106,N_2253,N_1191);
xor U4107 (N_4107,N_988,N_1322);
nor U4108 (N_4108,N_1138,N_2783);
and U4109 (N_4109,N_1917,N_1274);
and U4110 (N_4110,N_2686,N_298);
nor U4111 (N_4111,N_2476,N_1902);
or U4112 (N_4112,N_2054,N_2980);
nand U4113 (N_4113,N_2489,N_824);
nor U4114 (N_4114,N_1537,N_865);
and U4115 (N_4115,N_610,N_178);
nand U4116 (N_4116,N_1377,N_2268);
and U4117 (N_4117,N_1060,N_290);
xnor U4118 (N_4118,N_375,N_920);
or U4119 (N_4119,N_581,N_913);
nor U4120 (N_4120,N_2150,N_1341);
nand U4121 (N_4121,N_2533,N_813);
xor U4122 (N_4122,N_2167,N_2128);
nor U4123 (N_4123,N_2598,N_1990);
xor U4124 (N_4124,N_2134,N_912);
or U4125 (N_4125,N_1773,N_2681);
and U4126 (N_4126,N_2036,N_1729);
and U4127 (N_4127,N_1984,N_2087);
or U4128 (N_4128,N_1004,N_506);
nor U4129 (N_4129,N_220,N_1081);
xnor U4130 (N_4130,N_2105,N_2860);
and U4131 (N_4131,N_985,N_2238);
or U4132 (N_4132,N_851,N_2468);
xnor U4133 (N_4133,N_802,N_1866);
and U4134 (N_4134,N_123,N_1440);
nand U4135 (N_4135,N_1640,N_2123);
nor U4136 (N_4136,N_235,N_2132);
or U4137 (N_4137,N_1282,N_2487);
nor U4138 (N_4138,N_1613,N_1443);
or U4139 (N_4139,N_775,N_0);
nor U4140 (N_4140,N_2440,N_1497);
xnor U4141 (N_4141,N_1232,N_1863);
nand U4142 (N_4142,N_2379,N_1439);
nor U4143 (N_4143,N_259,N_642);
or U4144 (N_4144,N_903,N_1898);
nand U4145 (N_4145,N_649,N_2647);
and U4146 (N_4146,N_2098,N_780);
nor U4147 (N_4147,N_2295,N_772);
nor U4148 (N_4148,N_798,N_1876);
nor U4149 (N_4149,N_1762,N_931);
and U4150 (N_4150,N_827,N_2560);
and U4151 (N_4151,N_1801,N_373);
or U4152 (N_4152,N_857,N_2842);
nand U4153 (N_4153,N_753,N_1143);
and U4154 (N_4154,N_663,N_1637);
nor U4155 (N_4155,N_647,N_1142);
xor U4156 (N_4156,N_898,N_2209);
nand U4157 (N_4157,N_2190,N_2310);
nand U4158 (N_4158,N_2502,N_606);
and U4159 (N_4159,N_1991,N_860);
nand U4160 (N_4160,N_200,N_2500);
nor U4161 (N_4161,N_2360,N_2582);
nand U4162 (N_4162,N_2759,N_2622);
and U4163 (N_4163,N_383,N_1110);
xnor U4164 (N_4164,N_351,N_2051);
xor U4165 (N_4165,N_643,N_108);
or U4166 (N_4166,N_422,N_1923);
and U4167 (N_4167,N_976,N_2541);
xor U4168 (N_4168,N_446,N_2321);
and U4169 (N_4169,N_2293,N_1948);
or U4170 (N_4170,N_630,N_784);
and U4171 (N_4171,N_205,N_699);
or U4172 (N_4172,N_266,N_257);
nor U4173 (N_4173,N_1583,N_2948);
and U4174 (N_4174,N_279,N_2804);
nor U4175 (N_4175,N_718,N_1625);
or U4176 (N_4176,N_2661,N_945);
or U4177 (N_4177,N_61,N_2503);
or U4178 (N_4178,N_2536,N_1861);
nand U4179 (N_4179,N_515,N_935);
or U4180 (N_4180,N_1829,N_2183);
or U4181 (N_4181,N_1953,N_1955);
and U4182 (N_4182,N_2200,N_204);
and U4183 (N_4183,N_1452,N_239);
nand U4184 (N_4184,N_392,N_688);
or U4185 (N_4185,N_1044,N_2232);
or U4186 (N_4186,N_2663,N_1442);
and U4187 (N_4187,N_499,N_1310);
nand U4188 (N_4188,N_1478,N_1797);
nor U4189 (N_4189,N_2192,N_2969);
xor U4190 (N_4190,N_2849,N_166);
xor U4191 (N_4191,N_1840,N_2835);
xnor U4192 (N_4192,N_793,N_587);
or U4193 (N_4193,N_2447,N_1629);
and U4194 (N_4194,N_2762,N_187);
xor U4195 (N_4195,N_1802,N_1287);
xor U4196 (N_4196,N_2815,N_959);
or U4197 (N_4197,N_226,N_2387);
nor U4198 (N_4198,N_1580,N_2682);
nand U4199 (N_4199,N_1713,N_413);
xnor U4200 (N_4200,N_2889,N_1949);
or U4201 (N_4201,N_1343,N_285);
xnor U4202 (N_4202,N_435,N_2289);
nand U4203 (N_4203,N_1336,N_2340);
or U4204 (N_4204,N_899,N_2438);
nor U4205 (N_4205,N_1936,N_86);
nand U4206 (N_4206,N_2809,N_1842);
nand U4207 (N_4207,N_267,N_372);
xor U4208 (N_4208,N_1783,N_2828);
nand U4209 (N_4209,N_65,N_490);
or U4210 (N_4210,N_890,N_652);
nand U4211 (N_4211,N_2021,N_1481);
or U4212 (N_4212,N_1856,N_525);
or U4213 (N_4213,N_348,N_1733);
or U4214 (N_4214,N_400,N_1771);
xor U4215 (N_4215,N_60,N_480);
or U4216 (N_4216,N_327,N_1887);
or U4217 (N_4217,N_2547,N_1845);
and U4218 (N_4218,N_2758,N_888);
xnor U4219 (N_4219,N_26,N_2519);
xnor U4220 (N_4220,N_2638,N_2820);
xnor U4221 (N_4221,N_176,N_1155);
or U4222 (N_4222,N_1105,N_185);
xor U4223 (N_4223,N_1815,N_1209);
or U4224 (N_4224,N_2713,N_2592);
and U4225 (N_4225,N_1753,N_169);
nand U4226 (N_4226,N_822,N_867);
nand U4227 (N_4227,N_2491,N_1635);
and U4228 (N_4228,N_1030,N_368);
and U4229 (N_4229,N_2994,N_2692);
or U4230 (N_4230,N_1109,N_1451);
xor U4231 (N_4231,N_1406,N_2645);
xnor U4232 (N_4232,N_1665,N_657);
and U4233 (N_4233,N_1685,N_1204);
and U4234 (N_4234,N_2819,N_1351);
nor U4235 (N_4235,N_2170,N_1169);
nand U4236 (N_4236,N_1899,N_314);
and U4237 (N_4237,N_2637,N_1492);
nor U4238 (N_4238,N_520,N_2916);
nor U4239 (N_4239,N_1021,N_2058);
nor U4240 (N_4240,N_1828,N_1272);
and U4241 (N_4241,N_836,N_414);
nand U4242 (N_4242,N_12,N_2785);
xor U4243 (N_4243,N_337,N_481);
nand U4244 (N_4244,N_2210,N_1779);
or U4245 (N_4245,N_2859,N_345);
nor U4246 (N_4246,N_1752,N_2083);
nor U4247 (N_4247,N_2768,N_2129);
or U4248 (N_4248,N_2262,N_2260);
nor U4249 (N_4249,N_2294,N_63);
xnor U4250 (N_4250,N_2636,N_2354);
or U4251 (N_4251,N_2331,N_704);
nand U4252 (N_4252,N_2357,N_2997);
or U4253 (N_4253,N_1388,N_1892);
and U4254 (N_4254,N_1261,N_2029);
and U4255 (N_4255,N_1927,N_1523);
nor U4256 (N_4256,N_1880,N_18);
and U4257 (N_4257,N_906,N_1166);
xor U4258 (N_4258,N_1047,N_1764);
xor U4259 (N_4259,N_111,N_1108);
xor U4260 (N_4260,N_1968,N_67);
nand U4261 (N_4261,N_1767,N_1011);
xor U4262 (N_4262,N_622,N_787);
xnor U4263 (N_4263,N_2887,N_1039);
nand U4264 (N_4264,N_607,N_54);
xor U4265 (N_4265,N_807,N_2684);
and U4266 (N_4266,N_2342,N_1877);
nand U4267 (N_4267,N_409,N_1624);
or U4268 (N_4268,N_2148,N_2601);
nor U4269 (N_4269,N_2403,N_2855);
nor U4270 (N_4270,N_2159,N_803);
nand U4271 (N_4271,N_1152,N_2765);
or U4272 (N_4272,N_2109,N_2135);
and U4273 (N_4273,N_2228,N_1313);
xor U4274 (N_4274,N_1995,N_2012);
nor U4275 (N_4275,N_99,N_315);
nand U4276 (N_4276,N_613,N_304);
nor U4277 (N_4277,N_2535,N_1076);
xnor U4278 (N_4278,N_634,N_1760);
or U4279 (N_4279,N_22,N_1471);
or U4280 (N_4280,N_2943,N_552);
and U4281 (N_4281,N_1846,N_1118);
xor U4282 (N_4282,N_1747,N_1642);
nor U4283 (N_4283,N_995,N_2985);
and U4284 (N_4284,N_1883,N_2717);
and U4285 (N_4285,N_171,N_2401);
or U4286 (N_4286,N_2208,N_1323);
nand U4287 (N_4287,N_1291,N_1236);
or U4288 (N_4288,N_1254,N_491);
xor U4289 (N_4289,N_353,N_2619);
nor U4290 (N_4290,N_1317,N_2166);
nor U4291 (N_4291,N_1623,N_142);
nor U4292 (N_4292,N_714,N_810);
and U4293 (N_4293,N_242,N_1738);
xnor U4294 (N_4294,N_2261,N_2841);
nor U4295 (N_4295,N_2545,N_1449);
xnor U4296 (N_4296,N_425,N_1122);
or U4297 (N_4297,N_2241,N_580);
or U4298 (N_4298,N_1638,N_2413);
xnor U4299 (N_4299,N_1671,N_2967);
nor U4300 (N_4300,N_302,N_1541);
nand U4301 (N_4301,N_415,N_1270);
and U4302 (N_4302,N_672,N_1370);
nor U4303 (N_4303,N_1103,N_969);
and U4304 (N_4304,N_2479,N_1250);
nor U4305 (N_4305,N_876,N_2161);
nand U4306 (N_4306,N_1896,N_1000);
and U4307 (N_4307,N_1201,N_664);
and U4308 (N_4308,N_1784,N_1235);
or U4309 (N_4309,N_1900,N_1858);
nand U4310 (N_4310,N_629,N_1776);
xor U4311 (N_4311,N_1438,N_2774);
or U4312 (N_4312,N_1615,N_1989);
xor U4313 (N_4313,N_758,N_561);
xor U4314 (N_4314,N_2169,N_2565);
nand U4315 (N_4315,N_2441,N_1554);
and U4316 (N_4316,N_823,N_1657);
or U4317 (N_4317,N_1423,N_2648);
nand U4318 (N_4318,N_921,N_206);
xnor U4319 (N_4319,N_1594,N_1969);
nor U4320 (N_4320,N_2498,N_1348);
nor U4321 (N_4321,N_2960,N_2116);
xor U4322 (N_4322,N_280,N_2155);
nand U4323 (N_4323,N_1053,N_329);
and U4324 (N_4324,N_2504,N_1895);
or U4325 (N_4325,N_644,N_1602);
xor U4326 (N_4326,N_2028,N_1253);
nor U4327 (N_4327,N_1827,N_2891);
xnor U4328 (N_4328,N_2472,N_2623);
xor U4329 (N_4329,N_252,N_550);
xor U4330 (N_4330,N_1651,N_1412);
nor U4331 (N_4331,N_2643,N_2867);
nand U4332 (N_4332,N_407,N_394);
xnor U4333 (N_4333,N_624,N_819);
or U4334 (N_4334,N_1188,N_1681);
xnor U4335 (N_4335,N_2067,N_118);
and U4336 (N_4336,N_628,N_2888);
and U4337 (N_4337,N_2521,N_1884);
and U4338 (N_4338,N_459,N_1668);
or U4339 (N_4339,N_2180,N_1396);
and U4340 (N_4340,N_1158,N_1993);
nor U4341 (N_4341,N_2674,N_1473);
or U4342 (N_4342,N_485,N_1791);
or U4343 (N_4343,N_845,N_458);
nor U4344 (N_4344,N_971,N_1960);
or U4345 (N_4345,N_1121,N_1933);
nand U4346 (N_4346,N_1673,N_2591);
nand U4347 (N_4347,N_2409,N_1697);
or U4348 (N_4348,N_2490,N_498);
xnor U4349 (N_4349,N_2127,N_717);
xor U4350 (N_4350,N_2898,N_1970);
nand U4351 (N_4351,N_1385,N_74);
nand U4352 (N_4352,N_1751,N_2154);
and U4353 (N_4353,N_2723,N_544);
or U4354 (N_4354,N_2983,N_2654);
or U4355 (N_4355,N_583,N_2988);
nor U4356 (N_4356,N_150,N_1487);
or U4357 (N_4357,N_2644,N_2457);
or U4358 (N_4358,N_2861,N_195);
xnor U4359 (N_4359,N_237,N_334);
nand U4360 (N_4360,N_603,N_2019);
nand U4361 (N_4361,N_2095,N_2299);
nor U4362 (N_4362,N_1890,N_2540);
nor U4363 (N_4363,N_1470,N_2612);
nor U4364 (N_4364,N_2657,N_17);
and U4365 (N_4365,N_2121,N_439);
or U4366 (N_4366,N_2719,N_2254);
and U4367 (N_4367,N_747,N_2033);
nand U4368 (N_4368,N_159,N_2225);
and U4369 (N_4369,N_223,N_20);
nand U4370 (N_4370,N_1020,N_2950);
nor U4371 (N_4371,N_308,N_2416);
xnor U4372 (N_4372,N_2972,N_967);
nand U4373 (N_4373,N_2885,N_1544);
nand U4374 (N_4374,N_2040,N_21);
xnor U4375 (N_4375,N_173,N_1536);
nor U4376 (N_4376,N_165,N_1966);
and U4377 (N_4377,N_1321,N_1818);
nor U4378 (N_4378,N_2556,N_918);
or U4379 (N_4379,N_294,N_1765);
or U4380 (N_4380,N_2651,N_905);
nand U4381 (N_4381,N_19,N_1705);
and U4382 (N_4382,N_596,N_197);
and U4383 (N_4383,N_2928,N_763);
and U4384 (N_4384,N_1964,N_1549);
nand U4385 (N_4385,N_1257,N_421);
xor U4386 (N_4386,N_2966,N_1728);
or U4387 (N_4387,N_1140,N_2775);
and U4388 (N_4388,N_1803,N_1154);
and U4389 (N_4389,N_2395,N_2729);
and U4390 (N_4390,N_1806,N_1763);
nand U4391 (N_4391,N_2080,N_42);
and U4392 (N_4392,N_788,N_162);
xor U4393 (N_4393,N_528,N_2567);
nor U4394 (N_4394,N_1686,N_2112);
nor U4395 (N_4395,N_357,N_1357);
and U4396 (N_4396,N_234,N_2157);
xor U4397 (N_4397,N_1086,N_1857);
nand U4398 (N_4398,N_379,N_2625);
nand U4399 (N_4399,N_136,N_612);
xnor U4400 (N_4400,N_1735,N_1046);
or U4401 (N_4401,N_1644,N_2777);
or U4402 (N_4402,N_382,N_765);
and U4403 (N_4403,N_1476,N_1290);
nand U4404 (N_4404,N_57,N_2938);
nor U4405 (N_4405,N_542,N_1741);
and U4406 (N_4406,N_1242,N_2824);
and U4407 (N_4407,N_2290,N_2057);
or U4408 (N_4408,N_659,N_1087);
xor U4409 (N_4409,N_1215,N_932);
nor U4410 (N_4410,N_2018,N_2978);
nand U4411 (N_4411,N_1680,N_147);
nor U4412 (N_4412,N_1136,N_2620);
nand U4413 (N_4413,N_2038,N_419);
nand U4414 (N_4414,N_2524,N_270);
or U4415 (N_4415,N_859,N_457);
nand U4416 (N_4416,N_2724,N_352);
or U4417 (N_4417,N_1181,N_2430);
nor U4418 (N_4418,N_2981,N_1743);
xor U4419 (N_4419,N_25,N_1222);
or U4420 (N_4420,N_1798,N_2024);
xnor U4421 (N_4421,N_2703,N_1850);
nor U4422 (N_4422,N_1778,N_964);
or U4423 (N_4423,N_1277,N_2823);
or U4424 (N_4424,N_1495,N_2470);
or U4425 (N_4425,N_1639,N_1708);
xnor U4426 (N_4426,N_989,N_1045);
and U4427 (N_4427,N_1982,N_322);
nand U4428 (N_4428,N_1568,N_1391);
nor U4429 (N_4429,N_483,N_1484);
xor U4430 (N_4430,N_1598,N_1447);
and U4431 (N_4431,N_1107,N_460);
or U4432 (N_4432,N_1361,N_2146);
or U4433 (N_4433,N_2798,N_2436);
xor U4434 (N_4434,N_749,N_420);
xor U4435 (N_4435,N_1119,N_2089);
xnor U4436 (N_4436,N_2892,N_990);
xor U4437 (N_4437,N_846,N_1575);
nor U4438 (N_4438,N_779,N_230);
or U4439 (N_4439,N_2396,N_2270);
nor U4440 (N_4440,N_1775,N_639);
and U4441 (N_4441,N_94,N_152);
or U4442 (N_4442,N_2695,N_2453);
and U4443 (N_4443,N_815,N_2626);
or U4444 (N_4444,N_2875,N_87);
nor U4445 (N_4445,N_1114,N_2473);
nor U4446 (N_4446,N_745,N_1712);
and U4447 (N_4447,N_364,N_2558);
nor U4448 (N_4448,N_2163,N_2996);
and U4449 (N_4449,N_2925,N_1730);
xnor U4450 (N_4450,N_1832,N_1330);
or U4451 (N_4451,N_1183,N_452);
xnor U4452 (N_4452,N_1262,N_2845);
and U4453 (N_4453,N_241,N_2780);
nand U4454 (N_4454,N_708,N_2324);
and U4455 (N_4455,N_1926,N_1976);
or U4456 (N_4456,N_1689,N_484);
nand U4457 (N_4457,N_1059,N_11);
xor U4458 (N_4458,N_2776,N_1329);
xnor U4459 (N_4459,N_363,N_2296);
xor U4460 (N_4460,N_15,N_2811);
or U4461 (N_4461,N_1144,N_125);
and U4462 (N_4462,N_172,N_2267);
nand U4463 (N_4463,N_594,N_2077);
nand U4464 (N_4464,N_1631,N_1363);
xnor U4465 (N_4465,N_655,N_1132);
or U4466 (N_4466,N_2313,N_1048);
xor U4467 (N_4467,N_1360,N_1605);
xnor U4468 (N_4468,N_564,N_916);
and U4469 (N_4469,N_424,N_1980);
xor U4470 (N_4470,N_511,N_546);
nor U4471 (N_4471,N_2833,N_1337);
and U4472 (N_4472,N_1975,N_1816);
xor U4473 (N_4473,N_2818,N_2068);
and U4474 (N_4474,N_1418,N_1395);
and U4475 (N_4475,N_761,N_2614);
nor U4476 (N_4476,N_1813,N_2691);
and U4477 (N_4477,N_2305,N_1950);
nor U4478 (N_4478,N_2581,N_791);
xnor U4479 (N_4479,N_955,N_477);
nor U4480 (N_4480,N_151,N_1971);
nand U4481 (N_4481,N_1259,N_1432);
nor U4482 (N_4482,N_2616,N_1134);
nor U4483 (N_4483,N_2079,N_2327);
and U4484 (N_4484,N_2275,N_258);
and U4485 (N_4485,N_402,N_2566);
nand U4486 (N_4486,N_982,N_849);
nand U4487 (N_4487,N_1758,N_536);
nor U4488 (N_4488,N_1302,N_645);
and U4489 (N_4489,N_1042,N_1849);
nor U4490 (N_4490,N_1587,N_1002);
and U4491 (N_4491,N_2802,N_1224);
nor U4492 (N_4492,N_1986,N_265);
xor U4493 (N_4493,N_2001,N_2927);
nand U4494 (N_4494,N_683,N_1660);
and U4495 (N_4495,N_1305,N_1617);
or U4496 (N_4496,N_2229,N_2376);
xor U4497 (N_4497,N_1300,N_1350);
and U4498 (N_4498,N_1911,N_2602);
nand U4499 (N_4499,N_1401,N_2767);
nor U4500 (N_4500,N_1033,N_21);
and U4501 (N_4501,N_1680,N_2133);
xor U4502 (N_4502,N_302,N_2207);
and U4503 (N_4503,N_581,N_2029);
xnor U4504 (N_4504,N_2400,N_1318);
xnor U4505 (N_4505,N_1655,N_1885);
xnor U4506 (N_4506,N_1915,N_1773);
and U4507 (N_4507,N_581,N_20);
nand U4508 (N_4508,N_1342,N_1475);
xnor U4509 (N_4509,N_664,N_77);
or U4510 (N_4510,N_2756,N_1993);
xnor U4511 (N_4511,N_735,N_2025);
and U4512 (N_4512,N_1288,N_2150);
nor U4513 (N_4513,N_2646,N_2580);
or U4514 (N_4514,N_2533,N_1165);
nor U4515 (N_4515,N_315,N_826);
and U4516 (N_4516,N_547,N_896);
or U4517 (N_4517,N_2585,N_2394);
nor U4518 (N_4518,N_2999,N_2922);
nor U4519 (N_4519,N_1473,N_2299);
and U4520 (N_4520,N_1150,N_1726);
nor U4521 (N_4521,N_2529,N_1019);
nor U4522 (N_4522,N_276,N_686);
xor U4523 (N_4523,N_1996,N_801);
nor U4524 (N_4524,N_1373,N_234);
nand U4525 (N_4525,N_2198,N_1872);
nand U4526 (N_4526,N_2845,N_2160);
or U4527 (N_4527,N_230,N_61);
xnor U4528 (N_4528,N_657,N_163);
nand U4529 (N_4529,N_2410,N_222);
and U4530 (N_4530,N_22,N_602);
xor U4531 (N_4531,N_1749,N_412);
xor U4532 (N_4532,N_1642,N_1228);
nand U4533 (N_4533,N_506,N_2020);
nand U4534 (N_4534,N_1669,N_2470);
nand U4535 (N_4535,N_1816,N_329);
nor U4536 (N_4536,N_2410,N_2188);
and U4537 (N_4537,N_2164,N_849);
or U4538 (N_4538,N_1503,N_2189);
or U4539 (N_4539,N_2576,N_78);
nand U4540 (N_4540,N_74,N_1950);
nand U4541 (N_4541,N_1068,N_1647);
xnor U4542 (N_4542,N_591,N_1115);
xnor U4543 (N_4543,N_2557,N_1615);
nor U4544 (N_4544,N_2405,N_16);
nor U4545 (N_4545,N_1190,N_1700);
or U4546 (N_4546,N_1513,N_2398);
nand U4547 (N_4547,N_2460,N_60);
or U4548 (N_4548,N_1395,N_889);
or U4549 (N_4549,N_2361,N_1945);
and U4550 (N_4550,N_215,N_1932);
nand U4551 (N_4551,N_32,N_1604);
and U4552 (N_4552,N_1874,N_1979);
xnor U4553 (N_4553,N_283,N_267);
xor U4554 (N_4554,N_2873,N_2778);
nand U4555 (N_4555,N_153,N_1472);
or U4556 (N_4556,N_1339,N_742);
xor U4557 (N_4557,N_259,N_1046);
nor U4558 (N_4558,N_69,N_2392);
xnor U4559 (N_4559,N_1236,N_2602);
and U4560 (N_4560,N_2400,N_2085);
nor U4561 (N_4561,N_151,N_697);
and U4562 (N_4562,N_2501,N_2189);
nor U4563 (N_4563,N_1618,N_1131);
or U4564 (N_4564,N_1708,N_228);
or U4565 (N_4565,N_440,N_326);
nand U4566 (N_4566,N_2932,N_838);
nand U4567 (N_4567,N_1539,N_2506);
nor U4568 (N_4568,N_422,N_2569);
nor U4569 (N_4569,N_2397,N_2592);
and U4570 (N_4570,N_1338,N_2975);
nand U4571 (N_4571,N_1486,N_2091);
and U4572 (N_4572,N_2680,N_1746);
nand U4573 (N_4573,N_2176,N_1027);
and U4574 (N_4574,N_1664,N_2555);
nand U4575 (N_4575,N_1024,N_1043);
and U4576 (N_4576,N_1441,N_2076);
and U4577 (N_4577,N_300,N_93);
xor U4578 (N_4578,N_2773,N_1012);
xor U4579 (N_4579,N_2057,N_1139);
xor U4580 (N_4580,N_2599,N_451);
and U4581 (N_4581,N_443,N_794);
nor U4582 (N_4582,N_1252,N_2541);
or U4583 (N_4583,N_2333,N_2273);
and U4584 (N_4584,N_2229,N_2946);
xor U4585 (N_4585,N_1333,N_2689);
and U4586 (N_4586,N_1440,N_418);
xnor U4587 (N_4587,N_2157,N_1849);
and U4588 (N_4588,N_836,N_9);
nand U4589 (N_4589,N_212,N_2005);
and U4590 (N_4590,N_1329,N_29);
nand U4591 (N_4591,N_824,N_2981);
xor U4592 (N_4592,N_477,N_650);
or U4593 (N_4593,N_302,N_2217);
xnor U4594 (N_4594,N_1258,N_2112);
nor U4595 (N_4595,N_1225,N_1771);
and U4596 (N_4596,N_1614,N_819);
nor U4597 (N_4597,N_1089,N_2295);
nor U4598 (N_4598,N_173,N_2805);
nand U4599 (N_4599,N_484,N_160);
and U4600 (N_4600,N_2505,N_969);
and U4601 (N_4601,N_2591,N_2795);
nor U4602 (N_4602,N_2316,N_576);
and U4603 (N_4603,N_2785,N_2239);
or U4604 (N_4604,N_763,N_2478);
and U4605 (N_4605,N_1637,N_262);
nor U4606 (N_4606,N_2590,N_1320);
nor U4607 (N_4607,N_2416,N_1403);
nor U4608 (N_4608,N_1331,N_1539);
nor U4609 (N_4609,N_20,N_1844);
and U4610 (N_4610,N_2920,N_215);
nor U4611 (N_4611,N_1673,N_938);
nand U4612 (N_4612,N_2168,N_1682);
and U4613 (N_4613,N_2021,N_874);
xnor U4614 (N_4614,N_137,N_2444);
xnor U4615 (N_4615,N_2630,N_409);
and U4616 (N_4616,N_728,N_1912);
or U4617 (N_4617,N_2677,N_987);
nand U4618 (N_4618,N_2071,N_226);
xnor U4619 (N_4619,N_609,N_1351);
and U4620 (N_4620,N_2304,N_1589);
nor U4621 (N_4621,N_2657,N_1995);
nand U4622 (N_4622,N_1818,N_2563);
and U4623 (N_4623,N_2636,N_2383);
or U4624 (N_4624,N_1178,N_1767);
or U4625 (N_4625,N_1696,N_2085);
nand U4626 (N_4626,N_1120,N_1043);
or U4627 (N_4627,N_2001,N_2366);
or U4628 (N_4628,N_1203,N_2740);
nor U4629 (N_4629,N_1597,N_230);
nor U4630 (N_4630,N_2106,N_394);
nor U4631 (N_4631,N_1960,N_330);
nand U4632 (N_4632,N_1445,N_2337);
and U4633 (N_4633,N_2599,N_1606);
or U4634 (N_4634,N_279,N_2250);
nor U4635 (N_4635,N_978,N_2863);
xor U4636 (N_4636,N_909,N_1481);
nand U4637 (N_4637,N_1131,N_2160);
and U4638 (N_4638,N_150,N_1568);
nor U4639 (N_4639,N_915,N_1698);
nand U4640 (N_4640,N_822,N_2266);
and U4641 (N_4641,N_2019,N_706);
and U4642 (N_4642,N_2073,N_1417);
nand U4643 (N_4643,N_2655,N_1472);
nand U4644 (N_4644,N_1353,N_2413);
or U4645 (N_4645,N_1789,N_807);
and U4646 (N_4646,N_800,N_2163);
nor U4647 (N_4647,N_182,N_1714);
xnor U4648 (N_4648,N_1969,N_2677);
nand U4649 (N_4649,N_1444,N_2413);
nand U4650 (N_4650,N_2777,N_2155);
and U4651 (N_4651,N_2764,N_1578);
nand U4652 (N_4652,N_1302,N_1687);
xor U4653 (N_4653,N_193,N_474);
nor U4654 (N_4654,N_2077,N_1356);
nor U4655 (N_4655,N_2836,N_79);
and U4656 (N_4656,N_664,N_1890);
and U4657 (N_4657,N_2343,N_941);
nor U4658 (N_4658,N_443,N_1819);
xnor U4659 (N_4659,N_1469,N_1047);
nor U4660 (N_4660,N_2017,N_595);
and U4661 (N_4661,N_1195,N_2990);
nor U4662 (N_4662,N_270,N_2103);
and U4663 (N_4663,N_613,N_197);
or U4664 (N_4664,N_1312,N_1902);
nor U4665 (N_4665,N_1213,N_1024);
xor U4666 (N_4666,N_2410,N_2888);
and U4667 (N_4667,N_1292,N_35);
and U4668 (N_4668,N_2578,N_2205);
nand U4669 (N_4669,N_918,N_247);
nand U4670 (N_4670,N_608,N_1988);
or U4671 (N_4671,N_2101,N_2082);
nand U4672 (N_4672,N_1318,N_1506);
nor U4673 (N_4673,N_1300,N_446);
nand U4674 (N_4674,N_35,N_1109);
nand U4675 (N_4675,N_1582,N_320);
xor U4676 (N_4676,N_1265,N_316);
nor U4677 (N_4677,N_76,N_698);
xnor U4678 (N_4678,N_1658,N_2448);
nand U4679 (N_4679,N_1958,N_144);
nor U4680 (N_4680,N_1152,N_446);
nor U4681 (N_4681,N_2762,N_2344);
xnor U4682 (N_4682,N_676,N_2362);
nor U4683 (N_4683,N_1821,N_1361);
or U4684 (N_4684,N_1096,N_1204);
xor U4685 (N_4685,N_292,N_2188);
xnor U4686 (N_4686,N_85,N_2000);
xor U4687 (N_4687,N_2395,N_1450);
xor U4688 (N_4688,N_701,N_1386);
and U4689 (N_4689,N_1392,N_2926);
nand U4690 (N_4690,N_1962,N_1867);
nor U4691 (N_4691,N_1297,N_1621);
nor U4692 (N_4692,N_195,N_313);
or U4693 (N_4693,N_143,N_2150);
nor U4694 (N_4694,N_1206,N_1040);
xnor U4695 (N_4695,N_735,N_1997);
and U4696 (N_4696,N_395,N_1425);
or U4697 (N_4697,N_357,N_1056);
and U4698 (N_4698,N_1034,N_613);
and U4699 (N_4699,N_1703,N_896);
or U4700 (N_4700,N_69,N_1039);
and U4701 (N_4701,N_1749,N_1708);
nor U4702 (N_4702,N_1693,N_2461);
and U4703 (N_4703,N_495,N_1469);
nand U4704 (N_4704,N_303,N_1020);
nand U4705 (N_4705,N_493,N_691);
nor U4706 (N_4706,N_550,N_2478);
nor U4707 (N_4707,N_2834,N_345);
nand U4708 (N_4708,N_530,N_1662);
and U4709 (N_4709,N_1384,N_455);
nand U4710 (N_4710,N_1364,N_1207);
nor U4711 (N_4711,N_1474,N_462);
xnor U4712 (N_4712,N_567,N_14);
xor U4713 (N_4713,N_1121,N_2525);
nand U4714 (N_4714,N_371,N_2295);
and U4715 (N_4715,N_2202,N_823);
nor U4716 (N_4716,N_2028,N_2197);
xor U4717 (N_4717,N_306,N_107);
and U4718 (N_4718,N_758,N_1363);
or U4719 (N_4719,N_424,N_45);
nor U4720 (N_4720,N_2525,N_244);
nor U4721 (N_4721,N_403,N_2113);
and U4722 (N_4722,N_158,N_1898);
and U4723 (N_4723,N_1104,N_1353);
xor U4724 (N_4724,N_1663,N_444);
nand U4725 (N_4725,N_2193,N_107);
and U4726 (N_4726,N_1524,N_1195);
nor U4727 (N_4727,N_1605,N_605);
xor U4728 (N_4728,N_631,N_913);
or U4729 (N_4729,N_1439,N_1918);
and U4730 (N_4730,N_2573,N_2525);
nand U4731 (N_4731,N_865,N_393);
or U4732 (N_4732,N_2395,N_800);
nor U4733 (N_4733,N_1769,N_2363);
nand U4734 (N_4734,N_718,N_796);
nand U4735 (N_4735,N_2445,N_965);
nand U4736 (N_4736,N_445,N_914);
nor U4737 (N_4737,N_1598,N_1305);
and U4738 (N_4738,N_1044,N_2060);
and U4739 (N_4739,N_2986,N_812);
and U4740 (N_4740,N_718,N_2887);
nand U4741 (N_4741,N_2048,N_1261);
xor U4742 (N_4742,N_931,N_1311);
xnor U4743 (N_4743,N_2316,N_1532);
nand U4744 (N_4744,N_1542,N_1549);
or U4745 (N_4745,N_2174,N_696);
and U4746 (N_4746,N_794,N_1338);
or U4747 (N_4747,N_2904,N_2484);
nor U4748 (N_4748,N_1987,N_2619);
nor U4749 (N_4749,N_2846,N_1441);
xor U4750 (N_4750,N_75,N_25);
xnor U4751 (N_4751,N_2113,N_2772);
and U4752 (N_4752,N_2196,N_1191);
and U4753 (N_4753,N_2890,N_295);
or U4754 (N_4754,N_2741,N_1932);
and U4755 (N_4755,N_1071,N_377);
or U4756 (N_4756,N_1339,N_2853);
or U4757 (N_4757,N_2483,N_1764);
and U4758 (N_4758,N_888,N_1643);
xor U4759 (N_4759,N_457,N_1595);
nor U4760 (N_4760,N_2853,N_891);
and U4761 (N_4761,N_2261,N_1839);
and U4762 (N_4762,N_1110,N_2245);
nand U4763 (N_4763,N_2826,N_1202);
xor U4764 (N_4764,N_569,N_2155);
and U4765 (N_4765,N_2141,N_2189);
or U4766 (N_4766,N_1872,N_1538);
and U4767 (N_4767,N_52,N_456);
and U4768 (N_4768,N_1155,N_1152);
nand U4769 (N_4769,N_474,N_1837);
and U4770 (N_4770,N_1074,N_898);
nand U4771 (N_4771,N_355,N_2847);
nor U4772 (N_4772,N_1675,N_2342);
or U4773 (N_4773,N_359,N_1737);
nand U4774 (N_4774,N_1504,N_1270);
nor U4775 (N_4775,N_2112,N_1815);
nand U4776 (N_4776,N_507,N_1990);
nor U4777 (N_4777,N_1022,N_605);
xnor U4778 (N_4778,N_2521,N_1803);
or U4779 (N_4779,N_2193,N_787);
nand U4780 (N_4780,N_2486,N_272);
or U4781 (N_4781,N_1353,N_974);
xor U4782 (N_4782,N_43,N_2695);
xnor U4783 (N_4783,N_1822,N_400);
nor U4784 (N_4784,N_2018,N_1330);
xor U4785 (N_4785,N_583,N_2855);
xnor U4786 (N_4786,N_2956,N_2694);
xor U4787 (N_4787,N_2152,N_1202);
and U4788 (N_4788,N_2555,N_991);
nor U4789 (N_4789,N_1494,N_1671);
nand U4790 (N_4790,N_1776,N_980);
nand U4791 (N_4791,N_567,N_1854);
xor U4792 (N_4792,N_1665,N_2887);
or U4793 (N_4793,N_1257,N_1715);
or U4794 (N_4794,N_1073,N_494);
nor U4795 (N_4795,N_658,N_2289);
or U4796 (N_4796,N_2990,N_1464);
and U4797 (N_4797,N_2567,N_1591);
nand U4798 (N_4798,N_1095,N_2334);
nand U4799 (N_4799,N_1461,N_2774);
xor U4800 (N_4800,N_1187,N_2242);
and U4801 (N_4801,N_1949,N_2389);
nand U4802 (N_4802,N_2568,N_909);
nor U4803 (N_4803,N_2710,N_2252);
nand U4804 (N_4804,N_1803,N_365);
nor U4805 (N_4805,N_1198,N_159);
nor U4806 (N_4806,N_1346,N_2488);
and U4807 (N_4807,N_1563,N_172);
nor U4808 (N_4808,N_2605,N_289);
nand U4809 (N_4809,N_951,N_2920);
nand U4810 (N_4810,N_1601,N_1205);
xnor U4811 (N_4811,N_1623,N_2776);
xor U4812 (N_4812,N_657,N_1735);
nand U4813 (N_4813,N_2535,N_645);
xor U4814 (N_4814,N_49,N_747);
nor U4815 (N_4815,N_1218,N_2842);
nor U4816 (N_4816,N_990,N_401);
xnor U4817 (N_4817,N_243,N_1919);
nand U4818 (N_4818,N_1271,N_824);
nand U4819 (N_4819,N_779,N_2726);
xor U4820 (N_4820,N_1820,N_2581);
and U4821 (N_4821,N_2695,N_2416);
xnor U4822 (N_4822,N_481,N_655);
and U4823 (N_4823,N_830,N_2576);
nor U4824 (N_4824,N_1458,N_1468);
or U4825 (N_4825,N_432,N_2975);
and U4826 (N_4826,N_417,N_345);
and U4827 (N_4827,N_2914,N_1043);
or U4828 (N_4828,N_2888,N_1693);
and U4829 (N_4829,N_1028,N_804);
nor U4830 (N_4830,N_1526,N_884);
or U4831 (N_4831,N_122,N_1260);
and U4832 (N_4832,N_451,N_296);
and U4833 (N_4833,N_873,N_2506);
and U4834 (N_4834,N_1304,N_1265);
nand U4835 (N_4835,N_1590,N_795);
nor U4836 (N_4836,N_245,N_64);
and U4837 (N_4837,N_626,N_462);
or U4838 (N_4838,N_2478,N_2138);
or U4839 (N_4839,N_723,N_2685);
xnor U4840 (N_4840,N_2111,N_2804);
or U4841 (N_4841,N_2087,N_2258);
xor U4842 (N_4842,N_2799,N_2968);
nor U4843 (N_4843,N_398,N_1699);
xnor U4844 (N_4844,N_701,N_1042);
nand U4845 (N_4845,N_1079,N_2009);
xnor U4846 (N_4846,N_2251,N_2914);
and U4847 (N_4847,N_649,N_740);
and U4848 (N_4848,N_1340,N_416);
or U4849 (N_4849,N_805,N_234);
nor U4850 (N_4850,N_667,N_2200);
xor U4851 (N_4851,N_235,N_1964);
nor U4852 (N_4852,N_2510,N_2737);
nor U4853 (N_4853,N_732,N_1282);
nand U4854 (N_4854,N_444,N_357);
nor U4855 (N_4855,N_7,N_1012);
nand U4856 (N_4856,N_1613,N_732);
nor U4857 (N_4857,N_47,N_53);
nor U4858 (N_4858,N_75,N_547);
and U4859 (N_4859,N_56,N_1796);
and U4860 (N_4860,N_1684,N_1028);
xnor U4861 (N_4861,N_802,N_2412);
or U4862 (N_4862,N_2218,N_2948);
nand U4863 (N_4863,N_2603,N_1618);
xnor U4864 (N_4864,N_1432,N_294);
nor U4865 (N_4865,N_2314,N_1701);
nand U4866 (N_4866,N_1265,N_1802);
nor U4867 (N_4867,N_725,N_1730);
nand U4868 (N_4868,N_1152,N_380);
nor U4869 (N_4869,N_1738,N_2738);
or U4870 (N_4870,N_656,N_2694);
xor U4871 (N_4871,N_1158,N_1491);
nor U4872 (N_4872,N_1749,N_426);
nor U4873 (N_4873,N_2254,N_1950);
nor U4874 (N_4874,N_2504,N_1038);
or U4875 (N_4875,N_2655,N_2744);
nor U4876 (N_4876,N_952,N_1359);
nor U4877 (N_4877,N_2922,N_1622);
xor U4878 (N_4878,N_1401,N_646);
xnor U4879 (N_4879,N_2377,N_734);
nor U4880 (N_4880,N_920,N_1205);
and U4881 (N_4881,N_1996,N_2569);
nand U4882 (N_4882,N_1384,N_266);
or U4883 (N_4883,N_272,N_1844);
or U4884 (N_4884,N_1569,N_1425);
xnor U4885 (N_4885,N_1524,N_1483);
or U4886 (N_4886,N_1914,N_855);
xnor U4887 (N_4887,N_250,N_2458);
xor U4888 (N_4888,N_1628,N_2830);
nor U4889 (N_4889,N_1179,N_961);
nor U4890 (N_4890,N_190,N_497);
nor U4891 (N_4891,N_2841,N_2677);
and U4892 (N_4892,N_1060,N_199);
or U4893 (N_4893,N_615,N_2093);
and U4894 (N_4894,N_1424,N_1305);
xnor U4895 (N_4895,N_2561,N_2936);
nand U4896 (N_4896,N_1658,N_177);
nor U4897 (N_4897,N_2196,N_226);
or U4898 (N_4898,N_2736,N_279);
or U4899 (N_4899,N_690,N_1592);
or U4900 (N_4900,N_1251,N_2905);
nor U4901 (N_4901,N_1065,N_1913);
and U4902 (N_4902,N_2033,N_1318);
and U4903 (N_4903,N_1395,N_1416);
nor U4904 (N_4904,N_870,N_162);
and U4905 (N_4905,N_2334,N_2043);
xor U4906 (N_4906,N_1661,N_508);
nand U4907 (N_4907,N_1367,N_821);
nor U4908 (N_4908,N_2616,N_1486);
or U4909 (N_4909,N_281,N_2032);
or U4910 (N_4910,N_1874,N_2140);
nand U4911 (N_4911,N_2054,N_1117);
and U4912 (N_4912,N_1963,N_361);
and U4913 (N_4913,N_938,N_1408);
or U4914 (N_4914,N_2728,N_2676);
nor U4915 (N_4915,N_780,N_2478);
nor U4916 (N_4916,N_1010,N_1435);
nand U4917 (N_4917,N_2225,N_940);
xnor U4918 (N_4918,N_2598,N_1861);
xnor U4919 (N_4919,N_261,N_2847);
nand U4920 (N_4920,N_2041,N_2746);
nand U4921 (N_4921,N_1775,N_267);
and U4922 (N_4922,N_1930,N_867);
xnor U4923 (N_4923,N_2675,N_2504);
xor U4924 (N_4924,N_1451,N_803);
or U4925 (N_4925,N_2600,N_2019);
nor U4926 (N_4926,N_1135,N_408);
or U4927 (N_4927,N_958,N_996);
and U4928 (N_4928,N_1548,N_2675);
nor U4929 (N_4929,N_528,N_2560);
xnor U4930 (N_4930,N_762,N_2197);
nand U4931 (N_4931,N_882,N_50);
nor U4932 (N_4932,N_1864,N_2397);
nor U4933 (N_4933,N_1410,N_78);
xnor U4934 (N_4934,N_2793,N_1552);
nand U4935 (N_4935,N_1132,N_1839);
or U4936 (N_4936,N_2142,N_251);
or U4937 (N_4937,N_1953,N_1770);
or U4938 (N_4938,N_2811,N_2877);
or U4939 (N_4939,N_51,N_1386);
and U4940 (N_4940,N_284,N_1951);
xnor U4941 (N_4941,N_2984,N_2112);
and U4942 (N_4942,N_1805,N_15);
or U4943 (N_4943,N_2063,N_625);
nor U4944 (N_4944,N_932,N_1864);
and U4945 (N_4945,N_451,N_2255);
xor U4946 (N_4946,N_2822,N_1142);
nor U4947 (N_4947,N_2596,N_753);
or U4948 (N_4948,N_586,N_1771);
or U4949 (N_4949,N_1692,N_1647);
nand U4950 (N_4950,N_2681,N_1658);
or U4951 (N_4951,N_1645,N_1381);
nor U4952 (N_4952,N_2312,N_2228);
or U4953 (N_4953,N_1608,N_1361);
nand U4954 (N_4954,N_691,N_850);
nand U4955 (N_4955,N_1817,N_2056);
and U4956 (N_4956,N_774,N_1628);
nor U4957 (N_4957,N_122,N_2691);
nor U4958 (N_4958,N_2753,N_247);
and U4959 (N_4959,N_2643,N_2591);
nor U4960 (N_4960,N_119,N_2108);
nand U4961 (N_4961,N_1464,N_1174);
nor U4962 (N_4962,N_456,N_2176);
xnor U4963 (N_4963,N_848,N_162);
nor U4964 (N_4964,N_2379,N_2975);
nor U4965 (N_4965,N_2505,N_354);
nand U4966 (N_4966,N_2453,N_504);
nand U4967 (N_4967,N_1452,N_1678);
nand U4968 (N_4968,N_580,N_37);
nand U4969 (N_4969,N_949,N_321);
xor U4970 (N_4970,N_2450,N_939);
xor U4971 (N_4971,N_1872,N_2335);
nand U4972 (N_4972,N_967,N_1600);
nand U4973 (N_4973,N_1444,N_2998);
and U4974 (N_4974,N_2047,N_1723);
or U4975 (N_4975,N_1383,N_643);
or U4976 (N_4976,N_629,N_942);
xnor U4977 (N_4977,N_395,N_2644);
nand U4978 (N_4978,N_666,N_1965);
or U4979 (N_4979,N_1561,N_1334);
or U4980 (N_4980,N_2845,N_692);
or U4981 (N_4981,N_2798,N_1624);
nand U4982 (N_4982,N_2570,N_218);
and U4983 (N_4983,N_2160,N_130);
nor U4984 (N_4984,N_2798,N_2467);
and U4985 (N_4985,N_374,N_1811);
nand U4986 (N_4986,N_1048,N_166);
nand U4987 (N_4987,N_34,N_1678);
nand U4988 (N_4988,N_2835,N_1349);
and U4989 (N_4989,N_2762,N_608);
nand U4990 (N_4990,N_2396,N_2463);
and U4991 (N_4991,N_554,N_1861);
nand U4992 (N_4992,N_1000,N_2918);
and U4993 (N_4993,N_2139,N_2801);
and U4994 (N_4994,N_1924,N_547);
nand U4995 (N_4995,N_2290,N_476);
xnor U4996 (N_4996,N_1217,N_642);
xnor U4997 (N_4997,N_452,N_2730);
and U4998 (N_4998,N_1595,N_2218);
nor U4999 (N_4999,N_1658,N_2372);
nor U5000 (N_5000,N_1466,N_2736);
nor U5001 (N_5001,N_244,N_1442);
and U5002 (N_5002,N_1471,N_1989);
nor U5003 (N_5003,N_2603,N_679);
nor U5004 (N_5004,N_702,N_1108);
nand U5005 (N_5005,N_1712,N_1266);
nor U5006 (N_5006,N_1882,N_5);
and U5007 (N_5007,N_2764,N_1674);
nor U5008 (N_5008,N_503,N_407);
nor U5009 (N_5009,N_169,N_2826);
nor U5010 (N_5010,N_961,N_2960);
nand U5011 (N_5011,N_2929,N_568);
or U5012 (N_5012,N_1595,N_2482);
nor U5013 (N_5013,N_2932,N_1730);
nor U5014 (N_5014,N_1505,N_2778);
xnor U5015 (N_5015,N_50,N_2867);
or U5016 (N_5016,N_1480,N_195);
xor U5017 (N_5017,N_2365,N_608);
nor U5018 (N_5018,N_723,N_598);
and U5019 (N_5019,N_2324,N_2758);
or U5020 (N_5020,N_260,N_1146);
or U5021 (N_5021,N_1561,N_1432);
nand U5022 (N_5022,N_1940,N_1765);
xor U5023 (N_5023,N_551,N_33);
nand U5024 (N_5024,N_549,N_1452);
xor U5025 (N_5025,N_1573,N_284);
or U5026 (N_5026,N_2505,N_473);
xor U5027 (N_5027,N_1378,N_2488);
nor U5028 (N_5028,N_2310,N_2560);
or U5029 (N_5029,N_1513,N_1389);
and U5030 (N_5030,N_1933,N_2155);
nand U5031 (N_5031,N_456,N_939);
nor U5032 (N_5032,N_2155,N_2762);
or U5033 (N_5033,N_633,N_172);
or U5034 (N_5034,N_2538,N_1247);
nor U5035 (N_5035,N_1540,N_1355);
and U5036 (N_5036,N_2855,N_2315);
xor U5037 (N_5037,N_2173,N_164);
xnor U5038 (N_5038,N_65,N_2565);
xnor U5039 (N_5039,N_1040,N_1257);
xnor U5040 (N_5040,N_2172,N_567);
or U5041 (N_5041,N_231,N_1269);
nand U5042 (N_5042,N_2174,N_1660);
nand U5043 (N_5043,N_2938,N_525);
and U5044 (N_5044,N_63,N_17);
xor U5045 (N_5045,N_2254,N_2531);
and U5046 (N_5046,N_2989,N_695);
and U5047 (N_5047,N_2670,N_1259);
nor U5048 (N_5048,N_1352,N_1913);
nand U5049 (N_5049,N_937,N_2801);
or U5050 (N_5050,N_1921,N_270);
and U5051 (N_5051,N_2795,N_2358);
xnor U5052 (N_5052,N_2966,N_1290);
nor U5053 (N_5053,N_2239,N_1623);
xnor U5054 (N_5054,N_194,N_1036);
xnor U5055 (N_5055,N_1897,N_1180);
nand U5056 (N_5056,N_2825,N_1807);
and U5057 (N_5057,N_2371,N_478);
and U5058 (N_5058,N_2283,N_526);
nand U5059 (N_5059,N_531,N_1098);
nor U5060 (N_5060,N_1949,N_834);
and U5061 (N_5061,N_752,N_27);
nor U5062 (N_5062,N_2887,N_1363);
and U5063 (N_5063,N_936,N_1970);
and U5064 (N_5064,N_2370,N_2843);
nor U5065 (N_5065,N_1891,N_2372);
nor U5066 (N_5066,N_1606,N_1217);
and U5067 (N_5067,N_1942,N_2869);
and U5068 (N_5068,N_1859,N_1);
xnor U5069 (N_5069,N_2687,N_1835);
and U5070 (N_5070,N_317,N_1321);
or U5071 (N_5071,N_1525,N_1712);
nor U5072 (N_5072,N_538,N_2585);
nand U5073 (N_5073,N_944,N_812);
and U5074 (N_5074,N_367,N_840);
xnor U5075 (N_5075,N_1611,N_680);
or U5076 (N_5076,N_905,N_2289);
nand U5077 (N_5077,N_1104,N_272);
and U5078 (N_5078,N_2816,N_6);
or U5079 (N_5079,N_1477,N_2637);
nand U5080 (N_5080,N_1657,N_1748);
nor U5081 (N_5081,N_2889,N_1306);
nand U5082 (N_5082,N_440,N_2926);
xor U5083 (N_5083,N_479,N_2431);
and U5084 (N_5084,N_1057,N_736);
xnor U5085 (N_5085,N_405,N_1185);
xnor U5086 (N_5086,N_312,N_120);
and U5087 (N_5087,N_1530,N_1509);
nor U5088 (N_5088,N_387,N_1339);
and U5089 (N_5089,N_2021,N_273);
xor U5090 (N_5090,N_2360,N_804);
or U5091 (N_5091,N_1658,N_2796);
xnor U5092 (N_5092,N_2643,N_736);
and U5093 (N_5093,N_2960,N_1700);
xor U5094 (N_5094,N_747,N_2736);
xnor U5095 (N_5095,N_553,N_2671);
and U5096 (N_5096,N_846,N_64);
nor U5097 (N_5097,N_2343,N_1355);
xnor U5098 (N_5098,N_2955,N_1788);
xnor U5099 (N_5099,N_268,N_1348);
nor U5100 (N_5100,N_469,N_1572);
nor U5101 (N_5101,N_2990,N_2852);
nor U5102 (N_5102,N_1017,N_1237);
and U5103 (N_5103,N_1585,N_2178);
nand U5104 (N_5104,N_629,N_377);
and U5105 (N_5105,N_1244,N_1383);
and U5106 (N_5106,N_96,N_728);
or U5107 (N_5107,N_2252,N_109);
and U5108 (N_5108,N_124,N_940);
and U5109 (N_5109,N_1327,N_2108);
or U5110 (N_5110,N_2354,N_1357);
or U5111 (N_5111,N_2967,N_1601);
nor U5112 (N_5112,N_407,N_106);
xnor U5113 (N_5113,N_718,N_1581);
and U5114 (N_5114,N_1230,N_1191);
nand U5115 (N_5115,N_2567,N_475);
nor U5116 (N_5116,N_534,N_1157);
nand U5117 (N_5117,N_2923,N_2937);
or U5118 (N_5118,N_2181,N_2405);
nand U5119 (N_5119,N_1308,N_2458);
nor U5120 (N_5120,N_2768,N_2176);
nand U5121 (N_5121,N_2109,N_2190);
nor U5122 (N_5122,N_225,N_1499);
nor U5123 (N_5123,N_1978,N_1937);
nor U5124 (N_5124,N_699,N_2107);
and U5125 (N_5125,N_1684,N_1295);
and U5126 (N_5126,N_628,N_1985);
xnor U5127 (N_5127,N_2610,N_1420);
and U5128 (N_5128,N_1431,N_1865);
nor U5129 (N_5129,N_1144,N_1894);
and U5130 (N_5130,N_2667,N_262);
nand U5131 (N_5131,N_1010,N_631);
and U5132 (N_5132,N_1099,N_1096);
or U5133 (N_5133,N_559,N_2810);
or U5134 (N_5134,N_1690,N_521);
or U5135 (N_5135,N_1176,N_2776);
or U5136 (N_5136,N_2261,N_106);
and U5137 (N_5137,N_1138,N_1744);
xnor U5138 (N_5138,N_1926,N_1122);
nor U5139 (N_5139,N_1453,N_627);
and U5140 (N_5140,N_106,N_2752);
nand U5141 (N_5141,N_468,N_1739);
nand U5142 (N_5142,N_2152,N_203);
nor U5143 (N_5143,N_1966,N_548);
and U5144 (N_5144,N_230,N_976);
xor U5145 (N_5145,N_1843,N_2679);
and U5146 (N_5146,N_261,N_2871);
or U5147 (N_5147,N_1759,N_533);
xnor U5148 (N_5148,N_2789,N_2218);
nor U5149 (N_5149,N_2756,N_2288);
and U5150 (N_5150,N_2050,N_2614);
and U5151 (N_5151,N_2892,N_1179);
nor U5152 (N_5152,N_951,N_2798);
nand U5153 (N_5153,N_649,N_1430);
xor U5154 (N_5154,N_2646,N_1755);
xnor U5155 (N_5155,N_41,N_2);
and U5156 (N_5156,N_2653,N_2892);
nand U5157 (N_5157,N_870,N_1391);
nand U5158 (N_5158,N_1566,N_192);
nor U5159 (N_5159,N_2521,N_2444);
nor U5160 (N_5160,N_1485,N_1675);
nand U5161 (N_5161,N_1458,N_2929);
nand U5162 (N_5162,N_2770,N_1933);
and U5163 (N_5163,N_220,N_2255);
nand U5164 (N_5164,N_2090,N_726);
nor U5165 (N_5165,N_1370,N_114);
or U5166 (N_5166,N_364,N_2746);
nand U5167 (N_5167,N_2024,N_1050);
and U5168 (N_5168,N_1087,N_2191);
nand U5169 (N_5169,N_1947,N_606);
nand U5170 (N_5170,N_953,N_685);
xnor U5171 (N_5171,N_1128,N_715);
nand U5172 (N_5172,N_827,N_95);
and U5173 (N_5173,N_703,N_633);
and U5174 (N_5174,N_1704,N_1353);
xor U5175 (N_5175,N_2897,N_191);
or U5176 (N_5176,N_2817,N_1183);
or U5177 (N_5177,N_687,N_368);
xor U5178 (N_5178,N_2090,N_1123);
or U5179 (N_5179,N_301,N_556);
nand U5180 (N_5180,N_1288,N_885);
nor U5181 (N_5181,N_712,N_1676);
xnor U5182 (N_5182,N_1119,N_2790);
nor U5183 (N_5183,N_2278,N_321);
xnor U5184 (N_5184,N_2319,N_545);
nor U5185 (N_5185,N_1902,N_865);
nand U5186 (N_5186,N_1810,N_2253);
nor U5187 (N_5187,N_473,N_1557);
nor U5188 (N_5188,N_554,N_2028);
nand U5189 (N_5189,N_1318,N_2131);
and U5190 (N_5190,N_2279,N_1617);
and U5191 (N_5191,N_1403,N_1902);
xnor U5192 (N_5192,N_2536,N_2571);
or U5193 (N_5193,N_1852,N_1886);
nand U5194 (N_5194,N_2408,N_1002);
xnor U5195 (N_5195,N_1134,N_1464);
xor U5196 (N_5196,N_1608,N_1586);
xnor U5197 (N_5197,N_2345,N_1297);
nand U5198 (N_5198,N_791,N_1436);
and U5199 (N_5199,N_1045,N_1404);
and U5200 (N_5200,N_2804,N_63);
nor U5201 (N_5201,N_925,N_914);
xnor U5202 (N_5202,N_2647,N_2095);
and U5203 (N_5203,N_2672,N_1296);
and U5204 (N_5204,N_367,N_2308);
xnor U5205 (N_5205,N_947,N_761);
and U5206 (N_5206,N_2559,N_946);
nor U5207 (N_5207,N_1699,N_302);
or U5208 (N_5208,N_777,N_2598);
xnor U5209 (N_5209,N_2838,N_2023);
nor U5210 (N_5210,N_2519,N_881);
xor U5211 (N_5211,N_1261,N_1990);
nand U5212 (N_5212,N_2214,N_2265);
and U5213 (N_5213,N_2882,N_2026);
or U5214 (N_5214,N_744,N_2847);
xor U5215 (N_5215,N_726,N_2480);
or U5216 (N_5216,N_1763,N_109);
xnor U5217 (N_5217,N_2662,N_527);
xnor U5218 (N_5218,N_364,N_1423);
or U5219 (N_5219,N_1734,N_1356);
and U5220 (N_5220,N_416,N_2515);
nand U5221 (N_5221,N_2754,N_1912);
nor U5222 (N_5222,N_1996,N_1953);
and U5223 (N_5223,N_1425,N_2319);
or U5224 (N_5224,N_662,N_2415);
and U5225 (N_5225,N_2316,N_334);
xnor U5226 (N_5226,N_40,N_260);
and U5227 (N_5227,N_2344,N_128);
xor U5228 (N_5228,N_1994,N_283);
and U5229 (N_5229,N_2900,N_246);
nand U5230 (N_5230,N_2935,N_2986);
and U5231 (N_5231,N_1051,N_808);
and U5232 (N_5232,N_375,N_1323);
or U5233 (N_5233,N_525,N_719);
nor U5234 (N_5234,N_1744,N_96);
nand U5235 (N_5235,N_1173,N_1611);
xor U5236 (N_5236,N_739,N_1380);
nand U5237 (N_5237,N_483,N_2480);
or U5238 (N_5238,N_1446,N_2464);
nor U5239 (N_5239,N_555,N_1538);
and U5240 (N_5240,N_835,N_45);
and U5241 (N_5241,N_2333,N_697);
or U5242 (N_5242,N_2605,N_1128);
nand U5243 (N_5243,N_134,N_308);
nand U5244 (N_5244,N_2701,N_2342);
or U5245 (N_5245,N_2112,N_1223);
nor U5246 (N_5246,N_2363,N_2716);
and U5247 (N_5247,N_813,N_2690);
xor U5248 (N_5248,N_2233,N_1523);
nor U5249 (N_5249,N_1813,N_178);
xnor U5250 (N_5250,N_236,N_1297);
xor U5251 (N_5251,N_1097,N_1083);
and U5252 (N_5252,N_996,N_422);
and U5253 (N_5253,N_730,N_729);
nor U5254 (N_5254,N_668,N_1330);
xnor U5255 (N_5255,N_532,N_385);
nand U5256 (N_5256,N_176,N_462);
or U5257 (N_5257,N_1830,N_202);
or U5258 (N_5258,N_2430,N_2699);
and U5259 (N_5259,N_389,N_686);
nand U5260 (N_5260,N_1740,N_1565);
or U5261 (N_5261,N_1416,N_2487);
or U5262 (N_5262,N_1224,N_878);
nor U5263 (N_5263,N_2531,N_342);
xor U5264 (N_5264,N_2549,N_490);
and U5265 (N_5265,N_2515,N_2758);
nor U5266 (N_5266,N_1040,N_1332);
xor U5267 (N_5267,N_638,N_215);
nor U5268 (N_5268,N_916,N_2313);
and U5269 (N_5269,N_1660,N_1404);
nor U5270 (N_5270,N_834,N_2141);
and U5271 (N_5271,N_2005,N_470);
nand U5272 (N_5272,N_1545,N_2919);
and U5273 (N_5273,N_211,N_1225);
and U5274 (N_5274,N_1115,N_1238);
and U5275 (N_5275,N_371,N_593);
and U5276 (N_5276,N_748,N_1035);
nand U5277 (N_5277,N_2625,N_1579);
or U5278 (N_5278,N_2526,N_673);
and U5279 (N_5279,N_926,N_2012);
nor U5280 (N_5280,N_1717,N_1853);
and U5281 (N_5281,N_2568,N_309);
xnor U5282 (N_5282,N_1981,N_312);
xnor U5283 (N_5283,N_1678,N_312);
nand U5284 (N_5284,N_2852,N_396);
xnor U5285 (N_5285,N_271,N_2113);
nor U5286 (N_5286,N_2395,N_835);
xnor U5287 (N_5287,N_1448,N_2230);
or U5288 (N_5288,N_598,N_1693);
nand U5289 (N_5289,N_2770,N_1458);
and U5290 (N_5290,N_2962,N_1520);
nand U5291 (N_5291,N_851,N_1829);
xor U5292 (N_5292,N_118,N_2007);
or U5293 (N_5293,N_902,N_1960);
or U5294 (N_5294,N_2898,N_1719);
or U5295 (N_5295,N_1804,N_2239);
nor U5296 (N_5296,N_1505,N_1732);
and U5297 (N_5297,N_2472,N_2876);
xor U5298 (N_5298,N_2419,N_1355);
nor U5299 (N_5299,N_925,N_1434);
nand U5300 (N_5300,N_23,N_762);
xor U5301 (N_5301,N_1863,N_1792);
or U5302 (N_5302,N_834,N_2930);
or U5303 (N_5303,N_2312,N_2368);
and U5304 (N_5304,N_3,N_1565);
and U5305 (N_5305,N_1790,N_2970);
nor U5306 (N_5306,N_1896,N_1153);
nand U5307 (N_5307,N_1092,N_340);
or U5308 (N_5308,N_2894,N_328);
xnor U5309 (N_5309,N_1718,N_2036);
nor U5310 (N_5310,N_1438,N_2975);
xnor U5311 (N_5311,N_2156,N_969);
or U5312 (N_5312,N_173,N_1749);
and U5313 (N_5313,N_127,N_2360);
nor U5314 (N_5314,N_221,N_2980);
nor U5315 (N_5315,N_2138,N_1473);
and U5316 (N_5316,N_931,N_1028);
xnor U5317 (N_5317,N_2288,N_2748);
nor U5318 (N_5318,N_1482,N_1378);
xnor U5319 (N_5319,N_1342,N_1309);
nand U5320 (N_5320,N_2337,N_1214);
or U5321 (N_5321,N_771,N_950);
nand U5322 (N_5322,N_838,N_2971);
and U5323 (N_5323,N_574,N_496);
and U5324 (N_5324,N_1071,N_233);
nand U5325 (N_5325,N_1575,N_336);
xor U5326 (N_5326,N_2242,N_477);
and U5327 (N_5327,N_2863,N_675);
nor U5328 (N_5328,N_1159,N_2928);
nor U5329 (N_5329,N_2343,N_1198);
nor U5330 (N_5330,N_591,N_164);
xnor U5331 (N_5331,N_497,N_141);
nand U5332 (N_5332,N_1724,N_1718);
or U5333 (N_5333,N_1063,N_1956);
and U5334 (N_5334,N_2869,N_2136);
or U5335 (N_5335,N_2914,N_1961);
nor U5336 (N_5336,N_2320,N_2934);
nor U5337 (N_5337,N_2816,N_975);
and U5338 (N_5338,N_2071,N_2741);
and U5339 (N_5339,N_2063,N_656);
xor U5340 (N_5340,N_316,N_1018);
or U5341 (N_5341,N_2849,N_2533);
and U5342 (N_5342,N_97,N_736);
and U5343 (N_5343,N_2924,N_2270);
or U5344 (N_5344,N_278,N_2921);
nor U5345 (N_5345,N_2012,N_940);
nor U5346 (N_5346,N_2239,N_1586);
nor U5347 (N_5347,N_142,N_776);
nand U5348 (N_5348,N_2484,N_1880);
nand U5349 (N_5349,N_913,N_771);
xor U5350 (N_5350,N_1744,N_459);
and U5351 (N_5351,N_2628,N_125);
and U5352 (N_5352,N_1600,N_2407);
or U5353 (N_5353,N_2089,N_217);
nand U5354 (N_5354,N_2270,N_1107);
and U5355 (N_5355,N_314,N_302);
xor U5356 (N_5356,N_1613,N_2544);
xor U5357 (N_5357,N_309,N_717);
or U5358 (N_5358,N_2271,N_638);
nor U5359 (N_5359,N_2125,N_2652);
or U5360 (N_5360,N_1738,N_1051);
nor U5361 (N_5361,N_1461,N_2818);
nand U5362 (N_5362,N_2408,N_498);
nor U5363 (N_5363,N_1713,N_343);
nor U5364 (N_5364,N_1939,N_2905);
xor U5365 (N_5365,N_91,N_2620);
or U5366 (N_5366,N_2980,N_212);
nand U5367 (N_5367,N_1848,N_2903);
and U5368 (N_5368,N_1473,N_413);
and U5369 (N_5369,N_2934,N_628);
or U5370 (N_5370,N_2421,N_575);
nor U5371 (N_5371,N_220,N_1505);
xor U5372 (N_5372,N_490,N_1094);
or U5373 (N_5373,N_645,N_2123);
or U5374 (N_5374,N_165,N_41);
xor U5375 (N_5375,N_1994,N_2675);
nor U5376 (N_5376,N_1680,N_1489);
nor U5377 (N_5377,N_2595,N_2825);
nor U5378 (N_5378,N_1434,N_425);
or U5379 (N_5379,N_426,N_1547);
and U5380 (N_5380,N_1150,N_1427);
nand U5381 (N_5381,N_1624,N_2358);
xnor U5382 (N_5382,N_58,N_2585);
nand U5383 (N_5383,N_2593,N_2843);
nand U5384 (N_5384,N_2584,N_2534);
and U5385 (N_5385,N_1585,N_2331);
nor U5386 (N_5386,N_186,N_1586);
or U5387 (N_5387,N_1158,N_421);
or U5388 (N_5388,N_403,N_1014);
and U5389 (N_5389,N_2060,N_1291);
or U5390 (N_5390,N_952,N_1030);
nand U5391 (N_5391,N_2955,N_450);
nor U5392 (N_5392,N_2866,N_2024);
or U5393 (N_5393,N_874,N_718);
and U5394 (N_5394,N_304,N_2304);
nand U5395 (N_5395,N_1433,N_2641);
nand U5396 (N_5396,N_475,N_1197);
nor U5397 (N_5397,N_1372,N_785);
nor U5398 (N_5398,N_1600,N_346);
or U5399 (N_5399,N_2013,N_906);
nor U5400 (N_5400,N_2810,N_481);
xor U5401 (N_5401,N_1813,N_1144);
xor U5402 (N_5402,N_475,N_1742);
or U5403 (N_5403,N_589,N_1777);
or U5404 (N_5404,N_244,N_1588);
nor U5405 (N_5405,N_2479,N_693);
nand U5406 (N_5406,N_1502,N_29);
nor U5407 (N_5407,N_555,N_1370);
or U5408 (N_5408,N_504,N_293);
xor U5409 (N_5409,N_149,N_2855);
nor U5410 (N_5410,N_1993,N_2124);
nand U5411 (N_5411,N_2058,N_2789);
or U5412 (N_5412,N_1099,N_1840);
nor U5413 (N_5413,N_2819,N_738);
xor U5414 (N_5414,N_2182,N_2689);
xnor U5415 (N_5415,N_2229,N_549);
xnor U5416 (N_5416,N_624,N_1567);
nor U5417 (N_5417,N_1233,N_1152);
and U5418 (N_5418,N_51,N_1737);
nand U5419 (N_5419,N_1686,N_2032);
nor U5420 (N_5420,N_1120,N_1595);
xor U5421 (N_5421,N_1416,N_389);
nor U5422 (N_5422,N_2308,N_2494);
nor U5423 (N_5423,N_840,N_2968);
nor U5424 (N_5424,N_2851,N_2342);
nor U5425 (N_5425,N_1367,N_2911);
nand U5426 (N_5426,N_661,N_2302);
or U5427 (N_5427,N_2501,N_1914);
and U5428 (N_5428,N_2571,N_504);
or U5429 (N_5429,N_2366,N_2009);
nor U5430 (N_5430,N_1978,N_506);
nor U5431 (N_5431,N_2720,N_1916);
and U5432 (N_5432,N_2206,N_1879);
or U5433 (N_5433,N_2420,N_2107);
xnor U5434 (N_5434,N_263,N_478);
and U5435 (N_5435,N_2954,N_689);
and U5436 (N_5436,N_1377,N_2964);
or U5437 (N_5437,N_1354,N_488);
or U5438 (N_5438,N_2691,N_401);
or U5439 (N_5439,N_2962,N_2190);
nor U5440 (N_5440,N_1520,N_2154);
nor U5441 (N_5441,N_2034,N_1928);
or U5442 (N_5442,N_2705,N_2380);
or U5443 (N_5443,N_2997,N_1759);
or U5444 (N_5444,N_1325,N_263);
xor U5445 (N_5445,N_380,N_316);
nand U5446 (N_5446,N_2568,N_2309);
or U5447 (N_5447,N_2262,N_1715);
and U5448 (N_5448,N_98,N_1111);
nor U5449 (N_5449,N_2726,N_2368);
nand U5450 (N_5450,N_1419,N_1105);
nand U5451 (N_5451,N_13,N_393);
nand U5452 (N_5452,N_224,N_636);
xnor U5453 (N_5453,N_311,N_843);
nor U5454 (N_5454,N_2249,N_2168);
xor U5455 (N_5455,N_988,N_524);
or U5456 (N_5456,N_955,N_972);
nand U5457 (N_5457,N_1443,N_1082);
or U5458 (N_5458,N_163,N_616);
or U5459 (N_5459,N_941,N_1148);
and U5460 (N_5460,N_1488,N_928);
and U5461 (N_5461,N_2889,N_2007);
or U5462 (N_5462,N_2706,N_180);
and U5463 (N_5463,N_758,N_1115);
xor U5464 (N_5464,N_1409,N_258);
nor U5465 (N_5465,N_1072,N_903);
xor U5466 (N_5466,N_1633,N_2177);
and U5467 (N_5467,N_131,N_951);
nand U5468 (N_5468,N_2060,N_994);
xor U5469 (N_5469,N_1794,N_2919);
xnor U5470 (N_5470,N_1966,N_1143);
nor U5471 (N_5471,N_694,N_1707);
nor U5472 (N_5472,N_2956,N_2334);
nand U5473 (N_5473,N_2750,N_1023);
nor U5474 (N_5474,N_1672,N_1692);
and U5475 (N_5475,N_1091,N_2255);
xnor U5476 (N_5476,N_335,N_2340);
nand U5477 (N_5477,N_1778,N_1459);
nand U5478 (N_5478,N_107,N_1995);
nand U5479 (N_5479,N_2352,N_1395);
xnor U5480 (N_5480,N_819,N_2206);
nand U5481 (N_5481,N_1744,N_2899);
xor U5482 (N_5482,N_827,N_695);
nor U5483 (N_5483,N_1977,N_1618);
xnor U5484 (N_5484,N_2082,N_1504);
or U5485 (N_5485,N_586,N_640);
nor U5486 (N_5486,N_2028,N_2878);
or U5487 (N_5487,N_903,N_408);
nand U5488 (N_5488,N_2771,N_1703);
xor U5489 (N_5489,N_770,N_1298);
or U5490 (N_5490,N_2919,N_769);
xor U5491 (N_5491,N_2242,N_1564);
nand U5492 (N_5492,N_2249,N_2027);
xnor U5493 (N_5493,N_1247,N_2670);
nor U5494 (N_5494,N_2751,N_862);
xor U5495 (N_5495,N_1275,N_563);
nand U5496 (N_5496,N_1270,N_1715);
and U5497 (N_5497,N_967,N_152);
nor U5498 (N_5498,N_549,N_744);
nor U5499 (N_5499,N_1670,N_1061);
xor U5500 (N_5500,N_682,N_1459);
xor U5501 (N_5501,N_2440,N_2992);
nand U5502 (N_5502,N_766,N_2274);
or U5503 (N_5503,N_2754,N_2995);
and U5504 (N_5504,N_2239,N_2550);
nand U5505 (N_5505,N_2790,N_2011);
nor U5506 (N_5506,N_2880,N_16);
xor U5507 (N_5507,N_0,N_438);
nor U5508 (N_5508,N_2528,N_730);
nor U5509 (N_5509,N_2338,N_1404);
or U5510 (N_5510,N_466,N_1980);
nand U5511 (N_5511,N_2960,N_1166);
xor U5512 (N_5512,N_1207,N_2279);
nand U5513 (N_5513,N_2629,N_17);
nor U5514 (N_5514,N_757,N_1261);
nand U5515 (N_5515,N_638,N_1072);
nand U5516 (N_5516,N_1045,N_1998);
xnor U5517 (N_5517,N_443,N_2862);
xor U5518 (N_5518,N_2178,N_1391);
nand U5519 (N_5519,N_1048,N_1087);
xor U5520 (N_5520,N_1528,N_402);
and U5521 (N_5521,N_2371,N_2863);
nand U5522 (N_5522,N_521,N_105);
xor U5523 (N_5523,N_1477,N_442);
or U5524 (N_5524,N_404,N_1360);
nand U5525 (N_5525,N_239,N_1574);
nor U5526 (N_5526,N_526,N_2789);
and U5527 (N_5527,N_654,N_1113);
nand U5528 (N_5528,N_2242,N_2370);
nand U5529 (N_5529,N_2675,N_2281);
nand U5530 (N_5530,N_2172,N_57);
or U5531 (N_5531,N_2945,N_476);
nor U5532 (N_5532,N_644,N_858);
and U5533 (N_5533,N_2927,N_340);
and U5534 (N_5534,N_435,N_2794);
nand U5535 (N_5535,N_846,N_2064);
and U5536 (N_5536,N_134,N_2695);
xnor U5537 (N_5537,N_1225,N_2093);
or U5538 (N_5538,N_1134,N_1410);
and U5539 (N_5539,N_654,N_281);
xnor U5540 (N_5540,N_1803,N_1104);
xnor U5541 (N_5541,N_2949,N_351);
xnor U5542 (N_5542,N_1134,N_958);
xor U5543 (N_5543,N_2805,N_2258);
and U5544 (N_5544,N_2861,N_519);
xor U5545 (N_5545,N_2507,N_1206);
xnor U5546 (N_5546,N_924,N_1467);
xnor U5547 (N_5547,N_1995,N_1040);
nor U5548 (N_5548,N_2915,N_1146);
nand U5549 (N_5549,N_725,N_1015);
nor U5550 (N_5550,N_1310,N_934);
or U5551 (N_5551,N_816,N_1508);
nand U5552 (N_5552,N_2996,N_273);
xor U5553 (N_5553,N_115,N_2712);
nand U5554 (N_5554,N_625,N_1340);
or U5555 (N_5555,N_2251,N_1121);
and U5556 (N_5556,N_2228,N_361);
nand U5557 (N_5557,N_2009,N_1852);
nor U5558 (N_5558,N_901,N_316);
nand U5559 (N_5559,N_2839,N_945);
nand U5560 (N_5560,N_2532,N_2779);
xor U5561 (N_5561,N_677,N_1268);
nand U5562 (N_5562,N_748,N_1943);
or U5563 (N_5563,N_2077,N_2218);
or U5564 (N_5564,N_2459,N_2015);
nand U5565 (N_5565,N_2350,N_743);
and U5566 (N_5566,N_462,N_2892);
xor U5567 (N_5567,N_1826,N_2174);
nor U5568 (N_5568,N_1820,N_2090);
xor U5569 (N_5569,N_910,N_126);
nor U5570 (N_5570,N_2369,N_1040);
or U5571 (N_5571,N_1495,N_1421);
and U5572 (N_5572,N_309,N_141);
xnor U5573 (N_5573,N_1590,N_1752);
nor U5574 (N_5574,N_2016,N_1824);
or U5575 (N_5575,N_2168,N_334);
or U5576 (N_5576,N_2190,N_933);
or U5577 (N_5577,N_183,N_1989);
nand U5578 (N_5578,N_1317,N_608);
nand U5579 (N_5579,N_2099,N_1288);
or U5580 (N_5580,N_1534,N_1258);
and U5581 (N_5581,N_1697,N_1647);
xor U5582 (N_5582,N_1698,N_2499);
xor U5583 (N_5583,N_1184,N_2314);
and U5584 (N_5584,N_39,N_2471);
nand U5585 (N_5585,N_2534,N_2331);
xnor U5586 (N_5586,N_2483,N_2821);
and U5587 (N_5587,N_1438,N_865);
nor U5588 (N_5588,N_483,N_2992);
nand U5589 (N_5589,N_1183,N_243);
nor U5590 (N_5590,N_381,N_842);
nand U5591 (N_5591,N_1092,N_1148);
or U5592 (N_5592,N_2984,N_1629);
xor U5593 (N_5593,N_19,N_2680);
xor U5594 (N_5594,N_484,N_1116);
nand U5595 (N_5595,N_2984,N_493);
and U5596 (N_5596,N_566,N_2899);
and U5597 (N_5597,N_492,N_2475);
nor U5598 (N_5598,N_675,N_2154);
xnor U5599 (N_5599,N_1375,N_2674);
nand U5600 (N_5600,N_156,N_2186);
or U5601 (N_5601,N_2694,N_1561);
nor U5602 (N_5602,N_465,N_2746);
nor U5603 (N_5603,N_2871,N_385);
nor U5604 (N_5604,N_2211,N_201);
xor U5605 (N_5605,N_1338,N_693);
xnor U5606 (N_5606,N_1654,N_13);
xnor U5607 (N_5607,N_1539,N_393);
and U5608 (N_5608,N_2803,N_2346);
xnor U5609 (N_5609,N_2644,N_1624);
nand U5610 (N_5610,N_2423,N_202);
and U5611 (N_5611,N_2992,N_2094);
nor U5612 (N_5612,N_2316,N_2013);
xor U5613 (N_5613,N_451,N_2314);
nand U5614 (N_5614,N_997,N_453);
nand U5615 (N_5615,N_1624,N_2676);
nand U5616 (N_5616,N_474,N_2026);
or U5617 (N_5617,N_1018,N_2129);
nor U5618 (N_5618,N_1395,N_2580);
nor U5619 (N_5619,N_2985,N_656);
nand U5620 (N_5620,N_2193,N_1314);
xor U5621 (N_5621,N_2588,N_1166);
nand U5622 (N_5622,N_713,N_11);
xnor U5623 (N_5623,N_10,N_2808);
xnor U5624 (N_5624,N_2795,N_1430);
xor U5625 (N_5625,N_2803,N_1700);
and U5626 (N_5626,N_595,N_312);
nand U5627 (N_5627,N_2935,N_199);
xor U5628 (N_5628,N_2425,N_265);
xor U5629 (N_5629,N_1931,N_516);
nor U5630 (N_5630,N_2071,N_962);
or U5631 (N_5631,N_2873,N_2673);
and U5632 (N_5632,N_1349,N_2113);
or U5633 (N_5633,N_2932,N_1362);
nor U5634 (N_5634,N_691,N_2556);
nor U5635 (N_5635,N_2784,N_1375);
or U5636 (N_5636,N_2437,N_1981);
and U5637 (N_5637,N_2066,N_1195);
xnor U5638 (N_5638,N_352,N_926);
and U5639 (N_5639,N_2000,N_1129);
or U5640 (N_5640,N_1538,N_361);
nand U5641 (N_5641,N_947,N_453);
nor U5642 (N_5642,N_2037,N_256);
and U5643 (N_5643,N_1516,N_436);
nor U5644 (N_5644,N_624,N_616);
xnor U5645 (N_5645,N_1017,N_1401);
nand U5646 (N_5646,N_2764,N_2934);
and U5647 (N_5647,N_977,N_948);
nand U5648 (N_5648,N_99,N_497);
nand U5649 (N_5649,N_2233,N_2471);
or U5650 (N_5650,N_977,N_733);
and U5651 (N_5651,N_455,N_1213);
nor U5652 (N_5652,N_587,N_1924);
nor U5653 (N_5653,N_2411,N_2142);
xnor U5654 (N_5654,N_1962,N_2997);
or U5655 (N_5655,N_756,N_1573);
nor U5656 (N_5656,N_1103,N_1869);
nor U5657 (N_5657,N_1414,N_1763);
or U5658 (N_5658,N_2468,N_1803);
nor U5659 (N_5659,N_2222,N_1304);
or U5660 (N_5660,N_1234,N_797);
nand U5661 (N_5661,N_2573,N_1957);
or U5662 (N_5662,N_333,N_1102);
or U5663 (N_5663,N_525,N_1201);
xnor U5664 (N_5664,N_984,N_565);
and U5665 (N_5665,N_614,N_668);
or U5666 (N_5666,N_471,N_190);
xor U5667 (N_5667,N_1645,N_1436);
and U5668 (N_5668,N_2668,N_185);
nand U5669 (N_5669,N_1691,N_1463);
nor U5670 (N_5670,N_2100,N_89);
and U5671 (N_5671,N_1854,N_2709);
nand U5672 (N_5672,N_2992,N_76);
xor U5673 (N_5673,N_1193,N_2779);
nor U5674 (N_5674,N_553,N_991);
or U5675 (N_5675,N_1387,N_1945);
and U5676 (N_5676,N_296,N_2709);
nand U5677 (N_5677,N_2337,N_2204);
nor U5678 (N_5678,N_1236,N_1845);
nor U5679 (N_5679,N_955,N_1475);
and U5680 (N_5680,N_1656,N_2473);
nor U5681 (N_5681,N_1532,N_239);
xor U5682 (N_5682,N_1101,N_2936);
or U5683 (N_5683,N_780,N_1269);
nand U5684 (N_5684,N_1841,N_2726);
nand U5685 (N_5685,N_1409,N_1685);
and U5686 (N_5686,N_1105,N_506);
and U5687 (N_5687,N_2870,N_730);
nand U5688 (N_5688,N_1707,N_177);
nor U5689 (N_5689,N_198,N_495);
nor U5690 (N_5690,N_2749,N_1910);
xor U5691 (N_5691,N_341,N_1496);
xor U5692 (N_5692,N_1344,N_2983);
xor U5693 (N_5693,N_2569,N_1816);
xnor U5694 (N_5694,N_1682,N_1232);
and U5695 (N_5695,N_1862,N_1048);
or U5696 (N_5696,N_83,N_2076);
or U5697 (N_5697,N_2903,N_318);
nor U5698 (N_5698,N_1160,N_2904);
and U5699 (N_5699,N_2379,N_2023);
nand U5700 (N_5700,N_1285,N_1722);
and U5701 (N_5701,N_1405,N_1916);
and U5702 (N_5702,N_2756,N_2457);
nor U5703 (N_5703,N_2839,N_105);
and U5704 (N_5704,N_1942,N_937);
nand U5705 (N_5705,N_354,N_2761);
nor U5706 (N_5706,N_9,N_1852);
nand U5707 (N_5707,N_997,N_1396);
xor U5708 (N_5708,N_2549,N_365);
and U5709 (N_5709,N_1715,N_1571);
xnor U5710 (N_5710,N_2643,N_2252);
or U5711 (N_5711,N_2370,N_1050);
xor U5712 (N_5712,N_2408,N_2587);
xor U5713 (N_5713,N_463,N_647);
or U5714 (N_5714,N_1919,N_1667);
and U5715 (N_5715,N_434,N_207);
or U5716 (N_5716,N_1054,N_1076);
nand U5717 (N_5717,N_2589,N_2656);
nand U5718 (N_5718,N_2283,N_1197);
nor U5719 (N_5719,N_952,N_1872);
nand U5720 (N_5720,N_1667,N_761);
and U5721 (N_5721,N_1347,N_469);
nand U5722 (N_5722,N_2504,N_586);
xor U5723 (N_5723,N_1144,N_2930);
xnor U5724 (N_5724,N_1874,N_1688);
nand U5725 (N_5725,N_1629,N_2593);
nor U5726 (N_5726,N_1619,N_2959);
or U5727 (N_5727,N_1250,N_2036);
and U5728 (N_5728,N_398,N_2756);
xnor U5729 (N_5729,N_1484,N_1098);
and U5730 (N_5730,N_2139,N_2833);
xor U5731 (N_5731,N_1359,N_1426);
nand U5732 (N_5732,N_1021,N_2827);
xor U5733 (N_5733,N_2454,N_1953);
xor U5734 (N_5734,N_249,N_312);
or U5735 (N_5735,N_1454,N_1464);
and U5736 (N_5736,N_1565,N_1287);
nor U5737 (N_5737,N_2403,N_498);
nand U5738 (N_5738,N_148,N_748);
and U5739 (N_5739,N_1029,N_2283);
xnor U5740 (N_5740,N_2142,N_1526);
or U5741 (N_5741,N_2190,N_1025);
nand U5742 (N_5742,N_46,N_2186);
or U5743 (N_5743,N_1462,N_441);
or U5744 (N_5744,N_519,N_223);
nand U5745 (N_5745,N_2323,N_345);
and U5746 (N_5746,N_2856,N_2616);
nand U5747 (N_5747,N_1381,N_1666);
xor U5748 (N_5748,N_2052,N_715);
and U5749 (N_5749,N_254,N_2953);
and U5750 (N_5750,N_493,N_2490);
nor U5751 (N_5751,N_302,N_297);
nor U5752 (N_5752,N_557,N_21);
xor U5753 (N_5753,N_1063,N_2618);
or U5754 (N_5754,N_675,N_772);
nand U5755 (N_5755,N_1821,N_1747);
and U5756 (N_5756,N_2890,N_1335);
nor U5757 (N_5757,N_1225,N_1101);
xnor U5758 (N_5758,N_151,N_2144);
or U5759 (N_5759,N_853,N_2594);
or U5760 (N_5760,N_591,N_2886);
or U5761 (N_5761,N_1498,N_633);
and U5762 (N_5762,N_777,N_1745);
nor U5763 (N_5763,N_1920,N_2667);
nand U5764 (N_5764,N_114,N_885);
nor U5765 (N_5765,N_2320,N_1089);
or U5766 (N_5766,N_524,N_309);
or U5767 (N_5767,N_1480,N_106);
and U5768 (N_5768,N_2407,N_1703);
nand U5769 (N_5769,N_1125,N_2713);
nand U5770 (N_5770,N_2743,N_642);
or U5771 (N_5771,N_780,N_1555);
or U5772 (N_5772,N_2531,N_2598);
nand U5773 (N_5773,N_1012,N_1700);
xor U5774 (N_5774,N_914,N_1882);
and U5775 (N_5775,N_706,N_1044);
nor U5776 (N_5776,N_2926,N_2246);
nand U5777 (N_5777,N_1981,N_2195);
or U5778 (N_5778,N_1959,N_2583);
xor U5779 (N_5779,N_750,N_1807);
xor U5780 (N_5780,N_2158,N_1751);
nand U5781 (N_5781,N_2329,N_1615);
or U5782 (N_5782,N_135,N_397);
and U5783 (N_5783,N_1443,N_2417);
nor U5784 (N_5784,N_39,N_578);
and U5785 (N_5785,N_1781,N_1366);
nor U5786 (N_5786,N_1372,N_2850);
or U5787 (N_5787,N_289,N_2531);
or U5788 (N_5788,N_2453,N_537);
or U5789 (N_5789,N_2396,N_2331);
nor U5790 (N_5790,N_995,N_434);
nand U5791 (N_5791,N_318,N_1374);
and U5792 (N_5792,N_2597,N_825);
or U5793 (N_5793,N_407,N_1287);
or U5794 (N_5794,N_1181,N_1208);
xor U5795 (N_5795,N_2425,N_626);
and U5796 (N_5796,N_227,N_2196);
nand U5797 (N_5797,N_17,N_2736);
xor U5798 (N_5798,N_835,N_1930);
and U5799 (N_5799,N_1127,N_1578);
and U5800 (N_5800,N_994,N_62);
or U5801 (N_5801,N_1205,N_1916);
nand U5802 (N_5802,N_2799,N_2852);
nor U5803 (N_5803,N_2818,N_281);
nor U5804 (N_5804,N_2231,N_766);
or U5805 (N_5805,N_571,N_591);
nand U5806 (N_5806,N_776,N_1650);
and U5807 (N_5807,N_2541,N_821);
and U5808 (N_5808,N_527,N_2538);
nand U5809 (N_5809,N_378,N_1775);
nor U5810 (N_5810,N_670,N_795);
nor U5811 (N_5811,N_2427,N_727);
nor U5812 (N_5812,N_39,N_2472);
nor U5813 (N_5813,N_2475,N_2645);
xnor U5814 (N_5814,N_1436,N_297);
or U5815 (N_5815,N_1916,N_1734);
and U5816 (N_5816,N_2421,N_869);
or U5817 (N_5817,N_2024,N_1414);
nand U5818 (N_5818,N_1823,N_2346);
and U5819 (N_5819,N_1638,N_888);
and U5820 (N_5820,N_2134,N_94);
or U5821 (N_5821,N_775,N_551);
nand U5822 (N_5822,N_1224,N_1162);
xnor U5823 (N_5823,N_612,N_2117);
nor U5824 (N_5824,N_2603,N_243);
and U5825 (N_5825,N_988,N_1127);
or U5826 (N_5826,N_925,N_2200);
or U5827 (N_5827,N_2501,N_1516);
nand U5828 (N_5828,N_1182,N_1920);
or U5829 (N_5829,N_2747,N_1742);
nor U5830 (N_5830,N_2530,N_2857);
xnor U5831 (N_5831,N_2878,N_1866);
and U5832 (N_5832,N_87,N_1489);
or U5833 (N_5833,N_1846,N_1617);
nand U5834 (N_5834,N_1880,N_249);
xor U5835 (N_5835,N_1530,N_1357);
nor U5836 (N_5836,N_2661,N_195);
or U5837 (N_5837,N_241,N_402);
or U5838 (N_5838,N_2356,N_2899);
and U5839 (N_5839,N_1473,N_1380);
xnor U5840 (N_5840,N_2477,N_316);
nand U5841 (N_5841,N_1728,N_824);
nor U5842 (N_5842,N_2847,N_202);
nand U5843 (N_5843,N_1815,N_2806);
nor U5844 (N_5844,N_1530,N_1956);
nand U5845 (N_5845,N_2905,N_2497);
nand U5846 (N_5846,N_2895,N_1172);
nor U5847 (N_5847,N_2782,N_69);
xnor U5848 (N_5848,N_1085,N_2434);
or U5849 (N_5849,N_2370,N_944);
nand U5850 (N_5850,N_2509,N_286);
or U5851 (N_5851,N_1860,N_2949);
and U5852 (N_5852,N_2364,N_246);
nand U5853 (N_5853,N_1828,N_1113);
and U5854 (N_5854,N_983,N_770);
and U5855 (N_5855,N_2577,N_2703);
and U5856 (N_5856,N_1520,N_1032);
nand U5857 (N_5857,N_1947,N_1899);
and U5858 (N_5858,N_853,N_1638);
xnor U5859 (N_5859,N_1523,N_1518);
xnor U5860 (N_5860,N_2109,N_1113);
nand U5861 (N_5861,N_1284,N_1288);
and U5862 (N_5862,N_578,N_2217);
nand U5863 (N_5863,N_2892,N_2559);
or U5864 (N_5864,N_861,N_1509);
nor U5865 (N_5865,N_2162,N_1206);
or U5866 (N_5866,N_1388,N_739);
nand U5867 (N_5867,N_2034,N_2605);
and U5868 (N_5868,N_2776,N_1282);
xnor U5869 (N_5869,N_1924,N_76);
and U5870 (N_5870,N_1356,N_377);
nor U5871 (N_5871,N_1391,N_1816);
nand U5872 (N_5872,N_2677,N_2014);
nand U5873 (N_5873,N_2058,N_1878);
or U5874 (N_5874,N_494,N_1087);
and U5875 (N_5875,N_2936,N_602);
or U5876 (N_5876,N_790,N_1545);
and U5877 (N_5877,N_873,N_2080);
nor U5878 (N_5878,N_2523,N_41);
and U5879 (N_5879,N_1549,N_125);
and U5880 (N_5880,N_1335,N_2459);
nand U5881 (N_5881,N_841,N_613);
nor U5882 (N_5882,N_1233,N_1869);
or U5883 (N_5883,N_2344,N_2026);
nor U5884 (N_5884,N_2873,N_1643);
nand U5885 (N_5885,N_1156,N_1330);
nor U5886 (N_5886,N_516,N_238);
and U5887 (N_5887,N_2881,N_2143);
nand U5888 (N_5888,N_1278,N_558);
nand U5889 (N_5889,N_2885,N_321);
nor U5890 (N_5890,N_47,N_141);
and U5891 (N_5891,N_1177,N_2712);
xor U5892 (N_5892,N_958,N_2516);
nand U5893 (N_5893,N_2615,N_1036);
or U5894 (N_5894,N_2362,N_1389);
nor U5895 (N_5895,N_2578,N_2454);
or U5896 (N_5896,N_660,N_178);
nor U5897 (N_5897,N_2522,N_1796);
nor U5898 (N_5898,N_317,N_1232);
nand U5899 (N_5899,N_832,N_2498);
nor U5900 (N_5900,N_482,N_1515);
nor U5901 (N_5901,N_753,N_1319);
xor U5902 (N_5902,N_358,N_2320);
and U5903 (N_5903,N_2477,N_2320);
and U5904 (N_5904,N_1960,N_2268);
nand U5905 (N_5905,N_1200,N_1964);
nand U5906 (N_5906,N_2876,N_2484);
nand U5907 (N_5907,N_153,N_367);
xor U5908 (N_5908,N_890,N_2385);
nand U5909 (N_5909,N_2872,N_2064);
nor U5910 (N_5910,N_569,N_2699);
nand U5911 (N_5911,N_380,N_1098);
nand U5912 (N_5912,N_1957,N_326);
nor U5913 (N_5913,N_874,N_2950);
nor U5914 (N_5914,N_1039,N_1114);
nor U5915 (N_5915,N_689,N_948);
nor U5916 (N_5916,N_257,N_1495);
nor U5917 (N_5917,N_1638,N_2406);
or U5918 (N_5918,N_670,N_2668);
nand U5919 (N_5919,N_972,N_318);
nor U5920 (N_5920,N_2836,N_888);
nand U5921 (N_5921,N_1326,N_771);
or U5922 (N_5922,N_259,N_1347);
nor U5923 (N_5923,N_1622,N_1327);
or U5924 (N_5924,N_1067,N_2506);
nor U5925 (N_5925,N_1576,N_2019);
and U5926 (N_5926,N_1450,N_1553);
nor U5927 (N_5927,N_2624,N_1178);
nor U5928 (N_5928,N_1556,N_513);
and U5929 (N_5929,N_1938,N_1256);
nand U5930 (N_5930,N_58,N_2324);
nor U5931 (N_5931,N_2329,N_348);
nand U5932 (N_5932,N_1370,N_71);
or U5933 (N_5933,N_670,N_1989);
nand U5934 (N_5934,N_1261,N_1918);
xor U5935 (N_5935,N_1414,N_2287);
nor U5936 (N_5936,N_2752,N_975);
nand U5937 (N_5937,N_296,N_1916);
xor U5938 (N_5938,N_349,N_2511);
nor U5939 (N_5939,N_412,N_1999);
or U5940 (N_5940,N_2783,N_2115);
nand U5941 (N_5941,N_2370,N_1808);
or U5942 (N_5942,N_1094,N_2145);
nand U5943 (N_5943,N_2530,N_2314);
nor U5944 (N_5944,N_1831,N_2954);
nor U5945 (N_5945,N_2776,N_18);
nand U5946 (N_5946,N_1107,N_1285);
or U5947 (N_5947,N_30,N_1847);
nor U5948 (N_5948,N_502,N_2421);
or U5949 (N_5949,N_706,N_141);
or U5950 (N_5950,N_2381,N_655);
nand U5951 (N_5951,N_828,N_1710);
or U5952 (N_5952,N_797,N_1169);
or U5953 (N_5953,N_787,N_1268);
or U5954 (N_5954,N_2461,N_885);
nand U5955 (N_5955,N_2312,N_2255);
nor U5956 (N_5956,N_2021,N_156);
xor U5957 (N_5957,N_1697,N_2009);
or U5958 (N_5958,N_148,N_1349);
and U5959 (N_5959,N_1329,N_1402);
and U5960 (N_5960,N_1351,N_733);
nor U5961 (N_5961,N_2798,N_894);
nor U5962 (N_5962,N_983,N_2047);
nor U5963 (N_5963,N_2061,N_683);
or U5964 (N_5964,N_400,N_759);
nor U5965 (N_5965,N_454,N_654);
or U5966 (N_5966,N_2418,N_2133);
nor U5967 (N_5967,N_1042,N_2991);
nand U5968 (N_5968,N_697,N_1546);
or U5969 (N_5969,N_1377,N_1792);
and U5970 (N_5970,N_2145,N_2630);
nor U5971 (N_5971,N_643,N_656);
or U5972 (N_5972,N_1544,N_1999);
or U5973 (N_5973,N_747,N_423);
or U5974 (N_5974,N_1706,N_2860);
xor U5975 (N_5975,N_1826,N_592);
or U5976 (N_5976,N_1945,N_916);
or U5977 (N_5977,N_2737,N_938);
xnor U5978 (N_5978,N_585,N_2570);
nand U5979 (N_5979,N_1687,N_843);
xor U5980 (N_5980,N_1065,N_1654);
nor U5981 (N_5981,N_1244,N_2450);
nor U5982 (N_5982,N_293,N_2681);
and U5983 (N_5983,N_2490,N_302);
nor U5984 (N_5984,N_328,N_145);
or U5985 (N_5985,N_96,N_145);
nor U5986 (N_5986,N_1649,N_1436);
and U5987 (N_5987,N_2010,N_299);
or U5988 (N_5988,N_1305,N_1705);
xor U5989 (N_5989,N_1742,N_1003);
or U5990 (N_5990,N_167,N_2364);
nand U5991 (N_5991,N_607,N_2936);
xnor U5992 (N_5992,N_2468,N_2922);
nor U5993 (N_5993,N_2361,N_1120);
or U5994 (N_5994,N_2422,N_814);
nand U5995 (N_5995,N_300,N_281);
or U5996 (N_5996,N_982,N_1682);
and U5997 (N_5997,N_2504,N_1647);
nand U5998 (N_5998,N_2959,N_1367);
nor U5999 (N_5999,N_2111,N_2057);
xor U6000 (N_6000,N_4578,N_3061);
nand U6001 (N_6001,N_4453,N_4925);
or U6002 (N_6002,N_5638,N_4900);
or U6003 (N_6003,N_4146,N_4889);
xor U6004 (N_6004,N_4892,N_5843);
nor U6005 (N_6005,N_4445,N_4316);
xor U6006 (N_6006,N_5018,N_4426);
and U6007 (N_6007,N_3319,N_3308);
and U6008 (N_6008,N_5025,N_4518);
xor U6009 (N_6009,N_3307,N_4456);
xor U6010 (N_6010,N_3444,N_4959);
xor U6011 (N_6011,N_4147,N_3321);
nor U6012 (N_6012,N_5789,N_5862);
or U6013 (N_6013,N_3610,N_5469);
or U6014 (N_6014,N_4512,N_5016);
and U6015 (N_6015,N_5803,N_4415);
or U6016 (N_6016,N_5474,N_4034);
and U6017 (N_6017,N_4565,N_5711);
and U6018 (N_6018,N_4843,N_4582);
and U6019 (N_6019,N_3630,N_4602);
and U6020 (N_6020,N_5952,N_5491);
nand U6021 (N_6021,N_4036,N_5530);
and U6022 (N_6022,N_5221,N_5657);
or U6023 (N_6023,N_5747,N_4965);
xnor U6024 (N_6024,N_5217,N_3130);
and U6025 (N_6025,N_3121,N_4293);
xor U6026 (N_6026,N_5886,N_3210);
and U6027 (N_6027,N_5556,N_4651);
and U6028 (N_6028,N_4035,N_4947);
or U6029 (N_6029,N_4044,N_4401);
nand U6030 (N_6030,N_3769,N_5997);
or U6031 (N_6031,N_3903,N_4275);
nand U6032 (N_6032,N_5623,N_3374);
and U6033 (N_6033,N_5444,N_5204);
nor U6034 (N_6034,N_4066,N_5580);
and U6035 (N_6035,N_5620,N_3571);
xor U6036 (N_6036,N_3552,N_4150);
nand U6037 (N_6037,N_5526,N_4761);
xor U6038 (N_6038,N_3506,N_3486);
nor U6039 (N_6039,N_4144,N_4438);
or U6040 (N_6040,N_4698,N_4295);
xnor U6041 (N_6041,N_4680,N_4118);
nand U6042 (N_6042,N_5695,N_5356);
and U6043 (N_6043,N_5980,N_3100);
xnor U6044 (N_6044,N_3489,N_4733);
nand U6045 (N_6045,N_3084,N_3186);
and U6046 (N_6046,N_4519,N_4233);
nand U6047 (N_6047,N_5929,N_5168);
or U6048 (N_6048,N_5908,N_5285);
or U6049 (N_6049,N_3395,N_4672);
or U6050 (N_6050,N_3007,N_3836);
nand U6051 (N_6051,N_4259,N_4175);
nor U6052 (N_6052,N_3668,N_3793);
nand U6053 (N_6053,N_3142,N_5702);
xnor U6054 (N_6054,N_4523,N_4385);
xor U6055 (N_6055,N_4835,N_5738);
nor U6056 (N_6056,N_5978,N_3901);
or U6057 (N_6057,N_5933,N_4514);
or U6058 (N_6058,N_4483,N_3752);
nand U6059 (N_6059,N_4967,N_4158);
and U6060 (N_6060,N_5107,N_3697);
nand U6061 (N_6061,N_5960,N_3895);
xnor U6062 (N_6062,N_3956,N_3298);
or U6063 (N_6063,N_3010,N_4466);
nand U6064 (N_6064,N_3365,N_5449);
nor U6065 (N_6065,N_5874,N_4422);
or U6066 (N_6066,N_5673,N_3200);
nor U6067 (N_6067,N_3382,N_3429);
and U6068 (N_6068,N_4719,N_5034);
xnor U6069 (N_6069,N_4740,N_3348);
nor U6070 (N_6070,N_3952,N_3314);
xnor U6071 (N_6071,N_5312,N_3999);
and U6072 (N_6072,N_3774,N_4319);
nand U6073 (N_6073,N_3137,N_3612);
and U6074 (N_6074,N_4349,N_5727);
xor U6075 (N_6075,N_3928,N_3768);
nor U6076 (N_6076,N_5201,N_5195);
nor U6077 (N_6077,N_5541,N_4802);
and U6078 (N_6078,N_4223,N_3068);
xnor U6079 (N_6079,N_3112,N_5257);
nor U6080 (N_6080,N_5077,N_3251);
xor U6081 (N_6081,N_3450,N_4591);
or U6082 (N_6082,N_3286,N_3110);
xor U6083 (N_6083,N_5684,N_4559);
nand U6084 (N_6084,N_5480,N_5968);
xor U6085 (N_6085,N_3115,N_3270);
and U6086 (N_6086,N_4992,N_4720);
nand U6087 (N_6087,N_4945,N_4928);
nor U6088 (N_6088,N_3215,N_4291);
nand U6089 (N_6089,N_4267,N_5639);
nand U6090 (N_6090,N_4944,N_3234);
nor U6091 (N_6091,N_4963,N_3476);
and U6092 (N_6092,N_3898,N_5887);
xnor U6093 (N_6093,N_5409,N_3811);
nor U6094 (N_6094,N_5872,N_4503);
or U6095 (N_6095,N_4244,N_5280);
xnor U6096 (N_6096,N_5004,N_3759);
nor U6097 (N_6097,N_3954,N_5850);
nor U6098 (N_6098,N_5764,N_5563);
or U6099 (N_6099,N_4728,N_5687);
or U6100 (N_6100,N_3977,N_3619);
xor U6101 (N_6101,N_3247,N_4722);
or U6102 (N_6102,N_3771,N_4762);
xor U6103 (N_6103,N_3767,N_3177);
or U6104 (N_6104,N_5050,N_3713);
xnor U6105 (N_6105,N_3704,N_3322);
or U6106 (N_6106,N_4297,N_4330);
nor U6107 (N_6107,N_4791,N_3248);
nor U6108 (N_6108,N_5425,N_5589);
nand U6109 (N_6109,N_4739,N_5058);
nand U6110 (N_6110,N_3568,N_4999);
nor U6111 (N_6111,N_4713,N_4235);
xnor U6112 (N_6112,N_4723,N_5760);
and U6113 (N_6113,N_5600,N_4557);
xnor U6114 (N_6114,N_4792,N_3710);
nand U6115 (N_6115,N_3970,N_4051);
nand U6116 (N_6116,N_3180,N_5860);
or U6117 (N_6117,N_3035,N_5609);
nor U6118 (N_6118,N_5650,N_4725);
or U6119 (N_6119,N_4902,N_4696);
and U6120 (N_6120,N_3955,N_3896);
or U6121 (N_6121,N_3030,N_4757);
xnor U6122 (N_6122,N_4987,N_4822);
and U6123 (N_6123,N_3468,N_5691);
nand U6124 (N_6124,N_4904,N_3449);
nor U6125 (N_6125,N_5694,N_4619);
nand U6126 (N_6126,N_4564,N_4601);
nand U6127 (N_6127,N_4727,N_4594);
and U6128 (N_6128,N_5642,N_4343);
nand U6129 (N_6129,N_3492,N_5259);
xnor U6130 (N_6130,N_5141,N_5538);
or U6131 (N_6131,N_4803,N_4638);
or U6132 (N_6132,N_3926,N_4229);
xnor U6133 (N_6133,N_3364,N_5818);
nand U6134 (N_6134,N_4833,N_3245);
or U6135 (N_6135,N_5410,N_5547);
nand U6136 (N_6136,N_5636,N_4002);
or U6137 (N_6137,N_3566,N_3516);
or U6138 (N_6138,N_5110,N_3338);
or U6139 (N_6139,N_4962,N_3812);
and U6140 (N_6140,N_4299,N_3995);
xor U6141 (N_6141,N_5357,N_4756);
and U6142 (N_6142,N_3602,N_5436);
nor U6143 (N_6143,N_3257,N_3734);
nor U6144 (N_6144,N_5767,N_4510);
and U6145 (N_6145,N_5721,N_3191);
or U6146 (N_6146,N_5975,N_4093);
xor U6147 (N_6147,N_4227,N_5385);
and U6148 (N_6148,N_4442,N_4394);
or U6149 (N_6149,N_4825,N_4921);
nor U6150 (N_6150,N_3949,N_4853);
xnor U6151 (N_6151,N_3343,N_3885);
nand U6152 (N_6152,N_4377,N_5641);
and U6153 (N_6153,N_4260,N_5535);
nand U6154 (N_6154,N_5696,N_4521);
and U6155 (N_6155,N_4481,N_5473);
nand U6156 (N_6156,N_5942,N_4841);
and U6157 (N_6157,N_4779,N_4480);
and U6158 (N_6158,N_3262,N_4540);
or U6159 (N_6159,N_5967,N_3665);
or U6160 (N_6160,N_5136,N_4750);
or U6161 (N_6161,N_4972,N_5174);
nand U6162 (N_6162,N_5607,N_5699);
nand U6163 (N_6163,N_3376,N_4817);
and U6164 (N_6164,N_5038,N_4073);
nor U6165 (N_6165,N_3466,N_5379);
nand U6166 (N_6166,N_3876,N_5742);
xnor U6167 (N_6167,N_4671,N_5194);
or U6168 (N_6168,N_5234,N_5082);
nand U6169 (N_6169,N_3854,N_5779);
nand U6170 (N_6170,N_3782,N_5307);
xnor U6171 (N_6171,N_5670,N_5640);
nor U6172 (N_6172,N_5878,N_5811);
and U6173 (N_6173,N_5730,N_3375);
and U6174 (N_6174,N_3608,N_4242);
or U6175 (N_6175,N_4501,N_3853);
nor U6176 (N_6176,N_5889,N_3523);
nand U6177 (N_6177,N_5121,N_5938);
nand U6178 (N_6178,N_4289,N_5111);
nor U6179 (N_6179,N_4606,N_4829);
xnor U6180 (N_6180,N_4149,N_3139);
xnor U6181 (N_6181,N_4212,N_5712);
nand U6182 (N_6182,N_3134,N_3138);
nand U6183 (N_6183,N_4771,N_3992);
or U6184 (N_6184,N_4101,N_3507);
nor U6185 (N_6185,N_3776,N_3047);
xnor U6186 (N_6186,N_5987,N_4169);
nand U6187 (N_6187,N_5891,N_3436);
nor U6188 (N_6188,N_3185,N_3118);
and U6189 (N_6189,N_3543,N_4133);
xor U6190 (N_6190,N_4855,N_4734);
nand U6191 (N_6191,N_5261,N_3501);
xnor U6192 (N_6192,N_5506,N_4443);
or U6193 (N_6193,N_3742,N_5070);
and U6194 (N_6194,N_5052,N_3260);
nand U6195 (N_6195,N_4243,N_5880);
nor U6196 (N_6196,N_3154,N_3554);
nor U6197 (N_6197,N_5296,N_5153);
and U6198 (N_6198,N_5635,N_4737);
or U6199 (N_6199,N_4917,N_4552);
nor U6200 (N_6200,N_5899,N_5163);
nor U6201 (N_6201,N_4524,N_3276);
xor U6202 (N_6202,N_3086,N_3421);
and U6203 (N_6203,N_4745,N_5983);
and U6204 (N_6204,N_5840,N_4359);
and U6205 (N_6205,N_4626,N_3760);
nand U6206 (N_6206,N_5821,N_5910);
or U6207 (N_6207,N_5315,N_5578);
nor U6208 (N_6208,N_4842,N_5715);
and U6209 (N_6209,N_3062,N_3743);
and U6210 (N_6210,N_5233,N_3336);
nand U6211 (N_6211,N_5800,N_4074);
xor U6212 (N_6212,N_5505,N_5970);
xnor U6213 (N_6213,N_3117,N_5842);
and U6214 (N_6214,N_5736,N_5906);
and U6215 (N_6215,N_3494,N_4020);
xnor U6216 (N_6216,N_3419,N_5515);
and U6217 (N_6217,N_4577,N_5355);
and U6218 (N_6218,N_5778,N_5043);
xnor U6219 (N_6219,N_3575,N_3269);
nand U6220 (N_6220,N_4136,N_5446);
or U6221 (N_6221,N_4382,N_3093);
nor U6222 (N_6222,N_4048,N_5180);
nor U6223 (N_6223,N_5301,N_4414);
xnor U6224 (N_6224,N_3477,N_4386);
nor U6225 (N_6225,N_3461,N_5722);
nand U6226 (N_6226,N_5713,N_5406);
nor U6227 (N_6227,N_5277,N_4971);
and U6228 (N_6228,N_3306,N_5901);
xnor U6229 (N_6229,N_5571,N_4449);
nand U6230 (N_6230,N_3726,N_3073);
nor U6231 (N_6231,N_4166,N_4079);
xnor U6232 (N_6232,N_4605,N_3667);
nor U6233 (N_6233,N_3018,N_5661);
or U6234 (N_6234,N_5788,N_4588);
xnor U6235 (N_6235,N_3266,N_5830);
nand U6236 (N_6236,N_5314,N_4274);
and U6237 (N_6237,N_3255,N_4189);
and U6238 (N_6238,N_5513,N_4590);
and U6239 (N_6239,N_5591,N_4256);
nor U6240 (N_6240,N_5400,N_3109);
nor U6241 (N_6241,N_4247,N_3039);
or U6242 (N_6242,N_3478,N_5187);
or U6243 (N_6243,N_5698,N_4946);
nor U6244 (N_6244,N_4840,N_4642);
nand U6245 (N_6245,N_5158,N_3106);
nor U6246 (N_6246,N_3405,N_3317);
or U6247 (N_6247,N_4758,N_5316);
or U6248 (N_6248,N_3606,N_3821);
and U6249 (N_6249,N_5371,N_3125);
nand U6250 (N_6250,N_5274,N_3379);
nand U6251 (N_6251,N_5834,N_4464);
or U6252 (N_6252,N_4883,N_3224);
xor U6253 (N_6253,N_3629,N_5304);
xor U6254 (N_6254,N_4773,N_3385);
xnor U6255 (N_6255,N_4535,N_5598);
nor U6256 (N_6256,N_5423,N_5318);
nor U6257 (N_6257,N_3409,N_5492);
xor U6258 (N_6258,N_4918,N_5593);
and U6259 (N_6259,N_4615,N_4024);
or U6260 (N_6260,N_4208,N_4860);
and U6261 (N_6261,N_5615,N_4789);
xor U6262 (N_6262,N_4864,N_5990);
and U6263 (N_6263,N_4203,N_4441);
nand U6264 (N_6264,N_5869,N_4106);
nand U6265 (N_6265,N_4954,N_5909);
and U6266 (N_6266,N_5300,N_3238);
or U6267 (N_6267,N_3529,N_3615);
nand U6268 (N_6268,N_5823,N_5440);
and U6269 (N_6269,N_3179,N_4652);
xnor U6270 (N_6270,N_5757,N_3809);
and U6271 (N_6271,N_5197,N_3691);
and U6272 (N_6272,N_3867,N_5054);
nor U6273 (N_6273,N_4681,N_4184);
nand U6274 (N_6274,N_4217,N_4978);
or U6275 (N_6275,N_5857,N_4703);
nor U6276 (N_6276,N_5498,N_3623);
nor U6277 (N_6277,N_4873,N_3864);
xnor U6278 (N_6278,N_5030,N_4811);
xnor U6279 (N_6279,N_4796,N_3387);
and U6280 (N_6280,N_3611,N_5617);
or U6281 (N_6281,N_5710,N_4950);
or U6282 (N_6282,N_4327,N_3886);
or U6283 (N_6283,N_5948,N_3786);
xor U6284 (N_6284,N_4931,N_4163);
nand U6285 (N_6285,N_4225,N_5585);
xnor U6286 (N_6286,N_5267,N_3880);
and U6287 (N_6287,N_5214,N_5922);
nor U6288 (N_6288,N_3806,N_4526);
and U6289 (N_6289,N_5572,N_3924);
xor U6290 (N_6290,N_4751,N_3750);
or U6291 (N_6291,N_5175,N_5483);
nand U6292 (N_6292,N_4455,N_4831);
nor U6293 (N_6293,N_5338,N_5130);
nand U6294 (N_6294,N_4286,N_5524);
xnor U6295 (N_6295,N_5555,N_5202);
nor U6296 (N_6296,N_3242,N_4354);
nor U6297 (N_6297,N_3301,N_5472);
nor U6298 (N_6298,N_3846,N_4539);
nor U6299 (N_6299,N_4387,N_5605);
nand U6300 (N_6300,N_4492,N_5391);
nor U6301 (N_6301,N_5051,N_4974);
nand U6302 (N_6302,N_5348,N_3295);
nor U6303 (N_6303,N_4272,N_5424);
or U6304 (N_6304,N_5218,N_5614);
nor U6305 (N_6305,N_4300,N_3646);
xor U6306 (N_6306,N_4092,N_5648);
and U6307 (N_6307,N_5069,N_4104);
and U6308 (N_6308,N_4870,N_3650);
nand U6309 (N_6309,N_5509,N_5795);
and U6310 (N_6310,N_4909,N_3881);
and U6311 (N_6311,N_3985,N_5140);
nor U6312 (N_6312,N_5705,N_3335);
nand U6313 (N_6313,N_5629,N_5005);
and U6314 (N_6314,N_5374,N_4744);
xnor U6315 (N_6315,N_3442,N_3899);
xnor U6316 (N_6316,N_4111,N_4391);
nor U6317 (N_6317,N_4040,N_3016);
nand U6318 (N_6318,N_3239,N_3531);
or U6319 (N_6319,N_4365,N_4576);
nand U6320 (N_6320,N_5903,N_4957);
and U6321 (N_6321,N_3280,N_5522);
xnor U6322 (N_6322,N_3290,N_3254);
or U6323 (N_6323,N_4311,N_3856);
nor U6324 (N_6324,N_3350,N_5588);
nand U6325 (N_6325,N_5819,N_3916);
nor U6326 (N_6326,N_5667,N_4029);
or U6327 (N_6327,N_5561,N_3085);
nand U6328 (N_6328,N_4433,N_5323);
nor U6329 (N_6329,N_3017,N_3647);
and U6330 (N_6330,N_4821,N_4643);
xor U6331 (N_6331,N_5086,N_4699);
xnor U6332 (N_6332,N_5414,N_4436);
xnor U6333 (N_6333,N_3683,N_5476);
nand U6334 (N_6334,N_3528,N_4923);
xor U6335 (N_6335,N_5709,N_3712);
or U6336 (N_6336,N_4255,N_5965);
nand U6337 (N_6337,N_4325,N_4228);
nand U6338 (N_6338,N_4419,N_3435);
nor U6339 (N_6339,N_5403,N_5637);
xnor U6340 (N_6340,N_3252,N_4746);
or U6341 (N_6341,N_4198,N_5991);
nor U6342 (N_6342,N_3320,N_4383);
or U6343 (N_6343,N_4583,N_3063);
nand U6344 (N_6344,N_4350,N_4905);
or U6345 (N_6345,N_3192,N_3340);
or U6346 (N_6346,N_5949,N_5003);
xor U6347 (N_6347,N_5943,N_4669);
nand U6348 (N_6348,N_3563,N_3043);
nand U6349 (N_6349,N_5962,N_5036);
xor U6350 (N_6350,N_3493,N_3099);
and U6351 (N_6351,N_3512,N_3082);
and U6352 (N_6352,N_4099,N_4213);
nand U6353 (N_6353,N_4209,N_4096);
nor U6354 (N_6354,N_3631,N_5162);
nand U6355 (N_6355,N_4961,N_5604);
and U6356 (N_6356,N_5241,N_5870);
or U6357 (N_6357,N_5809,N_5311);
nor U6358 (N_6358,N_4710,N_3877);
nor U6359 (N_6359,N_5227,N_4375);
xnor U6360 (N_6360,N_4834,N_4780);
nand U6361 (N_6361,N_5359,N_3076);
xnor U6362 (N_6362,N_5010,N_5981);
xnor U6363 (N_6363,N_5876,N_5115);
and U6364 (N_6364,N_3300,N_4566);
nor U6365 (N_6365,N_5279,N_3979);
and U6366 (N_6366,N_5595,N_5184);
nand U6367 (N_6367,N_4875,N_4384);
and U6368 (N_6368,N_3406,N_5366);
nand U6369 (N_6369,N_4714,N_4660);
or U6370 (N_6370,N_3678,N_4986);
and U6371 (N_6371,N_3469,N_4997);
xnor U6372 (N_6372,N_5254,N_5930);
nor U6373 (N_6373,N_5724,N_5845);
nand U6374 (N_6374,N_5014,N_4795);
and U6375 (N_6375,N_4425,N_4673);
and U6376 (N_6376,N_3441,N_4505);
xor U6377 (N_6377,N_5408,N_3324);
xor U6378 (N_6378,N_5185,N_3538);
nor U6379 (N_6379,N_3588,N_4207);
xor U6380 (N_6380,N_3232,N_5758);
xor U6381 (N_6381,N_3176,N_4257);
or U6382 (N_6382,N_5507,N_4115);
nand U6383 (N_6383,N_4323,N_5065);
or U6384 (N_6384,N_3887,N_3859);
or U6385 (N_6385,N_4537,N_4078);
and U6386 (N_6386,N_3371,N_5288);
nor U6387 (N_6387,N_3359,N_3948);
nand U6388 (N_6388,N_3488,N_3246);
nand U6389 (N_6389,N_3312,N_5131);
xor U6390 (N_6390,N_4121,N_4194);
or U6391 (N_6391,N_3508,N_4894);
xnor U6392 (N_6392,N_4326,N_4684);
xor U6393 (N_6393,N_4258,N_3598);
nor U6394 (N_6394,N_3637,N_3624);
nand U6395 (N_6395,N_3694,N_3869);
or U6396 (N_6396,N_4312,N_3504);
nand U6397 (N_6397,N_5810,N_5389);
xor U6398 (N_6398,N_3475,N_5461);
and U6399 (N_6399,N_4388,N_5203);
and U6400 (N_6400,N_4374,N_5468);
nand U6401 (N_6401,N_3780,N_5192);
nor U6402 (N_6402,N_3613,N_4340);
nand U6403 (N_6403,N_5861,N_4743);
or U6404 (N_6404,N_4711,N_5717);
xor U6405 (N_6405,N_4649,N_5404);
xnor U6406 (N_6406,N_5019,N_3594);
and U6407 (N_6407,N_3959,N_4276);
xnor U6408 (N_6408,N_5208,N_5791);
nor U6409 (N_6409,N_4161,N_3513);
nand U6410 (N_6410,N_5766,N_5976);
xor U6411 (N_6411,N_4494,N_5139);
xnor U6412 (N_6412,N_5841,N_3119);
nand U6413 (N_6413,N_3349,N_3041);
xor U6414 (N_6414,N_4117,N_5049);
nor U6415 (N_6415,N_3431,N_5856);
xnor U6416 (N_6416,N_3820,N_5294);
nand U6417 (N_6417,N_5033,N_5848);
and U6418 (N_6418,N_3527,N_3929);
nor U6419 (N_6419,N_4434,N_5450);
or U6420 (N_6420,N_5319,N_5675);
or U6421 (N_6421,N_5776,N_5682);
nor U6422 (N_6422,N_3014,N_3582);
nand U6423 (N_6423,N_4181,N_4620);
xnor U6424 (N_6424,N_3840,N_4416);
nor U6425 (N_6425,N_5740,N_5807);
xnor U6426 (N_6426,N_3465,N_4690);
and U6427 (N_6427,N_5814,N_3194);
nor U6428 (N_6428,N_5630,N_3454);
or U6429 (N_6429,N_4645,N_3445);
nor U6430 (N_6430,N_5542,N_5146);
nand U6431 (N_6431,N_4333,N_3763);
nand U6432 (N_6432,N_4609,N_5243);
and U6433 (N_6433,N_3092,N_5060);
and U6434 (N_6434,N_3794,N_3236);
xnor U6435 (N_6435,N_4955,N_5240);
or U6436 (N_6436,N_5616,N_5027);
xor U6437 (N_6437,N_5466,N_3221);
nor U6438 (N_6438,N_3590,N_5517);
nand U6439 (N_6439,N_5100,N_4336);
or U6440 (N_6440,N_4162,N_3370);
nand U6441 (N_6441,N_3751,N_4785);
and U6442 (N_6442,N_3744,N_5351);
and U6443 (N_6443,N_4232,N_4774);
nor U6444 (N_6444,N_3762,N_5704);
nand U6445 (N_6445,N_4580,N_5774);
and U6446 (N_6446,N_4482,N_3622);
nor U6447 (N_6447,N_4065,N_4995);
nand U6448 (N_6448,N_3577,N_5612);
or U6449 (N_6449,N_4741,N_3603);
or U6450 (N_6450,N_5752,N_4731);
nand U6451 (N_6451,N_4653,N_4630);
or U6452 (N_6452,N_5292,N_5448);
nor U6453 (N_6453,N_3366,N_3277);
or U6454 (N_6454,N_3748,N_3243);
or U6455 (N_6455,N_5432,N_3229);
and U6456 (N_6456,N_3964,N_4689);
or U6457 (N_6457,N_4807,N_4472);
or U6458 (N_6458,N_3329,N_5482);
or U6459 (N_6459,N_4406,N_3573);
and U6460 (N_6460,N_3651,N_5134);
and U6461 (N_6461,N_4216,N_4520);
and U6462 (N_6462,N_5370,N_5502);
and U6463 (N_6463,N_4427,N_3167);
nand U6464 (N_6464,N_3211,N_4246);
xnor U6465 (N_6465,N_4898,N_3635);
nand U6466 (N_6466,N_5006,N_3173);
or U6467 (N_6467,N_4554,N_5282);
or U6468 (N_6468,N_5714,N_5112);
nor U6469 (N_6469,N_4663,N_4471);
or U6470 (N_6470,N_4567,N_4876);
xnor U6471 (N_6471,N_4279,N_4052);
xor U6472 (N_6472,N_5944,N_3111);
and U6473 (N_6473,N_4888,N_5677);
or U6474 (N_6474,N_5781,N_3196);
nand U6475 (N_6475,N_3005,N_3911);
and U6476 (N_6476,N_3330,N_4852);
nor U6477 (N_6477,N_4417,N_4534);
nand U6478 (N_6478,N_3988,N_3618);
nand U6479 (N_6479,N_4125,N_5171);
nor U6480 (N_6480,N_3968,N_5854);
xor U6481 (N_6481,N_5905,N_3599);
and U6482 (N_6482,N_4597,N_5177);
nor U6483 (N_6483,N_5592,N_3932);
and U6484 (N_6484,N_4625,N_3264);
xor U6485 (N_6485,N_3534,N_4462);
xor U6486 (N_6486,N_5864,N_5737);
nand U6487 (N_6487,N_5388,N_4160);
xor U6488 (N_6488,N_3593,N_5678);
or U6489 (N_6489,N_4315,N_5128);
xnor U6490 (N_6490,N_5665,N_4805);
xor U6491 (N_6491,N_3051,N_5386);
xor U6492 (N_6492,N_5354,N_4430);
nor U6493 (N_6493,N_5471,N_5836);
or U6494 (N_6494,N_5418,N_4584);
nor U6495 (N_6495,N_4799,N_3747);
xor U6496 (N_6496,N_3228,N_3957);
nand U6497 (N_6497,N_5299,N_4265);
nor U6498 (N_6498,N_4879,N_3075);
and U6499 (N_6499,N_5289,N_3787);
nor U6500 (N_6500,N_4236,N_3866);
nand U6501 (N_6501,N_4054,N_3060);
nor U6502 (N_6502,N_3050,N_5368);
nor U6503 (N_6503,N_3672,N_5120);
or U6504 (N_6504,N_5215,N_4485);
nor U6505 (N_6505,N_5516,N_4362);
or U6506 (N_6506,N_4479,N_5377);
and U6507 (N_6507,N_4116,N_3059);
and U6508 (N_6508,N_3273,N_3556);
nor U6509 (N_6509,N_5164,N_5264);
xor U6510 (N_6510,N_4983,N_4061);
xor U6511 (N_6511,N_3907,N_3023);
nand U6512 (N_6512,N_4013,N_4709);
or U6513 (N_6513,N_5701,N_4516);
nor U6514 (N_6514,N_4041,N_5963);
nand U6515 (N_6515,N_4358,N_5884);
nor U6516 (N_6516,N_3914,N_3855);
and U6517 (N_6517,N_5902,N_3391);
nor U6518 (N_6518,N_5759,N_4662);
nand U6519 (N_6519,N_3249,N_3116);
nand U6520 (N_6520,N_4551,N_5108);
xnor U6521 (N_6521,N_3164,N_5305);
or U6522 (N_6522,N_4753,N_5925);
nor U6523 (N_6523,N_5117,N_5888);
or U6524 (N_6524,N_4623,N_4185);
and U6525 (N_6525,N_3827,N_3567);
nand U6526 (N_6526,N_3161,N_5647);
and U6527 (N_6527,N_4555,N_3605);
xor U6528 (N_6528,N_5161,N_4527);
nor U6529 (N_6529,N_4976,N_5999);
nor U6530 (N_6530,N_4344,N_4199);
xor U6531 (N_6531,N_3019,N_3562);
or U6532 (N_6532,N_4657,N_3189);
or U6533 (N_6533,N_4887,N_5594);
nand U6534 (N_6534,N_4129,N_5831);
and U6535 (N_6535,N_5055,N_4668);
nand U6536 (N_6536,N_4956,N_3656);
or U6537 (N_6537,N_4230,N_4907);
nor U6538 (N_6538,N_4655,N_4607);
nand U6539 (N_6539,N_4778,N_4515);
xor U6540 (N_6540,N_3334,N_3497);
or U6541 (N_6541,N_5559,N_3231);
nor U6542 (N_6542,N_3716,N_5336);
nor U6543 (N_6543,N_3700,N_3345);
nand U6544 (N_6544,N_5835,N_5602);
xnor U6545 (N_6545,N_4282,N_3020);
and U6546 (N_6546,N_3772,N_5936);
and U6547 (N_6547,N_3094,N_4105);
nor U6548 (N_6548,N_4793,N_5654);
nand U6549 (N_6549,N_5923,N_3717);
xor U6550 (N_6550,N_4575,N_4084);
xor U6551 (N_6551,N_5302,N_3945);
or U6552 (N_6552,N_4820,N_3352);
nor U6553 (N_6553,N_3408,N_5839);
and U6554 (N_6554,N_5283,N_3845);
or U6555 (N_6555,N_4068,N_5534);
and U6556 (N_6556,N_5504,N_5995);
xor U6557 (N_6557,N_4355,N_5935);
xnor U6558 (N_6558,N_5690,N_5228);
xnor U6559 (N_6559,N_4476,N_3660);
nand U6560 (N_6560,N_5478,N_3218);
xnor U6561 (N_6561,N_3514,N_3775);
xor U6562 (N_6562,N_3576,N_4431);
nand U6563 (N_6563,N_3052,N_4882);
xor U6564 (N_6564,N_5383,N_5753);
nor U6565 (N_6565,N_5587,N_4755);
or U6566 (N_6566,N_5871,N_3058);
and U6567 (N_6567,N_4599,N_5239);
and U6568 (N_6568,N_3626,N_5806);
or U6569 (N_6569,N_3146,N_3559);
and U6570 (N_6570,N_4808,N_5080);
and U6571 (N_6571,N_3833,N_4919);
nor U6572 (N_6572,N_4893,N_5531);
or U6573 (N_6573,N_4990,N_3415);
nor U6574 (N_6574,N_3294,N_3947);
or U6575 (N_6575,N_4528,N_5734);
xnor U6576 (N_6576,N_4646,N_5022);
nand U6577 (N_6577,N_3511,N_4191);
nand U6578 (N_6578,N_3396,N_5552);
nand U6579 (N_6579,N_4484,N_3484);
nor U6580 (N_6580,N_3399,N_3162);
nor U6581 (N_6581,N_3682,N_4670);
xnor U6582 (N_6582,N_4083,N_4317);
or U6583 (N_6583,N_5532,N_3757);
nor U6584 (N_6584,N_4342,N_5493);
xor U6585 (N_6585,N_4592,N_3012);
nor U6586 (N_6586,N_5570,N_5392);
or U6587 (N_6587,N_3299,N_4784);
or U6588 (N_6588,N_5102,N_4953);
nor U6589 (N_6589,N_5335,N_4459);
xnor U6590 (N_6590,N_5953,N_4939);
nor U6591 (N_6591,N_4263,N_4221);
nor U6592 (N_6592,N_5456,N_3908);
xnor U6593 (N_6593,N_4183,N_4049);
and U6594 (N_6594,N_3532,N_4428);
nor U6595 (N_6595,N_5295,N_3487);
nor U6596 (N_6596,N_4007,N_5907);
nor U6597 (N_6597,N_3526,N_5001);
xnor U6598 (N_6598,N_5892,N_4975);
or U6599 (N_6599,N_3420,N_4752);
xor U6600 (N_6600,N_3939,N_5969);
nand U6601 (N_6601,N_4461,N_4448);
nor U6602 (N_6602,N_5275,N_4991);
nand U6603 (N_6603,N_4826,N_3288);
nor U6604 (N_6604,N_5863,N_5401);
and U6605 (N_6605,N_3363,N_5852);
and U6606 (N_6606,N_3578,N_3381);
xnor U6607 (N_6607,N_5276,N_3510);
nor U6608 (N_6608,N_5166,N_4866);
nand U6609 (N_6609,N_5007,N_4122);
and U6610 (N_6610,N_3090,N_3392);
or U6611 (N_6611,N_5268,N_3356);
xnor U6612 (N_6612,N_3936,N_4716);
nand U6613 (N_6613,N_5236,N_5618);
or U6614 (N_6614,N_5674,N_5873);
and U6615 (N_6615,N_5927,N_3858);
nand U6616 (N_6616,N_5365,N_5653);
nand U6617 (N_6617,N_3861,N_4574);
nand U6618 (N_6618,N_4872,N_5106);
nand U6619 (N_6619,N_3457,N_4827);
and U6620 (N_6620,N_3166,N_5959);
and U6621 (N_6621,N_4691,N_3781);
and U6622 (N_6622,N_4878,N_5947);
nor U6623 (N_6623,N_5745,N_3437);
xnor U6624 (N_6624,N_5769,N_4968);
or U6625 (N_6625,N_4563,N_3297);
xor U6626 (N_6626,N_4451,N_3986);
or U6627 (N_6627,N_4318,N_3580);
xnor U6628 (N_6628,N_5971,N_4287);
and U6629 (N_6629,N_5105,N_3798);
and U6630 (N_6630,N_3265,N_3460);
nand U6631 (N_6631,N_4846,N_3223);
or U6632 (N_6632,N_5340,N_4542);
or U6633 (N_6633,N_5692,N_5877);
and U6634 (N_6634,N_4298,N_5364);
nand U6635 (N_6635,N_4786,N_3805);
or U6636 (N_6636,N_3940,N_4429);
nand U6637 (N_6637,N_3158,N_5361);
nand U6638 (N_6638,N_4151,N_3407);
nor U6639 (N_6639,N_3558,N_3434);
and U6640 (N_6640,N_3098,N_5083);
nand U6641 (N_6641,N_5039,N_5985);
and U6642 (N_6642,N_3944,N_3912);
xor U6643 (N_6643,N_5394,N_4487);
xnor U6644 (N_6644,N_4969,N_4307);
and U6645 (N_6645,N_5415,N_4393);
nand U6646 (N_6646,N_3551,N_5142);
nor U6647 (N_6647,N_3730,N_4338);
xnor U6648 (N_6648,N_4139,N_4610);
xnor U6649 (N_6649,N_4214,N_3692);
nand U6650 (N_6650,N_3498,N_5633);
and U6651 (N_6651,N_4794,N_5875);
and U6652 (N_6652,N_3097,N_4403);
and U6653 (N_6653,N_3208,N_4765);
nor U6654 (N_6654,N_3910,N_5726);
or U6655 (N_6655,N_5544,N_4390);
or U6656 (N_6656,N_5501,N_3789);
nor U6657 (N_6657,N_5660,N_4392);
nor U6658 (N_6658,N_5244,N_5265);
nand U6659 (N_6659,N_3709,N_5567);
and U6660 (N_6660,N_3801,N_5896);
nor U6661 (N_6661,N_4172,N_4844);
or U6662 (N_6662,N_5475,N_5116);
xnor U6663 (N_6663,N_4767,N_3021);
or U6664 (N_6664,N_5209,N_5237);
xnor U6665 (N_6665,N_4581,N_5095);
or U6666 (N_6666,N_3817,N_5123);
nand U6667 (N_6667,N_3394,N_5281);
or U6668 (N_6668,N_5979,N_5762);
nand U6669 (N_6669,N_3384,N_4131);
and U6670 (N_6670,N_5763,N_3641);
or U6671 (N_6671,N_5148,N_3796);
nand U6672 (N_6672,N_5287,N_4254);
or U6673 (N_6673,N_5984,N_5242);
nand U6674 (N_6674,N_4130,N_3152);
or U6675 (N_6675,N_3733,N_5865);
nand U6676 (N_6676,N_5645,N_4748);
nor U6677 (N_6677,N_4200,N_3272);
and U6678 (N_6678,N_3416,N_5619);
xor U6679 (N_6679,N_5632,N_4364);
xnor U6680 (N_6680,N_4869,N_3184);
or U6681 (N_6681,N_3874,N_3969);
nand U6682 (N_6682,N_3398,N_5467);
and U6683 (N_6683,N_5255,N_5780);
or U6684 (N_6684,N_4371,N_4290);
and U6685 (N_6685,N_4964,N_4556);
nand U6686 (N_6686,N_5145,N_5113);
and U6687 (N_6687,N_5231,N_3378);
nor U6688 (N_6688,N_3155,N_4418);
or U6689 (N_6689,N_5453,N_5331);
nor U6690 (N_6690,N_5460,N_4148);
and U6691 (N_6691,N_3207,N_3346);
nor U6692 (N_6692,N_3711,N_4334);
or U6693 (N_6693,N_5119,N_4749);
nand U6694 (N_6694,N_4863,N_3105);
nand U6695 (N_6695,N_3024,N_3731);
nand U6696 (N_6696,N_3706,N_5367);
xnor U6697 (N_6697,N_5178,N_4376);
nor U6698 (N_6698,N_3621,N_3707);
and U6699 (N_6699,N_5804,N_4569);
nand U6700 (N_6700,N_5939,N_3669);
nor U6701 (N_6701,N_5099,N_4628);
or U6702 (N_6702,N_5576,N_5973);
and U6703 (N_6703,N_3686,N_4446);
or U6704 (N_6704,N_5062,N_4174);
nand U6705 (N_6705,N_5782,N_4324);
or U6706 (N_6706,N_4050,N_3347);
and U6707 (N_6707,N_4294,N_3337);
nand U6708 (N_6708,N_4814,N_4706);
and U6709 (N_6709,N_4192,N_5372);
and U6710 (N_6710,N_4621,N_4123);
and U6711 (N_6711,N_5230,N_5805);
and U6712 (N_6712,N_4941,N_4182);
and U6713 (N_6713,N_5041,N_5373);
xnor U6714 (N_6714,N_5672,N_3729);
and U6715 (N_6715,N_5376,N_3057);
or U6716 (N_6716,N_4292,N_3261);
xor U6717 (N_6717,N_4637,N_5773);
xnor U6718 (N_6718,N_3813,N_3841);
nor U6719 (N_6719,N_5459,N_3857);
and U6720 (N_6720,N_5622,N_4650);
nor U6721 (N_6721,N_5219,N_4372);
and U6722 (N_6722,N_3104,N_5829);
and U6723 (N_6723,N_3323,N_5345);
or U6724 (N_6724,N_5545,N_3927);
nor U6725 (N_6725,N_4124,N_3333);
nor U6726 (N_6726,N_5838,N_5510);
and U6727 (N_6727,N_5008,N_3963);
xnor U6728 (N_6728,N_3696,N_4560);
nand U6729 (N_6729,N_3203,N_3727);
xnor U6730 (N_6730,N_3909,N_4145);
and U6731 (N_6731,N_3547,N_3077);
and U6732 (N_6732,N_3915,N_5439);
nand U6733 (N_6733,N_3193,N_3026);
or U6734 (N_6734,N_5813,N_4220);
and U6735 (N_6735,N_5462,N_3042);
nand U6736 (N_6736,N_5347,N_5756);
nand U6737 (N_6737,N_4687,N_5352);
and U6738 (N_6738,N_3745,N_4090);
xor U6739 (N_6739,N_4369,N_5611);
xor U6740 (N_6740,N_3755,N_5610);
nand U6741 (N_6741,N_4100,N_3883);
and U6742 (N_6742,N_3636,N_4231);
and U6743 (N_6743,N_3009,N_5771);
nor U6744 (N_6744,N_5042,N_5138);
nand U6745 (N_6745,N_4211,N_5103);
nand U6746 (N_6746,N_4631,N_3803);
xor U6747 (N_6747,N_4988,N_4395);
and U6748 (N_6748,N_5081,N_4586);
and U6749 (N_6749,N_5741,N_5579);
nand U6750 (N_6750,N_3209,N_4009);
and U6751 (N_6751,N_3481,N_4399);
nor U6752 (N_6752,N_5085,N_5437);
nand U6753 (N_6753,N_4037,N_5308);
nor U6754 (N_6754,N_4469,N_3289);
xor U6755 (N_6755,N_4465,N_5429);
nand U6756 (N_6756,N_4088,N_5998);
nand U6757 (N_6757,N_4304,N_4787);
and U6758 (N_6758,N_4460,N_3373);
and U6759 (N_6759,N_4708,N_4134);
nand U6760 (N_6760,N_4110,N_3275);
nand U6761 (N_6761,N_3975,N_5390);
nand U6762 (N_6762,N_3027,N_4913);
xor U6763 (N_6763,N_4156,N_3604);
nand U6764 (N_6764,N_4940,N_4138);
nand U6765 (N_6765,N_4943,N_4611);
nand U6766 (N_6766,N_4960,N_3591);
or U6767 (N_6767,N_3482,N_4022);
xor U6768 (N_6768,N_5735,N_3546);
and U6769 (N_6769,N_3227,N_3123);
or U6770 (N_6770,N_5057,N_5431);
nor U6771 (N_6771,N_3816,N_5247);
or U6772 (N_6772,N_3735,N_4187);
xnor U6773 (N_6773,N_5056,N_3509);
xnor U6774 (N_6774,N_3171,N_4823);
and U6775 (N_6775,N_5317,N_4015);
nand U6776 (N_6776,N_5853,N_3088);
nor U6777 (N_6777,N_3432,N_5603);
and U6778 (N_6778,N_4202,N_3617);
and U6779 (N_6779,N_5298,N_4296);
and U6780 (N_6780,N_4458,N_3046);
or U6781 (N_6781,N_3736,N_3217);
xnor U6782 (N_6782,N_3520,N_5744);
xnor U6783 (N_6783,N_3502,N_4253);
nor U6784 (N_6784,N_4573,N_4153);
and U6785 (N_6785,N_3982,N_3518);
nand U6786 (N_6786,N_3922,N_3135);
nand U6787 (N_6787,N_3754,N_4966);
nor U6788 (N_6788,N_5271,N_4306);
and U6789 (N_6789,N_5601,N_4411);
xnor U6790 (N_6790,N_5866,N_4081);
xor U6791 (N_6791,N_5796,N_3430);
or U6792 (N_6792,N_5329,N_5344);
xnor U6793 (N_6793,N_3721,N_3723);
xor U6794 (N_6794,N_5911,N_4568);
or U6795 (N_6795,N_3607,N_3640);
nor U6796 (N_6796,N_3868,N_3412);
nor U6797 (N_6797,N_3632,N_5822);
nand U6798 (N_6798,N_5586,N_3078);
xor U6799 (N_6799,N_4686,N_5723);
and U6800 (N_6800,N_5560,N_3136);
and U6801 (N_6801,N_3553,N_4782);
nand U6802 (N_6802,N_4204,N_4721);
nand U6803 (N_6803,N_3674,N_5118);
and U6804 (N_6804,N_4618,N_4381);
or U6805 (N_6805,N_3971,N_3839);
xor U6806 (N_6806,N_3521,N_3807);
or U6807 (N_6807,N_3875,N_3783);
or U6808 (N_6808,N_5519,N_5179);
or U6809 (N_6809,N_3006,N_4280);
nor U6810 (N_6810,N_3779,N_3725);
and U6811 (N_6811,N_5172,N_3560);
xor U6812 (N_6812,N_5897,N_5837);
nor U6813 (N_6813,N_3595,N_4178);
and U6814 (N_6814,N_3600,N_4032);
nand U6815 (N_6815,N_3339,N_4884);
nor U6816 (N_6816,N_5225,N_3225);
xor U6817 (N_6817,N_3377,N_3074);
and U6818 (N_6818,N_3677,N_5728);
xor U6819 (N_6819,N_4437,N_4128);
nand U6820 (N_6820,N_4109,N_5920);
nand U6821 (N_6821,N_5855,N_5787);
and U6822 (N_6822,N_3648,N_4938);
and U6823 (N_6823,N_5235,N_5679);
xnor U6824 (N_6824,N_4571,N_4781);
xnor U6825 (N_6825,N_5032,N_4850);
nor U6826 (N_6826,N_5982,N_4353);
nand U6827 (N_6827,N_4404,N_3067);
xor U6828 (N_6828,N_5253,N_5749);
nand U6829 (N_6829,N_4911,N_4847);
nand U6830 (N_6830,N_3401,N_5369);
xor U6831 (N_6831,N_3525,N_3756);
nand U6832 (N_6832,N_4018,N_5224);
nor U6833 (N_6833,N_5992,N_3541);
xor U6834 (N_6834,N_5291,N_3069);
nor U6835 (N_6835,N_3888,N_4874);
nor U6836 (N_6836,N_3549,N_5026);
nor U6837 (N_6837,N_4475,N_3291);
nand U6838 (N_6838,N_3654,N_3095);
nand U6839 (N_6839,N_3284,N_3778);
xor U6840 (N_6840,N_5293,N_3427);
nor U6841 (N_6841,N_3860,N_5977);
or U6842 (N_6842,N_3950,N_5489);
and U6843 (N_6843,N_4454,N_4837);
and U6844 (N_6844,N_3202,N_4768);
nand U6845 (N_6845,N_5859,N_3358);
nor U6846 (N_6846,N_3351,N_3183);
or U6847 (N_6847,N_5303,N_4903);
nand U6848 (N_6848,N_4705,N_4730);
xor U6849 (N_6849,N_5708,N_3851);
nor U6850 (N_6850,N_3372,N_3244);
and U6851 (N_6851,N_3749,N_5511);
xor U6852 (N_6852,N_5849,N_3362);
xor U6853 (N_6853,N_4447,N_4858);
or U6854 (N_6854,N_4634,N_4026);
or U6855 (N_6855,N_3921,N_4815);
xor U6856 (N_6856,N_4797,N_4838);
and U6857 (N_6857,N_5720,N_5941);
xnor U6858 (N_6858,N_4360,N_3080);
and U6859 (N_6859,N_3681,N_5387);
and U6860 (N_6860,N_4320,N_3884);
and U6861 (N_6861,N_3285,N_4132);
and U6862 (N_6862,N_4589,N_3539);
nor U6863 (N_6863,N_5739,N_5216);
xnor U6864 (N_6864,N_5820,N_3832);
nand U6865 (N_6865,N_4284,N_4937);
or U6866 (N_6866,N_4547,N_5067);
nand U6867 (N_6867,N_3129,N_4219);
xor U6868 (N_6868,N_4329,N_3800);
xor U6869 (N_6869,N_4729,N_4868);
or U6870 (N_6870,N_3662,N_3838);
or U6871 (N_6871,N_3746,N_3585);
nand U6872 (N_6872,N_3182,N_3096);
or U6873 (N_6873,N_3467,N_3271);
or U6874 (N_6874,N_3474,N_4980);
or U6875 (N_6875,N_5101,N_4249);
and U6876 (N_6876,N_4570,N_4097);
nor U6877 (N_6877,N_4989,N_4763);
nand U6878 (N_6878,N_4656,N_3263);
nand U6879 (N_6879,N_3989,N_4828);
and U6880 (N_6880,N_4511,N_4608);
and U6881 (N_6881,N_5064,N_5416);
xor U6882 (N_6882,N_3542,N_5490);
nand U6883 (N_6883,N_5321,N_4622);
or U6884 (N_6884,N_4165,N_3972);
and U6885 (N_6885,N_3175,N_3601);
and U6886 (N_6886,N_4977,N_5210);
nor U6887 (N_6887,N_3657,N_4337);
or U6888 (N_6888,N_3149,N_4210);
nor U6889 (N_6889,N_4936,N_3879);
and U6890 (N_6890,N_4558,N_4091);
nor U6891 (N_6891,N_5137,N_4985);
xor U6892 (N_6892,N_3850,N_4085);
nand U6893 (N_6893,N_3443,N_3680);
xor U6894 (N_6894,N_5613,N_4738);
nand U6895 (N_6895,N_5912,N_4627);
nand U6896 (N_6896,N_4309,N_4405);
nand U6897 (N_6897,N_3418,N_3688);
xor U6898 (N_6898,N_4867,N_5183);
nand U6899 (N_6899,N_5144,N_4266);
xnor U6900 (N_6900,N_3628,N_3967);
nand U6901 (N_6901,N_5790,N_3831);
or U6902 (N_6902,N_3458,N_4979);
and U6903 (N_6903,N_5754,N_5226);
or U6904 (N_6904,N_3645,N_4766);
xnor U6905 (N_6905,N_5358,N_4341);
xnor U6906 (N_6906,N_4470,N_5427);
nor U6907 (N_6907,N_3837,N_3714);
or U6908 (N_6908,N_5824,N_3535);
and U6909 (N_6909,N_3653,N_3784);
nor U6910 (N_6910,N_5258,N_5914);
or U6911 (N_6911,N_3108,N_5797);
nand U6912 (N_6912,N_3897,N_5434);
or U6913 (N_6913,N_4926,N_4444);
xor U6914 (N_6914,N_3383,N_5273);
nand U6915 (N_6915,N_3819,N_5955);
nor U6916 (N_6916,N_5508,N_5706);
nor U6917 (N_6917,N_3033,N_4424);
xnor U6918 (N_6918,N_5212,N_4504);
and U6919 (N_6919,N_3011,N_5700);
nand U6920 (N_6920,N_4572,N_4532);
nor U6921 (N_6921,N_3483,N_5339);
nor U6922 (N_6922,N_3132,N_4193);
and U6923 (N_6923,N_4335,N_5537);
nor U6924 (N_6924,N_5190,N_4102);
xor U6925 (N_6925,N_5309,N_5825);
nand U6926 (N_6926,N_4043,N_5495);
xor U6927 (N_6927,N_4270,N_3400);
xnor U6928 (N_6928,N_4545,N_3655);
and U6929 (N_6929,N_3279,N_4973);
nand U6930 (N_6930,N_4019,N_5816);
or U6931 (N_6931,N_3946,N_4409);
xor U6932 (N_6932,N_3587,N_5104);
nand U6933 (N_6933,N_3089,N_5808);
and U6934 (N_6934,N_5514,N_4701);
or U6935 (N_6935,N_5332,N_4450);
nor U6936 (N_6936,N_5703,N_3823);
nand U6937 (N_6937,N_4474,N_3825);
or U6938 (N_6938,N_4076,N_4113);
nand U6939 (N_6939,N_3524,N_3169);
nor U6940 (N_6940,N_4396,N_5091);
or U6941 (N_6941,N_5313,N_3331);
xnor U6942 (N_6942,N_4717,N_3414);
nor U6943 (N_6943,N_5658,N_5890);
nand U6944 (N_6944,N_3361,N_5442);
xnor U6945 (N_6945,N_5550,N_5380);
or U6946 (N_6946,N_3739,N_3679);
nand U6947 (N_6947,N_4927,N_4432);
or U6948 (N_6948,N_5075,N_3670);
and U6949 (N_6949,N_3505,N_5919);
or U6950 (N_6950,N_4251,N_5958);
nand U6951 (N_6951,N_3519,N_5223);
and U6952 (N_6952,N_3165,N_3367);
xor U6953 (N_6953,N_4788,N_3942);
nand U6954 (N_6954,N_3127,N_4331);
nor U6955 (N_6955,N_4321,N_5479);
nor U6956 (N_6956,N_5792,N_3906);
and U6957 (N_6957,N_5523,N_4612);
nor U6958 (N_6958,N_3732,N_3205);
xor U6959 (N_6959,N_3045,N_4435);
nand U6960 (N_6960,N_5827,N_5229);
or U6961 (N_6961,N_4154,N_5031);
xor U6962 (N_6962,N_4982,N_5263);
nor U6963 (N_6963,N_3943,N_4142);
or U6964 (N_6964,N_4303,N_5046);
xnor U6965 (N_6965,N_4170,N_5147);
xnor U6966 (N_6966,N_5017,N_3274);
and U6967 (N_6967,N_4886,N_5306);
xor U6968 (N_6968,N_5152,N_4277);
or U6969 (N_6969,N_4598,N_5433);
nand U6970 (N_6970,N_5688,N_3788);
nor U6971 (N_6971,N_5554,N_3141);
and U6972 (N_6972,N_5088,N_5484);
nor U6973 (N_6973,N_4001,N_3159);
and U6974 (N_6974,N_5363,N_3984);
and U6975 (N_6975,N_3951,N_4861);
nand U6976 (N_6976,N_4021,N_4252);
and U6977 (N_6977,N_5411,N_3584);
xor U6978 (N_6978,N_4509,N_5548);
nor U6979 (N_6979,N_5733,N_4053);
or U6980 (N_6980,N_4206,N_4033);
or U6981 (N_6981,N_4885,N_4697);
nand U6982 (N_6982,N_3491,N_5072);
nor U6983 (N_6983,N_3545,N_4901);
xnor U6984 (N_6984,N_4155,N_5553);
or U6985 (N_6985,N_3530,N_5802);
nand U6986 (N_6986,N_5222,N_4288);
xor U6987 (N_6987,N_5037,N_4103);
and U6988 (N_6988,N_4525,N_3479);
and U6989 (N_6989,N_5384,N_5832);
nor U6990 (N_6990,N_3302,N_5015);
or U6991 (N_6991,N_5725,N_5422);
and U6992 (N_6992,N_4654,N_3724);
nor U6993 (N_6993,N_5915,N_5883);
nor U6994 (N_6994,N_5333,N_3240);
nand U6995 (N_6995,N_3572,N_5868);
xnor U6996 (N_6996,N_4764,N_4600);
xnor U6997 (N_6997,N_5486,N_4201);
nand U6998 (N_6998,N_3536,N_3728);
nand U6999 (N_6999,N_5045,N_5750);
or U7000 (N_7000,N_3071,N_4718);
nand U7001 (N_7001,N_4017,N_5529);
nand U7002 (N_7002,N_3197,N_4363);
nor U7003 (N_7003,N_5378,N_5847);
nor U7004 (N_7004,N_3087,N_3976);
xnor U7005 (N_7005,N_5631,N_5290);
or U7006 (N_7006,N_4659,N_5143);
xnor U7007 (N_7007,N_3638,N_4949);
nand U7008 (N_7008,N_4629,N_4818);
and U7009 (N_7009,N_5732,N_4452);
nor U7010 (N_7010,N_4543,N_5021);
or U7011 (N_7011,N_4087,N_4506);
xor U7012 (N_7012,N_5551,N_3326);
xnor U7013 (N_7013,N_4517,N_3145);
xnor U7014 (N_7014,N_3070,N_4045);
xnor U7015 (N_7015,N_4871,N_5176);
nor U7016 (N_7016,N_4140,N_3389);
or U7017 (N_7017,N_4224,N_5584);
nand U7018 (N_7018,N_5784,N_3423);
nand U7019 (N_7019,N_5173,N_5198);
or U7020 (N_7020,N_4268,N_5438);
nand U7021 (N_7021,N_3878,N_3495);
nor U7022 (N_7022,N_5413,N_3663);
or U7023 (N_7023,N_5028,N_4014);
or U7024 (N_7024,N_5353,N_5775);
or U7025 (N_7025,N_4011,N_3101);
nand U7026 (N_7026,N_4003,N_3643);
and U7027 (N_7027,N_3397,N_5481);
or U7028 (N_7028,N_3586,N_3962);
and U7029 (N_7029,N_5528,N_3303);
xnor U7030 (N_7030,N_3037,N_4830);
and U7031 (N_7031,N_3318,N_4067);
or U7032 (N_7032,N_4930,N_3705);
xor U7033 (N_7033,N_3404,N_5188);
xnor U7034 (N_7034,N_3327,N_4849);
xnor U7035 (N_7035,N_3464,N_5071);
nand U7036 (N_7036,N_3126,N_5350);
nor U7037 (N_7037,N_4042,N_5399);
and U7038 (N_7038,N_5098,N_5606);
and U7039 (N_7039,N_4635,N_3658);
nor U7040 (N_7040,N_5539,N_3411);
and U7041 (N_7041,N_3187,N_3201);
xor U7042 (N_7042,N_4538,N_4806);
xor U7043 (N_7043,N_3998,N_4038);
or U7044 (N_7044,N_5893,N_4440);
and U7045 (N_7045,N_4370,N_3214);
nor U7046 (N_7046,N_3792,N_3835);
or U7047 (N_7047,N_3353,N_4141);
nand U7048 (N_7048,N_5512,N_4502);
and U7049 (N_7049,N_4468,N_3644);
xnor U7050 (N_7050,N_3316,N_5232);
nor U7051 (N_7051,N_3890,N_5156);
or U7052 (N_7052,N_5447,N_3843);
nand U7053 (N_7053,N_5646,N_3703);
xor U7054 (N_7054,N_3456,N_3029);
or U7055 (N_7055,N_5346,N_3113);
and U7056 (N_7056,N_4880,N_3293);
and U7057 (N_7057,N_4916,N_3168);
or U7058 (N_7058,N_5089,N_4732);
nor U7059 (N_7059,N_3144,N_3847);
and U7060 (N_7060,N_5590,N_5426);
or U7061 (N_7061,N_3561,N_3128);
or U7062 (N_7062,N_5785,N_5488);
nor U7063 (N_7063,N_4477,N_5562);
xnor U7064 (N_7064,N_4077,N_5666);
nand U7065 (N_7065,N_4028,N_4675);
nor U7066 (N_7066,N_4707,N_5269);
nand U7067 (N_7067,N_5503,N_5349);
or U7068 (N_7068,N_3022,N_3673);
nor U7069 (N_7069,N_3496,N_4008);
xnor U7070 (N_7070,N_4367,N_4075);
or U7071 (N_7071,N_5882,N_3424);
nor U7072 (N_7072,N_3802,N_3533);
nor U7073 (N_7073,N_3206,N_4310);
and U7074 (N_7074,N_5669,N_5518);
nor U7075 (N_7075,N_5986,N_5521);
xor U7076 (N_7076,N_4948,N_5284);
nor U7077 (N_7077,N_3160,N_3740);
and U7078 (N_7078,N_5668,N_3564);
nor U7079 (N_7079,N_3720,N_5096);
nor U7080 (N_7080,N_3871,N_5109);
xnor U7081 (N_7081,N_3557,N_3548);
nand U7082 (N_7082,N_5685,N_3862);
nor U7083 (N_7083,N_3758,N_5904);
and U7084 (N_7084,N_3328,N_4777);
and U7085 (N_7085,N_3034,N_3157);
nand U7086 (N_7086,N_5465,N_4549);
and U7087 (N_7087,N_4747,N_3981);
nand U7088 (N_7088,N_3357,N_4301);
nor U7089 (N_7089,N_4759,N_4234);
nor U7090 (N_7090,N_4914,N_3428);
and U7091 (N_7091,N_4241,N_5655);
and U7092 (N_7092,N_4190,N_4715);
xnor U7093 (N_7093,N_4271,N_5485);
and U7094 (N_7094,N_3459,N_4595);
or U7095 (N_7095,N_4970,N_3230);
and U7096 (N_7096,N_4810,N_3500);
nor U7097 (N_7097,N_3790,N_3143);
nand U7098 (N_7098,N_5181,N_5199);
nor U7099 (N_7099,N_5337,N_3900);
or U7100 (N_7100,N_4379,N_5260);
nor U7101 (N_7101,N_3235,N_5951);
or U7102 (N_7102,N_4046,N_3025);
and U7103 (N_7103,N_4205,N_3708);
nand U7104 (N_7104,N_4693,N_3452);
and U7105 (N_7105,N_4674,N_5248);
xor U7106 (N_7106,N_3515,N_3049);
nand U7107 (N_7107,N_5718,N_3311);
nor U7108 (N_7108,N_4702,N_3008);
xor U7109 (N_7109,N_5249,N_3226);
or U7110 (N_7110,N_3814,N_3153);
xnor U7111 (N_7111,N_5937,N_5765);
or U7112 (N_7112,N_3719,N_3935);
and U7113 (N_7113,N_5916,N_5746);
nand U7114 (N_7114,N_4644,N_5628);
nand U7115 (N_7115,N_3451,N_5150);
xor U7116 (N_7116,N_4665,N_5213);
nand U7117 (N_7117,N_4025,N_3905);
nand U7118 (N_7118,N_3258,N_3310);
xnor U7119 (N_7119,N_5245,N_5396);
nor U7120 (N_7120,N_3738,N_3634);
nand U7121 (N_7121,N_3937,N_3369);
xor U7122 (N_7122,N_5833,N_3993);
xor U7123 (N_7123,N_4064,N_5155);
xnor U7124 (N_7124,N_3147,N_3828);
nand U7125 (N_7125,N_5167,N_3282);
and U7126 (N_7126,N_3589,N_5761);
and U7127 (N_7127,N_5246,N_3131);
or U7128 (N_7128,N_4677,N_3795);
xnor U7129 (N_7129,N_5238,N_4261);
or U7130 (N_7130,N_4240,N_3765);
or U7131 (N_7131,N_4226,N_3818);
or U7132 (N_7132,N_3973,N_5989);
and U7133 (N_7133,N_5342,N_3961);
xor U7134 (N_7134,N_3453,N_5044);
nor U7135 (N_7135,N_4062,N_4238);
nand U7136 (N_7136,N_3785,N_4057);
nand U7137 (N_7137,N_4775,N_3565);
nor U7138 (N_7138,N_5697,N_5801);
and U7139 (N_7139,N_5402,N_3863);
and U7140 (N_7140,N_4832,N_5191);
or U7141 (N_7141,N_3671,N_5659);
or U7142 (N_7142,N_4688,N_5325);
nand U7143 (N_7143,N_4389,N_5327);
or U7144 (N_7144,N_4593,N_5879);
xnor U7145 (N_7145,N_4023,N_4497);
nor U7146 (N_7146,N_4108,N_3390);
or U7147 (N_7147,N_3056,N_4890);
or U7148 (N_7148,N_4283,N_3597);
or U7149 (N_7149,N_4010,N_3195);
and U7150 (N_7150,N_4920,N_4877);
and U7151 (N_7151,N_5954,N_3055);
or U7152 (N_7152,N_3815,N_3004);
nor U7153 (N_7153,N_3689,N_4059);
and U7154 (N_7154,N_4531,N_4237);
and U7155 (N_7155,N_5608,N_3386);
nand U7156 (N_7156,N_3616,N_3919);
or U7157 (N_7157,N_3722,N_3253);
and U7158 (N_7158,N_4346,N_4790);
or U7159 (N_7159,N_5707,N_4726);
nor U7160 (N_7160,N_3313,N_5421);
nor U7161 (N_7161,N_5867,N_3675);
nor U7162 (N_7162,N_5812,N_4413);
nor U7163 (N_7163,N_5540,N_4676);
and U7164 (N_7164,N_4636,N_4197);
and U7165 (N_7165,N_3341,N_4529);
or U7166 (N_7166,N_4754,N_3174);
nor U7167 (N_7167,N_3148,N_3699);
xnor U7168 (N_7168,N_5652,N_5206);
and U7169 (N_7169,N_4624,N_5452);
nor U7170 (N_7170,N_5527,N_4159);
nand U7171 (N_7171,N_3517,N_3642);
nor U7172 (N_7172,N_4313,N_4314);
nor U7173 (N_7173,N_3188,N_4080);
and U7174 (N_7174,N_4016,N_4072);
or U7175 (N_7175,N_3388,N_3544);
or U7176 (N_7176,N_3873,N_4546);
xnor U7177 (N_7177,N_4137,N_5470);
nor U7178 (N_7178,N_4005,N_5957);
xor U7179 (N_7179,N_4486,N_3826);
and U7180 (N_7180,N_3808,N_3233);
xnor U7181 (N_7181,N_4089,N_3422);
or U7182 (N_7182,N_4801,N_4561);
and U7183 (N_7183,N_3256,N_4070);
nor U7184 (N_7184,N_5455,N_5533);
xor U7185 (N_7185,N_5159,N_3666);
xnor U7186 (N_7186,N_5793,N_4910);
and U7187 (N_7187,N_5783,N_5680);
or U7188 (N_7188,N_5557,N_4862);
or U7189 (N_7189,N_3685,N_4908);
nand U7190 (N_7190,N_3053,N_5964);
and U7191 (N_7191,N_5170,N_5068);
nand U7192 (N_7192,N_4420,N_3472);
or U7193 (N_7193,N_4107,N_5114);
and U7194 (N_7194,N_5165,N_4897);
nor U7195 (N_7195,N_5272,N_3609);
nor U7196 (N_7196,N_4180,N_3462);
nand U7197 (N_7197,N_3620,N_3824);
nand U7198 (N_7198,N_4500,N_3614);
and U7199 (N_7199,N_4173,N_5012);
xor U7200 (N_7200,N_3393,N_4328);
nor U7201 (N_7201,N_3579,N_4648);
and U7202 (N_7202,N_5211,N_3447);
nand U7203 (N_7203,N_3122,N_3413);
nor U7204 (N_7204,N_4463,N_5846);
nor U7205 (N_7205,N_5430,N_4682);
nor U7206 (N_7206,N_4380,N_3237);
nor U7207 (N_7207,N_3701,N_5972);
or U7208 (N_7208,N_3212,N_3003);
nor U7209 (N_7209,N_5048,N_3065);
xor U7210 (N_7210,N_3980,N_5626);
or U7211 (N_7211,N_3490,N_5597);
and U7212 (N_7212,N_4408,N_3773);
nand U7213 (N_7213,N_5932,N_3083);
nand U7214 (N_7214,N_5676,N_4994);
nand U7215 (N_7215,N_5794,N_5994);
and U7216 (N_7216,N_5496,N_4478);
or U7217 (N_7217,N_3676,N_5076);
nor U7218 (N_7218,N_3570,N_5079);
xnor U7219 (N_7219,N_5582,N_5000);
or U7220 (N_7220,N_5135,N_3891);
nor U7221 (N_7221,N_3693,N_5926);
xor U7222 (N_7222,N_3103,N_3870);
nand U7223 (N_7223,N_3965,N_3718);
xnor U7224 (N_7224,N_4457,N_5463);
or U7225 (N_7225,N_4683,N_4186);
xnor U7226 (N_7226,N_5950,N_4550);
or U7227 (N_7227,N_5094,N_4218);
or U7228 (N_7228,N_3639,N_5013);
or U7229 (N_7229,N_5828,N_5035);
or U7230 (N_7230,N_3190,N_3216);
and U7231 (N_7231,N_3797,N_5681);
nand U7232 (N_7232,N_3438,N_4856);
and U7233 (N_7233,N_4239,N_4616);
nor U7234 (N_7234,N_4499,N_3038);
and U7235 (N_7235,N_4533,N_5328);
xor U7236 (N_7236,N_4039,N_3120);
and U7237 (N_7237,N_5405,N_5066);
nor U7238 (N_7238,N_5266,N_5200);
nand U7239 (N_7239,N_3882,N_5092);
nand U7240 (N_7240,N_3140,N_5360);
xor U7241 (N_7241,N_4633,N_5693);
nor U7242 (N_7242,N_5053,N_4647);
or U7243 (N_7243,N_5683,N_4507);
and U7244 (N_7244,N_5428,N_4776);
xor U7245 (N_7245,N_5621,N_3355);
nor U7246 (N_7246,N_5913,N_3267);
and U7247 (N_7247,N_3305,N_5412);
or U7248 (N_7248,N_5084,N_5154);
nor U7249 (N_7249,N_5458,N_3522);
nor U7250 (N_7250,N_5719,N_4143);
or U7251 (N_7251,N_4548,N_5921);
or U7252 (N_7252,N_3463,N_5477);
and U7253 (N_7253,N_3659,N_4126);
or U7254 (N_7254,N_3555,N_4119);
nor U7255 (N_7255,N_3974,N_4489);
nand U7256 (N_7256,N_3178,N_5786);
or U7257 (N_7257,N_3550,N_4095);
nand U7258 (N_7258,N_3281,N_5169);
nor U7259 (N_7259,N_4854,N_4179);
nand U7260 (N_7260,N_5087,N_5934);
xor U7261 (N_7261,N_4915,N_3966);
and U7262 (N_7262,N_5464,N_5129);
and U7263 (N_7263,N_4857,N_4058);
nand U7264 (N_7264,N_4639,N_5063);
nand U7265 (N_7265,N_5320,N_5815);
or U7266 (N_7266,N_5624,N_3537);
xor U7267 (N_7267,N_5543,N_5748);
or U7268 (N_7268,N_3664,N_4922);
or U7269 (N_7269,N_4614,N_3766);
nor U7270 (N_7270,N_3151,N_5040);
and U7271 (N_7271,N_5407,N_4491);
xor U7272 (N_7272,N_5133,N_4398);
or U7273 (N_7273,N_5568,N_5671);
or U7274 (N_7274,N_3425,N_4553);
and U7275 (N_7275,N_5419,N_5565);
nand U7276 (N_7276,N_3569,N_5193);
and U7277 (N_7277,N_5002,N_4357);
nor U7278 (N_7278,N_4895,N_5940);
xor U7279 (N_7279,N_4735,N_3199);
xor U7280 (N_7280,N_5799,N_3991);
nand U7281 (N_7281,N_5743,N_5397);
nor U7282 (N_7282,N_4952,N_5581);
xor U7283 (N_7283,N_3304,N_5577);
nand U7284 (N_7284,N_5716,N_3001);
and U7285 (N_7285,N_5931,N_4742);
nor U7286 (N_7286,N_4530,N_5826);
nor U7287 (N_7287,N_5020,N_3315);
nor U7288 (N_7288,N_3156,N_5894);
nor U7289 (N_7289,N_3627,N_4772);
or U7290 (N_7290,N_5132,N_4929);
xor U7291 (N_7291,N_5127,N_4695);
xnor U7292 (N_7292,N_4112,N_4339);
xnor U7293 (N_7293,N_4783,N_3737);
and U7294 (N_7294,N_4932,N_4704);
nor U7295 (N_7295,N_5286,N_3842);
or U7296 (N_7296,N_5023,N_4167);
and U7297 (N_7297,N_3499,N_4410);
or U7298 (N_7298,N_5494,N_4177);
or U7299 (N_7299,N_5900,N_3250);
xor U7300 (N_7300,N_3941,N_3040);
or U7301 (N_7301,N_4804,N_3124);
nor U7302 (N_7302,N_4617,N_5729);
nand U7303 (N_7303,N_3687,N_3485);
or U7304 (N_7304,N_5073,N_3920);
and U7305 (N_7305,N_4397,N_3913);
xor U7306 (N_7306,N_5362,N_3777);
xnor U7307 (N_7307,N_3990,N_5186);
and U7308 (N_7308,N_4816,N_3770);
nor U7309 (N_7309,N_4285,N_5252);
and U7310 (N_7310,N_4664,N_3810);
and U7311 (N_7311,N_4060,N_5097);
nand U7312 (N_7312,N_4935,N_4496);
and U7313 (N_7313,N_3761,N_4724);
and U7314 (N_7314,N_3931,N_3402);
and U7315 (N_7315,N_4812,N_3829);
and U7316 (N_7316,N_3918,N_4848);
nand U7317 (N_7317,N_4215,N_5961);
nand U7318 (N_7318,N_3000,N_4604);
and U7319 (N_7319,N_4613,N_4281);
nor U7320 (N_7320,N_4836,N_4157);
xnor U7321 (N_7321,N_5297,N_5656);
or U7322 (N_7322,N_3996,N_4171);
xnor U7323 (N_7323,N_3309,N_5966);
nor U7324 (N_7324,N_3448,N_4488);
and U7325 (N_7325,N_3114,N_3072);
xnor U7326 (N_7326,N_4596,N_3830);
nor U7327 (N_7327,N_5924,N_3844);
and U7328 (N_7328,N_5946,N_5256);
or U7329 (N_7329,N_3695,N_3470);
and U7330 (N_7330,N_3433,N_3241);
or U7331 (N_7331,N_5417,N_3283);
nor U7332 (N_7332,N_5454,N_5009);
nor U7333 (N_7333,N_4587,N_4603);
and U7334 (N_7334,N_5251,N_4770);
nor U7335 (N_7335,N_5278,N_4906);
and U7336 (N_7336,N_5858,N_3661);
or U7337 (N_7337,N_4152,N_4027);
nand U7338 (N_7338,N_3997,N_3198);
nor U7339 (N_7339,N_4378,N_5334);
and U7340 (N_7340,N_3342,N_4086);
xnor U7341 (N_7341,N_3894,N_3403);
xor U7342 (N_7342,N_3994,N_3360);
and U7343 (N_7343,N_5596,N_5569);
nor U7344 (N_7344,N_4881,N_4562);
or U7345 (N_7345,N_5126,N_5122);
and U7346 (N_7346,N_4400,N_5047);
nand U7347 (N_7347,N_5160,N_4934);
nand U7348 (N_7348,N_4798,N_3417);
nand U7349 (N_7349,N_3064,N_5029);
xor U7350 (N_7350,N_3987,N_3540);
xor U7351 (N_7351,N_3133,N_3344);
nor U7352 (N_7352,N_5451,N_4899);
nor U7353 (N_7353,N_3804,N_3889);
xor U7354 (N_7354,N_5917,N_3480);
xnor U7355 (N_7355,N_4114,N_5583);
xor U7356 (N_7356,N_5956,N_4250);
nor U7357 (N_7357,N_4661,N_3455);
or U7358 (N_7358,N_4264,N_4063);
and U7359 (N_7359,N_3592,N_4135);
xor U7360 (N_7360,N_5625,N_3983);
nand U7361 (N_7361,N_4996,N_4006);
and U7362 (N_7362,N_5651,N_3066);
xor U7363 (N_7363,N_3439,N_4819);
and U7364 (N_7364,N_4769,N_4368);
or U7365 (N_7365,N_5250,N_3031);
nand U7366 (N_7366,N_5525,N_5644);
nand U7367 (N_7367,N_5011,N_4056);
and U7368 (N_7368,N_5575,N_3715);
xnor U7369 (N_7369,N_3044,N_5125);
and U7370 (N_7370,N_4641,N_4809);
nand U7371 (N_7371,N_5196,N_5024);
xor U7372 (N_7372,N_3698,N_3163);
and U7373 (N_7373,N_4098,N_5664);
nand U7374 (N_7374,N_3933,N_5751);
or U7375 (N_7375,N_5573,N_4541);
and U7376 (N_7376,N_3268,N_3292);
or U7377 (N_7377,N_5220,N_5599);
nor U7378 (N_7378,N_4984,N_4467);
nor U7379 (N_7379,N_5500,N_4958);
or U7380 (N_7380,N_3893,N_3354);
xnor U7381 (N_7381,N_4508,N_4760);
nor U7382 (N_7382,N_4498,N_5205);
or U7383 (N_7383,N_4439,N_4951);
and U7384 (N_7384,N_4993,N_4164);
xnor U7385 (N_7385,N_5270,N_3079);
nor U7386 (N_7386,N_4679,N_4356);
nand U7387 (N_7387,N_5395,N_4865);
nor U7388 (N_7388,N_3036,N_3102);
nor U7389 (N_7389,N_3172,N_3219);
xor U7390 (N_7390,N_3953,N_3649);
and U7391 (N_7391,N_5078,N_4196);
nand U7392 (N_7392,N_3426,N_4513);
nor U7393 (N_7393,N_5844,N_4348);
nor U7394 (N_7394,N_3923,N_4423);
nand U7395 (N_7395,N_5993,N_4579);
and U7396 (N_7396,N_4845,N_4495);
xnor U7397 (N_7397,N_3220,N_3741);
and U7398 (N_7398,N_4248,N_4407);
and U7399 (N_7399,N_3625,N_3849);
nand U7400 (N_7400,N_3410,N_4031);
nor U7401 (N_7401,N_4859,N_3325);
xor U7402 (N_7402,N_3684,N_5420);
and U7403 (N_7403,N_5059,N_4736);
or U7404 (N_7404,N_5996,N_5310);
and U7405 (N_7405,N_3503,N_4891);
and U7406 (N_7406,N_5326,N_3917);
nand U7407 (N_7407,N_5341,N_4176);
xnor U7408 (N_7408,N_3596,N_5393);
xnor U7409 (N_7409,N_4069,N_4030);
nand U7410 (N_7410,N_5445,N_3852);
nor U7411 (N_7411,N_5322,N_4473);
nand U7412 (N_7412,N_5093,N_3902);
nor U7413 (N_7413,N_3028,N_3213);
nor U7414 (N_7414,N_5770,N_4322);
xnor U7415 (N_7415,N_3978,N_5643);
or U7416 (N_7416,N_5928,N_5689);
xor U7417 (N_7417,N_4851,N_4127);
nor U7418 (N_7418,N_5546,N_3471);
or U7419 (N_7419,N_3574,N_5536);
xnor U7420 (N_7420,N_5435,N_3048);
nand U7421 (N_7421,N_3633,N_4332);
nor U7422 (N_7422,N_4345,N_4544);
and U7423 (N_7423,N_4352,N_3002);
or U7424 (N_7424,N_5798,N_4981);
nand U7425 (N_7425,N_5061,N_4273);
nor U7426 (N_7426,N_5945,N_4493);
nand U7427 (N_7427,N_4278,N_3296);
xor U7428 (N_7428,N_4896,N_3054);
or U7429 (N_7429,N_4262,N_5343);
xnor U7430 (N_7430,N_4942,N_5755);
or U7431 (N_7431,N_4222,N_4305);
xor U7432 (N_7432,N_4012,N_5549);
xnor U7433 (N_7433,N_3799,N_3583);
nand U7434 (N_7434,N_5817,N_5330);
nor U7435 (N_7435,N_5375,N_5885);
nand U7436 (N_7436,N_5566,N_3013);
nand U7437 (N_7437,N_5441,N_4678);
and U7438 (N_7438,N_4536,N_4800);
xnor U7439 (N_7439,N_5151,N_5487);
nor U7440 (N_7440,N_3753,N_5768);
or U7441 (N_7441,N_3473,N_4412);
and U7442 (N_7442,N_4361,N_5520);
or U7443 (N_7443,N_3925,N_3958);
xor U7444 (N_7444,N_4585,N_5207);
or U7445 (N_7445,N_3690,N_4712);
xor U7446 (N_7446,N_4047,N_3652);
nor U7447 (N_7447,N_3702,N_4351);
and U7448 (N_7448,N_4522,N_3960);
and U7449 (N_7449,N_5457,N_3581);
nand U7450 (N_7450,N_4071,N_3181);
nor U7451 (N_7451,N_4168,N_5663);
and U7452 (N_7452,N_5382,N_3259);
nand U7453 (N_7453,N_4839,N_5898);
xor U7454 (N_7454,N_4632,N_3150);
or U7455 (N_7455,N_5627,N_5731);
xnor U7456 (N_7456,N_5090,N_4813);
nand U7457 (N_7457,N_4082,N_5918);
nor U7458 (N_7458,N_5649,N_4694);
nand U7459 (N_7459,N_5574,N_5895);
and U7460 (N_7460,N_5634,N_5381);
nand U7461 (N_7461,N_4302,N_4347);
nand U7462 (N_7462,N_3107,N_3204);
nand U7463 (N_7463,N_5443,N_4004);
nor U7464 (N_7464,N_4055,N_3934);
or U7465 (N_7465,N_3848,N_4421);
or U7466 (N_7466,N_3222,N_3938);
nor U7467 (N_7467,N_4188,N_5881);
xor U7468 (N_7468,N_5499,N_4000);
nor U7469 (N_7469,N_5189,N_4700);
or U7470 (N_7470,N_5772,N_4490);
nand U7471 (N_7471,N_4933,N_5988);
nand U7472 (N_7472,N_5851,N_5686);
xor U7473 (N_7473,N_5497,N_3822);
and U7474 (N_7474,N_4685,N_4120);
and U7475 (N_7475,N_4658,N_5182);
or U7476 (N_7476,N_5157,N_3368);
xnor U7477 (N_7477,N_3764,N_5662);
and U7478 (N_7478,N_3091,N_5974);
nor U7479 (N_7479,N_3872,N_4924);
and U7480 (N_7480,N_5558,N_3834);
nor U7481 (N_7481,N_3332,N_4667);
or U7482 (N_7482,N_3446,N_4308);
or U7483 (N_7483,N_5777,N_3930);
xnor U7484 (N_7484,N_5324,N_4640);
nand U7485 (N_7485,N_3287,N_3440);
nand U7486 (N_7486,N_3170,N_4366);
xnor U7487 (N_7487,N_3081,N_3015);
nor U7488 (N_7488,N_3032,N_4094);
xor U7489 (N_7489,N_4824,N_4912);
and U7490 (N_7490,N_3380,N_4402);
nor U7491 (N_7491,N_4998,N_4269);
nor U7492 (N_7492,N_4692,N_3278);
xnor U7493 (N_7493,N_3892,N_4195);
nor U7494 (N_7494,N_5149,N_4666);
or U7495 (N_7495,N_3904,N_4373);
xnor U7496 (N_7496,N_3791,N_5398);
or U7497 (N_7497,N_4245,N_5262);
and U7498 (N_7498,N_5564,N_5124);
and U7499 (N_7499,N_5074,N_3865);
nand U7500 (N_7500,N_3399,N_4744);
or U7501 (N_7501,N_5535,N_3405);
nand U7502 (N_7502,N_5649,N_3140);
nor U7503 (N_7503,N_5713,N_3656);
nand U7504 (N_7504,N_5726,N_3120);
xor U7505 (N_7505,N_5777,N_3686);
nand U7506 (N_7506,N_5627,N_3168);
nand U7507 (N_7507,N_5135,N_4548);
nand U7508 (N_7508,N_5476,N_3850);
and U7509 (N_7509,N_4874,N_3942);
and U7510 (N_7510,N_4081,N_4353);
and U7511 (N_7511,N_3630,N_5775);
or U7512 (N_7512,N_3437,N_4529);
or U7513 (N_7513,N_4830,N_3655);
or U7514 (N_7514,N_3233,N_4074);
xnor U7515 (N_7515,N_5684,N_4436);
and U7516 (N_7516,N_5860,N_5913);
xor U7517 (N_7517,N_3937,N_5669);
or U7518 (N_7518,N_5925,N_5768);
or U7519 (N_7519,N_4473,N_5055);
or U7520 (N_7520,N_3534,N_4823);
or U7521 (N_7521,N_3911,N_3854);
or U7522 (N_7522,N_4492,N_3952);
nor U7523 (N_7523,N_3634,N_4551);
nor U7524 (N_7524,N_3194,N_3907);
nor U7525 (N_7525,N_3059,N_4837);
and U7526 (N_7526,N_3879,N_3516);
xnor U7527 (N_7527,N_5533,N_4427);
nor U7528 (N_7528,N_5427,N_3606);
or U7529 (N_7529,N_4527,N_3596);
nor U7530 (N_7530,N_3686,N_3983);
xnor U7531 (N_7531,N_5104,N_3843);
nor U7532 (N_7532,N_3653,N_5402);
nor U7533 (N_7533,N_3096,N_4247);
nand U7534 (N_7534,N_4953,N_4794);
xnor U7535 (N_7535,N_5065,N_5611);
nand U7536 (N_7536,N_3085,N_4909);
xnor U7537 (N_7537,N_5987,N_3430);
nor U7538 (N_7538,N_3433,N_3557);
xor U7539 (N_7539,N_3072,N_4800);
or U7540 (N_7540,N_3804,N_4350);
xor U7541 (N_7541,N_5006,N_3477);
nor U7542 (N_7542,N_3914,N_3479);
nand U7543 (N_7543,N_3517,N_5560);
nand U7544 (N_7544,N_5658,N_4541);
nand U7545 (N_7545,N_5058,N_4619);
nor U7546 (N_7546,N_5059,N_5838);
nor U7547 (N_7547,N_3483,N_3301);
and U7548 (N_7548,N_5832,N_5162);
nor U7549 (N_7549,N_5454,N_5767);
or U7550 (N_7550,N_4637,N_3169);
or U7551 (N_7551,N_4732,N_4314);
and U7552 (N_7552,N_3368,N_5800);
or U7553 (N_7553,N_4526,N_5303);
nand U7554 (N_7554,N_5205,N_3988);
nand U7555 (N_7555,N_3081,N_5109);
or U7556 (N_7556,N_4554,N_3048);
nand U7557 (N_7557,N_3052,N_3039);
nor U7558 (N_7558,N_4734,N_4391);
nor U7559 (N_7559,N_5522,N_4015);
nand U7560 (N_7560,N_3323,N_3030);
or U7561 (N_7561,N_3991,N_5187);
nand U7562 (N_7562,N_4215,N_4354);
and U7563 (N_7563,N_5264,N_5546);
xnor U7564 (N_7564,N_4886,N_5273);
xnor U7565 (N_7565,N_5803,N_4647);
or U7566 (N_7566,N_4219,N_3992);
nand U7567 (N_7567,N_4481,N_4691);
or U7568 (N_7568,N_5146,N_5935);
xnor U7569 (N_7569,N_3879,N_4041);
nor U7570 (N_7570,N_5523,N_4541);
or U7571 (N_7571,N_5108,N_5456);
nand U7572 (N_7572,N_4502,N_5906);
nand U7573 (N_7573,N_4260,N_3144);
xnor U7574 (N_7574,N_4710,N_3982);
or U7575 (N_7575,N_3294,N_3043);
and U7576 (N_7576,N_3216,N_4436);
nand U7577 (N_7577,N_3315,N_5914);
xor U7578 (N_7578,N_4909,N_3154);
xnor U7579 (N_7579,N_5162,N_4633);
nor U7580 (N_7580,N_3882,N_3854);
xor U7581 (N_7581,N_4545,N_5910);
nand U7582 (N_7582,N_4384,N_4205);
nor U7583 (N_7583,N_3223,N_3977);
nand U7584 (N_7584,N_3901,N_3621);
nor U7585 (N_7585,N_5879,N_5070);
nand U7586 (N_7586,N_5284,N_3910);
nor U7587 (N_7587,N_5649,N_3608);
xor U7588 (N_7588,N_4874,N_3964);
or U7589 (N_7589,N_4531,N_5218);
nand U7590 (N_7590,N_4520,N_3205);
or U7591 (N_7591,N_3867,N_3469);
xnor U7592 (N_7592,N_4666,N_4969);
or U7593 (N_7593,N_5071,N_3149);
nor U7594 (N_7594,N_5154,N_5386);
and U7595 (N_7595,N_3328,N_4838);
nor U7596 (N_7596,N_4621,N_4914);
nand U7597 (N_7597,N_4494,N_4532);
and U7598 (N_7598,N_5825,N_5371);
nand U7599 (N_7599,N_4082,N_3463);
xor U7600 (N_7600,N_5123,N_3105);
or U7601 (N_7601,N_3362,N_3696);
and U7602 (N_7602,N_3035,N_3510);
or U7603 (N_7603,N_3581,N_3322);
xor U7604 (N_7604,N_3514,N_3757);
nor U7605 (N_7605,N_3874,N_5397);
nand U7606 (N_7606,N_3747,N_3754);
xnor U7607 (N_7607,N_4625,N_3367);
nand U7608 (N_7608,N_4590,N_3351);
or U7609 (N_7609,N_3974,N_4431);
xnor U7610 (N_7610,N_4603,N_3010);
xnor U7611 (N_7611,N_4571,N_3302);
nand U7612 (N_7612,N_4727,N_5367);
and U7613 (N_7613,N_4530,N_5654);
or U7614 (N_7614,N_4132,N_3018);
nor U7615 (N_7615,N_4326,N_5975);
or U7616 (N_7616,N_4801,N_5481);
or U7617 (N_7617,N_4363,N_4808);
nor U7618 (N_7618,N_5327,N_5617);
nor U7619 (N_7619,N_4443,N_3172);
nand U7620 (N_7620,N_5863,N_4850);
nand U7621 (N_7621,N_3886,N_5422);
or U7622 (N_7622,N_5120,N_3774);
and U7623 (N_7623,N_5609,N_3189);
nor U7624 (N_7624,N_4495,N_3557);
nor U7625 (N_7625,N_4487,N_4266);
nor U7626 (N_7626,N_4516,N_4584);
or U7627 (N_7627,N_5702,N_5744);
nor U7628 (N_7628,N_3944,N_5680);
and U7629 (N_7629,N_5387,N_3379);
or U7630 (N_7630,N_5803,N_3740);
xor U7631 (N_7631,N_4395,N_4624);
xor U7632 (N_7632,N_5121,N_5931);
and U7633 (N_7633,N_3013,N_3071);
nor U7634 (N_7634,N_5198,N_3701);
nand U7635 (N_7635,N_4114,N_4587);
nand U7636 (N_7636,N_4080,N_3143);
or U7637 (N_7637,N_3880,N_5003);
xnor U7638 (N_7638,N_4183,N_3689);
and U7639 (N_7639,N_5432,N_4594);
nand U7640 (N_7640,N_4263,N_5643);
or U7641 (N_7641,N_5641,N_3345);
or U7642 (N_7642,N_5422,N_5693);
nand U7643 (N_7643,N_3266,N_4842);
nand U7644 (N_7644,N_4434,N_3973);
nor U7645 (N_7645,N_5411,N_5699);
nor U7646 (N_7646,N_3929,N_4511);
nor U7647 (N_7647,N_4916,N_5892);
and U7648 (N_7648,N_4400,N_5828);
nor U7649 (N_7649,N_5041,N_4464);
nand U7650 (N_7650,N_3904,N_5978);
xor U7651 (N_7651,N_5561,N_4848);
nor U7652 (N_7652,N_3181,N_4096);
nor U7653 (N_7653,N_4048,N_3561);
or U7654 (N_7654,N_4035,N_4894);
xor U7655 (N_7655,N_3734,N_3342);
and U7656 (N_7656,N_4781,N_5661);
nand U7657 (N_7657,N_5459,N_4475);
and U7658 (N_7658,N_3703,N_4019);
or U7659 (N_7659,N_4722,N_4807);
nor U7660 (N_7660,N_5902,N_3450);
and U7661 (N_7661,N_3890,N_5977);
nand U7662 (N_7662,N_4273,N_3603);
xor U7663 (N_7663,N_5452,N_5109);
xnor U7664 (N_7664,N_4049,N_5280);
and U7665 (N_7665,N_4238,N_4979);
xnor U7666 (N_7666,N_5846,N_5543);
xnor U7667 (N_7667,N_3511,N_4797);
xor U7668 (N_7668,N_4857,N_5909);
and U7669 (N_7669,N_5313,N_4864);
nor U7670 (N_7670,N_5986,N_3996);
and U7671 (N_7671,N_5700,N_4444);
or U7672 (N_7672,N_3472,N_5157);
xnor U7673 (N_7673,N_4929,N_5052);
or U7674 (N_7674,N_5440,N_5500);
and U7675 (N_7675,N_4098,N_5593);
or U7676 (N_7676,N_3850,N_4575);
or U7677 (N_7677,N_3856,N_3841);
and U7678 (N_7678,N_3852,N_5892);
and U7679 (N_7679,N_5920,N_3075);
and U7680 (N_7680,N_4515,N_3863);
nor U7681 (N_7681,N_4467,N_4034);
and U7682 (N_7682,N_5796,N_5635);
xnor U7683 (N_7683,N_3155,N_3654);
nand U7684 (N_7684,N_4550,N_4631);
and U7685 (N_7685,N_5072,N_3788);
xnor U7686 (N_7686,N_5596,N_3786);
and U7687 (N_7687,N_5999,N_5858);
and U7688 (N_7688,N_3431,N_4513);
xnor U7689 (N_7689,N_3946,N_4806);
and U7690 (N_7690,N_3474,N_4795);
and U7691 (N_7691,N_4644,N_4452);
xor U7692 (N_7692,N_5851,N_4231);
nor U7693 (N_7693,N_5557,N_3156);
xor U7694 (N_7694,N_5288,N_3753);
nor U7695 (N_7695,N_3308,N_3273);
or U7696 (N_7696,N_5578,N_4722);
nand U7697 (N_7697,N_5909,N_4026);
nor U7698 (N_7698,N_5025,N_3415);
and U7699 (N_7699,N_4119,N_4068);
and U7700 (N_7700,N_5278,N_4930);
xnor U7701 (N_7701,N_4112,N_3165);
and U7702 (N_7702,N_3911,N_3626);
and U7703 (N_7703,N_3817,N_5684);
nand U7704 (N_7704,N_3236,N_3890);
and U7705 (N_7705,N_5230,N_5977);
xnor U7706 (N_7706,N_5291,N_3024);
nand U7707 (N_7707,N_4142,N_4215);
and U7708 (N_7708,N_4336,N_5074);
xor U7709 (N_7709,N_3127,N_4036);
nor U7710 (N_7710,N_5454,N_4480);
and U7711 (N_7711,N_3515,N_5779);
xnor U7712 (N_7712,N_3688,N_5307);
nand U7713 (N_7713,N_4037,N_5791);
xnor U7714 (N_7714,N_4735,N_5059);
and U7715 (N_7715,N_4174,N_3390);
and U7716 (N_7716,N_4420,N_4559);
nand U7717 (N_7717,N_5977,N_4607);
and U7718 (N_7718,N_5372,N_5889);
or U7719 (N_7719,N_4948,N_3813);
nand U7720 (N_7720,N_5710,N_5599);
and U7721 (N_7721,N_5359,N_3816);
xor U7722 (N_7722,N_4693,N_5172);
xor U7723 (N_7723,N_3084,N_4529);
or U7724 (N_7724,N_4605,N_3597);
nor U7725 (N_7725,N_3769,N_3789);
xnor U7726 (N_7726,N_3361,N_3567);
nor U7727 (N_7727,N_3272,N_4577);
or U7728 (N_7728,N_4272,N_4826);
or U7729 (N_7729,N_4030,N_4757);
nand U7730 (N_7730,N_3336,N_5068);
and U7731 (N_7731,N_5416,N_3115);
or U7732 (N_7732,N_3758,N_5896);
xor U7733 (N_7733,N_5051,N_4948);
or U7734 (N_7734,N_3513,N_4607);
nand U7735 (N_7735,N_4353,N_4707);
nor U7736 (N_7736,N_5644,N_4496);
nand U7737 (N_7737,N_3148,N_5512);
xnor U7738 (N_7738,N_3143,N_5348);
nand U7739 (N_7739,N_4001,N_3061);
xnor U7740 (N_7740,N_4307,N_3016);
nand U7741 (N_7741,N_4606,N_4078);
xor U7742 (N_7742,N_5634,N_4219);
nor U7743 (N_7743,N_4367,N_5176);
nor U7744 (N_7744,N_4309,N_5856);
and U7745 (N_7745,N_3555,N_5486);
xor U7746 (N_7746,N_3767,N_5493);
and U7747 (N_7747,N_4244,N_5504);
and U7748 (N_7748,N_4006,N_5631);
and U7749 (N_7749,N_4297,N_5937);
xor U7750 (N_7750,N_3755,N_3211);
xnor U7751 (N_7751,N_5613,N_5845);
xnor U7752 (N_7752,N_4288,N_4555);
or U7753 (N_7753,N_5577,N_4331);
nor U7754 (N_7754,N_5197,N_4158);
xor U7755 (N_7755,N_5407,N_4525);
or U7756 (N_7756,N_5251,N_3590);
or U7757 (N_7757,N_3355,N_4900);
xnor U7758 (N_7758,N_5967,N_5469);
nor U7759 (N_7759,N_4761,N_4073);
nand U7760 (N_7760,N_4858,N_5622);
xnor U7761 (N_7761,N_3933,N_4709);
and U7762 (N_7762,N_4626,N_3603);
nand U7763 (N_7763,N_5771,N_4765);
nor U7764 (N_7764,N_3302,N_3482);
or U7765 (N_7765,N_4064,N_4512);
nor U7766 (N_7766,N_5303,N_3085);
xnor U7767 (N_7767,N_3654,N_4601);
and U7768 (N_7768,N_3786,N_4524);
nand U7769 (N_7769,N_3927,N_4415);
or U7770 (N_7770,N_5061,N_5130);
nand U7771 (N_7771,N_4738,N_3566);
or U7772 (N_7772,N_4286,N_4145);
nor U7773 (N_7773,N_4479,N_3040);
xor U7774 (N_7774,N_3243,N_4379);
or U7775 (N_7775,N_3647,N_5003);
nor U7776 (N_7776,N_5354,N_5046);
nand U7777 (N_7777,N_5941,N_5680);
xnor U7778 (N_7778,N_5473,N_5756);
xnor U7779 (N_7779,N_3866,N_5797);
nand U7780 (N_7780,N_4268,N_4376);
nor U7781 (N_7781,N_5958,N_3742);
and U7782 (N_7782,N_5260,N_3148);
nand U7783 (N_7783,N_5354,N_4018);
and U7784 (N_7784,N_4114,N_3293);
nand U7785 (N_7785,N_4982,N_5453);
xor U7786 (N_7786,N_5692,N_3032);
or U7787 (N_7787,N_5155,N_3566);
xnor U7788 (N_7788,N_4715,N_4144);
nand U7789 (N_7789,N_3513,N_4426);
and U7790 (N_7790,N_5224,N_4872);
and U7791 (N_7791,N_5363,N_4976);
nand U7792 (N_7792,N_4142,N_5994);
xor U7793 (N_7793,N_5720,N_3799);
and U7794 (N_7794,N_4434,N_4134);
or U7795 (N_7795,N_5063,N_5137);
nand U7796 (N_7796,N_4448,N_5627);
nand U7797 (N_7797,N_4000,N_4202);
and U7798 (N_7798,N_4453,N_3574);
xor U7799 (N_7799,N_5549,N_3171);
nand U7800 (N_7800,N_4027,N_3162);
nor U7801 (N_7801,N_5980,N_3222);
xnor U7802 (N_7802,N_3824,N_5777);
and U7803 (N_7803,N_3144,N_4724);
nand U7804 (N_7804,N_3906,N_4820);
nand U7805 (N_7805,N_5627,N_4424);
nor U7806 (N_7806,N_4115,N_5717);
or U7807 (N_7807,N_5448,N_3102);
xnor U7808 (N_7808,N_4414,N_3367);
or U7809 (N_7809,N_4927,N_3241);
xor U7810 (N_7810,N_4539,N_3331);
nand U7811 (N_7811,N_4292,N_5737);
xor U7812 (N_7812,N_3651,N_4187);
xor U7813 (N_7813,N_3025,N_4350);
nor U7814 (N_7814,N_5106,N_4258);
or U7815 (N_7815,N_4965,N_4273);
nand U7816 (N_7816,N_3055,N_3160);
and U7817 (N_7817,N_4611,N_3695);
or U7818 (N_7818,N_5255,N_3182);
or U7819 (N_7819,N_4171,N_5068);
and U7820 (N_7820,N_5055,N_4678);
and U7821 (N_7821,N_3815,N_5333);
xnor U7822 (N_7822,N_3903,N_4543);
xor U7823 (N_7823,N_3691,N_5374);
xor U7824 (N_7824,N_4436,N_5781);
and U7825 (N_7825,N_4928,N_5028);
xnor U7826 (N_7826,N_5942,N_4938);
nand U7827 (N_7827,N_3081,N_3804);
or U7828 (N_7828,N_3607,N_5526);
or U7829 (N_7829,N_4401,N_5506);
or U7830 (N_7830,N_4816,N_5247);
or U7831 (N_7831,N_5254,N_5672);
or U7832 (N_7832,N_4869,N_5421);
and U7833 (N_7833,N_5358,N_3466);
and U7834 (N_7834,N_4836,N_5592);
and U7835 (N_7835,N_3500,N_5420);
nand U7836 (N_7836,N_4369,N_3861);
and U7837 (N_7837,N_5113,N_5491);
xnor U7838 (N_7838,N_5781,N_3306);
xor U7839 (N_7839,N_4329,N_4464);
nand U7840 (N_7840,N_4683,N_4881);
nand U7841 (N_7841,N_5831,N_3013);
xnor U7842 (N_7842,N_3350,N_3359);
nand U7843 (N_7843,N_3230,N_4517);
xnor U7844 (N_7844,N_5953,N_3271);
nor U7845 (N_7845,N_3107,N_4932);
or U7846 (N_7846,N_3072,N_4172);
nor U7847 (N_7847,N_4374,N_3639);
and U7848 (N_7848,N_4115,N_3268);
nor U7849 (N_7849,N_3485,N_3156);
xnor U7850 (N_7850,N_3280,N_4730);
and U7851 (N_7851,N_4848,N_3477);
xnor U7852 (N_7852,N_5738,N_5769);
or U7853 (N_7853,N_4999,N_5115);
xnor U7854 (N_7854,N_4960,N_4179);
or U7855 (N_7855,N_4427,N_5734);
or U7856 (N_7856,N_4380,N_4526);
or U7857 (N_7857,N_4493,N_3544);
xnor U7858 (N_7858,N_5382,N_3713);
and U7859 (N_7859,N_3977,N_5478);
xor U7860 (N_7860,N_5011,N_5767);
or U7861 (N_7861,N_5006,N_5781);
or U7862 (N_7862,N_3739,N_3239);
nand U7863 (N_7863,N_3175,N_4826);
nor U7864 (N_7864,N_4743,N_3504);
nor U7865 (N_7865,N_5867,N_4537);
or U7866 (N_7866,N_5593,N_4005);
nor U7867 (N_7867,N_4065,N_4165);
or U7868 (N_7868,N_3585,N_4541);
and U7869 (N_7869,N_3206,N_4967);
nor U7870 (N_7870,N_5942,N_5874);
xor U7871 (N_7871,N_4205,N_3162);
and U7872 (N_7872,N_3681,N_5865);
xnor U7873 (N_7873,N_3608,N_3716);
or U7874 (N_7874,N_3999,N_3152);
nor U7875 (N_7875,N_3021,N_5345);
and U7876 (N_7876,N_4920,N_3490);
nand U7877 (N_7877,N_5211,N_5355);
nor U7878 (N_7878,N_5306,N_3640);
nor U7879 (N_7879,N_3411,N_3500);
nor U7880 (N_7880,N_4889,N_4809);
nand U7881 (N_7881,N_3065,N_3631);
and U7882 (N_7882,N_5323,N_4627);
and U7883 (N_7883,N_5486,N_4981);
nor U7884 (N_7884,N_4439,N_5371);
and U7885 (N_7885,N_5908,N_3222);
xnor U7886 (N_7886,N_3133,N_4315);
nor U7887 (N_7887,N_3741,N_5831);
and U7888 (N_7888,N_5587,N_4171);
nand U7889 (N_7889,N_4223,N_4024);
or U7890 (N_7890,N_3777,N_5020);
nand U7891 (N_7891,N_5442,N_4694);
nand U7892 (N_7892,N_3702,N_3958);
or U7893 (N_7893,N_5119,N_5329);
nor U7894 (N_7894,N_4750,N_3317);
and U7895 (N_7895,N_4046,N_5179);
or U7896 (N_7896,N_5140,N_4530);
nand U7897 (N_7897,N_5331,N_3953);
or U7898 (N_7898,N_5455,N_5900);
or U7899 (N_7899,N_5324,N_4107);
xor U7900 (N_7900,N_3458,N_5812);
or U7901 (N_7901,N_4698,N_3383);
or U7902 (N_7902,N_4429,N_3175);
or U7903 (N_7903,N_3393,N_3292);
or U7904 (N_7904,N_3745,N_4737);
and U7905 (N_7905,N_5098,N_4814);
nand U7906 (N_7906,N_5553,N_5608);
xor U7907 (N_7907,N_4649,N_5808);
nand U7908 (N_7908,N_5412,N_3533);
and U7909 (N_7909,N_5744,N_3458);
or U7910 (N_7910,N_5861,N_4031);
and U7911 (N_7911,N_4627,N_5586);
or U7912 (N_7912,N_3612,N_3213);
nand U7913 (N_7913,N_4153,N_4311);
or U7914 (N_7914,N_3181,N_3639);
xnor U7915 (N_7915,N_4586,N_3832);
nor U7916 (N_7916,N_4246,N_3160);
nand U7917 (N_7917,N_3913,N_4278);
or U7918 (N_7918,N_5152,N_5375);
xor U7919 (N_7919,N_5906,N_4683);
or U7920 (N_7920,N_4793,N_5987);
and U7921 (N_7921,N_5949,N_5956);
or U7922 (N_7922,N_5353,N_4850);
nor U7923 (N_7923,N_4917,N_3282);
nor U7924 (N_7924,N_4056,N_5066);
nor U7925 (N_7925,N_5372,N_3474);
nor U7926 (N_7926,N_4091,N_4820);
and U7927 (N_7927,N_3984,N_4130);
or U7928 (N_7928,N_5270,N_4226);
and U7929 (N_7929,N_3188,N_5794);
nand U7930 (N_7930,N_5393,N_5542);
or U7931 (N_7931,N_5583,N_3704);
or U7932 (N_7932,N_4866,N_3094);
or U7933 (N_7933,N_5047,N_4989);
nor U7934 (N_7934,N_5321,N_3672);
xnor U7935 (N_7935,N_5833,N_3094);
or U7936 (N_7936,N_4411,N_4943);
or U7937 (N_7937,N_5673,N_3036);
and U7938 (N_7938,N_4646,N_3628);
nand U7939 (N_7939,N_3124,N_3286);
or U7940 (N_7940,N_3448,N_5516);
xor U7941 (N_7941,N_5219,N_4746);
and U7942 (N_7942,N_4240,N_4728);
nor U7943 (N_7943,N_3703,N_4693);
nand U7944 (N_7944,N_3081,N_4180);
xor U7945 (N_7945,N_3559,N_5414);
and U7946 (N_7946,N_4840,N_5872);
or U7947 (N_7947,N_4989,N_4094);
and U7948 (N_7948,N_3330,N_3644);
xnor U7949 (N_7949,N_5652,N_3607);
xnor U7950 (N_7950,N_4959,N_5593);
nor U7951 (N_7951,N_5178,N_3810);
nor U7952 (N_7952,N_3093,N_5519);
or U7953 (N_7953,N_3937,N_5098);
nand U7954 (N_7954,N_3411,N_5658);
and U7955 (N_7955,N_5205,N_5672);
nor U7956 (N_7956,N_3635,N_5091);
nor U7957 (N_7957,N_3675,N_4403);
and U7958 (N_7958,N_5455,N_3130);
nand U7959 (N_7959,N_4031,N_3219);
and U7960 (N_7960,N_4690,N_5053);
or U7961 (N_7961,N_4369,N_5117);
nor U7962 (N_7962,N_3845,N_3199);
and U7963 (N_7963,N_3977,N_5264);
xnor U7964 (N_7964,N_3708,N_5970);
nor U7965 (N_7965,N_4582,N_3583);
and U7966 (N_7966,N_5632,N_3237);
nand U7967 (N_7967,N_4174,N_4018);
nand U7968 (N_7968,N_3237,N_3535);
or U7969 (N_7969,N_5414,N_5777);
xnor U7970 (N_7970,N_4922,N_3638);
xnor U7971 (N_7971,N_5619,N_3873);
nor U7972 (N_7972,N_5802,N_5381);
xnor U7973 (N_7973,N_4504,N_5558);
nor U7974 (N_7974,N_4244,N_5235);
xnor U7975 (N_7975,N_5059,N_4954);
and U7976 (N_7976,N_4512,N_5958);
xor U7977 (N_7977,N_5049,N_5811);
and U7978 (N_7978,N_3681,N_3705);
nor U7979 (N_7979,N_5522,N_5815);
nand U7980 (N_7980,N_3845,N_3120);
xnor U7981 (N_7981,N_4690,N_5888);
nor U7982 (N_7982,N_5875,N_3922);
nand U7983 (N_7983,N_5831,N_4207);
or U7984 (N_7984,N_4813,N_4644);
xnor U7985 (N_7985,N_4325,N_3962);
xor U7986 (N_7986,N_3303,N_4888);
or U7987 (N_7987,N_3520,N_5854);
nor U7988 (N_7988,N_4393,N_4509);
and U7989 (N_7989,N_5262,N_3322);
or U7990 (N_7990,N_5243,N_4635);
xor U7991 (N_7991,N_4301,N_4430);
nand U7992 (N_7992,N_4171,N_3596);
and U7993 (N_7993,N_5297,N_4030);
and U7994 (N_7994,N_5593,N_5794);
and U7995 (N_7995,N_3179,N_3639);
or U7996 (N_7996,N_4758,N_3467);
nor U7997 (N_7997,N_3077,N_3153);
nand U7998 (N_7998,N_4574,N_4155);
xnor U7999 (N_7999,N_3349,N_4963);
nand U8000 (N_8000,N_5931,N_3651);
xor U8001 (N_8001,N_3143,N_5416);
and U8002 (N_8002,N_4545,N_5933);
and U8003 (N_8003,N_4350,N_5209);
or U8004 (N_8004,N_3268,N_3588);
nor U8005 (N_8005,N_3049,N_4941);
xnor U8006 (N_8006,N_4460,N_4024);
nand U8007 (N_8007,N_5716,N_5761);
xnor U8008 (N_8008,N_3853,N_5987);
and U8009 (N_8009,N_5646,N_5128);
nand U8010 (N_8010,N_3113,N_5968);
and U8011 (N_8011,N_3625,N_3101);
nor U8012 (N_8012,N_5881,N_3823);
and U8013 (N_8013,N_3935,N_3026);
and U8014 (N_8014,N_3585,N_5369);
and U8015 (N_8015,N_5810,N_5224);
nor U8016 (N_8016,N_5115,N_3181);
and U8017 (N_8017,N_5365,N_4505);
nor U8018 (N_8018,N_5990,N_4107);
nand U8019 (N_8019,N_5885,N_3114);
nor U8020 (N_8020,N_3810,N_5814);
nand U8021 (N_8021,N_4432,N_3644);
nor U8022 (N_8022,N_5148,N_5811);
or U8023 (N_8023,N_5063,N_4085);
or U8024 (N_8024,N_4404,N_5621);
or U8025 (N_8025,N_4553,N_3036);
and U8026 (N_8026,N_3801,N_5754);
xor U8027 (N_8027,N_5377,N_5302);
and U8028 (N_8028,N_5928,N_3971);
xnor U8029 (N_8029,N_4297,N_3317);
nand U8030 (N_8030,N_5647,N_4215);
nor U8031 (N_8031,N_4969,N_4665);
xor U8032 (N_8032,N_4502,N_3189);
nor U8033 (N_8033,N_4871,N_5179);
xnor U8034 (N_8034,N_3010,N_4082);
and U8035 (N_8035,N_5346,N_5978);
nand U8036 (N_8036,N_4343,N_4098);
xnor U8037 (N_8037,N_3431,N_4190);
or U8038 (N_8038,N_5740,N_3466);
and U8039 (N_8039,N_5540,N_4375);
nor U8040 (N_8040,N_3433,N_5703);
nand U8041 (N_8041,N_5234,N_4823);
xnor U8042 (N_8042,N_4063,N_5999);
or U8043 (N_8043,N_3059,N_3405);
xor U8044 (N_8044,N_5228,N_5515);
nor U8045 (N_8045,N_5125,N_5526);
or U8046 (N_8046,N_4779,N_4277);
xor U8047 (N_8047,N_5391,N_5077);
and U8048 (N_8048,N_4349,N_3630);
or U8049 (N_8049,N_5546,N_4869);
or U8050 (N_8050,N_4052,N_3945);
nand U8051 (N_8051,N_4411,N_3518);
xnor U8052 (N_8052,N_5765,N_4162);
nand U8053 (N_8053,N_5660,N_4098);
nand U8054 (N_8054,N_4413,N_3564);
or U8055 (N_8055,N_4652,N_5146);
nor U8056 (N_8056,N_5514,N_4240);
or U8057 (N_8057,N_4249,N_5211);
nand U8058 (N_8058,N_5304,N_3519);
or U8059 (N_8059,N_4740,N_3938);
and U8060 (N_8060,N_4208,N_4191);
or U8061 (N_8061,N_4287,N_5862);
and U8062 (N_8062,N_4338,N_4549);
nor U8063 (N_8063,N_4653,N_5317);
nand U8064 (N_8064,N_4547,N_4983);
or U8065 (N_8065,N_5194,N_4644);
nor U8066 (N_8066,N_5285,N_3502);
nand U8067 (N_8067,N_3225,N_4463);
xor U8068 (N_8068,N_3574,N_4814);
xnor U8069 (N_8069,N_4818,N_5189);
and U8070 (N_8070,N_5928,N_3181);
nand U8071 (N_8071,N_3916,N_4244);
nor U8072 (N_8072,N_5466,N_3176);
nand U8073 (N_8073,N_3674,N_3715);
or U8074 (N_8074,N_4548,N_4975);
xor U8075 (N_8075,N_4352,N_4835);
nand U8076 (N_8076,N_3117,N_5953);
or U8077 (N_8077,N_3248,N_4495);
and U8078 (N_8078,N_3388,N_3807);
xnor U8079 (N_8079,N_4747,N_5258);
xor U8080 (N_8080,N_3036,N_4074);
nand U8081 (N_8081,N_5783,N_4441);
nor U8082 (N_8082,N_5999,N_5852);
and U8083 (N_8083,N_5711,N_5562);
and U8084 (N_8084,N_4032,N_4343);
xor U8085 (N_8085,N_3319,N_3582);
nand U8086 (N_8086,N_5760,N_4612);
or U8087 (N_8087,N_5476,N_5607);
nor U8088 (N_8088,N_5330,N_4731);
nand U8089 (N_8089,N_5717,N_5795);
nand U8090 (N_8090,N_4660,N_4375);
nand U8091 (N_8091,N_5634,N_4430);
nor U8092 (N_8092,N_5306,N_3174);
nand U8093 (N_8093,N_4607,N_3001);
xor U8094 (N_8094,N_5390,N_3504);
nor U8095 (N_8095,N_4592,N_3328);
nand U8096 (N_8096,N_4510,N_4951);
nor U8097 (N_8097,N_4242,N_3463);
nand U8098 (N_8098,N_5472,N_5937);
or U8099 (N_8099,N_4105,N_4089);
nor U8100 (N_8100,N_4673,N_3051);
and U8101 (N_8101,N_4974,N_5398);
nor U8102 (N_8102,N_4962,N_3918);
xnor U8103 (N_8103,N_3958,N_4051);
nor U8104 (N_8104,N_4244,N_4856);
nand U8105 (N_8105,N_3585,N_4107);
or U8106 (N_8106,N_3821,N_3682);
and U8107 (N_8107,N_3305,N_3099);
and U8108 (N_8108,N_5925,N_3071);
xor U8109 (N_8109,N_5926,N_3256);
nand U8110 (N_8110,N_3399,N_3934);
xor U8111 (N_8111,N_3569,N_5862);
xor U8112 (N_8112,N_5691,N_4254);
or U8113 (N_8113,N_3630,N_4135);
and U8114 (N_8114,N_5317,N_4274);
xnor U8115 (N_8115,N_3141,N_5461);
xor U8116 (N_8116,N_4259,N_5012);
nor U8117 (N_8117,N_5791,N_3880);
and U8118 (N_8118,N_5851,N_3628);
and U8119 (N_8119,N_4145,N_3264);
xnor U8120 (N_8120,N_3688,N_4607);
nor U8121 (N_8121,N_4516,N_3547);
xor U8122 (N_8122,N_3775,N_4357);
xor U8123 (N_8123,N_3372,N_4443);
nand U8124 (N_8124,N_5815,N_3808);
xnor U8125 (N_8125,N_3571,N_4619);
and U8126 (N_8126,N_4313,N_3495);
nand U8127 (N_8127,N_5164,N_5631);
or U8128 (N_8128,N_3849,N_4916);
nor U8129 (N_8129,N_5856,N_5731);
nor U8130 (N_8130,N_4976,N_5340);
or U8131 (N_8131,N_4594,N_4800);
nand U8132 (N_8132,N_5427,N_5751);
nor U8133 (N_8133,N_4135,N_5144);
or U8134 (N_8134,N_3141,N_4353);
xor U8135 (N_8135,N_3354,N_3112);
or U8136 (N_8136,N_3272,N_4312);
nand U8137 (N_8137,N_5337,N_3430);
nor U8138 (N_8138,N_5719,N_3470);
or U8139 (N_8139,N_5594,N_5940);
xor U8140 (N_8140,N_3671,N_3107);
nand U8141 (N_8141,N_3458,N_3368);
or U8142 (N_8142,N_5463,N_5055);
nand U8143 (N_8143,N_5754,N_5589);
and U8144 (N_8144,N_3119,N_4228);
nor U8145 (N_8145,N_4409,N_5111);
xor U8146 (N_8146,N_4280,N_3180);
nor U8147 (N_8147,N_3863,N_3914);
or U8148 (N_8148,N_3770,N_3735);
xnor U8149 (N_8149,N_5163,N_4216);
nand U8150 (N_8150,N_5447,N_5548);
nand U8151 (N_8151,N_5378,N_4886);
xor U8152 (N_8152,N_3187,N_4779);
xnor U8153 (N_8153,N_4802,N_3466);
and U8154 (N_8154,N_4253,N_5848);
and U8155 (N_8155,N_4530,N_3813);
nand U8156 (N_8156,N_3378,N_4623);
nor U8157 (N_8157,N_3371,N_4090);
and U8158 (N_8158,N_3574,N_5199);
nor U8159 (N_8159,N_3291,N_5311);
nor U8160 (N_8160,N_4678,N_4791);
nand U8161 (N_8161,N_3543,N_3370);
xnor U8162 (N_8162,N_4306,N_3078);
nor U8163 (N_8163,N_3488,N_4115);
or U8164 (N_8164,N_5094,N_4765);
and U8165 (N_8165,N_5904,N_5035);
nand U8166 (N_8166,N_4923,N_3113);
or U8167 (N_8167,N_3786,N_3960);
nor U8168 (N_8168,N_3166,N_3042);
and U8169 (N_8169,N_5696,N_3853);
xnor U8170 (N_8170,N_5565,N_3776);
nor U8171 (N_8171,N_5526,N_3555);
nand U8172 (N_8172,N_3131,N_4850);
xnor U8173 (N_8173,N_3397,N_3067);
and U8174 (N_8174,N_3630,N_4703);
or U8175 (N_8175,N_4785,N_3444);
nor U8176 (N_8176,N_4236,N_3900);
nand U8177 (N_8177,N_3454,N_3371);
nor U8178 (N_8178,N_3881,N_4367);
and U8179 (N_8179,N_3169,N_3981);
and U8180 (N_8180,N_4413,N_3227);
nor U8181 (N_8181,N_5956,N_3945);
and U8182 (N_8182,N_4699,N_5217);
nand U8183 (N_8183,N_5337,N_4886);
or U8184 (N_8184,N_5643,N_4204);
and U8185 (N_8185,N_4454,N_4729);
and U8186 (N_8186,N_4118,N_5919);
nand U8187 (N_8187,N_4402,N_5171);
and U8188 (N_8188,N_4199,N_4328);
xor U8189 (N_8189,N_5918,N_4836);
nor U8190 (N_8190,N_4734,N_5172);
and U8191 (N_8191,N_5824,N_3501);
or U8192 (N_8192,N_3109,N_5424);
or U8193 (N_8193,N_5206,N_5711);
and U8194 (N_8194,N_5898,N_5496);
xor U8195 (N_8195,N_3351,N_5314);
and U8196 (N_8196,N_5213,N_4496);
or U8197 (N_8197,N_3606,N_3871);
nor U8198 (N_8198,N_4131,N_3242);
or U8199 (N_8199,N_4368,N_3246);
and U8200 (N_8200,N_4579,N_4029);
or U8201 (N_8201,N_4247,N_4325);
nor U8202 (N_8202,N_4719,N_5633);
nand U8203 (N_8203,N_5999,N_5748);
or U8204 (N_8204,N_3261,N_4060);
or U8205 (N_8205,N_3300,N_3308);
nor U8206 (N_8206,N_3586,N_5840);
and U8207 (N_8207,N_4726,N_4091);
nor U8208 (N_8208,N_4792,N_5601);
nand U8209 (N_8209,N_3682,N_4445);
or U8210 (N_8210,N_3187,N_5192);
or U8211 (N_8211,N_3174,N_5051);
nor U8212 (N_8212,N_4050,N_4092);
and U8213 (N_8213,N_4166,N_3613);
and U8214 (N_8214,N_4355,N_5940);
xnor U8215 (N_8215,N_5737,N_4188);
and U8216 (N_8216,N_4453,N_4536);
and U8217 (N_8217,N_5739,N_5241);
nor U8218 (N_8218,N_3483,N_4215);
xnor U8219 (N_8219,N_5840,N_4437);
and U8220 (N_8220,N_5129,N_4739);
nor U8221 (N_8221,N_3054,N_5195);
nand U8222 (N_8222,N_5243,N_5452);
xnor U8223 (N_8223,N_4619,N_5582);
nor U8224 (N_8224,N_5781,N_4475);
or U8225 (N_8225,N_3560,N_5050);
or U8226 (N_8226,N_3175,N_3124);
or U8227 (N_8227,N_5364,N_4818);
xor U8228 (N_8228,N_4718,N_5900);
and U8229 (N_8229,N_5514,N_3950);
xor U8230 (N_8230,N_4091,N_5412);
nor U8231 (N_8231,N_5007,N_3145);
xnor U8232 (N_8232,N_4622,N_5445);
nand U8233 (N_8233,N_4997,N_4147);
or U8234 (N_8234,N_4659,N_4874);
xor U8235 (N_8235,N_4848,N_3428);
and U8236 (N_8236,N_4483,N_4251);
xnor U8237 (N_8237,N_5217,N_5461);
or U8238 (N_8238,N_4278,N_4609);
nand U8239 (N_8239,N_5962,N_5704);
or U8240 (N_8240,N_3842,N_4206);
or U8241 (N_8241,N_4663,N_4778);
nand U8242 (N_8242,N_3917,N_4570);
nor U8243 (N_8243,N_3030,N_5223);
or U8244 (N_8244,N_5937,N_5011);
nor U8245 (N_8245,N_5199,N_3932);
or U8246 (N_8246,N_4942,N_5690);
or U8247 (N_8247,N_4953,N_4839);
xor U8248 (N_8248,N_4499,N_5608);
xor U8249 (N_8249,N_4287,N_4143);
nor U8250 (N_8250,N_5720,N_3376);
or U8251 (N_8251,N_5909,N_3905);
nand U8252 (N_8252,N_3610,N_4520);
xnor U8253 (N_8253,N_3095,N_4283);
nand U8254 (N_8254,N_5937,N_5202);
nor U8255 (N_8255,N_3318,N_5505);
nor U8256 (N_8256,N_5525,N_5662);
and U8257 (N_8257,N_3623,N_3311);
or U8258 (N_8258,N_4039,N_4095);
nand U8259 (N_8259,N_3044,N_3094);
xor U8260 (N_8260,N_3917,N_3185);
and U8261 (N_8261,N_4868,N_4497);
nand U8262 (N_8262,N_3539,N_4348);
xor U8263 (N_8263,N_5046,N_3421);
or U8264 (N_8264,N_4086,N_4353);
xnor U8265 (N_8265,N_4645,N_3499);
and U8266 (N_8266,N_3675,N_4936);
or U8267 (N_8267,N_4501,N_5509);
or U8268 (N_8268,N_4485,N_4745);
nand U8269 (N_8269,N_5307,N_4004);
or U8270 (N_8270,N_4621,N_5666);
nor U8271 (N_8271,N_5751,N_3857);
and U8272 (N_8272,N_5788,N_5204);
xor U8273 (N_8273,N_4850,N_5002);
nor U8274 (N_8274,N_4169,N_4441);
xor U8275 (N_8275,N_4104,N_3663);
or U8276 (N_8276,N_5432,N_3377);
nand U8277 (N_8277,N_5261,N_3654);
nor U8278 (N_8278,N_3373,N_3813);
nand U8279 (N_8279,N_3557,N_4391);
nor U8280 (N_8280,N_4237,N_5904);
nand U8281 (N_8281,N_4502,N_3837);
nand U8282 (N_8282,N_3410,N_4514);
and U8283 (N_8283,N_5583,N_4948);
or U8284 (N_8284,N_3122,N_4125);
and U8285 (N_8285,N_4486,N_4265);
nor U8286 (N_8286,N_5406,N_3370);
nor U8287 (N_8287,N_4837,N_5684);
nor U8288 (N_8288,N_3244,N_5453);
and U8289 (N_8289,N_4185,N_5045);
nor U8290 (N_8290,N_5743,N_4217);
nor U8291 (N_8291,N_5814,N_4089);
and U8292 (N_8292,N_3632,N_4026);
and U8293 (N_8293,N_5460,N_4443);
and U8294 (N_8294,N_4347,N_3442);
nand U8295 (N_8295,N_3112,N_3808);
xor U8296 (N_8296,N_5133,N_3699);
nor U8297 (N_8297,N_4364,N_5317);
nor U8298 (N_8298,N_4142,N_4876);
or U8299 (N_8299,N_5592,N_4278);
xor U8300 (N_8300,N_3543,N_4456);
nand U8301 (N_8301,N_4755,N_3980);
and U8302 (N_8302,N_3530,N_3876);
xnor U8303 (N_8303,N_3121,N_3537);
and U8304 (N_8304,N_3659,N_4244);
and U8305 (N_8305,N_5387,N_4487);
xnor U8306 (N_8306,N_5885,N_5453);
nand U8307 (N_8307,N_4100,N_4869);
and U8308 (N_8308,N_3630,N_5616);
nor U8309 (N_8309,N_5003,N_5492);
xnor U8310 (N_8310,N_3992,N_3092);
or U8311 (N_8311,N_5472,N_3697);
xnor U8312 (N_8312,N_4822,N_4943);
xnor U8313 (N_8313,N_4348,N_5761);
and U8314 (N_8314,N_4228,N_3383);
and U8315 (N_8315,N_3447,N_4741);
and U8316 (N_8316,N_3498,N_5397);
xnor U8317 (N_8317,N_3285,N_3872);
xnor U8318 (N_8318,N_3214,N_3867);
xor U8319 (N_8319,N_4181,N_5696);
or U8320 (N_8320,N_3567,N_5680);
nor U8321 (N_8321,N_3934,N_4133);
or U8322 (N_8322,N_3502,N_5650);
xor U8323 (N_8323,N_3730,N_4886);
nor U8324 (N_8324,N_3811,N_5930);
nand U8325 (N_8325,N_4101,N_4184);
xor U8326 (N_8326,N_5582,N_4958);
xnor U8327 (N_8327,N_5812,N_4859);
nor U8328 (N_8328,N_4418,N_5532);
nand U8329 (N_8329,N_3560,N_4110);
and U8330 (N_8330,N_5536,N_4975);
nand U8331 (N_8331,N_3583,N_3721);
nand U8332 (N_8332,N_5816,N_5881);
nand U8333 (N_8333,N_3843,N_3967);
nor U8334 (N_8334,N_3716,N_5636);
xor U8335 (N_8335,N_5542,N_5546);
nand U8336 (N_8336,N_3058,N_5233);
nor U8337 (N_8337,N_3955,N_3617);
or U8338 (N_8338,N_5303,N_3514);
and U8339 (N_8339,N_4333,N_4852);
nand U8340 (N_8340,N_4979,N_3140);
nand U8341 (N_8341,N_5063,N_5503);
nor U8342 (N_8342,N_5141,N_4876);
nor U8343 (N_8343,N_5287,N_3813);
nor U8344 (N_8344,N_5887,N_5108);
xor U8345 (N_8345,N_5931,N_5505);
xor U8346 (N_8346,N_4789,N_4085);
or U8347 (N_8347,N_4202,N_5650);
nand U8348 (N_8348,N_4601,N_5325);
or U8349 (N_8349,N_5463,N_4069);
xor U8350 (N_8350,N_4960,N_3589);
and U8351 (N_8351,N_4084,N_4983);
nor U8352 (N_8352,N_5927,N_5856);
and U8353 (N_8353,N_5350,N_4924);
nor U8354 (N_8354,N_4490,N_5491);
nand U8355 (N_8355,N_4465,N_4312);
xnor U8356 (N_8356,N_5760,N_4731);
and U8357 (N_8357,N_3473,N_3349);
nor U8358 (N_8358,N_3799,N_3875);
or U8359 (N_8359,N_4006,N_4260);
and U8360 (N_8360,N_5072,N_3843);
and U8361 (N_8361,N_3256,N_3281);
xor U8362 (N_8362,N_5544,N_3620);
or U8363 (N_8363,N_4520,N_3594);
nor U8364 (N_8364,N_3274,N_4801);
nor U8365 (N_8365,N_5383,N_4231);
nor U8366 (N_8366,N_4193,N_4290);
xor U8367 (N_8367,N_4246,N_3747);
nand U8368 (N_8368,N_5653,N_4001);
xnor U8369 (N_8369,N_4273,N_4684);
xnor U8370 (N_8370,N_4663,N_4828);
nand U8371 (N_8371,N_5777,N_3533);
nor U8372 (N_8372,N_4524,N_5863);
or U8373 (N_8373,N_5364,N_5062);
nor U8374 (N_8374,N_5142,N_4249);
nor U8375 (N_8375,N_4712,N_3899);
or U8376 (N_8376,N_3793,N_5816);
or U8377 (N_8377,N_3365,N_5773);
xnor U8378 (N_8378,N_5967,N_3559);
or U8379 (N_8379,N_4203,N_3198);
or U8380 (N_8380,N_3227,N_5133);
nand U8381 (N_8381,N_4338,N_4873);
nor U8382 (N_8382,N_5096,N_3643);
nand U8383 (N_8383,N_5739,N_3141);
nand U8384 (N_8384,N_3667,N_3468);
nor U8385 (N_8385,N_4544,N_5885);
nor U8386 (N_8386,N_5426,N_4530);
or U8387 (N_8387,N_5446,N_5530);
nor U8388 (N_8388,N_3880,N_4344);
and U8389 (N_8389,N_5972,N_5644);
or U8390 (N_8390,N_3136,N_4571);
and U8391 (N_8391,N_4273,N_4235);
or U8392 (N_8392,N_3863,N_3626);
or U8393 (N_8393,N_4720,N_5693);
xnor U8394 (N_8394,N_4285,N_3671);
xnor U8395 (N_8395,N_3944,N_3257);
or U8396 (N_8396,N_3074,N_3471);
or U8397 (N_8397,N_5292,N_4683);
or U8398 (N_8398,N_4580,N_4386);
xor U8399 (N_8399,N_5950,N_5979);
xnor U8400 (N_8400,N_3531,N_4198);
nand U8401 (N_8401,N_4613,N_5931);
nor U8402 (N_8402,N_5855,N_4328);
and U8403 (N_8403,N_4545,N_5763);
nor U8404 (N_8404,N_3386,N_5157);
xnor U8405 (N_8405,N_3781,N_5700);
nor U8406 (N_8406,N_3279,N_4161);
and U8407 (N_8407,N_3494,N_4985);
nor U8408 (N_8408,N_5963,N_4346);
xor U8409 (N_8409,N_5504,N_3865);
xor U8410 (N_8410,N_4621,N_5791);
or U8411 (N_8411,N_5645,N_3469);
nor U8412 (N_8412,N_4259,N_5666);
xnor U8413 (N_8413,N_3964,N_4386);
and U8414 (N_8414,N_4623,N_4749);
and U8415 (N_8415,N_4455,N_3528);
or U8416 (N_8416,N_3062,N_3187);
or U8417 (N_8417,N_4008,N_3582);
nand U8418 (N_8418,N_4830,N_3461);
nor U8419 (N_8419,N_4717,N_4444);
or U8420 (N_8420,N_5491,N_5159);
and U8421 (N_8421,N_3603,N_4313);
and U8422 (N_8422,N_4721,N_3233);
or U8423 (N_8423,N_3820,N_5486);
and U8424 (N_8424,N_4303,N_4198);
xnor U8425 (N_8425,N_4211,N_4515);
and U8426 (N_8426,N_3917,N_4652);
or U8427 (N_8427,N_3799,N_3071);
xor U8428 (N_8428,N_4002,N_3867);
and U8429 (N_8429,N_3498,N_3314);
nor U8430 (N_8430,N_4688,N_4462);
and U8431 (N_8431,N_5178,N_5906);
or U8432 (N_8432,N_3928,N_5931);
xor U8433 (N_8433,N_4388,N_3312);
nand U8434 (N_8434,N_5184,N_4890);
xor U8435 (N_8435,N_4776,N_4260);
xor U8436 (N_8436,N_5984,N_4898);
or U8437 (N_8437,N_3557,N_3071);
nor U8438 (N_8438,N_4508,N_4278);
nand U8439 (N_8439,N_5276,N_5740);
nand U8440 (N_8440,N_5528,N_4311);
or U8441 (N_8441,N_5133,N_5745);
xor U8442 (N_8442,N_3813,N_4833);
and U8443 (N_8443,N_4737,N_4779);
nand U8444 (N_8444,N_3385,N_4677);
or U8445 (N_8445,N_5905,N_3261);
nand U8446 (N_8446,N_3491,N_3576);
xnor U8447 (N_8447,N_5074,N_4036);
nor U8448 (N_8448,N_5512,N_4279);
xnor U8449 (N_8449,N_4842,N_5426);
nand U8450 (N_8450,N_4737,N_5901);
xnor U8451 (N_8451,N_4810,N_4548);
or U8452 (N_8452,N_3916,N_4548);
and U8453 (N_8453,N_5758,N_3862);
and U8454 (N_8454,N_3304,N_5637);
xor U8455 (N_8455,N_3789,N_5200);
nor U8456 (N_8456,N_3812,N_4998);
nor U8457 (N_8457,N_4264,N_3829);
xnor U8458 (N_8458,N_3916,N_3879);
nor U8459 (N_8459,N_3570,N_4117);
or U8460 (N_8460,N_3796,N_4645);
nor U8461 (N_8461,N_4642,N_4476);
or U8462 (N_8462,N_3547,N_3777);
nand U8463 (N_8463,N_3650,N_4255);
nor U8464 (N_8464,N_3793,N_5651);
nor U8465 (N_8465,N_5115,N_4033);
xor U8466 (N_8466,N_4529,N_3697);
nand U8467 (N_8467,N_4836,N_3617);
xnor U8468 (N_8468,N_5296,N_5111);
and U8469 (N_8469,N_3730,N_3894);
and U8470 (N_8470,N_3957,N_5353);
or U8471 (N_8471,N_3823,N_4863);
or U8472 (N_8472,N_4176,N_5991);
and U8473 (N_8473,N_3940,N_4234);
and U8474 (N_8474,N_3057,N_4932);
xnor U8475 (N_8475,N_5832,N_5788);
xnor U8476 (N_8476,N_5984,N_3777);
xor U8477 (N_8477,N_3088,N_3415);
nand U8478 (N_8478,N_3165,N_4017);
or U8479 (N_8479,N_3855,N_3670);
nand U8480 (N_8480,N_3273,N_3794);
and U8481 (N_8481,N_4751,N_5587);
nor U8482 (N_8482,N_5476,N_3619);
nor U8483 (N_8483,N_5689,N_3047);
or U8484 (N_8484,N_3788,N_4542);
nand U8485 (N_8485,N_3646,N_5259);
nor U8486 (N_8486,N_5253,N_4679);
nor U8487 (N_8487,N_4767,N_4915);
nand U8488 (N_8488,N_5223,N_4695);
or U8489 (N_8489,N_4635,N_5879);
xnor U8490 (N_8490,N_3243,N_4521);
nor U8491 (N_8491,N_3453,N_4190);
xnor U8492 (N_8492,N_4709,N_5694);
or U8493 (N_8493,N_3457,N_4702);
or U8494 (N_8494,N_3971,N_4352);
xor U8495 (N_8495,N_3401,N_5041);
or U8496 (N_8496,N_5506,N_4373);
xor U8497 (N_8497,N_4132,N_3260);
xnor U8498 (N_8498,N_3653,N_3964);
nor U8499 (N_8499,N_3378,N_5817);
and U8500 (N_8500,N_5172,N_4349);
nor U8501 (N_8501,N_5462,N_4721);
nor U8502 (N_8502,N_4221,N_5196);
nand U8503 (N_8503,N_5723,N_5663);
nand U8504 (N_8504,N_5493,N_3671);
or U8505 (N_8505,N_4331,N_4201);
and U8506 (N_8506,N_5104,N_3877);
nor U8507 (N_8507,N_3465,N_3525);
and U8508 (N_8508,N_5827,N_4429);
xnor U8509 (N_8509,N_4786,N_5817);
or U8510 (N_8510,N_4137,N_4742);
nand U8511 (N_8511,N_5176,N_5883);
xor U8512 (N_8512,N_3000,N_3513);
or U8513 (N_8513,N_4137,N_4355);
and U8514 (N_8514,N_5498,N_5605);
or U8515 (N_8515,N_4200,N_4278);
or U8516 (N_8516,N_3934,N_3753);
nor U8517 (N_8517,N_5480,N_3451);
xor U8518 (N_8518,N_3070,N_3269);
nor U8519 (N_8519,N_3819,N_4826);
nor U8520 (N_8520,N_5869,N_5535);
xnor U8521 (N_8521,N_4640,N_4725);
nor U8522 (N_8522,N_5505,N_3467);
nand U8523 (N_8523,N_3532,N_5489);
or U8524 (N_8524,N_3224,N_3190);
or U8525 (N_8525,N_4033,N_3513);
and U8526 (N_8526,N_3163,N_5876);
or U8527 (N_8527,N_5810,N_4595);
nand U8528 (N_8528,N_4904,N_3991);
and U8529 (N_8529,N_5278,N_3631);
nor U8530 (N_8530,N_4728,N_5020);
nand U8531 (N_8531,N_3932,N_5307);
xnor U8532 (N_8532,N_5273,N_5071);
or U8533 (N_8533,N_3876,N_4439);
and U8534 (N_8534,N_4354,N_5972);
or U8535 (N_8535,N_5296,N_4010);
and U8536 (N_8536,N_3999,N_5889);
or U8537 (N_8537,N_4109,N_4848);
nand U8538 (N_8538,N_4098,N_3802);
xor U8539 (N_8539,N_4730,N_5270);
xnor U8540 (N_8540,N_5094,N_4311);
nand U8541 (N_8541,N_3905,N_3720);
or U8542 (N_8542,N_5835,N_3733);
nand U8543 (N_8543,N_5103,N_3879);
xnor U8544 (N_8544,N_5675,N_4548);
nor U8545 (N_8545,N_3157,N_4689);
and U8546 (N_8546,N_3191,N_3148);
nand U8547 (N_8547,N_3029,N_5921);
xnor U8548 (N_8548,N_4061,N_4749);
and U8549 (N_8549,N_3567,N_3515);
xnor U8550 (N_8550,N_3174,N_4461);
and U8551 (N_8551,N_5836,N_4465);
nor U8552 (N_8552,N_3175,N_3311);
nor U8553 (N_8553,N_4136,N_5534);
nand U8554 (N_8554,N_3613,N_4163);
xnor U8555 (N_8555,N_3515,N_3460);
and U8556 (N_8556,N_5888,N_5999);
nand U8557 (N_8557,N_5340,N_5102);
xor U8558 (N_8558,N_5068,N_4433);
nor U8559 (N_8559,N_5324,N_3568);
or U8560 (N_8560,N_5281,N_4323);
nand U8561 (N_8561,N_3054,N_4930);
nor U8562 (N_8562,N_3811,N_5742);
or U8563 (N_8563,N_5754,N_5222);
xor U8564 (N_8564,N_3525,N_5301);
and U8565 (N_8565,N_5092,N_5136);
nor U8566 (N_8566,N_3632,N_4386);
xnor U8567 (N_8567,N_3798,N_5169);
nor U8568 (N_8568,N_3806,N_5289);
or U8569 (N_8569,N_3480,N_4561);
nand U8570 (N_8570,N_3409,N_3311);
and U8571 (N_8571,N_3011,N_4805);
xor U8572 (N_8572,N_4405,N_5189);
xnor U8573 (N_8573,N_5129,N_5760);
nor U8574 (N_8574,N_4239,N_5693);
xnor U8575 (N_8575,N_5327,N_5932);
nand U8576 (N_8576,N_3957,N_5853);
or U8577 (N_8577,N_3809,N_4985);
nor U8578 (N_8578,N_3801,N_5817);
and U8579 (N_8579,N_5731,N_3049);
xor U8580 (N_8580,N_4590,N_3080);
nor U8581 (N_8581,N_3081,N_4307);
xor U8582 (N_8582,N_3624,N_3379);
nor U8583 (N_8583,N_5932,N_4697);
xnor U8584 (N_8584,N_3985,N_5850);
and U8585 (N_8585,N_3313,N_4327);
xor U8586 (N_8586,N_4958,N_5212);
and U8587 (N_8587,N_3459,N_3600);
nor U8588 (N_8588,N_5095,N_4807);
or U8589 (N_8589,N_5642,N_3273);
xor U8590 (N_8590,N_3151,N_5056);
xnor U8591 (N_8591,N_3350,N_5072);
nor U8592 (N_8592,N_5231,N_4193);
or U8593 (N_8593,N_4606,N_5567);
nor U8594 (N_8594,N_4988,N_3606);
or U8595 (N_8595,N_3213,N_5017);
xnor U8596 (N_8596,N_3072,N_4242);
and U8597 (N_8597,N_5389,N_3327);
nand U8598 (N_8598,N_3528,N_3917);
nor U8599 (N_8599,N_3768,N_5604);
or U8600 (N_8600,N_3269,N_5903);
nand U8601 (N_8601,N_3245,N_4481);
and U8602 (N_8602,N_5467,N_5526);
and U8603 (N_8603,N_4653,N_5187);
nor U8604 (N_8604,N_3421,N_4522);
nor U8605 (N_8605,N_3709,N_4323);
xor U8606 (N_8606,N_5069,N_5412);
xor U8607 (N_8607,N_3371,N_4977);
nor U8608 (N_8608,N_4524,N_4520);
xnor U8609 (N_8609,N_4151,N_5168);
nor U8610 (N_8610,N_5579,N_3480);
or U8611 (N_8611,N_3908,N_4110);
nor U8612 (N_8612,N_3645,N_4270);
nand U8613 (N_8613,N_5805,N_4187);
nor U8614 (N_8614,N_5948,N_5149);
or U8615 (N_8615,N_3969,N_5278);
or U8616 (N_8616,N_4245,N_3918);
nand U8617 (N_8617,N_3469,N_4965);
nand U8618 (N_8618,N_4133,N_5116);
and U8619 (N_8619,N_3792,N_5541);
nand U8620 (N_8620,N_4808,N_3567);
xor U8621 (N_8621,N_5995,N_3348);
nand U8622 (N_8622,N_3964,N_5573);
or U8623 (N_8623,N_3340,N_5693);
xnor U8624 (N_8624,N_3361,N_3077);
and U8625 (N_8625,N_4569,N_3757);
or U8626 (N_8626,N_3495,N_5295);
nor U8627 (N_8627,N_4625,N_5958);
and U8628 (N_8628,N_3736,N_4429);
nand U8629 (N_8629,N_3601,N_4512);
or U8630 (N_8630,N_4106,N_5694);
nand U8631 (N_8631,N_5262,N_5963);
or U8632 (N_8632,N_5753,N_4714);
nor U8633 (N_8633,N_4787,N_5699);
xor U8634 (N_8634,N_4707,N_5248);
or U8635 (N_8635,N_3729,N_5424);
and U8636 (N_8636,N_5685,N_4070);
and U8637 (N_8637,N_4776,N_4009);
nor U8638 (N_8638,N_4657,N_5149);
xnor U8639 (N_8639,N_3005,N_3583);
nand U8640 (N_8640,N_5637,N_5943);
and U8641 (N_8641,N_4947,N_5908);
xor U8642 (N_8642,N_4582,N_4889);
and U8643 (N_8643,N_4599,N_4746);
xor U8644 (N_8644,N_4226,N_5669);
nor U8645 (N_8645,N_3252,N_5033);
and U8646 (N_8646,N_4191,N_5941);
nand U8647 (N_8647,N_3910,N_5420);
nor U8648 (N_8648,N_3363,N_4627);
or U8649 (N_8649,N_3104,N_4461);
xnor U8650 (N_8650,N_5573,N_3409);
nand U8651 (N_8651,N_5019,N_4459);
xnor U8652 (N_8652,N_5053,N_3045);
nor U8653 (N_8653,N_4491,N_5876);
or U8654 (N_8654,N_5663,N_5248);
nand U8655 (N_8655,N_3624,N_4223);
nand U8656 (N_8656,N_4478,N_5485);
and U8657 (N_8657,N_3830,N_5855);
nand U8658 (N_8658,N_5761,N_4148);
and U8659 (N_8659,N_4741,N_3286);
or U8660 (N_8660,N_4702,N_4038);
nor U8661 (N_8661,N_5854,N_5209);
nor U8662 (N_8662,N_5658,N_3235);
or U8663 (N_8663,N_4791,N_3013);
xor U8664 (N_8664,N_4455,N_3698);
nor U8665 (N_8665,N_3803,N_4364);
and U8666 (N_8666,N_5633,N_4560);
or U8667 (N_8667,N_3120,N_4058);
xnor U8668 (N_8668,N_4543,N_5196);
nand U8669 (N_8669,N_5539,N_5093);
nor U8670 (N_8670,N_3217,N_5416);
and U8671 (N_8671,N_3041,N_3885);
xnor U8672 (N_8672,N_3641,N_3819);
nand U8673 (N_8673,N_5316,N_3745);
and U8674 (N_8674,N_4186,N_3723);
or U8675 (N_8675,N_3481,N_4700);
and U8676 (N_8676,N_5462,N_3244);
nand U8677 (N_8677,N_3453,N_5620);
nor U8678 (N_8678,N_5651,N_3708);
nor U8679 (N_8679,N_3328,N_5752);
nand U8680 (N_8680,N_5990,N_3666);
or U8681 (N_8681,N_4360,N_5405);
nand U8682 (N_8682,N_4274,N_3464);
and U8683 (N_8683,N_4457,N_3124);
nand U8684 (N_8684,N_4397,N_3150);
or U8685 (N_8685,N_3882,N_5334);
nor U8686 (N_8686,N_4931,N_4540);
or U8687 (N_8687,N_5632,N_4158);
xor U8688 (N_8688,N_5685,N_3733);
xnor U8689 (N_8689,N_4501,N_5318);
or U8690 (N_8690,N_5407,N_4960);
and U8691 (N_8691,N_4073,N_5409);
or U8692 (N_8692,N_5755,N_3716);
nand U8693 (N_8693,N_4488,N_5778);
or U8694 (N_8694,N_5629,N_3869);
xor U8695 (N_8695,N_5159,N_4020);
nand U8696 (N_8696,N_4519,N_3018);
and U8697 (N_8697,N_5756,N_4392);
nor U8698 (N_8698,N_3032,N_3490);
nand U8699 (N_8699,N_3140,N_4779);
or U8700 (N_8700,N_5071,N_5446);
nand U8701 (N_8701,N_5284,N_5385);
xnor U8702 (N_8702,N_4148,N_5695);
and U8703 (N_8703,N_5801,N_5131);
nor U8704 (N_8704,N_3546,N_5191);
or U8705 (N_8705,N_3837,N_3910);
or U8706 (N_8706,N_3321,N_3360);
and U8707 (N_8707,N_4348,N_4718);
nand U8708 (N_8708,N_4340,N_3255);
xnor U8709 (N_8709,N_4962,N_4211);
xnor U8710 (N_8710,N_3310,N_5498);
nand U8711 (N_8711,N_5619,N_4705);
nand U8712 (N_8712,N_5558,N_5182);
nor U8713 (N_8713,N_3230,N_5537);
nand U8714 (N_8714,N_4496,N_5335);
and U8715 (N_8715,N_4661,N_4259);
nand U8716 (N_8716,N_3135,N_5369);
and U8717 (N_8717,N_4436,N_3648);
and U8718 (N_8718,N_4614,N_5000);
and U8719 (N_8719,N_4832,N_5548);
nand U8720 (N_8720,N_5354,N_4067);
nand U8721 (N_8721,N_4509,N_5918);
nand U8722 (N_8722,N_4439,N_4762);
and U8723 (N_8723,N_4274,N_3873);
or U8724 (N_8724,N_4550,N_4424);
xor U8725 (N_8725,N_4798,N_4926);
xor U8726 (N_8726,N_5281,N_3316);
nand U8727 (N_8727,N_5716,N_3689);
xnor U8728 (N_8728,N_3318,N_5186);
nor U8729 (N_8729,N_5936,N_5307);
or U8730 (N_8730,N_3975,N_3138);
xnor U8731 (N_8731,N_4263,N_5814);
nand U8732 (N_8732,N_5171,N_3777);
nor U8733 (N_8733,N_5077,N_5697);
and U8734 (N_8734,N_5057,N_3886);
nand U8735 (N_8735,N_3317,N_5596);
or U8736 (N_8736,N_5512,N_3583);
or U8737 (N_8737,N_5676,N_5327);
nand U8738 (N_8738,N_3011,N_5705);
or U8739 (N_8739,N_5856,N_4158);
nand U8740 (N_8740,N_4030,N_5104);
and U8741 (N_8741,N_5954,N_3738);
and U8742 (N_8742,N_4974,N_3141);
or U8743 (N_8743,N_4982,N_5709);
nor U8744 (N_8744,N_5374,N_5733);
and U8745 (N_8745,N_5975,N_5520);
and U8746 (N_8746,N_5039,N_3118);
nor U8747 (N_8747,N_4730,N_3003);
nor U8748 (N_8748,N_3670,N_5482);
and U8749 (N_8749,N_3885,N_5166);
nor U8750 (N_8750,N_4342,N_3862);
or U8751 (N_8751,N_5381,N_4555);
nor U8752 (N_8752,N_5181,N_3008);
nand U8753 (N_8753,N_5831,N_3060);
nor U8754 (N_8754,N_5930,N_3944);
and U8755 (N_8755,N_3597,N_5778);
nor U8756 (N_8756,N_5605,N_5995);
xor U8757 (N_8757,N_3582,N_5284);
nand U8758 (N_8758,N_4831,N_4604);
xnor U8759 (N_8759,N_4298,N_3774);
nor U8760 (N_8760,N_5219,N_5108);
and U8761 (N_8761,N_4903,N_4566);
xnor U8762 (N_8762,N_3986,N_4001);
and U8763 (N_8763,N_3493,N_5154);
or U8764 (N_8764,N_4924,N_3981);
xor U8765 (N_8765,N_4031,N_4261);
nand U8766 (N_8766,N_5836,N_4827);
xnor U8767 (N_8767,N_4728,N_4332);
and U8768 (N_8768,N_4704,N_4894);
and U8769 (N_8769,N_5736,N_5144);
nand U8770 (N_8770,N_4580,N_4697);
nor U8771 (N_8771,N_5178,N_4060);
nand U8772 (N_8772,N_5717,N_5235);
or U8773 (N_8773,N_5014,N_3999);
nand U8774 (N_8774,N_5601,N_5549);
nor U8775 (N_8775,N_5794,N_3812);
nor U8776 (N_8776,N_5833,N_4183);
nor U8777 (N_8777,N_5585,N_5159);
or U8778 (N_8778,N_5280,N_3526);
and U8779 (N_8779,N_5596,N_4653);
xor U8780 (N_8780,N_5884,N_5466);
or U8781 (N_8781,N_4533,N_3368);
and U8782 (N_8782,N_3729,N_5359);
nor U8783 (N_8783,N_3395,N_3887);
xnor U8784 (N_8784,N_3525,N_3780);
nor U8785 (N_8785,N_4398,N_4938);
nand U8786 (N_8786,N_3229,N_4796);
nand U8787 (N_8787,N_5548,N_3704);
nor U8788 (N_8788,N_4182,N_5166);
nand U8789 (N_8789,N_4718,N_4006);
nand U8790 (N_8790,N_4482,N_3295);
or U8791 (N_8791,N_4578,N_4348);
xnor U8792 (N_8792,N_4815,N_5826);
nor U8793 (N_8793,N_3014,N_5596);
nand U8794 (N_8794,N_5835,N_5440);
nand U8795 (N_8795,N_3284,N_4016);
or U8796 (N_8796,N_5508,N_3605);
or U8797 (N_8797,N_3503,N_3147);
xnor U8798 (N_8798,N_4299,N_5114);
nand U8799 (N_8799,N_3622,N_3779);
or U8800 (N_8800,N_4396,N_5829);
and U8801 (N_8801,N_5707,N_5899);
xnor U8802 (N_8802,N_5658,N_5766);
or U8803 (N_8803,N_3598,N_4175);
nand U8804 (N_8804,N_3000,N_5778);
and U8805 (N_8805,N_5538,N_3299);
or U8806 (N_8806,N_3940,N_4577);
and U8807 (N_8807,N_4539,N_3325);
nor U8808 (N_8808,N_3705,N_3606);
nand U8809 (N_8809,N_3046,N_5491);
nor U8810 (N_8810,N_3672,N_4441);
xnor U8811 (N_8811,N_5844,N_5397);
or U8812 (N_8812,N_3277,N_4434);
or U8813 (N_8813,N_4803,N_5587);
nor U8814 (N_8814,N_3680,N_4006);
or U8815 (N_8815,N_5401,N_4667);
nor U8816 (N_8816,N_3881,N_3915);
and U8817 (N_8817,N_5456,N_3484);
nor U8818 (N_8818,N_4065,N_3876);
or U8819 (N_8819,N_5245,N_4027);
nand U8820 (N_8820,N_3656,N_4644);
nor U8821 (N_8821,N_5300,N_3359);
xor U8822 (N_8822,N_5132,N_4102);
xnor U8823 (N_8823,N_3873,N_4361);
xnor U8824 (N_8824,N_5805,N_5958);
and U8825 (N_8825,N_3166,N_3060);
or U8826 (N_8826,N_3542,N_5825);
and U8827 (N_8827,N_5955,N_4974);
nand U8828 (N_8828,N_5502,N_5489);
nor U8829 (N_8829,N_3105,N_4824);
nor U8830 (N_8830,N_4485,N_3186);
xor U8831 (N_8831,N_4211,N_5120);
and U8832 (N_8832,N_5484,N_4803);
or U8833 (N_8833,N_3440,N_5456);
and U8834 (N_8834,N_4667,N_5971);
nor U8835 (N_8835,N_3223,N_3595);
nand U8836 (N_8836,N_3317,N_5488);
nand U8837 (N_8837,N_3142,N_5648);
nand U8838 (N_8838,N_5922,N_5237);
nor U8839 (N_8839,N_4130,N_3697);
or U8840 (N_8840,N_4340,N_5098);
nand U8841 (N_8841,N_3208,N_3416);
or U8842 (N_8842,N_3059,N_3874);
and U8843 (N_8843,N_4376,N_5004);
or U8844 (N_8844,N_4554,N_4681);
xor U8845 (N_8845,N_3804,N_3631);
and U8846 (N_8846,N_5180,N_4621);
nor U8847 (N_8847,N_5683,N_5583);
nand U8848 (N_8848,N_5783,N_5775);
nand U8849 (N_8849,N_3455,N_5103);
and U8850 (N_8850,N_4372,N_5273);
and U8851 (N_8851,N_3368,N_4583);
nor U8852 (N_8852,N_4778,N_5600);
and U8853 (N_8853,N_3252,N_5693);
or U8854 (N_8854,N_4257,N_3231);
nand U8855 (N_8855,N_5770,N_3974);
nand U8856 (N_8856,N_5308,N_4653);
nor U8857 (N_8857,N_5725,N_4914);
nor U8858 (N_8858,N_3727,N_5222);
nor U8859 (N_8859,N_5648,N_5541);
nand U8860 (N_8860,N_5139,N_5699);
xnor U8861 (N_8861,N_5534,N_3078);
nor U8862 (N_8862,N_3148,N_3249);
nand U8863 (N_8863,N_5988,N_4780);
or U8864 (N_8864,N_3512,N_3341);
nor U8865 (N_8865,N_5137,N_4107);
and U8866 (N_8866,N_3880,N_4321);
nor U8867 (N_8867,N_3246,N_3951);
nor U8868 (N_8868,N_5870,N_5167);
and U8869 (N_8869,N_4330,N_4993);
nand U8870 (N_8870,N_4010,N_4563);
nand U8871 (N_8871,N_3218,N_4045);
xnor U8872 (N_8872,N_5785,N_3555);
and U8873 (N_8873,N_3341,N_5781);
nand U8874 (N_8874,N_5091,N_3386);
xor U8875 (N_8875,N_3974,N_3334);
or U8876 (N_8876,N_5865,N_4748);
or U8877 (N_8877,N_4220,N_3844);
or U8878 (N_8878,N_3484,N_4298);
nor U8879 (N_8879,N_5955,N_5520);
nand U8880 (N_8880,N_4195,N_4304);
nor U8881 (N_8881,N_5796,N_4712);
xnor U8882 (N_8882,N_5518,N_4456);
and U8883 (N_8883,N_3886,N_3171);
nor U8884 (N_8884,N_3690,N_5468);
or U8885 (N_8885,N_3717,N_5037);
xnor U8886 (N_8886,N_5164,N_4762);
and U8887 (N_8887,N_5969,N_3204);
and U8888 (N_8888,N_5494,N_3073);
nand U8889 (N_8889,N_4943,N_4173);
and U8890 (N_8890,N_4154,N_5345);
and U8891 (N_8891,N_5663,N_3104);
nor U8892 (N_8892,N_4198,N_5772);
or U8893 (N_8893,N_4857,N_4628);
nor U8894 (N_8894,N_3891,N_3051);
or U8895 (N_8895,N_4664,N_3152);
nor U8896 (N_8896,N_5766,N_5127);
xor U8897 (N_8897,N_3515,N_5061);
nand U8898 (N_8898,N_3928,N_3717);
and U8899 (N_8899,N_5485,N_4431);
and U8900 (N_8900,N_3903,N_5756);
or U8901 (N_8901,N_5346,N_5204);
xnor U8902 (N_8902,N_3482,N_3322);
nor U8903 (N_8903,N_4313,N_4436);
or U8904 (N_8904,N_4040,N_3811);
xor U8905 (N_8905,N_5675,N_3164);
nor U8906 (N_8906,N_4596,N_3343);
xnor U8907 (N_8907,N_5804,N_3078);
nand U8908 (N_8908,N_5097,N_5159);
xnor U8909 (N_8909,N_5506,N_4472);
or U8910 (N_8910,N_5028,N_4910);
and U8911 (N_8911,N_5217,N_3630);
xor U8912 (N_8912,N_4007,N_4637);
xnor U8913 (N_8913,N_4117,N_5142);
nand U8914 (N_8914,N_5911,N_4380);
xnor U8915 (N_8915,N_4018,N_5985);
nor U8916 (N_8916,N_4191,N_5923);
xor U8917 (N_8917,N_4745,N_5658);
and U8918 (N_8918,N_4248,N_5179);
nor U8919 (N_8919,N_4338,N_5776);
nand U8920 (N_8920,N_5054,N_4294);
nor U8921 (N_8921,N_4594,N_4190);
xor U8922 (N_8922,N_3113,N_3927);
nand U8923 (N_8923,N_3681,N_5005);
nand U8924 (N_8924,N_4032,N_5573);
or U8925 (N_8925,N_5159,N_4337);
nand U8926 (N_8926,N_5101,N_4952);
or U8927 (N_8927,N_3954,N_3141);
nor U8928 (N_8928,N_4059,N_5269);
or U8929 (N_8929,N_3638,N_5325);
nand U8930 (N_8930,N_5717,N_3353);
nand U8931 (N_8931,N_3299,N_5286);
or U8932 (N_8932,N_3383,N_3974);
or U8933 (N_8933,N_5326,N_3758);
or U8934 (N_8934,N_3357,N_3348);
nand U8935 (N_8935,N_5210,N_3747);
xor U8936 (N_8936,N_4779,N_5434);
nor U8937 (N_8937,N_5756,N_4520);
nand U8938 (N_8938,N_4725,N_4502);
or U8939 (N_8939,N_3204,N_5825);
nor U8940 (N_8940,N_4806,N_4862);
or U8941 (N_8941,N_5657,N_3213);
nand U8942 (N_8942,N_3267,N_4448);
nand U8943 (N_8943,N_4829,N_4732);
nor U8944 (N_8944,N_5751,N_5692);
or U8945 (N_8945,N_4138,N_5370);
xnor U8946 (N_8946,N_4186,N_4978);
nor U8947 (N_8947,N_5973,N_5829);
and U8948 (N_8948,N_3029,N_3901);
and U8949 (N_8949,N_3934,N_4833);
or U8950 (N_8950,N_5260,N_5986);
or U8951 (N_8951,N_3822,N_3838);
or U8952 (N_8952,N_5430,N_4933);
nand U8953 (N_8953,N_4233,N_5825);
and U8954 (N_8954,N_4999,N_4273);
and U8955 (N_8955,N_4387,N_5441);
and U8956 (N_8956,N_3787,N_3973);
nand U8957 (N_8957,N_3272,N_4149);
xor U8958 (N_8958,N_5154,N_5143);
nand U8959 (N_8959,N_5794,N_3847);
or U8960 (N_8960,N_5392,N_3557);
or U8961 (N_8961,N_3289,N_5661);
or U8962 (N_8962,N_4781,N_4003);
nand U8963 (N_8963,N_4790,N_5817);
and U8964 (N_8964,N_5131,N_3685);
or U8965 (N_8965,N_5842,N_4369);
xnor U8966 (N_8966,N_4174,N_4881);
or U8967 (N_8967,N_3212,N_5817);
nor U8968 (N_8968,N_5413,N_4782);
and U8969 (N_8969,N_3140,N_3792);
xnor U8970 (N_8970,N_3778,N_4577);
nand U8971 (N_8971,N_3635,N_5885);
xnor U8972 (N_8972,N_5764,N_4792);
or U8973 (N_8973,N_3811,N_5474);
or U8974 (N_8974,N_4937,N_5643);
nor U8975 (N_8975,N_5192,N_5259);
and U8976 (N_8976,N_5555,N_3776);
xnor U8977 (N_8977,N_4438,N_3435);
nor U8978 (N_8978,N_5350,N_3456);
xor U8979 (N_8979,N_4916,N_3815);
or U8980 (N_8980,N_4374,N_4348);
nand U8981 (N_8981,N_4169,N_4677);
xnor U8982 (N_8982,N_5477,N_5561);
nor U8983 (N_8983,N_5830,N_3665);
nand U8984 (N_8984,N_3831,N_4578);
and U8985 (N_8985,N_3391,N_3067);
nor U8986 (N_8986,N_5947,N_5928);
nor U8987 (N_8987,N_3050,N_3076);
or U8988 (N_8988,N_3414,N_5888);
xor U8989 (N_8989,N_4784,N_4335);
and U8990 (N_8990,N_4766,N_4555);
xor U8991 (N_8991,N_5468,N_5175);
and U8992 (N_8992,N_3125,N_3290);
xnor U8993 (N_8993,N_5499,N_5064);
xor U8994 (N_8994,N_4264,N_3556);
and U8995 (N_8995,N_4074,N_4179);
and U8996 (N_8996,N_5259,N_3179);
xnor U8997 (N_8997,N_3884,N_4326);
nand U8998 (N_8998,N_4450,N_3725);
or U8999 (N_8999,N_5706,N_3900);
xnor U9000 (N_9000,N_7042,N_8427);
xnor U9001 (N_9001,N_7810,N_8050);
xnor U9002 (N_9002,N_7441,N_6503);
nor U9003 (N_9003,N_7669,N_6667);
and U9004 (N_9004,N_6666,N_8950);
nand U9005 (N_9005,N_8967,N_7646);
and U9006 (N_9006,N_8863,N_6432);
nand U9007 (N_9007,N_6349,N_7733);
nor U9008 (N_9008,N_8291,N_8083);
xor U9009 (N_9009,N_6431,N_8959);
or U9010 (N_9010,N_7590,N_6661);
xor U9011 (N_9011,N_6880,N_7652);
xor U9012 (N_9012,N_7852,N_6485);
or U9013 (N_9013,N_8743,N_8750);
nor U9014 (N_9014,N_7535,N_7162);
nand U9015 (N_9015,N_6972,N_7099);
nand U9016 (N_9016,N_8136,N_6738);
or U9017 (N_9017,N_7465,N_6149);
xor U9018 (N_9018,N_7292,N_6071);
or U9019 (N_9019,N_7489,N_6148);
xnor U9020 (N_9020,N_7354,N_8847);
nand U9021 (N_9021,N_7897,N_8511);
or U9022 (N_9022,N_6652,N_8957);
nor U9023 (N_9023,N_7755,N_6933);
xor U9024 (N_9024,N_8092,N_8554);
xor U9025 (N_9025,N_8032,N_6935);
nand U9026 (N_9026,N_7629,N_6466);
xnor U9027 (N_9027,N_8824,N_6787);
nand U9028 (N_9028,N_8503,N_6082);
nor U9029 (N_9029,N_6608,N_7152);
or U9030 (N_9030,N_6792,N_8691);
or U9031 (N_9031,N_7018,N_8297);
nand U9032 (N_9032,N_8405,N_8848);
nor U9033 (N_9033,N_8197,N_8025);
xor U9034 (N_9034,N_7604,N_8949);
nand U9035 (N_9035,N_7155,N_7447);
nand U9036 (N_9036,N_7185,N_7355);
and U9037 (N_9037,N_8986,N_6087);
or U9038 (N_9038,N_7278,N_6470);
nor U9039 (N_9039,N_8714,N_8692);
or U9040 (N_9040,N_7095,N_8971);
nor U9041 (N_9041,N_6109,N_6521);
nor U9042 (N_9042,N_6379,N_8550);
nor U9043 (N_9043,N_7218,N_6258);
xnor U9044 (N_9044,N_8732,N_7221);
nand U9045 (N_9045,N_6386,N_7421);
or U9046 (N_9046,N_8107,N_8482);
xnor U9047 (N_9047,N_8505,N_7645);
or U9048 (N_9048,N_8239,N_6014);
or U9049 (N_9049,N_6140,N_8839);
and U9050 (N_9050,N_7051,N_6657);
nand U9051 (N_9051,N_7873,N_8854);
nor U9052 (N_9052,N_7937,N_6088);
and U9053 (N_9053,N_8140,N_8281);
or U9054 (N_9054,N_6736,N_7160);
nor U9055 (N_9055,N_7675,N_7188);
xor U9056 (N_9056,N_8320,N_7667);
nand U9057 (N_9057,N_7213,N_7343);
nand U9058 (N_9058,N_7148,N_8819);
or U9059 (N_9059,N_6823,N_6511);
nand U9060 (N_9060,N_8984,N_7439);
xnor U9061 (N_9061,N_7934,N_8703);
nor U9062 (N_9062,N_7577,N_8346);
or U9063 (N_9063,N_7472,N_8577);
xnor U9064 (N_9064,N_8471,N_7158);
nor U9065 (N_9065,N_7466,N_6984);
and U9066 (N_9066,N_8173,N_8319);
or U9067 (N_9067,N_8308,N_7593);
nor U9068 (N_9068,N_6436,N_7938);
or U9069 (N_9069,N_6942,N_7026);
nor U9070 (N_9070,N_8061,N_8566);
nand U9071 (N_9071,N_7723,N_6969);
nor U9072 (N_9072,N_6085,N_8288);
and U9073 (N_9073,N_6439,N_6094);
xnor U9074 (N_9074,N_6453,N_7971);
and U9075 (N_9075,N_6978,N_8335);
nor U9076 (N_9076,N_8290,N_8868);
nor U9077 (N_9077,N_6651,N_6514);
nand U9078 (N_9078,N_6421,N_7484);
nor U9079 (N_9079,N_8418,N_8029);
nor U9080 (N_9080,N_7431,N_8610);
xor U9081 (N_9081,N_7620,N_7970);
and U9082 (N_9082,N_8027,N_8857);
nand U9083 (N_9083,N_8240,N_8227);
nor U9084 (N_9084,N_8120,N_8101);
or U9085 (N_9085,N_6126,N_8499);
nor U9086 (N_9086,N_7144,N_8474);
nand U9087 (N_9087,N_6245,N_7333);
nor U9088 (N_9088,N_7528,N_7920);
xnor U9089 (N_9089,N_8416,N_7956);
nor U9090 (N_9090,N_7556,N_8300);
or U9091 (N_9091,N_7692,N_7109);
or U9092 (N_9092,N_8135,N_8406);
nor U9093 (N_9093,N_8070,N_6851);
nand U9094 (N_9094,N_8338,N_8768);
or U9095 (N_9095,N_8574,N_7836);
nand U9096 (N_9096,N_8008,N_7068);
or U9097 (N_9097,N_7178,N_7508);
and U9098 (N_9098,N_8560,N_8054);
nor U9099 (N_9099,N_7706,N_8496);
nand U9100 (N_9100,N_6417,N_6357);
and U9101 (N_9101,N_6817,N_7861);
or U9102 (N_9102,N_8347,N_7444);
xnor U9103 (N_9103,N_7210,N_6291);
and U9104 (N_9104,N_8634,N_8589);
nor U9105 (N_9105,N_6315,N_7949);
or U9106 (N_9106,N_7828,N_7731);
and U9107 (N_9107,N_7300,N_6873);
and U9108 (N_9108,N_8461,N_8313);
or U9109 (N_9109,N_8475,N_6610);
and U9110 (N_9110,N_8463,N_8830);
nand U9111 (N_9111,N_6264,N_7673);
and U9112 (N_9112,N_7850,N_7941);
and U9113 (N_9113,N_6958,N_7027);
nand U9114 (N_9114,N_8422,N_7690);
nand U9115 (N_9115,N_7778,N_6306);
and U9116 (N_9116,N_7437,N_7151);
xor U9117 (N_9117,N_6323,N_6102);
and U9118 (N_9118,N_7559,N_7182);
xor U9119 (N_9119,N_6639,N_7392);
nor U9120 (N_9120,N_7291,N_8219);
or U9121 (N_9121,N_6352,N_6504);
or U9122 (N_9122,N_6536,N_8758);
and U9123 (N_9123,N_6189,N_6027);
nor U9124 (N_9124,N_6856,N_7075);
xnor U9125 (N_9125,N_7043,N_7341);
or U9126 (N_9126,N_6412,N_6227);
xnor U9127 (N_9127,N_8097,N_6004);
and U9128 (N_9128,N_8642,N_6695);
nand U9129 (N_9129,N_7543,N_7927);
xor U9130 (N_9130,N_7180,N_6107);
and U9131 (N_9131,N_7262,N_6354);
or U9132 (N_9132,N_6546,N_6335);
or U9133 (N_9133,N_6911,N_6212);
nor U9134 (N_9134,N_8425,N_6670);
and U9135 (N_9135,N_8960,N_7693);
nor U9136 (N_9136,N_7174,N_6310);
xor U9137 (N_9137,N_7896,N_8127);
xor U9138 (N_9138,N_6635,N_6206);
nand U9139 (N_9139,N_7251,N_6089);
and U9140 (N_9140,N_7425,N_8798);
nand U9141 (N_9141,N_8433,N_7791);
nand U9142 (N_9142,N_8675,N_6685);
xnor U9143 (N_9143,N_6782,N_7924);
and U9144 (N_9144,N_7183,N_7638);
nor U9145 (N_9145,N_6325,N_8771);
xor U9146 (N_9146,N_8987,N_8039);
nor U9147 (N_9147,N_8075,N_6897);
and U9148 (N_9148,N_6960,N_8552);
or U9149 (N_9149,N_8722,N_7056);
nor U9150 (N_9150,N_8343,N_6717);
nand U9151 (N_9151,N_6114,N_6816);
xor U9152 (N_9152,N_7224,N_8063);
and U9153 (N_9153,N_8294,N_7812);
xor U9154 (N_9154,N_6876,N_7476);
xor U9155 (N_9155,N_8139,N_8792);
xor U9156 (N_9156,N_7594,N_7967);
xor U9157 (N_9157,N_6401,N_8782);
and U9158 (N_9158,N_8753,N_8316);
nor U9159 (N_9159,N_8924,N_7928);
nand U9160 (N_9160,N_7513,N_6831);
nand U9161 (N_9161,N_6518,N_6414);
nand U9162 (N_9162,N_6300,N_7222);
and U9163 (N_9163,N_8181,N_7790);
and U9164 (N_9164,N_6739,N_8390);
xnor U9165 (N_9165,N_7579,N_8966);
nand U9166 (N_9166,N_7602,N_6619);
xor U9167 (N_9167,N_7096,N_6205);
or U9168 (N_9168,N_6139,N_6026);
xor U9169 (N_9169,N_6266,N_8440);
nand U9170 (N_9170,N_8664,N_8146);
nor U9171 (N_9171,N_6865,N_6128);
xor U9172 (N_9172,N_8869,N_6679);
xnor U9173 (N_9173,N_6195,N_8177);
or U9174 (N_9174,N_6975,N_7592);
nor U9175 (N_9175,N_8669,N_7900);
and U9176 (N_9176,N_6533,N_6901);
xnor U9177 (N_9177,N_8270,N_7584);
xor U9178 (N_9178,N_7858,N_7655);
and U9179 (N_9179,N_7003,N_6309);
nor U9180 (N_9180,N_7798,N_6598);
and U9181 (N_9181,N_6735,N_6424);
and U9182 (N_9182,N_8866,N_8677);
nor U9183 (N_9183,N_8943,N_6721);
or U9184 (N_9184,N_6484,N_6479);
and U9185 (N_9185,N_7914,N_8815);
nand U9186 (N_9186,N_6725,N_6103);
and U9187 (N_9187,N_6429,N_8588);
nand U9188 (N_9188,N_7101,N_8807);
or U9189 (N_9189,N_7912,N_7512);
xor U9190 (N_9190,N_6776,N_6192);
or U9191 (N_9191,N_6364,N_8906);
and U9192 (N_9192,N_8538,N_8769);
nand U9193 (N_9193,N_8018,N_8658);
nand U9194 (N_9194,N_7232,N_8614);
nor U9195 (N_9195,N_7076,N_7752);
or U9196 (N_9196,N_6864,N_8805);
xnor U9197 (N_9197,N_7795,N_8071);
nand U9198 (N_9198,N_7377,N_6902);
and U9199 (N_9199,N_6037,N_8233);
or U9200 (N_9200,N_7371,N_7277);
and U9201 (N_9201,N_7611,N_7560);
and U9202 (N_9202,N_8752,N_7407);
or U9203 (N_9203,N_6395,N_8582);
nand U9204 (N_9204,N_8615,N_6755);
nor U9205 (N_9205,N_7997,N_6908);
and U9206 (N_9206,N_8251,N_8021);
nand U9207 (N_9207,N_6003,N_7127);
xnor U9208 (N_9208,N_8689,N_6146);
nor U9209 (N_9209,N_6572,N_6832);
and U9210 (N_9210,N_7568,N_8145);
nor U9211 (N_9211,N_7084,N_7697);
and U9212 (N_9212,N_8829,N_7236);
nor U9213 (N_9213,N_6222,N_8043);
or U9214 (N_9214,N_7793,N_6450);
and U9215 (N_9215,N_7954,N_8843);
xnor U9216 (N_9216,N_6279,N_8555);
or U9217 (N_9217,N_8502,N_8653);
xnor U9218 (N_9218,N_6813,N_8913);
xnor U9219 (N_9219,N_6059,N_6575);
xor U9220 (N_9220,N_6790,N_8572);
and U9221 (N_9221,N_7695,N_7086);
or U9222 (N_9222,N_6100,N_7618);
xor U9223 (N_9223,N_7478,N_6030);
nor U9224 (N_9224,N_7302,N_6815);
nor U9225 (N_9225,N_8019,N_6369);
nor U9226 (N_9226,N_7394,N_7662);
and U9227 (N_9227,N_7321,N_7996);
xor U9228 (N_9228,N_6034,N_8549);
or U9229 (N_9229,N_6645,N_6111);
or U9230 (N_9230,N_6091,N_7811);
and U9231 (N_9231,N_8404,N_6616);
nand U9232 (N_9232,N_8275,N_8383);
nor U9233 (N_9233,N_7973,N_8804);
xor U9234 (N_9234,N_7708,N_8944);
or U9235 (N_9235,N_8414,N_7890);
or U9236 (N_9236,N_6256,N_7619);
or U9237 (N_9237,N_7913,N_6550);
nor U9238 (N_9238,N_6664,N_8309);
nand U9239 (N_9239,N_6384,N_7322);
or U9240 (N_9240,N_8336,N_7936);
or U9241 (N_9241,N_6872,N_6544);
xor U9242 (N_9242,N_8413,N_6804);
and U9243 (N_9243,N_8800,N_6957);
nand U9244 (N_9244,N_6791,N_6543);
or U9245 (N_9245,N_7907,N_7044);
nand U9246 (N_9246,N_6631,N_7814);
or U9247 (N_9247,N_6185,N_6548);
nor U9248 (N_9248,N_8277,N_8933);
xnor U9249 (N_9249,N_7610,N_8153);
or U9250 (N_9250,N_6442,N_7600);
or U9251 (N_9251,N_8640,N_7758);
and U9252 (N_9252,N_7588,N_7265);
xnor U9253 (N_9253,N_6438,N_8081);
xor U9254 (N_9254,N_7782,N_8174);
and U9255 (N_9255,N_7124,N_8236);
nand U9256 (N_9256,N_6233,N_7868);
nand U9257 (N_9257,N_8789,N_7682);
or U9258 (N_9258,N_7903,N_6637);
nor U9259 (N_9259,N_6927,N_8108);
or U9260 (N_9260,N_7768,N_8485);
and U9261 (N_9261,N_7862,N_6702);
xor U9262 (N_9262,N_7062,N_8838);
nand U9263 (N_9263,N_6563,N_6886);
or U9264 (N_9264,N_8084,N_6951);
nor U9265 (N_9265,N_7589,N_6096);
nand U9266 (N_9266,N_8392,N_6783);
xor U9267 (N_9267,N_8702,N_8776);
xnor U9268 (N_9268,N_7209,N_7743);
and U9269 (N_9269,N_6799,N_6579);
nand U9270 (N_9270,N_7889,N_6105);
or U9271 (N_9271,N_7440,N_8668);
xor U9272 (N_9272,N_7073,N_7507);
or U9273 (N_9273,N_7331,N_8875);
nand U9274 (N_9274,N_8410,N_6780);
and U9275 (N_9275,N_7179,N_8852);
or U9276 (N_9276,N_7296,N_6440);
and U9277 (N_9277,N_7865,N_6242);
or U9278 (N_9278,N_8059,N_6928);
xnor U9279 (N_9279,N_8911,N_6081);
and U9280 (N_9280,N_8927,N_7734);
or U9281 (N_9281,N_8565,N_6964);
and U9282 (N_9282,N_7035,N_6696);
xnor U9283 (N_9283,N_6072,N_6896);
and U9284 (N_9284,N_7855,N_8030);
and U9285 (N_9285,N_7069,N_7842);
nor U9286 (N_9286,N_7367,N_6508);
and U9287 (N_9287,N_6983,N_6122);
nor U9288 (N_9288,N_8573,N_8352);
nor U9289 (N_9289,N_8730,N_7665);
nor U9290 (N_9290,N_7819,N_8199);
nand U9291 (N_9291,N_7966,N_8431);
xnor U9292 (N_9292,N_7411,N_7376);
nor U9293 (N_9293,N_8564,N_8686);
and U9294 (N_9294,N_8129,N_6058);
xor U9295 (N_9295,N_6493,N_6768);
nor U9296 (N_9296,N_7882,N_8882);
nand U9297 (N_9297,N_7736,N_6643);
nor U9298 (N_9298,N_8327,N_8515);
or U9299 (N_9299,N_8939,N_8417);
xnor U9300 (N_9300,N_7995,N_8131);
or U9301 (N_9301,N_7931,N_7844);
nand U9302 (N_9302,N_6729,N_7306);
nand U9303 (N_9303,N_7930,N_8473);
or U9304 (N_9304,N_7244,N_7651);
and U9305 (N_9305,N_7766,N_7194);
or U9306 (N_9306,N_7316,N_7516);
nand U9307 (N_9307,N_8783,N_7517);
nand U9308 (N_9308,N_7678,N_8072);
or U9309 (N_9309,N_7351,N_8304);
xnor U9310 (N_9310,N_6870,N_6853);
nor U9311 (N_9311,N_8516,N_8157);
or U9312 (N_9312,N_8749,N_6904);
xor U9313 (N_9313,N_8657,N_7837);
or U9314 (N_9314,N_8881,N_8729);
nor U9315 (N_9315,N_7356,N_7338);
or U9316 (N_9316,N_6333,N_6991);
or U9317 (N_9317,N_7202,N_6557);
and U9318 (N_9318,N_6118,N_8909);
nand U9319 (N_9319,N_6237,N_7252);
and U9320 (N_9320,N_7420,N_8213);
or U9321 (N_9321,N_8429,N_6952);
xor U9322 (N_9322,N_8231,N_8331);
and U9323 (N_9323,N_6298,N_7279);
and U9324 (N_9324,N_6177,N_8919);
and U9325 (N_9325,N_8188,N_6859);
or U9326 (N_9326,N_6270,N_6419);
xor U9327 (N_9327,N_7456,N_7985);
nand U9328 (N_9328,N_8643,N_8481);
xor U9329 (N_9329,N_6934,N_7036);
nand U9330 (N_9330,N_7840,N_8898);
nor U9331 (N_9331,N_8522,N_7114);
nor U9332 (N_9332,N_6658,N_8712);
xnor U9333 (N_9333,N_7267,N_8823);
nand U9334 (N_9334,N_8611,N_6130);
nand U9335 (N_9335,N_6181,N_8479);
and U9336 (N_9336,N_6962,N_7198);
and U9337 (N_9337,N_7091,N_7130);
xnor U9338 (N_9338,N_8625,N_8649);
or U9339 (N_9339,N_6948,N_8850);
and U9340 (N_9340,N_6216,N_6158);
nor U9341 (N_9341,N_8841,N_8631);
and U9342 (N_9342,N_6630,N_6372);
or U9343 (N_9343,N_8785,N_8598);
nand U9344 (N_9344,N_7094,N_8969);
nand U9345 (N_9345,N_8684,N_6527);
or U9346 (N_9346,N_8916,N_6673);
nand U9347 (N_9347,N_8619,N_8215);
nand U9348 (N_9348,N_6537,N_7845);
nor U9349 (N_9349,N_8604,N_6744);
nor U9350 (N_9350,N_7348,N_7546);
nand U9351 (N_9351,N_8500,N_8818);
nor U9352 (N_9352,N_7683,N_7770);
nor U9353 (N_9353,N_8076,N_6690);
and U9354 (N_9354,N_8263,N_6207);
and U9355 (N_9355,N_7090,N_7515);
nand U9356 (N_9356,N_6239,N_7403);
or U9357 (N_9357,N_7497,N_6775);
or U9358 (N_9358,N_6640,N_7181);
or U9359 (N_9359,N_8756,N_8133);
and U9360 (N_9360,N_6973,N_6737);
nand U9361 (N_9361,N_6510,N_7237);
xor U9362 (N_9362,N_7243,N_7963);
nand U9363 (N_9363,N_8370,N_6211);
nor U9364 (N_9364,N_7848,N_7370);
xor U9365 (N_9365,N_6506,N_6191);
nand U9366 (N_9366,N_7635,N_8261);
xnor U9367 (N_9367,N_8864,N_6993);
nand U9368 (N_9368,N_8015,N_6324);
xnor U9369 (N_9369,N_7072,N_8055);
and U9370 (N_9370,N_7360,N_8583);
or U9371 (N_9371,N_7040,N_7113);
and U9372 (N_9372,N_8531,N_6407);
or U9373 (N_9373,N_6376,N_7541);
nand U9374 (N_9374,N_6476,N_8045);
and U9375 (N_9375,N_7303,N_6663);
xnor U9376 (N_9376,N_8917,N_6293);
and U9377 (N_9377,N_8895,N_8813);
or U9378 (N_9378,N_8034,N_6743);
and U9379 (N_9379,N_6774,N_8945);
or U9380 (N_9380,N_7245,N_7741);
and U9381 (N_9381,N_8685,N_6634);
or U9382 (N_9382,N_6649,N_6019);
or U9383 (N_9383,N_6405,N_8925);
nor U9384 (N_9384,N_6621,N_6194);
or U9385 (N_9385,N_8205,N_8036);
nand U9386 (N_9386,N_8662,N_7459);
or U9387 (N_9387,N_6924,N_8058);
nand U9388 (N_9388,N_6779,N_6998);
xnor U9389 (N_9389,N_8698,N_8301);
nand U9390 (N_9390,N_7728,N_6229);
xnor U9391 (N_9391,N_6068,N_6187);
and U9392 (N_9392,N_8374,N_6892);
nand U9393 (N_9393,N_8575,N_6017);
and U9394 (N_9394,N_8530,N_7382);
and U9395 (N_9395,N_7942,N_7872);
or U9396 (N_9396,N_6127,N_6327);
nor U9397 (N_9397,N_7491,N_7779);
or U9398 (N_9398,N_8412,N_6628);
or U9399 (N_9399,N_8033,N_6841);
or U9400 (N_9400,N_8764,N_7052);
nand U9401 (N_9401,N_7305,N_6767);
xnor U9402 (N_9402,N_8477,N_6562);
xnor U9403 (N_9403,N_7234,N_7603);
nand U9404 (N_9404,N_7999,N_7984);
nor U9405 (N_9405,N_8062,N_6837);
or U9406 (N_9406,N_7353,N_7193);
and U9407 (N_9407,N_8194,N_6223);
nand U9408 (N_9408,N_6588,N_7197);
or U9409 (N_9409,N_7994,N_8525);
xnor U9410 (N_9410,N_7529,N_8437);
xnor U9411 (N_9411,N_7294,N_7521);
or U9412 (N_9412,N_8734,N_7415);
and U9413 (N_9413,N_7640,N_7263);
nor U9414 (N_9414,N_8394,N_7961);
or U9415 (N_9415,N_8355,N_7867);
xor U9416 (N_9416,N_8638,N_7328);
nor U9417 (N_9417,N_8393,N_8627);
nand U9418 (N_9418,N_7481,N_6342);
and U9419 (N_9419,N_7548,N_6715);
nor U9420 (N_9420,N_8468,N_6273);
or U9421 (N_9421,N_8371,N_8968);
nand U9422 (N_9422,N_6574,N_8727);
and U9423 (N_9423,N_7346,N_7668);
xor U9424 (N_9424,N_6701,N_7166);
or U9425 (N_9425,N_6750,N_7434);
and U9426 (N_9426,N_7694,N_7164);
xor U9427 (N_9427,N_6974,N_6764);
and U9428 (N_9428,N_7864,N_8624);
xor U9429 (N_9429,N_8144,N_6977);
nand U9430 (N_9430,N_6923,N_6362);
or U9431 (N_9431,N_7974,N_7396);
and U9432 (N_9432,N_6806,N_6997);
or U9433 (N_9433,N_6938,N_6117);
nand U9434 (N_9434,N_8469,N_6238);
and U9435 (N_9435,N_6408,N_7034);
xor U9436 (N_9436,N_6077,N_6818);
xor U9437 (N_9437,N_7945,N_7225);
xnor U9438 (N_9438,N_8321,N_7064);
nand U9439 (N_9439,N_8149,N_6252);
and U9440 (N_9440,N_7223,N_8628);
xor U9441 (N_9441,N_7313,N_8935);
nor U9442 (N_9442,N_8249,N_8951);
xor U9443 (N_9443,N_7835,N_8187);
and U9444 (N_9444,N_6219,N_7575);
and U9445 (N_9445,N_8781,N_8773);
nand U9446 (N_9446,N_7979,N_8138);
nand U9447 (N_9447,N_7813,N_8360);
and U9448 (N_9448,N_6013,N_8762);
or U9449 (N_9449,N_6677,N_7080);
and U9450 (N_9450,N_8623,N_7659);
xnor U9451 (N_9451,N_7550,N_6836);
nor U9452 (N_9452,N_7599,N_7270);
nor U9453 (N_9453,N_6009,N_8837);
nor U9454 (N_9454,N_8232,N_7312);
or U9455 (N_9455,N_6980,N_6542);
or U9456 (N_9456,N_6012,N_7388);
or U9457 (N_9457,N_7247,N_8533);
and U9458 (N_9458,N_8535,N_8467);
nor U9459 (N_9459,N_6553,N_7774);
and U9460 (N_9460,N_7473,N_8570);
nand U9461 (N_9461,N_8150,N_7772);
nand U9462 (N_9462,N_6937,N_6008);
and U9463 (N_9463,N_7686,N_7977);
and U9464 (N_9464,N_7275,N_8717);
nor U9465 (N_9465,N_7991,N_7192);
nand U9466 (N_9466,N_6204,N_7029);
and U9467 (N_9467,N_7171,N_7688);
or U9468 (N_9468,N_8885,N_7239);
xor U9469 (N_9469,N_6530,N_7750);
or U9470 (N_9470,N_7827,N_6294);
nand U9471 (N_9471,N_8497,N_7429);
and U9472 (N_9472,N_8681,N_7884);
and U9473 (N_9473,N_7137,N_7014);
xor U9474 (N_9474,N_7187,N_7413);
xor U9475 (N_9475,N_6602,N_7627);
and U9476 (N_9476,N_6752,N_8774);
and U9477 (N_9477,N_7039,N_7136);
nor U9478 (N_9478,N_7710,N_6501);
nor U9479 (N_9479,N_6040,N_8388);
nand U9480 (N_9480,N_6312,N_8521);
xor U9481 (N_9481,N_8652,N_7820);
nand U9482 (N_9482,N_6692,N_8910);
or U9483 (N_9483,N_7764,N_8472);
and U9484 (N_9484,N_7060,N_8715);
xor U9485 (N_9485,N_8341,N_7940);
nor U9486 (N_9486,N_7121,N_8286);
and U9487 (N_9487,N_6878,N_6581);
nand U9488 (N_9488,N_6397,N_8078);
nand U9489 (N_9489,N_6618,N_7045);
nand U9490 (N_9490,N_8465,N_7511);
or U9491 (N_9491,N_6474,N_6808);
xnor U9492 (N_9492,N_7280,N_8845);
nor U9493 (N_9493,N_8218,N_7740);
or U9494 (N_9494,N_8733,N_6910);
or U9495 (N_9495,N_8886,N_6035);
or U9496 (N_9496,N_8400,N_8825);
xnor U9497 (N_9497,N_6093,N_7266);
or U9498 (N_9498,N_8920,N_6883);
and U9499 (N_9499,N_6796,N_8606);
or U9500 (N_9500,N_6269,N_8526);
or U9501 (N_9501,N_8376,N_6344);
nor U9502 (N_9502,N_7735,N_8013);
xor U9503 (N_9503,N_6731,N_8047);
or U9504 (N_9504,N_7796,N_6490);
xor U9505 (N_9505,N_6918,N_8183);
nor U9506 (N_9506,N_8965,N_8123);
or U9507 (N_9507,N_7832,N_6489);
xor U9508 (N_9508,N_8849,N_8247);
xnor U9509 (N_9509,N_8802,N_8322);
or U9510 (N_9510,N_6593,N_8736);
or U9511 (N_9511,N_7424,N_7079);
or U9512 (N_9512,N_8840,N_7038);
nor U9513 (N_9513,N_7493,N_8994);
and U9514 (N_9514,N_8889,N_6567);
nand U9515 (N_9515,N_6039,N_7165);
and U9516 (N_9516,N_6578,N_8086);
nand U9517 (N_9517,N_6404,N_8591);
nor U9518 (N_9518,N_8922,N_7061);
xor U9519 (N_9519,N_6164,N_8141);
or U9520 (N_9520,N_7107,N_7962);
nand U9521 (N_9521,N_6084,N_6175);
and U9522 (N_9522,N_6794,N_6316);
nand U9523 (N_9523,N_8048,N_6263);
nand U9524 (N_9524,N_7551,N_8586);
nand U9525 (N_9525,N_6171,N_7345);
xnor U9526 (N_9526,N_7500,N_6531);
and U9527 (N_9527,N_7946,N_8861);
nor U9528 (N_9528,N_8244,N_6587);
or U9529 (N_9529,N_6547,N_6966);
xnor U9530 (N_9530,N_6512,N_8407);
and U9531 (N_9531,N_7057,N_6698);
xnor U9532 (N_9532,N_8432,N_6576);
nor U9533 (N_9533,N_6820,N_7358);
and U9534 (N_9534,N_8532,N_7537);
xor U9535 (N_9535,N_8763,N_7077);
xnor U9536 (N_9536,N_7721,N_8038);
or U9537 (N_9537,N_8613,N_6410);
nand U9538 (N_9538,N_8787,N_6329);
nor U9539 (N_9539,N_6193,N_8833);
nand U9540 (N_9540,N_6970,N_7326);
nand U9541 (N_9541,N_6538,N_8793);
and U9542 (N_9542,N_7738,N_7909);
or U9543 (N_9543,N_6929,N_8246);
xnor U9544 (N_9544,N_8650,N_8937);
nor U9545 (N_9545,N_7704,N_7825);
nor U9546 (N_9546,N_8741,N_6622);
or U9547 (N_9547,N_7253,N_7859);
xnor U9548 (N_9548,N_6104,N_7587);
or U9549 (N_9549,N_6110,N_7526);
xnor U9550 (N_9550,N_6788,N_7111);
or U9551 (N_9551,N_7958,N_6064);
nand U9552 (N_9552,N_7159,N_7965);
nand U9553 (N_9553,N_7536,N_6341);
nor U9554 (N_9554,N_6625,N_7561);
or U9555 (N_9555,N_6320,N_7432);
xor U9556 (N_9556,N_6825,N_7916);
or U9557 (N_9557,N_8444,N_6488);
and U9558 (N_9558,N_7074,N_6370);
nand U9559 (N_9559,N_6683,N_8009);
or U9560 (N_9560,N_7830,N_6250);
nand U9561 (N_9561,N_6704,N_8867);
xnor U9562 (N_9562,N_8723,N_6125);
or U9563 (N_9563,N_6433,N_8186);
or U9564 (N_9564,N_8912,N_8524);
or U9565 (N_9565,N_7104,N_6778);
xnor U9566 (N_9566,N_8095,N_6525);
and U9567 (N_9567,N_8216,N_8373);
nor U9568 (N_9568,N_7910,N_6711);
xor U9569 (N_9569,N_7625,N_7059);
and U9570 (N_9570,N_7332,N_8822);
nor U9571 (N_9571,N_8639,N_6772);
nor U9572 (N_9572,N_6385,N_8104);
and U9573 (N_9573,N_8720,N_7480);
or U9574 (N_9574,N_6360,N_6044);
nand U9575 (N_9575,N_6340,N_8602);
and U9576 (N_9576,N_8545,N_7482);
nor U9577 (N_9577,N_6838,N_7430);
nand U9578 (N_9578,N_6707,N_8165);
nor U9579 (N_9579,N_6914,N_6083);
nor U9580 (N_9580,N_6287,N_8980);
nor U9581 (N_9581,N_7661,N_8234);
and U9582 (N_9582,N_6671,N_7401);
nand U9583 (N_9583,N_8222,N_6373);
nand U9584 (N_9584,N_6319,N_6786);
nor U9585 (N_9585,N_7339,N_6422);
or U9586 (N_9586,N_8963,N_8459);
nor U9587 (N_9587,N_6693,N_8991);
or U9588 (N_9588,N_8509,N_7379);
xor U9589 (N_9589,N_8484,N_8243);
nand U9590 (N_9590,N_6604,N_8399);
xor U9591 (N_9591,N_6852,N_7047);
xnor U9592 (N_9592,N_7423,N_8452);
and U9593 (N_9593,N_6654,N_6168);
nand U9594 (N_9594,N_8827,N_8274);
xor U9595 (N_9595,N_7381,N_7499);
nand U9596 (N_9596,N_8656,N_7639);
or U9597 (N_9597,N_6495,N_7450);
and U9598 (N_9598,N_6116,N_7446);
xor U9599 (N_9599,N_8035,N_6653);
nand U9600 (N_9600,N_6172,N_8421);
and U9601 (N_9601,N_7334,N_8042);
nor U9602 (N_9602,N_7642,N_6353);
xnor U9603 (N_9603,N_7570,N_6151);
nor U9604 (N_9604,N_8816,N_8790);
nand U9605 (N_9605,N_7011,N_8988);
or U9606 (N_9606,N_6748,N_6443);
nand U9607 (N_9607,N_8871,N_6720);
or U9608 (N_9608,N_6515,N_8812);
or U9609 (N_9609,N_8637,N_6160);
nand U9610 (N_9610,N_7871,N_8934);
xor U9611 (N_9611,N_7238,N_6023);
xnor U9612 (N_9612,N_7032,N_6762);
or U9613 (N_9613,N_8000,N_6028);
nor U9614 (N_9614,N_7250,N_6979);
nor U9615 (N_9615,N_7255,N_6002);
or U9616 (N_9616,N_8620,N_6284);
and U9617 (N_9617,N_6459,N_7801);
or U9618 (N_9618,N_8630,N_7458);
nand U9619 (N_9619,N_7065,N_8193);
xnor U9620 (N_9620,N_7899,N_7953);
nor U9621 (N_9621,N_7081,N_7295);
xor U9622 (N_9622,N_6680,N_7847);
or U9623 (N_9623,N_8109,N_7426);
nand U9624 (N_9624,N_8896,N_6260);
or U9625 (N_9625,N_8160,N_6569);
nor U9626 (N_9626,N_6272,N_6015);
nand U9627 (N_9627,N_6871,N_8085);
and U9628 (N_9628,N_6090,N_7744);
and U9629 (N_9629,N_8434,N_8491);
nand U9630 (N_9630,N_6423,N_6461);
xnor U9631 (N_9631,N_8184,N_8080);
xor U9632 (N_9632,N_7319,N_7126);
or U9633 (N_9633,N_6482,N_6051);
nand U9634 (N_9634,N_6766,N_6697);
xor U9635 (N_9635,N_8894,N_6699);
nand U9636 (N_9636,N_6464,N_8143);
or U9637 (N_9637,N_8455,N_6170);
and U9638 (N_9638,N_8476,N_8259);
nor U9639 (N_9639,N_6347,N_7007);
or U9640 (N_9640,N_7630,N_7598);
nor U9641 (N_9641,N_6304,N_6332);
nand U9642 (N_9642,N_6981,N_7140);
or U9643 (N_9643,N_6848,N_8674);
nor U9644 (N_9644,N_8384,N_7374);
nor U9645 (N_9645,N_6789,N_7176);
or U9646 (N_9646,N_8273,N_6903);
nor U9647 (N_9647,N_7874,N_8266);
nand U9648 (N_9648,N_7384,N_7988);
nor U9649 (N_9649,N_7474,N_7142);
nor U9650 (N_9650,N_8151,N_6967);
nor U9651 (N_9651,N_7133,N_7654);
nor U9652 (N_9652,N_7976,N_6611);
and U9653 (N_9653,N_6947,N_8651);
or U9654 (N_9654,N_8398,N_6295);
or U9655 (N_9655,N_6339,N_7103);
nor U9656 (N_9656,N_6157,N_7408);
nand U9657 (N_9657,N_8292,N_6142);
xor U9658 (N_9658,N_7623,N_7992);
xor U9659 (N_9659,N_6594,N_6235);
and U9660 (N_9660,N_7259,N_8494);
or U9661 (N_9661,N_6571,N_6054);
nand U9662 (N_9662,N_8954,N_8207);
nand U9663 (N_9663,N_6770,N_6060);
nor U9664 (N_9664,N_6894,N_6392);
nand U9665 (N_9665,N_6159,N_8523);
nor U9666 (N_9666,N_8103,N_8661);
nand U9667 (N_9667,N_7856,N_7893);
and U9668 (N_9668,N_7048,N_6828);
nand U9669 (N_9669,N_7621,N_6468);
nand U9670 (N_9670,N_7248,N_7317);
nor U9671 (N_9671,N_6123,N_7925);
nand U9672 (N_9672,N_7921,N_8710);
and U9673 (N_9673,N_8453,N_6773);
xor U9674 (N_9674,N_8609,N_7699);
nand U9675 (N_9675,N_8245,N_8325);
xnor U9676 (N_9676,N_7097,N_6497);
nor U9677 (N_9677,N_8357,N_7622);
and U9678 (N_9678,N_6491,N_8719);
nand U9679 (N_9679,N_7019,N_7718);
xnor U9680 (N_9680,N_7205,N_7514);
nor U9681 (N_9681,N_6945,N_7713);
nand U9682 (N_9682,N_7116,N_7299);
and U9683 (N_9683,N_7046,N_8351);
nand U9684 (N_9684,N_7657,N_6383);
nor U9685 (N_9685,N_6596,N_7211);
nor U9686 (N_9686,N_7748,N_8046);
nand U9687 (N_9687,N_8017,N_7745);
and U9688 (N_9688,N_7617,N_6730);
nor U9689 (N_9689,N_8704,N_8527);
nor U9690 (N_9690,N_8470,N_8809);
and U9691 (N_9691,N_6198,N_7083);
nand U9692 (N_9692,N_6907,N_8587);
or U9693 (N_9693,N_7824,N_6334);
nand U9694 (N_9694,N_6555,N_7714);
and U9695 (N_9695,N_6277,N_7443);
nand U9696 (N_9696,N_6708,N_6124);
and U9697 (N_9697,N_6154,N_6632);
or U9698 (N_9698,N_8578,N_6247);
or U9699 (N_9699,N_7455,N_8411);
nand U9700 (N_9700,N_6156,N_8821);
nor U9701 (N_9701,N_6188,N_7853);
nor U9702 (N_9702,N_7063,N_7787);
xnor U9703 (N_9703,N_7643,N_7416);
xnor U9704 (N_9704,N_6812,N_7919);
nand U9705 (N_9705,N_8731,N_6275);
xor U9706 (N_9706,N_6337,N_8212);
nand U9707 (N_9707,N_6393,N_6522);
nand U9708 (N_9708,N_6868,N_7800);
or U9709 (N_9709,N_6798,N_8303);
and U9710 (N_9710,N_7908,N_7866);
or U9711 (N_9711,N_6426,N_7428);
or U9712 (N_9712,N_6655,N_7823);
nand U9713 (N_9713,N_7542,N_6819);
nand U9714 (N_9714,N_6590,N_8056);
or U9715 (N_9715,N_8788,N_6763);
or U9716 (N_9716,N_7632,N_8961);
nand U9717 (N_9717,N_8716,N_8449);
or U9718 (N_9718,N_8093,N_8345);
nand U9719 (N_9719,N_7696,N_8483);
nor U9720 (N_9720,N_7849,N_6437);
xnor U9721 (N_9721,N_7947,N_8022);
or U9722 (N_9722,N_6824,N_6609);
nor U9723 (N_9723,N_6940,N_7301);
nor U9724 (N_9724,N_8632,N_6351);
nor U9725 (N_9725,N_7150,N_7709);
and U9726 (N_9726,N_8167,N_7722);
nand U9727 (N_9727,N_8999,N_6668);
or U9728 (N_9728,N_8893,N_8220);
or U9729 (N_9729,N_6220,N_8419);
xnor U9730 (N_9730,N_6108,N_8176);
and U9731 (N_9731,N_6931,N_6046);
xnor U9732 (N_9732,N_7402,N_8377);
xnor U9733 (N_9733,N_8817,N_7939);
nor U9734 (N_9734,N_8952,N_7049);
nand U9735 (N_9735,N_8814,N_6186);
or U9736 (N_9736,N_6165,N_7555);
or U9737 (N_9737,N_8880,N_8460);
and U9738 (N_9738,N_7705,N_6190);
nand U9739 (N_9739,N_7843,N_6867);
nor U9740 (N_9740,N_8978,N_8673);
nand U9741 (N_9741,N_8512,N_8507);
nand U9742 (N_9742,N_7664,N_8581);
and U9743 (N_9743,N_8116,N_8264);
nor U9744 (N_9744,N_6452,N_6881);
nor U9745 (N_9745,N_7106,N_6056);
xor U9746 (N_9746,N_7269,N_8799);
or U9747 (N_9747,N_7539,N_6888);
nand U9748 (N_9748,N_7666,N_8958);
nor U9749 (N_9749,N_8326,N_7540);
and U9750 (N_9750,N_8592,N_8102);
and U9751 (N_9751,N_8744,N_6467);
or U9752 (N_9752,N_7031,N_8659);
xor U9753 (N_9753,N_6016,N_6182);
xor U9754 (N_9754,N_6753,N_7763);
nand U9755 (N_9755,N_8279,N_7214);
nor U9756 (N_9756,N_8010,N_7204);
and U9757 (N_9757,N_8024,N_7118);
nand U9758 (N_9758,N_8340,N_7254);
and U9759 (N_9759,N_7955,N_6318);
xor U9760 (N_9760,N_7463,N_7352);
xor U9761 (N_9761,N_8887,N_6595);
xor U9762 (N_9762,N_7993,N_6135);
or U9763 (N_9763,N_7329,N_8998);
nor U9764 (N_9764,N_7172,N_6221);
nand U9765 (N_9765,N_6827,N_7405);
nor U9766 (N_9766,N_7271,N_7229);
nand U9767 (N_9767,N_7576,N_6863);
xor U9768 (N_9768,N_6153,N_7404);
or U9769 (N_9769,N_7672,N_7131);
and U9770 (N_9770,N_8899,N_8040);
xnor U9771 (N_9771,N_6274,N_8990);
and U9772 (N_9772,N_8458,N_7684);
xor U9773 (N_9773,N_8112,N_7167);
nor U9774 (N_9774,N_8997,N_7510);
xor U9775 (N_9775,N_7717,N_7342);
nand U9776 (N_9776,N_8683,N_8299);
nor U9777 (N_9777,N_8617,N_7730);
nand U9778 (N_9778,N_6719,N_7324);
or U9779 (N_9779,N_8923,N_8621);
xnor U9780 (N_9780,N_7315,N_7451);
nor U9781 (N_9781,N_7711,N_8077);
nand U9782 (N_9782,N_7902,N_8278);
and U9783 (N_9783,N_8682,N_7146);
xor U9784 (N_9784,N_7981,N_7207);
nand U9785 (N_9785,N_7490,N_7002);
or U9786 (N_9786,N_8385,N_7505);
xnor U9787 (N_9787,N_8540,N_8645);
nand U9788 (N_9788,N_8446,N_8096);
nor U9789 (N_9789,N_6617,N_7479);
nor U9790 (N_9790,N_6874,N_7904);
nand U9791 (N_9791,N_7799,N_8890);
xnor U9792 (N_9792,N_8439,N_8065);
nor U9793 (N_9793,N_8551,N_7477);
nor U9794 (N_9794,N_7534,N_7707);
or U9795 (N_9795,N_6196,N_7102);
and U9796 (N_9796,N_6709,N_8295);
nor U9797 (N_9797,N_6201,N_8114);
nand U9798 (N_9798,N_6636,N_6714);
and U9799 (N_9799,N_6112,N_7530);
or U9800 (N_9800,N_6502,N_6650);
nor U9801 (N_9801,N_7760,N_6943);
nor U9802 (N_9802,N_7361,N_7948);
nand U9803 (N_9803,N_7742,N_8751);
xnor U9804 (N_9804,N_8772,N_7242);
or U9805 (N_9805,N_6416,N_7390);
and U9806 (N_9806,N_7287,N_7634);
xor U9807 (N_9807,N_7691,N_6292);
or U9808 (N_9808,N_8725,N_6313);
and U9809 (N_9809,N_8011,N_6218);
or U9810 (N_9810,N_8330,N_8835);
nor U9811 (N_9811,N_8663,N_8172);
or U9812 (N_9812,N_7869,N_6167);
or U9813 (N_9813,N_6913,N_6010);
xnor U9814 (N_9814,N_6570,N_6202);
xor U9815 (N_9815,N_8369,N_8348);
nor U9816 (N_9816,N_6687,N_7671);
nor U9817 (N_9817,N_7241,N_7147);
nand U9818 (N_9818,N_6742,N_7877);
and U9819 (N_9819,N_6282,N_7807);
or U9820 (N_9820,N_8152,N_7935);
xor U9821 (N_9821,N_6759,N_6358);
nor U9822 (N_9822,N_6932,N_6532);
or U9823 (N_9823,N_6672,N_8430);
xor U9824 (N_9824,N_6173,N_8903);
nand U9825 (N_9825,N_8700,N_6477);
and U9826 (N_9826,N_8955,N_8618);
xnor U9827 (N_9827,N_8190,N_6866);
nor U9828 (N_9828,N_7105,N_6529);
nand U9829 (N_9829,N_7574,N_6965);
or U9830 (N_9830,N_8831,N_8438);
nand U9831 (N_9831,N_7990,N_7389);
nand U9832 (N_9832,N_6771,N_7829);
xnor U9833 (N_9833,N_7933,N_8450);
nor U9834 (N_9834,N_6254,N_6001);
xnor U9835 (N_9835,N_8546,N_6845);
nor U9836 (N_9836,N_8626,N_8169);
xor U9837 (N_9837,N_6080,N_7739);
xnor U9838 (N_9838,N_8806,N_7566);
nand U9839 (N_9839,N_8576,N_7433);
nor U9840 (N_9840,N_7132,N_8794);
nand U9841 (N_9841,N_6380,N_6063);
or U9842 (N_9842,N_7041,N_6740);
xnor U9843 (N_9843,N_7344,N_6183);
nor U9844 (N_9844,N_6471,N_7289);
xnor U9845 (N_9845,N_6891,N_8445);
or U9846 (N_9846,N_7591,N_8122);
and U9847 (N_9847,N_8293,N_8254);
xor U9848 (N_9848,N_6356,N_6612);
and U9849 (N_9849,N_7318,N_8711);
xnor U9850 (N_9850,N_6539,N_7487);
nor U9851 (N_9851,N_6826,N_8358);
nor U9852 (N_9852,N_8088,N_6062);
nor U9853 (N_9853,N_7020,N_7464);
and U9854 (N_9854,N_6152,N_7751);
and U9855 (N_9855,N_7161,N_6255);
nand U9856 (N_9856,N_6633,N_6987);
and U9857 (N_9857,N_8601,N_6208);
or U9858 (N_9858,N_8436,N_6345);
nor U9859 (N_9859,N_6733,N_7327);
nand U9860 (N_9860,N_8189,N_7274);
or U9861 (N_9861,N_7553,N_6920);
or U9862 (N_9862,N_6906,N_7397);
or U9863 (N_9863,N_7506,N_6627);
and U9864 (N_9864,N_7347,N_8784);
nand U9865 (N_9865,N_8622,N_6231);
xor U9866 (N_9866,N_7380,N_7545);
nand U9867 (N_9867,N_8766,N_8306);
or U9868 (N_9868,N_7637,N_8599);
nand U9869 (N_9869,N_8907,N_7952);
or U9870 (N_9870,N_6936,N_7788);
or U9871 (N_9871,N_6811,N_8745);
nor U9872 (N_9872,N_6849,N_7395);
nand U9873 (N_9873,N_6830,N_8087);
and U9874 (N_9874,N_8694,N_6810);
and U9875 (N_9875,N_7297,N_7391);
xnor U9876 (N_9876,N_6716,N_6784);
and U9877 (N_9877,N_6496,N_8915);
nor U9878 (N_9878,N_8302,N_8031);
xor U9879 (N_9879,N_6996,N_6517);
and U9880 (N_9880,N_6359,N_8982);
xnor U9881 (N_9881,N_7438,N_7771);
and U9882 (N_9882,N_7915,N_6528);
and U9883 (N_9883,N_6603,N_8519);
or U9884 (N_9884,N_8296,N_8687);
nand U9885 (N_9885,N_7834,N_8801);
nand U9886 (N_9886,N_6577,N_8049);
and U9887 (N_9887,N_8230,N_6785);
or U9888 (N_9888,N_8111,N_6558);
and U9889 (N_9889,N_6399,N_6469);
and U9890 (N_9890,N_8761,N_6656);
xnor U9891 (N_9891,N_8182,N_8211);
nor U9892 (N_9892,N_8580,N_6475);
nor U9893 (N_9893,N_6814,N_8367);
nor U9894 (N_9894,N_8853,N_7201);
and U9895 (N_9895,N_7365,N_8217);
or U9896 (N_9896,N_6289,N_8976);
nor U9897 (N_9897,N_8158,N_7323);
nor U9898 (N_9898,N_8644,N_6197);
nand U9899 (N_9899,N_6133,N_8175);
and U9900 (N_9900,N_7372,N_8334);
xnor U9901 (N_9901,N_8778,N_7607);
or U9902 (N_9902,N_7596,N_8386);
nand U9903 (N_9903,N_7917,N_7776);
and U9904 (N_9904,N_7217,N_7724);
xor U9905 (N_9905,N_7154,N_7016);
nand U9906 (N_9906,N_8562,N_8020);
nor U9907 (N_9907,N_6243,N_7792);
xnor U9908 (N_9908,N_6802,N_8237);
or U9909 (N_9909,N_8435,N_7950);
nor U9910 (N_9910,N_7055,N_8159);
nand U9911 (N_9911,N_8359,N_7518);
or U9912 (N_9912,N_8543,N_8770);
and U9913 (N_9913,N_6303,N_6069);
or U9914 (N_9914,N_7230,N_8765);
nor U9915 (N_9915,N_6162,N_6494);
and U9916 (N_9916,N_7822,N_6047);
and U9917 (N_9917,N_7892,N_8828);
nor U9918 (N_9918,N_7228,N_8797);
and U9919 (N_9919,N_7100,N_8099);
xor U9920 (N_9920,N_6076,N_7870);
nand U9921 (N_9921,N_6749,N_6694);
and U9922 (N_9922,N_8391,N_7880);
xnor U9923 (N_9923,N_6226,N_8128);
xnor U9924 (N_9924,N_6857,N_8311);
and U9925 (N_9925,N_7067,N_8379);
xor U9926 (N_9926,N_7375,N_8214);
nand U9927 (N_9927,N_8826,N_8541);
and U9928 (N_9928,N_7258,N_7839);
nand U9929 (N_9929,N_8571,N_7605);
nor U9930 (N_9930,N_6005,N_8660);
or U9931 (N_9931,N_8196,N_8462);
and U9932 (N_9932,N_8738,N_7887);
xor U9933 (N_9933,N_6199,N_8100);
nand U9934 (N_9934,N_6296,N_6953);
or U9935 (N_9935,N_8121,N_7926);
nor U9936 (N_9936,N_8892,N_6070);
xor U9937 (N_9937,N_7304,N_8490);
xor U9938 (N_9938,N_8993,N_6834);
nor U9939 (N_9939,N_7078,N_8028);
xor U9940 (N_9940,N_7364,N_7399);
or U9941 (N_9941,N_8612,N_6454);
nor U9942 (N_9942,N_6321,N_6994);
and U9943 (N_9943,N_8728,N_6455);
xor U9944 (N_9944,N_7761,N_8670);
or U9945 (N_9945,N_6074,N_7944);
nand U9946 (N_9946,N_7175,N_7951);
xnor U9947 (N_9947,N_7648,N_6746);
and U9948 (N_9948,N_8520,N_6809);
nand U9949 (N_9949,N_7186,N_7261);
nand U9950 (N_9950,N_8168,N_7544);
or U9951 (N_9951,N_6734,N_6458);
nor U9952 (N_9952,N_6065,N_7885);
nand U9953 (N_9953,N_8079,N_7578);
nand U9954 (N_9954,N_7340,N_8365);
or U9955 (N_9955,N_7523,N_8811);
nor U9956 (N_9956,N_7486,N_6705);
xor U9957 (N_9957,N_6747,N_7663);
nand U9958 (N_9958,N_7362,N_7157);
xnor U9959 (N_9959,N_8068,N_6033);
xnor U9960 (N_9960,N_6150,N_7082);
nand U9961 (N_9961,N_8709,N_8655);
or U9962 (N_9962,N_7785,N_8282);
nand U9963 (N_9963,N_8718,N_8198);
nand U9964 (N_9964,N_7461,N_7803);
or U9965 (N_9965,N_8872,N_8884);
or U9966 (N_9966,N_8836,N_7058);
and U9967 (N_9967,N_7905,N_8106);
and U9968 (N_9968,N_7808,N_8584);
nor U9969 (N_9969,N_7460,N_8258);
nor U9970 (N_9970,N_6552,N_6248);
nor U9971 (N_9971,N_6688,N_6434);
and U9972 (N_9972,N_6781,N_8688);
and U9973 (N_9973,N_6520,N_6297);
xnor U9974 (N_9974,N_8777,N_8260);
xnor U9975 (N_9975,N_8271,N_8701);
nor U9976 (N_9976,N_6513,N_7585);
and U9977 (N_9977,N_8257,N_6445);
nand U9978 (N_9978,N_8905,N_6000);
xor U9979 (N_9979,N_8403,N_6884);
or U9980 (N_9980,N_8557,N_6042);
nor U9981 (N_9981,N_6885,N_6642);
and U9982 (N_9982,N_6597,N_8447);
xnor U9983 (N_9983,N_8155,N_8992);
nor U9984 (N_9984,N_6230,N_7982);
and U9985 (N_9985,N_6137,N_7298);
or U9986 (N_9986,N_7427,N_7359);
nor U9987 (N_9987,N_7017,N_8364);
and U9988 (N_9988,N_8124,N_8972);
or U9989 (N_9989,N_6161,N_7385);
nand U9990 (N_9990,N_7613,N_6620);
nand U9991 (N_9991,N_6803,N_8423);
and U9992 (N_9992,N_6573,N_7092);
xnor U9993 (N_9993,N_6253,N_8635);
xor U9994 (N_9994,N_6299,N_6540);
nand U9995 (N_9995,N_6141,N_8269);
nor U9996 (N_9996,N_8366,N_8529);
nand U9997 (N_9997,N_6022,N_6916);
nand U9998 (N_9998,N_6147,N_6326);
and U9999 (N_9999,N_7557,N_7190);
and U10000 (N_10000,N_8671,N_8113);
and U10001 (N_10001,N_7249,N_6726);
xor U10002 (N_10002,N_8202,N_6890);
and U10003 (N_10003,N_7726,N_6700);
or U10004 (N_10004,N_8052,N_7453);
or U10005 (N_10005,N_6646,N_7288);
and U10006 (N_10006,N_6648,N_6586);
nand U10007 (N_10007,N_7000,N_6241);
nor U10008 (N_10008,N_6516,N_7206);
nand U10009 (N_10009,N_6665,N_7773);
nand U10010 (N_10010,N_8874,N_7448);
or U10011 (N_10011,N_6676,N_8844);
nand U10012 (N_10012,N_8558,N_6251);
nand U10013 (N_10013,N_6092,N_8420);
and U10014 (N_10014,N_7115,N_8534);
nand U10015 (N_10015,N_8931,N_7644);
or U10016 (N_10016,N_6101,N_6869);
and U10017 (N_10017,N_8223,N_8832);
nor U10018 (N_10018,N_7492,N_7071);
or U10019 (N_10019,N_8415,N_6232);
xnor U10020 (N_10020,N_6184,N_6995);
nor U10021 (N_10021,N_8119,N_6283);
nand U10022 (N_10022,N_6134,N_8206);
nand U10023 (N_10023,N_6712,N_6225);
or U10024 (N_10024,N_6847,N_8256);
xnor U10025 (N_10025,N_6200,N_6224);
nor U10026 (N_10026,N_8349,N_6959);
xnor U10027 (N_10027,N_6758,N_6999);
or U10028 (N_10028,N_6675,N_6057);
nor U10029 (N_10029,N_8289,N_8180);
nor U10030 (N_10030,N_6839,N_6899);
or U10031 (N_10031,N_8779,N_6052);
or U10032 (N_10032,N_7786,N_8105);
or U10033 (N_10033,N_8117,N_6580);
nor U10034 (N_10034,N_8082,N_7729);
nor U10035 (N_10035,N_8001,N_6213);
nand U10036 (N_10036,N_8115,N_7320);
nor U10037 (N_10037,N_6681,N_8930);
xor U10038 (N_10038,N_8699,N_6381);
and U10039 (N_10039,N_8888,N_6055);
or U10040 (N_10040,N_8929,N_6025);
or U10041 (N_10041,N_7501,N_6278);
xor U10042 (N_10042,N_6944,N_6968);
xor U10043 (N_10043,N_8185,N_6435);
and U10044 (N_10044,N_8210,N_7110);
xnor U10045 (N_10045,N_7285,N_8979);
nor U10046 (N_10046,N_6411,N_8478);
nand U10047 (N_10047,N_6754,N_7272);
nor U10048 (N_10048,N_7538,N_7571);
or U10049 (N_10049,N_6829,N_6568);
xor U10050 (N_10050,N_8547,N_7894);
nand U10051 (N_10051,N_7231,N_8690);
xor U10052 (N_10052,N_6457,N_7246);
xor U10053 (N_10053,N_8918,N_6842);
nor U10054 (N_10054,N_6099,N_6350);
nor U10055 (N_10055,N_8755,N_6163);
or U10056 (N_10056,N_8865,N_8002);
or U10057 (N_10057,N_6366,N_6259);
nor U10058 (N_10058,N_6387,N_7143);
nor U10059 (N_10059,N_7398,N_6368);
and U10060 (N_10060,N_7720,N_7498);
nor U10061 (N_10061,N_8767,N_8518);
xor U10062 (N_10062,N_7549,N_7732);
or U10063 (N_10063,N_7189,N_6174);
xnor U10064 (N_10064,N_7177,N_7633);
nand U10065 (N_10065,N_8203,N_6336);
nand U10066 (N_10066,N_6115,N_7418);
or U10067 (N_10067,N_7414,N_6500);
and U10068 (N_10068,N_7454,N_6583);
nor U10069 (N_10069,N_6946,N_7276);
or U10070 (N_10070,N_8859,N_7108);
and U10071 (N_10071,N_6722,N_8252);
xnor U10072 (N_10072,N_8250,N_7616);
and U10073 (N_10073,N_7208,N_6121);
xnor U10074 (N_10074,N_6367,N_7050);
xor U10075 (N_10075,N_8544,N_6441);
nand U10076 (N_10076,N_7702,N_8742);
and U10077 (N_10077,N_8314,N_8596);
nor U10078 (N_10078,N_8361,N_7054);
xor U10079 (N_10079,N_8053,N_7658);
xor U10080 (N_10080,N_6097,N_8125);
or U10081 (N_10081,N_6073,N_8464);
nand U10082 (N_10082,N_6209,N_7030);
or U10083 (N_10083,N_6724,N_7959);
and U10084 (N_10084,N_6486,N_6343);
and U10085 (N_10085,N_8110,N_8713);
nor U10086 (N_10086,N_7129,N_8317);
and U10087 (N_10087,N_6307,N_7624);
xnor U10088 (N_10088,N_7469,N_7670);
or U10089 (N_10089,N_8746,N_7781);
or U10090 (N_10090,N_8996,N_8280);
or U10091 (N_10091,N_7886,N_8006);
or U10092 (N_10092,N_8757,N_7975);
or U10093 (N_10093,N_6403,N_8489);
or U10094 (N_10094,N_6396,N_8023);
nor U10095 (N_10095,N_7685,N_8283);
or U10096 (N_10096,N_7818,N_7906);
xnor U10097 (N_10097,N_8693,N_6447);
nand U10098 (N_10098,N_7522,N_7494);
and U10099 (N_10099,N_8090,N_8375);
nor U10100 (N_10100,N_6565,N_7631);
nor U10101 (N_10101,N_7562,N_8879);
and U10102 (N_10102,N_6605,N_7088);
or U10103 (N_10103,N_6950,N_6889);
and U10104 (N_10104,N_8678,N_7212);
nor U10105 (N_10105,N_8938,N_6976);
and U10106 (N_10106,N_7226,N_8162);
nand U10107 (N_10107,N_7689,N_8737);
and U10108 (N_10108,N_8877,N_8735);
xor U10109 (N_10109,N_6045,N_6249);
xnor U10110 (N_10110,N_6955,N_7001);
nor U10111 (N_10111,N_7227,N_8488);
nand U10112 (N_10112,N_6246,N_7552);
xnor U10113 (N_10113,N_8803,N_7422);
xnor U10114 (N_10114,N_7826,N_8248);
nor U10115 (N_10115,N_7888,N_6854);
nor U10116 (N_10116,N_7215,N_6564);
nor U10117 (N_10117,N_7488,N_8426);
nor U10118 (N_10118,N_7712,N_7163);
xor U10119 (N_10119,N_7021,N_8284);
xor U10120 (N_10120,N_8200,N_8648);
xnor U10121 (N_10121,N_8228,N_8229);
nor U10122 (N_10122,N_8748,N_7567);
xnor U10123 (N_10123,N_7615,N_7216);
nor U10124 (N_10124,N_7200,N_7112);
xor U10125 (N_10125,N_6041,N_6613);
and U10126 (N_10126,N_7943,N_6276);
nand U10127 (N_10127,N_7273,N_8666);
xor U10128 (N_10128,N_6939,N_8616);
nand U10129 (N_10129,N_7998,N_6481);
xnor U10130 (N_10130,N_7601,N_6682);
or U10131 (N_10131,N_7817,N_8561);
nor U10132 (N_10132,N_7727,N_8897);
xor U10133 (N_10133,N_8328,N_8695);
nand U10134 (N_10134,N_7863,N_6281);
nor U10135 (N_10135,N_8016,N_8724);
and U10136 (N_10136,N_8672,N_6877);
and U10137 (N_10137,N_6561,N_6723);
nand U10138 (N_10138,N_8942,N_7804);
nand U10139 (N_10139,N_8667,N_8372);
nand U10140 (N_10140,N_6756,N_6390);
nand U10141 (N_10141,N_8810,N_8498);
and U10142 (N_10142,N_7286,N_6949);
nand U10143 (N_10143,N_6144,N_8094);
nor U10144 (N_10144,N_7475,N_8593);
or U10145 (N_10145,N_6132,N_7656);
xnor U10146 (N_10146,N_6822,N_8791);
xnor U10147 (N_10147,N_8985,N_7009);
xor U10148 (N_10148,N_6930,N_7281);
nand U10149 (N_10149,N_6807,N_6425);
and U10150 (N_10150,N_6898,N_8633);
or U10151 (N_10151,N_8926,N_8569);
and U10152 (N_10152,N_8350,N_8508);
xor U10153 (N_10153,N_6732,N_8936);
xnor U10154 (N_10154,N_7314,N_7120);
and U10155 (N_10155,N_8209,N_8409);
or U10156 (N_10156,N_8654,N_6261);
or U10157 (N_10157,N_6420,N_7554);
nor U10158 (N_10158,N_6095,N_6559);
or U10159 (N_10159,N_7879,N_7769);
or U10160 (N_10160,N_6601,N_8970);
and U10161 (N_10161,N_8312,N_7268);
nor U10162 (N_10162,N_8147,N_8556);
or U10163 (N_10163,N_6214,N_7649);
nand U10164 (N_10164,N_6363,N_6413);
nand U10165 (N_10165,N_7293,N_8568);
nor U10166 (N_10166,N_8679,N_6355);
xnor U10167 (N_10167,N_6795,N_7307);
nor U10168 (N_10168,N_8536,N_6331);
nor U10169 (N_10169,N_6378,N_6346);
nand U10170 (N_10170,N_8224,N_8705);
xnor U10171 (N_10171,N_7746,N_6860);
and U10172 (N_10172,N_7929,N_7128);
xor U10173 (N_10173,N_7024,N_8590);
and U10174 (N_10174,N_8567,N_7533);
and U10175 (N_10175,N_6727,N_7070);
nor U10176 (N_10176,N_7308,N_6179);
xor U10177 (N_10177,N_8740,N_7901);
nor U10178 (N_10178,N_7282,N_6887);
nor U10179 (N_10179,N_8870,N_8064);
or U10180 (N_10180,N_6460,N_6718);
nor U10181 (N_10181,N_7350,N_8454);
or U10182 (N_10182,N_6409,N_7650);
nand U10183 (N_10183,N_7911,N_7028);
xor U10184 (N_10184,N_8708,N_7895);
nand U10185 (N_10185,N_8204,N_8595);
nand U10186 (N_10186,N_7532,N_6757);
nor U10187 (N_10187,N_6113,N_6988);
nand U10188 (N_10188,N_8265,N_8597);
xor U10189 (N_10189,N_6406,N_6624);
xnor U10190 (N_10190,N_7968,N_7156);
or U10191 (N_10191,N_6478,N_8241);
nand U10192 (N_10192,N_7435,N_8073);
nor U10193 (N_10193,N_7653,N_6240);
xnor U10194 (N_10194,N_8069,N_8605);
or U10195 (N_10195,N_6024,N_7806);
nand U10196 (N_10196,N_6963,N_6840);
nor U10197 (N_10197,N_6921,N_8820);
xnor U10198 (N_10198,N_8067,N_6893);
xnor U10199 (N_10199,N_7445,N_8759);
xnor U10200 (N_10200,N_8142,N_6038);
nand U10201 (N_10201,N_8956,N_8680);
or U10202 (N_10202,N_8276,N_8480);
and U10203 (N_10203,N_7851,N_6922);
nor U10204 (N_10204,N_6371,N_8585);
and U10205 (N_10205,N_7470,N_7386);
xnor U10206 (N_10206,N_8796,N_6509);
or U10207 (N_10207,N_6492,N_8226);
nor U10208 (N_10208,N_8636,N_8037);
and U10209 (N_10209,N_8760,N_6079);
nor U10210 (N_10210,N_6234,N_7563);
or U10211 (N_10211,N_7677,N_6462);
xnor U10212 (N_10212,N_7565,N_8154);
and U10213 (N_10213,N_6430,N_7980);
xor U10214 (N_10214,N_6505,N_6833);
or U10215 (N_10215,N_7703,N_8665);
and U10216 (N_10216,N_8487,N_6961);
nand U10217 (N_10217,N_6591,N_6317);
nand U10218 (N_10218,N_7719,N_7195);
nand U10219 (N_10219,N_6761,N_6882);
nand U10220 (N_10220,N_6850,N_7972);
xor U10221 (N_10221,N_6741,N_8387);
nand U10222 (N_10222,N_6290,N_8513);
xor U10223 (N_10223,N_6456,N_6879);
nand U10224 (N_10224,N_6472,N_7986);
nand U10225 (N_10225,N_6136,N_8007);
or U10226 (N_10226,N_6526,N_6728);
nand U10227 (N_10227,N_8272,N_7010);
nand U10228 (N_10228,N_7134,N_6710);
and U10229 (N_10229,N_8941,N_8307);
nand U10230 (N_10230,N_6760,N_7357);
and U10231 (N_10231,N_8170,N_8381);
nand U10232 (N_10232,N_6007,N_7725);
nor U10233 (N_10233,N_7520,N_7467);
nor U10234 (N_10234,N_6534,N_8786);
and U10235 (N_10235,N_8166,N_6267);
xnor U10236 (N_10236,N_8221,N_8983);
or U10237 (N_10237,N_6846,N_7547);
nor U10238 (N_10238,N_8441,N_7138);
nand U10239 (N_10239,N_6236,N_8856);
or U10240 (N_10240,N_8044,N_8389);
or U10241 (N_10241,N_7586,N_7582);
nand U10242 (N_10242,N_6444,N_6449);
xor U10243 (N_10243,N_7483,N_8179);
nand U10244 (N_10244,N_7168,N_8253);
nand U10245 (N_10245,N_7989,N_7833);
and U10246 (N_10246,N_8255,N_6180);
and U10247 (N_10247,N_8098,N_6745);
nor U10248 (N_10248,N_8242,N_7647);
nor U10249 (N_10249,N_8517,N_8973);
xor U10250 (N_10250,N_6280,N_6203);
nand U10251 (N_10251,N_6769,N_6043);
nor U10252 (N_10252,N_7821,N_7191);
or U10253 (N_10253,N_6348,N_6900);
nand U10254 (N_10254,N_7008,N_7089);
or U10255 (N_10255,N_8780,N_6684);
or U10256 (N_10256,N_8285,N_8362);
nor U10257 (N_10257,N_8380,N_7679);
nor U10258 (N_10258,N_6427,N_6011);
xnor U10259 (N_10259,N_7409,N_8542);
nand U10260 (N_10260,N_7759,N_6905);
nand U10261 (N_10261,N_8208,N_6986);
nor U10262 (N_10262,N_6048,N_6330);
nor U10263 (N_10263,N_7775,N_7898);
nand U10264 (N_10264,N_7716,N_8267);
xor U10265 (N_10265,N_7383,N_7125);
xor U10266 (N_10266,N_8156,N_6415);
xnor U10267 (N_10267,N_6554,N_7004);
xor U10268 (N_10268,N_7923,N_7753);
nor U10269 (N_10269,N_8902,N_8921);
and U10270 (N_10270,N_8315,N_7509);
nor U10271 (N_10271,N_7066,N_7199);
xor U10272 (N_10272,N_7337,N_7816);
xnor U10273 (N_10273,N_6322,N_8235);
xor U10274 (N_10274,N_7325,N_7737);
xor U10275 (N_10275,N_7698,N_7283);
xor U10276 (N_10276,N_8539,N_6541);
nor U10277 (N_10277,N_7969,N_7378);
or U10278 (N_10278,N_8201,N_7015);
xor U10279 (N_10279,N_7196,N_6895);
or U10280 (N_10280,N_6793,N_7442);
xor U10281 (N_10281,N_8946,N_8148);
nand U10282 (N_10282,N_6629,N_8721);
and U10283 (N_10283,N_8323,N_7119);
or U10284 (N_10284,N_7597,N_6765);
nand U10285 (N_10285,N_8646,N_8457);
nand U10286 (N_10286,N_6551,N_8192);
and U10287 (N_10287,N_8948,N_8842);
nand U10288 (N_10288,N_6560,N_6777);
nand U10289 (N_10289,N_7960,N_6031);
nor U10290 (N_10290,N_7311,N_7674);
nand U10291 (N_10291,N_6119,N_7233);
or U10292 (N_10292,N_6519,N_8873);
nor U10293 (N_10293,N_8118,N_7747);
nand U10294 (N_10294,N_6262,N_6155);
nor U10295 (N_10295,N_7525,N_7680);
xnor U10296 (N_10296,N_8451,N_7700);
and U10297 (N_10297,N_7330,N_7794);
or U10298 (N_10298,N_7572,N_8163);
nor U10299 (N_10299,N_6067,N_6061);
nor U10300 (N_10300,N_6659,N_8161);
xor U10301 (N_10301,N_6985,N_6098);
nand U10302 (N_10302,N_7173,N_8354);
nand U10303 (N_10303,N_8238,N_8395);
and U10304 (N_10304,N_7366,N_7922);
nor U10305 (N_10305,N_8344,N_7641);
nor U10306 (N_10306,N_7033,N_8553);
nand U10307 (N_10307,N_8947,N_6463);
xnor U10308 (N_10308,N_7417,N_8676);
nand U10309 (N_10309,N_8074,N_6751);
or U10310 (N_10310,N_8378,N_8504);
nand U10311 (N_10311,N_8132,N_8057);
nor U10312 (N_10312,N_7749,N_6217);
xnor U10313 (N_10313,N_8456,N_6302);
xor U10314 (N_10314,N_6971,N_7580);
nand U10315 (N_10315,N_7098,N_7628);
xor U10316 (N_10316,N_8962,N_7676);
or U10317 (N_10317,N_6623,N_6797);
nand U10318 (N_10318,N_7891,N_6843);
and U10319 (N_10319,N_7290,N_6271);
xnor U10320 (N_10320,N_8329,N_6660);
or U10321 (N_10321,N_8026,N_8495);
or U10322 (N_10322,N_6050,N_6498);
and U10323 (N_10323,N_7087,N_7495);
xor U10324 (N_10324,N_8012,N_8559);
nor U10325 (N_10325,N_7614,N_7203);
or U10326 (N_10326,N_6361,N_6689);
xor U10327 (N_10327,N_6394,N_6917);
nand U10328 (N_10328,N_6265,N_7841);
and U10329 (N_10329,N_8401,N_7504);
nand U10330 (N_10330,N_7681,N_7802);
nand U10331 (N_10331,N_7784,N_8858);
nor U10332 (N_10332,N_8164,N_6592);
nand U10333 (N_10333,N_8171,N_6641);
and U10334 (N_10334,N_8137,N_6992);
and U10335 (N_10335,N_7145,N_8492);
xnor U10336 (N_10336,N_6228,N_6138);
nand U10337 (N_10337,N_7240,N_6166);
nand U10338 (N_10338,N_7368,N_6662);
xor U10339 (N_10339,N_7987,N_6606);
nor U10340 (N_10340,N_6989,N_7608);
and U10341 (N_10341,N_8066,N_6480);
xnor U10342 (N_10342,N_8975,N_8191);
nand U10343 (N_10343,N_6844,N_7123);
or U10344 (N_10344,N_6545,N_7519);
nand U10345 (N_10345,N_8914,N_8397);
nor U10346 (N_10346,N_8754,N_7754);
and U10347 (N_10347,N_7569,N_8318);
or U10348 (N_10348,N_8739,N_6078);
or U10349 (N_10349,N_6145,N_8268);
nor U10350 (N_10350,N_7857,N_6982);
and U10351 (N_10351,N_6446,N_8408);
and U10352 (N_10352,N_7184,N_6483);
and U10353 (N_10353,N_6858,N_6535);
or U10354 (N_10354,N_6402,N_8396);
and U10355 (N_10355,N_8977,N_7410);
nand U10356 (N_10356,N_7387,N_8603);
nand U10357 (N_10357,N_6678,N_7135);
and U10358 (N_10358,N_7715,N_6391);
nor U10359 (N_10359,N_7310,N_7256);
and U10360 (N_10360,N_6066,N_7349);
or U10361 (N_10361,N_8908,N_6169);
nor U10362 (N_10362,N_7838,N_7022);
or U10363 (N_10363,N_8795,N_6801);
nand U10364 (N_10364,N_7037,N_8989);
nand U10365 (N_10365,N_7609,N_6669);
xor U10366 (N_10366,N_7468,N_8339);
nand U10367 (N_10367,N_6941,N_8608);
nand U10368 (N_10368,N_7449,N_8514);
and U10369 (N_10369,N_7558,N_6909);
and U10370 (N_10370,N_6053,N_6644);
or U10371 (N_10371,N_7626,N_7369);
or U10372 (N_10372,N_7264,N_8928);
or U10373 (N_10373,N_7583,N_7406);
and U10374 (N_10374,N_6861,N_8563);
nand U10375 (N_10375,N_6398,N_7531);
and U10376 (N_10376,N_7765,N_8629);
or U10377 (N_10377,N_8004,N_7687);
xor U10378 (N_10378,N_8178,N_6032);
xnor U10379 (N_10379,N_8808,N_6919);
nand U10380 (N_10380,N_6821,N_8932);
or U10381 (N_10381,N_6713,N_7284);
or U10382 (N_10382,N_7860,N_8005);
xor U10383 (N_10383,N_8443,N_7220);
and U10384 (N_10384,N_6301,N_7756);
and U10385 (N_10385,N_6451,N_7606);
nand U10386 (N_10386,N_8402,N_7436);
nor U10387 (N_10387,N_8342,N_8707);
or U10388 (N_10388,N_8878,N_8726);
or U10389 (N_10389,N_8003,N_7462);
nand U10390 (N_10390,N_6805,N_8298);
and U10391 (N_10391,N_8641,N_6549);
nor U10392 (N_10392,N_8855,N_7169);
xnor U10393 (N_10393,N_7983,N_7013);
xor U10394 (N_10394,N_8862,N_6507);
or U10395 (N_10395,N_6006,N_6614);
nor U10396 (N_10396,N_6862,N_7373);
and U10397 (N_10397,N_6465,N_7757);
xor U10398 (N_10398,N_7485,N_6049);
nand U10399 (N_10399,N_7025,N_6582);
or U10400 (N_10400,N_7831,N_7878);
nor U10401 (N_10401,N_8528,N_7117);
nor U10402 (N_10402,N_7978,N_8014);
nor U10403 (N_10403,N_8448,N_6382);
nor U10404 (N_10404,N_8091,N_8747);
nand U10405 (N_10405,N_8964,N_8594);
or U10406 (N_10406,N_7573,N_6308);
xor U10407 (N_10407,N_6086,N_7524);
nand U10408 (N_10408,N_7400,N_6314);
or U10409 (N_10409,N_7612,N_6638);
nand U10410 (N_10410,N_6244,N_8940);
nand U10411 (N_10411,N_8134,N_6129);
nor U10412 (N_10412,N_8846,N_7918);
nand U10413 (N_10413,N_6626,N_8647);
nor U10414 (N_10414,N_6305,N_6400);
and U10415 (N_10415,N_8126,N_7141);
xnor U10416 (N_10416,N_7660,N_6106);
nor U10417 (N_10417,N_6448,N_7564);
xor U10418 (N_10418,N_8305,N_6365);
or U10419 (N_10419,N_8995,N_6926);
xor U10420 (N_10420,N_6120,N_8051);
nand U10421 (N_10421,N_8600,N_7527);
and U10422 (N_10422,N_8368,N_7854);
or U10423 (N_10423,N_8225,N_7235);
xnor U10424 (N_10424,N_8466,N_6388);
or U10425 (N_10425,N_7393,N_7957);
nor U10426 (N_10426,N_8510,N_7335);
nor U10427 (N_10427,N_6556,N_7846);
nand U10428 (N_10428,N_8876,N_8548);
and U10429 (N_10429,N_7122,N_8382);
nand U10430 (N_10430,N_8775,N_8424);
and U10431 (N_10431,N_8363,N_8696);
and U10432 (N_10432,N_6286,N_6018);
nor U10433 (N_10433,N_8501,N_6021);
xnor U10434 (N_10434,N_7876,N_6855);
nand U10435 (N_10435,N_6428,N_8262);
xnor U10436 (N_10436,N_6674,N_6800);
nand U10437 (N_10437,N_6375,N_7412);
or U10438 (N_10438,N_8901,N_8981);
and U10439 (N_10439,N_7883,N_6036);
nand U10440 (N_10440,N_7005,N_7581);
nand U10441 (N_10441,N_6487,N_8883);
or U10442 (N_10442,N_6389,N_6523);
nor U10443 (N_10443,N_6131,N_7701);
nor U10444 (N_10444,N_7767,N_8607);
nor U10445 (N_10445,N_8860,N_6990);
nand U10446 (N_10446,N_6875,N_6215);
nor U10447 (N_10447,N_7932,N_6912);
nor U10448 (N_10448,N_7093,N_6176);
nand U10449 (N_10449,N_8493,N_7762);
and U10450 (N_10450,N_6075,N_8442);
nand U10451 (N_10451,N_7012,N_7471);
and U10452 (N_10452,N_6647,N_6020);
xnor U10453 (N_10453,N_7336,N_8891);
and U10454 (N_10454,N_6210,N_8579);
nor U10455 (N_10455,N_6585,N_7964);
nand U10456 (N_10456,N_8506,N_6925);
nor U10457 (N_10457,N_6599,N_8195);
xor U10458 (N_10458,N_6473,N_6029);
nand U10459 (N_10459,N_8356,N_8130);
nand U10460 (N_10460,N_6288,N_7777);
nor U10461 (N_10461,N_7053,N_6418);
xor U10462 (N_10462,N_7309,N_7875);
nor U10463 (N_10463,N_7636,N_8697);
xor U10464 (N_10464,N_7139,N_8089);
and U10465 (N_10465,N_7457,N_6338);
nand U10466 (N_10466,N_6268,N_7789);
or U10467 (N_10467,N_6691,N_7419);
nor U10468 (N_10468,N_6566,N_8953);
nor U10469 (N_10469,N_6524,N_8834);
or U10470 (N_10470,N_7502,N_6285);
xor U10471 (N_10471,N_8974,N_7805);
nor U10472 (N_10472,N_8486,N_8041);
and U10473 (N_10473,N_7149,N_8428);
xnor U10474 (N_10474,N_6915,N_8332);
or U10475 (N_10475,N_7503,N_7780);
xnor U10476 (N_10476,N_6257,N_8353);
xor U10477 (N_10477,N_7260,N_6954);
xnor U10478 (N_10478,N_8706,N_6956);
nor U10479 (N_10479,N_8904,N_7783);
or U10480 (N_10480,N_8324,N_8310);
nor U10481 (N_10481,N_8333,N_6178);
or U10482 (N_10482,N_6703,N_6374);
nor U10483 (N_10483,N_7809,N_7797);
nand U10484 (N_10484,N_6328,N_6835);
nor U10485 (N_10485,N_6143,N_7153);
and U10486 (N_10486,N_6600,N_7257);
xor U10487 (N_10487,N_6499,N_8060);
or U10488 (N_10488,N_7170,N_6607);
nand U10489 (N_10489,N_6615,N_7452);
nor U10490 (N_10490,N_7085,N_6706);
and U10491 (N_10491,N_7815,N_6311);
nand U10492 (N_10492,N_7595,N_7023);
and U10493 (N_10493,N_8337,N_6686);
nand U10494 (N_10494,N_6589,N_6377);
nand U10495 (N_10495,N_7496,N_8851);
nor U10496 (N_10496,N_7006,N_6584);
xnor U10497 (N_10497,N_8900,N_7881);
nor U10498 (N_10498,N_7363,N_8537);
and U10499 (N_10499,N_8287,N_7219);
or U10500 (N_10500,N_6666,N_7615);
or U10501 (N_10501,N_8678,N_7731);
and U10502 (N_10502,N_7780,N_7188);
nor U10503 (N_10503,N_8443,N_8030);
and U10504 (N_10504,N_7317,N_7731);
nand U10505 (N_10505,N_7640,N_8449);
xnor U10506 (N_10506,N_6519,N_7716);
nor U10507 (N_10507,N_6279,N_6926);
nand U10508 (N_10508,N_6697,N_6449);
or U10509 (N_10509,N_8493,N_6906);
or U10510 (N_10510,N_8418,N_6496);
or U10511 (N_10511,N_8281,N_6814);
or U10512 (N_10512,N_6135,N_6454);
nor U10513 (N_10513,N_7336,N_8617);
nand U10514 (N_10514,N_6110,N_8885);
or U10515 (N_10515,N_6083,N_7065);
nor U10516 (N_10516,N_6819,N_6431);
nor U10517 (N_10517,N_8603,N_6090);
and U10518 (N_10518,N_7572,N_7792);
xnor U10519 (N_10519,N_7621,N_6499);
or U10520 (N_10520,N_8041,N_8284);
and U10521 (N_10521,N_6483,N_6789);
or U10522 (N_10522,N_6614,N_8097);
or U10523 (N_10523,N_8783,N_8270);
and U10524 (N_10524,N_8895,N_7382);
and U10525 (N_10525,N_6990,N_6984);
nor U10526 (N_10526,N_7206,N_7682);
nand U10527 (N_10527,N_8814,N_7952);
nor U10528 (N_10528,N_7554,N_7829);
nor U10529 (N_10529,N_8122,N_6552);
and U10530 (N_10530,N_6727,N_7524);
xnor U10531 (N_10531,N_7142,N_7617);
nor U10532 (N_10532,N_8775,N_7902);
nand U10533 (N_10533,N_8799,N_6366);
or U10534 (N_10534,N_6100,N_6214);
nand U10535 (N_10535,N_8754,N_8831);
nor U10536 (N_10536,N_7914,N_8708);
nand U10537 (N_10537,N_6269,N_7714);
nor U10538 (N_10538,N_6203,N_8308);
or U10539 (N_10539,N_6084,N_7913);
xnor U10540 (N_10540,N_8018,N_6719);
or U10541 (N_10541,N_6577,N_8434);
nand U10542 (N_10542,N_6123,N_7078);
and U10543 (N_10543,N_7445,N_8701);
or U10544 (N_10544,N_8286,N_6522);
xnor U10545 (N_10545,N_7483,N_6065);
or U10546 (N_10546,N_7290,N_8312);
nand U10547 (N_10547,N_6364,N_7248);
or U10548 (N_10548,N_8666,N_7565);
and U10549 (N_10549,N_8775,N_7593);
nand U10550 (N_10550,N_8948,N_6338);
nand U10551 (N_10551,N_8748,N_6502);
and U10552 (N_10552,N_7015,N_6653);
nor U10553 (N_10553,N_6815,N_7805);
nor U10554 (N_10554,N_8307,N_7787);
and U10555 (N_10555,N_6825,N_6720);
nand U10556 (N_10556,N_8714,N_7590);
nand U10557 (N_10557,N_8125,N_7489);
nand U10558 (N_10558,N_8930,N_6013);
xnor U10559 (N_10559,N_7693,N_8747);
nor U10560 (N_10560,N_7593,N_8147);
nand U10561 (N_10561,N_7323,N_6862);
nand U10562 (N_10562,N_7276,N_8433);
xnor U10563 (N_10563,N_8479,N_7586);
xnor U10564 (N_10564,N_8188,N_7973);
and U10565 (N_10565,N_7877,N_7019);
or U10566 (N_10566,N_6665,N_6216);
and U10567 (N_10567,N_8480,N_6174);
xor U10568 (N_10568,N_6426,N_7551);
and U10569 (N_10569,N_7008,N_6166);
or U10570 (N_10570,N_8540,N_7295);
or U10571 (N_10571,N_8484,N_7404);
and U10572 (N_10572,N_7234,N_8406);
or U10573 (N_10573,N_8814,N_6528);
xnor U10574 (N_10574,N_7382,N_7298);
nor U10575 (N_10575,N_8720,N_8301);
or U10576 (N_10576,N_6036,N_7857);
xnor U10577 (N_10577,N_7106,N_8635);
xor U10578 (N_10578,N_7271,N_7265);
and U10579 (N_10579,N_8328,N_7766);
nor U10580 (N_10580,N_6243,N_7655);
nor U10581 (N_10581,N_8173,N_8769);
nor U10582 (N_10582,N_6115,N_7318);
nand U10583 (N_10583,N_6145,N_7103);
nand U10584 (N_10584,N_6158,N_6553);
xnor U10585 (N_10585,N_6440,N_8901);
or U10586 (N_10586,N_7606,N_6586);
xnor U10587 (N_10587,N_7951,N_6780);
xnor U10588 (N_10588,N_6736,N_6804);
xor U10589 (N_10589,N_7755,N_6429);
nand U10590 (N_10590,N_6831,N_7618);
and U10591 (N_10591,N_7337,N_8298);
and U10592 (N_10592,N_7238,N_8113);
xor U10593 (N_10593,N_7279,N_8650);
nand U10594 (N_10594,N_6528,N_8543);
xnor U10595 (N_10595,N_6456,N_6720);
or U10596 (N_10596,N_7160,N_8585);
and U10597 (N_10597,N_6027,N_8097);
nand U10598 (N_10598,N_6892,N_7277);
nor U10599 (N_10599,N_7015,N_6645);
nand U10600 (N_10600,N_7789,N_6253);
xnor U10601 (N_10601,N_6894,N_8478);
and U10602 (N_10602,N_6125,N_7210);
and U10603 (N_10603,N_7101,N_8298);
nand U10604 (N_10604,N_8652,N_6253);
nand U10605 (N_10605,N_6346,N_8597);
or U10606 (N_10606,N_7550,N_7998);
nand U10607 (N_10607,N_8609,N_7690);
xnor U10608 (N_10608,N_7172,N_8150);
nor U10609 (N_10609,N_7331,N_7232);
nand U10610 (N_10610,N_7159,N_6217);
or U10611 (N_10611,N_8696,N_8323);
or U10612 (N_10612,N_6495,N_6172);
or U10613 (N_10613,N_7279,N_8041);
and U10614 (N_10614,N_6547,N_8257);
nor U10615 (N_10615,N_8426,N_7767);
nor U10616 (N_10616,N_6893,N_7515);
xnor U10617 (N_10617,N_8825,N_6501);
and U10618 (N_10618,N_6360,N_7729);
nand U10619 (N_10619,N_6845,N_6968);
nand U10620 (N_10620,N_6819,N_7816);
nand U10621 (N_10621,N_6399,N_7389);
nor U10622 (N_10622,N_8812,N_6777);
or U10623 (N_10623,N_7793,N_6675);
nand U10624 (N_10624,N_8374,N_8325);
nand U10625 (N_10625,N_8049,N_8414);
xnor U10626 (N_10626,N_6160,N_7885);
or U10627 (N_10627,N_6872,N_7663);
nor U10628 (N_10628,N_7098,N_6627);
xnor U10629 (N_10629,N_6662,N_7728);
xor U10630 (N_10630,N_6710,N_7151);
nand U10631 (N_10631,N_8967,N_7260);
nor U10632 (N_10632,N_6229,N_8556);
nor U10633 (N_10633,N_7911,N_8341);
nor U10634 (N_10634,N_6902,N_6684);
nand U10635 (N_10635,N_7359,N_8779);
nor U10636 (N_10636,N_6560,N_7973);
xnor U10637 (N_10637,N_6651,N_6073);
nand U10638 (N_10638,N_8454,N_8016);
nand U10639 (N_10639,N_8573,N_6869);
nor U10640 (N_10640,N_6728,N_8299);
or U10641 (N_10641,N_6283,N_8163);
xnor U10642 (N_10642,N_6368,N_6966);
nor U10643 (N_10643,N_7781,N_8903);
nand U10644 (N_10644,N_7690,N_6724);
nor U10645 (N_10645,N_7544,N_7352);
xor U10646 (N_10646,N_8981,N_8963);
nor U10647 (N_10647,N_7850,N_6736);
xor U10648 (N_10648,N_6579,N_8396);
or U10649 (N_10649,N_7342,N_8548);
and U10650 (N_10650,N_6783,N_7428);
and U10651 (N_10651,N_6911,N_8515);
nor U10652 (N_10652,N_7211,N_6342);
nand U10653 (N_10653,N_8142,N_8357);
or U10654 (N_10654,N_6168,N_6139);
nand U10655 (N_10655,N_7471,N_6117);
nor U10656 (N_10656,N_7726,N_7219);
or U10657 (N_10657,N_6911,N_7376);
or U10658 (N_10658,N_6178,N_7394);
xnor U10659 (N_10659,N_7279,N_7185);
and U10660 (N_10660,N_7622,N_8912);
and U10661 (N_10661,N_7797,N_7588);
or U10662 (N_10662,N_6868,N_7101);
nand U10663 (N_10663,N_7125,N_6385);
nand U10664 (N_10664,N_6324,N_6506);
nor U10665 (N_10665,N_6371,N_6639);
nand U10666 (N_10666,N_7860,N_7255);
or U10667 (N_10667,N_8232,N_6377);
xnor U10668 (N_10668,N_6583,N_8564);
nand U10669 (N_10669,N_6662,N_7827);
or U10670 (N_10670,N_8724,N_6014);
and U10671 (N_10671,N_6627,N_7580);
xnor U10672 (N_10672,N_6881,N_6961);
xnor U10673 (N_10673,N_6075,N_6206);
nand U10674 (N_10674,N_7242,N_6838);
or U10675 (N_10675,N_6478,N_7884);
or U10676 (N_10676,N_6739,N_8948);
nor U10677 (N_10677,N_7107,N_7284);
and U10678 (N_10678,N_7936,N_6505);
or U10679 (N_10679,N_6339,N_7054);
nor U10680 (N_10680,N_8688,N_7211);
and U10681 (N_10681,N_6778,N_8913);
xor U10682 (N_10682,N_7232,N_8883);
nor U10683 (N_10683,N_6169,N_8622);
xor U10684 (N_10684,N_8685,N_8307);
and U10685 (N_10685,N_7211,N_6437);
and U10686 (N_10686,N_7876,N_7708);
nor U10687 (N_10687,N_6727,N_8941);
xor U10688 (N_10688,N_8837,N_7537);
nand U10689 (N_10689,N_6844,N_7336);
and U10690 (N_10690,N_8478,N_6536);
nor U10691 (N_10691,N_7636,N_7968);
nor U10692 (N_10692,N_7553,N_8332);
or U10693 (N_10693,N_6600,N_7053);
nand U10694 (N_10694,N_8367,N_8472);
and U10695 (N_10695,N_7383,N_6078);
nor U10696 (N_10696,N_8147,N_8858);
or U10697 (N_10697,N_7540,N_8759);
and U10698 (N_10698,N_6112,N_8857);
nor U10699 (N_10699,N_6253,N_6674);
or U10700 (N_10700,N_6996,N_8563);
nand U10701 (N_10701,N_7037,N_7920);
xnor U10702 (N_10702,N_8431,N_6597);
nand U10703 (N_10703,N_7794,N_7298);
nor U10704 (N_10704,N_6799,N_7208);
xnor U10705 (N_10705,N_6766,N_7111);
nor U10706 (N_10706,N_8168,N_6831);
nand U10707 (N_10707,N_8549,N_8405);
nor U10708 (N_10708,N_7567,N_7693);
nand U10709 (N_10709,N_8240,N_8665);
xor U10710 (N_10710,N_8231,N_6382);
nor U10711 (N_10711,N_8493,N_8649);
nor U10712 (N_10712,N_6295,N_6026);
nand U10713 (N_10713,N_6127,N_6995);
nand U10714 (N_10714,N_8179,N_7767);
nor U10715 (N_10715,N_7082,N_7909);
and U10716 (N_10716,N_8746,N_6417);
xor U10717 (N_10717,N_8137,N_7757);
xor U10718 (N_10718,N_8326,N_8604);
or U10719 (N_10719,N_7665,N_6673);
and U10720 (N_10720,N_7804,N_6052);
or U10721 (N_10721,N_8490,N_8892);
and U10722 (N_10722,N_6065,N_6395);
nor U10723 (N_10723,N_6116,N_8808);
and U10724 (N_10724,N_6724,N_7970);
nor U10725 (N_10725,N_7400,N_6566);
or U10726 (N_10726,N_8215,N_8320);
or U10727 (N_10727,N_8518,N_7483);
nor U10728 (N_10728,N_8717,N_8542);
xnor U10729 (N_10729,N_7579,N_8272);
or U10730 (N_10730,N_7872,N_8754);
xor U10731 (N_10731,N_8808,N_6321);
nor U10732 (N_10732,N_7828,N_8586);
and U10733 (N_10733,N_8517,N_7281);
nor U10734 (N_10734,N_6960,N_6577);
nand U10735 (N_10735,N_7167,N_7820);
or U10736 (N_10736,N_8365,N_7804);
xnor U10737 (N_10737,N_7287,N_7871);
and U10738 (N_10738,N_8648,N_8286);
and U10739 (N_10739,N_6061,N_6549);
and U10740 (N_10740,N_7743,N_6822);
nor U10741 (N_10741,N_8533,N_8106);
or U10742 (N_10742,N_8693,N_8719);
nand U10743 (N_10743,N_8931,N_8788);
nand U10744 (N_10744,N_8684,N_6357);
and U10745 (N_10745,N_8870,N_7508);
xnor U10746 (N_10746,N_8001,N_6944);
or U10747 (N_10747,N_7825,N_8800);
or U10748 (N_10748,N_7312,N_8465);
or U10749 (N_10749,N_6297,N_8614);
nand U10750 (N_10750,N_8716,N_7741);
or U10751 (N_10751,N_7172,N_6452);
xnor U10752 (N_10752,N_7269,N_6035);
nand U10753 (N_10753,N_7700,N_6867);
or U10754 (N_10754,N_7866,N_6887);
nor U10755 (N_10755,N_8150,N_7027);
or U10756 (N_10756,N_7133,N_7579);
or U10757 (N_10757,N_6189,N_8434);
xnor U10758 (N_10758,N_7179,N_7490);
nand U10759 (N_10759,N_7454,N_7037);
or U10760 (N_10760,N_8868,N_8267);
nand U10761 (N_10761,N_8652,N_6749);
and U10762 (N_10762,N_8625,N_8800);
nand U10763 (N_10763,N_8413,N_7756);
xor U10764 (N_10764,N_8127,N_8410);
nand U10765 (N_10765,N_6207,N_7644);
nand U10766 (N_10766,N_8963,N_6997);
xor U10767 (N_10767,N_6368,N_8029);
nand U10768 (N_10768,N_6987,N_6292);
and U10769 (N_10769,N_7279,N_7871);
nand U10770 (N_10770,N_8048,N_6873);
or U10771 (N_10771,N_7996,N_8036);
nand U10772 (N_10772,N_6052,N_6561);
nand U10773 (N_10773,N_7884,N_6939);
nand U10774 (N_10774,N_8264,N_7222);
nor U10775 (N_10775,N_7273,N_6506);
nor U10776 (N_10776,N_8851,N_8449);
or U10777 (N_10777,N_8750,N_7342);
xor U10778 (N_10778,N_6657,N_6557);
nor U10779 (N_10779,N_6245,N_8098);
xor U10780 (N_10780,N_7339,N_8863);
and U10781 (N_10781,N_8427,N_6006);
xnor U10782 (N_10782,N_8592,N_8275);
and U10783 (N_10783,N_8178,N_6780);
xnor U10784 (N_10784,N_8598,N_8966);
and U10785 (N_10785,N_6982,N_6729);
or U10786 (N_10786,N_8982,N_7988);
nor U10787 (N_10787,N_7917,N_7076);
and U10788 (N_10788,N_6340,N_8051);
nand U10789 (N_10789,N_8020,N_7763);
nor U10790 (N_10790,N_8192,N_7420);
nor U10791 (N_10791,N_7139,N_8234);
nand U10792 (N_10792,N_8034,N_6219);
nand U10793 (N_10793,N_7070,N_6471);
and U10794 (N_10794,N_6115,N_7259);
nand U10795 (N_10795,N_8132,N_8526);
or U10796 (N_10796,N_7942,N_8782);
nand U10797 (N_10797,N_6131,N_8167);
nor U10798 (N_10798,N_8594,N_8428);
nand U10799 (N_10799,N_6132,N_6694);
and U10800 (N_10800,N_8132,N_7497);
nor U10801 (N_10801,N_6468,N_6769);
and U10802 (N_10802,N_8721,N_6253);
or U10803 (N_10803,N_8657,N_6317);
xor U10804 (N_10804,N_6955,N_7828);
or U10805 (N_10805,N_7100,N_6783);
or U10806 (N_10806,N_7694,N_7006);
or U10807 (N_10807,N_8295,N_7342);
xor U10808 (N_10808,N_6881,N_7375);
and U10809 (N_10809,N_6355,N_6455);
xnor U10810 (N_10810,N_8931,N_8580);
or U10811 (N_10811,N_6832,N_6070);
nor U10812 (N_10812,N_6111,N_7074);
or U10813 (N_10813,N_7179,N_8505);
and U10814 (N_10814,N_7509,N_6963);
nor U10815 (N_10815,N_7956,N_8679);
nor U10816 (N_10816,N_6923,N_6797);
xnor U10817 (N_10817,N_8690,N_8815);
xnor U10818 (N_10818,N_6522,N_6977);
nand U10819 (N_10819,N_6537,N_6265);
nand U10820 (N_10820,N_8651,N_6474);
xor U10821 (N_10821,N_8364,N_8265);
or U10822 (N_10822,N_6192,N_7941);
nand U10823 (N_10823,N_8642,N_8796);
xnor U10824 (N_10824,N_8295,N_7642);
nand U10825 (N_10825,N_8372,N_7595);
and U10826 (N_10826,N_8186,N_8965);
nand U10827 (N_10827,N_6104,N_7075);
and U10828 (N_10828,N_7428,N_6132);
nor U10829 (N_10829,N_6479,N_8522);
and U10830 (N_10830,N_6505,N_7655);
nor U10831 (N_10831,N_8221,N_7708);
nor U10832 (N_10832,N_7628,N_6878);
and U10833 (N_10833,N_7316,N_6167);
or U10834 (N_10834,N_6541,N_7785);
or U10835 (N_10835,N_8195,N_8893);
or U10836 (N_10836,N_6866,N_6189);
and U10837 (N_10837,N_7010,N_8283);
and U10838 (N_10838,N_8925,N_7357);
and U10839 (N_10839,N_6511,N_6972);
and U10840 (N_10840,N_8705,N_8219);
and U10841 (N_10841,N_8795,N_7716);
xor U10842 (N_10842,N_7972,N_8109);
or U10843 (N_10843,N_8534,N_6685);
nand U10844 (N_10844,N_6044,N_6096);
nor U10845 (N_10845,N_8445,N_8950);
and U10846 (N_10846,N_6361,N_6830);
nand U10847 (N_10847,N_7756,N_8762);
xnor U10848 (N_10848,N_7805,N_7002);
or U10849 (N_10849,N_6695,N_6787);
xnor U10850 (N_10850,N_8029,N_6790);
xnor U10851 (N_10851,N_6354,N_7236);
nand U10852 (N_10852,N_8716,N_6367);
and U10853 (N_10853,N_7997,N_6283);
and U10854 (N_10854,N_7456,N_7391);
nor U10855 (N_10855,N_7935,N_8178);
and U10856 (N_10856,N_6418,N_7262);
nand U10857 (N_10857,N_7157,N_7713);
xor U10858 (N_10858,N_7016,N_6858);
xor U10859 (N_10859,N_7975,N_7120);
and U10860 (N_10860,N_7781,N_6374);
nor U10861 (N_10861,N_6218,N_6183);
xnor U10862 (N_10862,N_6700,N_8600);
nand U10863 (N_10863,N_6496,N_7101);
nor U10864 (N_10864,N_8778,N_6759);
nand U10865 (N_10865,N_6328,N_8209);
or U10866 (N_10866,N_6326,N_7797);
xnor U10867 (N_10867,N_6283,N_7674);
and U10868 (N_10868,N_8887,N_7729);
and U10869 (N_10869,N_7936,N_6993);
nand U10870 (N_10870,N_6367,N_6954);
or U10871 (N_10871,N_6885,N_6558);
xnor U10872 (N_10872,N_7162,N_8475);
nor U10873 (N_10873,N_7039,N_8728);
nor U10874 (N_10874,N_8977,N_8472);
nor U10875 (N_10875,N_6100,N_8538);
nor U10876 (N_10876,N_6468,N_8240);
nand U10877 (N_10877,N_7448,N_6849);
and U10878 (N_10878,N_8003,N_8516);
nor U10879 (N_10879,N_8351,N_8671);
xor U10880 (N_10880,N_8909,N_8728);
nand U10881 (N_10881,N_8166,N_8886);
nand U10882 (N_10882,N_6103,N_6847);
or U10883 (N_10883,N_7433,N_7817);
nand U10884 (N_10884,N_6506,N_8164);
xnor U10885 (N_10885,N_7436,N_7402);
nand U10886 (N_10886,N_8960,N_6508);
nand U10887 (N_10887,N_7360,N_8493);
nor U10888 (N_10888,N_6261,N_7917);
xnor U10889 (N_10889,N_8037,N_8406);
or U10890 (N_10890,N_8912,N_6618);
or U10891 (N_10891,N_7476,N_6886);
or U10892 (N_10892,N_7814,N_8981);
xor U10893 (N_10893,N_7169,N_8718);
nand U10894 (N_10894,N_8021,N_7203);
or U10895 (N_10895,N_6880,N_7264);
nor U10896 (N_10896,N_7115,N_8034);
nor U10897 (N_10897,N_6245,N_6819);
nor U10898 (N_10898,N_6120,N_8690);
nor U10899 (N_10899,N_8846,N_6523);
or U10900 (N_10900,N_7390,N_7901);
xor U10901 (N_10901,N_8502,N_8204);
and U10902 (N_10902,N_8355,N_7509);
nand U10903 (N_10903,N_7135,N_6715);
nor U10904 (N_10904,N_7506,N_7117);
or U10905 (N_10905,N_8296,N_6898);
or U10906 (N_10906,N_7633,N_8451);
or U10907 (N_10907,N_6963,N_6234);
nor U10908 (N_10908,N_8845,N_7950);
nand U10909 (N_10909,N_8398,N_6676);
nor U10910 (N_10910,N_7393,N_7032);
nor U10911 (N_10911,N_8507,N_8190);
xor U10912 (N_10912,N_7225,N_6398);
nor U10913 (N_10913,N_8201,N_8895);
and U10914 (N_10914,N_6751,N_8895);
nand U10915 (N_10915,N_8733,N_7508);
nand U10916 (N_10916,N_6639,N_6664);
nand U10917 (N_10917,N_7970,N_6601);
xnor U10918 (N_10918,N_7221,N_7648);
nor U10919 (N_10919,N_6204,N_7277);
xor U10920 (N_10920,N_7873,N_7284);
or U10921 (N_10921,N_8358,N_7903);
or U10922 (N_10922,N_8498,N_7248);
and U10923 (N_10923,N_8742,N_7397);
or U10924 (N_10924,N_7274,N_6873);
nand U10925 (N_10925,N_8389,N_8336);
or U10926 (N_10926,N_6226,N_8137);
and U10927 (N_10927,N_6434,N_6176);
nand U10928 (N_10928,N_7235,N_8296);
and U10929 (N_10929,N_6702,N_7318);
or U10930 (N_10930,N_7509,N_6585);
nor U10931 (N_10931,N_8665,N_6104);
nor U10932 (N_10932,N_7618,N_8613);
and U10933 (N_10933,N_8914,N_8995);
nand U10934 (N_10934,N_8166,N_8067);
and U10935 (N_10935,N_6390,N_7757);
nor U10936 (N_10936,N_8352,N_6375);
xor U10937 (N_10937,N_7980,N_8743);
xnor U10938 (N_10938,N_7701,N_8146);
nor U10939 (N_10939,N_6192,N_6432);
or U10940 (N_10940,N_8033,N_7353);
xor U10941 (N_10941,N_7795,N_7484);
or U10942 (N_10942,N_6904,N_8490);
xnor U10943 (N_10943,N_7722,N_8978);
nor U10944 (N_10944,N_6489,N_8974);
nand U10945 (N_10945,N_6956,N_6991);
xnor U10946 (N_10946,N_7486,N_7735);
nor U10947 (N_10947,N_7588,N_8248);
and U10948 (N_10948,N_6579,N_8324);
nand U10949 (N_10949,N_7568,N_8637);
nand U10950 (N_10950,N_8323,N_8857);
xnor U10951 (N_10951,N_6443,N_6558);
or U10952 (N_10952,N_7218,N_8763);
and U10953 (N_10953,N_8755,N_6020);
and U10954 (N_10954,N_7986,N_6458);
nand U10955 (N_10955,N_6731,N_8645);
or U10956 (N_10956,N_6375,N_7270);
or U10957 (N_10957,N_6740,N_8569);
nor U10958 (N_10958,N_8325,N_6772);
or U10959 (N_10959,N_7179,N_6540);
or U10960 (N_10960,N_6143,N_8831);
nor U10961 (N_10961,N_7334,N_7645);
xnor U10962 (N_10962,N_8171,N_6369);
nand U10963 (N_10963,N_7789,N_6156);
nor U10964 (N_10964,N_8577,N_7644);
or U10965 (N_10965,N_7667,N_7702);
xnor U10966 (N_10966,N_6778,N_6741);
nor U10967 (N_10967,N_8206,N_6465);
and U10968 (N_10968,N_6268,N_8829);
xnor U10969 (N_10969,N_6833,N_7979);
nand U10970 (N_10970,N_6061,N_6625);
or U10971 (N_10971,N_8901,N_8595);
or U10972 (N_10972,N_8360,N_6064);
nor U10973 (N_10973,N_8581,N_8359);
nor U10974 (N_10974,N_6750,N_8153);
nand U10975 (N_10975,N_8648,N_8816);
xor U10976 (N_10976,N_6319,N_7214);
nor U10977 (N_10977,N_8751,N_8103);
nand U10978 (N_10978,N_7799,N_6120);
nand U10979 (N_10979,N_6116,N_8844);
and U10980 (N_10980,N_6962,N_8358);
or U10981 (N_10981,N_8348,N_8839);
xor U10982 (N_10982,N_7307,N_8274);
or U10983 (N_10983,N_6859,N_7826);
and U10984 (N_10984,N_8660,N_7811);
and U10985 (N_10985,N_8783,N_6866);
xor U10986 (N_10986,N_6599,N_8126);
or U10987 (N_10987,N_6083,N_6354);
and U10988 (N_10988,N_8079,N_6464);
or U10989 (N_10989,N_6114,N_7642);
nand U10990 (N_10990,N_8219,N_6296);
nor U10991 (N_10991,N_8671,N_7835);
nand U10992 (N_10992,N_8444,N_7621);
nand U10993 (N_10993,N_6509,N_8592);
and U10994 (N_10994,N_8670,N_7407);
nor U10995 (N_10995,N_7344,N_7594);
and U10996 (N_10996,N_8698,N_8526);
or U10997 (N_10997,N_6260,N_6500);
or U10998 (N_10998,N_6082,N_8310);
xor U10999 (N_10999,N_8835,N_6943);
nor U11000 (N_11000,N_7927,N_6797);
and U11001 (N_11001,N_7269,N_7288);
xor U11002 (N_11002,N_7145,N_6307);
nor U11003 (N_11003,N_8668,N_8357);
nor U11004 (N_11004,N_6356,N_6740);
nor U11005 (N_11005,N_8706,N_6868);
and U11006 (N_11006,N_6559,N_7081);
nor U11007 (N_11007,N_8500,N_6122);
xor U11008 (N_11008,N_6987,N_8170);
nor U11009 (N_11009,N_7542,N_6042);
nor U11010 (N_11010,N_8755,N_7762);
or U11011 (N_11011,N_7595,N_7126);
nor U11012 (N_11012,N_7783,N_7138);
nand U11013 (N_11013,N_6742,N_7868);
nand U11014 (N_11014,N_8621,N_8622);
nand U11015 (N_11015,N_6357,N_6599);
and U11016 (N_11016,N_6057,N_6058);
xnor U11017 (N_11017,N_6040,N_6696);
or U11018 (N_11018,N_8303,N_7377);
xor U11019 (N_11019,N_7904,N_6665);
and U11020 (N_11020,N_7159,N_6628);
xor U11021 (N_11021,N_7127,N_7286);
xnor U11022 (N_11022,N_6073,N_8628);
nand U11023 (N_11023,N_8466,N_7384);
nand U11024 (N_11024,N_8230,N_7904);
xnor U11025 (N_11025,N_7925,N_7834);
nor U11026 (N_11026,N_6431,N_7213);
nand U11027 (N_11027,N_6166,N_6887);
nand U11028 (N_11028,N_7483,N_6484);
nand U11029 (N_11029,N_6533,N_7021);
nor U11030 (N_11030,N_8208,N_7611);
nor U11031 (N_11031,N_7522,N_8400);
nand U11032 (N_11032,N_7575,N_8898);
xor U11033 (N_11033,N_7443,N_6280);
xnor U11034 (N_11034,N_6321,N_7319);
nor U11035 (N_11035,N_6326,N_7997);
nor U11036 (N_11036,N_6576,N_7113);
nand U11037 (N_11037,N_7749,N_8881);
xnor U11038 (N_11038,N_6964,N_6006);
and U11039 (N_11039,N_6784,N_7175);
xor U11040 (N_11040,N_6354,N_8180);
or U11041 (N_11041,N_8913,N_8914);
nand U11042 (N_11042,N_7237,N_7967);
nand U11043 (N_11043,N_7537,N_7038);
nor U11044 (N_11044,N_8399,N_8929);
and U11045 (N_11045,N_8688,N_8929);
and U11046 (N_11046,N_7619,N_8028);
or U11047 (N_11047,N_8057,N_8810);
nor U11048 (N_11048,N_7494,N_6434);
xor U11049 (N_11049,N_6651,N_8168);
and U11050 (N_11050,N_6389,N_8771);
xnor U11051 (N_11051,N_6557,N_6451);
or U11052 (N_11052,N_7746,N_8497);
and U11053 (N_11053,N_8726,N_7019);
and U11054 (N_11054,N_6131,N_8033);
xnor U11055 (N_11055,N_7941,N_7024);
nor U11056 (N_11056,N_7648,N_7880);
xnor U11057 (N_11057,N_6717,N_6339);
or U11058 (N_11058,N_6301,N_6198);
xnor U11059 (N_11059,N_7049,N_6738);
xor U11060 (N_11060,N_6834,N_6663);
nand U11061 (N_11061,N_8683,N_6255);
nand U11062 (N_11062,N_8253,N_8659);
or U11063 (N_11063,N_6226,N_7296);
nor U11064 (N_11064,N_8606,N_7185);
and U11065 (N_11065,N_7602,N_6701);
or U11066 (N_11066,N_7533,N_8119);
xor U11067 (N_11067,N_8712,N_6135);
nand U11068 (N_11068,N_8061,N_7814);
nand U11069 (N_11069,N_7018,N_6907);
nor U11070 (N_11070,N_7538,N_7707);
and U11071 (N_11071,N_7184,N_7150);
nor U11072 (N_11072,N_7827,N_6755);
xnor U11073 (N_11073,N_6778,N_6234);
nor U11074 (N_11074,N_6189,N_7132);
and U11075 (N_11075,N_7195,N_7247);
xnor U11076 (N_11076,N_7168,N_8226);
nor U11077 (N_11077,N_7334,N_7045);
or U11078 (N_11078,N_6128,N_6623);
nand U11079 (N_11079,N_6439,N_7532);
xor U11080 (N_11080,N_8872,N_7461);
and U11081 (N_11081,N_6026,N_8962);
xnor U11082 (N_11082,N_7713,N_6954);
and U11083 (N_11083,N_6626,N_6301);
nor U11084 (N_11084,N_7446,N_6965);
nand U11085 (N_11085,N_6344,N_8319);
and U11086 (N_11086,N_7525,N_7791);
xor U11087 (N_11087,N_7579,N_8217);
nand U11088 (N_11088,N_7463,N_7450);
nand U11089 (N_11089,N_6089,N_6641);
nor U11090 (N_11090,N_6900,N_6967);
nor U11091 (N_11091,N_7700,N_7452);
xnor U11092 (N_11092,N_8708,N_8154);
xor U11093 (N_11093,N_8350,N_6518);
nor U11094 (N_11094,N_6645,N_8106);
or U11095 (N_11095,N_6714,N_7608);
nand U11096 (N_11096,N_6784,N_8166);
nand U11097 (N_11097,N_7332,N_7759);
and U11098 (N_11098,N_6959,N_7047);
and U11099 (N_11099,N_7855,N_6808);
and U11100 (N_11100,N_7947,N_7367);
nand U11101 (N_11101,N_8722,N_7857);
nor U11102 (N_11102,N_8568,N_7030);
and U11103 (N_11103,N_7431,N_6568);
or U11104 (N_11104,N_7849,N_6040);
xnor U11105 (N_11105,N_6587,N_7527);
nand U11106 (N_11106,N_6994,N_8152);
nand U11107 (N_11107,N_6460,N_6457);
xor U11108 (N_11108,N_8552,N_6326);
nor U11109 (N_11109,N_8384,N_8770);
nand U11110 (N_11110,N_6041,N_6252);
nand U11111 (N_11111,N_6408,N_6740);
and U11112 (N_11112,N_8288,N_6153);
nor U11113 (N_11113,N_7723,N_8963);
and U11114 (N_11114,N_6802,N_6704);
or U11115 (N_11115,N_8056,N_7985);
nand U11116 (N_11116,N_7943,N_7793);
and U11117 (N_11117,N_6573,N_7111);
xnor U11118 (N_11118,N_7039,N_8993);
xnor U11119 (N_11119,N_8783,N_8700);
xnor U11120 (N_11120,N_7683,N_6155);
or U11121 (N_11121,N_6686,N_8503);
xnor U11122 (N_11122,N_7673,N_7232);
and U11123 (N_11123,N_6719,N_8546);
or U11124 (N_11124,N_8071,N_7814);
nor U11125 (N_11125,N_8739,N_8700);
xnor U11126 (N_11126,N_6673,N_6403);
xor U11127 (N_11127,N_6786,N_6975);
or U11128 (N_11128,N_7106,N_7563);
or U11129 (N_11129,N_7789,N_6925);
and U11130 (N_11130,N_8735,N_8568);
and U11131 (N_11131,N_7362,N_7828);
nand U11132 (N_11132,N_8353,N_7051);
xor U11133 (N_11133,N_6329,N_8398);
or U11134 (N_11134,N_6217,N_7231);
xor U11135 (N_11135,N_6868,N_6617);
and U11136 (N_11136,N_8018,N_6806);
xnor U11137 (N_11137,N_8437,N_8042);
nor U11138 (N_11138,N_6144,N_7097);
or U11139 (N_11139,N_8563,N_8183);
and U11140 (N_11140,N_6831,N_6696);
nand U11141 (N_11141,N_6858,N_7254);
xnor U11142 (N_11142,N_6093,N_7473);
and U11143 (N_11143,N_6694,N_8929);
nand U11144 (N_11144,N_8708,N_6102);
or U11145 (N_11145,N_6154,N_7074);
and U11146 (N_11146,N_8300,N_7416);
nand U11147 (N_11147,N_7292,N_7871);
or U11148 (N_11148,N_7094,N_8864);
or U11149 (N_11149,N_7919,N_8897);
and U11150 (N_11150,N_6904,N_8309);
xor U11151 (N_11151,N_6207,N_6010);
nor U11152 (N_11152,N_8256,N_8393);
nand U11153 (N_11153,N_7214,N_6803);
and U11154 (N_11154,N_7653,N_8522);
xnor U11155 (N_11155,N_7662,N_8793);
or U11156 (N_11156,N_7396,N_8125);
xnor U11157 (N_11157,N_6321,N_8303);
and U11158 (N_11158,N_6551,N_8425);
and U11159 (N_11159,N_8959,N_7399);
nor U11160 (N_11160,N_7981,N_6583);
xor U11161 (N_11161,N_6753,N_7841);
and U11162 (N_11162,N_6765,N_6805);
and U11163 (N_11163,N_6086,N_8629);
and U11164 (N_11164,N_6300,N_8105);
and U11165 (N_11165,N_7457,N_6191);
xor U11166 (N_11166,N_7423,N_6729);
nand U11167 (N_11167,N_8997,N_7375);
and U11168 (N_11168,N_6801,N_8354);
nor U11169 (N_11169,N_8717,N_8748);
nand U11170 (N_11170,N_7308,N_6075);
nor U11171 (N_11171,N_6237,N_6186);
or U11172 (N_11172,N_6161,N_7182);
nand U11173 (N_11173,N_8221,N_8477);
nor U11174 (N_11174,N_8515,N_6007);
nor U11175 (N_11175,N_8047,N_7843);
nor U11176 (N_11176,N_8571,N_7088);
xnor U11177 (N_11177,N_7183,N_8494);
nand U11178 (N_11178,N_6613,N_6456);
nor U11179 (N_11179,N_7714,N_7031);
nor U11180 (N_11180,N_8181,N_7853);
or U11181 (N_11181,N_7984,N_7691);
xor U11182 (N_11182,N_6346,N_8399);
and U11183 (N_11183,N_8176,N_7523);
or U11184 (N_11184,N_8232,N_8821);
or U11185 (N_11185,N_7206,N_6520);
and U11186 (N_11186,N_8885,N_7334);
or U11187 (N_11187,N_8353,N_6324);
xor U11188 (N_11188,N_7244,N_7510);
or U11189 (N_11189,N_8676,N_7885);
or U11190 (N_11190,N_7897,N_8890);
nor U11191 (N_11191,N_7713,N_6152);
nor U11192 (N_11192,N_7656,N_6540);
and U11193 (N_11193,N_6507,N_7908);
and U11194 (N_11194,N_6339,N_7029);
nor U11195 (N_11195,N_8988,N_6379);
nor U11196 (N_11196,N_7208,N_7359);
and U11197 (N_11197,N_8972,N_6648);
nor U11198 (N_11198,N_8086,N_7394);
or U11199 (N_11199,N_7997,N_7550);
xnor U11200 (N_11200,N_7346,N_6751);
nand U11201 (N_11201,N_8378,N_8746);
xor U11202 (N_11202,N_6255,N_8305);
and U11203 (N_11203,N_6693,N_7601);
nand U11204 (N_11204,N_6052,N_8381);
or U11205 (N_11205,N_7352,N_8114);
xor U11206 (N_11206,N_6297,N_8161);
nand U11207 (N_11207,N_6190,N_7963);
or U11208 (N_11208,N_7377,N_8453);
and U11209 (N_11209,N_8803,N_6909);
or U11210 (N_11210,N_6430,N_7710);
or U11211 (N_11211,N_6578,N_8756);
xor U11212 (N_11212,N_6345,N_7848);
xnor U11213 (N_11213,N_6702,N_8341);
nand U11214 (N_11214,N_8449,N_6575);
and U11215 (N_11215,N_7125,N_6912);
and U11216 (N_11216,N_6467,N_8289);
and U11217 (N_11217,N_7396,N_6974);
and U11218 (N_11218,N_6263,N_7154);
or U11219 (N_11219,N_6165,N_8749);
nand U11220 (N_11220,N_7380,N_7017);
or U11221 (N_11221,N_7953,N_6708);
nor U11222 (N_11222,N_7380,N_7614);
nand U11223 (N_11223,N_8466,N_7675);
nor U11224 (N_11224,N_7130,N_8320);
nor U11225 (N_11225,N_6793,N_6370);
xor U11226 (N_11226,N_6677,N_6989);
and U11227 (N_11227,N_7788,N_7157);
xnor U11228 (N_11228,N_8474,N_7838);
nor U11229 (N_11229,N_6817,N_8533);
or U11230 (N_11230,N_8660,N_7929);
nand U11231 (N_11231,N_6601,N_8099);
nand U11232 (N_11232,N_8062,N_6936);
nor U11233 (N_11233,N_7456,N_6726);
and U11234 (N_11234,N_6385,N_6787);
xor U11235 (N_11235,N_6053,N_6757);
and U11236 (N_11236,N_8380,N_6527);
xor U11237 (N_11237,N_8479,N_6865);
xnor U11238 (N_11238,N_7937,N_7359);
nand U11239 (N_11239,N_6573,N_6162);
xor U11240 (N_11240,N_8819,N_6698);
nand U11241 (N_11241,N_8433,N_6824);
nand U11242 (N_11242,N_6431,N_8591);
xnor U11243 (N_11243,N_8864,N_7965);
nor U11244 (N_11244,N_7535,N_7530);
nand U11245 (N_11245,N_7452,N_8601);
or U11246 (N_11246,N_7305,N_8254);
nor U11247 (N_11247,N_7476,N_6460);
nor U11248 (N_11248,N_8753,N_7213);
nand U11249 (N_11249,N_7291,N_6746);
and U11250 (N_11250,N_6019,N_7052);
or U11251 (N_11251,N_7892,N_6854);
xnor U11252 (N_11252,N_7893,N_7419);
nand U11253 (N_11253,N_8995,N_7299);
xor U11254 (N_11254,N_6728,N_8371);
xnor U11255 (N_11255,N_7384,N_6460);
nand U11256 (N_11256,N_6205,N_8735);
xnor U11257 (N_11257,N_6696,N_8716);
nand U11258 (N_11258,N_6710,N_6821);
or U11259 (N_11259,N_8445,N_7703);
or U11260 (N_11260,N_8678,N_7293);
nor U11261 (N_11261,N_6069,N_8908);
nand U11262 (N_11262,N_7953,N_7271);
nor U11263 (N_11263,N_7388,N_7414);
nor U11264 (N_11264,N_7329,N_7799);
or U11265 (N_11265,N_6348,N_7941);
and U11266 (N_11266,N_6432,N_7537);
nand U11267 (N_11267,N_6871,N_6612);
nand U11268 (N_11268,N_7035,N_6171);
nor U11269 (N_11269,N_8785,N_7687);
nor U11270 (N_11270,N_7161,N_6230);
and U11271 (N_11271,N_7423,N_7943);
nor U11272 (N_11272,N_6521,N_7166);
and U11273 (N_11273,N_6838,N_8339);
or U11274 (N_11274,N_6412,N_6031);
or U11275 (N_11275,N_8220,N_7620);
or U11276 (N_11276,N_8829,N_8370);
or U11277 (N_11277,N_8020,N_7880);
nand U11278 (N_11278,N_8335,N_6294);
nor U11279 (N_11279,N_8666,N_7748);
nand U11280 (N_11280,N_7524,N_8184);
or U11281 (N_11281,N_6900,N_8102);
nor U11282 (N_11282,N_7359,N_6243);
nand U11283 (N_11283,N_6089,N_8020);
nor U11284 (N_11284,N_8584,N_7001);
nand U11285 (N_11285,N_8865,N_7878);
and U11286 (N_11286,N_6816,N_8127);
xnor U11287 (N_11287,N_7258,N_6786);
or U11288 (N_11288,N_6182,N_8850);
and U11289 (N_11289,N_7148,N_8150);
nand U11290 (N_11290,N_6029,N_8837);
nor U11291 (N_11291,N_7009,N_8354);
and U11292 (N_11292,N_6029,N_6026);
nor U11293 (N_11293,N_6409,N_8914);
nor U11294 (N_11294,N_7499,N_6251);
nand U11295 (N_11295,N_7692,N_6315);
nor U11296 (N_11296,N_7393,N_6345);
and U11297 (N_11297,N_6194,N_6610);
and U11298 (N_11298,N_8621,N_6461);
or U11299 (N_11299,N_8579,N_6436);
xor U11300 (N_11300,N_8926,N_8128);
xnor U11301 (N_11301,N_8891,N_8825);
xnor U11302 (N_11302,N_6750,N_8592);
xnor U11303 (N_11303,N_8694,N_7668);
or U11304 (N_11304,N_7015,N_8928);
and U11305 (N_11305,N_8944,N_7423);
and U11306 (N_11306,N_6281,N_6792);
nand U11307 (N_11307,N_8025,N_6548);
and U11308 (N_11308,N_8131,N_8271);
or U11309 (N_11309,N_7968,N_7264);
or U11310 (N_11310,N_6898,N_6772);
xnor U11311 (N_11311,N_6221,N_7341);
xnor U11312 (N_11312,N_6335,N_7901);
xor U11313 (N_11313,N_6313,N_7000);
nor U11314 (N_11314,N_6145,N_6311);
or U11315 (N_11315,N_8401,N_8153);
xnor U11316 (N_11316,N_6385,N_7465);
nor U11317 (N_11317,N_6868,N_7929);
nand U11318 (N_11318,N_7355,N_6007);
nand U11319 (N_11319,N_7597,N_8062);
nand U11320 (N_11320,N_8358,N_7414);
nor U11321 (N_11321,N_7956,N_7299);
xnor U11322 (N_11322,N_6947,N_7710);
or U11323 (N_11323,N_6343,N_6958);
or U11324 (N_11324,N_6193,N_6841);
or U11325 (N_11325,N_8572,N_8413);
nor U11326 (N_11326,N_6948,N_7115);
or U11327 (N_11327,N_6329,N_7160);
or U11328 (N_11328,N_6635,N_8638);
nor U11329 (N_11329,N_6413,N_8935);
and U11330 (N_11330,N_7791,N_6660);
xor U11331 (N_11331,N_8090,N_7449);
or U11332 (N_11332,N_6183,N_8163);
and U11333 (N_11333,N_8680,N_8237);
or U11334 (N_11334,N_6201,N_7901);
nand U11335 (N_11335,N_6858,N_7256);
or U11336 (N_11336,N_6004,N_7380);
and U11337 (N_11337,N_8169,N_6136);
nor U11338 (N_11338,N_7597,N_6292);
or U11339 (N_11339,N_7212,N_7816);
nand U11340 (N_11340,N_7561,N_8075);
xnor U11341 (N_11341,N_7633,N_7394);
nor U11342 (N_11342,N_6156,N_6071);
or U11343 (N_11343,N_7970,N_8423);
and U11344 (N_11344,N_8791,N_7234);
nor U11345 (N_11345,N_7467,N_8543);
or U11346 (N_11346,N_8938,N_6074);
nand U11347 (N_11347,N_7509,N_8717);
xnor U11348 (N_11348,N_7986,N_8196);
nand U11349 (N_11349,N_8768,N_7011);
xnor U11350 (N_11350,N_6063,N_8389);
nand U11351 (N_11351,N_7095,N_7098);
nand U11352 (N_11352,N_8835,N_6626);
nand U11353 (N_11353,N_7892,N_6329);
or U11354 (N_11354,N_7718,N_8979);
nand U11355 (N_11355,N_7267,N_6848);
nand U11356 (N_11356,N_6919,N_6060);
and U11357 (N_11357,N_7778,N_6203);
nand U11358 (N_11358,N_6835,N_8621);
xnor U11359 (N_11359,N_7008,N_7789);
nor U11360 (N_11360,N_7845,N_8549);
nand U11361 (N_11361,N_6221,N_8419);
or U11362 (N_11362,N_7119,N_7820);
or U11363 (N_11363,N_7242,N_8216);
and U11364 (N_11364,N_6490,N_8837);
nor U11365 (N_11365,N_7879,N_7487);
and U11366 (N_11366,N_7601,N_7196);
nor U11367 (N_11367,N_8056,N_8799);
xnor U11368 (N_11368,N_8855,N_8934);
or U11369 (N_11369,N_6385,N_6382);
or U11370 (N_11370,N_7957,N_7412);
xor U11371 (N_11371,N_6468,N_6217);
nor U11372 (N_11372,N_7903,N_6437);
nor U11373 (N_11373,N_8751,N_7445);
xor U11374 (N_11374,N_7130,N_8604);
xor U11375 (N_11375,N_7644,N_7187);
xor U11376 (N_11376,N_8697,N_6526);
xnor U11377 (N_11377,N_7209,N_6230);
or U11378 (N_11378,N_6265,N_6425);
or U11379 (N_11379,N_6386,N_8568);
nand U11380 (N_11380,N_7433,N_8368);
nor U11381 (N_11381,N_6632,N_8319);
nand U11382 (N_11382,N_7653,N_8337);
nor U11383 (N_11383,N_7165,N_7852);
nand U11384 (N_11384,N_7982,N_7370);
and U11385 (N_11385,N_6809,N_6683);
or U11386 (N_11386,N_7752,N_6939);
and U11387 (N_11387,N_8547,N_7784);
nor U11388 (N_11388,N_8052,N_7608);
xnor U11389 (N_11389,N_8702,N_8779);
or U11390 (N_11390,N_8322,N_7382);
and U11391 (N_11391,N_6409,N_8669);
or U11392 (N_11392,N_6150,N_8111);
nor U11393 (N_11393,N_6764,N_8349);
or U11394 (N_11394,N_8070,N_8977);
xor U11395 (N_11395,N_8004,N_8407);
xor U11396 (N_11396,N_8689,N_8617);
xor U11397 (N_11397,N_8825,N_8349);
xnor U11398 (N_11398,N_8000,N_6840);
nand U11399 (N_11399,N_8202,N_6994);
nor U11400 (N_11400,N_8251,N_6495);
xnor U11401 (N_11401,N_8101,N_6381);
nand U11402 (N_11402,N_8417,N_7338);
and U11403 (N_11403,N_7431,N_8903);
or U11404 (N_11404,N_6881,N_6157);
or U11405 (N_11405,N_8151,N_7472);
or U11406 (N_11406,N_7259,N_7966);
nand U11407 (N_11407,N_7013,N_8403);
xor U11408 (N_11408,N_6840,N_7692);
xnor U11409 (N_11409,N_7664,N_7347);
or U11410 (N_11410,N_8952,N_7075);
and U11411 (N_11411,N_7730,N_7075);
nor U11412 (N_11412,N_6385,N_7165);
or U11413 (N_11413,N_8040,N_6316);
and U11414 (N_11414,N_6218,N_8962);
nor U11415 (N_11415,N_8819,N_8935);
nor U11416 (N_11416,N_7362,N_7518);
or U11417 (N_11417,N_8866,N_6974);
nand U11418 (N_11418,N_6861,N_7404);
or U11419 (N_11419,N_6611,N_6410);
xnor U11420 (N_11420,N_8688,N_6350);
nand U11421 (N_11421,N_7017,N_8792);
and U11422 (N_11422,N_6396,N_8327);
or U11423 (N_11423,N_7848,N_8845);
and U11424 (N_11424,N_6173,N_6829);
nor U11425 (N_11425,N_8542,N_8825);
nor U11426 (N_11426,N_6480,N_8833);
nand U11427 (N_11427,N_8834,N_8665);
or U11428 (N_11428,N_6398,N_8717);
or U11429 (N_11429,N_7308,N_6033);
nor U11430 (N_11430,N_7344,N_8815);
xnor U11431 (N_11431,N_7872,N_6927);
xnor U11432 (N_11432,N_8050,N_6186);
xor U11433 (N_11433,N_7199,N_7347);
nand U11434 (N_11434,N_7164,N_6593);
nor U11435 (N_11435,N_7020,N_8239);
nor U11436 (N_11436,N_7364,N_6906);
or U11437 (N_11437,N_7414,N_8692);
xnor U11438 (N_11438,N_6302,N_8561);
xnor U11439 (N_11439,N_6075,N_6231);
or U11440 (N_11440,N_7105,N_7044);
nand U11441 (N_11441,N_6974,N_8455);
nor U11442 (N_11442,N_8250,N_7375);
nand U11443 (N_11443,N_6940,N_7189);
nor U11444 (N_11444,N_7736,N_8770);
or U11445 (N_11445,N_6716,N_7261);
and U11446 (N_11446,N_7517,N_7093);
xnor U11447 (N_11447,N_8790,N_6484);
and U11448 (N_11448,N_7195,N_8288);
or U11449 (N_11449,N_6618,N_6767);
xnor U11450 (N_11450,N_6893,N_8238);
nor U11451 (N_11451,N_6539,N_7093);
or U11452 (N_11452,N_8796,N_6535);
nor U11453 (N_11453,N_8726,N_6662);
and U11454 (N_11454,N_6003,N_8269);
or U11455 (N_11455,N_8741,N_7317);
and U11456 (N_11456,N_6222,N_8096);
nor U11457 (N_11457,N_8250,N_8445);
nand U11458 (N_11458,N_8412,N_8383);
or U11459 (N_11459,N_7014,N_8921);
xnor U11460 (N_11460,N_8455,N_7588);
nand U11461 (N_11461,N_6694,N_7218);
nor U11462 (N_11462,N_7165,N_7314);
or U11463 (N_11463,N_7367,N_6134);
and U11464 (N_11464,N_6473,N_7431);
nand U11465 (N_11465,N_7442,N_6432);
and U11466 (N_11466,N_8505,N_7873);
and U11467 (N_11467,N_6901,N_6725);
nor U11468 (N_11468,N_7320,N_7561);
nand U11469 (N_11469,N_8397,N_8558);
xor U11470 (N_11470,N_6002,N_7425);
or U11471 (N_11471,N_8492,N_7519);
or U11472 (N_11472,N_8686,N_7802);
nor U11473 (N_11473,N_6466,N_6100);
nand U11474 (N_11474,N_6079,N_6330);
or U11475 (N_11475,N_8602,N_6172);
xnor U11476 (N_11476,N_8695,N_8680);
and U11477 (N_11477,N_6284,N_6854);
nand U11478 (N_11478,N_7577,N_6592);
nand U11479 (N_11479,N_8807,N_8682);
nand U11480 (N_11480,N_8853,N_7051);
nor U11481 (N_11481,N_6092,N_8183);
nor U11482 (N_11482,N_7791,N_8833);
or U11483 (N_11483,N_8488,N_7042);
or U11484 (N_11484,N_7331,N_8338);
nor U11485 (N_11485,N_8175,N_8569);
or U11486 (N_11486,N_7961,N_6013);
xnor U11487 (N_11487,N_7379,N_8366);
or U11488 (N_11488,N_7631,N_6715);
and U11489 (N_11489,N_7898,N_6514);
and U11490 (N_11490,N_6082,N_8953);
and U11491 (N_11491,N_7925,N_6932);
and U11492 (N_11492,N_7819,N_8610);
nor U11493 (N_11493,N_8522,N_8597);
nand U11494 (N_11494,N_6949,N_8549);
xnor U11495 (N_11495,N_8846,N_6972);
nand U11496 (N_11496,N_7152,N_7040);
nor U11497 (N_11497,N_7667,N_8469);
nor U11498 (N_11498,N_7688,N_6218);
and U11499 (N_11499,N_6023,N_7776);
nor U11500 (N_11500,N_6351,N_7006);
nor U11501 (N_11501,N_8319,N_7999);
or U11502 (N_11502,N_8202,N_8723);
xor U11503 (N_11503,N_7419,N_6308);
or U11504 (N_11504,N_6239,N_6955);
xnor U11505 (N_11505,N_7438,N_7656);
or U11506 (N_11506,N_6546,N_7702);
nor U11507 (N_11507,N_6216,N_8568);
or U11508 (N_11508,N_8922,N_7536);
xor U11509 (N_11509,N_7293,N_7590);
or U11510 (N_11510,N_8959,N_6744);
and U11511 (N_11511,N_6885,N_6305);
xnor U11512 (N_11512,N_6772,N_6638);
or U11513 (N_11513,N_6566,N_8469);
or U11514 (N_11514,N_6318,N_7991);
nand U11515 (N_11515,N_7126,N_8965);
nor U11516 (N_11516,N_7124,N_7841);
nand U11517 (N_11517,N_7389,N_6612);
or U11518 (N_11518,N_8356,N_8518);
and U11519 (N_11519,N_6991,N_8768);
xor U11520 (N_11520,N_7682,N_7783);
nor U11521 (N_11521,N_6387,N_6366);
xnor U11522 (N_11522,N_6407,N_7902);
nor U11523 (N_11523,N_7933,N_6629);
nand U11524 (N_11524,N_7698,N_7670);
and U11525 (N_11525,N_8217,N_8861);
or U11526 (N_11526,N_7595,N_7296);
nand U11527 (N_11527,N_6561,N_8863);
or U11528 (N_11528,N_6094,N_8067);
xnor U11529 (N_11529,N_7787,N_6378);
or U11530 (N_11530,N_8473,N_7370);
xnor U11531 (N_11531,N_7348,N_6237);
or U11532 (N_11532,N_7360,N_6664);
xnor U11533 (N_11533,N_8845,N_7737);
and U11534 (N_11534,N_7476,N_8778);
and U11535 (N_11535,N_8108,N_6680);
and U11536 (N_11536,N_7316,N_6229);
and U11537 (N_11537,N_8309,N_8567);
xor U11538 (N_11538,N_8474,N_8361);
or U11539 (N_11539,N_8457,N_7071);
and U11540 (N_11540,N_6475,N_7369);
xnor U11541 (N_11541,N_8082,N_8221);
or U11542 (N_11542,N_8741,N_7417);
or U11543 (N_11543,N_7030,N_6828);
nand U11544 (N_11544,N_6174,N_6202);
nand U11545 (N_11545,N_7568,N_7889);
xor U11546 (N_11546,N_6645,N_7600);
nand U11547 (N_11547,N_6080,N_8196);
nor U11548 (N_11548,N_6973,N_8958);
xnor U11549 (N_11549,N_7574,N_6209);
and U11550 (N_11550,N_8740,N_8134);
and U11551 (N_11551,N_6722,N_7732);
nand U11552 (N_11552,N_8173,N_6690);
xnor U11553 (N_11553,N_8469,N_7476);
nor U11554 (N_11554,N_8269,N_8861);
nand U11555 (N_11555,N_8591,N_8049);
xnor U11556 (N_11556,N_7279,N_8077);
nor U11557 (N_11557,N_7955,N_6292);
nor U11558 (N_11558,N_8397,N_7889);
nand U11559 (N_11559,N_8685,N_6368);
nand U11560 (N_11560,N_6555,N_8055);
or U11561 (N_11561,N_8498,N_7225);
nand U11562 (N_11562,N_7011,N_7068);
nand U11563 (N_11563,N_7604,N_7938);
xnor U11564 (N_11564,N_6150,N_7422);
nand U11565 (N_11565,N_6707,N_7636);
and U11566 (N_11566,N_8758,N_7343);
nand U11567 (N_11567,N_7183,N_8079);
xnor U11568 (N_11568,N_7348,N_7180);
nand U11569 (N_11569,N_8385,N_6128);
nand U11570 (N_11570,N_7241,N_8016);
and U11571 (N_11571,N_6146,N_7058);
and U11572 (N_11572,N_6468,N_7050);
xor U11573 (N_11573,N_7969,N_6994);
or U11574 (N_11574,N_8458,N_8950);
nand U11575 (N_11575,N_8973,N_6292);
xor U11576 (N_11576,N_6293,N_7354);
nor U11577 (N_11577,N_8661,N_7810);
or U11578 (N_11578,N_7145,N_7783);
xor U11579 (N_11579,N_7685,N_6479);
and U11580 (N_11580,N_6963,N_6489);
and U11581 (N_11581,N_8364,N_6910);
and U11582 (N_11582,N_6608,N_7631);
or U11583 (N_11583,N_8279,N_8196);
and U11584 (N_11584,N_7771,N_6249);
xnor U11585 (N_11585,N_7379,N_6087);
and U11586 (N_11586,N_6590,N_6444);
nor U11587 (N_11587,N_8000,N_6224);
and U11588 (N_11588,N_7378,N_8956);
or U11589 (N_11589,N_8955,N_6447);
nor U11590 (N_11590,N_8429,N_6946);
nor U11591 (N_11591,N_6416,N_6479);
and U11592 (N_11592,N_6639,N_7910);
nor U11593 (N_11593,N_7170,N_7435);
xnor U11594 (N_11594,N_7437,N_8317);
nor U11595 (N_11595,N_6925,N_8772);
xor U11596 (N_11596,N_7675,N_7521);
nand U11597 (N_11597,N_8123,N_8085);
nand U11598 (N_11598,N_8088,N_8494);
nand U11599 (N_11599,N_6267,N_8932);
or U11600 (N_11600,N_7912,N_8623);
and U11601 (N_11601,N_7715,N_8869);
nor U11602 (N_11602,N_8179,N_8774);
nand U11603 (N_11603,N_7038,N_8587);
or U11604 (N_11604,N_7249,N_8118);
xnor U11605 (N_11605,N_7295,N_8268);
or U11606 (N_11606,N_7313,N_7525);
and U11607 (N_11607,N_6722,N_6421);
or U11608 (N_11608,N_6095,N_8834);
nand U11609 (N_11609,N_8401,N_7316);
xor U11610 (N_11610,N_7210,N_8072);
and U11611 (N_11611,N_6833,N_8797);
and U11612 (N_11612,N_8966,N_6313);
or U11613 (N_11613,N_7142,N_7419);
and U11614 (N_11614,N_7628,N_7152);
and U11615 (N_11615,N_6896,N_7222);
nand U11616 (N_11616,N_8481,N_6791);
or U11617 (N_11617,N_6554,N_8783);
and U11618 (N_11618,N_8511,N_6713);
or U11619 (N_11619,N_6666,N_8630);
or U11620 (N_11620,N_6647,N_8423);
nand U11621 (N_11621,N_6348,N_8331);
nor U11622 (N_11622,N_7004,N_7116);
and U11623 (N_11623,N_8049,N_8847);
xnor U11624 (N_11624,N_6171,N_6176);
or U11625 (N_11625,N_7364,N_6967);
nor U11626 (N_11626,N_8130,N_8169);
or U11627 (N_11627,N_7050,N_6047);
nor U11628 (N_11628,N_6454,N_7220);
nand U11629 (N_11629,N_8642,N_6259);
nand U11630 (N_11630,N_6840,N_7065);
xor U11631 (N_11631,N_8520,N_8981);
and U11632 (N_11632,N_6707,N_8335);
or U11633 (N_11633,N_8611,N_8390);
nand U11634 (N_11634,N_7210,N_8996);
or U11635 (N_11635,N_6169,N_7902);
and U11636 (N_11636,N_8328,N_7573);
nand U11637 (N_11637,N_6213,N_7771);
nor U11638 (N_11638,N_7287,N_7259);
or U11639 (N_11639,N_6768,N_6935);
or U11640 (N_11640,N_8543,N_7940);
nand U11641 (N_11641,N_7475,N_7569);
nand U11642 (N_11642,N_8512,N_8690);
xor U11643 (N_11643,N_7998,N_7699);
nand U11644 (N_11644,N_8847,N_7751);
or U11645 (N_11645,N_6868,N_8013);
nor U11646 (N_11646,N_8074,N_7540);
nand U11647 (N_11647,N_8107,N_7506);
or U11648 (N_11648,N_7801,N_7053);
nand U11649 (N_11649,N_7825,N_6094);
nor U11650 (N_11650,N_8269,N_7969);
or U11651 (N_11651,N_8540,N_6642);
xor U11652 (N_11652,N_6087,N_7154);
or U11653 (N_11653,N_7762,N_6409);
or U11654 (N_11654,N_6413,N_8549);
xor U11655 (N_11655,N_7651,N_7797);
or U11656 (N_11656,N_7200,N_6357);
or U11657 (N_11657,N_6693,N_7949);
nand U11658 (N_11658,N_7283,N_6582);
and U11659 (N_11659,N_8175,N_7648);
or U11660 (N_11660,N_8831,N_7224);
nand U11661 (N_11661,N_6265,N_6988);
nor U11662 (N_11662,N_7375,N_7698);
nor U11663 (N_11663,N_8885,N_8461);
xor U11664 (N_11664,N_7171,N_6425);
xor U11665 (N_11665,N_6849,N_6764);
nand U11666 (N_11666,N_6393,N_6080);
or U11667 (N_11667,N_7120,N_6586);
nand U11668 (N_11668,N_7329,N_7439);
nand U11669 (N_11669,N_6774,N_7124);
nor U11670 (N_11670,N_8159,N_8769);
nand U11671 (N_11671,N_6845,N_7792);
nor U11672 (N_11672,N_7680,N_6735);
nand U11673 (N_11673,N_8064,N_8755);
nor U11674 (N_11674,N_8232,N_6652);
and U11675 (N_11675,N_7007,N_6190);
and U11676 (N_11676,N_8653,N_7546);
or U11677 (N_11677,N_6746,N_8096);
xor U11678 (N_11678,N_6765,N_6210);
nor U11679 (N_11679,N_8082,N_6819);
nor U11680 (N_11680,N_8165,N_8171);
and U11681 (N_11681,N_8728,N_8480);
xor U11682 (N_11682,N_8787,N_6351);
nand U11683 (N_11683,N_6576,N_8545);
or U11684 (N_11684,N_6744,N_8635);
nor U11685 (N_11685,N_6145,N_6189);
xor U11686 (N_11686,N_8318,N_8901);
nand U11687 (N_11687,N_8992,N_8938);
nand U11688 (N_11688,N_8528,N_8278);
nor U11689 (N_11689,N_8803,N_8206);
nor U11690 (N_11690,N_8301,N_7729);
or U11691 (N_11691,N_6360,N_6643);
or U11692 (N_11692,N_7446,N_8783);
nand U11693 (N_11693,N_8177,N_7120);
xor U11694 (N_11694,N_6166,N_6304);
or U11695 (N_11695,N_7801,N_6341);
and U11696 (N_11696,N_7018,N_8219);
xnor U11697 (N_11697,N_7344,N_8991);
xor U11698 (N_11698,N_7031,N_8882);
and U11699 (N_11699,N_8822,N_8867);
nand U11700 (N_11700,N_6499,N_8816);
and U11701 (N_11701,N_6542,N_7168);
nor U11702 (N_11702,N_8996,N_8086);
nand U11703 (N_11703,N_6398,N_7587);
nor U11704 (N_11704,N_7674,N_7028);
and U11705 (N_11705,N_6659,N_6650);
nand U11706 (N_11706,N_6140,N_6582);
nand U11707 (N_11707,N_8753,N_8566);
and U11708 (N_11708,N_7409,N_6083);
or U11709 (N_11709,N_7041,N_7706);
or U11710 (N_11710,N_6670,N_8245);
nor U11711 (N_11711,N_6182,N_8127);
xnor U11712 (N_11712,N_6554,N_8905);
or U11713 (N_11713,N_8862,N_8393);
nand U11714 (N_11714,N_7057,N_7874);
or U11715 (N_11715,N_7627,N_7879);
or U11716 (N_11716,N_8182,N_7383);
xor U11717 (N_11717,N_7217,N_7882);
xor U11718 (N_11718,N_7662,N_6134);
xnor U11719 (N_11719,N_8537,N_6688);
nand U11720 (N_11720,N_7496,N_6194);
nor U11721 (N_11721,N_6529,N_6353);
and U11722 (N_11722,N_8098,N_6639);
xnor U11723 (N_11723,N_7573,N_6516);
or U11724 (N_11724,N_8112,N_8476);
nand U11725 (N_11725,N_6900,N_8011);
xor U11726 (N_11726,N_8779,N_6146);
nand U11727 (N_11727,N_6528,N_7984);
xor U11728 (N_11728,N_6991,N_6112);
nand U11729 (N_11729,N_6635,N_8384);
nor U11730 (N_11730,N_6793,N_7425);
or U11731 (N_11731,N_6118,N_7905);
xnor U11732 (N_11732,N_6511,N_6734);
and U11733 (N_11733,N_8970,N_8132);
or U11734 (N_11734,N_8276,N_8305);
and U11735 (N_11735,N_8436,N_7050);
xnor U11736 (N_11736,N_8450,N_8343);
xor U11737 (N_11737,N_6313,N_8911);
and U11738 (N_11738,N_6281,N_8209);
nand U11739 (N_11739,N_6582,N_7583);
nor U11740 (N_11740,N_7619,N_7768);
or U11741 (N_11741,N_7002,N_6873);
and U11742 (N_11742,N_6884,N_8059);
nand U11743 (N_11743,N_6242,N_8003);
nand U11744 (N_11744,N_7432,N_6624);
nor U11745 (N_11745,N_7877,N_7393);
or U11746 (N_11746,N_6802,N_6184);
nor U11747 (N_11747,N_6080,N_6985);
xnor U11748 (N_11748,N_8735,N_7581);
xor U11749 (N_11749,N_8114,N_6752);
nor U11750 (N_11750,N_6795,N_8942);
and U11751 (N_11751,N_6465,N_6178);
xnor U11752 (N_11752,N_8855,N_7799);
and U11753 (N_11753,N_6445,N_7976);
nor U11754 (N_11754,N_8867,N_7536);
and U11755 (N_11755,N_7953,N_6412);
and U11756 (N_11756,N_6220,N_7323);
nor U11757 (N_11757,N_6096,N_8853);
nand U11758 (N_11758,N_6363,N_8292);
xnor U11759 (N_11759,N_7513,N_7119);
or U11760 (N_11760,N_6483,N_8758);
xnor U11761 (N_11761,N_6426,N_7936);
or U11762 (N_11762,N_6528,N_7775);
or U11763 (N_11763,N_8029,N_7103);
nand U11764 (N_11764,N_6858,N_7967);
nand U11765 (N_11765,N_7150,N_8104);
and U11766 (N_11766,N_7156,N_7936);
nand U11767 (N_11767,N_7249,N_7589);
nor U11768 (N_11768,N_7853,N_8259);
nand U11769 (N_11769,N_6215,N_8633);
nor U11770 (N_11770,N_8888,N_8266);
and U11771 (N_11771,N_7819,N_8118);
xnor U11772 (N_11772,N_7672,N_7604);
nand U11773 (N_11773,N_8904,N_8710);
and U11774 (N_11774,N_7076,N_8954);
xor U11775 (N_11775,N_7647,N_6322);
nand U11776 (N_11776,N_8650,N_8744);
xor U11777 (N_11777,N_7659,N_8835);
or U11778 (N_11778,N_6577,N_7591);
and U11779 (N_11779,N_8197,N_7276);
xor U11780 (N_11780,N_8294,N_8832);
and U11781 (N_11781,N_6915,N_8192);
nand U11782 (N_11782,N_7053,N_7741);
nand U11783 (N_11783,N_7450,N_7186);
or U11784 (N_11784,N_8276,N_8581);
xor U11785 (N_11785,N_6171,N_8315);
nand U11786 (N_11786,N_8958,N_8741);
nor U11787 (N_11787,N_6534,N_7051);
xor U11788 (N_11788,N_6626,N_8328);
nor U11789 (N_11789,N_6134,N_8009);
and U11790 (N_11790,N_6107,N_6645);
xnor U11791 (N_11791,N_7283,N_6904);
nand U11792 (N_11792,N_7502,N_6150);
or U11793 (N_11793,N_7496,N_6479);
or U11794 (N_11794,N_8800,N_6392);
nor U11795 (N_11795,N_7413,N_7753);
xnor U11796 (N_11796,N_6636,N_6823);
or U11797 (N_11797,N_6024,N_7639);
and U11798 (N_11798,N_8757,N_8724);
nor U11799 (N_11799,N_7453,N_7327);
nand U11800 (N_11800,N_8374,N_6077);
and U11801 (N_11801,N_8186,N_6041);
nor U11802 (N_11802,N_8233,N_7334);
and U11803 (N_11803,N_8045,N_7009);
and U11804 (N_11804,N_8420,N_7170);
or U11805 (N_11805,N_6008,N_6671);
and U11806 (N_11806,N_8588,N_8681);
xnor U11807 (N_11807,N_8389,N_7643);
and U11808 (N_11808,N_7436,N_7430);
nor U11809 (N_11809,N_8259,N_8786);
or U11810 (N_11810,N_6581,N_8734);
nor U11811 (N_11811,N_7562,N_8561);
or U11812 (N_11812,N_6370,N_6322);
and U11813 (N_11813,N_8925,N_6348);
nand U11814 (N_11814,N_8944,N_7455);
xor U11815 (N_11815,N_7816,N_7971);
nand U11816 (N_11816,N_8847,N_7062);
nor U11817 (N_11817,N_8594,N_7054);
nand U11818 (N_11818,N_6859,N_7641);
nor U11819 (N_11819,N_8722,N_7231);
nand U11820 (N_11820,N_7495,N_6270);
nand U11821 (N_11821,N_6428,N_6670);
nand U11822 (N_11822,N_8738,N_6936);
nor U11823 (N_11823,N_7235,N_6336);
nor U11824 (N_11824,N_8890,N_6397);
xor U11825 (N_11825,N_8335,N_6446);
and U11826 (N_11826,N_7095,N_6569);
and U11827 (N_11827,N_6846,N_7285);
nor U11828 (N_11828,N_7908,N_8675);
nand U11829 (N_11829,N_8976,N_6717);
nand U11830 (N_11830,N_8124,N_8158);
xnor U11831 (N_11831,N_7597,N_8789);
or U11832 (N_11832,N_8083,N_8730);
or U11833 (N_11833,N_7429,N_8354);
or U11834 (N_11834,N_8983,N_6803);
or U11835 (N_11835,N_8793,N_6277);
or U11836 (N_11836,N_6323,N_8507);
and U11837 (N_11837,N_8810,N_7306);
and U11838 (N_11838,N_7117,N_6052);
or U11839 (N_11839,N_8266,N_6068);
nand U11840 (N_11840,N_7556,N_7293);
or U11841 (N_11841,N_7692,N_6921);
xnor U11842 (N_11842,N_8427,N_6439);
nor U11843 (N_11843,N_8923,N_7351);
and U11844 (N_11844,N_8070,N_7141);
nand U11845 (N_11845,N_7306,N_6233);
and U11846 (N_11846,N_6355,N_6127);
xor U11847 (N_11847,N_6691,N_8562);
nor U11848 (N_11848,N_7166,N_6664);
nand U11849 (N_11849,N_6211,N_6763);
xor U11850 (N_11850,N_7723,N_8437);
and U11851 (N_11851,N_6633,N_7506);
and U11852 (N_11852,N_6311,N_7472);
nor U11853 (N_11853,N_6869,N_8841);
nor U11854 (N_11854,N_6195,N_8952);
nand U11855 (N_11855,N_8767,N_7447);
or U11856 (N_11856,N_7307,N_8045);
nand U11857 (N_11857,N_6492,N_8467);
or U11858 (N_11858,N_8561,N_8508);
and U11859 (N_11859,N_8947,N_8340);
and U11860 (N_11860,N_7847,N_6494);
nor U11861 (N_11861,N_6846,N_8495);
xor U11862 (N_11862,N_6067,N_8324);
and U11863 (N_11863,N_6910,N_7658);
or U11864 (N_11864,N_7651,N_7993);
nand U11865 (N_11865,N_8430,N_6635);
and U11866 (N_11866,N_8205,N_7687);
nor U11867 (N_11867,N_8690,N_7620);
and U11868 (N_11868,N_8494,N_8330);
nor U11869 (N_11869,N_8952,N_8571);
and U11870 (N_11870,N_7663,N_8095);
xor U11871 (N_11871,N_8279,N_8234);
and U11872 (N_11872,N_7894,N_8415);
and U11873 (N_11873,N_6646,N_7627);
xor U11874 (N_11874,N_8303,N_7380);
nor U11875 (N_11875,N_7635,N_6374);
xor U11876 (N_11876,N_6806,N_8263);
nor U11877 (N_11877,N_6447,N_7158);
nor U11878 (N_11878,N_8335,N_6689);
nor U11879 (N_11879,N_6944,N_8504);
xor U11880 (N_11880,N_7069,N_6633);
xor U11881 (N_11881,N_8980,N_8257);
xor U11882 (N_11882,N_7759,N_8302);
xnor U11883 (N_11883,N_6773,N_8996);
and U11884 (N_11884,N_7861,N_8932);
xnor U11885 (N_11885,N_7203,N_8357);
nor U11886 (N_11886,N_7292,N_7802);
or U11887 (N_11887,N_6664,N_6521);
xor U11888 (N_11888,N_7984,N_7944);
nand U11889 (N_11889,N_6069,N_6005);
or U11890 (N_11890,N_8644,N_7877);
or U11891 (N_11891,N_7492,N_6190);
nor U11892 (N_11892,N_7562,N_8548);
nand U11893 (N_11893,N_8743,N_7414);
nand U11894 (N_11894,N_8856,N_7274);
nand U11895 (N_11895,N_8154,N_8117);
xnor U11896 (N_11896,N_6177,N_8431);
nand U11897 (N_11897,N_6594,N_8066);
nor U11898 (N_11898,N_7684,N_6450);
nand U11899 (N_11899,N_8575,N_6628);
or U11900 (N_11900,N_7048,N_7023);
nand U11901 (N_11901,N_6806,N_7900);
xnor U11902 (N_11902,N_8934,N_6794);
or U11903 (N_11903,N_6226,N_6723);
xnor U11904 (N_11904,N_8073,N_8025);
nor U11905 (N_11905,N_6987,N_6699);
or U11906 (N_11906,N_6481,N_7827);
and U11907 (N_11907,N_7028,N_7228);
nor U11908 (N_11908,N_7432,N_8707);
xor U11909 (N_11909,N_7036,N_6268);
nand U11910 (N_11910,N_7738,N_6124);
nor U11911 (N_11911,N_6356,N_7704);
nor U11912 (N_11912,N_6193,N_7273);
nand U11913 (N_11913,N_8000,N_7237);
nand U11914 (N_11914,N_8353,N_7987);
or U11915 (N_11915,N_8726,N_6092);
xor U11916 (N_11916,N_6703,N_8655);
xor U11917 (N_11917,N_8190,N_6125);
nor U11918 (N_11918,N_6564,N_8662);
nor U11919 (N_11919,N_7307,N_6439);
nor U11920 (N_11920,N_7222,N_8619);
nor U11921 (N_11921,N_7893,N_8074);
nor U11922 (N_11922,N_6668,N_7396);
nor U11923 (N_11923,N_7126,N_6306);
or U11924 (N_11924,N_8350,N_6452);
or U11925 (N_11925,N_7038,N_7897);
nand U11926 (N_11926,N_6300,N_7752);
and U11927 (N_11927,N_8328,N_8719);
and U11928 (N_11928,N_6378,N_6480);
or U11929 (N_11929,N_8246,N_6781);
nor U11930 (N_11930,N_7270,N_6147);
nand U11931 (N_11931,N_8790,N_6362);
nor U11932 (N_11932,N_7506,N_7916);
nand U11933 (N_11933,N_6732,N_6708);
nand U11934 (N_11934,N_7368,N_7293);
and U11935 (N_11935,N_8641,N_8236);
xnor U11936 (N_11936,N_7263,N_7974);
nand U11937 (N_11937,N_7682,N_6224);
xnor U11938 (N_11938,N_8569,N_8280);
or U11939 (N_11939,N_6186,N_7634);
nand U11940 (N_11940,N_7793,N_6520);
xnor U11941 (N_11941,N_7050,N_6548);
and U11942 (N_11942,N_8765,N_8363);
and U11943 (N_11943,N_6403,N_8039);
nand U11944 (N_11944,N_6395,N_8441);
and U11945 (N_11945,N_8681,N_6096);
or U11946 (N_11946,N_6485,N_7803);
nand U11947 (N_11947,N_8827,N_7180);
xnor U11948 (N_11948,N_8151,N_6639);
xnor U11949 (N_11949,N_7369,N_6936);
or U11950 (N_11950,N_8375,N_6557);
and U11951 (N_11951,N_7376,N_8164);
and U11952 (N_11952,N_6746,N_7912);
nand U11953 (N_11953,N_8474,N_6881);
nand U11954 (N_11954,N_6201,N_8250);
and U11955 (N_11955,N_7085,N_6403);
or U11956 (N_11956,N_8269,N_8327);
and U11957 (N_11957,N_7908,N_8440);
and U11958 (N_11958,N_6880,N_6682);
or U11959 (N_11959,N_7229,N_8074);
or U11960 (N_11960,N_8396,N_6770);
nor U11961 (N_11961,N_7542,N_8265);
or U11962 (N_11962,N_6620,N_8065);
nand U11963 (N_11963,N_8824,N_7188);
nand U11964 (N_11964,N_8952,N_6738);
and U11965 (N_11965,N_8994,N_6871);
or U11966 (N_11966,N_8858,N_7297);
xnor U11967 (N_11967,N_8176,N_8265);
and U11968 (N_11968,N_7744,N_6218);
and U11969 (N_11969,N_6955,N_7029);
and U11970 (N_11970,N_6961,N_7915);
nand U11971 (N_11971,N_8181,N_7008);
or U11972 (N_11972,N_6634,N_6654);
xor U11973 (N_11973,N_8465,N_8954);
nor U11974 (N_11974,N_8691,N_6293);
nand U11975 (N_11975,N_8256,N_6898);
xor U11976 (N_11976,N_8984,N_7295);
nor U11977 (N_11977,N_8175,N_8489);
or U11978 (N_11978,N_8456,N_8884);
xnor U11979 (N_11979,N_8384,N_6719);
or U11980 (N_11980,N_6990,N_8198);
nand U11981 (N_11981,N_6299,N_8829);
nor U11982 (N_11982,N_8627,N_6355);
nor U11983 (N_11983,N_7532,N_7319);
nor U11984 (N_11984,N_8091,N_8113);
nand U11985 (N_11985,N_7840,N_7452);
xor U11986 (N_11986,N_6833,N_7904);
or U11987 (N_11987,N_6666,N_8291);
nor U11988 (N_11988,N_8604,N_8148);
xor U11989 (N_11989,N_7698,N_8269);
or U11990 (N_11990,N_7659,N_7013);
nand U11991 (N_11991,N_7178,N_8179);
and U11992 (N_11992,N_6452,N_7029);
nand U11993 (N_11993,N_6111,N_6090);
and U11994 (N_11994,N_7331,N_6177);
or U11995 (N_11995,N_8110,N_7674);
or U11996 (N_11996,N_8988,N_7629);
nor U11997 (N_11997,N_6043,N_7210);
nor U11998 (N_11998,N_7377,N_6919);
nand U11999 (N_11999,N_6674,N_8187);
nor U12000 (N_12000,N_10313,N_10326);
or U12001 (N_12001,N_11345,N_9401);
nor U12002 (N_12002,N_9189,N_9122);
xnor U12003 (N_12003,N_9225,N_11287);
and U12004 (N_12004,N_11024,N_9001);
or U12005 (N_12005,N_11384,N_11239);
xor U12006 (N_12006,N_10893,N_11919);
or U12007 (N_12007,N_10422,N_11255);
or U12008 (N_12008,N_10700,N_9452);
and U12009 (N_12009,N_10290,N_11774);
or U12010 (N_12010,N_11839,N_11124);
nor U12011 (N_12011,N_9118,N_11265);
and U12012 (N_12012,N_10607,N_10726);
nand U12013 (N_12013,N_9781,N_10357);
nand U12014 (N_12014,N_11521,N_9424);
nand U12015 (N_12015,N_11565,N_9346);
nor U12016 (N_12016,N_10333,N_11967);
xnor U12017 (N_12017,N_9187,N_11496);
or U12018 (N_12018,N_10033,N_11787);
nand U12019 (N_12019,N_11566,N_9921);
and U12020 (N_12020,N_11497,N_11708);
or U12021 (N_12021,N_11146,N_10072);
nand U12022 (N_12022,N_9762,N_10104);
nand U12023 (N_12023,N_10111,N_10904);
xor U12024 (N_12024,N_10585,N_10858);
nor U12025 (N_12025,N_11102,N_9653);
xor U12026 (N_12026,N_11554,N_11508);
or U12027 (N_12027,N_9635,N_10289);
nand U12028 (N_12028,N_9787,N_10828);
nand U12029 (N_12029,N_11529,N_11025);
and U12030 (N_12030,N_10991,N_9940);
or U12031 (N_12031,N_11625,N_11023);
nand U12032 (N_12032,N_11151,N_11224);
nor U12033 (N_12033,N_11471,N_9736);
or U12034 (N_12034,N_10508,N_10261);
and U12035 (N_12035,N_10322,N_11792);
and U12036 (N_12036,N_10186,N_9568);
nand U12037 (N_12037,N_11030,N_9768);
nand U12038 (N_12038,N_11322,N_11998);
and U12039 (N_12039,N_10952,N_11600);
xnor U12040 (N_12040,N_9116,N_10910);
and U12041 (N_12041,N_11428,N_11973);
or U12042 (N_12042,N_9528,N_10778);
or U12043 (N_12043,N_10579,N_9987);
xnor U12044 (N_12044,N_9851,N_10405);
nor U12045 (N_12045,N_10716,N_11658);
and U12046 (N_12046,N_10065,N_10757);
nand U12047 (N_12047,N_10773,N_11890);
xor U12048 (N_12048,N_10601,N_9922);
xor U12049 (N_12049,N_11988,N_11573);
or U12050 (N_12050,N_10349,N_11002);
or U12051 (N_12051,N_9429,N_11835);
or U12052 (N_12052,N_9703,N_9780);
and U12053 (N_12053,N_9980,N_10399);
or U12054 (N_12054,N_9010,N_10285);
xor U12055 (N_12055,N_10783,N_10061);
xnor U12056 (N_12056,N_9302,N_10552);
nand U12057 (N_12057,N_9510,N_10701);
or U12058 (N_12058,N_9735,N_9591);
and U12059 (N_12059,N_9869,N_11810);
nor U12060 (N_12060,N_9953,N_11088);
nor U12061 (N_12061,N_9173,N_9976);
and U12062 (N_12062,N_10846,N_9821);
nor U12063 (N_12063,N_10721,N_10587);
or U12064 (N_12064,N_10990,N_11164);
or U12065 (N_12065,N_9795,N_11041);
or U12066 (N_12066,N_9998,N_9504);
nand U12067 (N_12067,N_11672,N_10613);
nand U12068 (N_12068,N_11905,N_11781);
or U12069 (N_12069,N_10364,N_9737);
nor U12070 (N_12070,N_9501,N_10791);
nand U12071 (N_12071,N_10424,N_11756);
or U12072 (N_12072,N_9517,N_11376);
xnor U12073 (N_12073,N_11409,N_9358);
or U12074 (N_12074,N_11270,N_9476);
nor U12075 (N_12075,N_9878,N_10848);
xnor U12076 (N_12076,N_9624,N_10831);
and U12077 (N_12077,N_9601,N_9293);
and U12078 (N_12078,N_9321,N_9607);
nor U12079 (N_12079,N_9082,N_9299);
xor U12080 (N_12080,N_10220,N_10095);
or U12081 (N_12081,N_11156,N_9433);
or U12082 (N_12082,N_10907,N_11033);
nand U12083 (N_12083,N_9563,N_10949);
or U12084 (N_12084,N_9551,N_10435);
or U12085 (N_12085,N_9755,N_9988);
xnor U12086 (N_12086,N_9231,N_9221);
or U12087 (N_12087,N_9718,N_11056);
nor U12088 (N_12088,N_11414,N_11811);
nor U12089 (N_12089,N_10666,N_10837);
or U12090 (N_12090,N_11460,N_11140);
and U12091 (N_12091,N_11558,N_11855);
xnor U12092 (N_12092,N_9398,N_9388);
nor U12093 (N_12093,N_9954,N_10488);
or U12094 (N_12094,N_10170,N_10352);
and U12095 (N_12095,N_11451,N_11216);
nand U12096 (N_12096,N_11609,N_9806);
nor U12097 (N_12097,N_9372,N_9005);
nor U12098 (N_12098,N_9628,N_10255);
nand U12099 (N_12099,N_10808,N_9532);
nor U12100 (N_12100,N_10087,N_10180);
nor U12101 (N_12101,N_11860,N_10648);
or U12102 (N_12102,N_10854,N_10473);
nand U12103 (N_12103,N_9909,N_9838);
nand U12104 (N_12104,N_11344,N_10015);
nor U12105 (N_12105,N_11116,N_9678);
and U12106 (N_12106,N_9746,N_11805);
nor U12107 (N_12107,N_10943,N_11780);
xor U12108 (N_12108,N_10630,N_10467);
and U12109 (N_12109,N_9468,N_10489);
xnor U12110 (N_12110,N_9195,N_11010);
and U12111 (N_12111,N_11858,N_9884);
or U12112 (N_12112,N_10679,N_9769);
or U12113 (N_12113,N_9182,N_10169);
and U12114 (N_12114,N_10525,N_11570);
nand U12115 (N_12115,N_11346,N_11293);
or U12116 (N_12116,N_11433,N_9114);
nor U12117 (N_12117,N_9232,N_11831);
and U12118 (N_12118,N_11739,N_9077);
nand U12119 (N_12119,N_9576,N_9169);
nor U12120 (N_12120,N_9991,N_9667);
and U12121 (N_12121,N_10766,N_11348);
nand U12122 (N_12122,N_9101,N_9334);
nand U12123 (N_12123,N_10271,N_9380);
or U12124 (N_12124,N_11753,N_9257);
nor U12125 (N_12125,N_11992,N_9471);
xnor U12126 (N_12126,N_9417,N_10076);
nand U12127 (N_12127,N_11013,N_10763);
nor U12128 (N_12128,N_11142,N_9212);
nor U12129 (N_12129,N_10542,N_11371);
nor U12130 (N_12130,N_11418,N_11581);
nand U12131 (N_12131,N_9125,N_10785);
or U12132 (N_12132,N_10121,N_11583);
or U12133 (N_12133,N_11877,N_9834);
xnor U12134 (N_12134,N_10363,N_10671);
and U12135 (N_12135,N_10284,N_9845);
and U12136 (N_12136,N_9920,N_10479);
or U12137 (N_12137,N_9885,N_10491);
xnor U12138 (N_12138,N_9801,N_11368);
or U12139 (N_12139,N_10674,N_10761);
nand U12140 (N_12140,N_10970,N_10400);
and U12141 (N_12141,N_10633,N_9274);
or U12142 (N_12142,N_11136,N_11706);
or U12143 (N_12143,N_10862,N_10042);
nand U12144 (N_12144,N_11607,N_10030);
xnor U12145 (N_12145,N_9606,N_10737);
nor U12146 (N_12146,N_9547,N_10518);
nand U12147 (N_12147,N_10299,N_9590);
or U12148 (N_12148,N_9758,N_10682);
and U12149 (N_12149,N_10870,N_9013);
xor U12150 (N_12150,N_9712,N_9587);
and U12151 (N_12151,N_10090,N_9081);
xor U12152 (N_12152,N_9461,N_9256);
and U12153 (N_12153,N_11203,N_10138);
or U12154 (N_12154,N_10233,N_9665);
nand U12155 (N_12155,N_9295,N_11982);
and U12156 (N_12156,N_9854,N_11684);
xnor U12157 (N_12157,N_11685,N_11430);
nor U12158 (N_12158,N_11489,N_9642);
nand U12159 (N_12159,N_9196,N_9670);
nor U12160 (N_12160,N_9032,N_10523);
or U12161 (N_12161,N_9155,N_10824);
or U12162 (N_12162,N_11107,N_10063);
or U12163 (N_12163,N_11511,N_10227);
nor U12164 (N_12164,N_10654,N_11734);
xor U12165 (N_12165,N_11037,N_10114);
and U12166 (N_12166,N_10342,N_9350);
or U12167 (N_12167,N_10845,N_9278);
xnor U12168 (N_12168,N_11655,N_11021);
nand U12169 (N_12169,N_11372,N_10484);
nor U12170 (N_12170,N_9638,N_9457);
and U12171 (N_12171,N_9098,N_10146);
and U12172 (N_12172,N_11411,N_11777);
or U12173 (N_12173,N_10698,N_11130);
xor U12174 (N_12174,N_11507,N_11247);
nand U12175 (N_12175,N_10296,N_9965);
xnor U12176 (N_12176,N_9719,N_9259);
nand U12177 (N_12177,N_10964,N_9338);
xnor U12178 (N_12178,N_11246,N_11909);
and U12179 (N_12179,N_10101,N_9695);
or U12180 (N_12180,N_10141,N_11165);
and U12181 (N_12181,N_9161,N_10059);
nand U12182 (N_12182,N_9156,N_10250);
or U12183 (N_12183,N_10989,N_9199);
nand U12184 (N_12184,N_9031,N_11343);
nand U12185 (N_12185,N_9033,N_10971);
nand U12186 (N_12186,N_11606,N_10834);
nand U12187 (N_12187,N_9109,N_10126);
nor U12188 (N_12188,N_11269,N_11532);
and U12189 (N_12189,N_11485,N_10743);
nand U12190 (N_12190,N_9558,N_11274);
and U12191 (N_12191,N_9876,N_11957);
nor U12192 (N_12192,N_9798,N_11044);
and U12193 (N_12193,N_11398,N_11744);
nand U12194 (N_12194,N_11481,N_10093);
nor U12195 (N_12195,N_11280,N_11295);
xor U12196 (N_12196,N_11822,N_10890);
nand U12197 (N_12197,N_9222,N_11564);
or U12198 (N_12198,N_11236,N_11561);
nor U12199 (N_12199,N_10177,N_9400);
nor U12200 (N_12200,N_9102,N_11468);
xor U12201 (N_12201,N_9023,N_11079);
nor U12202 (N_12202,N_9577,N_9469);
and U12203 (N_12203,N_11784,N_11159);
nand U12204 (N_12204,N_11050,N_11148);
or U12205 (N_12205,N_11878,N_11965);
nand U12206 (N_12206,N_10041,N_11986);
nor U12207 (N_12207,N_10874,N_11698);
xnor U12208 (N_12208,N_9272,N_11046);
or U12209 (N_12209,N_9201,N_11580);
and U12210 (N_12210,N_11198,N_11456);
or U12211 (N_12211,N_11557,N_9121);
nand U12212 (N_12212,N_11892,N_11347);
xnor U12213 (N_12213,N_10639,N_10925);
nor U12214 (N_12214,N_10811,N_11197);
nor U12215 (N_12215,N_9766,N_10641);
xnor U12216 (N_12216,N_10549,N_10018);
xnor U12217 (N_12217,N_9773,N_9849);
nor U12218 (N_12218,N_9608,N_9038);
or U12219 (N_12219,N_10591,N_11796);
xnor U12220 (N_12220,N_10206,N_9213);
xor U12221 (N_12221,N_9880,N_11874);
and U12222 (N_12222,N_9068,N_9206);
xnor U12223 (N_12223,N_10440,N_9680);
xor U12224 (N_12224,N_11066,N_11168);
nand U12225 (N_12225,N_11183,N_10691);
nand U12226 (N_12226,N_10600,N_9453);
or U12227 (N_12227,N_10764,N_9713);
and U12228 (N_12228,N_9062,N_10596);
nand U12229 (N_12229,N_11128,N_11331);
or U12230 (N_12230,N_11989,N_10779);
nor U12231 (N_12231,N_9384,N_9145);
and U12232 (N_12232,N_11445,N_9085);
nor U12233 (N_12233,N_11305,N_10071);
nand U12234 (N_12234,N_10175,N_11918);
and U12235 (N_12235,N_10280,N_9464);
nand U12236 (N_12236,N_9345,N_10000);
nor U12237 (N_12237,N_10781,N_9333);
nor U12238 (N_12238,N_9900,N_10684);
nor U12239 (N_12239,N_9552,N_10362);
nand U12240 (N_12240,N_11432,N_11826);
nand U12241 (N_12241,N_9675,N_10960);
nand U12242 (N_12242,N_10941,N_10835);
and U12243 (N_12243,N_9809,N_11427);
xor U12244 (N_12244,N_10643,N_9726);
or U12245 (N_12245,N_10911,N_11782);
xor U12246 (N_12246,N_9579,N_9767);
or U12247 (N_12247,N_9414,N_10192);
nor U12248 (N_12248,N_10324,N_10618);
nor U12249 (N_12249,N_11632,N_9438);
nand U12250 (N_12250,N_11263,N_9743);
xnor U12251 (N_12251,N_9306,N_9390);
xnor U12252 (N_12252,N_11399,N_10795);
or U12253 (N_12253,N_10096,N_9721);
nor U12254 (N_12254,N_10912,N_9336);
or U12255 (N_12255,N_9915,N_11424);
nand U12256 (N_12256,N_10133,N_11127);
or U12257 (N_12257,N_11902,N_11184);
nand U12258 (N_12258,N_10210,N_9616);
nand U12259 (N_12259,N_10117,N_11995);
nor U12260 (N_12260,N_9679,N_9699);
nor U12261 (N_12261,N_9725,N_9403);
or U12262 (N_12262,N_9454,N_9430);
and U12263 (N_12263,N_11061,N_10305);
or U12264 (N_12264,N_11549,N_11326);
nand U12265 (N_12265,N_9382,N_9238);
or U12266 (N_12266,N_10401,N_9111);
or U12267 (N_12267,N_10985,N_10199);
or U12268 (N_12268,N_9513,N_10021);
and U12269 (N_12269,N_11644,N_11610);
xor U12270 (N_12270,N_10026,N_11555);
or U12271 (N_12271,N_11611,N_10200);
nand U12272 (N_12272,N_10685,N_9506);
or U12273 (N_12273,N_11510,N_9378);
xor U12274 (N_12274,N_9979,N_11334);
or U12275 (N_12275,N_10724,N_11694);
nand U12276 (N_12276,N_9701,N_11426);
or U12277 (N_12277,N_9054,N_9439);
or U12278 (N_12278,N_10526,N_11891);
nor U12279 (N_12279,N_10827,N_10244);
and U12280 (N_12280,N_11517,N_11300);
xnor U12281 (N_12281,N_11117,N_10487);
nand U12282 (N_12282,N_9200,N_10900);
nor U12283 (N_12283,N_9738,N_9782);
xnor U12284 (N_12284,N_11009,N_11111);
xor U12285 (N_12285,N_9441,N_11126);
nand U12286 (N_12286,N_9927,N_10856);
or U12287 (N_12287,N_11962,N_10775);
nor U12288 (N_12288,N_9727,N_11930);
nand U12289 (N_12289,N_10547,N_10536);
or U12290 (N_12290,N_10664,N_11803);
and U12291 (N_12291,N_9749,N_10988);
xor U12292 (N_12292,N_11390,N_9599);
or U12293 (N_12293,N_10201,N_11543);
xor U12294 (N_12294,N_10798,N_10570);
xor U12295 (N_12295,N_11848,N_9947);
xor U12296 (N_12296,N_10036,N_11923);
nor U12297 (N_12297,N_9300,N_9648);
nand U12298 (N_12298,N_10646,N_10402);
nand U12299 (N_12299,N_10888,N_9170);
xor U12300 (N_12300,N_9202,N_9567);
and U12301 (N_12301,N_10350,N_9126);
or U12302 (N_12302,N_9919,N_10564);
nor U12303 (N_12303,N_10413,N_10656);
xor U12304 (N_12304,N_11463,N_9765);
nor U12305 (N_12305,N_10094,N_11022);
nor U12306 (N_12306,N_9522,N_9264);
and U12307 (N_12307,N_10840,N_10476);
nand U12308 (N_12308,N_10575,N_9741);
and U12309 (N_12309,N_10797,N_11642);
xnor U12310 (N_12310,N_10441,N_9584);
and U12311 (N_12311,N_9561,N_9818);
nor U12312 (N_12312,N_11700,N_10754);
xnor U12313 (N_12313,N_11048,N_9764);
nor U12314 (N_12314,N_10158,N_9562);
and U12315 (N_12315,N_10876,N_11656);
nor U12316 (N_12316,N_9978,N_9381);
xor U12317 (N_12317,N_10624,N_10038);
and U12318 (N_12318,N_11400,N_11181);
or U12319 (N_12319,N_10493,N_10092);
or U12320 (N_12320,N_9520,N_11571);
nor U12321 (N_12321,N_11940,N_10696);
or U12322 (N_12322,N_10729,N_10875);
or U12323 (N_12323,N_11683,N_11211);
nand U12324 (N_12324,N_9369,N_10714);
or U12325 (N_12325,N_9158,N_10332);
or U12326 (N_12326,N_10687,N_11219);
nand U12327 (N_12327,N_11171,N_9269);
nor U12328 (N_12328,N_10728,N_10617);
xor U12329 (N_12329,N_10431,N_9630);
and U12330 (N_12330,N_10360,N_11604);
nand U12331 (N_12331,N_11779,N_9024);
nor U12332 (N_12332,N_11064,N_10712);
and U12333 (N_12333,N_9009,N_11568);
nand U12334 (N_12334,N_9941,N_10892);
nand U12335 (N_12335,N_10753,N_9324);
or U12336 (N_12336,N_9949,N_11636);
xor U12337 (N_12337,N_11282,N_10468);
and U12338 (N_12338,N_9950,N_10164);
and U12339 (N_12339,N_11804,N_9545);
and U12340 (N_12340,N_11715,N_10527);
nand U12341 (N_12341,N_11546,N_11473);
nand U12342 (N_12342,N_9308,N_9497);
xor U12343 (N_12343,N_11985,N_10241);
nand U12344 (N_12344,N_11824,N_10385);
nor U12345 (N_12345,N_9004,N_10514);
or U12346 (N_12346,N_10788,N_11693);
or U12347 (N_12347,N_10436,N_9487);
nand U12348 (N_12348,N_11383,N_11394);
nor U12349 (N_12349,N_10929,N_10913);
nor U12350 (N_12350,N_9794,N_11846);
nand U12351 (N_12351,N_9602,N_10512);
or U12352 (N_12352,N_10669,N_11603);
nand U12353 (N_12353,N_9135,N_11089);
or U12354 (N_12354,N_9825,N_11264);
or U12355 (N_12355,N_10995,N_10558);
or U12356 (N_12356,N_11637,N_10833);
nor U12357 (N_12357,N_9808,N_10389);
xnor U12358 (N_12358,N_10474,N_11078);
or U12359 (N_12359,N_11155,N_11526);
xor U12360 (N_12360,N_9582,N_9003);
xnor U12361 (N_12361,N_11752,N_11338);
or U12362 (N_12362,N_11647,N_9219);
nor U12363 (N_12363,N_9759,N_9152);
xor U12364 (N_12364,N_11360,N_10454);
and U12365 (N_12365,N_10667,N_11340);
nor U12366 (N_12366,N_9788,N_10231);
xor U12367 (N_12367,N_9347,N_9143);
and U12368 (N_12368,N_10425,N_11235);
or U12369 (N_12369,N_9373,N_11385);
and U12370 (N_12370,N_11240,N_11416);
or U12371 (N_12371,N_9702,N_9053);
nand U12372 (N_12372,N_10377,N_11429);
or U12373 (N_12373,N_10166,N_10148);
and U12374 (N_12374,N_9374,N_11776);
xor U12375 (N_12375,N_9756,N_11868);
nor U12376 (N_12376,N_11733,N_11315);
nor U12377 (N_12377,N_9521,N_9227);
nor U12378 (N_12378,N_10823,N_9249);
xor U12379 (N_12379,N_11873,N_10309);
nor U12380 (N_12380,N_9783,N_10394);
or U12381 (N_12381,N_9981,N_11916);
and U12382 (N_12382,N_9681,N_11243);
or U12383 (N_12383,N_11951,N_9907);
nor U12384 (N_12384,N_11178,N_9511);
and U12385 (N_12385,N_10242,N_10722);
and U12386 (N_12386,N_9750,N_11807);
or U12387 (N_12387,N_9828,N_9729);
and U12388 (N_12388,N_11289,N_9399);
nand U12389 (N_12389,N_11176,N_11623);
and U12390 (N_12390,N_11323,N_10275);
nand U12391 (N_12391,N_10403,N_10125);
nand U12392 (N_12392,N_11249,N_9140);
or U12393 (N_12393,N_9811,N_10608);
nor U12394 (N_12394,N_10992,N_9856);
or U12395 (N_12395,N_9619,N_9816);
xnor U12396 (N_12396,N_9903,N_10713);
nand U12397 (N_12397,N_11195,N_10356);
nor U12398 (N_12398,N_11585,N_10909);
nor U12399 (N_12399,N_9254,N_10532);
nand U12400 (N_12400,N_11727,N_9252);
nor U12401 (N_12401,N_11038,N_9641);
nor U12402 (N_12402,N_10216,N_9436);
or U12403 (N_12403,N_10872,N_10237);
or U12404 (N_12404,N_11370,N_10588);
and U12405 (N_12405,N_9803,N_9659);
and U12406 (N_12406,N_10062,N_10168);
xor U12407 (N_12407,N_10611,N_11053);
or U12408 (N_12408,N_11129,N_11936);
or U12409 (N_12409,N_9560,N_11169);
and U12410 (N_12410,N_10853,N_10122);
or U12411 (N_12411,N_9644,N_10470);
xnor U12412 (N_12412,N_11499,N_10940);
nand U12413 (N_12413,N_10882,N_10083);
and U12414 (N_12414,N_11039,N_9315);
or U12415 (N_12415,N_10478,N_11791);
nor U12416 (N_12416,N_10595,N_9847);
nor U12417 (N_12417,N_11761,N_9385);
xnor U12418 (N_12418,N_11045,N_10129);
xor U12419 (N_12419,N_11864,N_10963);
nand U12420 (N_12420,N_10054,N_10822);
xor U12421 (N_12421,N_10139,N_9993);
xor U12422 (N_12422,N_9757,N_9533);
nand U12423 (N_12423,N_9419,N_10393);
and U12424 (N_12424,N_10844,N_9105);
xor U12425 (N_12425,N_9181,N_9508);
xnor U12426 (N_12426,N_9117,N_10272);
and U12427 (N_12427,N_11968,N_10770);
nand U12428 (N_12428,N_10746,N_10965);
nand U12429 (N_12429,N_11457,N_10251);
nand U12430 (N_12430,N_9610,N_9831);
nor U12431 (N_12431,N_10723,N_11929);
xor U12432 (N_12432,N_9914,N_10477);
or U12433 (N_12433,N_9198,N_11579);
or U12434 (N_12434,N_9583,N_10293);
nor U12435 (N_12435,N_10418,N_10014);
nand U12436 (N_12436,N_11448,N_11705);
nand U12437 (N_12437,N_9214,N_11477);
nand U12438 (N_12438,N_10359,N_9556);
nor U12439 (N_12439,N_9074,N_11339);
xnor U12440 (N_12440,N_9050,N_11505);
or U12441 (N_12441,N_9128,N_9039);
xor U12442 (N_12442,N_9800,N_11987);
or U12443 (N_12443,N_9890,N_11087);
xor U12444 (N_12444,N_9790,N_9844);
or U12445 (N_12445,N_10632,N_10548);
xnor U12446 (N_12446,N_10453,N_10456);
xor U12447 (N_12447,N_11091,N_11072);
xnor U12448 (N_12448,N_11185,N_11498);
and U12449 (N_12449,N_9444,N_9580);
and U12450 (N_12450,N_10442,N_11302);
and U12451 (N_12451,N_9744,N_11110);
nor U12452 (N_12452,N_9985,N_10123);
xnor U12453 (N_12453,N_10005,N_10416);
nor U12454 (N_12454,N_10124,N_10306);
or U12455 (N_12455,N_11166,N_9633);
and U12456 (N_12456,N_9426,N_10528);
or U12457 (N_12457,N_9715,N_9804);
and U12458 (N_12458,N_9925,N_10673);
and U12459 (N_12459,N_11530,N_9326);
xor U12460 (N_12460,N_10957,N_10246);
nand U12461 (N_12461,N_9011,N_10612);
xnor U12462 (N_12462,N_11248,N_11365);
nand U12463 (N_12463,N_11054,N_11502);
nand U12464 (N_12464,N_9605,N_10860);
xnor U12465 (N_12465,N_10850,N_11643);
nor U12466 (N_12466,N_11098,N_9711);
and U12467 (N_12467,N_9184,N_11308);
nor U12468 (N_12468,N_10173,N_9311);
nor U12469 (N_12469,N_10006,N_11225);
nand U12470 (N_12470,N_9867,N_9923);
or U12471 (N_12471,N_9029,N_11258);
xnor U12472 (N_12472,N_10353,N_9281);
nand U12473 (N_12473,N_9056,N_10559);
and U12474 (N_12474,N_10574,N_9945);
nand U12475 (N_12475,N_10278,N_10247);
or U12476 (N_12476,N_9028,N_9176);
or U12477 (N_12477,N_10144,N_9707);
or U12478 (N_12478,N_9643,N_11093);
nor U12479 (N_12479,N_11139,N_9622);
nor U12480 (N_12480,N_11619,N_10235);
nand U12481 (N_12481,N_9594,N_11482);
nor U12482 (N_12482,N_11844,N_11194);
nor U12483 (N_12483,N_9215,N_9770);
xnor U12484 (N_12484,N_11267,N_11653);
and U12485 (N_12485,N_11153,N_11682);
xnor U12486 (N_12486,N_9304,N_10942);
nand U12487 (N_12487,N_9217,N_10610);
and U12488 (N_12488,N_9428,N_9518);
or U12489 (N_12489,N_10398,N_9708);
xor U12490 (N_12490,N_9686,N_11931);
nand U12491 (N_12491,N_9629,N_9235);
xnor U12492 (N_12492,N_9955,N_9022);
nor U12493 (N_12493,N_10603,N_11335);
or U12494 (N_12494,N_9422,N_10908);
nand U12495 (N_12495,N_11837,N_10543);
xor U12496 (N_12496,N_11336,N_10919);
nand U12497 (N_12497,N_9442,N_11057);
or U12498 (N_12498,N_11944,N_11309);
nor U12499 (N_12499,N_9065,N_11108);
nor U12500 (N_12500,N_9070,N_9246);
nor U12501 (N_12501,N_9134,N_9092);
nor U12502 (N_12502,N_11605,N_9455);
or U12503 (N_12503,N_11677,N_10259);
or U12504 (N_12504,N_10939,N_11541);
nor U12505 (N_12505,N_10501,N_10039);
nor U12506 (N_12506,N_9443,N_11884);
or U12507 (N_12507,N_10510,N_9097);
and U12508 (N_12508,N_9110,N_11516);
and U12509 (N_12509,N_11154,N_11217);
xor U12510 (N_12510,N_10159,N_9078);
xor U12511 (N_12511,N_9984,N_10819);
or U12512 (N_12512,N_10650,N_9971);
nand U12513 (N_12513,N_9992,N_11567);
nor U12514 (N_12514,N_11205,N_9185);
nor U12515 (N_12515,N_11620,N_10719);
xor U12516 (N_12516,N_9833,N_11645);
and U12517 (N_12517,N_11597,N_10787);
and U12518 (N_12518,N_10924,N_11459);
nand U12519 (N_12519,N_10735,N_11068);
xnor U12520 (N_12520,N_11696,N_9674);
xor U12521 (N_12521,N_10215,N_10914);
xor U12522 (N_12522,N_10580,N_10218);
nor U12523 (N_12523,N_9019,N_10590);
nand U12524 (N_12524,N_10937,N_10695);
xor U12525 (N_12525,N_10013,N_10162);
nand U12526 (N_12526,N_9413,N_10024);
and U12527 (N_12527,N_10706,N_10681);
xnor U12528 (N_12528,N_10652,N_9353);
xnor U12529 (N_12529,N_11035,N_10708);
or U12530 (N_12530,N_10145,N_11651);
and U12531 (N_12531,N_11147,N_10931);
nand U12532 (N_12532,N_9309,N_9625);
or U12533 (N_12533,N_9855,N_10738);
nor U12534 (N_12534,N_9975,N_9516);
or U12535 (N_12535,N_9935,N_10154);
nand U12536 (N_12536,N_11589,N_11230);
or U12537 (N_12537,N_10756,N_11578);
nand U12538 (N_12538,N_9409,N_11330);
nand U12539 (N_12539,N_9450,N_10704);
nand U12540 (N_12540,N_11547,N_10131);
xor U12541 (N_12541,N_9244,N_11577);
or U12542 (N_12542,N_11404,N_11362);
and U12543 (N_12543,N_9073,N_11865);
xnor U12544 (N_12544,N_9323,N_9911);
nor U12545 (N_12545,N_9230,N_10774);
and U12546 (N_12546,N_10046,N_11717);
or U12547 (N_12547,N_9906,N_10115);
nand U12548 (N_12548,N_9015,N_10816);
nand U12549 (N_12549,N_10081,N_11621);
nand U12550 (N_12550,N_10986,N_9046);
nand U12551 (N_12551,N_9229,N_10460);
or U12552 (N_12552,N_10376,N_10283);
nand U12553 (N_12553,N_9723,N_10439);
and U12554 (N_12554,N_10449,N_11832);
xor U12555 (N_12555,N_10560,N_11245);
nor U12556 (N_12556,N_9127,N_11545);
or U12557 (N_12557,N_9676,N_9328);
xnor U12558 (N_12558,N_10609,N_10873);
and U12559 (N_12559,N_11823,N_10500);
nand U12560 (N_12560,N_11680,N_10602);
nor U12561 (N_12561,N_11062,N_9211);
and U12562 (N_12562,N_9456,N_9682);
nor U12563 (N_12563,N_11020,N_10814);
or U12564 (N_12564,N_11304,N_9440);
and U12565 (N_12565,N_11190,N_10171);
nor U12566 (N_12566,N_9331,N_10052);
or U12567 (N_12567,N_10507,N_11228);
and U12568 (N_12568,N_9448,N_11073);
or U12569 (N_12569,N_9258,N_11679);
or U12570 (N_12570,N_11149,N_11983);
nand U12571 (N_12571,N_11450,N_10744);
or U12572 (N_12572,N_9327,N_11437);
xnor U12573 (N_12573,N_11018,N_9864);
nor U12574 (N_12574,N_11821,N_11144);
xnor U12575 (N_12575,N_10796,N_11378);
or U12576 (N_12576,N_9509,N_10291);
xor U12577 (N_12577,N_11979,N_9093);
and U12578 (N_12578,N_11749,N_11524);
nand U12579 (N_12579,N_10926,N_9537);
and U12580 (N_12580,N_9434,N_10644);
nor U12581 (N_12581,N_10181,N_10371);
nand U12582 (N_12582,N_11350,N_10268);
or U12583 (N_12583,N_11012,N_9179);
and U12584 (N_12584,N_10813,N_11317);
nor U12585 (N_12585,N_9872,N_11283);
xnor U12586 (N_12586,N_11748,N_10881);
xor U12587 (N_12587,N_10140,N_9524);
nand U12588 (N_12588,N_10167,N_11681);
nor U12589 (N_12589,N_11687,N_10414);
nor U12590 (N_12590,N_11652,N_9389);
nor U12591 (N_12591,N_9843,N_9929);
nor U12592 (N_12592,N_10849,N_10142);
nand U12593 (N_12593,N_9188,N_11080);
or U12594 (N_12594,N_9728,N_10187);
nor U12595 (N_12595,N_9650,N_11536);
and U12596 (N_12596,N_10343,N_9491);
xor U12597 (N_12597,N_11667,N_11082);
nand U12598 (N_12598,N_10107,N_11440);
and U12599 (N_12599,N_11997,N_11766);
nor U12600 (N_12600,N_9411,N_11598);
and U12601 (N_12601,N_11083,N_10745);
or U12602 (N_12602,N_11052,N_11513);
nand U12603 (N_12603,N_10105,N_11506);
or U12604 (N_12604,N_11431,N_10903);
and U12605 (N_12605,N_10338,N_9335);
xnor U12606 (N_12606,N_11834,N_11556);
or U12607 (N_12607,N_11273,N_11937);
nand U12608 (N_12608,N_9251,N_9042);
xnor U12609 (N_12609,N_9930,N_11917);
nand U12610 (N_12610,N_10011,N_10517);
or U12611 (N_12611,N_9820,N_10969);
nand U12612 (N_12612,N_9600,N_10070);
xnor U12613 (N_12613,N_9329,N_9530);
xor U12614 (N_12614,N_10583,N_10747);
or U12615 (N_12615,N_11588,N_9901);
and U12616 (N_12616,N_9239,N_9797);
or U12617 (N_12617,N_10327,N_10444);
xnor U12618 (N_12618,N_9236,N_9063);
nor U12619 (N_12619,N_10534,N_9645);
or U12620 (N_12620,N_11889,N_11707);
and U12621 (N_12621,N_11639,N_10053);
nand U12622 (N_12622,N_9823,N_10492);
xnor U12623 (N_12623,N_11109,N_11898);
and U12624 (N_12624,N_11233,N_10150);
xnor U12625 (N_12625,N_9714,N_11363);
nor U12626 (N_12626,N_11419,N_9483);
and U12627 (N_12627,N_11872,N_9360);
and U12628 (N_12628,N_9362,N_9282);
nor U12629 (N_12629,N_10803,N_10051);
xor U12630 (N_12630,N_9585,N_11838);
nor U12631 (N_12631,N_10503,N_11279);
or U12632 (N_12632,N_9696,N_10772);
or U12633 (N_12633,N_11816,N_10623);
xnor U12634 (N_12634,N_9944,N_10137);
or U12635 (N_12635,N_11005,N_10035);
nand U12636 (N_12636,N_10273,N_10034);
or U12637 (N_12637,N_9091,N_11187);
nor U12638 (N_12638,N_9640,N_11461);
xor U12639 (N_12639,N_11442,N_10196);
xnor U12640 (N_12640,N_11969,N_10298);
nand U12641 (N_12641,N_10927,N_9478);
nand U12642 (N_12642,N_10204,N_10573);
nand U12643 (N_12643,N_10688,N_10485);
nor U12644 (N_12644,N_9939,N_10286);
and U12645 (N_12645,N_9402,N_9037);
nand U12646 (N_12646,N_10794,N_11096);
and U12647 (N_12647,N_10857,N_10683);
nand U12648 (N_12648,N_11934,N_11152);
or U12649 (N_12649,N_11560,N_10040);
xnor U12650 (N_12650,N_10482,N_9131);
nor U12651 (N_12651,N_9862,N_11857);
nor U12652 (N_12652,N_10640,N_10236);
or U12653 (N_12653,N_9934,N_11266);
nor U12654 (N_12654,N_11312,N_10465);
xor U12655 (N_12655,N_10584,N_9512);
nor U12656 (N_12656,N_9802,N_10620);
xnor U12657 (N_12657,N_10516,N_9722);
xor U12658 (N_12658,N_9964,N_11789);
xor U12659 (N_12659,N_9942,N_9666);
nand U12660 (N_12660,N_11288,N_9226);
nand U12661 (N_12661,N_9612,N_10225);
nand U12662 (N_12662,N_10048,N_11841);
nand U12663 (N_12663,N_9449,N_11963);
nand U12664 (N_12664,N_9026,N_11757);
xnor U12665 (N_12665,N_11903,N_9410);
nand U12666 (N_12666,N_9507,N_11436);
xnor U12667 (N_12667,N_10020,N_10996);
nor U12668 (N_12668,N_10212,N_9310);
xnor U12669 (N_12669,N_11664,N_10281);
and U12670 (N_12670,N_10529,N_11590);
nand U12671 (N_12671,N_9059,N_11410);
xor U12672 (N_12672,N_11624,N_10759);
and U12673 (N_12673,N_10546,N_11192);
and U12674 (N_12674,N_10635,N_10068);
nand U12675 (N_12675,N_9754,N_9086);
nand U12676 (N_12676,N_9564,N_9870);
nand U12677 (N_12677,N_11867,N_10452);
nor U12678 (N_12678,N_11017,N_9761);
or U12679 (N_12679,N_11342,N_11351);
xor U12680 (N_12680,N_9277,N_10692);
and U12681 (N_12681,N_9748,N_10842);
nand U12682 (N_12682,N_10836,N_10189);
nand U12683 (N_12683,N_9348,N_9733);
and U12684 (N_12684,N_11281,N_11472);
xnor U12685 (N_12685,N_9569,N_10193);
or U12686 (N_12686,N_11276,N_9529);
nor U12687 (N_12687,N_11635,N_10861);
and U12688 (N_12688,N_10367,N_9325);
or U12689 (N_12689,N_10676,N_11559);
nand U12690 (N_12690,N_10366,N_11075);
nand U12691 (N_12691,N_10504,N_9623);
nand U12692 (N_12692,N_9910,N_9021);
nand U12693 (N_12693,N_10576,N_9163);
or U12694 (N_12694,N_9099,N_11818);
nor U12695 (N_12695,N_10029,N_10116);
nand U12696 (N_12696,N_11671,N_9375);
and U12697 (N_12697,N_11070,N_9242);
and U12698 (N_12698,N_11793,N_9489);
nor U12699 (N_12699,N_11215,N_10866);
xnor U12700 (N_12700,N_9879,N_11332);
and U12701 (N_12701,N_11801,N_9432);
nor U12702 (N_12702,N_11767,N_10975);
or U12703 (N_12703,N_10234,N_11220);
nand U12704 (N_12704,N_10176,N_10207);
nor U12705 (N_12705,N_10445,N_10337);
xor U12706 (N_12706,N_10197,N_10384);
nor U12707 (N_12707,N_10545,N_11134);
or U12708 (N_12708,N_9492,N_9275);
xor U12709 (N_12709,N_10417,N_11047);
nor U12710 (N_12710,N_10852,N_9990);
nor U12711 (N_12711,N_11994,N_11392);
xor U12712 (N_12712,N_9977,N_11221);
nor U12713 (N_12713,N_11851,N_9420);
and U12714 (N_12714,N_10195,N_10689);
nor U12715 (N_12715,N_11938,N_9371);
nor U12716 (N_12716,N_9871,N_10742);
xor U12717 (N_12717,N_11125,N_11799);
or U12718 (N_12718,N_11065,N_11942);
and U12719 (N_12719,N_11975,N_11158);
and U12720 (N_12720,N_9280,N_9697);
nor U12721 (N_12721,N_11949,N_10895);
and U12722 (N_12722,N_11366,N_10315);
nor U12723 (N_12723,N_9663,N_9192);
nand U12724 (N_12724,N_11722,N_9690);
nand U12725 (N_12725,N_10025,N_10522);
and U12726 (N_12726,N_11259,N_9171);
nor U12727 (N_12727,N_11850,N_9810);
nor U12728 (N_12728,N_11019,N_11812);
or U12729 (N_12729,N_11956,N_9540);
and U12730 (N_12730,N_10027,N_11303);
or U12731 (N_12731,N_10135,N_10923);
xnor U12732 (N_12732,N_10381,N_9262);
or U12733 (N_12733,N_11633,N_11768);
or U12734 (N_12734,N_9357,N_10078);
and U12735 (N_12735,N_10172,N_11945);
nor U12736 (N_12736,N_10977,N_11423);
xnor U12737 (N_12737,N_11806,N_11397);
nand U12738 (N_12738,N_11553,N_9652);
and U12739 (N_12739,N_11191,N_10288);
and U12740 (N_12740,N_10341,N_10106);
xnor U12741 (N_12741,N_9427,N_10330);
nor U12742 (N_12742,N_9034,N_9266);
xor U12743 (N_12743,N_9000,N_11719);
or U12744 (N_12744,N_10917,N_10365);
or U12745 (N_12745,N_10443,N_9496);
nor U12746 (N_12746,N_11209,N_11991);
or U12747 (N_12747,N_10944,N_11097);
or U12748 (N_12748,N_11692,N_9615);
or U12749 (N_12749,N_9205,N_10279);
xnor U12750 (N_12750,N_11031,N_11138);
nor U12751 (N_12751,N_10373,N_11765);
nor U12752 (N_12752,N_9435,N_9902);
or U12753 (N_12753,N_9095,N_11290);
or U12754 (N_12754,N_9064,N_9079);
and U12755 (N_12755,N_10511,N_11750);
or U12756 (N_12756,N_9421,N_9888);
nand U12757 (N_12757,N_10829,N_10276);
nand U12758 (N_12758,N_9165,N_11514);
or U12759 (N_12759,N_10877,N_9832);
or U12760 (N_12760,N_10392,N_10841);
and U12761 (N_12761,N_9322,N_9108);
nand U12762 (N_12762,N_10638,N_10537);
nor U12763 (N_12763,N_9318,N_9088);
and U12764 (N_12764,N_9292,N_11746);
nand U12765 (N_12765,N_10163,N_9283);
xor U12766 (N_12766,N_11256,N_11897);
nand U12767 (N_12767,N_11301,N_9525);
nand U12768 (N_12768,N_10252,N_10165);
xor U12769 (N_12769,N_10132,N_10731);
nand U12770 (N_12770,N_11234,N_10655);
and U12771 (N_12771,N_10209,N_11167);
or U12772 (N_12772,N_10457,N_10678);
nand U12773 (N_12773,N_9129,N_9397);
or U12774 (N_12774,N_10486,N_9203);
nand U12775 (N_12775,N_10886,N_10428);
nor U12776 (N_12776,N_10463,N_11550);
and U12777 (N_12777,N_10657,N_10270);
nand U12778 (N_12778,N_10768,N_11180);
or U12779 (N_12779,N_11843,N_9462);
xor U12780 (N_12780,N_10022,N_11214);
nand U12781 (N_12781,N_10191,N_10659);
nor U12782 (N_12782,N_9190,N_11519);
nor U12783 (N_12783,N_9912,N_11137);
nor U12784 (N_12784,N_9951,N_9534);
nand U12785 (N_12785,N_11173,N_9233);
nand U12786 (N_12786,N_9636,N_11405);
xor U12787 (N_12787,N_9180,N_10804);
nand U12788 (N_12788,N_9210,N_11101);
nor U12789 (N_12789,N_11594,N_11172);
and U12790 (N_12790,N_10818,N_11003);
nor U12791 (N_12791,N_11401,N_11381);
nand U12792 (N_12792,N_11354,N_9043);
nand U12793 (N_12793,N_11000,N_10254);
xor U12794 (N_12794,N_10031,N_9848);
or U12795 (N_12795,N_9351,N_9763);
or U12796 (N_12796,N_9661,N_11520);
xor U12797 (N_12797,N_11709,N_9146);
xnor U12798 (N_12798,N_11853,N_10325);
xnor U12799 (N_12799,N_11775,N_9157);
nor U12800 (N_12800,N_9893,N_10586);
or U12801 (N_12801,N_10055,N_9866);
nand U12802 (N_12802,N_10755,N_11329);
or U12803 (N_12803,N_11990,N_11830);
nor U12804 (N_12804,N_11493,N_11809);
xnor U12805 (N_12805,N_10184,N_10032);
and U12806 (N_12806,N_10049,N_10649);
xnor U12807 (N_12807,N_11601,N_9288);
xnor U12808 (N_12808,N_9614,N_9057);
or U12809 (N_12809,N_11391,N_10515);
xnor U12810 (N_12810,N_9793,N_11189);
nor U12811 (N_12811,N_10113,N_10319);
xnor U12812 (N_12812,N_9463,N_11026);
and U12813 (N_12813,N_10152,N_9760);
or U12814 (N_12814,N_11504,N_9730);
xnor U12815 (N_12815,N_9815,N_11641);
xor U12816 (N_12816,N_9377,N_9732);
nand U12817 (N_12817,N_10801,N_9995);
nand U12818 (N_12818,N_10614,N_11479);
xor U12819 (N_12819,N_11310,N_11356);
nor U12820 (N_12820,N_9120,N_11425);
nor U12821 (N_12821,N_11721,N_10734);
or U12822 (N_12822,N_9051,N_9359);
or U12823 (N_12823,N_10898,N_9159);
nand U12824 (N_12824,N_9164,N_9753);
xnor U12825 (N_12825,N_11413,N_10037);
or U12826 (N_12826,N_11491,N_10217);
or U12827 (N_12827,N_10981,N_10642);
nand U12828 (N_12828,N_11307,N_10003);
nor U12829 (N_12829,N_10752,N_10524);
nor U12830 (N_12830,N_9654,N_9151);
or U12831 (N_12831,N_11920,N_11893);
nand U12832 (N_12832,N_11913,N_10481);
nand U12833 (N_12833,N_9136,N_11540);
or U12834 (N_12834,N_9356,N_9094);
nor U12835 (N_12835,N_9405,N_11675);
nor U12836 (N_12836,N_9071,N_9812);
nand U12837 (N_12837,N_11071,N_11434);
xor U12838 (N_12838,N_9224,N_10368);
or U12839 (N_12839,N_11114,N_9027);
xnor U12840 (N_12840,N_11534,N_10519);
xnor U12841 (N_12841,N_11008,N_9926);
or U12842 (N_12842,N_9894,N_9603);
xor U12843 (N_12843,N_10832,N_11745);
and U12844 (N_12844,N_9361,N_10219);
and U12845 (N_12845,N_9112,N_11458);
xor U12846 (N_12846,N_9550,N_10407);
and U12847 (N_12847,N_11141,N_10765);
or U12848 (N_12848,N_11747,N_10625);
xor U12849 (N_12849,N_11999,N_11059);
nand U12850 (N_12850,N_11977,N_9581);
and U12851 (N_12851,N_9655,N_9514);
or U12852 (N_12852,N_9052,N_9330);
xnor U12853 (N_12853,N_9096,N_11320);
and U12854 (N_12854,N_9394,N_11627);
nand U12855 (N_12855,N_11286,N_9799);
nor U12856 (N_12856,N_11352,N_10019);
or U12857 (N_12857,N_11455,N_9554);
xnor U12858 (N_12858,N_11518,N_10974);
nor U12859 (N_12859,N_9989,N_9379);
or U12860 (N_12860,N_10863,N_10901);
nor U12861 (N_12861,N_9243,N_11596);
nor U12862 (N_12862,N_11638,N_9166);
nand U12863 (N_12863,N_9957,N_11689);
or U12864 (N_12864,N_11260,N_11972);
nand U12865 (N_12865,N_11879,N_9431);
nor U12866 (N_12866,N_9541,N_10815);
xor U12867 (N_12867,N_11654,N_11663);
or U12868 (N_12868,N_11882,N_9363);
nor U12869 (N_12869,N_10419,N_9393);
nand U12870 (N_12870,N_11608,N_11251);
and U12871 (N_12871,N_10727,N_10188);
and U12872 (N_12872,N_11648,N_11118);
or U12873 (N_12873,N_11703,N_10631);
nor U12874 (N_12874,N_10820,N_11375);
nand U12875 (N_12875,N_11542,N_10447);
nor U12876 (N_12876,N_10361,N_10348);
nand U12877 (N_12877,N_9553,N_9535);
and U12878 (N_12878,N_10086,N_11927);
and U12879 (N_12879,N_11595,N_9807);
nand U12880 (N_12880,N_10718,N_10099);
xnor U12881 (N_12881,N_9407,N_9777);
or U12882 (N_12882,N_11976,N_10075);
or U12883 (N_12883,N_9572,N_10634);
or U12884 (N_12884,N_9882,N_9298);
nor U12885 (N_12885,N_10567,N_11380);
or U12886 (N_12886,N_10069,N_10258);
and U12887 (N_12887,N_10582,N_10979);
nor U12888 (N_12888,N_11845,N_11786);
nor U12889 (N_12889,N_10790,N_10748);
xor U12890 (N_12890,N_9466,N_11820);
and U12891 (N_12891,N_10889,N_9297);
or U12892 (N_12892,N_9089,N_11699);
nor U12893 (N_12893,N_9596,N_10715);
xnor U12894 (N_12894,N_11474,N_10495);
nand U12895 (N_12895,N_11629,N_11970);
nand U12896 (N_12896,N_9589,N_9857);
nor U12897 (N_12897,N_9191,N_10947);
xor U12898 (N_12898,N_11123,N_9228);
xnor U12899 (N_12899,N_11241,N_9137);
and U12900 (N_12900,N_11486,N_9482);
or U12901 (N_12901,N_9694,N_9937);
nand U12902 (N_12902,N_11327,N_10983);
xnor U12903 (N_12903,N_10505,N_10404);
and U12904 (N_12904,N_9824,N_9341);
nor U12905 (N_12905,N_11525,N_9932);
and U12906 (N_12906,N_9041,N_11121);
or U12907 (N_12907,N_11769,N_11503);
nand U12908 (N_12908,N_9956,N_10314);
or U12909 (N_12909,N_11077,N_9792);
or U12910 (N_12910,N_9671,N_11028);
xnor U12911 (N_12911,N_9928,N_11728);
or U12912 (N_12912,N_11422,N_9090);
or U12913 (N_12913,N_9688,N_9687);
nor U12914 (N_12914,N_10079,N_10249);
nor U12915 (N_12915,N_9933,N_9084);
xnor U12916 (N_12916,N_11819,N_11885);
nand U12917 (N_12917,N_9035,N_9692);
or U12918 (N_12918,N_9963,N_10945);
xor U12919 (N_12919,N_10329,N_9776);
and U12920 (N_12920,N_10578,N_9012);
nor U12921 (N_12921,N_11562,N_9208);
or U12922 (N_12922,N_10429,N_11896);
and U12923 (N_12923,N_10415,N_9148);
nand U12924 (N_12924,N_10108,N_11535);
and U12925 (N_12925,N_9354,N_10267);
or U12926 (N_12926,N_11755,N_10073);
nor U12927 (N_12927,N_10760,N_10594);
nor U12928 (N_12928,N_10561,N_9415);
nand U12929 (N_12929,N_9447,N_10396);
nor U12930 (N_12930,N_9877,N_9343);
xor U12931 (N_12931,N_9391,N_10920);
nor U12932 (N_12932,N_10799,N_9775);
nor U12933 (N_12933,N_11665,N_11901);
or U12934 (N_12934,N_11412,N_10112);
or U12935 (N_12935,N_11132,N_10213);
nor U12936 (N_12936,N_9404,N_11948);
nor U12937 (N_12937,N_11933,N_9488);
nor U12938 (N_12938,N_11758,N_11718);
nor U12939 (N_12939,N_10346,N_10382);
or U12940 (N_12940,N_11908,N_11421);
xnor U12941 (N_12941,N_11599,N_9693);
xnor U12942 (N_12942,N_11318,N_10421);
nand U12943 (N_12943,N_9364,N_11626);
or U12944 (N_12944,N_10344,N_10023);
or U12945 (N_12945,N_10777,N_10156);
or U12946 (N_12946,N_9285,N_10946);
or U12947 (N_12947,N_10707,N_9745);
nand U12948 (N_12948,N_10432,N_10606);
and U12949 (N_12949,N_9237,N_10395);
xor U12950 (N_12950,N_9006,N_9586);
nand U12951 (N_12951,N_9961,N_9853);
nor U12952 (N_12952,N_10702,N_9366);
or U12953 (N_12953,N_11015,N_11364);
nor U12954 (N_12954,N_11895,N_9526);
and U12955 (N_12955,N_11886,N_10262);
nand U12956 (N_12956,N_10067,N_11271);
nor U12957 (N_12957,N_10539,N_10520);
nand U12958 (N_12958,N_11712,N_10089);
nor U12959 (N_12959,N_11840,N_10380);
xor U12960 (N_12960,N_10265,N_11257);
and U12961 (N_12961,N_9265,N_9892);
nor U12962 (N_12962,N_11741,N_9387);
or U12963 (N_12963,N_9836,N_9045);
xnor U12964 (N_12964,N_9830,N_10826);
or U12965 (N_12965,N_11754,N_10450);
xnor U12966 (N_12966,N_11016,N_9425);
xnor U12967 (N_12967,N_11095,N_9649);
or U12968 (N_12968,N_9700,N_11162);
xnor U12969 (N_12969,N_11449,N_11495);
xnor U12970 (N_12970,N_10374,N_10906);
nand U12971 (N_12971,N_9850,N_11509);
and U12972 (N_12972,N_11716,N_9486);
xor U12973 (N_12973,N_11695,N_11112);
nor U12974 (N_12974,N_9014,N_10934);
nor U12975 (N_12975,N_10462,N_11145);
nor U12976 (N_12976,N_9657,N_9669);
nor U12977 (N_12977,N_9982,N_11453);
nor U12978 (N_12978,N_11771,N_11911);
nand U12979 (N_12979,N_11447,N_11231);
and U12980 (N_12980,N_11004,N_11593);
and U12981 (N_12981,N_11325,N_10253);
and U12982 (N_12982,N_11538,N_9717);
and U12983 (N_12983,N_10316,N_11725);
or U12984 (N_12984,N_9319,N_10553);
and U12985 (N_12985,N_9075,N_10300);
nor U12986 (N_12986,N_9412,N_11622);
or U12987 (N_12987,N_11113,N_11268);
or U12988 (N_12988,N_11186,N_9573);
and U12989 (N_12989,N_11253,N_9383);
or U12990 (N_12990,N_11828,N_11852);
and U12991 (N_12991,N_9367,N_10948);
nand U12992 (N_12992,N_9113,N_10865);
nand U12993 (N_12993,N_11592,N_9588);
xnor U12994 (N_12994,N_9887,N_11697);
xor U12995 (N_12995,N_10780,N_11961);
and U12996 (N_12996,N_10936,N_10007);
nor U12997 (N_12997,N_9475,N_10933);
nor U12998 (N_12998,N_10932,N_10130);
and U12999 (N_12999,N_10328,N_10883);
nor U13000 (N_13000,N_11337,N_10675);
or U13001 (N_13001,N_11888,N_10264);
and U13002 (N_13002,N_11959,N_11063);
nor U13003 (N_13003,N_9631,N_9997);
nand U13004 (N_13004,N_11357,N_10459);
and U13005 (N_13005,N_10238,N_11043);
nand U13006 (N_13006,N_9193,N_11494);
and U13007 (N_13007,N_9575,N_11690);
and U13008 (N_13008,N_11875,N_9048);
nor U13009 (N_13009,N_10993,N_10878);
nor U13010 (N_13010,N_10800,N_10592);
xor U13011 (N_13011,N_9859,N_11759);
and U13012 (N_13012,N_10455,N_10709);
xnor U13013 (N_13013,N_9030,N_10226);
xnor U13014 (N_13014,N_10260,N_9066);
nand U13015 (N_13015,N_9007,N_10157);
nor U13016 (N_13016,N_11086,N_10810);
nor U13017 (N_13017,N_10257,N_11226);
nand U13018 (N_13018,N_10521,N_10012);
and U13019 (N_13019,N_10628,N_9119);
nand U13020 (N_13020,N_10263,N_9734);
or U13021 (N_13021,N_11914,N_11904);
and U13022 (N_13022,N_9100,N_9519);
xor U13023 (N_13023,N_10615,N_10228);
nand U13024 (N_13024,N_9852,N_11798);
nand U13025 (N_13025,N_11115,N_11574);
or U13026 (N_13026,N_10464,N_9918);
and U13027 (N_13027,N_9747,N_11711);
nand U13028 (N_13028,N_9974,N_11196);
nor U13029 (N_13029,N_9595,N_10426);
and U13030 (N_13030,N_10438,N_9865);
nand U13031 (N_13031,N_9634,N_9499);
nand U13032 (N_13032,N_10136,N_11388);
nor U13033 (N_13033,N_11862,N_10544);
nor U13034 (N_13034,N_11361,N_9683);
nor U13035 (N_13035,N_11569,N_9837);
and U13036 (N_13036,N_11306,N_10017);
or U13037 (N_13037,N_10149,N_10879);
nor U13038 (N_13038,N_11674,N_11912);
or U13039 (N_13039,N_10155,N_11210);
or U13040 (N_13040,N_11242,N_10513);
and U13041 (N_13041,N_9503,N_9194);
nand U13042 (N_13042,N_11760,N_11292);
nand U13043 (N_13043,N_9303,N_10767);
nand U13044 (N_13044,N_10077,N_9209);
and U13045 (N_13045,N_10956,N_9881);
and U13046 (N_13046,N_9494,N_10103);
and U13047 (N_13047,N_11034,N_11029);
xnor U13048 (N_13048,N_10506,N_9392);
nor U13049 (N_13049,N_11106,N_9255);
nand U13050 (N_13050,N_11373,N_11032);
and U13051 (N_13051,N_10894,N_10334);
nand U13052 (N_13052,N_11261,N_10232);
nand U13053 (N_13053,N_10976,N_9543);
nor U13054 (N_13054,N_10496,N_11591);
xnor U13055 (N_13055,N_9970,N_11476);
nand U13056 (N_13056,N_9597,N_11212);
and U13057 (N_13057,N_10248,N_11182);
xor U13058 (N_13058,N_10224,N_9495);
nor U13059 (N_13059,N_11408,N_11058);
or U13060 (N_13060,N_10670,N_9523);
nand U13061 (N_13061,N_10997,N_11980);
nor U13062 (N_13062,N_9660,N_10812);
xnor U13063 (N_13063,N_9133,N_9817);
or U13064 (N_13064,N_9875,N_10884);
nand U13065 (N_13065,N_11539,N_11011);
and U13066 (N_13066,N_11612,N_9500);
nand U13067 (N_13067,N_10185,N_9897);
nand U13068 (N_13068,N_10347,N_10311);
xnor U13069 (N_13069,N_11814,N_10720);
or U13070 (N_13070,N_9423,N_11660);
xnor U13071 (N_13071,N_10058,N_10962);
nand U13072 (N_13072,N_9899,N_9317);
xor U13073 (N_13073,N_11469,N_11379);
and U13074 (N_13074,N_10758,N_11713);
or U13075 (N_13075,N_11122,N_10509);
or U13076 (N_13076,N_10057,N_10308);
nor U13077 (N_13077,N_10060,N_9973);
nand U13078 (N_13078,N_11795,N_9966);
and U13079 (N_13079,N_9080,N_11670);
or U13080 (N_13080,N_10789,N_10554);
or U13081 (N_13081,N_11817,N_10008);
and U13082 (N_13082,N_10223,N_9861);
nor U13083 (N_13083,N_9220,N_10653);
nor U13084 (N_13084,N_11763,N_9784);
nand U13085 (N_13085,N_9445,N_11407);
nand U13086 (N_13086,N_9290,N_9863);
and U13087 (N_13087,N_10239,N_10110);
and U13088 (N_13088,N_10677,N_10494);
nand U13089 (N_13089,N_9774,N_10699);
nor U13090 (N_13090,N_10143,N_10002);
xor U13091 (N_13091,N_9883,N_9617);
and U13092 (N_13092,N_9938,N_10102);
xnor U13093 (N_13093,N_9477,N_10109);
or U13094 (N_13094,N_9340,N_11815);
nand U13095 (N_13095,N_10458,N_9611);
or U13096 (N_13096,N_11958,N_9609);
and U13097 (N_13097,N_9779,N_9104);
xnor U13098 (N_13098,N_10569,N_10179);
nand U13099 (N_13099,N_11353,N_10408);
and U13100 (N_13100,N_11762,N_10867);
nor U13101 (N_13101,N_11470,N_9958);
nor U13102 (N_13102,N_9672,N_10080);
xnor U13103 (N_13103,N_9141,N_11100);
or U13104 (N_13104,N_9473,N_9273);
and U13105 (N_13105,N_10498,N_11349);
nand U13106 (N_13106,N_9578,N_10269);
nand U13107 (N_13107,N_11321,N_9291);
or U13108 (N_13108,N_11157,N_11935);
xor U13109 (N_13109,N_9036,N_11993);
nor U13110 (N_13110,N_11669,N_11794);
and U13111 (N_13111,N_9936,N_9241);
and U13112 (N_13112,N_10599,N_11926);
xor U13113 (N_13113,N_9739,N_11081);
xor U13114 (N_13114,N_9395,N_11673);
and U13115 (N_13115,N_10118,N_11615);
nor U13116 (N_13116,N_10672,N_10050);
xor U13117 (N_13117,N_10161,N_11444);
and U13118 (N_13118,N_9972,N_11150);
nor U13119 (N_13119,N_9055,N_11238);
nand U13120 (N_13120,N_9253,N_11237);
and U13121 (N_13121,N_9983,N_9067);
and U13122 (N_13122,N_11042,N_9437);
nor U13123 (N_13123,N_11551,N_11724);
nor U13124 (N_13124,N_11634,N_10098);
and U13125 (N_13125,N_10045,N_10703);
xnor U13126 (N_13126,N_9673,N_11403);
xor U13127 (N_13127,N_10423,N_11484);
nand U13128 (N_13128,N_11439,N_11783);
nor U13129 (N_13129,N_9132,N_9555);
nand U13130 (N_13130,N_11910,N_11454);
nor U13131 (N_13131,N_10955,N_9827);
nand U13132 (N_13132,N_11174,N_9574);
and U13133 (N_13133,N_9948,N_10880);
nor U13134 (N_13134,N_10411,N_11105);
nand U13135 (N_13135,N_10336,N_9841);
xnor U13136 (N_13136,N_9962,N_10972);
nand U13137 (N_13137,N_11714,N_10959);
nor U13138 (N_13138,N_10208,N_9287);
nand U13139 (N_13139,N_9826,N_10953);
nand U13140 (N_13140,N_11199,N_11358);
or U13141 (N_13141,N_11480,N_10551);
xor U13142 (N_13142,N_11871,N_9868);
xnor U13143 (N_13143,N_10295,N_10461);
xor U13144 (N_13144,N_9268,N_11659);
xor U13145 (N_13145,N_11387,N_10710);
nor U13146 (N_13146,N_10741,N_11202);
nand U13147 (N_13147,N_11227,N_11922);
or U13148 (N_13148,N_11614,N_10378);
nand U13149 (N_13149,N_9498,N_11515);
nand U13150 (N_13150,N_9771,N_9474);
xnor U13151 (N_13151,N_9458,N_9724);
xnor U13152 (N_13152,N_10119,N_9480);
and U13153 (N_13153,N_11001,N_10771);
nand U13154 (N_13154,N_10556,N_11232);
nand U13155 (N_13155,N_11103,N_11284);
xor U13156 (N_13156,N_9153,N_11772);
and U13157 (N_13157,N_9905,N_9546);
or U13158 (N_13158,N_11007,N_10016);
or U13159 (N_13159,N_11313,N_11027);
or U13160 (N_13160,N_11584,N_10088);
or U13161 (N_13161,N_10128,N_10230);
nand U13162 (N_13162,N_10375,N_9835);
xnor U13163 (N_13163,N_11955,N_9709);
nand U13164 (N_13164,N_10918,N_11296);
nand U13165 (N_13165,N_11069,N_11544);
or U13166 (N_13166,N_11943,N_10028);
or U13167 (N_13167,N_11946,N_9946);
and U13168 (N_13168,N_11797,N_9662);
nor U13169 (N_13169,N_11389,N_11964);
and U13170 (N_13170,N_11602,N_11163);
xor U13171 (N_13171,N_9593,N_9349);
nor U13172 (N_13172,N_11899,N_10318);
nor U13173 (N_13173,N_10668,N_10535);
nand U13174 (N_13174,N_10792,N_9592);
nor U13175 (N_13175,N_9786,N_10297);
nand U13176 (N_13176,N_10190,N_10645);
and U13177 (N_13177,N_11866,N_10183);
and U13178 (N_13178,N_9952,N_9549);
nor U13179 (N_13179,N_11788,N_9204);
nand U13180 (N_13180,N_11743,N_11778);
nor U13181 (N_13181,N_9805,N_11406);
nor U13182 (N_13182,N_9352,N_10471);
or U13183 (N_13183,N_11869,N_11764);
nand U13184 (N_13184,N_9689,N_10446);
nor U13185 (N_13185,N_11984,N_11084);
xor U13186 (N_13186,N_10379,N_10961);
or U13187 (N_13187,N_11085,N_11735);
or U13188 (N_13188,N_10434,N_10998);
nor U13189 (N_13189,N_10851,N_10821);
or U13190 (N_13190,N_11177,N_10605);
and U13191 (N_13191,N_11881,N_11616);
nand U13192 (N_13192,N_9994,N_9175);
and U13193 (N_13193,N_11333,N_11417);
or U13194 (N_13194,N_9598,N_11572);
xnor U13195 (N_13195,N_11576,N_9376);
or U13196 (N_13196,N_10762,N_11500);
nand U13197 (N_13197,N_10843,N_9446);
xnor U13198 (N_13198,N_11206,N_9270);
xnor U13199 (N_13199,N_11971,N_10572);
and U13200 (N_13200,N_9368,N_11966);
nand U13201 (N_13201,N_10151,N_10905);
xor U13202 (N_13202,N_10830,N_9742);
or U13203 (N_13203,N_10621,N_10954);
nor U13204 (N_13204,N_11328,N_10951);
or U13205 (N_13205,N_9895,N_11014);
nor U13206 (N_13206,N_11736,N_10497);
or U13207 (N_13207,N_9570,N_11252);
nand U13208 (N_13208,N_9470,N_10499);
nand U13209 (N_13209,N_9123,N_9566);
nand U13210 (N_13210,N_11661,N_10793);
or U13211 (N_13211,N_11204,N_9286);
nor U13212 (N_13212,N_10358,N_11825);
and U13213 (N_13213,N_11298,N_11036);
xor U13214 (N_13214,N_11907,N_10383);
nor U13215 (N_13215,N_11446,N_10541);
nand U13216 (N_13216,N_11466,N_11462);
or U13217 (N_13217,N_10317,N_9320);
nand U13218 (N_13218,N_10490,N_10321);
nor U13219 (N_13219,N_11836,N_11522);
nor U13220 (N_13220,N_9479,N_9160);
nand U13221 (N_13221,N_9261,N_11691);
xor U13222 (N_13222,N_10619,N_11894);
or U13223 (N_13223,N_11678,N_11179);
xnor U13224 (N_13224,N_10825,N_11161);
nor U13225 (N_13225,N_9168,N_11668);
and U13226 (N_13226,N_11040,N_11377);
or U13227 (N_13227,N_10531,N_10550);
xnor U13228 (N_13228,N_10420,N_11701);
nand U13229 (N_13229,N_9627,N_10871);
xor U13230 (N_13230,N_10604,N_10968);
xor U13231 (N_13231,N_11941,N_10597);
xor U13232 (N_13232,N_10725,N_11582);
nor U13233 (N_13233,N_11207,N_11369);
nor U13234 (N_13234,N_10202,N_9138);
and U13235 (N_13235,N_10662,N_10807);
nor U13236 (N_13236,N_11386,N_10740);
nand U13237 (N_13237,N_10571,N_10354);
xnor U13238 (N_13238,N_11887,N_10935);
nor U13239 (N_13239,N_10390,N_9813);
nor U13240 (N_13240,N_10915,N_9344);
xnor U13241 (N_13241,N_9720,N_10412);
nor U13242 (N_13242,N_11244,N_9107);
nor U13243 (N_13243,N_10047,N_10973);
xor U13244 (N_13244,N_10627,N_10966);
nor U13245 (N_13245,N_9186,N_9691);
and U13246 (N_13246,N_9337,N_9858);
and U13247 (N_13247,N_11200,N_11395);
or U13248 (N_13248,N_11487,N_11299);
nand U13249 (N_13249,N_9467,N_11374);
nor U13250 (N_13250,N_9891,N_11640);
xor U13251 (N_13251,N_9706,N_9969);
xnor U13252 (N_13252,N_10730,N_9819);
or U13253 (N_13253,N_11587,N_11060);
nor U13254 (N_13254,N_11527,N_11563);
or U13255 (N_13255,N_9313,N_10502);
nand U13256 (N_13256,N_9677,N_10266);
nand U13257 (N_13257,N_9651,N_11119);
nor U13258 (N_13258,N_10660,N_10469);
nor U13259 (N_13259,N_10203,N_9571);
and U13260 (N_13260,N_11731,N_10806);
xnor U13261 (N_13261,N_11657,N_11537);
nor U13262 (N_13262,N_9465,N_9040);
and U13263 (N_13263,N_11133,N_11649);
nand U13264 (N_13264,N_9710,N_11175);
or U13265 (N_13265,N_10307,N_9025);
or U13266 (N_13266,N_9839,N_11297);
nor U13267 (N_13267,N_10887,N_10651);
and U13268 (N_13268,N_10839,N_10663);
or U13269 (N_13269,N_9740,N_10980);
nand U13270 (N_13270,N_10896,N_11790);
nand U13271 (N_13271,N_10287,N_9924);
nand U13272 (N_13272,N_10769,N_10809);
or U13273 (N_13273,N_10097,N_11996);
nand U13274 (N_13274,N_10897,N_9017);
or U13275 (N_13275,N_10693,N_11049);
xnor U13276 (N_13276,N_11094,N_11732);
nand U13277 (N_13277,N_11981,N_11382);
xnor U13278 (N_13278,N_10994,N_9752);
and U13279 (N_13279,N_10147,N_9789);
or U13280 (N_13280,N_10451,N_10292);
and U13281 (N_13281,N_9874,N_11876);
and U13282 (N_13282,N_9931,N_10174);
nor U13283 (N_13283,N_10958,N_10391);
xor U13284 (N_13284,N_9076,N_11723);
or U13285 (N_13285,N_10312,N_10134);
nor U13286 (N_13286,N_10472,N_9106);
nor U13287 (N_13287,N_9943,N_10658);
and U13288 (N_13288,N_11250,N_11729);
and U13289 (N_13289,N_9846,N_11170);
or U13290 (N_13290,N_11218,N_10540);
nand U13291 (N_13291,N_9999,N_9301);
and U13292 (N_13292,N_11618,N_9791);
nand U13293 (N_13293,N_9960,N_10294);
xnor U13294 (N_13294,N_10085,N_10004);
nand U13295 (N_13295,N_10555,N_10448);
xor U13296 (N_13296,N_10697,N_11441);
and U13297 (N_13297,N_11213,N_11055);
or U13298 (N_13298,N_10369,N_10869);
or U13299 (N_13299,N_10010,N_9814);
xor U13300 (N_13300,N_9996,N_9016);
or U13301 (N_13301,N_9183,N_9646);
and U13302 (N_13302,N_10211,N_9162);
and U13303 (N_13303,N_10091,N_10240);
and U13304 (N_13304,N_11950,N_11849);
xor U13305 (N_13305,N_9460,N_10066);
xnor U13306 (N_13306,N_10950,N_9860);
and U13307 (N_13307,N_10885,N_9621);
xor U13308 (N_13308,N_9481,N_10409);
nor U13309 (N_13309,N_11883,N_10577);
xnor U13310 (N_13310,N_10930,N_10680);
nand U13311 (N_13311,N_10009,N_9044);
or U13312 (N_13312,N_11925,N_9967);
nor U13313 (N_13313,N_9751,N_11802);
xnor U13314 (N_13314,N_11928,N_10274);
nand U13315 (N_13315,N_11978,N_9406);
or U13316 (N_13316,N_9245,N_11906);
xor U13317 (N_13317,N_10786,N_10717);
or U13318 (N_13318,N_9247,N_9559);
xor U13319 (N_13319,N_11465,N_10339);
and U13320 (N_13320,N_11617,N_11646);
xnor U13321 (N_13321,N_9314,N_10589);
and U13322 (N_13322,N_11686,N_10530);
nor U13323 (N_13323,N_11915,N_10868);
xor U13324 (N_13324,N_10750,N_11478);
and U13325 (N_13325,N_9822,N_11201);
nand U13326 (N_13326,N_10483,N_11631);
or U13327 (N_13327,N_9539,N_10302);
xnor U13328 (N_13328,N_9538,N_9250);
and U13329 (N_13329,N_9296,N_9626);
and U13330 (N_13330,N_11932,N_10222);
nor U13331 (N_13331,N_11808,N_11710);
or U13332 (N_13332,N_9130,N_11488);
nor U13333 (N_13333,N_11947,N_11954);
nor U13334 (N_13334,N_10310,N_10562);
xor U13335 (N_13335,N_11939,N_10855);
or U13336 (N_13336,N_10563,N_10301);
or U13337 (N_13337,N_11842,N_11953);
nand U13338 (N_13338,N_11813,N_9685);
and U13339 (N_13339,N_10565,N_9968);
and U13340 (N_13340,N_10043,N_10705);
or U13341 (N_13341,N_9177,N_9305);
xnor U13342 (N_13342,N_11131,N_9632);
nor U13343 (N_13343,N_9149,N_10320);
nor U13344 (N_13344,N_9271,N_9124);
xnor U13345 (N_13345,N_9472,N_10100);
and U13346 (N_13346,N_11974,N_11090);
nand U13347 (N_13347,N_11666,N_11393);
xnor U13348 (N_13348,N_9772,N_11120);
or U13349 (N_13349,N_11720,N_10776);
and U13350 (N_13350,N_9418,N_9502);
and U13351 (N_13351,N_11475,N_10427);
or U13352 (N_13352,N_9668,N_9049);
nand U13353 (N_13353,N_10661,N_11751);
nor U13354 (N_13354,N_10665,N_11076);
or U13355 (N_13355,N_11548,N_11420);
nor U13356 (N_13356,N_10984,N_10736);
xor U13357 (N_13357,N_11730,N_10629);
nor U13358 (N_13358,N_10690,N_11452);
xnor U13359 (N_13359,N_9637,N_11921);
nand U13360 (N_13360,N_10304,N_11324);
or U13361 (N_13361,N_9408,N_10733);
and U13362 (N_13362,N_10466,N_11523);
or U13363 (N_13363,N_11650,N_11193);
nor U13364 (N_13364,N_11785,N_11359);
nor U13365 (N_13365,N_9332,N_9284);
nand U13366 (N_13366,N_10566,N_11512);
nand U13367 (N_13367,N_9139,N_10214);
nand U13368 (N_13368,N_9536,N_11285);
nand U13369 (N_13369,N_10044,N_9240);
nor U13370 (N_13370,N_9916,N_11859);
nand U13371 (N_13371,N_9115,N_11135);
nand U13372 (N_13372,N_11104,N_11188);
or U13373 (N_13373,N_11160,N_9840);
nand U13374 (N_13374,N_10397,N_9886);
or U13375 (N_13375,N_9778,N_11464);
xor U13376 (N_13376,N_9316,N_9248);
nand U13377 (N_13377,N_9716,N_10732);
and U13378 (N_13378,N_10538,N_10370);
xnor U13379 (N_13379,N_9276,N_10277);
and U13380 (N_13380,N_9986,N_11316);
nand U13381 (N_13381,N_10340,N_10581);
and U13382 (N_13382,N_9142,N_9908);
xor U13383 (N_13383,N_10074,N_11067);
or U13384 (N_13384,N_11278,N_9531);
or U13385 (N_13385,N_10533,N_11262);
nand U13386 (N_13386,N_9396,N_10056);
or U13387 (N_13387,N_11275,N_9873);
nor U13388 (N_13388,N_9312,N_11396);
nand U13389 (N_13389,N_11586,N_11319);
nand U13390 (N_13390,N_10987,N_9218);
nand U13391 (N_13391,N_9658,N_11341);
xor U13392 (N_13392,N_9459,N_9370);
nand U13393 (N_13393,N_9172,N_11630);
xor U13394 (N_13394,N_11402,N_11143);
and U13395 (N_13395,N_9557,N_9527);
nor U13396 (N_13396,N_9493,N_9020);
or U13397 (N_13397,N_9451,N_9490);
nor U13398 (N_13398,N_10922,N_9355);
nand U13399 (N_13399,N_10430,N_9103);
nor U13400 (N_13400,N_10406,N_9485);
nor U13401 (N_13401,N_10967,N_10335);
nor U13402 (N_13402,N_10711,N_10616);
nor U13403 (N_13403,N_11952,N_10636);
xor U13404 (N_13404,N_11662,N_9704);
or U13405 (N_13405,N_10221,N_11552);
xor U13406 (N_13406,N_11738,N_9178);
xnor U13407 (N_13407,N_11737,N_9842);
nor U13408 (N_13408,N_9898,N_9144);
nor U13409 (N_13409,N_11528,N_9829);
and U13410 (N_13410,N_9339,N_9959);
xnor U13411 (N_13411,N_10345,N_11277);
and U13412 (N_13412,N_10410,N_9147);
nand U13413 (N_13413,N_9260,N_10480);
or U13414 (N_13414,N_10838,N_11314);
or U13415 (N_13415,N_10351,N_9263);
nor U13416 (N_13416,N_9913,N_10784);
and U13417 (N_13417,N_11415,N_9684);
xor U13418 (N_13418,N_9604,N_10120);
or U13419 (N_13419,N_11880,N_11960);
xnor U13420 (N_13420,N_10355,N_11854);
xnor U13421 (N_13421,N_9565,N_9083);
xnor U13422 (N_13422,N_9234,N_10928);
and U13423 (N_13423,N_9548,N_10387);
or U13424 (N_13424,N_9889,N_10999);
and U13425 (N_13425,N_10749,N_10437);
nand U13426 (N_13426,N_10194,N_11827);
xor U13427 (N_13427,N_10802,N_9904);
and U13428 (N_13428,N_10938,N_11613);
nor U13429 (N_13429,N_9207,N_11222);
xor U13430 (N_13430,N_10891,N_11435);
nor U13431 (N_13431,N_11467,N_10182);
nand U13432 (N_13432,N_10127,N_9785);
nand U13433 (N_13433,N_11294,N_11492);
xor U13434 (N_13434,N_9174,N_10598);
nor U13435 (N_13435,N_11229,N_10388);
nor U13436 (N_13436,N_10978,N_9018);
xnor U13437 (N_13437,N_10372,N_10475);
xor U13438 (N_13438,N_9647,N_10916);
or U13439 (N_13439,N_10160,N_11924);
or U13440 (N_13440,N_10751,N_9279);
or U13441 (N_13441,N_9656,N_11438);
or U13442 (N_13442,N_11847,N_11726);
or U13443 (N_13443,N_11740,N_9167);
or U13444 (N_13444,N_9416,N_11311);
xor U13445 (N_13445,N_9061,N_11676);
xnor U13446 (N_13446,N_10739,N_10243);
and U13447 (N_13447,N_10245,N_10902);
and U13448 (N_13448,N_11483,N_10864);
nor U13449 (N_13449,N_9542,N_9047);
or U13450 (N_13450,N_10178,N_9639);
nand U13451 (N_13451,N_9731,N_9058);
or U13452 (N_13452,N_9896,N_11254);
xor U13453 (N_13453,N_10847,N_10805);
and U13454 (N_13454,N_9223,N_11006);
or U13455 (N_13455,N_11863,N_9342);
nor U13456 (N_13456,N_11531,N_11533);
and U13457 (N_13457,N_11501,N_9365);
or U13458 (N_13458,N_9294,N_9072);
or U13459 (N_13459,N_11628,N_10557);
xor U13460 (N_13460,N_9505,N_11702);
nand U13461 (N_13461,N_9620,N_9267);
or U13462 (N_13462,N_9917,N_10323);
xor U13463 (N_13463,N_11829,N_10064);
or U13464 (N_13464,N_11490,N_10817);
nor U13465 (N_13465,N_10899,N_11092);
xor U13466 (N_13466,N_11208,N_11291);
nand U13467 (N_13467,N_10568,N_10229);
nor U13468 (N_13468,N_10386,N_11272);
nand U13469 (N_13469,N_9618,N_11833);
or U13470 (N_13470,N_10205,N_9197);
or U13471 (N_13471,N_11443,N_9289);
nand U13472 (N_13472,N_10256,N_9544);
and U13473 (N_13473,N_11800,N_10982);
xor U13474 (N_13474,N_9307,N_9613);
xnor U13475 (N_13475,N_11355,N_10001);
nor U13476 (N_13476,N_10782,N_11900);
and U13477 (N_13477,N_10593,N_10859);
and U13478 (N_13478,N_11575,N_11099);
and U13479 (N_13479,N_11051,N_9150);
nand U13480 (N_13480,N_9705,N_10198);
or U13481 (N_13481,N_10331,N_10637);
xnor U13482 (N_13482,N_9154,N_11870);
or U13483 (N_13483,N_10153,N_11688);
or U13484 (N_13484,N_9008,N_11074);
or U13485 (N_13485,N_9069,N_11223);
or U13486 (N_13486,N_10282,N_9087);
xor U13487 (N_13487,N_10694,N_10647);
nand U13488 (N_13488,N_10084,N_9060);
nor U13489 (N_13489,N_10433,N_11770);
and U13490 (N_13490,N_11856,N_11861);
and U13491 (N_13491,N_10082,N_10303);
and U13492 (N_13492,N_10686,N_9002);
nand U13493 (N_13493,N_9796,N_10626);
nor U13494 (N_13494,N_9386,N_10921);
and U13495 (N_13495,N_9698,N_11742);
and U13496 (N_13496,N_9484,N_10622);
nor U13497 (N_13497,N_9515,N_11704);
nor U13498 (N_13498,N_11773,N_9216);
xor U13499 (N_13499,N_9664,N_11367);
nor U13500 (N_13500,N_10112,N_9409);
xnor U13501 (N_13501,N_11364,N_9677);
and U13502 (N_13502,N_11312,N_9898);
or U13503 (N_13503,N_9003,N_11302);
nor U13504 (N_13504,N_9958,N_11034);
xor U13505 (N_13505,N_9207,N_11982);
xor U13506 (N_13506,N_11959,N_10143);
xnor U13507 (N_13507,N_10745,N_11257);
nand U13508 (N_13508,N_10409,N_11695);
or U13509 (N_13509,N_11085,N_10290);
xor U13510 (N_13510,N_10806,N_9231);
and U13511 (N_13511,N_10740,N_9812);
xor U13512 (N_13512,N_9712,N_9879);
nand U13513 (N_13513,N_10510,N_10496);
nor U13514 (N_13514,N_11738,N_9050);
nor U13515 (N_13515,N_10673,N_9516);
nand U13516 (N_13516,N_10891,N_11867);
xor U13517 (N_13517,N_9506,N_9038);
nand U13518 (N_13518,N_10866,N_9826);
nor U13519 (N_13519,N_10954,N_11718);
nor U13520 (N_13520,N_9457,N_9546);
nand U13521 (N_13521,N_10478,N_10771);
or U13522 (N_13522,N_11989,N_9337);
nand U13523 (N_13523,N_9969,N_9515);
nor U13524 (N_13524,N_9763,N_9686);
and U13525 (N_13525,N_9891,N_10920);
or U13526 (N_13526,N_10627,N_10693);
or U13527 (N_13527,N_9662,N_9964);
nand U13528 (N_13528,N_9873,N_9819);
xor U13529 (N_13529,N_10706,N_11822);
and U13530 (N_13530,N_10751,N_9188);
or U13531 (N_13531,N_10045,N_10636);
and U13532 (N_13532,N_10930,N_11070);
xor U13533 (N_13533,N_9713,N_11540);
or U13534 (N_13534,N_11299,N_11849);
nand U13535 (N_13535,N_10401,N_11140);
or U13536 (N_13536,N_11743,N_9651);
or U13537 (N_13537,N_10810,N_10721);
or U13538 (N_13538,N_11098,N_10446);
or U13539 (N_13539,N_11273,N_9532);
xnor U13540 (N_13540,N_11525,N_9506);
nand U13541 (N_13541,N_10743,N_9548);
nand U13542 (N_13542,N_10130,N_10005);
and U13543 (N_13543,N_9938,N_9520);
nand U13544 (N_13544,N_10654,N_11764);
and U13545 (N_13545,N_11745,N_10102);
nor U13546 (N_13546,N_9782,N_11851);
nand U13547 (N_13547,N_10110,N_9121);
nor U13548 (N_13548,N_10882,N_9408);
xnor U13549 (N_13549,N_11733,N_11755);
xor U13550 (N_13550,N_11560,N_10192);
xor U13551 (N_13551,N_11349,N_11620);
xor U13552 (N_13552,N_9322,N_11059);
xor U13553 (N_13553,N_10091,N_11161);
nand U13554 (N_13554,N_10543,N_11038);
nor U13555 (N_13555,N_11429,N_11515);
nand U13556 (N_13556,N_9058,N_9504);
nand U13557 (N_13557,N_10755,N_10973);
xnor U13558 (N_13558,N_9430,N_11753);
xor U13559 (N_13559,N_9462,N_9855);
or U13560 (N_13560,N_11597,N_9988);
nand U13561 (N_13561,N_10017,N_10165);
nand U13562 (N_13562,N_9638,N_11473);
and U13563 (N_13563,N_10198,N_11185);
and U13564 (N_13564,N_9905,N_9070);
nor U13565 (N_13565,N_9782,N_9191);
nor U13566 (N_13566,N_9064,N_11673);
or U13567 (N_13567,N_10383,N_10728);
nor U13568 (N_13568,N_11163,N_10823);
nor U13569 (N_13569,N_9224,N_11200);
or U13570 (N_13570,N_10511,N_11532);
or U13571 (N_13571,N_9935,N_10246);
xnor U13572 (N_13572,N_9309,N_11553);
nor U13573 (N_13573,N_9604,N_11502);
nand U13574 (N_13574,N_11790,N_9439);
or U13575 (N_13575,N_10145,N_10033);
or U13576 (N_13576,N_10698,N_11552);
xor U13577 (N_13577,N_10282,N_10029);
or U13578 (N_13578,N_9598,N_9551);
nor U13579 (N_13579,N_11413,N_9744);
or U13580 (N_13580,N_9880,N_9211);
or U13581 (N_13581,N_11260,N_9250);
and U13582 (N_13582,N_10438,N_11249);
nor U13583 (N_13583,N_11595,N_11833);
nand U13584 (N_13584,N_9301,N_10354);
nor U13585 (N_13585,N_11549,N_10216);
nand U13586 (N_13586,N_10538,N_11294);
and U13587 (N_13587,N_10603,N_9095);
nor U13588 (N_13588,N_10711,N_11513);
or U13589 (N_13589,N_10629,N_11080);
nand U13590 (N_13590,N_9210,N_11071);
nand U13591 (N_13591,N_9700,N_10480);
nand U13592 (N_13592,N_9844,N_10875);
nor U13593 (N_13593,N_11559,N_10087);
and U13594 (N_13594,N_11037,N_10967);
nand U13595 (N_13595,N_9466,N_10152);
and U13596 (N_13596,N_11233,N_9009);
xor U13597 (N_13597,N_9873,N_11010);
nor U13598 (N_13598,N_11953,N_11206);
xnor U13599 (N_13599,N_11310,N_9448);
xor U13600 (N_13600,N_9586,N_11663);
xor U13601 (N_13601,N_10221,N_10926);
and U13602 (N_13602,N_9561,N_10754);
xnor U13603 (N_13603,N_10744,N_11573);
or U13604 (N_13604,N_10473,N_11325);
nand U13605 (N_13605,N_11604,N_10267);
nand U13606 (N_13606,N_10510,N_10731);
nand U13607 (N_13607,N_9154,N_10826);
or U13608 (N_13608,N_10975,N_11977);
or U13609 (N_13609,N_9416,N_9348);
nand U13610 (N_13610,N_10970,N_11764);
nand U13611 (N_13611,N_11179,N_11352);
nor U13612 (N_13612,N_11226,N_9701);
or U13613 (N_13613,N_9002,N_9796);
nor U13614 (N_13614,N_11132,N_11593);
nor U13615 (N_13615,N_11786,N_9089);
nor U13616 (N_13616,N_10776,N_10107);
or U13617 (N_13617,N_9321,N_9789);
and U13618 (N_13618,N_11018,N_11357);
or U13619 (N_13619,N_10231,N_9307);
nor U13620 (N_13620,N_10443,N_10641);
nand U13621 (N_13621,N_10265,N_9701);
xor U13622 (N_13622,N_9190,N_10217);
xor U13623 (N_13623,N_9170,N_9896);
and U13624 (N_13624,N_9954,N_10092);
nor U13625 (N_13625,N_11548,N_11679);
xnor U13626 (N_13626,N_10181,N_9955);
and U13627 (N_13627,N_9548,N_10155);
nand U13628 (N_13628,N_9477,N_11637);
xnor U13629 (N_13629,N_10665,N_9250);
nand U13630 (N_13630,N_9012,N_11749);
xnor U13631 (N_13631,N_11071,N_9913);
nor U13632 (N_13632,N_9081,N_9256);
and U13633 (N_13633,N_10213,N_9707);
nor U13634 (N_13634,N_9886,N_10623);
nor U13635 (N_13635,N_9338,N_10361);
or U13636 (N_13636,N_11323,N_10770);
xor U13637 (N_13637,N_9757,N_11712);
and U13638 (N_13638,N_11397,N_11786);
or U13639 (N_13639,N_11629,N_9784);
and U13640 (N_13640,N_9966,N_9932);
xor U13641 (N_13641,N_10269,N_11411);
nor U13642 (N_13642,N_10107,N_11077);
or U13643 (N_13643,N_9658,N_10796);
or U13644 (N_13644,N_11159,N_10547);
or U13645 (N_13645,N_9585,N_9718);
nor U13646 (N_13646,N_11548,N_10750);
nand U13647 (N_13647,N_9535,N_10058);
and U13648 (N_13648,N_9520,N_10569);
nor U13649 (N_13649,N_11538,N_11224);
nor U13650 (N_13650,N_11272,N_9580);
nor U13651 (N_13651,N_10002,N_9355);
nand U13652 (N_13652,N_11736,N_11743);
or U13653 (N_13653,N_11619,N_10743);
nor U13654 (N_13654,N_11056,N_10573);
and U13655 (N_13655,N_9735,N_11657);
nand U13656 (N_13656,N_10473,N_11442);
xor U13657 (N_13657,N_11275,N_10825);
and U13658 (N_13658,N_11502,N_10139);
nand U13659 (N_13659,N_10962,N_9116);
nand U13660 (N_13660,N_10774,N_11582);
or U13661 (N_13661,N_9188,N_11518);
xnor U13662 (N_13662,N_9209,N_9198);
and U13663 (N_13663,N_10930,N_10065);
nor U13664 (N_13664,N_9507,N_9545);
or U13665 (N_13665,N_10830,N_10163);
and U13666 (N_13666,N_11238,N_11350);
nor U13667 (N_13667,N_10572,N_9408);
or U13668 (N_13668,N_11619,N_10836);
and U13669 (N_13669,N_10990,N_11630);
and U13670 (N_13670,N_11237,N_9859);
xor U13671 (N_13671,N_9065,N_11456);
and U13672 (N_13672,N_11135,N_11266);
nor U13673 (N_13673,N_11126,N_11480);
nor U13674 (N_13674,N_10499,N_10693);
nor U13675 (N_13675,N_11590,N_11754);
nor U13676 (N_13676,N_9319,N_10819);
xnor U13677 (N_13677,N_11230,N_9649);
and U13678 (N_13678,N_10600,N_9575);
xnor U13679 (N_13679,N_9503,N_9102);
xor U13680 (N_13680,N_10577,N_10802);
and U13681 (N_13681,N_9814,N_11121);
or U13682 (N_13682,N_9737,N_9838);
or U13683 (N_13683,N_11034,N_10016);
xor U13684 (N_13684,N_9640,N_10753);
nor U13685 (N_13685,N_10281,N_11886);
nor U13686 (N_13686,N_11565,N_9942);
and U13687 (N_13687,N_9775,N_9513);
nand U13688 (N_13688,N_11963,N_10873);
or U13689 (N_13689,N_10074,N_10328);
xor U13690 (N_13690,N_11651,N_10137);
nor U13691 (N_13691,N_10452,N_9638);
xor U13692 (N_13692,N_10659,N_10947);
nand U13693 (N_13693,N_10525,N_9510);
nand U13694 (N_13694,N_10785,N_11599);
and U13695 (N_13695,N_9648,N_9198);
or U13696 (N_13696,N_10757,N_10963);
or U13697 (N_13697,N_9900,N_11405);
nand U13698 (N_13698,N_11685,N_11639);
or U13699 (N_13699,N_11058,N_10858);
nand U13700 (N_13700,N_11099,N_10680);
and U13701 (N_13701,N_10466,N_11398);
xnor U13702 (N_13702,N_10358,N_9152);
nand U13703 (N_13703,N_11624,N_11882);
nor U13704 (N_13704,N_10772,N_10318);
xor U13705 (N_13705,N_11893,N_10599);
nand U13706 (N_13706,N_9935,N_11453);
nor U13707 (N_13707,N_11653,N_10621);
or U13708 (N_13708,N_11599,N_9208);
or U13709 (N_13709,N_11253,N_11604);
nor U13710 (N_13710,N_10865,N_9479);
xnor U13711 (N_13711,N_10704,N_9122);
or U13712 (N_13712,N_10460,N_9818);
and U13713 (N_13713,N_10664,N_9733);
and U13714 (N_13714,N_9392,N_11774);
and U13715 (N_13715,N_10361,N_11974);
nand U13716 (N_13716,N_11354,N_10721);
and U13717 (N_13717,N_10758,N_10179);
and U13718 (N_13718,N_10982,N_10918);
nor U13719 (N_13719,N_11439,N_10318);
nand U13720 (N_13720,N_11442,N_10851);
xnor U13721 (N_13721,N_11482,N_9540);
xor U13722 (N_13722,N_11985,N_11619);
or U13723 (N_13723,N_11381,N_9420);
and U13724 (N_13724,N_10025,N_11297);
or U13725 (N_13725,N_9068,N_11949);
and U13726 (N_13726,N_11509,N_10566);
and U13727 (N_13727,N_9778,N_11859);
nor U13728 (N_13728,N_10888,N_9167);
or U13729 (N_13729,N_9354,N_10014);
and U13730 (N_13730,N_10782,N_9147);
or U13731 (N_13731,N_10528,N_11751);
and U13732 (N_13732,N_11025,N_11103);
and U13733 (N_13733,N_9432,N_11500);
and U13734 (N_13734,N_11199,N_9035);
nor U13735 (N_13735,N_11567,N_9689);
nor U13736 (N_13736,N_10163,N_11546);
nand U13737 (N_13737,N_11169,N_9216);
nor U13738 (N_13738,N_11722,N_10486);
nor U13739 (N_13739,N_9620,N_11397);
nor U13740 (N_13740,N_10504,N_10515);
xnor U13741 (N_13741,N_11045,N_11503);
nand U13742 (N_13742,N_10474,N_11817);
or U13743 (N_13743,N_11273,N_10667);
nand U13744 (N_13744,N_9768,N_11020);
or U13745 (N_13745,N_9389,N_11913);
and U13746 (N_13746,N_10175,N_11436);
and U13747 (N_13747,N_9227,N_10364);
and U13748 (N_13748,N_9946,N_9500);
or U13749 (N_13749,N_10347,N_10517);
nor U13750 (N_13750,N_11499,N_11567);
nor U13751 (N_13751,N_10626,N_10969);
xnor U13752 (N_13752,N_9780,N_10657);
and U13753 (N_13753,N_11208,N_9363);
or U13754 (N_13754,N_9657,N_10826);
nor U13755 (N_13755,N_10564,N_11432);
and U13756 (N_13756,N_10017,N_10390);
and U13757 (N_13757,N_10253,N_11665);
or U13758 (N_13758,N_9924,N_9947);
and U13759 (N_13759,N_9258,N_11255);
and U13760 (N_13760,N_10918,N_11971);
nand U13761 (N_13761,N_10510,N_9225);
xor U13762 (N_13762,N_11953,N_9797);
xnor U13763 (N_13763,N_10097,N_9581);
xor U13764 (N_13764,N_9922,N_10072);
nand U13765 (N_13765,N_10903,N_11493);
nor U13766 (N_13766,N_9609,N_11444);
xor U13767 (N_13767,N_9337,N_9072);
and U13768 (N_13768,N_11995,N_11424);
and U13769 (N_13769,N_11521,N_10174);
xor U13770 (N_13770,N_10935,N_11359);
or U13771 (N_13771,N_10955,N_10690);
or U13772 (N_13772,N_9904,N_9837);
or U13773 (N_13773,N_9937,N_10815);
xnor U13774 (N_13774,N_10940,N_9426);
nor U13775 (N_13775,N_11750,N_11859);
nor U13776 (N_13776,N_10235,N_9217);
and U13777 (N_13777,N_10442,N_10612);
or U13778 (N_13778,N_11137,N_11432);
nand U13779 (N_13779,N_10530,N_9153);
xor U13780 (N_13780,N_11358,N_10817);
or U13781 (N_13781,N_11340,N_11855);
and U13782 (N_13782,N_10623,N_11009);
or U13783 (N_13783,N_9728,N_9780);
nor U13784 (N_13784,N_10574,N_9677);
nand U13785 (N_13785,N_9857,N_10982);
xor U13786 (N_13786,N_11489,N_11530);
or U13787 (N_13787,N_11450,N_10524);
nor U13788 (N_13788,N_9354,N_9382);
xnor U13789 (N_13789,N_10369,N_9651);
nand U13790 (N_13790,N_9446,N_11859);
nor U13791 (N_13791,N_9562,N_9165);
nand U13792 (N_13792,N_10190,N_11142);
nor U13793 (N_13793,N_11003,N_10721);
or U13794 (N_13794,N_11737,N_10274);
or U13795 (N_13795,N_11798,N_10041);
nor U13796 (N_13796,N_11073,N_10662);
or U13797 (N_13797,N_11989,N_11440);
xnor U13798 (N_13798,N_11877,N_10595);
nand U13799 (N_13799,N_10917,N_11184);
nor U13800 (N_13800,N_11674,N_11603);
and U13801 (N_13801,N_11948,N_11047);
nor U13802 (N_13802,N_9251,N_10395);
and U13803 (N_13803,N_9415,N_10372);
nand U13804 (N_13804,N_9664,N_10622);
nand U13805 (N_13805,N_9038,N_10641);
and U13806 (N_13806,N_11549,N_9709);
nand U13807 (N_13807,N_10847,N_10563);
or U13808 (N_13808,N_10297,N_10702);
xnor U13809 (N_13809,N_11741,N_10807);
or U13810 (N_13810,N_9773,N_9701);
and U13811 (N_13811,N_9937,N_10153);
nand U13812 (N_13812,N_10816,N_10475);
xor U13813 (N_13813,N_9797,N_11738);
xor U13814 (N_13814,N_11653,N_11713);
xnor U13815 (N_13815,N_10078,N_9181);
nand U13816 (N_13816,N_10080,N_10569);
or U13817 (N_13817,N_11589,N_10076);
nor U13818 (N_13818,N_9253,N_11472);
and U13819 (N_13819,N_9705,N_11243);
or U13820 (N_13820,N_9947,N_9892);
or U13821 (N_13821,N_9834,N_11137);
or U13822 (N_13822,N_9229,N_11380);
or U13823 (N_13823,N_11694,N_9740);
nor U13824 (N_13824,N_9315,N_10843);
xor U13825 (N_13825,N_10803,N_11270);
or U13826 (N_13826,N_9829,N_10006);
nand U13827 (N_13827,N_10062,N_11801);
nand U13828 (N_13828,N_9589,N_10094);
xor U13829 (N_13829,N_9127,N_10841);
nor U13830 (N_13830,N_9376,N_9460);
xor U13831 (N_13831,N_9751,N_10399);
nand U13832 (N_13832,N_9203,N_11192);
nor U13833 (N_13833,N_10712,N_10065);
nand U13834 (N_13834,N_9779,N_10932);
xor U13835 (N_13835,N_11050,N_9418);
nand U13836 (N_13836,N_10425,N_11930);
and U13837 (N_13837,N_9307,N_10465);
nand U13838 (N_13838,N_9908,N_11440);
or U13839 (N_13839,N_10369,N_10156);
or U13840 (N_13840,N_9197,N_10639);
and U13841 (N_13841,N_9743,N_10075);
xor U13842 (N_13842,N_10700,N_10233);
nand U13843 (N_13843,N_11061,N_11887);
nor U13844 (N_13844,N_11199,N_11974);
nand U13845 (N_13845,N_9819,N_11576);
or U13846 (N_13846,N_10191,N_9715);
nand U13847 (N_13847,N_10469,N_11319);
nand U13848 (N_13848,N_11738,N_11776);
nor U13849 (N_13849,N_10762,N_11627);
nand U13850 (N_13850,N_10687,N_9131);
or U13851 (N_13851,N_11057,N_9568);
nor U13852 (N_13852,N_10814,N_9247);
nor U13853 (N_13853,N_9226,N_11838);
and U13854 (N_13854,N_9890,N_10398);
nor U13855 (N_13855,N_9242,N_9914);
xnor U13856 (N_13856,N_11749,N_10885);
or U13857 (N_13857,N_11586,N_11054);
or U13858 (N_13858,N_11222,N_9593);
or U13859 (N_13859,N_10950,N_9863);
nand U13860 (N_13860,N_11019,N_9154);
nor U13861 (N_13861,N_10537,N_11361);
nor U13862 (N_13862,N_11840,N_11801);
xor U13863 (N_13863,N_11767,N_10994);
or U13864 (N_13864,N_9226,N_11094);
xnor U13865 (N_13865,N_10726,N_11257);
xor U13866 (N_13866,N_9341,N_9491);
nor U13867 (N_13867,N_10229,N_10526);
or U13868 (N_13868,N_9025,N_10707);
and U13869 (N_13869,N_10286,N_11186);
xnor U13870 (N_13870,N_10108,N_9854);
nand U13871 (N_13871,N_11167,N_10141);
nand U13872 (N_13872,N_10499,N_11854);
nor U13873 (N_13873,N_11217,N_11876);
nand U13874 (N_13874,N_10362,N_10510);
nand U13875 (N_13875,N_9901,N_9093);
nor U13876 (N_13876,N_9338,N_10839);
xor U13877 (N_13877,N_11943,N_11597);
or U13878 (N_13878,N_10965,N_11890);
nand U13879 (N_13879,N_10813,N_11529);
and U13880 (N_13880,N_10332,N_10221);
and U13881 (N_13881,N_9528,N_11890);
xor U13882 (N_13882,N_9466,N_11386);
nor U13883 (N_13883,N_10396,N_9854);
xor U13884 (N_13884,N_11230,N_9089);
nand U13885 (N_13885,N_11540,N_9340);
or U13886 (N_13886,N_9735,N_9517);
xnor U13887 (N_13887,N_11576,N_11544);
nor U13888 (N_13888,N_9862,N_9941);
xor U13889 (N_13889,N_11093,N_10235);
xor U13890 (N_13890,N_10642,N_9569);
nor U13891 (N_13891,N_10034,N_9602);
nor U13892 (N_13892,N_9877,N_9920);
xnor U13893 (N_13893,N_11297,N_9666);
nor U13894 (N_13894,N_11475,N_11312);
nor U13895 (N_13895,N_10886,N_10912);
nand U13896 (N_13896,N_11689,N_9602);
and U13897 (N_13897,N_9561,N_10702);
or U13898 (N_13898,N_11453,N_11643);
nand U13899 (N_13899,N_11638,N_11691);
and U13900 (N_13900,N_11767,N_11138);
or U13901 (N_13901,N_10967,N_10370);
nor U13902 (N_13902,N_9970,N_10493);
and U13903 (N_13903,N_11563,N_11675);
nor U13904 (N_13904,N_10387,N_10786);
and U13905 (N_13905,N_9360,N_11155);
or U13906 (N_13906,N_10384,N_10991);
nand U13907 (N_13907,N_10220,N_9126);
nor U13908 (N_13908,N_9769,N_10677);
xor U13909 (N_13909,N_10122,N_10344);
xor U13910 (N_13910,N_10171,N_11110);
nand U13911 (N_13911,N_10938,N_9266);
nand U13912 (N_13912,N_9949,N_11311);
nor U13913 (N_13913,N_10169,N_9032);
xor U13914 (N_13914,N_10487,N_10674);
or U13915 (N_13915,N_9947,N_11329);
and U13916 (N_13916,N_9130,N_11091);
nand U13917 (N_13917,N_10643,N_9163);
nand U13918 (N_13918,N_9027,N_10173);
nor U13919 (N_13919,N_10356,N_9660);
nor U13920 (N_13920,N_11253,N_9109);
nor U13921 (N_13921,N_10040,N_9068);
nor U13922 (N_13922,N_11292,N_9889);
and U13923 (N_13923,N_9730,N_10168);
nor U13924 (N_13924,N_11076,N_10916);
xnor U13925 (N_13925,N_11670,N_10491);
nor U13926 (N_13926,N_10219,N_11022);
nor U13927 (N_13927,N_11161,N_9522);
and U13928 (N_13928,N_11360,N_9431);
or U13929 (N_13929,N_11850,N_11912);
or U13930 (N_13930,N_11941,N_10418);
nor U13931 (N_13931,N_11609,N_10258);
and U13932 (N_13932,N_11783,N_10827);
nor U13933 (N_13933,N_9512,N_9421);
xor U13934 (N_13934,N_9710,N_11097);
nand U13935 (N_13935,N_10480,N_9328);
and U13936 (N_13936,N_9388,N_11113);
nand U13937 (N_13937,N_9869,N_9353);
and U13938 (N_13938,N_11025,N_9015);
and U13939 (N_13939,N_9537,N_9061);
or U13940 (N_13940,N_10428,N_9197);
and U13941 (N_13941,N_11556,N_11152);
or U13942 (N_13942,N_10468,N_10447);
or U13943 (N_13943,N_11529,N_9305);
or U13944 (N_13944,N_10443,N_10260);
xor U13945 (N_13945,N_9929,N_11988);
and U13946 (N_13946,N_9808,N_11220);
nand U13947 (N_13947,N_10261,N_9895);
xnor U13948 (N_13948,N_10439,N_9454);
or U13949 (N_13949,N_9579,N_9571);
and U13950 (N_13950,N_10428,N_11382);
nand U13951 (N_13951,N_10711,N_11292);
and U13952 (N_13952,N_11402,N_9182);
nor U13953 (N_13953,N_11983,N_9376);
nand U13954 (N_13954,N_9776,N_11180);
or U13955 (N_13955,N_11497,N_10445);
and U13956 (N_13956,N_10751,N_11628);
and U13957 (N_13957,N_10950,N_11410);
nor U13958 (N_13958,N_11083,N_11346);
nor U13959 (N_13959,N_11959,N_9210);
nand U13960 (N_13960,N_11687,N_9907);
and U13961 (N_13961,N_11317,N_9028);
nand U13962 (N_13962,N_11269,N_11576);
and U13963 (N_13963,N_10973,N_10730);
xor U13964 (N_13964,N_9521,N_9829);
and U13965 (N_13965,N_10858,N_9977);
and U13966 (N_13966,N_11674,N_10849);
nand U13967 (N_13967,N_9994,N_9309);
xnor U13968 (N_13968,N_10086,N_11234);
nand U13969 (N_13969,N_9460,N_10748);
xnor U13970 (N_13970,N_10555,N_11103);
xor U13971 (N_13971,N_9554,N_11303);
nor U13972 (N_13972,N_11729,N_10515);
nand U13973 (N_13973,N_10849,N_11273);
and U13974 (N_13974,N_10016,N_10150);
and U13975 (N_13975,N_10167,N_11458);
nor U13976 (N_13976,N_11051,N_10066);
or U13977 (N_13977,N_10710,N_9642);
and U13978 (N_13978,N_9913,N_11381);
xnor U13979 (N_13979,N_10521,N_9566);
xnor U13980 (N_13980,N_10460,N_9874);
or U13981 (N_13981,N_9503,N_10916);
or U13982 (N_13982,N_10002,N_11389);
nand U13983 (N_13983,N_10462,N_10583);
or U13984 (N_13984,N_11664,N_10950);
nor U13985 (N_13985,N_11390,N_9263);
xnor U13986 (N_13986,N_11270,N_9898);
nand U13987 (N_13987,N_9711,N_11183);
xor U13988 (N_13988,N_9064,N_9737);
nand U13989 (N_13989,N_10084,N_11842);
and U13990 (N_13990,N_10269,N_10851);
and U13991 (N_13991,N_11099,N_10874);
xnor U13992 (N_13992,N_10010,N_11913);
xor U13993 (N_13993,N_11245,N_10512);
nor U13994 (N_13994,N_10181,N_10166);
nand U13995 (N_13995,N_11763,N_9985);
and U13996 (N_13996,N_9615,N_9708);
xor U13997 (N_13997,N_9102,N_10358);
nor U13998 (N_13998,N_11168,N_9700);
nand U13999 (N_13999,N_9502,N_10512);
xnor U14000 (N_14000,N_9548,N_10576);
nor U14001 (N_14001,N_10476,N_9243);
and U14002 (N_14002,N_11613,N_10806);
nor U14003 (N_14003,N_9704,N_10525);
xnor U14004 (N_14004,N_9833,N_9700);
and U14005 (N_14005,N_11857,N_9090);
and U14006 (N_14006,N_11413,N_11162);
nor U14007 (N_14007,N_10037,N_11128);
xor U14008 (N_14008,N_11402,N_9423);
xnor U14009 (N_14009,N_9796,N_10158);
and U14010 (N_14010,N_11243,N_11950);
and U14011 (N_14011,N_10486,N_9824);
nor U14012 (N_14012,N_9078,N_11783);
nor U14013 (N_14013,N_11686,N_10368);
xor U14014 (N_14014,N_9197,N_10020);
nand U14015 (N_14015,N_10539,N_11505);
and U14016 (N_14016,N_11588,N_11095);
and U14017 (N_14017,N_11557,N_10064);
and U14018 (N_14018,N_11562,N_10409);
nand U14019 (N_14019,N_11818,N_10519);
and U14020 (N_14020,N_10402,N_11869);
xnor U14021 (N_14021,N_10847,N_9571);
or U14022 (N_14022,N_9568,N_9536);
or U14023 (N_14023,N_10065,N_11062);
nand U14024 (N_14024,N_10244,N_11569);
or U14025 (N_14025,N_9300,N_11617);
and U14026 (N_14026,N_10157,N_9489);
nand U14027 (N_14027,N_11387,N_11561);
nand U14028 (N_14028,N_9846,N_10620);
nand U14029 (N_14029,N_11883,N_10935);
xnor U14030 (N_14030,N_11036,N_9911);
xor U14031 (N_14031,N_9691,N_10011);
nor U14032 (N_14032,N_10016,N_10050);
or U14033 (N_14033,N_10807,N_10818);
nor U14034 (N_14034,N_9860,N_10115);
xnor U14035 (N_14035,N_10030,N_11363);
xor U14036 (N_14036,N_10054,N_10512);
nand U14037 (N_14037,N_9099,N_11748);
nor U14038 (N_14038,N_9423,N_9895);
xor U14039 (N_14039,N_11472,N_10689);
xnor U14040 (N_14040,N_11454,N_10179);
and U14041 (N_14041,N_11853,N_9536);
xor U14042 (N_14042,N_11694,N_10089);
xor U14043 (N_14043,N_10943,N_9975);
nand U14044 (N_14044,N_11862,N_9964);
and U14045 (N_14045,N_11941,N_10485);
nor U14046 (N_14046,N_10829,N_11464);
nor U14047 (N_14047,N_9518,N_11726);
or U14048 (N_14048,N_11724,N_10771);
and U14049 (N_14049,N_10708,N_9064);
nand U14050 (N_14050,N_9015,N_10582);
and U14051 (N_14051,N_11910,N_9883);
and U14052 (N_14052,N_10247,N_11431);
nand U14053 (N_14053,N_11761,N_11299);
nor U14054 (N_14054,N_9913,N_11003);
and U14055 (N_14055,N_9660,N_10069);
xnor U14056 (N_14056,N_10599,N_9829);
xnor U14057 (N_14057,N_10242,N_10853);
nand U14058 (N_14058,N_9028,N_9252);
xor U14059 (N_14059,N_9485,N_10890);
xnor U14060 (N_14060,N_10605,N_10216);
nor U14061 (N_14061,N_10494,N_10398);
xnor U14062 (N_14062,N_11944,N_10685);
nor U14063 (N_14063,N_9238,N_11041);
or U14064 (N_14064,N_9884,N_9154);
xor U14065 (N_14065,N_9812,N_9529);
xor U14066 (N_14066,N_9238,N_9930);
nor U14067 (N_14067,N_10239,N_10473);
and U14068 (N_14068,N_9382,N_9228);
nor U14069 (N_14069,N_10449,N_9545);
xnor U14070 (N_14070,N_11139,N_11282);
and U14071 (N_14071,N_11589,N_10527);
or U14072 (N_14072,N_11505,N_10124);
nand U14073 (N_14073,N_11794,N_9057);
and U14074 (N_14074,N_11088,N_9747);
and U14075 (N_14075,N_10667,N_9474);
nand U14076 (N_14076,N_11186,N_9313);
xor U14077 (N_14077,N_10224,N_9403);
or U14078 (N_14078,N_11177,N_10431);
xnor U14079 (N_14079,N_10334,N_10792);
xor U14080 (N_14080,N_10420,N_9951);
xor U14081 (N_14081,N_10575,N_9545);
and U14082 (N_14082,N_11073,N_9689);
nor U14083 (N_14083,N_11652,N_10799);
and U14084 (N_14084,N_9566,N_10419);
nor U14085 (N_14085,N_9520,N_10638);
or U14086 (N_14086,N_9486,N_11965);
and U14087 (N_14087,N_10865,N_9850);
or U14088 (N_14088,N_11613,N_9996);
or U14089 (N_14089,N_10914,N_9644);
nor U14090 (N_14090,N_10500,N_9930);
and U14091 (N_14091,N_11387,N_10703);
nand U14092 (N_14092,N_11836,N_10394);
xnor U14093 (N_14093,N_9601,N_11830);
xnor U14094 (N_14094,N_11294,N_10124);
nor U14095 (N_14095,N_11745,N_11786);
nor U14096 (N_14096,N_10829,N_11979);
and U14097 (N_14097,N_10625,N_11444);
nand U14098 (N_14098,N_11874,N_9266);
and U14099 (N_14099,N_9092,N_11187);
or U14100 (N_14100,N_10833,N_9308);
and U14101 (N_14101,N_10709,N_10844);
and U14102 (N_14102,N_11057,N_11863);
or U14103 (N_14103,N_11260,N_10935);
and U14104 (N_14104,N_9788,N_9369);
nor U14105 (N_14105,N_11579,N_10660);
nand U14106 (N_14106,N_11087,N_11858);
xor U14107 (N_14107,N_9739,N_9939);
nand U14108 (N_14108,N_10626,N_10488);
xnor U14109 (N_14109,N_10416,N_9434);
nand U14110 (N_14110,N_10903,N_11057);
or U14111 (N_14111,N_10888,N_9505);
xor U14112 (N_14112,N_10326,N_9001);
and U14113 (N_14113,N_9221,N_11952);
nor U14114 (N_14114,N_10691,N_10388);
and U14115 (N_14115,N_11501,N_10995);
or U14116 (N_14116,N_10749,N_11041);
xnor U14117 (N_14117,N_11598,N_11033);
nor U14118 (N_14118,N_9143,N_10622);
nand U14119 (N_14119,N_10748,N_11012);
or U14120 (N_14120,N_10539,N_10025);
nor U14121 (N_14121,N_10575,N_11395);
or U14122 (N_14122,N_11669,N_9738);
xor U14123 (N_14123,N_11496,N_10806);
nand U14124 (N_14124,N_10579,N_10042);
nor U14125 (N_14125,N_9204,N_11764);
nand U14126 (N_14126,N_11107,N_9435);
and U14127 (N_14127,N_10800,N_11151);
nand U14128 (N_14128,N_9033,N_9836);
nor U14129 (N_14129,N_11396,N_9200);
xnor U14130 (N_14130,N_9619,N_10813);
nand U14131 (N_14131,N_10875,N_10281);
or U14132 (N_14132,N_11322,N_9077);
nand U14133 (N_14133,N_11690,N_9153);
nor U14134 (N_14134,N_11702,N_11157);
and U14135 (N_14135,N_11337,N_10472);
nor U14136 (N_14136,N_11933,N_10682);
nand U14137 (N_14137,N_9307,N_10563);
nand U14138 (N_14138,N_10553,N_9327);
and U14139 (N_14139,N_10353,N_10134);
xor U14140 (N_14140,N_9104,N_9493);
nor U14141 (N_14141,N_10360,N_11060);
nor U14142 (N_14142,N_9054,N_9324);
and U14143 (N_14143,N_9411,N_11204);
nor U14144 (N_14144,N_9557,N_9371);
nor U14145 (N_14145,N_11056,N_9201);
or U14146 (N_14146,N_11043,N_10974);
and U14147 (N_14147,N_10600,N_10249);
xor U14148 (N_14148,N_9220,N_11745);
nor U14149 (N_14149,N_11388,N_9883);
and U14150 (N_14150,N_10349,N_9196);
xor U14151 (N_14151,N_10655,N_11452);
or U14152 (N_14152,N_10014,N_10845);
and U14153 (N_14153,N_10680,N_11751);
nor U14154 (N_14154,N_10735,N_11101);
nand U14155 (N_14155,N_11846,N_9522);
nand U14156 (N_14156,N_10099,N_11807);
and U14157 (N_14157,N_11788,N_11625);
or U14158 (N_14158,N_10943,N_10730);
nor U14159 (N_14159,N_10380,N_9369);
and U14160 (N_14160,N_9465,N_9932);
or U14161 (N_14161,N_11919,N_9652);
xor U14162 (N_14162,N_11913,N_11220);
xor U14163 (N_14163,N_11485,N_9658);
nor U14164 (N_14164,N_9981,N_10947);
nand U14165 (N_14165,N_10869,N_9060);
nand U14166 (N_14166,N_9929,N_9107);
nand U14167 (N_14167,N_10540,N_9581);
nor U14168 (N_14168,N_9608,N_10858);
nor U14169 (N_14169,N_10836,N_10041);
nor U14170 (N_14170,N_11841,N_9358);
and U14171 (N_14171,N_9753,N_10867);
nand U14172 (N_14172,N_10111,N_11367);
or U14173 (N_14173,N_11998,N_9028);
and U14174 (N_14174,N_11535,N_10257);
xnor U14175 (N_14175,N_9847,N_9005);
nand U14176 (N_14176,N_9020,N_11549);
xnor U14177 (N_14177,N_10265,N_9056);
or U14178 (N_14178,N_9768,N_11068);
nand U14179 (N_14179,N_10125,N_9292);
xnor U14180 (N_14180,N_10733,N_10098);
and U14181 (N_14181,N_10491,N_9451);
and U14182 (N_14182,N_10805,N_10267);
or U14183 (N_14183,N_9221,N_10986);
or U14184 (N_14184,N_9923,N_10276);
xor U14185 (N_14185,N_10674,N_10309);
or U14186 (N_14186,N_10671,N_11695);
or U14187 (N_14187,N_10912,N_9475);
and U14188 (N_14188,N_9291,N_9315);
or U14189 (N_14189,N_9123,N_9319);
or U14190 (N_14190,N_11361,N_10383);
xnor U14191 (N_14191,N_10960,N_10231);
xnor U14192 (N_14192,N_9615,N_10590);
and U14193 (N_14193,N_10412,N_11300);
and U14194 (N_14194,N_11612,N_11195);
and U14195 (N_14195,N_9247,N_11279);
and U14196 (N_14196,N_11308,N_10338);
or U14197 (N_14197,N_11937,N_10142);
nor U14198 (N_14198,N_11309,N_11869);
nor U14199 (N_14199,N_11707,N_10027);
and U14200 (N_14200,N_11465,N_11316);
nand U14201 (N_14201,N_10223,N_9443);
nand U14202 (N_14202,N_9113,N_11087);
and U14203 (N_14203,N_10242,N_11755);
nand U14204 (N_14204,N_9908,N_10456);
or U14205 (N_14205,N_10217,N_11809);
nor U14206 (N_14206,N_9726,N_11758);
xor U14207 (N_14207,N_10550,N_10352);
xnor U14208 (N_14208,N_10099,N_10335);
nor U14209 (N_14209,N_10571,N_9700);
nand U14210 (N_14210,N_10148,N_11892);
nand U14211 (N_14211,N_11467,N_10232);
and U14212 (N_14212,N_9308,N_9753);
and U14213 (N_14213,N_9624,N_10102);
nor U14214 (N_14214,N_9921,N_10782);
nor U14215 (N_14215,N_10483,N_9296);
nor U14216 (N_14216,N_10124,N_11842);
or U14217 (N_14217,N_9131,N_11905);
nor U14218 (N_14218,N_9189,N_9279);
nor U14219 (N_14219,N_11412,N_11388);
and U14220 (N_14220,N_9809,N_9612);
nor U14221 (N_14221,N_11776,N_9666);
nor U14222 (N_14222,N_11442,N_10971);
xor U14223 (N_14223,N_11299,N_10707);
and U14224 (N_14224,N_11925,N_11337);
and U14225 (N_14225,N_11089,N_10163);
nand U14226 (N_14226,N_9654,N_10654);
and U14227 (N_14227,N_9761,N_11739);
xor U14228 (N_14228,N_10125,N_10322);
or U14229 (N_14229,N_10497,N_11404);
xor U14230 (N_14230,N_11347,N_9346);
nor U14231 (N_14231,N_10545,N_11828);
nor U14232 (N_14232,N_11963,N_11953);
xnor U14233 (N_14233,N_9397,N_10523);
nor U14234 (N_14234,N_10637,N_9447);
and U14235 (N_14235,N_9418,N_9725);
nand U14236 (N_14236,N_10266,N_9393);
or U14237 (N_14237,N_9119,N_10366);
nor U14238 (N_14238,N_9462,N_11422);
nand U14239 (N_14239,N_9005,N_11804);
nor U14240 (N_14240,N_9000,N_11709);
or U14241 (N_14241,N_9994,N_10635);
and U14242 (N_14242,N_9820,N_11880);
xor U14243 (N_14243,N_9418,N_10885);
and U14244 (N_14244,N_11500,N_9852);
xor U14245 (N_14245,N_10080,N_11484);
nand U14246 (N_14246,N_10822,N_9208);
and U14247 (N_14247,N_11075,N_9564);
or U14248 (N_14248,N_11142,N_11095);
nand U14249 (N_14249,N_11356,N_11149);
and U14250 (N_14250,N_11773,N_11248);
nand U14251 (N_14251,N_9506,N_10780);
nor U14252 (N_14252,N_9736,N_10889);
and U14253 (N_14253,N_11019,N_10898);
xnor U14254 (N_14254,N_11634,N_11883);
or U14255 (N_14255,N_9524,N_9882);
or U14256 (N_14256,N_10268,N_11671);
xor U14257 (N_14257,N_11355,N_10187);
xnor U14258 (N_14258,N_9202,N_11632);
nor U14259 (N_14259,N_10200,N_9408);
and U14260 (N_14260,N_10991,N_11841);
xnor U14261 (N_14261,N_9084,N_9969);
xor U14262 (N_14262,N_9968,N_10144);
xor U14263 (N_14263,N_11787,N_10221);
nor U14264 (N_14264,N_10882,N_11756);
nand U14265 (N_14265,N_11200,N_9486);
and U14266 (N_14266,N_9368,N_10926);
nand U14267 (N_14267,N_9694,N_11292);
and U14268 (N_14268,N_9730,N_9176);
nor U14269 (N_14269,N_9805,N_9708);
nand U14270 (N_14270,N_9004,N_10793);
or U14271 (N_14271,N_10363,N_9248);
nand U14272 (N_14272,N_9431,N_11041);
and U14273 (N_14273,N_10691,N_9372);
and U14274 (N_14274,N_11109,N_9900);
and U14275 (N_14275,N_11683,N_9034);
xnor U14276 (N_14276,N_11989,N_11303);
xor U14277 (N_14277,N_10966,N_9494);
or U14278 (N_14278,N_11215,N_9025);
xor U14279 (N_14279,N_11199,N_10376);
nor U14280 (N_14280,N_11170,N_10256);
and U14281 (N_14281,N_11469,N_11015);
or U14282 (N_14282,N_11654,N_9170);
nand U14283 (N_14283,N_9170,N_9733);
and U14284 (N_14284,N_10937,N_9272);
nor U14285 (N_14285,N_10026,N_11182);
nand U14286 (N_14286,N_10443,N_9246);
nand U14287 (N_14287,N_9186,N_11692);
or U14288 (N_14288,N_10063,N_10151);
nor U14289 (N_14289,N_11074,N_9047);
nor U14290 (N_14290,N_11786,N_11401);
and U14291 (N_14291,N_10447,N_11417);
and U14292 (N_14292,N_11284,N_10234);
xor U14293 (N_14293,N_11600,N_9240);
nand U14294 (N_14294,N_10822,N_11821);
nand U14295 (N_14295,N_11431,N_9589);
xnor U14296 (N_14296,N_9919,N_9720);
nand U14297 (N_14297,N_10832,N_11137);
nand U14298 (N_14298,N_11312,N_11038);
nand U14299 (N_14299,N_9845,N_10578);
nand U14300 (N_14300,N_9988,N_9274);
and U14301 (N_14301,N_11798,N_11398);
nor U14302 (N_14302,N_10775,N_11047);
nor U14303 (N_14303,N_10270,N_11384);
and U14304 (N_14304,N_10462,N_10452);
nor U14305 (N_14305,N_9296,N_11197);
xor U14306 (N_14306,N_10849,N_10248);
and U14307 (N_14307,N_9404,N_11469);
xor U14308 (N_14308,N_9664,N_9760);
xor U14309 (N_14309,N_10537,N_11340);
xnor U14310 (N_14310,N_10909,N_9602);
xor U14311 (N_14311,N_10873,N_11699);
and U14312 (N_14312,N_11638,N_9019);
nor U14313 (N_14313,N_9944,N_10269);
nand U14314 (N_14314,N_10871,N_11372);
or U14315 (N_14315,N_11303,N_10571);
nor U14316 (N_14316,N_10395,N_10363);
xor U14317 (N_14317,N_11780,N_11489);
and U14318 (N_14318,N_9167,N_11716);
or U14319 (N_14319,N_9458,N_11820);
nand U14320 (N_14320,N_9907,N_9376);
and U14321 (N_14321,N_9954,N_10759);
nor U14322 (N_14322,N_9187,N_11359);
nor U14323 (N_14323,N_9603,N_11603);
nand U14324 (N_14324,N_9079,N_9034);
and U14325 (N_14325,N_10462,N_10841);
or U14326 (N_14326,N_11068,N_10727);
or U14327 (N_14327,N_10667,N_9052);
xor U14328 (N_14328,N_10800,N_9615);
nand U14329 (N_14329,N_9828,N_9154);
xor U14330 (N_14330,N_10895,N_9891);
or U14331 (N_14331,N_11432,N_10342);
nand U14332 (N_14332,N_9128,N_10647);
or U14333 (N_14333,N_10291,N_11947);
or U14334 (N_14334,N_11867,N_11174);
nor U14335 (N_14335,N_10687,N_9948);
nor U14336 (N_14336,N_9382,N_10925);
and U14337 (N_14337,N_9422,N_11465);
or U14338 (N_14338,N_9601,N_11079);
or U14339 (N_14339,N_9086,N_9265);
and U14340 (N_14340,N_11371,N_10869);
nor U14341 (N_14341,N_10430,N_11721);
xnor U14342 (N_14342,N_11603,N_10987);
nand U14343 (N_14343,N_9638,N_11885);
and U14344 (N_14344,N_11298,N_10225);
nor U14345 (N_14345,N_10650,N_9222);
nand U14346 (N_14346,N_10280,N_10895);
nor U14347 (N_14347,N_10445,N_11979);
xnor U14348 (N_14348,N_9212,N_10398);
and U14349 (N_14349,N_11259,N_9317);
nand U14350 (N_14350,N_11970,N_10229);
nor U14351 (N_14351,N_9162,N_9793);
and U14352 (N_14352,N_9577,N_11622);
or U14353 (N_14353,N_9954,N_10064);
or U14354 (N_14354,N_10863,N_10913);
nand U14355 (N_14355,N_10351,N_9430);
and U14356 (N_14356,N_11570,N_10933);
xor U14357 (N_14357,N_11342,N_11271);
or U14358 (N_14358,N_10724,N_9751);
nand U14359 (N_14359,N_11127,N_10685);
nand U14360 (N_14360,N_10887,N_9100);
xnor U14361 (N_14361,N_9286,N_9023);
nor U14362 (N_14362,N_10016,N_11770);
nor U14363 (N_14363,N_9429,N_10349);
and U14364 (N_14364,N_9619,N_11908);
xor U14365 (N_14365,N_11340,N_9167);
xor U14366 (N_14366,N_10119,N_9344);
xnor U14367 (N_14367,N_10692,N_10068);
and U14368 (N_14368,N_10123,N_11660);
or U14369 (N_14369,N_11572,N_9504);
and U14370 (N_14370,N_11674,N_11896);
nor U14371 (N_14371,N_11964,N_9774);
or U14372 (N_14372,N_11431,N_10405);
nand U14373 (N_14373,N_9977,N_9085);
xnor U14374 (N_14374,N_11950,N_10791);
and U14375 (N_14375,N_9390,N_11865);
nor U14376 (N_14376,N_9516,N_11289);
nand U14377 (N_14377,N_10828,N_11191);
nand U14378 (N_14378,N_10921,N_9846);
nand U14379 (N_14379,N_10489,N_9655);
and U14380 (N_14380,N_11899,N_11747);
nand U14381 (N_14381,N_10535,N_11390);
nor U14382 (N_14382,N_9764,N_10240);
or U14383 (N_14383,N_11443,N_9717);
nand U14384 (N_14384,N_10309,N_10669);
or U14385 (N_14385,N_11252,N_10748);
xnor U14386 (N_14386,N_11306,N_11491);
and U14387 (N_14387,N_9876,N_11043);
xnor U14388 (N_14388,N_11857,N_10645);
nor U14389 (N_14389,N_11401,N_10199);
or U14390 (N_14390,N_11244,N_11231);
xnor U14391 (N_14391,N_11787,N_11019);
xor U14392 (N_14392,N_11231,N_9838);
and U14393 (N_14393,N_11018,N_11282);
nand U14394 (N_14394,N_10374,N_9533);
nor U14395 (N_14395,N_10382,N_10162);
or U14396 (N_14396,N_11586,N_11925);
nor U14397 (N_14397,N_10738,N_11647);
nand U14398 (N_14398,N_10761,N_9899);
nor U14399 (N_14399,N_9495,N_9592);
xor U14400 (N_14400,N_11057,N_9392);
xor U14401 (N_14401,N_9556,N_10340);
xnor U14402 (N_14402,N_11555,N_10865);
and U14403 (N_14403,N_9952,N_11797);
or U14404 (N_14404,N_10981,N_11681);
nor U14405 (N_14405,N_10746,N_11647);
nor U14406 (N_14406,N_9612,N_9877);
or U14407 (N_14407,N_9476,N_9774);
nand U14408 (N_14408,N_11835,N_11602);
nor U14409 (N_14409,N_10371,N_11883);
nor U14410 (N_14410,N_9866,N_9891);
xor U14411 (N_14411,N_10595,N_10918);
xnor U14412 (N_14412,N_11334,N_11997);
nor U14413 (N_14413,N_10745,N_10604);
nor U14414 (N_14414,N_11436,N_9649);
nor U14415 (N_14415,N_10166,N_9119);
nor U14416 (N_14416,N_11743,N_11745);
nor U14417 (N_14417,N_11197,N_10794);
xnor U14418 (N_14418,N_11452,N_9371);
nor U14419 (N_14419,N_9710,N_11583);
nand U14420 (N_14420,N_11768,N_11458);
or U14421 (N_14421,N_11595,N_11063);
nor U14422 (N_14422,N_10761,N_11961);
nor U14423 (N_14423,N_11919,N_9845);
or U14424 (N_14424,N_11316,N_10334);
xor U14425 (N_14425,N_10157,N_10957);
or U14426 (N_14426,N_10191,N_9126);
or U14427 (N_14427,N_11373,N_9726);
and U14428 (N_14428,N_10997,N_10498);
or U14429 (N_14429,N_10493,N_11098);
or U14430 (N_14430,N_11491,N_11671);
and U14431 (N_14431,N_10335,N_10167);
or U14432 (N_14432,N_11854,N_11536);
nand U14433 (N_14433,N_9024,N_10204);
nand U14434 (N_14434,N_9448,N_11913);
nor U14435 (N_14435,N_11074,N_10407);
xor U14436 (N_14436,N_11581,N_9160);
nor U14437 (N_14437,N_9686,N_11519);
and U14438 (N_14438,N_10520,N_11945);
or U14439 (N_14439,N_10507,N_10864);
nor U14440 (N_14440,N_10346,N_9413);
or U14441 (N_14441,N_10973,N_10283);
nand U14442 (N_14442,N_10272,N_10908);
or U14443 (N_14443,N_9271,N_11468);
or U14444 (N_14444,N_9719,N_9473);
xor U14445 (N_14445,N_11017,N_10552);
nor U14446 (N_14446,N_9901,N_11338);
or U14447 (N_14447,N_10427,N_10467);
or U14448 (N_14448,N_9997,N_10851);
nor U14449 (N_14449,N_9090,N_11269);
nand U14450 (N_14450,N_10403,N_11938);
and U14451 (N_14451,N_11265,N_9951);
xnor U14452 (N_14452,N_10186,N_9377);
or U14453 (N_14453,N_11327,N_10599);
and U14454 (N_14454,N_10854,N_11587);
and U14455 (N_14455,N_10004,N_9637);
and U14456 (N_14456,N_10671,N_11233);
xnor U14457 (N_14457,N_10263,N_11628);
nor U14458 (N_14458,N_10047,N_10313);
xnor U14459 (N_14459,N_10330,N_11556);
nand U14460 (N_14460,N_9199,N_9808);
nor U14461 (N_14461,N_10528,N_10050);
nand U14462 (N_14462,N_10283,N_11224);
and U14463 (N_14463,N_11229,N_9206);
and U14464 (N_14464,N_11781,N_9896);
or U14465 (N_14465,N_11336,N_11656);
and U14466 (N_14466,N_11411,N_11779);
nand U14467 (N_14467,N_11321,N_9477);
and U14468 (N_14468,N_11509,N_9450);
and U14469 (N_14469,N_11591,N_10855);
or U14470 (N_14470,N_10053,N_9188);
nand U14471 (N_14471,N_10155,N_9973);
and U14472 (N_14472,N_9451,N_11926);
xor U14473 (N_14473,N_10136,N_10206);
and U14474 (N_14474,N_10434,N_11781);
or U14475 (N_14475,N_9431,N_10825);
nand U14476 (N_14476,N_11796,N_11675);
nor U14477 (N_14477,N_10235,N_11113);
nor U14478 (N_14478,N_11156,N_10563);
xor U14479 (N_14479,N_10950,N_10845);
or U14480 (N_14480,N_10561,N_11557);
nor U14481 (N_14481,N_10868,N_11002);
and U14482 (N_14482,N_9105,N_11566);
xor U14483 (N_14483,N_9907,N_10610);
and U14484 (N_14484,N_9918,N_9216);
nand U14485 (N_14485,N_9304,N_11837);
and U14486 (N_14486,N_9962,N_9372);
or U14487 (N_14487,N_9942,N_9059);
or U14488 (N_14488,N_11616,N_10855);
nor U14489 (N_14489,N_11697,N_10891);
xor U14490 (N_14490,N_11245,N_9805);
xnor U14491 (N_14491,N_11296,N_10382);
nand U14492 (N_14492,N_10904,N_10636);
nand U14493 (N_14493,N_11057,N_9085);
xor U14494 (N_14494,N_11779,N_11334);
nand U14495 (N_14495,N_11670,N_10056);
nand U14496 (N_14496,N_10853,N_10641);
xor U14497 (N_14497,N_9338,N_10780);
nand U14498 (N_14498,N_10605,N_11021);
or U14499 (N_14499,N_9044,N_10765);
nand U14500 (N_14500,N_11465,N_11012);
xnor U14501 (N_14501,N_9748,N_10851);
nor U14502 (N_14502,N_9354,N_9100);
nand U14503 (N_14503,N_10984,N_11851);
and U14504 (N_14504,N_11715,N_10289);
xnor U14505 (N_14505,N_10139,N_10335);
or U14506 (N_14506,N_10441,N_10351);
nor U14507 (N_14507,N_10260,N_11578);
nand U14508 (N_14508,N_10505,N_11747);
xor U14509 (N_14509,N_11228,N_9970);
and U14510 (N_14510,N_10013,N_10188);
nand U14511 (N_14511,N_10816,N_11185);
xnor U14512 (N_14512,N_9299,N_11265);
or U14513 (N_14513,N_9568,N_11824);
and U14514 (N_14514,N_10098,N_9466);
nand U14515 (N_14515,N_9899,N_9457);
nor U14516 (N_14516,N_11745,N_10537);
or U14517 (N_14517,N_11778,N_10360);
or U14518 (N_14518,N_9711,N_9727);
nor U14519 (N_14519,N_11656,N_9625);
xor U14520 (N_14520,N_11271,N_9040);
nor U14521 (N_14521,N_9439,N_11796);
xnor U14522 (N_14522,N_9533,N_10524);
nand U14523 (N_14523,N_10226,N_9749);
nor U14524 (N_14524,N_11386,N_10525);
or U14525 (N_14525,N_10898,N_9466);
or U14526 (N_14526,N_10453,N_9151);
nor U14527 (N_14527,N_11661,N_11005);
nor U14528 (N_14528,N_10376,N_9944);
or U14529 (N_14529,N_11327,N_10182);
or U14530 (N_14530,N_10023,N_11219);
and U14531 (N_14531,N_11389,N_11088);
nand U14532 (N_14532,N_10001,N_10324);
nand U14533 (N_14533,N_9066,N_9619);
nand U14534 (N_14534,N_10275,N_11165);
nor U14535 (N_14535,N_9874,N_10658);
xnor U14536 (N_14536,N_11125,N_10506);
nor U14537 (N_14537,N_10990,N_9619);
and U14538 (N_14538,N_9615,N_10060);
or U14539 (N_14539,N_10499,N_9861);
and U14540 (N_14540,N_10652,N_11325);
nand U14541 (N_14541,N_11831,N_9219);
xnor U14542 (N_14542,N_9142,N_9415);
or U14543 (N_14543,N_10634,N_9224);
nor U14544 (N_14544,N_9540,N_11534);
nand U14545 (N_14545,N_10977,N_11300);
xnor U14546 (N_14546,N_10150,N_11514);
nor U14547 (N_14547,N_9949,N_10219);
nand U14548 (N_14548,N_10013,N_11429);
or U14549 (N_14549,N_10588,N_10231);
nor U14550 (N_14550,N_10519,N_10328);
or U14551 (N_14551,N_11180,N_10073);
nor U14552 (N_14552,N_10543,N_9023);
xnor U14553 (N_14553,N_10292,N_11058);
nand U14554 (N_14554,N_9534,N_10810);
or U14555 (N_14555,N_9426,N_9302);
and U14556 (N_14556,N_11850,N_10724);
and U14557 (N_14557,N_9415,N_11206);
or U14558 (N_14558,N_9083,N_9817);
nor U14559 (N_14559,N_10697,N_9721);
nand U14560 (N_14560,N_9958,N_11950);
nor U14561 (N_14561,N_9038,N_10776);
xnor U14562 (N_14562,N_11430,N_10138);
nor U14563 (N_14563,N_11196,N_11779);
and U14564 (N_14564,N_10731,N_10129);
xnor U14565 (N_14565,N_9809,N_9561);
xnor U14566 (N_14566,N_11280,N_9777);
or U14567 (N_14567,N_11151,N_11413);
xnor U14568 (N_14568,N_11979,N_9208);
nand U14569 (N_14569,N_10967,N_10226);
nor U14570 (N_14570,N_11109,N_10749);
xor U14571 (N_14571,N_11589,N_9420);
and U14572 (N_14572,N_10173,N_11659);
or U14573 (N_14573,N_10717,N_11555);
or U14574 (N_14574,N_11659,N_9377);
nor U14575 (N_14575,N_10706,N_9691);
or U14576 (N_14576,N_10274,N_10421);
and U14577 (N_14577,N_9233,N_10210);
nand U14578 (N_14578,N_11155,N_9192);
xor U14579 (N_14579,N_10750,N_9524);
or U14580 (N_14580,N_9503,N_9741);
and U14581 (N_14581,N_9320,N_10792);
xor U14582 (N_14582,N_9958,N_9528);
nor U14583 (N_14583,N_9547,N_11726);
nor U14584 (N_14584,N_10519,N_10584);
nand U14585 (N_14585,N_10065,N_9927);
or U14586 (N_14586,N_10167,N_9375);
nor U14587 (N_14587,N_10704,N_11617);
or U14588 (N_14588,N_10399,N_11753);
and U14589 (N_14589,N_9961,N_10133);
nor U14590 (N_14590,N_11615,N_11330);
nand U14591 (N_14591,N_10160,N_11442);
or U14592 (N_14592,N_11509,N_9602);
or U14593 (N_14593,N_10178,N_11572);
xor U14594 (N_14594,N_10910,N_9803);
and U14595 (N_14595,N_11577,N_11342);
xnor U14596 (N_14596,N_11609,N_10019);
or U14597 (N_14597,N_10944,N_9062);
and U14598 (N_14598,N_10207,N_11363);
xnor U14599 (N_14599,N_10784,N_11701);
nor U14600 (N_14600,N_10750,N_9885);
and U14601 (N_14601,N_9649,N_11802);
or U14602 (N_14602,N_11504,N_9232);
nor U14603 (N_14603,N_11522,N_10938);
and U14604 (N_14604,N_9495,N_9460);
and U14605 (N_14605,N_10247,N_11739);
and U14606 (N_14606,N_10571,N_9163);
nor U14607 (N_14607,N_10103,N_10557);
nor U14608 (N_14608,N_11357,N_9414);
nor U14609 (N_14609,N_10842,N_9109);
or U14610 (N_14610,N_9844,N_11085);
nor U14611 (N_14611,N_11198,N_10632);
nor U14612 (N_14612,N_10687,N_9202);
and U14613 (N_14613,N_9320,N_10870);
and U14614 (N_14614,N_9415,N_9762);
and U14615 (N_14615,N_11783,N_9645);
and U14616 (N_14616,N_10235,N_11026);
nor U14617 (N_14617,N_10547,N_10790);
nand U14618 (N_14618,N_10650,N_9536);
nand U14619 (N_14619,N_9058,N_9214);
nor U14620 (N_14620,N_9956,N_11286);
nor U14621 (N_14621,N_9888,N_11239);
and U14622 (N_14622,N_10255,N_9650);
and U14623 (N_14623,N_10354,N_11825);
and U14624 (N_14624,N_9026,N_9981);
and U14625 (N_14625,N_11189,N_11092);
nand U14626 (N_14626,N_10581,N_9281);
nor U14627 (N_14627,N_9525,N_11852);
or U14628 (N_14628,N_10353,N_11564);
or U14629 (N_14629,N_11996,N_9474);
nor U14630 (N_14630,N_9062,N_11607);
nor U14631 (N_14631,N_10938,N_9126);
or U14632 (N_14632,N_10291,N_11805);
nand U14633 (N_14633,N_11809,N_10273);
xnor U14634 (N_14634,N_10422,N_11529);
xor U14635 (N_14635,N_9975,N_10372);
or U14636 (N_14636,N_9529,N_11817);
nor U14637 (N_14637,N_10556,N_11841);
or U14638 (N_14638,N_11390,N_10419);
or U14639 (N_14639,N_10581,N_11997);
nand U14640 (N_14640,N_9705,N_9308);
nand U14641 (N_14641,N_9499,N_10551);
nand U14642 (N_14642,N_11409,N_11057);
or U14643 (N_14643,N_11923,N_9316);
and U14644 (N_14644,N_11369,N_9891);
nand U14645 (N_14645,N_9083,N_11896);
nor U14646 (N_14646,N_11806,N_11333);
or U14647 (N_14647,N_9645,N_10211);
and U14648 (N_14648,N_9097,N_9557);
xor U14649 (N_14649,N_11266,N_10622);
or U14650 (N_14650,N_10312,N_11422);
or U14651 (N_14651,N_10270,N_10576);
or U14652 (N_14652,N_11890,N_10683);
or U14653 (N_14653,N_9488,N_11930);
and U14654 (N_14654,N_10027,N_10510);
and U14655 (N_14655,N_9644,N_10930);
nor U14656 (N_14656,N_11854,N_10579);
and U14657 (N_14657,N_10079,N_10478);
or U14658 (N_14658,N_11611,N_11788);
and U14659 (N_14659,N_11299,N_11456);
nor U14660 (N_14660,N_9898,N_10836);
nand U14661 (N_14661,N_11371,N_11768);
or U14662 (N_14662,N_11057,N_11821);
or U14663 (N_14663,N_9443,N_11057);
and U14664 (N_14664,N_9378,N_10717);
or U14665 (N_14665,N_10585,N_9536);
and U14666 (N_14666,N_11891,N_10787);
nor U14667 (N_14667,N_10826,N_11855);
or U14668 (N_14668,N_9322,N_11198);
nor U14669 (N_14669,N_9974,N_10962);
nand U14670 (N_14670,N_11930,N_10589);
nand U14671 (N_14671,N_11300,N_11661);
nor U14672 (N_14672,N_10484,N_11092);
xor U14673 (N_14673,N_10211,N_11331);
nor U14674 (N_14674,N_10012,N_10923);
nand U14675 (N_14675,N_9173,N_11989);
xor U14676 (N_14676,N_10253,N_10667);
and U14677 (N_14677,N_10824,N_11894);
nor U14678 (N_14678,N_10707,N_9532);
nand U14679 (N_14679,N_10431,N_10110);
and U14680 (N_14680,N_9072,N_10770);
xnor U14681 (N_14681,N_11899,N_9668);
nand U14682 (N_14682,N_10883,N_11517);
xor U14683 (N_14683,N_11200,N_11879);
and U14684 (N_14684,N_10607,N_11205);
or U14685 (N_14685,N_11512,N_10220);
nor U14686 (N_14686,N_9887,N_11298);
and U14687 (N_14687,N_10560,N_9845);
nand U14688 (N_14688,N_11543,N_10689);
xor U14689 (N_14689,N_11245,N_11136);
or U14690 (N_14690,N_10070,N_9411);
nor U14691 (N_14691,N_10563,N_9852);
nor U14692 (N_14692,N_9079,N_11958);
xnor U14693 (N_14693,N_10677,N_10456);
xnor U14694 (N_14694,N_11806,N_10347);
or U14695 (N_14695,N_11119,N_9805);
or U14696 (N_14696,N_9628,N_11394);
or U14697 (N_14697,N_11957,N_10245);
nor U14698 (N_14698,N_11438,N_11536);
nand U14699 (N_14699,N_10832,N_10094);
or U14700 (N_14700,N_9501,N_11181);
nand U14701 (N_14701,N_10299,N_10801);
nor U14702 (N_14702,N_11977,N_11021);
nor U14703 (N_14703,N_9662,N_11837);
xor U14704 (N_14704,N_9924,N_9000);
nand U14705 (N_14705,N_11682,N_9851);
and U14706 (N_14706,N_9308,N_9564);
nand U14707 (N_14707,N_11758,N_9429);
xnor U14708 (N_14708,N_10996,N_9757);
and U14709 (N_14709,N_11928,N_10850);
or U14710 (N_14710,N_10702,N_10301);
xnor U14711 (N_14711,N_9371,N_10628);
or U14712 (N_14712,N_9375,N_10596);
or U14713 (N_14713,N_11195,N_10286);
or U14714 (N_14714,N_11345,N_11787);
nor U14715 (N_14715,N_10156,N_9851);
nor U14716 (N_14716,N_9844,N_11810);
xnor U14717 (N_14717,N_11373,N_10804);
or U14718 (N_14718,N_9371,N_10702);
nor U14719 (N_14719,N_11124,N_10017);
xnor U14720 (N_14720,N_9491,N_10687);
nor U14721 (N_14721,N_10685,N_9423);
and U14722 (N_14722,N_9928,N_9661);
xnor U14723 (N_14723,N_9877,N_11891);
or U14724 (N_14724,N_10811,N_11576);
nand U14725 (N_14725,N_9686,N_9789);
or U14726 (N_14726,N_9144,N_9119);
nand U14727 (N_14727,N_11623,N_11870);
and U14728 (N_14728,N_11761,N_9424);
xnor U14729 (N_14729,N_11307,N_9560);
or U14730 (N_14730,N_11903,N_9289);
or U14731 (N_14731,N_9254,N_10912);
nand U14732 (N_14732,N_9958,N_9231);
nor U14733 (N_14733,N_10815,N_11596);
xor U14734 (N_14734,N_10553,N_10843);
nand U14735 (N_14735,N_9923,N_10605);
nor U14736 (N_14736,N_10967,N_10750);
nor U14737 (N_14737,N_10834,N_11105);
nand U14738 (N_14738,N_9243,N_9100);
and U14739 (N_14739,N_11230,N_9131);
xnor U14740 (N_14740,N_9455,N_9410);
nor U14741 (N_14741,N_11444,N_11833);
or U14742 (N_14742,N_11454,N_11047);
xor U14743 (N_14743,N_9392,N_11749);
xor U14744 (N_14744,N_10468,N_10747);
xor U14745 (N_14745,N_10605,N_11710);
or U14746 (N_14746,N_9394,N_9145);
nor U14747 (N_14747,N_10830,N_9024);
nor U14748 (N_14748,N_11819,N_11052);
xnor U14749 (N_14749,N_9808,N_9459);
and U14750 (N_14750,N_10202,N_10915);
nand U14751 (N_14751,N_11506,N_9346);
or U14752 (N_14752,N_9605,N_10694);
nor U14753 (N_14753,N_9112,N_11549);
nor U14754 (N_14754,N_10442,N_11420);
nand U14755 (N_14755,N_9262,N_11114);
or U14756 (N_14756,N_11853,N_10116);
or U14757 (N_14757,N_10658,N_10730);
xor U14758 (N_14758,N_9203,N_11981);
and U14759 (N_14759,N_9335,N_11017);
xor U14760 (N_14760,N_10539,N_9718);
nor U14761 (N_14761,N_9833,N_11763);
nor U14762 (N_14762,N_10105,N_9165);
and U14763 (N_14763,N_9334,N_9272);
nand U14764 (N_14764,N_9794,N_10397);
and U14765 (N_14765,N_11668,N_11817);
nand U14766 (N_14766,N_9681,N_10019);
xnor U14767 (N_14767,N_11009,N_10618);
nor U14768 (N_14768,N_10239,N_9161);
xor U14769 (N_14769,N_11977,N_9524);
nand U14770 (N_14770,N_10642,N_11946);
nand U14771 (N_14771,N_11739,N_9476);
or U14772 (N_14772,N_11123,N_11360);
nor U14773 (N_14773,N_9452,N_11560);
and U14774 (N_14774,N_10103,N_10185);
and U14775 (N_14775,N_10584,N_9476);
xor U14776 (N_14776,N_9405,N_11362);
or U14777 (N_14777,N_9455,N_11887);
and U14778 (N_14778,N_10679,N_9013);
nand U14779 (N_14779,N_11368,N_10968);
xor U14780 (N_14780,N_11472,N_9036);
xnor U14781 (N_14781,N_11039,N_11091);
or U14782 (N_14782,N_11788,N_11123);
or U14783 (N_14783,N_10011,N_11608);
or U14784 (N_14784,N_11687,N_9996);
nand U14785 (N_14785,N_11715,N_11563);
or U14786 (N_14786,N_11294,N_10844);
xor U14787 (N_14787,N_9280,N_11479);
nor U14788 (N_14788,N_9456,N_11624);
nor U14789 (N_14789,N_9353,N_9887);
xnor U14790 (N_14790,N_10857,N_11013);
xor U14791 (N_14791,N_10534,N_11809);
and U14792 (N_14792,N_9319,N_9321);
xnor U14793 (N_14793,N_9408,N_11488);
nand U14794 (N_14794,N_11122,N_11254);
xnor U14795 (N_14795,N_9009,N_11736);
and U14796 (N_14796,N_10613,N_9726);
xor U14797 (N_14797,N_11383,N_11385);
xnor U14798 (N_14798,N_9828,N_9231);
nor U14799 (N_14799,N_11335,N_11735);
nor U14800 (N_14800,N_11759,N_11029);
nand U14801 (N_14801,N_11133,N_10369);
nand U14802 (N_14802,N_11619,N_10757);
nor U14803 (N_14803,N_11873,N_11226);
nand U14804 (N_14804,N_9227,N_9394);
and U14805 (N_14805,N_9521,N_11830);
nor U14806 (N_14806,N_9470,N_10073);
nand U14807 (N_14807,N_11717,N_11472);
nand U14808 (N_14808,N_11171,N_10744);
and U14809 (N_14809,N_10823,N_10108);
xnor U14810 (N_14810,N_9094,N_11952);
or U14811 (N_14811,N_10389,N_11434);
nor U14812 (N_14812,N_9975,N_9190);
xor U14813 (N_14813,N_9316,N_9874);
nor U14814 (N_14814,N_10453,N_11074);
and U14815 (N_14815,N_9413,N_10488);
nor U14816 (N_14816,N_9853,N_11103);
and U14817 (N_14817,N_11089,N_10204);
xnor U14818 (N_14818,N_9399,N_10483);
nor U14819 (N_14819,N_10242,N_10648);
xnor U14820 (N_14820,N_10016,N_10231);
nor U14821 (N_14821,N_10367,N_10813);
nor U14822 (N_14822,N_11188,N_11466);
or U14823 (N_14823,N_10261,N_11146);
or U14824 (N_14824,N_9267,N_11804);
or U14825 (N_14825,N_11933,N_9770);
and U14826 (N_14826,N_9876,N_11786);
nor U14827 (N_14827,N_9147,N_10706);
nor U14828 (N_14828,N_11021,N_10257);
nor U14829 (N_14829,N_9015,N_10390);
and U14830 (N_14830,N_11269,N_9777);
xor U14831 (N_14831,N_11780,N_10696);
xor U14832 (N_14832,N_10442,N_10656);
or U14833 (N_14833,N_11400,N_9983);
or U14834 (N_14834,N_10081,N_11018);
or U14835 (N_14835,N_9615,N_11026);
and U14836 (N_14836,N_9314,N_11761);
and U14837 (N_14837,N_9274,N_10985);
and U14838 (N_14838,N_9237,N_10640);
nand U14839 (N_14839,N_9474,N_10633);
xnor U14840 (N_14840,N_9103,N_11936);
nor U14841 (N_14841,N_9094,N_11097);
xnor U14842 (N_14842,N_11965,N_11952);
nand U14843 (N_14843,N_10514,N_11942);
nor U14844 (N_14844,N_10125,N_10257);
or U14845 (N_14845,N_9856,N_9759);
nand U14846 (N_14846,N_9501,N_10286);
nand U14847 (N_14847,N_11721,N_10407);
xnor U14848 (N_14848,N_11264,N_9699);
and U14849 (N_14849,N_9673,N_10486);
nand U14850 (N_14850,N_10101,N_10679);
or U14851 (N_14851,N_9031,N_10496);
nand U14852 (N_14852,N_11006,N_11324);
and U14853 (N_14853,N_9497,N_9105);
nand U14854 (N_14854,N_9776,N_9685);
nor U14855 (N_14855,N_9440,N_9204);
or U14856 (N_14856,N_11916,N_10399);
nand U14857 (N_14857,N_9313,N_11652);
nor U14858 (N_14858,N_10966,N_9202);
nor U14859 (N_14859,N_10501,N_9458);
or U14860 (N_14860,N_11529,N_9941);
xnor U14861 (N_14861,N_11867,N_9209);
or U14862 (N_14862,N_10963,N_10714);
xnor U14863 (N_14863,N_9370,N_10566);
and U14864 (N_14864,N_9013,N_9151);
nand U14865 (N_14865,N_11461,N_9149);
nor U14866 (N_14866,N_11027,N_11089);
and U14867 (N_14867,N_11372,N_9193);
xnor U14868 (N_14868,N_10245,N_10022);
nand U14869 (N_14869,N_11998,N_10746);
nor U14870 (N_14870,N_9719,N_9488);
nor U14871 (N_14871,N_10235,N_10526);
xnor U14872 (N_14872,N_10751,N_9354);
nand U14873 (N_14873,N_10476,N_11507);
and U14874 (N_14874,N_10320,N_10254);
nor U14875 (N_14875,N_9492,N_10641);
and U14876 (N_14876,N_9742,N_10698);
xor U14877 (N_14877,N_11045,N_11151);
nand U14878 (N_14878,N_9803,N_11385);
or U14879 (N_14879,N_9109,N_10855);
nand U14880 (N_14880,N_9791,N_11873);
or U14881 (N_14881,N_9812,N_10709);
nand U14882 (N_14882,N_10218,N_10424);
or U14883 (N_14883,N_9351,N_11128);
xnor U14884 (N_14884,N_11501,N_11408);
nand U14885 (N_14885,N_9502,N_10133);
xor U14886 (N_14886,N_11394,N_10364);
nor U14887 (N_14887,N_10722,N_11021);
nand U14888 (N_14888,N_11373,N_10029);
or U14889 (N_14889,N_9894,N_9796);
or U14890 (N_14890,N_9158,N_11971);
xnor U14891 (N_14891,N_11191,N_10531);
or U14892 (N_14892,N_9983,N_11676);
nand U14893 (N_14893,N_9548,N_11901);
and U14894 (N_14894,N_11576,N_9724);
and U14895 (N_14895,N_10730,N_10556);
xnor U14896 (N_14896,N_9991,N_9239);
and U14897 (N_14897,N_11328,N_9749);
xor U14898 (N_14898,N_9281,N_10728);
xor U14899 (N_14899,N_11963,N_11737);
and U14900 (N_14900,N_11839,N_11149);
or U14901 (N_14901,N_9864,N_9613);
and U14902 (N_14902,N_9749,N_10407);
or U14903 (N_14903,N_11059,N_9637);
or U14904 (N_14904,N_10536,N_10426);
nor U14905 (N_14905,N_9056,N_10457);
xnor U14906 (N_14906,N_9756,N_10938);
and U14907 (N_14907,N_11882,N_11602);
and U14908 (N_14908,N_10120,N_11452);
nand U14909 (N_14909,N_10844,N_10565);
nor U14910 (N_14910,N_11759,N_11003);
nand U14911 (N_14911,N_9006,N_10723);
xnor U14912 (N_14912,N_11917,N_11745);
nand U14913 (N_14913,N_9548,N_9367);
nand U14914 (N_14914,N_10626,N_9738);
and U14915 (N_14915,N_10970,N_9162);
nand U14916 (N_14916,N_11743,N_10925);
xnor U14917 (N_14917,N_11056,N_9478);
xnor U14918 (N_14918,N_9589,N_11506);
nand U14919 (N_14919,N_9907,N_9863);
nor U14920 (N_14920,N_9587,N_11338);
xor U14921 (N_14921,N_10768,N_9448);
nor U14922 (N_14922,N_11276,N_10722);
nand U14923 (N_14923,N_11257,N_9778);
nor U14924 (N_14924,N_9249,N_11850);
nor U14925 (N_14925,N_10974,N_10459);
and U14926 (N_14926,N_11251,N_9427);
nand U14927 (N_14927,N_11833,N_10481);
nor U14928 (N_14928,N_10837,N_10262);
xnor U14929 (N_14929,N_10903,N_9750);
or U14930 (N_14930,N_10198,N_11433);
nand U14931 (N_14931,N_11253,N_10708);
or U14932 (N_14932,N_9694,N_11036);
nor U14933 (N_14933,N_9517,N_11132);
or U14934 (N_14934,N_11236,N_9981);
xnor U14935 (N_14935,N_10355,N_11643);
and U14936 (N_14936,N_10398,N_10069);
nor U14937 (N_14937,N_10392,N_11730);
or U14938 (N_14938,N_11002,N_9579);
nor U14939 (N_14939,N_9127,N_9599);
and U14940 (N_14940,N_9719,N_11526);
xor U14941 (N_14941,N_10707,N_11895);
nor U14942 (N_14942,N_11628,N_11106);
nor U14943 (N_14943,N_9550,N_11816);
nor U14944 (N_14944,N_9598,N_10981);
nor U14945 (N_14945,N_10052,N_9779);
nor U14946 (N_14946,N_11729,N_11683);
or U14947 (N_14947,N_9008,N_10251);
and U14948 (N_14948,N_9221,N_9913);
nand U14949 (N_14949,N_11882,N_10091);
nand U14950 (N_14950,N_9323,N_10527);
or U14951 (N_14951,N_11505,N_9077);
xor U14952 (N_14952,N_10330,N_11474);
nand U14953 (N_14953,N_11699,N_11234);
nand U14954 (N_14954,N_11691,N_10845);
nor U14955 (N_14955,N_10793,N_11089);
nand U14956 (N_14956,N_10715,N_10523);
xor U14957 (N_14957,N_11283,N_9625);
xnor U14958 (N_14958,N_9106,N_10639);
nor U14959 (N_14959,N_9947,N_11874);
or U14960 (N_14960,N_9830,N_11237);
and U14961 (N_14961,N_11829,N_11577);
xnor U14962 (N_14962,N_11526,N_10535);
xnor U14963 (N_14963,N_9904,N_11670);
nand U14964 (N_14964,N_11407,N_11757);
and U14965 (N_14965,N_9438,N_10312);
and U14966 (N_14966,N_9447,N_9369);
nor U14967 (N_14967,N_9911,N_10131);
nand U14968 (N_14968,N_11365,N_11781);
nor U14969 (N_14969,N_11448,N_11357);
xnor U14970 (N_14970,N_10893,N_10070);
xor U14971 (N_14971,N_10593,N_9452);
or U14972 (N_14972,N_10558,N_9536);
or U14973 (N_14973,N_11627,N_11766);
and U14974 (N_14974,N_11751,N_11070);
nor U14975 (N_14975,N_9518,N_10554);
or U14976 (N_14976,N_9551,N_10305);
and U14977 (N_14977,N_11772,N_9709);
nor U14978 (N_14978,N_9682,N_11958);
nand U14979 (N_14979,N_10888,N_9024);
xnor U14980 (N_14980,N_10274,N_9026);
nor U14981 (N_14981,N_10631,N_10355);
or U14982 (N_14982,N_10671,N_10336);
or U14983 (N_14983,N_9515,N_9913);
nor U14984 (N_14984,N_9267,N_10174);
nand U14985 (N_14985,N_10455,N_9091);
nand U14986 (N_14986,N_10805,N_11829);
or U14987 (N_14987,N_11383,N_9468);
or U14988 (N_14988,N_9038,N_11715);
nor U14989 (N_14989,N_11710,N_11979);
nor U14990 (N_14990,N_10657,N_10658);
nand U14991 (N_14991,N_11343,N_9476);
nand U14992 (N_14992,N_11978,N_11848);
nand U14993 (N_14993,N_10904,N_9336);
xor U14994 (N_14994,N_10718,N_10281);
or U14995 (N_14995,N_9001,N_9389);
and U14996 (N_14996,N_9957,N_10063);
xnor U14997 (N_14997,N_9866,N_9807);
nor U14998 (N_14998,N_9002,N_9625);
nand U14999 (N_14999,N_10156,N_9794);
nand U15000 (N_15000,N_12903,N_12748);
xnor U15001 (N_15001,N_14862,N_12594);
or U15002 (N_15002,N_13837,N_14612);
or U15003 (N_15003,N_13714,N_13259);
xnor U15004 (N_15004,N_12252,N_13364);
and U15005 (N_15005,N_14257,N_14891);
nor U15006 (N_15006,N_12240,N_14263);
nor U15007 (N_15007,N_14213,N_13264);
or U15008 (N_15008,N_12328,N_14667);
nand U15009 (N_15009,N_13801,N_13836);
nand U15010 (N_15010,N_14985,N_14426);
nand U15011 (N_15011,N_13766,N_13570);
xnor U15012 (N_15012,N_14135,N_14723);
and U15013 (N_15013,N_13939,N_12869);
or U15014 (N_15014,N_14669,N_14077);
or U15015 (N_15015,N_14227,N_12637);
nand U15016 (N_15016,N_13527,N_14046);
xnor U15017 (N_15017,N_12756,N_12099);
nand U15018 (N_15018,N_12282,N_12368);
xnor U15019 (N_15019,N_14693,N_12627);
nand U15020 (N_15020,N_14228,N_13471);
xor U15021 (N_15021,N_14100,N_14501);
nand U15022 (N_15022,N_13686,N_14236);
nand U15023 (N_15023,N_12812,N_14929);
xnor U15024 (N_15024,N_12256,N_12035);
nor U15025 (N_15025,N_13752,N_14758);
nor U15026 (N_15026,N_14704,N_14418);
and U15027 (N_15027,N_12417,N_12208);
or U15028 (N_15028,N_14342,N_14869);
nand U15029 (N_15029,N_12217,N_14843);
nor U15030 (N_15030,N_13248,N_13954);
nand U15031 (N_15031,N_12411,N_12771);
xnor U15032 (N_15032,N_13340,N_14166);
and U15033 (N_15033,N_14247,N_13228);
xnor U15034 (N_15034,N_12286,N_13738);
and U15035 (N_15035,N_12258,N_12171);
nand U15036 (N_15036,N_13217,N_14207);
nand U15037 (N_15037,N_12062,N_12326);
or U15038 (N_15038,N_13549,N_12041);
or U15039 (N_15039,N_14543,N_13508);
nor U15040 (N_15040,N_12259,N_13150);
nand U15041 (N_15041,N_14975,N_13723);
nand U15042 (N_15042,N_14958,N_14103);
nand U15043 (N_15043,N_12969,N_13335);
or U15044 (N_15044,N_14281,N_14716);
nor U15045 (N_15045,N_13467,N_14494);
or U15046 (N_15046,N_13831,N_14392);
and U15047 (N_15047,N_13557,N_14846);
and U15048 (N_15048,N_13754,N_14686);
nand U15049 (N_15049,N_14559,N_13804);
xnor U15050 (N_15050,N_13692,N_13045);
xor U15051 (N_15051,N_14523,N_13143);
nand U15052 (N_15052,N_12151,N_12105);
and U15053 (N_15053,N_14911,N_12835);
nor U15054 (N_15054,N_14206,N_14607);
nand U15055 (N_15055,N_13255,N_12705);
nand U15056 (N_15056,N_13332,N_14382);
nand U15057 (N_15057,N_12810,N_14920);
and U15058 (N_15058,N_14783,N_13448);
or U15059 (N_15059,N_14199,N_14941);
xnor U15060 (N_15060,N_14503,N_13748);
or U15061 (N_15061,N_13936,N_14267);
and U15062 (N_15062,N_13604,N_12453);
xnor U15063 (N_15063,N_14456,N_13390);
nor U15064 (N_15064,N_13005,N_12264);
xor U15065 (N_15065,N_12459,N_12135);
or U15066 (N_15066,N_14613,N_12746);
or U15067 (N_15067,N_12842,N_13345);
nand U15068 (N_15068,N_14584,N_13652);
nand U15069 (N_15069,N_14972,N_14893);
or U15070 (N_15070,N_13744,N_13091);
and U15071 (N_15071,N_12095,N_14015);
nand U15072 (N_15072,N_13053,N_12593);
or U15073 (N_15073,N_14960,N_13629);
and U15074 (N_15074,N_14080,N_14966);
or U15075 (N_15075,N_12462,N_14579);
nand U15076 (N_15076,N_12441,N_13930);
xnor U15077 (N_15077,N_12938,N_13779);
or U15078 (N_15078,N_14362,N_12935);
xor U15079 (N_15079,N_13759,N_13132);
and U15080 (N_15080,N_13068,N_13239);
nor U15081 (N_15081,N_13808,N_14993);
and U15082 (N_15082,N_14526,N_13518);
or U15083 (N_15083,N_14041,N_13224);
or U15084 (N_15084,N_12031,N_14626);
nor U15085 (N_15085,N_12996,N_12981);
nor U15086 (N_15086,N_14666,N_14999);
or U15087 (N_15087,N_13167,N_13061);
and U15088 (N_15088,N_12028,N_13378);
nand U15089 (N_15089,N_12890,N_12340);
nand U15090 (N_15090,N_14379,N_12700);
and U15091 (N_15091,N_12821,N_12855);
nor U15092 (N_15092,N_12472,N_12854);
or U15093 (N_15093,N_12689,N_12487);
and U15094 (N_15094,N_14573,N_14443);
nand U15095 (N_15095,N_14630,N_14817);
xnor U15096 (N_15096,N_12691,N_12894);
or U15097 (N_15097,N_13070,N_13875);
or U15098 (N_15098,N_12735,N_13489);
and U15099 (N_15099,N_14542,N_13584);
and U15100 (N_15100,N_12281,N_13011);
nor U15101 (N_15101,N_12815,N_14295);
xor U15102 (N_15102,N_12589,N_12744);
or U15103 (N_15103,N_13298,N_13024);
xor U15104 (N_15104,N_13788,N_12428);
or U15105 (N_15105,N_14979,N_13796);
nor U15106 (N_15106,N_12829,N_14827);
or U15107 (N_15107,N_14126,N_14462);
xor U15108 (N_15108,N_14210,N_12361);
nor U15109 (N_15109,N_13777,N_14356);
and U15110 (N_15110,N_14971,N_12565);
nor U15111 (N_15111,N_13325,N_13092);
or U15112 (N_15112,N_13182,N_13493);
xnor U15113 (N_15113,N_13900,N_13140);
nand U15114 (N_15114,N_13880,N_12858);
and U15115 (N_15115,N_12283,N_14824);
or U15116 (N_15116,N_14685,N_13025);
or U15117 (N_15117,N_12685,N_13755);
nand U15118 (N_15118,N_12203,N_14388);
and U15119 (N_15119,N_12498,N_14528);
or U15120 (N_15120,N_14315,N_13855);
or U15121 (N_15121,N_13286,N_14132);
and U15122 (N_15122,N_13426,N_12864);
nand U15123 (N_15123,N_12574,N_12430);
and U15124 (N_15124,N_13680,N_14209);
nand U15125 (N_15125,N_14937,N_13594);
nand U15126 (N_15126,N_14609,N_12163);
nor U15127 (N_15127,N_13769,N_14300);
xnor U15128 (N_15128,N_12621,N_13934);
and U15129 (N_15129,N_12244,N_13597);
nor U15130 (N_15130,N_13751,N_13569);
nor U15131 (N_15131,N_14952,N_13810);
or U15132 (N_15132,N_13981,N_12350);
nand U15133 (N_15133,N_13268,N_13571);
or U15134 (N_15134,N_14026,N_13442);
or U15135 (N_15135,N_14049,N_13506);
nand U15136 (N_15136,N_13925,N_13216);
and U15137 (N_15137,N_14440,N_13459);
or U15138 (N_15138,N_14765,N_12611);
or U15139 (N_15139,N_14181,N_12481);
xnor U15140 (N_15140,N_14108,N_14953);
or U15141 (N_15141,N_13651,N_14880);
nor U15142 (N_15142,N_12630,N_12752);
nor U15143 (N_15143,N_13371,N_13116);
and U15144 (N_15144,N_13431,N_14286);
nor U15145 (N_15145,N_12362,N_13627);
and U15146 (N_15146,N_13389,N_14819);
nor U15147 (N_15147,N_12990,N_14718);
and U15148 (N_15148,N_12631,N_13343);
and U15149 (N_15149,N_13278,N_13658);
or U15150 (N_15150,N_14244,N_13118);
nor U15151 (N_15151,N_12440,N_14735);
or U15152 (N_15152,N_12180,N_12271);
nor U15153 (N_15153,N_14520,N_14033);
or U15154 (N_15154,N_12607,N_12658);
and U15155 (N_15155,N_13595,N_14073);
nor U15156 (N_15156,N_13990,N_13036);
and U15157 (N_15157,N_12051,N_12997);
xor U15158 (N_15158,N_12124,N_14238);
and U15159 (N_15159,N_14381,N_13186);
or U15160 (N_15160,N_12647,N_14334);
nand U15161 (N_15161,N_13030,N_12403);
nand U15162 (N_15162,N_12073,N_14738);
nor U15163 (N_15163,N_14914,N_14290);
or U15164 (N_15164,N_14470,N_13162);
nand U15165 (N_15165,N_14274,N_14296);
or U15166 (N_15166,N_12936,N_12918);
or U15167 (N_15167,N_14173,N_13410);
and U15168 (N_15168,N_12881,N_14742);
and U15169 (N_15169,N_13206,N_13358);
or U15170 (N_15170,N_14029,N_13122);
xnor U15171 (N_15171,N_14509,N_14143);
nand U15172 (N_15172,N_14570,N_13626);
nor U15173 (N_15173,N_14176,N_14245);
nand U15174 (N_15174,N_14679,N_13606);
nor U15175 (N_15175,N_12002,N_12976);
or U15176 (N_15176,N_14863,N_12220);
nand U15177 (N_15177,N_12108,N_13722);
or U15178 (N_15178,N_13137,N_14088);
nor U15179 (N_15179,N_12177,N_13912);
nand U15180 (N_15180,N_13585,N_14298);
nor U15181 (N_15181,N_14002,N_12770);
nor U15182 (N_15182,N_12040,N_13976);
nand U15183 (N_15183,N_12081,N_14899);
and U15184 (N_15184,N_13941,N_14039);
or U15185 (N_15185,N_12578,N_12473);
nand U15186 (N_15186,N_14662,N_12184);
xnor U15187 (N_15187,N_12531,N_13142);
xor U15188 (N_15188,N_13329,N_14389);
nor U15189 (N_15189,N_13641,N_12889);
nor U15190 (N_15190,N_14729,N_14347);
xor U15191 (N_15191,N_12353,N_14089);
nand U15192 (N_15192,N_14712,N_12921);
and U15193 (N_15193,N_13377,N_12169);
xor U15194 (N_15194,N_13402,N_13586);
xnor U15195 (N_15195,N_13640,N_14622);
xnor U15196 (N_15196,N_13180,N_12680);
and U15197 (N_15197,N_13603,N_12919);
or U15198 (N_15198,N_14183,N_14524);
nand U15199 (N_15199,N_12986,N_13156);
and U15200 (N_15200,N_13812,N_12788);
and U15201 (N_15201,N_12870,N_13795);
and U15202 (N_15202,N_12375,N_13399);
nor U15203 (N_15203,N_13512,N_13670);
xnor U15204 (N_15204,N_12486,N_14835);
and U15205 (N_15205,N_12093,N_12673);
xnor U15206 (N_15206,N_12910,N_13775);
and U15207 (N_15207,N_13850,N_12273);
and U15208 (N_15208,N_13684,N_13027);
nor U15209 (N_15209,N_12074,N_12939);
or U15210 (N_15210,N_12192,N_13819);
nand U15211 (N_15211,N_13873,N_12609);
and U15212 (N_15212,N_12933,N_13830);
xor U15213 (N_15213,N_14393,N_12954);
nor U15214 (N_15214,N_12674,N_14000);
xor U15215 (N_15215,N_13577,N_12765);
or U15216 (N_15216,N_12984,N_12070);
and U15217 (N_15217,N_13088,N_14232);
nor U15218 (N_15218,N_14991,N_13533);
nand U15219 (N_15219,N_12693,N_12551);
and U15220 (N_15220,N_14104,N_12964);
and U15221 (N_15221,N_12477,N_12659);
or U15222 (N_15222,N_14980,N_13681);
xnor U15223 (N_15223,N_13561,N_13073);
xnor U15224 (N_15224,N_14151,N_14567);
nor U15225 (N_15225,N_14569,N_14338);
and U15226 (N_15226,N_14438,N_14113);
xnor U15227 (N_15227,N_13672,N_12277);
and U15228 (N_15228,N_13896,N_13235);
nand U15229 (N_15229,N_12063,N_13120);
or U15230 (N_15230,N_13261,N_12737);
xor U15231 (N_15231,N_13632,N_12838);
nor U15232 (N_15232,N_14361,N_13428);
xnor U15233 (N_15233,N_14324,N_13477);
xnor U15234 (N_15234,N_13430,N_13064);
nand U15235 (N_15235,N_13948,N_14947);
nor U15236 (N_15236,N_14858,N_13885);
xor U15237 (N_15237,N_14777,N_14235);
xnor U15238 (N_15238,N_13950,N_13813);
xnor U15239 (N_15239,N_13565,N_13267);
or U15240 (N_15240,N_12597,N_13305);
and U15241 (N_15241,N_12072,N_14429);
xor U15242 (N_15242,N_12274,N_14106);
or U15243 (N_15243,N_12055,N_12956);
and U15244 (N_15244,N_14062,N_12335);
xor U15245 (N_15245,N_14022,N_12196);
nand U15246 (N_15246,N_13817,N_12129);
nor U15247 (N_15247,N_14353,N_12830);
nand U15248 (N_15248,N_13035,N_13805);
nor U15249 (N_15249,N_14994,N_14150);
nor U15250 (N_15250,N_12060,N_12468);
and U15251 (N_15251,N_14476,N_14156);
nor U15252 (N_15252,N_12882,N_14596);
or U15253 (N_15253,N_13820,N_13311);
nor U15254 (N_15254,N_12556,N_13336);
nand U15255 (N_15255,N_13094,N_14697);
nor U15256 (N_15256,N_12402,N_13136);
nor U15257 (N_15257,N_14511,N_14216);
and U15258 (N_15258,N_14517,N_12016);
xor U15259 (N_15259,N_12312,N_13520);
nand U15260 (N_15260,N_13676,N_12255);
xor U15261 (N_15261,N_13698,N_13409);
or U15262 (N_15262,N_14387,N_13274);
nand U15263 (N_15263,N_13272,N_12897);
nor U15264 (N_15264,N_14714,N_14936);
nand U15265 (N_15265,N_14482,N_12521);
or U15266 (N_15266,N_13152,N_12011);
xor U15267 (N_15267,N_13308,N_12644);
or U15268 (N_15268,N_13484,N_14877);
and U15269 (N_15269,N_12115,N_14024);
xor U15270 (N_15270,N_12497,N_12024);
nor U15271 (N_15271,N_13300,N_12851);
nand U15272 (N_15272,N_14593,N_13870);
and U15273 (N_15273,N_14924,N_12949);
or U15274 (N_15274,N_14252,N_13161);
and U15275 (N_15275,N_13974,N_14013);
and U15276 (N_15276,N_14316,N_14890);
nand U15277 (N_15277,N_13938,N_13620);
or U15278 (N_15278,N_13424,N_13840);
nor U15279 (N_15279,N_13101,N_12263);
nand U15280 (N_15280,N_12793,N_14842);
or U15281 (N_15281,N_12666,N_13087);
nand U15282 (N_15282,N_12583,N_14161);
nand U15283 (N_15283,N_14799,N_14654);
nand U15284 (N_15284,N_14745,N_14845);
xnor U15285 (N_15285,N_14873,N_12527);
nand U15286 (N_15286,N_13618,N_13968);
and U15287 (N_15287,N_13650,N_12065);
nor U15288 (N_15288,N_13104,N_14955);
xor U15289 (N_15289,N_12317,N_12699);
nor U15290 (N_15290,N_13514,N_12703);
nand U15291 (N_15291,N_14370,N_14795);
and U15292 (N_15292,N_14457,N_14726);
nand U15293 (N_15293,N_14722,N_13877);
or U15294 (N_15294,N_13729,N_14639);
and U15295 (N_15295,N_14778,N_14120);
nor U15296 (N_15296,N_14249,N_13794);
and U15297 (N_15297,N_13452,N_14606);
nor U15298 (N_15298,N_14036,N_13674);
nor U15299 (N_15299,N_13979,N_13806);
and U15300 (N_15300,N_14598,N_13382);
nor U15301 (N_15301,N_12270,N_12759);
nand U15302 (N_15302,N_12173,N_14284);
nand U15303 (N_15303,N_13465,N_12064);
or U15304 (N_15304,N_14492,N_14496);
or U15305 (N_15305,N_13176,N_13292);
or U15306 (N_15306,N_12057,N_13356);
nor U15307 (N_15307,N_14223,N_14028);
nand U15308 (N_15308,N_12107,N_12416);
xnor U15309 (N_15309,N_14921,N_12726);
xnor U15310 (N_15310,N_14988,N_12147);
nor U15311 (N_15311,N_13772,N_14906);
nor U15312 (N_15312,N_12648,N_14435);
and U15313 (N_15313,N_12702,N_14671);
xnor U15314 (N_15314,N_13083,N_13978);
nand U15315 (N_15315,N_12885,N_13170);
or U15316 (N_15316,N_13463,N_13709);
xnor U15317 (N_15317,N_13029,N_12853);
xor U15318 (N_15318,N_13482,N_12591);
nand U15319 (N_15319,N_14413,N_13636);
and U15320 (N_15320,N_13786,N_12331);
xnor U15321 (N_15321,N_12245,N_14097);
nor U15322 (N_15322,N_14696,N_13624);
nand U15323 (N_15323,N_12633,N_13852);
and U15324 (N_15324,N_13528,N_12710);
or U15325 (N_15325,N_14529,N_14403);
xnor U15326 (N_15326,N_13588,N_14264);
xor U15327 (N_15327,N_12021,N_14938);
nand U15328 (N_15328,N_12675,N_12837);
xor U15329 (N_15329,N_14532,N_12079);
nand U15330 (N_15330,N_12865,N_12360);
nor U15331 (N_15331,N_14060,N_12635);
nor U15332 (N_15332,N_14016,N_12983);
and U15333 (N_15333,N_12246,N_12846);
nand U15334 (N_15334,N_12747,N_13582);
or U15335 (N_15335,N_13711,N_14340);
xnor U15336 (N_15336,N_13917,N_12456);
nor U15337 (N_15337,N_12683,N_13758);
nor U15338 (N_15338,N_14963,N_12758);
or U15339 (N_15339,N_14871,N_14809);
nand U15340 (N_15340,N_13957,N_14390);
nor U15341 (N_15341,N_13450,N_13103);
xnor U15342 (N_15342,N_13370,N_12972);
nor U15343 (N_15343,N_13129,N_14887);
and U15344 (N_15344,N_12149,N_12823);
nor U15345 (N_15345,N_13200,N_12046);
and U15346 (N_15346,N_14449,N_14926);
or U15347 (N_15347,N_14273,N_13220);
or U15348 (N_15348,N_14304,N_13952);
nand U15349 (N_15349,N_13079,N_13572);
and U15350 (N_15350,N_12112,N_14085);
nand U15351 (N_15351,N_14056,N_13487);
nor U15352 (N_15352,N_12709,N_12701);
or U15353 (N_15353,N_13973,N_13591);
nand U15354 (N_15354,N_13147,N_14522);
and U15355 (N_15355,N_13907,N_13231);
nand U15356 (N_15356,N_14581,N_12886);
xnor U15357 (N_15357,N_12602,N_13853);
nand U15358 (N_15358,N_14260,N_14655);
xnor U15359 (N_15359,N_12304,N_14278);
nor U15360 (N_15360,N_13357,N_14701);
xor U15361 (N_15361,N_14650,N_14732);
nand U15362 (N_15362,N_14703,N_14757);
nand U15363 (N_15363,N_14432,N_14530);
nand U15364 (N_15364,N_13921,N_13634);
nand U15365 (N_15365,N_12447,N_14736);
and U15366 (N_15366,N_13633,N_12306);
nand U15367 (N_15367,N_14660,N_13997);
xor U15368 (N_15368,N_13552,N_13960);
nand U15369 (N_15369,N_14220,N_12457);
or U15370 (N_15370,N_12878,N_14762);
xnor U15371 (N_15371,N_13415,N_13432);
xor U15372 (N_15372,N_13710,N_12893);
nor U15373 (N_15373,N_12415,N_12628);
and U15374 (N_15374,N_14538,N_14774);
and U15375 (N_15375,N_13243,N_13622);
nor U15376 (N_15376,N_14325,N_13920);
or U15377 (N_15377,N_13730,N_14839);
or U15378 (N_15378,N_12210,N_12825);
xor U15379 (N_15379,N_12742,N_13532);
and U15380 (N_15380,N_14534,N_14146);
and U15381 (N_15381,N_13685,N_12776);
nor U15382 (N_15382,N_13271,N_12957);
xor U15383 (N_15383,N_14331,N_13888);
and U15384 (N_15384,N_14155,N_12143);
nor U15385 (N_15385,N_12959,N_14702);
and U15386 (N_15386,N_13384,N_12008);
xor U15387 (N_15387,N_13746,N_14825);
and U15388 (N_15388,N_13809,N_12238);
and U15389 (N_15389,N_14357,N_14805);
xor U15390 (N_15390,N_13368,N_13866);
nor U15391 (N_15391,N_13657,N_14625);
or U15392 (N_15392,N_14129,N_13720);
nor U15393 (N_15393,N_14759,N_14860);
nor U15394 (N_15394,N_14897,N_13944);
nand U15395 (N_15395,N_14711,N_13664);
and U15396 (N_15396,N_14190,N_14303);
and U15397 (N_15397,N_13998,N_14785);
or U15398 (N_15398,N_14321,N_12998);
xnor U15399 (N_15399,N_12339,N_14184);
xnor U15400 (N_15400,N_13906,N_12560);
nand U15401 (N_15401,N_12844,N_12723);
nand U15402 (N_15402,N_14967,N_12038);
nor U15403 (N_15403,N_14595,N_12087);
nor U15404 (N_15404,N_14527,N_13139);
xor U15405 (N_15405,N_13985,N_13196);
nand U15406 (N_15406,N_13937,N_12023);
nor U15407 (N_15407,N_12866,N_13980);
or U15408 (N_15408,N_12128,N_14329);
nor U15409 (N_15409,N_12315,N_13679);
xor U15410 (N_15410,N_14344,N_12506);
or U15411 (N_15411,N_12600,N_13691);
or U15412 (N_15412,N_14755,N_13352);
and U15413 (N_15413,N_14913,N_12961);
or U15414 (N_15414,N_12754,N_13212);
xor U15415 (N_15415,N_14204,N_14256);
or U15416 (N_15416,N_12197,N_13647);
nand U15417 (N_15417,N_12369,N_13443);
xnor U15418 (N_15418,N_14592,N_12017);
xor U15419 (N_15419,N_14261,N_13293);
nand U15420 (N_15420,N_13780,N_14317);
or U15421 (N_15421,N_12321,N_12704);
xnor U15422 (N_15422,N_13026,N_13822);
or U15423 (N_15423,N_13610,N_13965);
and U15424 (N_15424,N_13337,N_12899);
and U15425 (N_15425,N_12058,N_14351);
nor U15426 (N_15426,N_13219,N_14589);
or U15427 (N_15427,N_13910,N_12706);
xnor U15428 (N_15428,N_12785,N_12620);
and U15429 (N_15429,N_12424,N_13249);
nor U15430 (N_15430,N_14998,N_12279);
nor U15431 (N_15431,N_14445,N_12039);
or U15432 (N_15432,N_12109,N_13330);
nor U15433 (N_15433,N_13639,N_14467);
nand U15434 (N_15434,N_14208,N_13547);
nor U15435 (N_15435,N_12662,N_13057);
nor U15436 (N_15436,N_14657,N_13168);
nor U15437 (N_15437,N_13022,N_12618);
or U15438 (N_15438,N_14977,N_14250);
and U15439 (N_15439,N_14776,N_13943);
nand U15440 (N_15440,N_13656,N_14192);
xnor U15441 (N_15441,N_14731,N_14493);
and U15442 (N_15442,N_12158,N_14590);
or U15443 (N_15443,N_14756,N_13913);
and U15444 (N_15444,N_13833,N_14446);
nor U15445 (N_15445,N_12242,N_12059);
nand U15446 (N_15446,N_13111,N_12879);
nand U15447 (N_15447,N_14643,N_14480);
or U15448 (N_15448,N_14545,N_13114);
nor U15449 (N_15449,N_12533,N_12094);
xnor U15450 (N_15450,N_14694,N_13863);
xor U15451 (N_15451,N_14506,N_13551);
nor U15452 (N_15452,N_14222,N_13113);
nor U15453 (N_15453,N_13353,N_12679);
xor U15454 (N_15454,N_12117,N_12567);
and U15455 (N_15455,N_13559,N_13825);
and U15456 (N_15456,N_13225,N_12202);
nor U15457 (N_15457,N_14894,N_14337);
nor U15458 (N_15458,N_14961,N_13218);
or U15459 (N_15459,N_12420,N_13049);
nor U15460 (N_15460,N_13942,N_14883);
or U15461 (N_15461,N_14874,N_12982);
or U15462 (N_15462,N_14787,N_14747);
nand U15463 (N_15463,N_14554,N_12344);
xor U15464 (N_15464,N_12536,N_14063);
xnor U15465 (N_15465,N_12296,N_12206);
xor U15466 (N_15466,N_12750,N_13233);
and U15467 (N_15467,N_12963,N_12684);
nand U15468 (N_15468,N_12111,N_14583);
or U15469 (N_15469,N_14203,N_13517);
nand U15470 (N_15470,N_12558,N_13768);
or U15471 (N_15471,N_12407,N_13020);
xor U15472 (N_15472,N_14380,N_12048);
and U15473 (N_15473,N_14468,N_13964);
or U15474 (N_15474,N_12448,N_14107);
nand U15475 (N_15475,N_13902,N_12026);
and U15476 (N_15476,N_12346,N_12653);
and U15477 (N_15477,N_13909,N_13464);
xor U15478 (N_15478,N_12970,N_13718);
or U15479 (N_15479,N_13504,N_13495);
or U15480 (N_15480,N_14096,N_13181);
nor U15481 (N_15481,N_12412,N_13017);
nand U15482 (N_15482,N_14312,N_14995);
or U15483 (N_15483,N_12012,N_14591);
nor U15484 (N_15484,N_12366,N_13865);
nor U15485 (N_15485,N_12900,N_13770);
nand U15486 (N_15486,N_14868,N_12461);
nand U15487 (N_15487,N_14793,N_13398);
or U15488 (N_15488,N_12736,N_12225);
xnor U15489 (N_15489,N_13843,N_14363);
nor U15490 (N_15490,N_13468,N_12718);
xor U15491 (N_15491,N_14420,N_12032);
nand U15492 (N_15492,N_13229,N_12045);
or U15493 (N_15493,N_14214,N_14297);
or U15494 (N_15494,N_12397,N_14629);
or U15495 (N_15495,N_13787,N_13767);
nor U15496 (N_15496,N_12790,N_14744);
and U15497 (N_15497,N_14437,N_14659);
and U15498 (N_15498,N_14915,N_14647);
nand U15499 (N_15499,N_13546,N_12562);
xnor U15500 (N_15500,N_13972,N_13275);
nand U15501 (N_15501,N_13123,N_12843);
or U15502 (N_15502,N_14678,N_13953);
or U15503 (N_15503,N_12715,N_13749);
xnor U15504 (N_15504,N_14349,N_12388);
xnor U15505 (N_15505,N_12382,N_14571);
nor U15506 (N_15506,N_13187,N_12425);
and U15507 (N_15507,N_14441,N_12623);
and U15508 (N_15508,N_14067,N_14739);
or U15509 (N_15509,N_12189,N_13623);
nor U15510 (N_15510,N_14378,N_14651);
and U15511 (N_15511,N_14326,N_12934);
nor U15512 (N_15512,N_14069,N_14102);
nand U15513 (N_15513,N_14541,N_14838);
xnor U15514 (N_15514,N_14463,N_13935);
xnor U15515 (N_15515,N_13701,N_12349);
and U15516 (N_15516,N_12347,N_14352);
nor U15517 (N_15517,N_12050,N_12917);
xnor U15518 (N_15518,N_14763,N_13967);
and U15519 (N_15519,N_13778,N_12080);
or U15520 (N_15520,N_13625,N_13013);
nand U15521 (N_15521,N_14048,N_12389);
xnor U15522 (N_15522,N_13677,N_14875);
nand U15523 (N_15523,N_13310,N_12832);
and U15524 (N_15524,N_13062,N_12555);
nand U15525 (N_15525,N_12951,N_12019);
nor U15526 (N_15526,N_12614,N_12223);
or U15527 (N_15527,N_13899,N_12932);
and U15528 (N_15528,N_12187,N_12857);
nor U15529 (N_15529,N_12795,N_13446);
nor U15530 (N_15530,N_13494,N_12833);
nand U15531 (N_15531,N_13322,N_12122);
and U15532 (N_15532,N_14198,N_12401);
and U15533 (N_15533,N_13712,N_14027);
and U15534 (N_15534,N_14394,N_14453);
nand U15535 (N_15535,N_12626,N_12110);
xnor U15536 (N_15536,N_13349,N_14962);
and U15537 (N_15537,N_13879,N_14719);
nand U15538 (N_15538,N_12656,N_13303);
nor U15539 (N_15539,N_13177,N_14255);
and U15540 (N_15540,N_12546,N_14663);
or U15541 (N_15541,N_14137,N_14383);
xor U15542 (N_15542,N_12309,N_14856);
xor U15543 (N_15543,N_14631,N_13541);
nor U15544 (N_15544,N_12148,N_12325);
nand U15545 (N_15545,N_13166,N_13130);
xor U15546 (N_15546,N_13615,N_12582);
nand U15547 (N_15547,N_13066,N_13280);
xnor U15548 (N_15548,N_12826,N_12232);
or U15549 (N_15549,N_12342,N_13476);
and U15550 (N_15550,N_12234,N_14397);
xor U15551 (N_15551,N_12156,N_13522);
nand U15552 (N_15552,N_14052,N_12989);
nor U15553 (N_15553,N_13717,N_14644);
and U15554 (N_15554,N_13708,N_14117);
and U15555 (N_15555,N_13727,N_14535);
and U15556 (N_15556,N_14916,N_13251);
and U15557 (N_15557,N_12285,N_13385);
nand U15558 (N_15558,N_13056,N_12384);
xor U15559 (N_15559,N_12505,N_14125);
nand U15560 (N_15560,N_14710,N_13360);
and U15561 (N_15561,N_12280,N_14771);
nand U15562 (N_15562,N_12503,N_13080);
xor U15563 (N_15563,N_13673,N_12379);
nor U15564 (N_15564,N_14269,N_12446);
nor U15565 (N_15565,N_14101,N_12975);
xor U15566 (N_15566,N_14725,N_12181);
and U15567 (N_15567,N_14677,N_12671);
xnor U15568 (N_15568,N_12942,N_14045);
and U15569 (N_15569,N_14475,N_12444);
nand U15570 (N_15570,N_12272,N_12787);
and U15571 (N_15571,N_14642,N_14905);
nor U15572 (N_15572,N_13513,N_13175);
or U15573 (N_15573,N_12867,N_14428);
nand U15574 (N_15574,N_12717,N_12561);
xnor U15575 (N_15575,N_12792,N_13545);
and U15576 (N_15576,N_12138,N_13962);
xnor U15577 (N_15577,N_14674,N_14605);
nand U15578 (N_15578,N_13821,N_14105);
nor U15579 (N_15579,N_12807,N_13199);
xor U15580 (N_15580,N_13488,N_13728);
nor U15581 (N_15581,N_14949,N_14292);
and U15582 (N_15582,N_13050,N_13440);
xor U15583 (N_15583,N_13761,N_13126);
or U15584 (N_15584,N_14908,N_12332);
nand U15585 (N_15585,N_13047,N_13246);
and U15586 (N_15586,N_14603,N_12137);
xnor U15587 (N_15587,N_12153,N_14266);
or U15588 (N_15588,N_14018,N_14008);
and U15589 (N_15589,N_12423,N_12449);
or U15590 (N_15590,N_12014,N_13726);
nand U15591 (N_15591,N_13100,N_14189);
nor U15592 (N_15592,N_12528,N_13956);
or U15593 (N_15593,N_14810,N_13946);
nor U15594 (N_15594,N_13621,N_14130);
or U15595 (N_15595,N_13503,N_12883);
nand U15596 (N_15596,N_12977,N_13230);
or U15597 (N_15597,N_13285,N_12895);
and U15598 (N_15598,N_13406,N_13995);
nand U15599 (N_15599,N_12761,N_12818);
nor U15600 (N_15600,N_12469,N_14229);
or U15601 (N_15601,N_13660,N_13945);
nor U15602 (N_15602,N_13151,N_13745);
or U15603 (N_15603,N_12524,N_14037);
or U15604 (N_15604,N_13076,N_13887);
nand U15605 (N_15605,N_14237,N_13433);
or U15606 (N_15606,N_14345,N_12231);
xor U15607 (N_15607,N_12490,N_13250);
nor U15608 (N_15608,N_12436,N_12636);
and U15609 (N_15609,N_13171,N_13923);
nor U15610 (N_15610,N_12185,N_12925);
nor U15611 (N_15611,N_12371,N_13856);
xor U15612 (N_15612,N_14020,N_12733);
nand U15613 (N_15613,N_13454,N_14865);
nand U15614 (N_15614,N_12098,N_12037);
nand U15615 (N_15615,N_14400,N_13334);
nor U15616 (N_15616,N_13760,N_12711);
nor U15617 (N_15617,N_12027,N_13339);
or U15618 (N_15618,N_12452,N_14459);
xnor U15619 (N_15619,N_12845,N_14139);
and U15620 (N_15620,N_13619,N_13851);
nand U15621 (N_15621,N_12266,N_12141);
and U15622 (N_15622,N_13763,N_13302);
or U15623 (N_15623,N_12372,N_14375);
or U15624 (N_15624,N_14030,N_13816);
and U15625 (N_15625,N_13347,N_12322);
nor U15626 (N_15626,N_14162,N_12357);
and U15627 (N_15627,N_14930,N_13999);
nand U15628 (N_15628,N_14599,N_12649);
xnor U15629 (N_15629,N_12967,N_13736);
nand U15630 (N_15630,N_14202,N_13081);
and U15631 (N_15631,N_12025,N_12290);
and U15632 (N_15632,N_12617,N_14144);
and U15633 (N_15633,N_13413,N_14531);
xnor U15634 (N_15634,N_13849,N_13881);
xnor U15635 (N_15635,N_13098,N_12519);
or U15636 (N_15636,N_12378,N_13791);
or U15637 (N_15637,N_12356,N_14231);
xnor U15638 (N_15638,N_12213,N_14804);
nor U15639 (N_15639,N_12962,N_13498);
nor U15640 (N_15640,N_12175,N_12467);
nand U15641 (N_15641,N_12494,N_12955);
nand U15642 (N_15642,N_12029,N_12168);
and U15643 (N_15643,N_12809,N_12247);
xor U15644 (N_15644,N_13564,N_13529);
nor U15645 (N_15645,N_13580,N_12020);
xor U15646 (N_15646,N_13033,N_12454);
xor U15647 (N_15647,N_14167,N_12619);
xor U15648 (N_15648,N_14773,N_14857);
nor U15649 (N_15649,N_14861,N_14011);
nor U15650 (N_15650,N_13631,N_14852);
nand U15651 (N_15651,N_12249,N_14705);
nor U15652 (N_15652,N_14687,N_13189);
or U15653 (N_15653,N_12840,N_13046);
or U15654 (N_15654,N_13007,N_12393);
and U15655 (N_15655,N_12849,N_14623);
nand U15656 (N_15656,N_14123,N_14133);
nand U15657 (N_15657,N_13241,N_12517);
or U15658 (N_15658,N_12613,N_14092);
nor U15659 (N_15659,N_14925,N_14550);
xor U15660 (N_15660,N_13348,N_14709);
nor U15661 (N_15661,N_14055,N_12257);
nand U15662 (N_15662,N_13762,N_12140);
and U15663 (N_15663,N_12431,N_14093);
or U15664 (N_15664,N_13756,N_13688);
nor U15665 (N_15665,N_13500,N_12580);
nand U15666 (N_15666,N_13690,N_12096);
nand U15667 (N_15667,N_14772,N_13240);
nor U15668 (N_15668,N_14689,N_12753);
nor U15669 (N_15669,N_12928,N_14646);
nand U15670 (N_15670,N_14415,N_13781);
nor U15671 (N_15671,N_12937,N_14434);
nor U15672 (N_15672,N_13724,N_12267);
xor U15673 (N_15673,N_12599,N_12047);
and U15674 (N_15674,N_12590,N_12755);
or U15675 (N_15675,N_14059,N_14816);
and U15676 (N_15676,N_14280,N_14004);
or U15677 (N_15677,N_13237,N_12608);
or U15678 (N_15678,N_12732,N_12848);
xor U15679 (N_15679,N_14608,N_12493);
or U15680 (N_15680,N_12722,N_14734);
nand U15681 (N_15681,N_13544,N_12399);
nand U15682 (N_15682,N_14942,N_13872);
nand U15683 (N_15683,N_14536,N_14233);
or U15684 (N_15684,N_12953,N_13771);
or U15685 (N_15685,N_12345,N_12872);
and U15686 (N_15686,N_14323,N_12686);
or U15687 (N_15687,N_12884,N_14427);
xnor U15688 (N_15688,N_13198,N_14354);
and U15689 (N_15689,N_14043,N_12086);
nor U15690 (N_15690,N_12010,N_13593);
xnor U15691 (N_15691,N_12841,N_13157);
or U15692 (N_15692,N_12654,N_13307);
or U15693 (N_15693,N_13321,N_12078);
xor U15694 (N_15694,N_14614,N_14185);
or U15695 (N_15695,N_13519,N_12091);
or U15696 (N_15696,N_12999,N_14277);
nor U15697 (N_15697,N_13436,N_14811);
and U15698 (N_15698,N_14373,N_12367);
nand U15699 (N_15699,N_14813,N_14888);
xnor U15700 (N_15700,N_12483,N_12515);
and U15701 (N_15701,N_13739,N_13190);
or U15702 (N_15702,N_14841,N_13279);
and U15703 (N_15703,N_14328,N_13605);
nor U15704 (N_15704,N_14275,N_14489);
nand U15705 (N_15705,N_13531,N_14965);
nor U15706 (N_15706,N_12150,N_12941);
and U15707 (N_15707,N_12781,N_13014);
nor U15708 (N_15708,N_12394,N_12672);
nor U15709 (N_15709,N_12905,N_13437);
or U15710 (N_15710,N_14487,N_13562);
nor U15711 (N_15711,N_14945,N_13635);
xor U15712 (N_15712,N_14417,N_12772);
and U15713 (N_15713,N_12566,N_12170);
nor U15714 (N_15714,N_13173,N_12198);
xnor U15715 (N_15715,N_13648,N_14308);
xor U15716 (N_15716,N_13481,N_14989);
and U15717 (N_15717,N_12464,N_12655);
xnor U15718 (N_15718,N_12358,N_13324);
nor U15719 (N_15719,N_12525,N_14341);
xor U15720 (N_15720,N_14460,N_12154);
xnor U15721 (N_15721,N_14882,N_13653);
nand U15722 (N_15722,N_13209,N_12973);
nand U15723 (N_15723,N_13208,N_14750);
and U15724 (N_15724,N_12968,N_14411);
or U15725 (N_15725,N_13072,N_12887);
or U15726 (N_15726,N_12036,N_12355);
xor U15727 (N_15727,N_14201,N_12831);
xnor U15728 (N_15728,N_13179,N_13010);
nor U15729 (N_15729,N_13163,N_13993);
or U15730 (N_15730,N_14314,N_14330);
xnor U15731 (N_15731,N_13599,N_14006);
and U15732 (N_15732,N_13908,N_13869);
and U15733 (N_15733,N_14371,N_14454);
nor U15734 (N_15734,N_13195,N_13827);
nand U15735 (N_15735,N_12235,N_12404);
and U15736 (N_15736,N_14164,N_12912);
and U15737 (N_15737,N_14376,N_12496);
nor U15738 (N_15738,N_13444,N_13290);
or U15739 (N_15739,N_14230,N_13417);
nor U15740 (N_15740,N_13106,N_12365);
xor U15741 (N_15741,N_12119,N_12708);
nor U15742 (N_15742,N_14904,N_13721);
or U15743 (N_15743,N_12437,N_13333);
nand U15744 (N_15744,N_12100,N_13735);
nand U15745 (N_15745,N_14412,N_12164);
xor U15746 (N_15746,N_12634,N_14760);
xnor U15747 (N_15747,N_13502,N_12559);
and U15748 (N_15748,N_14017,N_12042);
nor U15749 (N_15749,N_14740,N_12924);
and U15750 (N_15750,N_13703,N_12791);
xor U15751 (N_15751,N_14367,N_14767);
and U15752 (N_15752,N_14940,N_14851);
and U15753 (N_15753,N_12302,N_14090);
and U15754 (N_15754,N_13458,N_13700);
or U15755 (N_15755,N_12200,N_13511);
nand U15756 (N_15756,N_14637,N_12387);
or U15757 (N_15757,N_14318,N_12373);
xnor U15758 (N_15758,N_12439,N_13882);
nor U15759 (N_15759,N_12022,N_14276);
nand U15760 (N_15760,N_14514,N_14163);
nand U15761 (N_15761,N_14169,N_13085);
nand U15762 (N_15762,N_12514,N_14472);
and U15763 (N_15763,N_13602,N_12904);
or U15764 (N_15764,N_13411,N_13099);
nand U15765 (N_15765,N_14692,N_14366);
nor U15766 (N_15766,N_13491,N_12987);
nor U15767 (N_15767,N_13835,N_14270);
xnor U15768 (N_15768,N_12261,N_13439);
nor U15769 (N_15769,N_12827,N_14188);
nand U15770 (N_15770,N_14766,N_13989);
and U15771 (N_15771,N_12125,N_12668);
and U15772 (N_15772,N_13844,N_13188);
xor U15773 (N_15773,N_13089,N_14684);
or U15774 (N_15774,N_12275,N_13742);
nand U15775 (N_15775,N_14934,N_14047);
xor U15776 (N_15776,N_14688,N_12061);
nand U15777 (N_15777,N_13608,N_14082);
xor U15778 (N_15778,N_12692,N_14486);
and U15779 (N_15779,N_12299,N_13270);
nand U15780 (N_15780,N_13153,N_13675);
or U15781 (N_15781,N_12670,N_14253);
xor U15782 (N_15782,N_12540,N_13455);
and U15783 (N_15783,N_14794,N_13327);
nor U15784 (N_15784,N_13226,N_14450);
nand U15785 (N_15785,N_14197,N_12174);
or U15786 (N_15786,N_14853,N_13876);
and U15787 (N_15787,N_13419,N_14552);
or U15788 (N_15788,N_14730,N_14698);
and U15789 (N_15789,N_14134,N_14768);
nand U15790 (N_15790,N_13003,N_12229);
xor U15791 (N_15791,N_12926,N_13987);
or U15792 (N_15792,N_14796,N_14119);
or U15793 (N_15793,N_14516,N_13596);
nand U15794 (N_15794,N_13792,N_13016);
or U15795 (N_15795,N_14481,N_13414);
nand U15796 (N_15796,N_13460,N_12898);
and U15797 (N_15797,N_12646,N_13515);
nor U15798 (N_15798,N_13699,N_14160);
or U15799 (N_15799,N_14444,N_12000);
or U15800 (N_15800,N_13154,N_13469);
nand U15801 (N_15801,N_13145,N_12056);
and U15802 (N_15802,N_14565,N_12165);
nand U15803 (N_15803,N_12862,N_14513);
and U15804 (N_15804,N_14038,N_14640);
and U15805 (N_15805,N_14782,N_13550);
or U15806 (N_15806,N_13655,N_12947);
xnor U15807 (N_15807,N_14850,N_13861);
nor U15808 (N_15808,N_14652,N_12297);
nand U15809 (N_15809,N_12584,N_12043);
xor U15810 (N_15810,N_12764,N_14604);
nor U15811 (N_15811,N_14140,N_12237);
and U15812 (N_15812,N_13932,N_13814);
or U15813 (N_15813,N_13018,N_12762);
xor U15814 (N_15814,N_13929,N_14551);
or U15815 (N_15815,N_14932,N_12092);
nand U15816 (N_15816,N_13916,N_14500);
nor U15817 (N_15817,N_13174,N_12908);
or U15818 (N_15818,N_12734,N_13367);
or U15819 (N_15819,N_13178,N_12698);
and U15820 (N_15820,N_13977,N_12538);
xnor U15821 (N_15821,N_13065,N_14884);
nor U15822 (N_15822,N_13802,N_12920);
or U15823 (N_15823,N_12577,N_14957);
nor U15824 (N_15824,N_12539,N_14675);
or U15825 (N_15825,N_12363,N_14479);
or U15826 (N_15826,N_13966,N_12660);
or U15827 (N_15827,N_14537,N_12629);
or U15828 (N_15828,N_12922,N_12712);
and U15829 (N_15829,N_14885,N_12132);
nand U15830 (N_15830,N_14896,N_13539);
or U15831 (N_15831,N_12901,N_14374);
nor U15832 (N_15832,N_13252,N_14748);
nor U15833 (N_15833,N_14784,N_13320);
xnor U15834 (N_15834,N_12508,N_12534);
or U15835 (N_15835,N_14272,N_12193);
nor U15836 (N_15836,N_13453,N_13093);
xor U15837 (N_15837,N_13601,N_14299);
nand U15838 (N_15838,N_13568,N_12233);
xor U15839 (N_15839,N_12511,N_14968);
and U15840 (N_15840,N_12814,N_14587);
and U15841 (N_15841,N_12421,N_14282);
xor U15842 (N_15842,N_14174,N_13257);
or U15843 (N_15843,N_14823,N_12856);
nand U15844 (N_15844,N_13750,N_12293);
and U15845 (N_15845,N_14539,N_13354);
or U15846 (N_15846,N_14939,N_13678);
nand U15847 (N_15847,N_13386,N_12643);
and U15848 (N_15848,N_13507,N_13846);
or U15849 (N_15849,N_14834,N_14497);
xnor U15850 (N_15850,N_13326,N_13051);
xnor U15851 (N_15851,N_13589,N_13203);
nor U15852 (N_15852,N_12385,N_12730);
or U15853 (N_15853,N_14798,N_13054);
xnor U15854 (N_15854,N_12839,N_13868);
nor U15855 (N_15855,N_14196,N_14749);
nor U15856 (N_15856,N_14248,N_14964);
nor U15857 (N_15857,N_13284,N_13716);
or U15858 (N_15858,N_13535,N_14800);
or U15859 (N_15859,N_12352,N_13304);
or U15860 (N_15860,N_14779,N_13105);
or U15861 (N_15861,N_14997,N_12544);
and U15862 (N_15862,N_13351,N_13687);
or U15863 (N_15863,N_13323,N_14111);
xnor U15864 (N_15864,N_12392,N_13903);
or U15865 (N_15865,N_13970,N_12859);
or U15866 (N_15866,N_14944,N_14491);
xor U15867 (N_15867,N_12318,N_14346);
xnor U15868 (N_15868,N_13764,N_12049);
nand U15869 (N_15869,N_13499,N_13915);
xnor U15870 (N_15870,N_12931,N_14665);
xor U15871 (N_15871,N_12336,N_14753);
nand U15872 (N_15872,N_14465,N_13159);
nor U15873 (N_15873,N_12606,N_14986);
and U15874 (N_15874,N_14582,N_13256);
or U15875 (N_15875,N_12236,N_12030);
nor U15876 (N_15876,N_13359,N_12786);
nor U15877 (N_15877,N_12380,N_12370);
nor U15878 (N_15878,N_12475,N_14658);
and U15879 (N_15879,N_13834,N_12877);
nand U15880 (N_15880,N_13645,N_13890);
nor U15881 (N_15881,N_12034,N_12808);
or U15882 (N_15882,N_12433,N_12638);
or U15883 (N_15883,N_12811,N_12640);
and U15884 (N_15884,N_13554,N_14970);
nand U15885 (N_15885,N_12518,N_12262);
or U15886 (N_15886,N_13457,N_14258);
xor U15887 (N_15887,N_14560,N_13363);
nor U15888 (N_15888,N_14305,N_14086);
nor U15889 (N_15889,N_14708,N_12913);
nor U15890 (N_15890,N_14781,N_12923);
nand U15891 (N_15891,N_13637,N_13994);
xnor U15892 (N_15892,N_12083,N_14336);
and U15893 (N_15893,N_12695,N_12557);
and U15894 (N_15894,N_12530,N_13617);
nand U15895 (N_15895,N_13008,N_14616);
and U15896 (N_15896,N_13540,N_12541);
or U15897 (N_15897,N_12311,N_14461);
xnor U15898 (N_15898,N_13075,N_13318);
or U15899 (N_15899,N_14620,N_14068);
nor U15900 (N_15900,N_12341,N_12343);
xor U15901 (N_15901,N_14408,N_13316);
nand U15902 (N_15902,N_14645,N_13612);
and U15903 (N_15903,N_14424,N_14791);
xor U15904 (N_15904,N_14803,N_14319);
nor U15905 (N_15905,N_14553,N_14826);
or U15906 (N_15906,N_13472,N_12657);
nand U15907 (N_15907,N_13291,N_12575);
nor U15908 (N_15908,N_14431,N_12268);
or U15909 (N_15909,N_12001,N_13451);
nand U15910 (N_15910,N_12950,N_12739);
xnor U15911 (N_15911,N_13164,N_14447);
nand U15912 (N_15912,N_12725,N_12409);
or U15913 (N_15913,N_13044,N_12015);
nor U15914 (N_15914,N_13799,N_12728);
and U15915 (N_15915,N_12927,N_12873);
nand U15916 (N_15916,N_13052,N_14661);
nand U15917 (N_15917,N_14395,N_14681);
or U15918 (N_15918,N_13269,N_12104);
xnor U15919 (N_15919,N_13350,N_12414);
or U15920 (N_15920,N_13201,N_14098);
nor U15921 (N_15921,N_12445,N_12585);
and U15922 (N_15922,N_14477,N_13213);
or U15923 (N_15923,N_13474,N_13124);
nor U15924 (N_15924,N_14398,N_13222);
or U15925 (N_15925,N_13665,N_13659);
xnor U15926 (N_15926,N_13215,N_14112);
or U15927 (N_15927,N_13933,N_12451);
and U15928 (N_15928,N_14064,N_13878);
nand U15929 (N_15929,N_14557,N_13982);
xor U15930 (N_15930,N_14670,N_12801);
nand U15931 (N_15931,N_12724,N_12167);
xor U15932 (N_15932,N_14399,N_12071);
and U15933 (N_15933,N_14870,N_14007);
nor U15934 (N_15934,N_14177,N_14577);
nor U15935 (N_15935,N_13734,N_14638);
or U15936 (N_15936,N_14455,N_13949);
nor U15937 (N_15937,N_12077,N_13172);
xnor U15938 (N_15938,N_13824,N_13071);
or U15939 (N_15939,N_14012,N_14558);
xor U15940 (N_15940,N_14032,N_14433);
nor U15941 (N_15941,N_13253,N_13223);
nand U15942 (N_15942,N_13847,N_12767);
xnor U15943 (N_15943,N_13785,N_13525);
nand U15944 (N_15944,N_12513,N_13574);
and U15945 (N_15945,N_12681,N_12224);
xor U15946 (N_15946,N_13628,N_12784);
nand U15947 (N_15947,N_14628,N_12512);
and U15948 (N_15948,N_14829,N_14118);
or U15949 (N_15949,N_12120,N_13289);
or U15950 (N_15950,N_12485,N_14525);
nand U15951 (N_15951,N_12875,N_14672);
nand U15952 (N_15952,N_13295,N_13396);
nand U15953 (N_15953,N_13060,N_12500);
nor U15954 (N_15954,N_12763,N_12696);
xnor U15955 (N_15955,N_14402,N_14586);
nor U15956 (N_15956,N_13395,N_12529);
or U15957 (N_15957,N_13109,N_12822);
and U15958 (N_15958,N_14830,N_13475);
nand U15959 (N_15959,N_14641,N_14892);
nor U15960 (N_15960,N_13084,N_13381);
nand U15961 (N_15961,N_14540,N_14576);
nand U15962 (N_15962,N_12993,N_13696);
and U15963 (N_15963,N_12896,N_12731);
or U15964 (N_15964,N_14673,N_14775);
nand U15965 (N_15965,N_14814,N_14294);
and U15966 (N_15966,N_14585,N_14458);
xnor U15967 (N_15967,N_12319,N_14180);
or U15968 (N_15968,N_12139,N_13666);
and U15969 (N_15969,N_13210,N_14490);
and U15970 (N_15970,N_12543,N_13563);
and U15971 (N_15971,N_14095,N_14855);
nor U15972 (N_15972,N_13379,N_12215);
and U15973 (N_15973,N_13019,N_12391);
and U15974 (N_15974,N_14876,N_12013);
nand U15975 (N_15975,N_12624,N_12480);
and U15976 (N_15976,N_13860,N_13315);
and U15977 (N_15977,N_13184,N_14279);
nor U15978 (N_15978,N_14488,N_13276);
or U15979 (N_15979,N_13001,N_12802);
xnor U15980 (N_15980,N_14676,N_12740);
or U15981 (N_15981,N_12676,N_13874);
and U15982 (N_15982,N_12222,N_12690);
nand U15983 (N_15983,N_14743,N_12176);
xnor U15984 (N_15984,N_14512,N_14075);
and U15985 (N_15985,N_12191,N_12819);
xor U15986 (N_15986,N_13383,N_12805);
xor U15987 (N_15987,N_14246,N_14680);
xnor U15988 (N_15988,N_14769,N_12721);
nor U15989 (N_15989,N_14301,N_13277);
or U15990 (N_15990,N_14886,N_12579);
nand U15991 (N_15991,N_13059,N_13919);
or U15992 (N_15992,N_12874,N_12250);
and U15993 (N_15993,N_13317,N_12009);
xor U15994 (N_15994,N_12960,N_13926);
xor U15995 (N_15995,N_14442,N_13227);
and U15996 (N_15996,N_14044,N_13095);
xor U15997 (N_15997,N_13889,N_13842);
xnor U15998 (N_15998,N_12642,N_14498);
and U15999 (N_15999,N_12526,N_14950);
xnor U16000 (N_16000,N_14355,N_12779);
or U16001 (N_16001,N_14265,N_12581);
xnor U16002 (N_16002,N_14061,N_12463);
nor U16003 (N_16003,N_14430,N_13362);
nand U16004 (N_16004,N_13119,N_14422);
xor U16005 (N_16005,N_14820,N_12478);
and U16006 (N_16006,N_13146,N_14306);
nand U16007 (N_16007,N_13845,N_13992);
nand U16008 (N_16008,N_12694,N_13380);
nand U16009 (N_16009,N_13614,N_13548);
and U16010 (N_16010,N_14724,N_12084);
nand U16011 (N_16011,N_14866,N_13516);
or U16012 (N_16012,N_14054,N_12323);
or U16013 (N_16013,N_14664,N_13671);
xor U16014 (N_16014,N_12276,N_12458);
or U16015 (N_16015,N_14307,N_12616);
nor U16016 (N_16016,N_13127,N_14014);
and U16017 (N_16017,N_12166,N_14138);
and U16018 (N_16018,N_12205,N_12488);
or U16019 (N_16019,N_13408,N_12294);
or U16020 (N_16020,N_13388,N_12201);
nand U16021 (N_16021,N_12314,N_13034);
or U16022 (N_16022,N_14801,N_12520);
xnor U16023 (N_16023,N_12604,N_12455);
nand U16024 (N_16024,N_12745,N_14168);
xor U16025 (N_16025,N_12871,N_12782);
nand U16026 (N_16026,N_14727,N_14518);
xnor U16027 (N_16027,N_13578,N_13638);
nand U16028 (N_16028,N_12965,N_14360);
xnor U16029 (N_16029,N_13798,N_14410);
and U16030 (N_16030,N_13221,N_13400);
and U16031 (N_16031,N_12850,N_14191);
xor U16032 (N_16032,N_14448,N_12354);
and U16033 (N_16033,N_14821,N_13859);
and U16034 (N_16034,N_13862,N_14243);
or U16035 (N_16035,N_13958,N_14469);
nand U16036 (N_16036,N_13811,N_14271);
nand U16037 (N_16037,N_13338,N_13534);
nor U16038 (N_16038,N_14343,N_13429);
nor U16039 (N_16039,N_14065,N_13683);
nand U16040 (N_16040,N_13486,N_14519);
nand U16041 (N_16041,N_12570,N_13041);
nand U16042 (N_16042,N_12418,N_14720);
and U16043 (N_16043,N_12383,N_14572);
and U16044 (N_16044,N_12227,N_14510);
or U16045 (N_16045,N_13258,N_13988);
nand U16046 (N_16046,N_12940,N_13815);
xnor U16047 (N_16047,N_12287,N_12716);
nor U16048 (N_16048,N_14484,N_12836);
or U16049 (N_16049,N_13940,N_12291);
nor U16050 (N_16050,N_14372,N_13447);
xnor U16051 (N_16051,N_12329,N_13244);
nor U16052 (N_16052,N_13197,N_14409);
nand U16053 (N_16053,N_12364,N_14600);
nand U16054 (N_16054,N_14556,N_13401);
nor U16055 (N_16055,N_13924,N_12860);
nor U16056 (N_16056,N_14832,N_12547);
or U16057 (N_16057,N_13449,N_12916);
xor U16058 (N_16058,N_13373,N_14339);
or U16059 (N_16059,N_14211,N_13895);
and U16060 (N_16060,N_14293,N_12615);
nand U16061 (N_16061,N_12146,N_12333);
and U16062 (N_16062,N_14548,N_14764);
and U16063 (N_16063,N_14574,N_13107);
or U16064 (N_16064,N_12054,N_13086);
xor U16065 (N_16065,N_14859,N_13069);
and U16066 (N_16066,N_14544,N_13420);
and U16067 (N_16067,N_14239,N_13743);
or U16068 (N_16068,N_13991,N_12310);
and U16069 (N_16069,N_12044,N_12713);
nand U16070 (N_16070,N_13892,N_14259);
nand U16071 (N_16071,N_13238,N_13630);
nor U16072 (N_16072,N_13530,N_14136);
or U16073 (N_16073,N_12419,N_13707);
xnor U16074 (N_16074,N_12550,N_14992);
nor U16075 (N_16075,N_13131,N_14788);
and U16076 (N_16076,N_12476,N_13185);
or U16077 (N_16077,N_14806,N_12303);
nand U16078 (N_16078,N_13435,N_14495);
nor U16079 (N_16079,N_12442,N_13818);
nor U16080 (N_16080,N_14087,N_14142);
nor U16081 (N_16081,N_14648,N_12930);
and U16082 (N_16082,N_12082,N_12535);
nand U16083 (N_16083,N_14287,N_14927);
nand U16084 (N_16084,N_12144,N_13102);
nor U16085 (N_16085,N_12824,N_14610);
xnor U16086 (N_16086,N_14746,N_13074);
nor U16087 (N_16087,N_14439,N_12183);
nand U16088 (N_16088,N_13783,N_12219);
nand U16089 (N_16089,N_12359,N_13996);
xnor U16090 (N_16090,N_12639,N_13774);
and U16091 (N_16091,N_14421,N_14194);
or U16092 (N_16092,N_12774,N_12804);
or U16093 (N_16093,N_14515,N_13505);
or U16094 (N_16094,N_13207,N_14369);
and U16095 (N_16095,N_14285,N_12123);
nand U16096 (N_16096,N_12587,N_13969);
or U16097 (N_16097,N_13682,N_12641);
xnor U16098 (N_16098,N_12852,N_14485);
nor U16099 (N_16099,N_14601,N_12195);
xnor U16100 (N_16100,N_14021,N_14717);
or U16101 (N_16101,N_12067,N_14147);
nand U16102 (N_16102,N_13553,N_14116);
or U16103 (N_16103,N_14931,N_14561);
nor U16104 (N_16104,N_12554,N_14240);
xor U16105 (N_16105,N_12650,N_13048);
nor U16106 (N_16106,N_13032,N_14611);
nor U16107 (N_16107,N_12239,N_13871);
and U16108 (N_16108,N_14262,N_13590);
nand U16109 (N_16109,N_12760,N_12749);
nand U16110 (N_16110,N_13392,N_13832);
and U16111 (N_16111,N_12005,N_12427);
xor U16112 (N_16112,N_12757,N_12207);
and U16113 (N_16113,N_13155,N_12101);
and U16114 (N_16114,N_14797,N_14051);
nor U16115 (N_16115,N_13616,N_13394);
nand U16116 (N_16116,N_14990,N_13807);
nor U16117 (N_16117,N_14451,N_12230);
xor U16118 (N_16118,N_14072,N_12783);
or U16119 (N_16119,N_14178,N_14291);
xor U16120 (N_16120,N_13121,N_14358);
nand U16121 (N_16121,N_14219,N_12313);
and U16122 (N_16122,N_14078,N_14700);
xor U16123 (N_16123,N_14836,N_13644);
nor U16124 (N_16124,N_14195,N_12160);
and U16125 (N_16125,N_12413,N_14844);
xor U16126 (N_16126,N_13893,N_14917);
or U16127 (N_16127,N_12817,N_12212);
or U16128 (N_16128,N_12460,N_13839);
nor U16129 (N_16129,N_13427,N_14691);
nor U16130 (N_16130,N_14332,N_14849);
and U16131 (N_16131,N_12214,N_12800);
or U16132 (N_16132,N_13911,N_12194);
and U16133 (N_16133,N_13165,N_14320);
nor U16134 (N_16134,N_12596,N_12632);
xor U16135 (N_16135,N_13387,N_14812);
and U16136 (N_16136,N_13922,N_12406);
nand U16137 (N_16137,N_14023,N_13192);
nand U16138 (N_16138,N_13983,N_12803);
nand U16139 (N_16139,N_13704,N_14170);
xor U16140 (N_16140,N_12226,N_12888);
or U16141 (N_16141,N_14715,N_13470);
or U16142 (N_16142,N_13282,N_12157);
nor U16143 (N_16143,N_12260,N_13984);
xnor U16144 (N_16144,N_14471,N_14154);
nor U16145 (N_16145,N_14309,N_12985);
and U16146 (N_16146,N_12327,N_13004);
and U16147 (N_16147,N_12426,N_14404);
and U16148 (N_16148,N_13705,N_14900);
xor U16149 (N_16149,N_12466,N_13299);
xor U16150 (N_16150,N_13848,N_12769);
nor U16151 (N_16151,N_13344,N_12988);
nor U16152 (N_16152,N_13897,N_13183);
nand U16153 (N_16153,N_13082,N_13273);
xnor U16154 (N_16154,N_13492,N_12443);
nor U16155 (N_16155,N_13613,N_12069);
and U16156 (N_16156,N_13611,N_13055);
nor U16157 (N_16157,N_14919,N_13521);
nor U16158 (N_16158,N_14205,N_14302);
nor U16159 (N_16159,N_13793,N_12395);
nand U16160 (N_16160,N_14928,N_13483);
nand U16161 (N_16161,N_13319,N_12216);
nor U16162 (N_16162,N_13575,N_14031);
and U16163 (N_16163,N_12789,N_12958);
or U16164 (N_16164,N_13695,N_13509);
xor U16165 (N_16165,N_14909,N_13927);
and U16166 (N_16166,N_12479,N_14364);
or U16167 (N_16167,N_12127,N_13797);
xnor U16168 (N_16168,N_13496,N_12777);
nand U16169 (N_16169,N_12470,N_12944);
and U16170 (N_16170,N_13043,N_12133);
nand U16171 (N_16171,N_13434,N_13287);
nand U16172 (N_16172,N_14854,N_13403);
nor U16173 (N_16173,N_14359,N_12510);
xor U16174 (N_16174,N_12743,N_14564);
xor U16175 (N_16175,N_14035,N_14881);
nand U16176 (N_16176,N_13296,N_12053);
xor U16177 (N_16177,N_13558,N_14602);
or U16178 (N_16178,N_13422,N_12102);
xor U16179 (N_16179,N_13829,N_12162);
xor U16180 (N_16180,N_14973,N_14547);
xor U16181 (N_16181,N_12502,N_13600);
xor U16182 (N_16182,N_13342,N_14555);
nand U16183 (N_16183,N_14502,N_13661);
xnor U16184 (N_16184,N_12465,N_14889);
or U16185 (N_16185,N_14121,N_13283);
and U16186 (N_16186,N_13063,N_13000);
or U16187 (N_16187,N_13375,N_14254);
nand U16188 (N_16188,N_14752,N_14053);
nand U16189 (N_16189,N_12351,N_12161);
nor U16190 (N_16190,N_14754,N_13784);
nand U16191 (N_16191,N_13854,N_12307);
nand U16192 (N_16192,N_13441,N_14706);
and U16193 (N_16193,N_14837,N_14071);
xor U16194 (N_16194,N_13254,N_13346);
nor U16195 (N_16195,N_12766,N_14621);
or U16196 (N_16196,N_12892,N_12828);
or U16197 (N_16197,N_12678,N_13077);
nor U16198 (N_16198,N_12211,N_13733);
xor U16199 (N_16199,N_13955,N_12945);
or U16200 (N_16200,N_13372,N_14699);
or U16201 (N_16201,N_12595,N_13376);
or U16202 (N_16202,N_14635,N_14242);
and U16203 (N_16203,N_12116,N_13478);
nand U16204 (N_16204,N_13538,N_12499);
xor U16205 (N_16205,N_12780,N_13112);
nor U16206 (N_16206,N_13397,N_14423);
and U16207 (N_16207,N_13587,N_14627);
or U16208 (N_16208,N_12688,N_14079);
xnor U16209 (N_16209,N_13841,N_13971);
xnor U16210 (N_16210,N_13125,N_12798);
nand U16211 (N_16211,N_12159,N_12324);
and U16212 (N_16212,N_14546,N_12553);
and U16213 (N_16213,N_12880,N_13236);
or U16214 (N_16214,N_12251,N_14234);
or U16215 (N_16215,N_14507,N_14983);
nand U16216 (N_16216,N_14597,N_14057);
nor U16217 (N_16217,N_12103,N_14005);
nor U16218 (N_16218,N_13643,N_12891);
nor U16219 (N_16219,N_13662,N_13898);
xor U16220 (N_16220,N_14157,N_14912);
xor U16221 (N_16221,N_14083,N_12188);
xor U16222 (N_16222,N_12228,N_13914);
nor U16223 (N_16223,N_13108,N_12813);
xnor U16224 (N_16224,N_12572,N_14001);
and U16225 (N_16225,N_14568,N_13418);
or U16226 (N_16226,N_12665,N_13294);
nand U16227 (N_16227,N_14867,N_14322);
nand U16228 (N_16228,N_13341,N_12278);
xnor U16229 (N_16229,N_13963,N_13021);
nor U16230 (N_16230,N_13193,N_13667);
nand U16231 (N_16231,N_14996,N_14401);
nor U16232 (N_16232,N_13609,N_14368);
or U16233 (N_16233,N_14580,N_12337);
xor U16234 (N_16234,N_14895,N_14241);
or U16235 (N_16235,N_13309,N_12172);
or U16236 (N_16236,N_13501,N_14864);
or U16237 (N_16237,N_14407,N_13523);
nand U16238 (N_16238,N_12834,N_14549);
and U16239 (N_16239,N_13931,N_14009);
or U16240 (N_16240,N_12492,N_14807);
nor U16241 (N_16241,N_14025,N_14419);
nand U16242 (N_16242,N_12066,N_12088);
and U16243 (N_16243,N_14978,N_13560);
nor U16244 (N_16244,N_12113,N_12943);
xor U16245 (N_16245,N_12542,N_12298);
or U16246 (N_16246,N_14653,N_13313);
xor U16247 (N_16247,N_13800,N_14770);
nor U16248 (N_16248,N_13134,N_12991);
xnor U16249 (N_16249,N_14416,N_13028);
or U16250 (N_16250,N_14903,N_12719);
and U16251 (N_16251,N_14217,N_13445);
nor U16252 (N_16252,N_13096,N_12720);
and U16253 (N_16253,N_12914,N_12484);
and U16254 (N_16254,N_14333,N_12265);
xor U16255 (N_16255,N_14040,N_12605);
and U16256 (N_16256,N_12284,N_13905);
xor U16257 (N_16257,N_14562,N_12661);
nand U16258 (N_16258,N_14109,N_12301);
nand U16259 (N_16259,N_13115,N_14384);
and U16260 (N_16260,N_14683,N_12847);
xor U16261 (N_16261,N_14058,N_14288);
and U16262 (N_16262,N_14984,N_14171);
nor U16263 (N_16263,N_14933,N_12075);
and U16264 (N_16264,N_13776,N_13158);
xnor U16265 (N_16265,N_14907,N_13928);
or U16266 (N_16266,N_13654,N_14464);
nor U16267 (N_16267,N_13040,N_12121);
nand U16268 (N_16268,N_14533,N_12974);
xnor U16269 (N_16269,N_12978,N_12482);
nand U16270 (N_16270,N_12295,N_12052);
and U16271 (N_16271,N_12269,N_13138);
nand U16272 (N_16272,N_13355,N_12241);
nor U16273 (N_16273,N_13479,N_14923);
xnor U16274 (N_16274,N_14396,N_13466);
and U16275 (N_16275,N_12405,N_13706);
nand U16276 (N_16276,N_14221,N_12697);
nand U16277 (N_16277,N_12741,N_13702);
or U16278 (N_16278,N_14350,N_14713);
nor U16279 (N_16279,N_14159,N_13009);
or U16280 (N_16280,N_14153,N_12450);
and U16281 (N_16281,N_12316,N_12569);
nand U16282 (N_16282,N_13456,N_13951);
or U16283 (N_16283,N_13689,N_14414);
nand U16284 (N_16284,N_14010,N_14879);
nor U16285 (N_16285,N_13959,N_13038);
xnor U16286 (N_16286,N_14212,N_14761);
nor U16287 (N_16287,N_12288,N_14365);
nand U16288 (N_16288,N_12495,N_12523);
xor U16289 (N_16289,N_13536,N_13773);
or U16290 (N_16290,N_14898,N_14128);
and U16291 (N_16291,N_13663,N_14226);
xnor U16292 (N_16292,N_14452,N_12522);
and U16293 (N_16293,N_13694,N_12545);
and U16294 (N_16294,N_12806,N_13015);
or U16295 (N_16295,N_12727,N_12552);
nand U16296 (N_16296,N_14283,N_12254);
and U16297 (N_16297,N_12909,N_13757);
nand U16298 (N_16298,N_14951,N_12738);
or U16299 (N_16299,N_14436,N_14578);
nor U16300 (N_16300,N_13365,N_14425);
nand U16301 (N_16301,N_13765,N_14649);
xnor U16302 (N_16302,N_12612,N_14737);
or U16303 (N_16303,N_12669,N_14974);
xnor U16304 (N_16304,N_14981,N_12778);
nand U16305 (N_16305,N_12861,N_13485);
xnor U16306 (N_16306,N_12243,N_12396);
xnor U16307 (N_16307,N_12221,N_12142);
nand U16308 (N_16308,N_13160,N_14508);
nand U16309 (N_16309,N_12707,N_13918);
and U16310 (N_16310,N_14200,N_13128);
xnor U16311 (N_16311,N_12966,N_13149);
xnor U16312 (N_16312,N_14070,N_14588);
and U16313 (N_16313,N_14707,N_13747);
nor U16314 (N_16314,N_13883,N_13141);
nor U16315 (N_16315,N_12645,N_12204);
xnor U16316 (N_16316,N_13462,N_14954);
nor U16317 (N_16317,N_14114,N_13369);
xnor U16318 (N_16318,N_12118,N_13693);
or U16319 (N_16319,N_13961,N_13314);
nand U16320 (N_16320,N_12610,N_12018);
or U16321 (N_16321,N_14165,N_13731);
or U16322 (N_16322,N_12209,N_13232);
xor U16323 (N_16323,N_14066,N_14959);
nand U16324 (N_16324,N_12902,N_14634);
nor U16325 (N_16325,N_14566,N_14987);
xor U16326 (N_16326,N_12334,N_13039);
and U16327 (N_16327,N_12474,N_12134);
xnor U16328 (N_16328,N_13668,N_13204);
xor U16329 (N_16329,N_12007,N_14172);
and U16330 (N_16330,N_12677,N_13715);
nor U16331 (N_16331,N_14152,N_13480);
xnor U16332 (N_16332,N_13202,N_12992);
nand U16333 (N_16333,N_12089,N_12489);
or U16334 (N_16334,N_14594,N_14385);
or U16335 (N_16335,N_13573,N_12603);
and U16336 (N_16336,N_14110,N_13117);
xnor U16337 (N_16337,N_13391,N_14563);
xor U16338 (N_16338,N_14131,N_14695);
or U16339 (N_16339,N_13135,N_12410);
nor U16340 (N_16340,N_13037,N_12714);
or U16341 (N_16341,N_12308,N_12907);
and U16342 (N_16342,N_14922,N_14348);
or U16343 (N_16343,N_14405,N_14878);
xnor U16344 (N_16344,N_13416,N_14218);
nand U16345 (N_16345,N_13838,N_14179);
xnor U16346 (N_16346,N_13260,N_13857);
nor U16347 (N_16347,N_14193,N_14377);
nor U16348 (N_16348,N_13012,N_14682);
nor U16349 (N_16349,N_12651,N_12438);
and U16350 (N_16350,N_13823,N_12471);
nand U16351 (N_16351,N_13461,N_13331);
nor U16352 (N_16352,N_12432,N_13194);
xor U16353 (N_16353,N_13753,N_12507);
nor U16354 (N_16354,N_14728,N_14391);
nand U16355 (N_16355,N_12868,N_13891);
nor U16356 (N_16356,N_12004,N_13583);
and U16357 (N_16357,N_14946,N_13067);
nor U16358 (N_16358,N_13732,N_12563);
nand U16359 (N_16359,N_14175,N_12126);
nor U16360 (N_16360,N_13374,N_12348);
or U16361 (N_16361,N_12179,N_13598);
and U16362 (N_16362,N_13740,N_12338);
nand U16363 (N_16363,N_12571,N_14224);
nand U16364 (N_16364,N_14081,N_14901);
or U16365 (N_16365,N_13556,N_13031);
nor U16366 (N_16366,N_12033,N_12131);
nor U16367 (N_16367,N_14327,N_12576);
and U16368 (N_16368,N_13211,N_14050);
or U16369 (N_16369,N_14034,N_14148);
xnor U16370 (N_16370,N_14918,N_13042);
nor U16371 (N_16371,N_14124,N_12682);
and U16372 (N_16372,N_13789,N_13262);
xor U16373 (N_16373,N_12876,N_14042);
and U16374 (N_16374,N_12568,N_13281);
nand U16375 (N_16375,N_12768,N_12130);
nand U16376 (N_16376,N_13510,N_14186);
and U16377 (N_16377,N_14976,N_12330);
nand U16378 (N_16378,N_13725,N_14289);
xor U16379 (N_16379,N_12820,N_14019);
nand U16380 (N_16380,N_14084,N_12501);
xnor U16381 (N_16381,N_13297,N_12422);
nor U16382 (N_16382,N_13425,N_12598);
xnor U16383 (N_16383,N_14310,N_13581);
nand U16384 (N_16384,N_14505,N_13205);
nor U16385 (N_16385,N_14668,N_14948);
nand U16386 (N_16386,N_13947,N_12532);
xnor U16387 (N_16387,N_13266,N_13328);
or U16388 (N_16388,N_12816,N_14636);
nor U16389 (N_16389,N_12586,N_13886);
or U16390 (N_16390,N_14902,N_12794);
xnor U16391 (N_16391,N_13148,N_12797);
xor U16392 (N_16392,N_12429,N_13894);
or U16393 (N_16393,N_12773,N_14633);
and U16394 (N_16394,N_12408,N_13555);
or U16395 (N_16395,N_13058,N_12178);
nand U16396 (N_16396,N_12199,N_13782);
xor U16397 (N_16397,N_14815,N_12667);
or U16398 (N_16398,N_14499,N_13473);
xor U16399 (N_16399,N_13975,N_14187);
nand U16400 (N_16400,N_12663,N_12097);
nor U16401 (N_16401,N_14313,N_13144);
nand U16402 (N_16402,N_12796,N_13828);
nor U16403 (N_16403,N_13312,N_12218);
xor U16404 (N_16404,N_12504,N_14483);
nand U16405 (N_16405,N_13524,N_12906);
and U16406 (N_16406,N_12664,N_13642);
nor U16407 (N_16407,N_12090,N_13412);
nand U16408 (N_16408,N_13006,N_13234);
or U16409 (N_16409,N_14158,N_12248);
nand U16410 (N_16410,N_13405,N_14848);
nor U16411 (N_16411,N_14076,N_13646);
xor U16412 (N_16412,N_12186,N_12622);
xnor U16413 (N_16413,N_12687,N_14474);
nor U16414 (N_16414,N_13407,N_13737);
nand U16415 (N_16415,N_14094,N_14251);
nor U16416 (N_16416,N_13078,N_12320);
and U16417 (N_16417,N_13741,N_12377);
and U16418 (N_16418,N_13867,N_13097);
nor U16419 (N_16419,N_12971,N_12911);
or U16420 (N_16420,N_13361,N_12573);
or U16421 (N_16421,N_13537,N_14268);
nor U16422 (N_16422,N_14619,N_14091);
nor U16423 (N_16423,N_12509,N_12289);
xor U16424 (N_16424,N_12106,N_12491);
nor U16425 (N_16425,N_14632,N_12145);
xor U16426 (N_16426,N_13543,N_13191);
xnor U16427 (N_16427,N_14792,N_14818);
nand U16428 (N_16428,N_13649,N_13497);
nor U16429 (N_16429,N_14311,N_12548);
xnor U16430 (N_16430,N_13803,N_14115);
nor U16431 (N_16431,N_12190,N_14504);
xor U16432 (N_16432,N_12995,N_14910);
and U16433 (N_16433,N_14786,N_14831);
nor U16434 (N_16434,N_14733,N_13904);
or U16435 (N_16435,N_13526,N_13090);
xor U16436 (N_16436,N_14943,N_13242);
nor U16437 (N_16437,N_14335,N_14751);
or U16438 (N_16438,N_12136,N_13263);
xor U16439 (N_16439,N_12003,N_13002);
xnor U16440 (N_16440,N_14141,N_14935);
nand U16441 (N_16441,N_12980,N_13576);
nor U16442 (N_16442,N_13592,N_14406);
xor U16443 (N_16443,N_12625,N_14074);
or U16444 (N_16444,N_13265,N_13393);
and U16445 (N_16445,N_12601,N_12915);
xor U16446 (N_16446,N_14122,N_14149);
nor U16447 (N_16447,N_12305,N_12253);
nor U16448 (N_16448,N_13713,N_12994);
nand U16449 (N_16449,N_12952,N_12979);
or U16450 (N_16450,N_12398,N_14956);
and U16451 (N_16451,N_13566,N_14225);
and U16452 (N_16452,N_13607,N_14127);
and U16453 (N_16453,N_13858,N_14182);
nor U16454 (N_16454,N_14840,N_13901);
and U16455 (N_16455,N_13864,N_13579);
xor U16456 (N_16456,N_13247,N_14808);
xor U16457 (N_16457,N_12068,N_12946);
nand U16458 (N_16458,N_12775,N_14656);
or U16459 (N_16459,N_12182,N_13490);
or U16460 (N_16460,N_14617,N_14822);
nand U16461 (N_16461,N_14473,N_14003);
xnor U16462 (N_16462,N_12376,N_14575);
or U16463 (N_16463,N_14872,N_14802);
or U16464 (N_16464,N_14386,N_13719);
and U16465 (N_16465,N_12386,N_12114);
and U16466 (N_16466,N_14478,N_14780);
xnor U16467 (N_16467,N_14690,N_12564);
nand U16468 (N_16468,N_12549,N_13133);
or U16469 (N_16469,N_13669,N_13366);
nand U16470 (N_16470,N_13110,N_12006);
nor U16471 (N_16471,N_12300,N_14618);
nand U16472 (N_16472,N_14145,N_13169);
nor U16473 (N_16473,N_12381,N_13404);
xor U16474 (N_16474,N_13214,N_13301);
or U16475 (N_16475,N_12948,N_12076);
nor U16476 (N_16476,N_14790,N_14215);
xnor U16477 (N_16477,N_12592,N_13306);
or U16478 (N_16478,N_14789,N_14466);
xor U16479 (N_16479,N_12516,N_13542);
and U16480 (N_16480,N_13826,N_13697);
or U16481 (N_16481,N_14721,N_13288);
nand U16482 (N_16482,N_14741,N_14969);
or U16483 (N_16483,N_13567,N_12374);
nand U16484 (N_16484,N_12152,N_12863);
and U16485 (N_16485,N_14615,N_14847);
nand U16486 (N_16486,N_12292,N_12652);
xor U16487 (N_16487,N_14982,N_13023);
and U16488 (N_16488,N_12434,N_12537);
and U16489 (N_16489,N_14833,N_12400);
and U16490 (N_16490,N_12929,N_12085);
xor U16491 (N_16491,N_14099,N_12799);
xor U16492 (N_16492,N_13438,N_13423);
and U16493 (N_16493,N_13884,N_13790);
or U16494 (N_16494,N_12729,N_13421);
nand U16495 (N_16495,N_14624,N_12155);
nor U16496 (N_16496,N_12588,N_14828);
xnor U16497 (N_16497,N_12390,N_12751);
nand U16498 (N_16498,N_13986,N_13245);
xnor U16499 (N_16499,N_14521,N_12435);
or U16500 (N_16500,N_14548,N_12235);
nand U16501 (N_16501,N_12013,N_13429);
xor U16502 (N_16502,N_13588,N_13835);
nor U16503 (N_16503,N_14012,N_14172);
and U16504 (N_16504,N_13148,N_12051);
nor U16505 (N_16505,N_14814,N_14577);
nand U16506 (N_16506,N_13892,N_14576);
nand U16507 (N_16507,N_14732,N_12795);
or U16508 (N_16508,N_12212,N_13923);
xnor U16509 (N_16509,N_14729,N_14085);
nand U16510 (N_16510,N_14491,N_14795);
or U16511 (N_16511,N_13455,N_14080);
nor U16512 (N_16512,N_12048,N_14697);
xor U16513 (N_16513,N_13778,N_12429);
nand U16514 (N_16514,N_14187,N_14013);
or U16515 (N_16515,N_13235,N_12107);
nor U16516 (N_16516,N_14955,N_12682);
nand U16517 (N_16517,N_13912,N_13939);
or U16518 (N_16518,N_13927,N_12992);
xor U16519 (N_16519,N_12694,N_14896);
or U16520 (N_16520,N_12765,N_13394);
nor U16521 (N_16521,N_14100,N_13969);
nor U16522 (N_16522,N_13708,N_13092);
xor U16523 (N_16523,N_12944,N_13994);
xnor U16524 (N_16524,N_14270,N_13485);
and U16525 (N_16525,N_13964,N_12616);
or U16526 (N_16526,N_14411,N_14935);
xnor U16527 (N_16527,N_13653,N_12876);
xnor U16528 (N_16528,N_14890,N_13875);
xor U16529 (N_16529,N_13241,N_13901);
nand U16530 (N_16530,N_13676,N_12184);
nor U16531 (N_16531,N_14712,N_12778);
nor U16532 (N_16532,N_12410,N_12037);
nand U16533 (N_16533,N_14860,N_13541);
or U16534 (N_16534,N_13875,N_12091);
xor U16535 (N_16535,N_12710,N_12594);
or U16536 (N_16536,N_13766,N_14953);
xnor U16537 (N_16537,N_14995,N_13588);
or U16538 (N_16538,N_12868,N_12609);
or U16539 (N_16539,N_14123,N_13097);
nand U16540 (N_16540,N_14988,N_13797);
xnor U16541 (N_16541,N_12230,N_12537);
nor U16542 (N_16542,N_13935,N_13235);
or U16543 (N_16543,N_14925,N_13612);
or U16544 (N_16544,N_13453,N_12148);
xor U16545 (N_16545,N_13548,N_14080);
xor U16546 (N_16546,N_14760,N_13398);
nor U16547 (N_16547,N_14354,N_13318);
or U16548 (N_16548,N_12164,N_12912);
and U16549 (N_16549,N_13953,N_14737);
and U16550 (N_16550,N_13453,N_14849);
xnor U16551 (N_16551,N_12726,N_13541);
nand U16552 (N_16552,N_14355,N_13597);
nor U16553 (N_16553,N_13116,N_14155);
and U16554 (N_16554,N_13435,N_12641);
or U16555 (N_16555,N_14316,N_12764);
nor U16556 (N_16556,N_12969,N_14770);
nand U16557 (N_16557,N_13554,N_14296);
nand U16558 (N_16558,N_13065,N_12806);
nor U16559 (N_16559,N_12823,N_12080);
and U16560 (N_16560,N_13784,N_13251);
nand U16561 (N_16561,N_13576,N_14162);
nand U16562 (N_16562,N_14279,N_14693);
or U16563 (N_16563,N_14631,N_13932);
or U16564 (N_16564,N_14589,N_13760);
or U16565 (N_16565,N_12194,N_14395);
xnor U16566 (N_16566,N_12076,N_13276);
xnor U16567 (N_16567,N_13237,N_12307);
or U16568 (N_16568,N_13841,N_13977);
or U16569 (N_16569,N_12851,N_12303);
nand U16570 (N_16570,N_13967,N_14740);
xor U16571 (N_16571,N_13525,N_13535);
nor U16572 (N_16572,N_14209,N_14158);
nand U16573 (N_16573,N_12875,N_12348);
or U16574 (N_16574,N_14900,N_12672);
xnor U16575 (N_16575,N_13496,N_14668);
or U16576 (N_16576,N_14069,N_14306);
and U16577 (N_16577,N_14715,N_12743);
xor U16578 (N_16578,N_13277,N_14555);
and U16579 (N_16579,N_12374,N_14708);
xnor U16580 (N_16580,N_12581,N_12867);
nor U16581 (N_16581,N_13687,N_12969);
nand U16582 (N_16582,N_13963,N_12679);
or U16583 (N_16583,N_13690,N_13598);
nand U16584 (N_16584,N_13127,N_13603);
and U16585 (N_16585,N_14035,N_14862);
nor U16586 (N_16586,N_13964,N_14141);
nor U16587 (N_16587,N_14259,N_13134);
nor U16588 (N_16588,N_12380,N_13638);
and U16589 (N_16589,N_13775,N_13203);
and U16590 (N_16590,N_13291,N_13330);
nand U16591 (N_16591,N_13597,N_13496);
and U16592 (N_16592,N_13466,N_14125);
xor U16593 (N_16593,N_12982,N_12794);
nand U16594 (N_16594,N_12382,N_14276);
nor U16595 (N_16595,N_14540,N_13668);
nand U16596 (N_16596,N_14325,N_12356);
nand U16597 (N_16597,N_13734,N_12595);
or U16598 (N_16598,N_13274,N_13927);
or U16599 (N_16599,N_14143,N_14674);
and U16600 (N_16600,N_14521,N_13412);
or U16601 (N_16601,N_14844,N_14576);
and U16602 (N_16602,N_12005,N_12192);
nand U16603 (N_16603,N_13269,N_13210);
nand U16604 (N_16604,N_13218,N_14066);
nand U16605 (N_16605,N_13603,N_14016);
nand U16606 (N_16606,N_13808,N_12458);
nor U16607 (N_16607,N_13682,N_14084);
nor U16608 (N_16608,N_13595,N_13011);
nor U16609 (N_16609,N_13804,N_12850);
nor U16610 (N_16610,N_14367,N_14728);
nor U16611 (N_16611,N_12338,N_13234);
xnor U16612 (N_16612,N_14919,N_14469);
and U16613 (N_16613,N_14754,N_14250);
nor U16614 (N_16614,N_12605,N_13566);
or U16615 (N_16615,N_14846,N_12338);
xnor U16616 (N_16616,N_12930,N_13377);
nand U16617 (N_16617,N_13673,N_13328);
nand U16618 (N_16618,N_12772,N_12085);
and U16619 (N_16619,N_13923,N_12785);
and U16620 (N_16620,N_14386,N_14619);
nor U16621 (N_16621,N_13023,N_14024);
xor U16622 (N_16622,N_12762,N_14167);
xor U16623 (N_16623,N_12972,N_12207);
nor U16624 (N_16624,N_14584,N_14896);
and U16625 (N_16625,N_12761,N_12216);
or U16626 (N_16626,N_13931,N_12673);
nor U16627 (N_16627,N_13656,N_13532);
and U16628 (N_16628,N_13810,N_13660);
and U16629 (N_16629,N_13199,N_12791);
nor U16630 (N_16630,N_13862,N_13471);
or U16631 (N_16631,N_14476,N_14338);
and U16632 (N_16632,N_14698,N_13821);
xor U16633 (N_16633,N_14424,N_14793);
or U16634 (N_16634,N_13578,N_12992);
and U16635 (N_16635,N_14837,N_13233);
xnor U16636 (N_16636,N_13101,N_12207);
nand U16637 (N_16637,N_14449,N_14487);
nor U16638 (N_16638,N_14820,N_13760);
nor U16639 (N_16639,N_12061,N_12580);
and U16640 (N_16640,N_14917,N_14645);
xor U16641 (N_16641,N_14337,N_12210);
nand U16642 (N_16642,N_13976,N_12696);
xnor U16643 (N_16643,N_14207,N_13589);
nand U16644 (N_16644,N_14895,N_14091);
or U16645 (N_16645,N_13710,N_14745);
and U16646 (N_16646,N_12101,N_12318);
nor U16647 (N_16647,N_14712,N_12066);
or U16648 (N_16648,N_13871,N_12423);
nand U16649 (N_16649,N_12247,N_13157);
xnor U16650 (N_16650,N_12388,N_14043);
or U16651 (N_16651,N_12339,N_12754);
or U16652 (N_16652,N_14747,N_13604);
or U16653 (N_16653,N_13266,N_12414);
xor U16654 (N_16654,N_14818,N_14537);
xnor U16655 (N_16655,N_13592,N_14107);
xnor U16656 (N_16656,N_12992,N_14592);
nor U16657 (N_16657,N_12374,N_12771);
or U16658 (N_16658,N_13109,N_12245);
xor U16659 (N_16659,N_13471,N_12272);
or U16660 (N_16660,N_14173,N_13219);
and U16661 (N_16661,N_12932,N_12672);
and U16662 (N_16662,N_12969,N_13753);
and U16663 (N_16663,N_14709,N_12363);
or U16664 (N_16664,N_13048,N_14668);
nor U16665 (N_16665,N_12443,N_13487);
xor U16666 (N_16666,N_14447,N_14966);
xor U16667 (N_16667,N_14383,N_13063);
nor U16668 (N_16668,N_12238,N_13093);
and U16669 (N_16669,N_13584,N_13192);
and U16670 (N_16670,N_13345,N_12395);
and U16671 (N_16671,N_13721,N_14625);
nor U16672 (N_16672,N_13406,N_14975);
nand U16673 (N_16673,N_14629,N_14408);
or U16674 (N_16674,N_12945,N_14826);
xor U16675 (N_16675,N_13499,N_13273);
and U16676 (N_16676,N_13607,N_13759);
or U16677 (N_16677,N_12200,N_12318);
nor U16678 (N_16678,N_12838,N_13662);
and U16679 (N_16679,N_14844,N_13951);
nand U16680 (N_16680,N_13272,N_12062);
xnor U16681 (N_16681,N_14043,N_13283);
and U16682 (N_16682,N_14088,N_13820);
xor U16683 (N_16683,N_14278,N_12066);
nand U16684 (N_16684,N_14770,N_12152);
nand U16685 (N_16685,N_12280,N_12124);
or U16686 (N_16686,N_13631,N_12844);
xor U16687 (N_16687,N_13684,N_13946);
and U16688 (N_16688,N_12951,N_14256);
and U16689 (N_16689,N_12767,N_13583);
or U16690 (N_16690,N_12823,N_14769);
or U16691 (N_16691,N_13617,N_12399);
or U16692 (N_16692,N_14980,N_14567);
nor U16693 (N_16693,N_12958,N_14060);
nand U16694 (N_16694,N_12802,N_13106);
nand U16695 (N_16695,N_13504,N_13178);
xnor U16696 (N_16696,N_13854,N_12840);
and U16697 (N_16697,N_12990,N_12732);
and U16698 (N_16698,N_12804,N_14747);
xnor U16699 (N_16699,N_12689,N_14771);
xor U16700 (N_16700,N_13613,N_13415);
and U16701 (N_16701,N_14318,N_12014);
xor U16702 (N_16702,N_13083,N_12679);
and U16703 (N_16703,N_14484,N_13597);
xnor U16704 (N_16704,N_13810,N_12065);
nor U16705 (N_16705,N_13066,N_14005);
nand U16706 (N_16706,N_14532,N_14217);
xor U16707 (N_16707,N_14022,N_13894);
nand U16708 (N_16708,N_12957,N_13392);
or U16709 (N_16709,N_13881,N_12793);
nor U16710 (N_16710,N_12307,N_13846);
nor U16711 (N_16711,N_12296,N_12114);
nor U16712 (N_16712,N_14824,N_12708);
or U16713 (N_16713,N_13059,N_13295);
xor U16714 (N_16714,N_13216,N_12068);
and U16715 (N_16715,N_14449,N_12488);
xnor U16716 (N_16716,N_13565,N_13935);
and U16717 (N_16717,N_12922,N_12862);
xnor U16718 (N_16718,N_13605,N_12969);
nand U16719 (N_16719,N_12713,N_12208);
and U16720 (N_16720,N_12987,N_12852);
nor U16721 (N_16721,N_13732,N_13299);
xnor U16722 (N_16722,N_13906,N_13146);
xor U16723 (N_16723,N_13045,N_13610);
xnor U16724 (N_16724,N_13611,N_13189);
xnor U16725 (N_16725,N_13444,N_14674);
and U16726 (N_16726,N_12062,N_13197);
xnor U16727 (N_16727,N_13983,N_12073);
nor U16728 (N_16728,N_14541,N_12191);
nor U16729 (N_16729,N_13915,N_12831);
and U16730 (N_16730,N_14763,N_12983);
nand U16731 (N_16731,N_13647,N_12975);
or U16732 (N_16732,N_12020,N_14947);
nor U16733 (N_16733,N_13400,N_13092);
nor U16734 (N_16734,N_14454,N_12665);
nand U16735 (N_16735,N_12879,N_14842);
nand U16736 (N_16736,N_14036,N_12857);
nand U16737 (N_16737,N_14398,N_12059);
nand U16738 (N_16738,N_12211,N_12344);
nor U16739 (N_16739,N_13569,N_14102);
and U16740 (N_16740,N_12505,N_13119);
nor U16741 (N_16741,N_12049,N_12016);
or U16742 (N_16742,N_14266,N_12255);
and U16743 (N_16743,N_14979,N_12884);
or U16744 (N_16744,N_13335,N_13297);
nand U16745 (N_16745,N_13681,N_12543);
nor U16746 (N_16746,N_13047,N_14801);
or U16747 (N_16747,N_14019,N_12703);
xor U16748 (N_16748,N_14305,N_13185);
nor U16749 (N_16749,N_12122,N_14845);
or U16750 (N_16750,N_14266,N_13001);
xnor U16751 (N_16751,N_13304,N_14838);
nor U16752 (N_16752,N_13310,N_13467);
nor U16753 (N_16753,N_12683,N_12016);
and U16754 (N_16754,N_13036,N_14023);
or U16755 (N_16755,N_12488,N_13053);
xnor U16756 (N_16756,N_12194,N_12877);
nand U16757 (N_16757,N_14844,N_14098);
and U16758 (N_16758,N_14581,N_14069);
xor U16759 (N_16759,N_12391,N_13224);
or U16760 (N_16760,N_14701,N_14647);
xor U16761 (N_16761,N_13889,N_12360);
xor U16762 (N_16762,N_13463,N_14776);
nor U16763 (N_16763,N_14004,N_14587);
nor U16764 (N_16764,N_13001,N_14842);
nor U16765 (N_16765,N_14208,N_14736);
xor U16766 (N_16766,N_13574,N_14374);
or U16767 (N_16767,N_13242,N_12399);
or U16768 (N_16768,N_14528,N_14955);
nor U16769 (N_16769,N_13029,N_14266);
or U16770 (N_16770,N_12406,N_14820);
xor U16771 (N_16771,N_14393,N_14127);
and U16772 (N_16772,N_13289,N_12739);
nand U16773 (N_16773,N_12385,N_13479);
nand U16774 (N_16774,N_14670,N_13438);
nand U16775 (N_16775,N_12434,N_13549);
xnor U16776 (N_16776,N_14357,N_13173);
nor U16777 (N_16777,N_13202,N_12705);
nand U16778 (N_16778,N_13462,N_13278);
nand U16779 (N_16779,N_12523,N_12598);
nand U16780 (N_16780,N_14581,N_13733);
nand U16781 (N_16781,N_13091,N_12727);
or U16782 (N_16782,N_12452,N_14094);
nor U16783 (N_16783,N_14519,N_13931);
nand U16784 (N_16784,N_14422,N_12641);
nand U16785 (N_16785,N_14250,N_13780);
or U16786 (N_16786,N_13079,N_14599);
nor U16787 (N_16787,N_13109,N_13610);
or U16788 (N_16788,N_13358,N_12891);
or U16789 (N_16789,N_12712,N_13097);
nand U16790 (N_16790,N_12366,N_12863);
nand U16791 (N_16791,N_13205,N_12931);
nand U16792 (N_16792,N_12490,N_12546);
nor U16793 (N_16793,N_12044,N_12369);
nor U16794 (N_16794,N_14094,N_14009);
xnor U16795 (N_16795,N_13710,N_14308);
nand U16796 (N_16796,N_12449,N_13342);
and U16797 (N_16797,N_13515,N_14019);
nand U16798 (N_16798,N_13129,N_14912);
and U16799 (N_16799,N_14977,N_13359);
nand U16800 (N_16800,N_14465,N_12684);
nand U16801 (N_16801,N_13559,N_13798);
and U16802 (N_16802,N_12377,N_14722);
xnor U16803 (N_16803,N_12534,N_14070);
or U16804 (N_16804,N_13765,N_13264);
nand U16805 (N_16805,N_13908,N_13294);
and U16806 (N_16806,N_13548,N_12634);
nand U16807 (N_16807,N_12993,N_12142);
or U16808 (N_16808,N_14827,N_13878);
nand U16809 (N_16809,N_13400,N_14693);
nor U16810 (N_16810,N_12324,N_12735);
and U16811 (N_16811,N_13678,N_14864);
nand U16812 (N_16812,N_14314,N_14759);
nand U16813 (N_16813,N_13640,N_14852);
nand U16814 (N_16814,N_14495,N_14961);
nor U16815 (N_16815,N_12724,N_13820);
or U16816 (N_16816,N_14439,N_14413);
or U16817 (N_16817,N_13436,N_12781);
or U16818 (N_16818,N_13911,N_14057);
xnor U16819 (N_16819,N_12929,N_14311);
and U16820 (N_16820,N_14838,N_12384);
nand U16821 (N_16821,N_14560,N_14847);
xnor U16822 (N_16822,N_12536,N_12184);
nand U16823 (N_16823,N_12795,N_13020);
nor U16824 (N_16824,N_14198,N_14119);
nand U16825 (N_16825,N_13917,N_14713);
or U16826 (N_16826,N_14438,N_12832);
or U16827 (N_16827,N_14865,N_13562);
nor U16828 (N_16828,N_12696,N_14476);
nor U16829 (N_16829,N_13015,N_13975);
nor U16830 (N_16830,N_14716,N_13266);
nand U16831 (N_16831,N_12554,N_13442);
nand U16832 (N_16832,N_13076,N_14198);
and U16833 (N_16833,N_12913,N_12504);
nor U16834 (N_16834,N_12194,N_13982);
and U16835 (N_16835,N_13180,N_14159);
nor U16836 (N_16836,N_13005,N_14295);
nand U16837 (N_16837,N_13904,N_13172);
and U16838 (N_16838,N_13108,N_14620);
xnor U16839 (N_16839,N_14381,N_12689);
and U16840 (N_16840,N_13391,N_13005);
xnor U16841 (N_16841,N_13662,N_12042);
or U16842 (N_16842,N_12870,N_12183);
nor U16843 (N_16843,N_12123,N_13251);
and U16844 (N_16844,N_12723,N_12604);
nor U16845 (N_16845,N_13955,N_14345);
and U16846 (N_16846,N_12410,N_13505);
and U16847 (N_16847,N_12259,N_13610);
or U16848 (N_16848,N_13504,N_13582);
nor U16849 (N_16849,N_13020,N_13802);
nor U16850 (N_16850,N_12027,N_13966);
and U16851 (N_16851,N_13426,N_12764);
and U16852 (N_16852,N_12990,N_14000);
and U16853 (N_16853,N_12276,N_13168);
and U16854 (N_16854,N_14447,N_13749);
xnor U16855 (N_16855,N_12583,N_12763);
nor U16856 (N_16856,N_12404,N_13464);
nor U16857 (N_16857,N_13659,N_12227);
nor U16858 (N_16858,N_14014,N_12521);
nand U16859 (N_16859,N_13559,N_14665);
nor U16860 (N_16860,N_14535,N_14069);
nor U16861 (N_16861,N_14468,N_12386);
and U16862 (N_16862,N_14746,N_12351);
or U16863 (N_16863,N_14203,N_14111);
or U16864 (N_16864,N_12111,N_13730);
and U16865 (N_16865,N_13969,N_13073);
nor U16866 (N_16866,N_13718,N_12475);
and U16867 (N_16867,N_14177,N_12981);
xor U16868 (N_16868,N_13397,N_12005);
nand U16869 (N_16869,N_14331,N_14600);
or U16870 (N_16870,N_14720,N_13960);
xnor U16871 (N_16871,N_12686,N_12862);
nand U16872 (N_16872,N_14516,N_14486);
or U16873 (N_16873,N_14060,N_12782);
xor U16874 (N_16874,N_12818,N_12132);
and U16875 (N_16875,N_12638,N_13660);
or U16876 (N_16876,N_12628,N_12033);
nor U16877 (N_16877,N_13078,N_12162);
nand U16878 (N_16878,N_13039,N_12283);
and U16879 (N_16879,N_14634,N_14153);
nor U16880 (N_16880,N_12591,N_12833);
nor U16881 (N_16881,N_13364,N_14791);
or U16882 (N_16882,N_14247,N_12835);
nor U16883 (N_16883,N_14887,N_14100);
xor U16884 (N_16884,N_13831,N_12125);
nor U16885 (N_16885,N_14915,N_14944);
nand U16886 (N_16886,N_14904,N_13406);
nand U16887 (N_16887,N_13347,N_14939);
xnor U16888 (N_16888,N_12178,N_13442);
nor U16889 (N_16889,N_13681,N_13706);
and U16890 (N_16890,N_14021,N_12761);
and U16891 (N_16891,N_13181,N_13327);
or U16892 (N_16892,N_13684,N_14234);
nand U16893 (N_16893,N_12383,N_13587);
or U16894 (N_16894,N_14456,N_14176);
and U16895 (N_16895,N_14443,N_13125);
xnor U16896 (N_16896,N_12186,N_13329);
xnor U16897 (N_16897,N_14707,N_13144);
nand U16898 (N_16898,N_12344,N_13061);
nand U16899 (N_16899,N_14594,N_13471);
nand U16900 (N_16900,N_13708,N_13409);
nand U16901 (N_16901,N_12114,N_14882);
nand U16902 (N_16902,N_13258,N_12647);
xnor U16903 (N_16903,N_12317,N_13851);
and U16904 (N_16904,N_13646,N_13059);
xor U16905 (N_16905,N_12458,N_14234);
and U16906 (N_16906,N_12300,N_12428);
xnor U16907 (N_16907,N_14165,N_13797);
nand U16908 (N_16908,N_14832,N_14067);
nor U16909 (N_16909,N_14834,N_14040);
nor U16910 (N_16910,N_13679,N_12794);
xnor U16911 (N_16911,N_14221,N_14172);
or U16912 (N_16912,N_14702,N_14427);
xor U16913 (N_16913,N_14587,N_14692);
and U16914 (N_16914,N_12676,N_13156);
and U16915 (N_16915,N_13205,N_14719);
nand U16916 (N_16916,N_13888,N_14679);
nor U16917 (N_16917,N_13520,N_12239);
nor U16918 (N_16918,N_12819,N_13994);
or U16919 (N_16919,N_12877,N_12436);
nor U16920 (N_16920,N_14349,N_14663);
xor U16921 (N_16921,N_12708,N_12529);
xnor U16922 (N_16922,N_13645,N_13221);
or U16923 (N_16923,N_14406,N_13184);
or U16924 (N_16924,N_13881,N_13552);
nor U16925 (N_16925,N_14746,N_12827);
or U16926 (N_16926,N_14132,N_12795);
nor U16927 (N_16927,N_12997,N_12515);
xor U16928 (N_16928,N_14181,N_12708);
nand U16929 (N_16929,N_14389,N_14644);
xor U16930 (N_16930,N_12759,N_12721);
xnor U16931 (N_16931,N_13866,N_12401);
xor U16932 (N_16932,N_13842,N_12467);
or U16933 (N_16933,N_12057,N_13040);
nand U16934 (N_16934,N_14712,N_13564);
or U16935 (N_16935,N_14703,N_12534);
nor U16936 (N_16936,N_13258,N_12293);
and U16937 (N_16937,N_13500,N_13050);
and U16938 (N_16938,N_12274,N_13430);
nand U16939 (N_16939,N_14101,N_13813);
nor U16940 (N_16940,N_14276,N_14027);
xor U16941 (N_16941,N_12381,N_13674);
xor U16942 (N_16942,N_12009,N_12760);
and U16943 (N_16943,N_13916,N_13250);
nor U16944 (N_16944,N_13286,N_14773);
nand U16945 (N_16945,N_12090,N_12467);
or U16946 (N_16946,N_13544,N_13027);
or U16947 (N_16947,N_14750,N_12852);
xor U16948 (N_16948,N_14154,N_14563);
and U16949 (N_16949,N_13429,N_14020);
nor U16950 (N_16950,N_14806,N_13987);
nor U16951 (N_16951,N_12953,N_13926);
and U16952 (N_16952,N_14298,N_12941);
and U16953 (N_16953,N_13879,N_12049);
or U16954 (N_16954,N_14619,N_12114);
and U16955 (N_16955,N_13056,N_14291);
xnor U16956 (N_16956,N_12991,N_14711);
nor U16957 (N_16957,N_13376,N_12685);
or U16958 (N_16958,N_14977,N_12145);
and U16959 (N_16959,N_14609,N_13638);
nor U16960 (N_16960,N_13053,N_12241);
and U16961 (N_16961,N_14701,N_12245);
and U16962 (N_16962,N_12248,N_12933);
nand U16963 (N_16963,N_12628,N_12382);
nand U16964 (N_16964,N_13095,N_12659);
nor U16965 (N_16965,N_12957,N_14384);
nor U16966 (N_16966,N_14016,N_12226);
and U16967 (N_16967,N_14154,N_13812);
nor U16968 (N_16968,N_14785,N_14821);
and U16969 (N_16969,N_13089,N_13301);
and U16970 (N_16970,N_13305,N_12379);
or U16971 (N_16971,N_12633,N_14138);
nor U16972 (N_16972,N_12438,N_14809);
and U16973 (N_16973,N_14124,N_12536);
nand U16974 (N_16974,N_12454,N_12559);
and U16975 (N_16975,N_12487,N_13147);
nor U16976 (N_16976,N_13181,N_14306);
or U16977 (N_16977,N_14696,N_13370);
nor U16978 (N_16978,N_12613,N_13909);
and U16979 (N_16979,N_13019,N_14429);
and U16980 (N_16980,N_14848,N_14929);
nor U16981 (N_16981,N_14760,N_13941);
nand U16982 (N_16982,N_14965,N_14724);
nor U16983 (N_16983,N_12888,N_14297);
and U16984 (N_16984,N_14535,N_13084);
and U16985 (N_16985,N_14138,N_12210);
or U16986 (N_16986,N_14713,N_12111);
nand U16987 (N_16987,N_12955,N_14049);
nand U16988 (N_16988,N_14082,N_12026);
nand U16989 (N_16989,N_13696,N_12883);
and U16990 (N_16990,N_14561,N_12350);
nor U16991 (N_16991,N_13621,N_13177);
nand U16992 (N_16992,N_12928,N_12578);
or U16993 (N_16993,N_13656,N_13772);
nor U16994 (N_16994,N_14085,N_12815);
xnor U16995 (N_16995,N_12889,N_12543);
or U16996 (N_16996,N_13858,N_14136);
nand U16997 (N_16997,N_12375,N_14965);
xor U16998 (N_16998,N_13783,N_13406);
or U16999 (N_16999,N_13223,N_14919);
or U17000 (N_17000,N_13788,N_12450);
nand U17001 (N_17001,N_14232,N_14099);
xnor U17002 (N_17002,N_14825,N_14647);
and U17003 (N_17003,N_14853,N_12480);
and U17004 (N_17004,N_12794,N_14076);
and U17005 (N_17005,N_14011,N_13612);
nand U17006 (N_17006,N_13188,N_13540);
nand U17007 (N_17007,N_14859,N_13472);
xnor U17008 (N_17008,N_14853,N_12255);
nor U17009 (N_17009,N_12500,N_12360);
and U17010 (N_17010,N_13574,N_13691);
nor U17011 (N_17011,N_14723,N_12045);
and U17012 (N_17012,N_13372,N_12749);
or U17013 (N_17013,N_12310,N_12102);
or U17014 (N_17014,N_14104,N_14031);
nor U17015 (N_17015,N_14205,N_12735);
nor U17016 (N_17016,N_13421,N_13214);
nor U17017 (N_17017,N_14328,N_14357);
and U17018 (N_17018,N_12673,N_12421);
nand U17019 (N_17019,N_12585,N_12956);
nor U17020 (N_17020,N_14299,N_13435);
and U17021 (N_17021,N_14778,N_14564);
nand U17022 (N_17022,N_14101,N_12458);
xor U17023 (N_17023,N_13088,N_13053);
nor U17024 (N_17024,N_12836,N_12268);
and U17025 (N_17025,N_12396,N_13168);
or U17026 (N_17026,N_14929,N_12099);
or U17027 (N_17027,N_14386,N_12623);
xor U17028 (N_17028,N_12123,N_13123);
or U17029 (N_17029,N_12821,N_14236);
or U17030 (N_17030,N_14146,N_12226);
nor U17031 (N_17031,N_12401,N_12549);
xnor U17032 (N_17032,N_12138,N_13153);
nor U17033 (N_17033,N_13329,N_14328);
or U17034 (N_17034,N_12669,N_12581);
nand U17035 (N_17035,N_12769,N_13402);
nand U17036 (N_17036,N_13836,N_13091);
xnor U17037 (N_17037,N_14977,N_14205);
or U17038 (N_17038,N_14720,N_14043);
nand U17039 (N_17039,N_13249,N_13310);
or U17040 (N_17040,N_12485,N_12398);
nand U17041 (N_17041,N_14596,N_12196);
nand U17042 (N_17042,N_13270,N_12301);
and U17043 (N_17043,N_13450,N_14522);
nor U17044 (N_17044,N_14518,N_13113);
and U17045 (N_17045,N_12001,N_13422);
nor U17046 (N_17046,N_12449,N_14359);
or U17047 (N_17047,N_14836,N_13025);
nand U17048 (N_17048,N_14163,N_13866);
and U17049 (N_17049,N_13036,N_14550);
nor U17050 (N_17050,N_13555,N_13699);
nor U17051 (N_17051,N_14743,N_12318);
and U17052 (N_17052,N_14239,N_12303);
xor U17053 (N_17053,N_12252,N_13747);
nand U17054 (N_17054,N_12779,N_12646);
xnor U17055 (N_17055,N_14801,N_12511);
xnor U17056 (N_17056,N_13831,N_14891);
or U17057 (N_17057,N_12983,N_13751);
xnor U17058 (N_17058,N_14885,N_13290);
nand U17059 (N_17059,N_13319,N_14449);
nand U17060 (N_17060,N_14474,N_13733);
nand U17061 (N_17061,N_14785,N_13357);
nor U17062 (N_17062,N_14278,N_12588);
xor U17063 (N_17063,N_14185,N_13399);
and U17064 (N_17064,N_12666,N_12025);
nand U17065 (N_17065,N_13405,N_12333);
or U17066 (N_17066,N_14277,N_12298);
nor U17067 (N_17067,N_13832,N_12494);
nand U17068 (N_17068,N_13444,N_12623);
nand U17069 (N_17069,N_14420,N_12970);
nor U17070 (N_17070,N_14804,N_14342);
nor U17071 (N_17071,N_14586,N_12147);
and U17072 (N_17072,N_13346,N_14494);
or U17073 (N_17073,N_14252,N_12985);
or U17074 (N_17074,N_12038,N_13804);
xor U17075 (N_17075,N_12968,N_12120);
nand U17076 (N_17076,N_13002,N_13641);
nand U17077 (N_17077,N_13608,N_14401);
nor U17078 (N_17078,N_13805,N_14726);
nor U17079 (N_17079,N_12837,N_12984);
nand U17080 (N_17080,N_14225,N_13025);
nand U17081 (N_17081,N_13439,N_14767);
nor U17082 (N_17082,N_12318,N_13509);
and U17083 (N_17083,N_14334,N_13404);
and U17084 (N_17084,N_13889,N_14172);
xnor U17085 (N_17085,N_12030,N_13373);
xor U17086 (N_17086,N_13200,N_12956);
or U17087 (N_17087,N_13323,N_14200);
and U17088 (N_17088,N_13267,N_13695);
nand U17089 (N_17089,N_14236,N_13136);
nor U17090 (N_17090,N_13750,N_14792);
and U17091 (N_17091,N_13752,N_13765);
and U17092 (N_17092,N_14852,N_14582);
nand U17093 (N_17093,N_13986,N_13867);
and U17094 (N_17094,N_13585,N_12945);
xor U17095 (N_17095,N_13956,N_13709);
or U17096 (N_17096,N_14282,N_13709);
and U17097 (N_17097,N_13917,N_12046);
or U17098 (N_17098,N_12294,N_14172);
nor U17099 (N_17099,N_12055,N_12596);
nand U17100 (N_17100,N_13610,N_12695);
nand U17101 (N_17101,N_12802,N_12993);
nand U17102 (N_17102,N_12043,N_14833);
nand U17103 (N_17103,N_14593,N_14542);
xor U17104 (N_17104,N_12240,N_14166);
nor U17105 (N_17105,N_12976,N_13391);
nor U17106 (N_17106,N_14310,N_14260);
nand U17107 (N_17107,N_13954,N_12779);
nand U17108 (N_17108,N_13083,N_14581);
and U17109 (N_17109,N_14974,N_14663);
and U17110 (N_17110,N_12799,N_14039);
nand U17111 (N_17111,N_14924,N_13103);
nor U17112 (N_17112,N_13370,N_13742);
and U17113 (N_17113,N_13751,N_12531);
nor U17114 (N_17114,N_13183,N_13845);
nor U17115 (N_17115,N_14383,N_12452);
and U17116 (N_17116,N_12424,N_12553);
xnor U17117 (N_17117,N_14446,N_13919);
or U17118 (N_17118,N_14669,N_13237);
nor U17119 (N_17119,N_14926,N_12599);
or U17120 (N_17120,N_12339,N_14074);
or U17121 (N_17121,N_13387,N_13308);
or U17122 (N_17122,N_12485,N_12727);
xor U17123 (N_17123,N_13773,N_13681);
or U17124 (N_17124,N_14734,N_12686);
or U17125 (N_17125,N_12449,N_12633);
nand U17126 (N_17126,N_12028,N_13478);
and U17127 (N_17127,N_12770,N_12205);
nor U17128 (N_17128,N_12762,N_13163);
nor U17129 (N_17129,N_14979,N_12464);
nand U17130 (N_17130,N_12357,N_13595);
nand U17131 (N_17131,N_14900,N_12594);
xnor U17132 (N_17132,N_13128,N_13756);
or U17133 (N_17133,N_13355,N_12019);
or U17134 (N_17134,N_12157,N_13335);
and U17135 (N_17135,N_13409,N_12397);
and U17136 (N_17136,N_12462,N_14308);
nor U17137 (N_17137,N_12589,N_12309);
nand U17138 (N_17138,N_12101,N_12817);
or U17139 (N_17139,N_14180,N_14891);
and U17140 (N_17140,N_12511,N_12307);
nand U17141 (N_17141,N_12200,N_14817);
nor U17142 (N_17142,N_13600,N_12127);
nand U17143 (N_17143,N_14544,N_13925);
and U17144 (N_17144,N_14871,N_14683);
or U17145 (N_17145,N_12973,N_12350);
and U17146 (N_17146,N_14073,N_14884);
and U17147 (N_17147,N_14753,N_12656);
nand U17148 (N_17148,N_12559,N_13550);
or U17149 (N_17149,N_14170,N_12391);
or U17150 (N_17150,N_12734,N_13267);
nand U17151 (N_17151,N_12590,N_14142);
or U17152 (N_17152,N_14340,N_14569);
and U17153 (N_17153,N_12535,N_12835);
or U17154 (N_17154,N_12386,N_14289);
and U17155 (N_17155,N_12633,N_13484);
nand U17156 (N_17156,N_13785,N_14113);
xor U17157 (N_17157,N_13808,N_14474);
and U17158 (N_17158,N_14462,N_13975);
or U17159 (N_17159,N_13561,N_12207);
nor U17160 (N_17160,N_12443,N_13907);
or U17161 (N_17161,N_14012,N_13992);
nand U17162 (N_17162,N_14195,N_12972);
and U17163 (N_17163,N_12512,N_14133);
nor U17164 (N_17164,N_13843,N_14776);
and U17165 (N_17165,N_12240,N_13117);
xor U17166 (N_17166,N_12286,N_12751);
xor U17167 (N_17167,N_14917,N_12431);
nor U17168 (N_17168,N_13976,N_12862);
nor U17169 (N_17169,N_14757,N_13326);
or U17170 (N_17170,N_13193,N_14517);
nor U17171 (N_17171,N_13768,N_13602);
and U17172 (N_17172,N_14381,N_14142);
nand U17173 (N_17173,N_13135,N_13141);
xor U17174 (N_17174,N_12501,N_14610);
and U17175 (N_17175,N_14656,N_13494);
nor U17176 (N_17176,N_14004,N_14287);
nor U17177 (N_17177,N_14160,N_13209);
nand U17178 (N_17178,N_12201,N_14136);
nor U17179 (N_17179,N_13085,N_13785);
and U17180 (N_17180,N_13253,N_12419);
nand U17181 (N_17181,N_14828,N_12317);
and U17182 (N_17182,N_13579,N_12737);
or U17183 (N_17183,N_14274,N_12643);
and U17184 (N_17184,N_14484,N_12214);
or U17185 (N_17185,N_12186,N_12698);
xnor U17186 (N_17186,N_12589,N_12070);
and U17187 (N_17187,N_14614,N_13799);
and U17188 (N_17188,N_14397,N_12007);
or U17189 (N_17189,N_12490,N_12682);
or U17190 (N_17190,N_13939,N_13640);
nor U17191 (N_17191,N_12267,N_12043);
nand U17192 (N_17192,N_12601,N_13021);
xor U17193 (N_17193,N_12659,N_13625);
xnor U17194 (N_17194,N_13000,N_14224);
or U17195 (N_17195,N_13375,N_12519);
nand U17196 (N_17196,N_14450,N_14835);
xnor U17197 (N_17197,N_12582,N_14077);
and U17198 (N_17198,N_13234,N_13257);
xnor U17199 (N_17199,N_14579,N_13135);
nor U17200 (N_17200,N_13187,N_13894);
nand U17201 (N_17201,N_14278,N_14795);
xnor U17202 (N_17202,N_13345,N_13006);
and U17203 (N_17203,N_12538,N_14904);
and U17204 (N_17204,N_14944,N_14996);
nand U17205 (N_17205,N_13491,N_14748);
xnor U17206 (N_17206,N_13130,N_12443);
or U17207 (N_17207,N_12901,N_14642);
and U17208 (N_17208,N_13294,N_14934);
and U17209 (N_17209,N_12366,N_14858);
or U17210 (N_17210,N_13232,N_12874);
and U17211 (N_17211,N_12038,N_14380);
and U17212 (N_17212,N_13132,N_14972);
or U17213 (N_17213,N_13596,N_12295);
nand U17214 (N_17214,N_12479,N_13780);
nand U17215 (N_17215,N_12782,N_13777);
and U17216 (N_17216,N_12608,N_13647);
or U17217 (N_17217,N_12754,N_14990);
or U17218 (N_17218,N_12389,N_13855);
or U17219 (N_17219,N_14728,N_12905);
and U17220 (N_17220,N_12954,N_12951);
xnor U17221 (N_17221,N_12222,N_14413);
or U17222 (N_17222,N_14710,N_14688);
nand U17223 (N_17223,N_14377,N_13622);
nor U17224 (N_17224,N_12483,N_14824);
and U17225 (N_17225,N_14595,N_14623);
nor U17226 (N_17226,N_12909,N_14542);
nand U17227 (N_17227,N_13943,N_12165);
nand U17228 (N_17228,N_13150,N_14048);
or U17229 (N_17229,N_13282,N_12429);
xnor U17230 (N_17230,N_14148,N_14279);
nand U17231 (N_17231,N_13596,N_13225);
and U17232 (N_17232,N_13435,N_12075);
nor U17233 (N_17233,N_12523,N_13256);
and U17234 (N_17234,N_13380,N_13565);
or U17235 (N_17235,N_13479,N_13807);
and U17236 (N_17236,N_12898,N_12613);
xnor U17237 (N_17237,N_14243,N_12577);
nand U17238 (N_17238,N_13954,N_12947);
nand U17239 (N_17239,N_14148,N_14116);
xor U17240 (N_17240,N_14771,N_13517);
xor U17241 (N_17241,N_12567,N_12954);
or U17242 (N_17242,N_12321,N_12769);
and U17243 (N_17243,N_13983,N_12354);
or U17244 (N_17244,N_14724,N_14760);
xnor U17245 (N_17245,N_12096,N_13288);
xnor U17246 (N_17246,N_12529,N_12184);
xnor U17247 (N_17247,N_13887,N_12394);
and U17248 (N_17248,N_13732,N_14891);
and U17249 (N_17249,N_13563,N_13393);
xor U17250 (N_17250,N_12643,N_13248);
nand U17251 (N_17251,N_13363,N_13245);
or U17252 (N_17252,N_13072,N_12286);
or U17253 (N_17253,N_14221,N_14999);
and U17254 (N_17254,N_12318,N_12925);
xnor U17255 (N_17255,N_14842,N_14343);
nor U17256 (N_17256,N_12945,N_12931);
xor U17257 (N_17257,N_14095,N_14762);
or U17258 (N_17258,N_13106,N_13768);
nor U17259 (N_17259,N_13260,N_14278);
and U17260 (N_17260,N_14937,N_14238);
or U17261 (N_17261,N_12447,N_13872);
or U17262 (N_17262,N_13400,N_12449);
nand U17263 (N_17263,N_12825,N_14005);
xnor U17264 (N_17264,N_12249,N_12774);
or U17265 (N_17265,N_13347,N_12532);
nand U17266 (N_17266,N_12245,N_12388);
xnor U17267 (N_17267,N_13966,N_13773);
and U17268 (N_17268,N_14223,N_14909);
xnor U17269 (N_17269,N_14636,N_14213);
and U17270 (N_17270,N_12920,N_12554);
or U17271 (N_17271,N_12205,N_12140);
or U17272 (N_17272,N_12854,N_13814);
or U17273 (N_17273,N_13944,N_12234);
xnor U17274 (N_17274,N_12951,N_14131);
and U17275 (N_17275,N_14847,N_13857);
and U17276 (N_17276,N_14453,N_13128);
and U17277 (N_17277,N_12865,N_14938);
or U17278 (N_17278,N_12821,N_13575);
and U17279 (N_17279,N_14084,N_12309);
nor U17280 (N_17280,N_14953,N_12855);
or U17281 (N_17281,N_13918,N_12615);
and U17282 (N_17282,N_14022,N_13524);
xnor U17283 (N_17283,N_12489,N_13000);
xnor U17284 (N_17284,N_12174,N_12237);
or U17285 (N_17285,N_12776,N_13510);
and U17286 (N_17286,N_12775,N_13320);
xnor U17287 (N_17287,N_12667,N_13744);
nand U17288 (N_17288,N_13989,N_14709);
nor U17289 (N_17289,N_14729,N_13750);
and U17290 (N_17290,N_14940,N_12864);
or U17291 (N_17291,N_12437,N_13711);
xor U17292 (N_17292,N_14422,N_13261);
and U17293 (N_17293,N_14020,N_14896);
nor U17294 (N_17294,N_13569,N_12175);
nor U17295 (N_17295,N_12913,N_13725);
nand U17296 (N_17296,N_12548,N_13108);
nand U17297 (N_17297,N_12880,N_12457);
xnor U17298 (N_17298,N_12013,N_14491);
nor U17299 (N_17299,N_13299,N_13382);
nor U17300 (N_17300,N_13760,N_14532);
nand U17301 (N_17301,N_14301,N_14101);
nand U17302 (N_17302,N_14272,N_13647);
or U17303 (N_17303,N_12973,N_12849);
and U17304 (N_17304,N_14376,N_13530);
xnor U17305 (N_17305,N_13129,N_14890);
and U17306 (N_17306,N_13929,N_12339);
or U17307 (N_17307,N_13346,N_13957);
or U17308 (N_17308,N_13156,N_12786);
nor U17309 (N_17309,N_13783,N_13606);
nand U17310 (N_17310,N_14755,N_14667);
and U17311 (N_17311,N_13999,N_12818);
nor U17312 (N_17312,N_14252,N_12560);
or U17313 (N_17313,N_13850,N_14222);
or U17314 (N_17314,N_13414,N_13479);
and U17315 (N_17315,N_13384,N_12915);
and U17316 (N_17316,N_14610,N_12623);
and U17317 (N_17317,N_12028,N_13262);
xor U17318 (N_17318,N_14614,N_12587);
nand U17319 (N_17319,N_12851,N_14585);
nand U17320 (N_17320,N_14605,N_13909);
nor U17321 (N_17321,N_12866,N_12133);
xnor U17322 (N_17322,N_14008,N_14708);
or U17323 (N_17323,N_13449,N_12660);
or U17324 (N_17324,N_13923,N_12598);
and U17325 (N_17325,N_14909,N_12104);
and U17326 (N_17326,N_14045,N_13031);
xnor U17327 (N_17327,N_13242,N_14392);
xnor U17328 (N_17328,N_12942,N_14586);
xor U17329 (N_17329,N_13678,N_14932);
nor U17330 (N_17330,N_14467,N_13953);
or U17331 (N_17331,N_12080,N_12904);
or U17332 (N_17332,N_12672,N_14860);
nand U17333 (N_17333,N_13706,N_14302);
and U17334 (N_17334,N_13712,N_12854);
and U17335 (N_17335,N_13099,N_14936);
xor U17336 (N_17336,N_12919,N_14949);
nor U17337 (N_17337,N_13583,N_12850);
nor U17338 (N_17338,N_13391,N_12910);
or U17339 (N_17339,N_12470,N_12163);
and U17340 (N_17340,N_13823,N_14904);
or U17341 (N_17341,N_13647,N_13139);
and U17342 (N_17342,N_12780,N_14452);
nand U17343 (N_17343,N_12609,N_13182);
or U17344 (N_17344,N_12560,N_13661);
and U17345 (N_17345,N_12471,N_13636);
and U17346 (N_17346,N_14384,N_12939);
nor U17347 (N_17347,N_12941,N_14526);
nor U17348 (N_17348,N_13421,N_13664);
and U17349 (N_17349,N_13443,N_12358);
and U17350 (N_17350,N_12610,N_14134);
xnor U17351 (N_17351,N_13013,N_12935);
nand U17352 (N_17352,N_12955,N_12673);
nor U17353 (N_17353,N_13712,N_14178);
xnor U17354 (N_17354,N_14603,N_13374);
and U17355 (N_17355,N_14081,N_12409);
and U17356 (N_17356,N_14665,N_14031);
nor U17357 (N_17357,N_12923,N_13751);
and U17358 (N_17358,N_12863,N_14601);
xor U17359 (N_17359,N_14190,N_13706);
xnor U17360 (N_17360,N_13292,N_12849);
nand U17361 (N_17361,N_12823,N_14542);
nor U17362 (N_17362,N_13020,N_13305);
xor U17363 (N_17363,N_14869,N_12780);
and U17364 (N_17364,N_14572,N_14104);
nand U17365 (N_17365,N_12081,N_13517);
and U17366 (N_17366,N_14162,N_12437);
and U17367 (N_17367,N_12653,N_13819);
and U17368 (N_17368,N_13731,N_12678);
xnor U17369 (N_17369,N_12662,N_12095);
or U17370 (N_17370,N_13456,N_13036);
or U17371 (N_17371,N_13417,N_14190);
or U17372 (N_17372,N_13880,N_14243);
xnor U17373 (N_17373,N_13221,N_14962);
xnor U17374 (N_17374,N_13073,N_14287);
and U17375 (N_17375,N_14949,N_14872);
nor U17376 (N_17376,N_12991,N_13809);
or U17377 (N_17377,N_14589,N_14069);
or U17378 (N_17378,N_14383,N_13916);
nand U17379 (N_17379,N_14787,N_14170);
nor U17380 (N_17380,N_12426,N_13600);
xor U17381 (N_17381,N_13704,N_14228);
or U17382 (N_17382,N_13417,N_12874);
xnor U17383 (N_17383,N_12374,N_12262);
nand U17384 (N_17384,N_13071,N_14804);
and U17385 (N_17385,N_14219,N_13016);
or U17386 (N_17386,N_14427,N_12800);
and U17387 (N_17387,N_12606,N_12613);
and U17388 (N_17388,N_14001,N_12641);
xor U17389 (N_17389,N_12094,N_14592);
xnor U17390 (N_17390,N_14473,N_12056);
or U17391 (N_17391,N_12960,N_12530);
nand U17392 (N_17392,N_14514,N_14919);
or U17393 (N_17393,N_12675,N_12133);
and U17394 (N_17394,N_13477,N_12232);
nor U17395 (N_17395,N_12278,N_12275);
nand U17396 (N_17396,N_14156,N_13267);
xnor U17397 (N_17397,N_14110,N_14546);
and U17398 (N_17398,N_14392,N_13889);
nor U17399 (N_17399,N_12845,N_14459);
and U17400 (N_17400,N_13683,N_13263);
nand U17401 (N_17401,N_14685,N_14285);
xnor U17402 (N_17402,N_12583,N_14309);
xor U17403 (N_17403,N_14638,N_13339);
or U17404 (N_17404,N_14201,N_13732);
nand U17405 (N_17405,N_13875,N_14215);
nor U17406 (N_17406,N_12527,N_12240);
and U17407 (N_17407,N_12390,N_12248);
nor U17408 (N_17408,N_12637,N_12194);
nor U17409 (N_17409,N_13911,N_14881);
nor U17410 (N_17410,N_14674,N_14647);
xor U17411 (N_17411,N_12779,N_14806);
and U17412 (N_17412,N_13141,N_14396);
nand U17413 (N_17413,N_14098,N_13032);
nand U17414 (N_17414,N_13479,N_12666);
xnor U17415 (N_17415,N_13427,N_14169);
nand U17416 (N_17416,N_13280,N_14269);
and U17417 (N_17417,N_13620,N_13305);
xnor U17418 (N_17418,N_12821,N_12795);
and U17419 (N_17419,N_13080,N_14683);
nand U17420 (N_17420,N_13228,N_14107);
xor U17421 (N_17421,N_12883,N_13838);
or U17422 (N_17422,N_12602,N_14729);
or U17423 (N_17423,N_12930,N_12209);
nor U17424 (N_17424,N_14363,N_12233);
nand U17425 (N_17425,N_13397,N_13253);
or U17426 (N_17426,N_14065,N_13685);
nand U17427 (N_17427,N_14623,N_13533);
nand U17428 (N_17428,N_13899,N_13432);
xor U17429 (N_17429,N_14789,N_14650);
or U17430 (N_17430,N_14137,N_12543);
or U17431 (N_17431,N_13453,N_13335);
nand U17432 (N_17432,N_13162,N_12513);
and U17433 (N_17433,N_12756,N_13060);
nand U17434 (N_17434,N_13513,N_14253);
nor U17435 (N_17435,N_12376,N_13222);
xor U17436 (N_17436,N_14722,N_13762);
xnor U17437 (N_17437,N_13656,N_14039);
xnor U17438 (N_17438,N_13277,N_14829);
and U17439 (N_17439,N_12919,N_13337);
and U17440 (N_17440,N_14538,N_13204);
and U17441 (N_17441,N_12091,N_12119);
and U17442 (N_17442,N_14740,N_13426);
xor U17443 (N_17443,N_13589,N_13848);
nand U17444 (N_17444,N_12621,N_13980);
nor U17445 (N_17445,N_13000,N_13025);
nor U17446 (N_17446,N_13326,N_12798);
nand U17447 (N_17447,N_14337,N_14588);
nor U17448 (N_17448,N_14621,N_13548);
or U17449 (N_17449,N_12639,N_13595);
nand U17450 (N_17450,N_13736,N_13882);
or U17451 (N_17451,N_13956,N_13186);
and U17452 (N_17452,N_12203,N_14810);
nand U17453 (N_17453,N_14854,N_13418);
nand U17454 (N_17454,N_14703,N_13264);
nor U17455 (N_17455,N_13314,N_12893);
xor U17456 (N_17456,N_13796,N_14541);
xnor U17457 (N_17457,N_12071,N_12684);
xor U17458 (N_17458,N_13426,N_12990);
xnor U17459 (N_17459,N_14923,N_14399);
xnor U17460 (N_17460,N_14591,N_14103);
xor U17461 (N_17461,N_13205,N_12400);
xnor U17462 (N_17462,N_13107,N_13579);
or U17463 (N_17463,N_13778,N_14692);
or U17464 (N_17464,N_13627,N_13322);
or U17465 (N_17465,N_13966,N_13816);
nor U17466 (N_17466,N_14124,N_14924);
and U17467 (N_17467,N_13434,N_13415);
xor U17468 (N_17468,N_14029,N_14358);
and U17469 (N_17469,N_14334,N_14677);
or U17470 (N_17470,N_14390,N_14455);
or U17471 (N_17471,N_12109,N_13531);
xnor U17472 (N_17472,N_13976,N_12026);
nand U17473 (N_17473,N_12475,N_12357);
and U17474 (N_17474,N_13791,N_13451);
and U17475 (N_17475,N_12374,N_13644);
xor U17476 (N_17476,N_12317,N_14427);
xor U17477 (N_17477,N_14001,N_12934);
nor U17478 (N_17478,N_13427,N_12330);
nor U17479 (N_17479,N_14641,N_14100);
nand U17480 (N_17480,N_14529,N_14324);
nor U17481 (N_17481,N_12966,N_12546);
or U17482 (N_17482,N_14055,N_13784);
and U17483 (N_17483,N_12552,N_14542);
nand U17484 (N_17484,N_12254,N_13587);
xor U17485 (N_17485,N_13603,N_13474);
and U17486 (N_17486,N_13154,N_14300);
xor U17487 (N_17487,N_12504,N_12941);
xor U17488 (N_17488,N_12508,N_13639);
nand U17489 (N_17489,N_14072,N_13675);
and U17490 (N_17490,N_12905,N_14883);
nand U17491 (N_17491,N_12556,N_14335);
nor U17492 (N_17492,N_12781,N_12241);
xnor U17493 (N_17493,N_12038,N_13677);
xnor U17494 (N_17494,N_14233,N_12197);
nor U17495 (N_17495,N_12472,N_12535);
or U17496 (N_17496,N_13493,N_12581);
nor U17497 (N_17497,N_14380,N_13034);
xor U17498 (N_17498,N_14598,N_14505);
nor U17499 (N_17499,N_14805,N_12979);
and U17500 (N_17500,N_13119,N_14369);
or U17501 (N_17501,N_14453,N_12782);
nand U17502 (N_17502,N_12439,N_12681);
nor U17503 (N_17503,N_14547,N_12833);
nor U17504 (N_17504,N_14908,N_12746);
or U17505 (N_17505,N_12860,N_13240);
nor U17506 (N_17506,N_12156,N_13907);
nand U17507 (N_17507,N_12236,N_12885);
nor U17508 (N_17508,N_14527,N_13321);
xor U17509 (N_17509,N_12304,N_13169);
and U17510 (N_17510,N_13825,N_12848);
xor U17511 (N_17511,N_12044,N_14733);
or U17512 (N_17512,N_13427,N_12520);
nor U17513 (N_17513,N_12070,N_14702);
xor U17514 (N_17514,N_13070,N_12304);
nor U17515 (N_17515,N_13969,N_12688);
xnor U17516 (N_17516,N_14366,N_13446);
or U17517 (N_17517,N_13526,N_13712);
xor U17518 (N_17518,N_13930,N_13615);
and U17519 (N_17519,N_13688,N_12916);
or U17520 (N_17520,N_14268,N_14055);
nand U17521 (N_17521,N_12464,N_12840);
xor U17522 (N_17522,N_12984,N_14936);
or U17523 (N_17523,N_14150,N_13426);
nor U17524 (N_17524,N_12030,N_12696);
xnor U17525 (N_17525,N_13860,N_13119);
nand U17526 (N_17526,N_12176,N_14693);
xor U17527 (N_17527,N_14647,N_13278);
nand U17528 (N_17528,N_13787,N_13328);
nor U17529 (N_17529,N_14188,N_14671);
nor U17530 (N_17530,N_13060,N_13554);
nand U17531 (N_17531,N_14409,N_12235);
nand U17532 (N_17532,N_13668,N_14647);
nand U17533 (N_17533,N_14123,N_13182);
nor U17534 (N_17534,N_13262,N_14011);
and U17535 (N_17535,N_12889,N_14194);
xnor U17536 (N_17536,N_14288,N_14426);
xnor U17537 (N_17537,N_12861,N_12484);
nor U17538 (N_17538,N_14864,N_14656);
nand U17539 (N_17539,N_14194,N_12839);
xnor U17540 (N_17540,N_13591,N_12536);
or U17541 (N_17541,N_13696,N_12006);
nand U17542 (N_17542,N_13079,N_12387);
nor U17543 (N_17543,N_13908,N_13540);
or U17544 (N_17544,N_14158,N_12401);
and U17545 (N_17545,N_14570,N_13390);
xnor U17546 (N_17546,N_14638,N_14368);
nand U17547 (N_17547,N_12392,N_14164);
and U17548 (N_17548,N_13952,N_13996);
and U17549 (N_17549,N_12048,N_13036);
nand U17550 (N_17550,N_12413,N_13772);
nor U17551 (N_17551,N_14609,N_12458);
and U17552 (N_17552,N_12441,N_13396);
xor U17553 (N_17553,N_13174,N_13265);
xnor U17554 (N_17554,N_13201,N_13975);
xnor U17555 (N_17555,N_14245,N_12592);
or U17556 (N_17556,N_14509,N_13307);
nor U17557 (N_17557,N_13100,N_14833);
nor U17558 (N_17558,N_13253,N_12661);
nor U17559 (N_17559,N_12310,N_13166);
nand U17560 (N_17560,N_13960,N_13822);
nor U17561 (N_17561,N_13381,N_13739);
or U17562 (N_17562,N_13852,N_13901);
nor U17563 (N_17563,N_12377,N_12620);
nand U17564 (N_17564,N_14707,N_12112);
nand U17565 (N_17565,N_13088,N_12992);
nor U17566 (N_17566,N_13052,N_12534);
nor U17567 (N_17567,N_14447,N_13100);
xor U17568 (N_17568,N_14479,N_14825);
nand U17569 (N_17569,N_14082,N_13902);
or U17570 (N_17570,N_13139,N_12080);
nor U17571 (N_17571,N_14062,N_12216);
or U17572 (N_17572,N_14761,N_12107);
nor U17573 (N_17573,N_12894,N_14248);
or U17574 (N_17574,N_14008,N_14019);
or U17575 (N_17575,N_14767,N_14437);
and U17576 (N_17576,N_12447,N_13361);
and U17577 (N_17577,N_13117,N_14731);
nand U17578 (N_17578,N_13234,N_14599);
nand U17579 (N_17579,N_12425,N_13049);
nand U17580 (N_17580,N_13904,N_14168);
nand U17581 (N_17581,N_12470,N_13789);
nand U17582 (N_17582,N_13569,N_12689);
nor U17583 (N_17583,N_14078,N_12807);
xor U17584 (N_17584,N_14849,N_12265);
or U17585 (N_17585,N_14097,N_14166);
and U17586 (N_17586,N_14234,N_13919);
nand U17587 (N_17587,N_12743,N_14595);
and U17588 (N_17588,N_14396,N_13594);
or U17589 (N_17589,N_12647,N_13221);
or U17590 (N_17590,N_14463,N_13646);
nor U17591 (N_17591,N_14557,N_14157);
or U17592 (N_17592,N_14575,N_14716);
or U17593 (N_17593,N_12508,N_12491);
nand U17594 (N_17594,N_12760,N_13870);
or U17595 (N_17595,N_12141,N_14038);
nor U17596 (N_17596,N_14614,N_13884);
and U17597 (N_17597,N_13149,N_13115);
and U17598 (N_17598,N_12871,N_12200);
and U17599 (N_17599,N_14378,N_13081);
nand U17600 (N_17600,N_12989,N_14004);
or U17601 (N_17601,N_12958,N_12353);
xnor U17602 (N_17602,N_13515,N_14604);
nor U17603 (N_17603,N_14896,N_12027);
or U17604 (N_17604,N_12672,N_13770);
xnor U17605 (N_17605,N_13382,N_14177);
or U17606 (N_17606,N_14610,N_12091);
nor U17607 (N_17607,N_14928,N_13500);
xnor U17608 (N_17608,N_14764,N_12877);
or U17609 (N_17609,N_13824,N_13762);
nand U17610 (N_17610,N_13432,N_14274);
xnor U17611 (N_17611,N_13701,N_12895);
xnor U17612 (N_17612,N_12650,N_14363);
or U17613 (N_17613,N_14323,N_14178);
xnor U17614 (N_17614,N_14777,N_12050);
or U17615 (N_17615,N_14375,N_13366);
xnor U17616 (N_17616,N_12461,N_14014);
nand U17617 (N_17617,N_12880,N_12592);
and U17618 (N_17618,N_12745,N_12803);
nand U17619 (N_17619,N_12399,N_12969);
and U17620 (N_17620,N_14780,N_13260);
and U17621 (N_17621,N_12990,N_14699);
xor U17622 (N_17622,N_12712,N_14570);
and U17623 (N_17623,N_12762,N_13607);
nor U17624 (N_17624,N_12562,N_12818);
or U17625 (N_17625,N_13443,N_12977);
xnor U17626 (N_17626,N_12859,N_13910);
nand U17627 (N_17627,N_13898,N_13033);
or U17628 (N_17628,N_12626,N_12579);
and U17629 (N_17629,N_13159,N_13621);
nor U17630 (N_17630,N_14736,N_14129);
or U17631 (N_17631,N_13560,N_14242);
and U17632 (N_17632,N_12647,N_12787);
nor U17633 (N_17633,N_13006,N_14493);
nor U17634 (N_17634,N_13579,N_14589);
xor U17635 (N_17635,N_12812,N_12559);
or U17636 (N_17636,N_13406,N_12150);
and U17637 (N_17637,N_14080,N_13235);
nand U17638 (N_17638,N_13759,N_12556);
xnor U17639 (N_17639,N_14796,N_14320);
or U17640 (N_17640,N_14361,N_13001);
xnor U17641 (N_17641,N_14262,N_14687);
nand U17642 (N_17642,N_14480,N_14777);
xnor U17643 (N_17643,N_13929,N_12516);
and U17644 (N_17644,N_13760,N_13835);
or U17645 (N_17645,N_13379,N_12762);
and U17646 (N_17646,N_13246,N_13269);
xnor U17647 (N_17647,N_14933,N_14478);
or U17648 (N_17648,N_13290,N_14924);
nor U17649 (N_17649,N_14430,N_13149);
and U17650 (N_17650,N_14827,N_12193);
nand U17651 (N_17651,N_12762,N_12804);
xor U17652 (N_17652,N_12960,N_13509);
nand U17653 (N_17653,N_13248,N_13678);
xnor U17654 (N_17654,N_13860,N_12428);
xnor U17655 (N_17655,N_13983,N_14726);
nor U17656 (N_17656,N_13596,N_12804);
or U17657 (N_17657,N_12369,N_12042);
xnor U17658 (N_17658,N_13648,N_13957);
xnor U17659 (N_17659,N_14443,N_13741);
xnor U17660 (N_17660,N_12890,N_14457);
or U17661 (N_17661,N_12962,N_12716);
xor U17662 (N_17662,N_13668,N_14076);
nor U17663 (N_17663,N_14025,N_14068);
nand U17664 (N_17664,N_12309,N_14797);
and U17665 (N_17665,N_14501,N_14398);
and U17666 (N_17666,N_13134,N_13297);
xor U17667 (N_17667,N_13272,N_13548);
nor U17668 (N_17668,N_14390,N_12940);
or U17669 (N_17669,N_13761,N_13915);
xor U17670 (N_17670,N_14879,N_14525);
and U17671 (N_17671,N_14191,N_12230);
or U17672 (N_17672,N_12035,N_13435);
or U17673 (N_17673,N_12523,N_12898);
nand U17674 (N_17674,N_13361,N_13592);
nor U17675 (N_17675,N_14870,N_12936);
and U17676 (N_17676,N_12859,N_14258);
nand U17677 (N_17677,N_14693,N_12158);
nand U17678 (N_17678,N_13477,N_13223);
nor U17679 (N_17679,N_14289,N_12983);
xnor U17680 (N_17680,N_13902,N_14306);
or U17681 (N_17681,N_13394,N_13381);
nand U17682 (N_17682,N_14216,N_13584);
and U17683 (N_17683,N_12426,N_12321);
nand U17684 (N_17684,N_14501,N_14172);
nor U17685 (N_17685,N_14946,N_14012);
xnor U17686 (N_17686,N_12124,N_13421);
or U17687 (N_17687,N_14766,N_14414);
or U17688 (N_17688,N_13713,N_12838);
nand U17689 (N_17689,N_13538,N_12472);
or U17690 (N_17690,N_12128,N_12405);
or U17691 (N_17691,N_14412,N_12161);
nand U17692 (N_17692,N_13237,N_13703);
xor U17693 (N_17693,N_13985,N_13595);
nand U17694 (N_17694,N_14584,N_14928);
xnor U17695 (N_17695,N_12160,N_13541);
and U17696 (N_17696,N_14412,N_12329);
or U17697 (N_17697,N_13665,N_14866);
nor U17698 (N_17698,N_14311,N_13855);
or U17699 (N_17699,N_14765,N_14729);
nor U17700 (N_17700,N_12152,N_13134);
nor U17701 (N_17701,N_14168,N_12478);
and U17702 (N_17702,N_14360,N_13106);
nand U17703 (N_17703,N_14829,N_14807);
xnor U17704 (N_17704,N_14351,N_12709);
or U17705 (N_17705,N_14464,N_13001);
or U17706 (N_17706,N_12402,N_12708);
or U17707 (N_17707,N_12417,N_13104);
or U17708 (N_17708,N_12498,N_14495);
or U17709 (N_17709,N_12754,N_12083);
nor U17710 (N_17710,N_13484,N_13429);
or U17711 (N_17711,N_14800,N_13609);
xnor U17712 (N_17712,N_12093,N_13030);
nand U17713 (N_17713,N_14655,N_13247);
or U17714 (N_17714,N_12936,N_14577);
and U17715 (N_17715,N_13698,N_14790);
nand U17716 (N_17716,N_14657,N_12230);
xnor U17717 (N_17717,N_13579,N_12452);
xnor U17718 (N_17718,N_14911,N_12202);
xnor U17719 (N_17719,N_13990,N_14192);
and U17720 (N_17720,N_14519,N_12922);
xnor U17721 (N_17721,N_12663,N_12738);
and U17722 (N_17722,N_14151,N_13990);
xor U17723 (N_17723,N_14787,N_12201);
nor U17724 (N_17724,N_12739,N_12362);
nor U17725 (N_17725,N_13814,N_12390);
or U17726 (N_17726,N_12015,N_12849);
nor U17727 (N_17727,N_14020,N_13855);
nor U17728 (N_17728,N_14261,N_13510);
xor U17729 (N_17729,N_12536,N_14283);
and U17730 (N_17730,N_14186,N_12871);
nor U17731 (N_17731,N_14760,N_12890);
and U17732 (N_17732,N_14721,N_14582);
xor U17733 (N_17733,N_14706,N_14459);
and U17734 (N_17734,N_12647,N_12084);
and U17735 (N_17735,N_12038,N_13415);
and U17736 (N_17736,N_13726,N_12312);
or U17737 (N_17737,N_14686,N_12607);
and U17738 (N_17738,N_12712,N_12430);
xor U17739 (N_17739,N_12019,N_13774);
or U17740 (N_17740,N_13858,N_13291);
nor U17741 (N_17741,N_13116,N_14522);
xnor U17742 (N_17742,N_12194,N_14321);
or U17743 (N_17743,N_14330,N_12107);
or U17744 (N_17744,N_13270,N_14627);
xor U17745 (N_17745,N_13161,N_12884);
or U17746 (N_17746,N_14501,N_13075);
xnor U17747 (N_17747,N_13395,N_14607);
nor U17748 (N_17748,N_14543,N_14361);
and U17749 (N_17749,N_14700,N_13619);
xnor U17750 (N_17750,N_14990,N_14965);
and U17751 (N_17751,N_14064,N_14712);
xnor U17752 (N_17752,N_12727,N_13928);
nand U17753 (N_17753,N_12643,N_13245);
and U17754 (N_17754,N_12830,N_14620);
xor U17755 (N_17755,N_12148,N_14157);
or U17756 (N_17756,N_12282,N_12197);
xor U17757 (N_17757,N_14206,N_13477);
nor U17758 (N_17758,N_12525,N_13417);
nand U17759 (N_17759,N_12301,N_13967);
nor U17760 (N_17760,N_14318,N_13262);
xnor U17761 (N_17761,N_12358,N_12496);
xor U17762 (N_17762,N_13200,N_13733);
and U17763 (N_17763,N_14435,N_13107);
xnor U17764 (N_17764,N_13900,N_14979);
nor U17765 (N_17765,N_12764,N_14611);
nor U17766 (N_17766,N_13876,N_12940);
xnor U17767 (N_17767,N_12316,N_14034);
and U17768 (N_17768,N_14889,N_12405);
nand U17769 (N_17769,N_12512,N_13499);
or U17770 (N_17770,N_13304,N_13418);
xnor U17771 (N_17771,N_12780,N_12697);
xor U17772 (N_17772,N_13142,N_14278);
or U17773 (N_17773,N_12039,N_13955);
or U17774 (N_17774,N_13785,N_14508);
xor U17775 (N_17775,N_14933,N_14222);
and U17776 (N_17776,N_14315,N_14422);
and U17777 (N_17777,N_12126,N_14614);
and U17778 (N_17778,N_14509,N_12128);
nor U17779 (N_17779,N_13857,N_13961);
nor U17780 (N_17780,N_12240,N_12836);
nor U17781 (N_17781,N_12401,N_12755);
xor U17782 (N_17782,N_14095,N_12754);
and U17783 (N_17783,N_14303,N_14180);
nor U17784 (N_17784,N_12139,N_14425);
nand U17785 (N_17785,N_14797,N_14306);
or U17786 (N_17786,N_14828,N_13963);
or U17787 (N_17787,N_12716,N_13229);
or U17788 (N_17788,N_13966,N_13436);
xor U17789 (N_17789,N_14585,N_13361);
or U17790 (N_17790,N_13456,N_13723);
and U17791 (N_17791,N_13085,N_14968);
nor U17792 (N_17792,N_13060,N_12392);
or U17793 (N_17793,N_14030,N_12557);
nand U17794 (N_17794,N_14492,N_12860);
and U17795 (N_17795,N_13107,N_12865);
or U17796 (N_17796,N_13804,N_14111);
xnor U17797 (N_17797,N_13597,N_12501);
xnor U17798 (N_17798,N_13883,N_14792);
nor U17799 (N_17799,N_13552,N_14221);
nand U17800 (N_17800,N_14740,N_14833);
or U17801 (N_17801,N_13343,N_14605);
nor U17802 (N_17802,N_14186,N_13536);
nand U17803 (N_17803,N_13431,N_14228);
xor U17804 (N_17804,N_14925,N_12749);
and U17805 (N_17805,N_14757,N_13296);
and U17806 (N_17806,N_14769,N_12408);
or U17807 (N_17807,N_14066,N_14269);
or U17808 (N_17808,N_12148,N_14954);
nor U17809 (N_17809,N_13154,N_14898);
xnor U17810 (N_17810,N_12991,N_12333);
xor U17811 (N_17811,N_14857,N_12142);
nor U17812 (N_17812,N_14567,N_13884);
nor U17813 (N_17813,N_14023,N_14898);
nand U17814 (N_17814,N_13272,N_12698);
xor U17815 (N_17815,N_12008,N_13976);
nand U17816 (N_17816,N_13941,N_13049);
xnor U17817 (N_17817,N_14922,N_13932);
nand U17818 (N_17818,N_14106,N_12359);
or U17819 (N_17819,N_13795,N_12690);
nand U17820 (N_17820,N_13546,N_13347);
xnor U17821 (N_17821,N_12114,N_12806);
nand U17822 (N_17822,N_12156,N_12707);
and U17823 (N_17823,N_13226,N_13508);
or U17824 (N_17824,N_12161,N_14346);
nor U17825 (N_17825,N_12267,N_14744);
or U17826 (N_17826,N_12986,N_12025);
xnor U17827 (N_17827,N_14154,N_14212);
nand U17828 (N_17828,N_13103,N_14223);
xor U17829 (N_17829,N_14537,N_12378);
xor U17830 (N_17830,N_14677,N_13523);
and U17831 (N_17831,N_14504,N_14342);
or U17832 (N_17832,N_12422,N_12538);
nor U17833 (N_17833,N_13503,N_14381);
and U17834 (N_17834,N_13970,N_12117);
xnor U17835 (N_17835,N_14152,N_13230);
xor U17836 (N_17836,N_14191,N_13203);
and U17837 (N_17837,N_14140,N_14110);
or U17838 (N_17838,N_14790,N_13981);
and U17839 (N_17839,N_14092,N_14278);
nor U17840 (N_17840,N_13548,N_14622);
and U17841 (N_17841,N_12911,N_13904);
and U17842 (N_17842,N_14341,N_13440);
or U17843 (N_17843,N_14175,N_12492);
nor U17844 (N_17844,N_14669,N_13419);
and U17845 (N_17845,N_13365,N_12548);
or U17846 (N_17846,N_12521,N_12025);
nor U17847 (N_17847,N_12471,N_14916);
xnor U17848 (N_17848,N_12962,N_14997);
nor U17849 (N_17849,N_12068,N_12797);
nand U17850 (N_17850,N_12501,N_12104);
nor U17851 (N_17851,N_13254,N_14209);
nor U17852 (N_17852,N_13630,N_14179);
nand U17853 (N_17853,N_12486,N_14567);
and U17854 (N_17854,N_13820,N_13342);
or U17855 (N_17855,N_12250,N_12107);
or U17856 (N_17856,N_14614,N_12517);
nor U17857 (N_17857,N_14005,N_14066);
and U17858 (N_17858,N_12302,N_13015);
xnor U17859 (N_17859,N_14566,N_12104);
nand U17860 (N_17860,N_14478,N_13981);
nand U17861 (N_17861,N_14624,N_14156);
or U17862 (N_17862,N_14974,N_14369);
nor U17863 (N_17863,N_13261,N_12897);
nor U17864 (N_17864,N_14971,N_13992);
nor U17865 (N_17865,N_14068,N_13141);
nand U17866 (N_17866,N_14079,N_13778);
xor U17867 (N_17867,N_12357,N_14975);
or U17868 (N_17868,N_14526,N_13707);
and U17869 (N_17869,N_12735,N_13660);
xnor U17870 (N_17870,N_14046,N_13721);
xnor U17871 (N_17871,N_14407,N_12651);
nor U17872 (N_17872,N_13755,N_14068);
xnor U17873 (N_17873,N_12662,N_13683);
and U17874 (N_17874,N_14665,N_14963);
xor U17875 (N_17875,N_14686,N_13324);
nand U17876 (N_17876,N_12679,N_13522);
and U17877 (N_17877,N_13345,N_13172);
and U17878 (N_17878,N_14716,N_14374);
or U17879 (N_17879,N_13517,N_12837);
xnor U17880 (N_17880,N_14928,N_14653);
nor U17881 (N_17881,N_13106,N_13581);
nor U17882 (N_17882,N_13215,N_12001);
nor U17883 (N_17883,N_12772,N_14275);
or U17884 (N_17884,N_14844,N_14759);
and U17885 (N_17885,N_12550,N_14318);
or U17886 (N_17886,N_14644,N_13590);
or U17887 (N_17887,N_13453,N_14531);
nand U17888 (N_17888,N_13920,N_12244);
nand U17889 (N_17889,N_12501,N_13882);
and U17890 (N_17890,N_13578,N_14119);
or U17891 (N_17891,N_12793,N_14155);
xor U17892 (N_17892,N_14284,N_12454);
nor U17893 (N_17893,N_14587,N_13033);
xnor U17894 (N_17894,N_12179,N_13655);
and U17895 (N_17895,N_13345,N_12089);
xor U17896 (N_17896,N_14543,N_14971);
and U17897 (N_17897,N_12672,N_14616);
or U17898 (N_17898,N_14090,N_12245);
xnor U17899 (N_17899,N_14006,N_13783);
or U17900 (N_17900,N_14693,N_13393);
or U17901 (N_17901,N_14923,N_12789);
or U17902 (N_17902,N_14902,N_13448);
xor U17903 (N_17903,N_12274,N_12542);
nor U17904 (N_17904,N_12160,N_14863);
and U17905 (N_17905,N_13453,N_13862);
or U17906 (N_17906,N_12877,N_14970);
and U17907 (N_17907,N_12883,N_14947);
and U17908 (N_17908,N_13848,N_13698);
nor U17909 (N_17909,N_14796,N_12160);
nor U17910 (N_17910,N_13559,N_13273);
and U17911 (N_17911,N_13792,N_13179);
xnor U17912 (N_17912,N_12847,N_14250);
nand U17913 (N_17913,N_12632,N_13918);
nand U17914 (N_17914,N_14463,N_13729);
nand U17915 (N_17915,N_12935,N_12068);
and U17916 (N_17916,N_14764,N_13493);
nand U17917 (N_17917,N_14236,N_13452);
xnor U17918 (N_17918,N_14945,N_12469);
xnor U17919 (N_17919,N_14854,N_12202);
nor U17920 (N_17920,N_14518,N_12500);
or U17921 (N_17921,N_12064,N_13934);
xnor U17922 (N_17922,N_13268,N_13212);
nand U17923 (N_17923,N_12755,N_12676);
or U17924 (N_17924,N_14223,N_13543);
nor U17925 (N_17925,N_12623,N_14704);
nand U17926 (N_17926,N_14821,N_13228);
and U17927 (N_17927,N_14186,N_12219);
nor U17928 (N_17928,N_13807,N_12834);
and U17929 (N_17929,N_14513,N_13614);
or U17930 (N_17930,N_12257,N_14794);
xor U17931 (N_17931,N_14037,N_14326);
xnor U17932 (N_17932,N_12841,N_13892);
nor U17933 (N_17933,N_12048,N_14463);
nor U17934 (N_17934,N_12822,N_12710);
nor U17935 (N_17935,N_13841,N_13883);
xnor U17936 (N_17936,N_13435,N_12703);
xnor U17937 (N_17937,N_14118,N_13923);
nor U17938 (N_17938,N_13984,N_12988);
xor U17939 (N_17939,N_12483,N_12812);
nor U17940 (N_17940,N_14466,N_14500);
nand U17941 (N_17941,N_14251,N_14435);
and U17942 (N_17942,N_13652,N_14059);
nor U17943 (N_17943,N_13126,N_14521);
nor U17944 (N_17944,N_13110,N_14914);
or U17945 (N_17945,N_12555,N_12876);
xnor U17946 (N_17946,N_14262,N_12180);
and U17947 (N_17947,N_14381,N_13098);
or U17948 (N_17948,N_14521,N_14741);
and U17949 (N_17949,N_12144,N_13391);
xnor U17950 (N_17950,N_14167,N_14462);
xor U17951 (N_17951,N_13760,N_12913);
or U17952 (N_17952,N_12955,N_12622);
xor U17953 (N_17953,N_14276,N_13642);
xor U17954 (N_17954,N_14454,N_14733);
nand U17955 (N_17955,N_12913,N_12845);
and U17956 (N_17956,N_14362,N_12423);
or U17957 (N_17957,N_13099,N_13851);
or U17958 (N_17958,N_14542,N_14732);
nor U17959 (N_17959,N_12082,N_12288);
nand U17960 (N_17960,N_13866,N_14180);
or U17961 (N_17961,N_14630,N_14224);
xnor U17962 (N_17962,N_14741,N_14791);
xor U17963 (N_17963,N_14735,N_13882);
or U17964 (N_17964,N_13371,N_12269);
or U17965 (N_17965,N_14461,N_14530);
or U17966 (N_17966,N_14574,N_14329);
nand U17967 (N_17967,N_12713,N_12711);
and U17968 (N_17968,N_12851,N_12124);
or U17969 (N_17969,N_14452,N_13541);
and U17970 (N_17970,N_14324,N_14185);
or U17971 (N_17971,N_13674,N_13463);
and U17972 (N_17972,N_14877,N_14824);
or U17973 (N_17973,N_13491,N_14832);
nor U17974 (N_17974,N_12675,N_14495);
nor U17975 (N_17975,N_14103,N_12087);
or U17976 (N_17976,N_13783,N_14485);
xnor U17977 (N_17977,N_14118,N_12152);
xnor U17978 (N_17978,N_12458,N_14232);
xnor U17979 (N_17979,N_12999,N_12459);
nor U17980 (N_17980,N_12061,N_12501);
or U17981 (N_17981,N_14320,N_13196);
or U17982 (N_17982,N_13736,N_13557);
and U17983 (N_17983,N_14133,N_13072);
and U17984 (N_17984,N_14063,N_13432);
and U17985 (N_17985,N_13103,N_13973);
or U17986 (N_17986,N_14979,N_14371);
nand U17987 (N_17987,N_13194,N_12858);
or U17988 (N_17988,N_13032,N_12805);
or U17989 (N_17989,N_13666,N_14414);
and U17990 (N_17990,N_13445,N_13954);
and U17991 (N_17991,N_12398,N_12007);
and U17992 (N_17992,N_12624,N_13492);
and U17993 (N_17993,N_12925,N_13568);
or U17994 (N_17994,N_13225,N_12896);
nand U17995 (N_17995,N_13192,N_13887);
nor U17996 (N_17996,N_14765,N_14479);
xnor U17997 (N_17997,N_12363,N_12757);
or U17998 (N_17998,N_14487,N_14940);
nor U17999 (N_17999,N_14494,N_13286);
nand U18000 (N_18000,N_15010,N_15667);
nand U18001 (N_18001,N_16843,N_17653);
xnor U18002 (N_18002,N_17537,N_15128);
or U18003 (N_18003,N_15066,N_16271);
xor U18004 (N_18004,N_16071,N_16155);
xor U18005 (N_18005,N_15473,N_17941);
nand U18006 (N_18006,N_15904,N_17367);
and U18007 (N_18007,N_16928,N_15651);
and U18008 (N_18008,N_16226,N_17202);
xnor U18009 (N_18009,N_16372,N_17519);
or U18010 (N_18010,N_16416,N_16799);
xnor U18011 (N_18011,N_16009,N_15301);
nand U18012 (N_18012,N_16542,N_17740);
nand U18013 (N_18013,N_17731,N_15238);
nand U18014 (N_18014,N_17961,N_16289);
nor U18015 (N_18015,N_15927,N_16350);
or U18016 (N_18016,N_16688,N_15071);
xnor U18017 (N_18017,N_17177,N_17084);
nand U18018 (N_18018,N_15877,N_15022);
or U18019 (N_18019,N_17021,N_15021);
xnor U18020 (N_18020,N_16726,N_15892);
and U18021 (N_18021,N_15724,N_16019);
nor U18022 (N_18022,N_16947,N_15858);
xnor U18023 (N_18023,N_17201,N_15767);
and U18024 (N_18024,N_17564,N_15034);
nand U18025 (N_18025,N_15109,N_16092);
nand U18026 (N_18026,N_16442,N_16180);
and U18027 (N_18027,N_16426,N_15910);
nor U18028 (N_18028,N_15084,N_15854);
xnor U18029 (N_18029,N_15100,N_17075);
and U18030 (N_18030,N_16079,N_17678);
and U18031 (N_18031,N_17701,N_17083);
nand U18032 (N_18032,N_16620,N_17390);
and U18033 (N_18033,N_16785,N_17280);
xor U18034 (N_18034,N_16411,N_15259);
xnor U18035 (N_18035,N_17078,N_16855);
or U18036 (N_18036,N_17552,N_17064);
nand U18037 (N_18037,N_16779,N_16508);
nor U18038 (N_18038,N_17873,N_15722);
nor U18039 (N_18039,N_15857,N_16388);
xnor U18040 (N_18040,N_15305,N_15993);
nand U18041 (N_18041,N_17425,N_17957);
or U18042 (N_18042,N_16266,N_16122);
and U18043 (N_18043,N_16057,N_15228);
and U18044 (N_18044,N_16607,N_16600);
nor U18045 (N_18045,N_16359,N_15578);
nand U18046 (N_18046,N_16356,N_17693);
xor U18047 (N_18047,N_16935,N_15367);
nor U18048 (N_18048,N_16588,N_17912);
nor U18049 (N_18049,N_17374,N_17560);
nor U18050 (N_18050,N_15064,N_17687);
nand U18051 (N_18051,N_17682,N_17447);
nand U18052 (N_18052,N_16938,N_16466);
and U18053 (N_18053,N_16351,N_15822);
nor U18054 (N_18054,N_17065,N_15374);
or U18055 (N_18055,N_16169,N_17484);
xor U18056 (N_18056,N_15634,N_15516);
xor U18057 (N_18057,N_17950,N_15496);
xnor U18058 (N_18058,N_17130,N_16500);
xor U18059 (N_18059,N_15011,N_15629);
nor U18060 (N_18060,N_16946,N_17115);
and U18061 (N_18061,N_17587,N_16605);
nor U18062 (N_18062,N_15918,N_16478);
or U18063 (N_18063,N_15658,N_16167);
xor U18064 (N_18064,N_16974,N_15221);
nand U18065 (N_18065,N_15354,N_16750);
nand U18066 (N_18066,N_17936,N_15674);
xor U18067 (N_18067,N_16433,N_15134);
xor U18068 (N_18068,N_17772,N_16247);
xor U18069 (N_18069,N_16093,N_16288);
or U18070 (N_18070,N_16677,N_16049);
nor U18071 (N_18071,N_16285,N_16082);
xor U18072 (N_18072,N_17755,N_15239);
nor U18073 (N_18073,N_15597,N_17306);
nor U18074 (N_18074,N_15984,N_17397);
xnor U18075 (N_18075,N_17190,N_17947);
or U18076 (N_18076,N_17145,N_17018);
and U18077 (N_18077,N_15944,N_15060);
and U18078 (N_18078,N_15465,N_16591);
and U18079 (N_18079,N_16203,N_17281);
xnor U18080 (N_18080,N_15309,N_16908);
nand U18081 (N_18081,N_15342,N_15535);
or U18082 (N_18082,N_17574,N_17795);
nand U18083 (N_18083,N_17316,N_15181);
or U18084 (N_18084,N_15958,N_16905);
xnor U18085 (N_18085,N_16526,N_16994);
nand U18086 (N_18086,N_16460,N_17747);
xor U18087 (N_18087,N_15205,N_16450);
and U18088 (N_18088,N_16875,N_15734);
nand U18089 (N_18089,N_16746,N_16244);
nand U18090 (N_18090,N_15498,N_15824);
nand U18091 (N_18091,N_17834,N_17315);
xor U18092 (N_18092,N_16457,N_17435);
or U18093 (N_18093,N_15063,N_17714);
nor U18094 (N_18094,N_15549,N_16102);
nor U18095 (N_18095,N_15188,N_15691);
xnor U18096 (N_18096,N_15726,N_16499);
nor U18097 (N_18097,N_16303,N_17489);
nand U18098 (N_18098,N_16566,N_16171);
nand U18099 (N_18099,N_15298,N_16486);
nor U18100 (N_18100,N_17467,N_15398);
xnor U18101 (N_18101,N_16116,N_17502);
or U18102 (N_18102,N_15540,N_16561);
xnor U18103 (N_18103,N_16802,N_15385);
nor U18104 (N_18104,N_16850,N_16780);
nor U18105 (N_18105,N_15326,N_16412);
and U18106 (N_18106,N_15056,N_17054);
or U18107 (N_18107,N_16624,N_15153);
nor U18108 (N_18108,N_15511,N_17840);
or U18109 (N_18109,N_15327,N_15289);
nor U18110 (N_18110,N_17407,N_15005);
xnor U18111 (N_18111,N_17849,N_17348);
nor U18112 (N_18112,N_16253,N_17762);
xnor U18113 (N_18113,N_16805,N_15121);
or U18114 (N_18114,N_15761,N_16212);
and U18115 (N_18115,N_16157,N_16306);
nor U18116 (N_18116,N_16282,N_15358);
xor U18117 (N_18117,N_17850,N_17010);
nand U18118 (N_18118,N_15210,N_15512);
or U18119 (N_18119,N_15889,N_15397);
nand U18120 (N_18120,N_15796,N_17480);
or U18121 (N_18121,N_16211,N_15423);
and U18122 (N_18122,N_15912,N_16518);
nand U18123 (N_18123,N_17323,N_17505);
and U18124 (N_18124,N_15092,N_16414);
nand U18125 (N_18125,N_17188,N_17392);
nand U18126 (N_18126,N_15303,N_17198);
or U18127 (N_18127,N_17784,N_17427);
xor U18128 (N_18128,N_15286,N_17800);
xor U18129 (N_18129,N_17943,N_15916);
and U18130 (N_18130,N_16208,N_15735);
xor U18131 (N_18131,N_17847,N_17210);
or U18132 (N_18132,N_15563,N_15365);
and U18133 (N_18133,N_16362,N_16047);
nor U18134 (N_18134,N_16503,N_16966);
or U18135 (N_18135,N_17458,N_15161);
and U18136 (N_18136,N_17883,N_15719);
xor U18137 (N_18137,N_17692,N_16610);
and U18138 (N_18138,N_15320,N_16309);
nor U18139 (N_18139,N_15001,N_16490);
nand U18140 (N_18140,N_16073,N_17462);
nand U18141 (N_18141,N_17414,N_17911);
and U18142 (N_18142,N_16926,N_16396);
or U18143 (N_18143,N_16196,N_16158);
xnor U18144 (N_18144,N_15567,N_16936);
nor U18145 (N_18145,N_16202,N_16817);
nand U18146 (N_18146,N_15560,N_17403);
and U18147 (N_18147,N_16540,N_17270);
or U18148 (N_18148,N_17142,N_16353);
nand U18149 (N_18149,N_17832,N_17421);
xor U18150 (N_18150,N_15452,N_15688);
or U18151 (N_18151,N_15939,N_16764);
or U18152 (N_18152,N_17454,N_16828);
or U18153 (N_18153,N_15720,N_15979);
nand U18154 (N_18154,N_15868,N_16614);
xor U18155 (N_18155,N_15584,N_15083);
nand U18156 (N_18156,N_16858,N_16280);
nand U18157 (N_18157,N_16962,N_17660);
nor U18158 (N_18158,N_16681,N_15282);
nand U18159 (N_18159,N_17120,N_17759);
nand U18160 (N_18160,N_15475,N_17944);
or U18161 (N_18161,N_15234,N_16618);
nor U18162 (N_18162,N_15368,N_16279);
and U18163 (N_18163,N_17684,N_17438);
and U18164 (N_18164,N_17758,N_16432);
nor U18165 (N_18165,N_16123,N_16434);
xnor U18166 (N_18166,N_15712,N_15410);
xor U18167 (N_18167,N_16492,N_17955);
nand U18168 (N_18168,N_17456,N_15055);
and U18169 (N_18169,N_15998,N_17196);
nand U18170 (N_18170,N_16842,N_16128);
nand U18171 (N_18171,N_16363,N_17636);
xor U18172 (N_18172,N_17634,N_17804);
or U18173 (N_18173,N_17650,N_17967);
or U18174 (N_18174,N_17624,N_16165);
nor U18175 (N_18175,N_15330,N_15631);
nor U18176 (N_18176,N_16734,N_17287);
or U18177 (N_18177,N_17540,N_16201);
nor U18178 (N_18178,N_16902,N_16330);
and U18179 (N_18179,N_17189,N_16653);
or U18180 (N_18180,N_15745,N_16277);
and U18181 (N_18181,N_16660,N_15522);
xor U18182 (N_18182,N_17426,N_15710);
and U18183 (N_18183,N_16294,N_15606);
or U18184 (N_18184,N_16172,N_16907);
or U18185 (N_18185,N_16596,N_15204);
or U18186 (N_18186,N_15569,N_16794);
xnor U18187 (N_18187,N_17872,N_16814);
xor U18188 (N_18188,N_17935,N_15002);
or U18189 (N_18189,N_16737,N_17289);
nand U18190 (N_18190,N_17016,N_15811);
xor U18191 (N_18191,N_15017,N_17530);
and U18192 (N_18192,N_16328,N_16404);
or U18193 (N_18193,N_16238,N_15896);
nand U18194 (N_18194,N_15448,N_17471);
or U18195 (N_18195,N_15028,N_17052);
or U18196 (N_18196,N_16455,N_17900);
nand U18197 (N_18197,N_17138,N_15440);
and U18198 (N_18198,N_16224,N_15510);
and U18199 (N_18199,N_15031,N_16872);
or U18200 (N_18200,N_16762,N_16704);
and U18201 (N_18201,N_15006,N_15400);
xor U18202 (N_18202,N_17495,N_16090);
xnor U18203 (N_18203,N_16844,N_17633);
nand U18204 (N_18204,N_16336,N_15463);
and U18205 (N_18205,N_15739,N_17193);
and U18206 (N_18206,N_15343,N_16945);
and U18207 (N_18207,N_16243,N_16748);
xor U18208 (N_18208,N_17441,N_16538);
nand U18209 (N_18209,N_17446,N_16340);
nand U18210 (N_18210,N_15237,N_16217);
nand U18211 (N_18211,N_15543,N_15494);
or U18212 (N_18212,N_17736,N_17744);
nor U18213 (N_18213,N_16106,N_15587);
nor U18214 (N_18214,N_17773,N_15786);
nor U18215 (N_18215,N_17350,N_16484);
and U18216 (N_18216,N_16459,N_16273);
xnor U18217 (N_18217,N_15191,N_17111);
and U18218 (N_18218,N_15319,N_17112);
xnor U18219 (N_18219,N_15190,N_17962);
nor U18220 (N_18220,N_16602,N_15633);
nor U18221 (N_18221,N_15808,N_16195);
nor U18222 (N_18222,N_16870,N_15257);
and U18223 (N_18223,N_17182,N_15247);
xnor U18224 (N_18224,N_15971,N_15997);
nand U18225 (N_18225,N_17924,N_16531);
xnor U18226 (N_18226,N_17014,N_16437);
nor U18227 (N_18227,N_15392,N_15794);
nand U18228 (N_18228,N_16925,N_17931);
and U18229 (N_18229,N_16310,N_17305);
nor U18230 (N_18230,N_16703,N_15758);
xor U18231 (N_18231,N_16581,N_16215);
nand U18232 (N_18232,N_15562,N_16701);
nor U18233 (N_18233,N_16996,N_15729);
or U18234 (N_18234,N_15533,N_17385);
nand U18235 (N_18235,N_17207,N_15402);
xnor U18236 (N_18236,N_16407,N_15603);
nor U18237 (N_18237,N_17308,N_17696);
nand U18238 (N_18238,N_17837,N_15447);
or U18239 (N_18239,N_16075,N_15050);
or U18240 (N_18240,N_17341,N_15474);
nand U18241 (N_18241,N_16747,N_17673);
xnor U18242 (N_18242,N_17139,N_15306);
or U18243 (N_18243,N_15941,N_15417);
xnor U18244 (N_18244,N_15746,N_17987);
and U18245 (N_18245,N_16707,N_15530);
nand U18246 (N_18246,N_17183,N_17585);
or U18247 (N_18247,N_15420,N_17171);
or U18248 (N_18248,N_16989,N_16237);
and U18249 (N_18249,N_16589,N_17160);
and U18250 (N_18250,N_15863,N_17365);
nand U18251 (N_18251,N_17137,N_15702);
nand U18252 (N_18252,N_16399,N_15509);
and U18253 (N_18253,N_17711,N_17806);
or U18254 (N_18254,N_17732,N_17440);
and U18255 (N_18255,N_17690,N_16101);
nor U18256 (N_18256,N_17117,N_16972);
nand U18257 (N_18257,N_15241,N_15311);
nor U18258 (N_18258,N_15831,N_16360);
nor U18259 (N_18259,N_15801,N_16326);
and U18260 (N_18260,N_15964,N_16252);
and U18261 (N_18261,N_17577,N_16213);
or U18262 (N_18262,N_17877,N_17321);
and U18263 (N_18263,N_17922,N_17284);
nand U18264 (N_18264,N_17251,N_17561);
nand U18265 (N_18265,N_15933,N_16804);
nand U18266 (N_18266,N_17702,N_17035);
nand U18267 (N_18267,N_15093,N_16862);
nor U18268 (N_18268,N_17878,N_16502);
nor U18269 (N_18269,N_17149,N_17179);
or U18270 (N_18270,N_17622,N_16942);
or U18271 (N_18271,N_16713,N_16959);
xor U18272 (N_18272,N_16118,N_15043);
nand U18273 (N_18273,N_15880,N_17896);
nor U18274 (N_18274,N_15192,N_15791);
nor U18275 (N_18275,N_15523,N_17663);
nor U18276 (N_18276,N_15037,N_15212);
xnor U18277 (N_18277,N_16173,N_16343);
and U18278 (N_18278,N_16002,N_17038);
or U18279 (N_18279,N_17356,N_17610);
or U18280 (N_18280,N_16772,N_17135);
and U18281 (N_18281,N_17897,N_16986);
nand U18282 (N_18282,N_15898,N_15125);
nand U18283 (N_18283,N_16714,N_17887);
or U18284 (N_18284,N_17646,N_16927);
or U18285 (N_18285,N_15159,N_15054);
nand U18286 (N_18286,N_16738,N_15390);
nor U18287 (N_18287,N_15931,N_16829);
nand U18288 (N_18288,N_16117,N_15682);
xnor U18289 (N_18289,N_17700,N_17378);
xnor U18290 (N_18290,N_16567,N_15577);
xnor U18291 (N_18291,N_15076,N_17158);
or U18292 (N_18292,N_16443,N_16394);
nand U18293 (N_18293,N_15980,N_16921);
or U18294 (N_18294,N_15271,N_16448);
nand U18295 (N_18295,N_15425,N_17531);
and U18296 (N_18296,N_16262,N_16633);
and U18297 (N_18297,N_17485,N_16022);
and U18298 (N_18298,N_17926,N_16979);
xor U18299 (N_18299,N_17580,N_16852);
xor U18300 (N_18300,N_15506,N_15059);
or U18301 (N_18301,N_15690,N_17890);
xor U18302 (N_18302,N_15936,N_16696);
and U18303 (N_18303,N_16819,N_16883);
nand U18304 (N_18304,N_15591,N_16788);
nand U18305 (N_18305,N_16191,N_15642);
or U18306 (N_18306,N_15777,N_15756);
or U18307 (N_18307,N_16899,N_16851);
nand U18308 (N_18308,N_15990,N_15748);
and U18309 (N_18309,N_15296,N_15278);
or U18310 (N_18310,N_15977,N_16425);
xnor U18311 (N_18311,N_15357,N_15950);
nor U18312 (N_18312,N_16291,N_16261);
xnor U18313 (N_18313,N_15760,N_17303);
xnor U18314 (N_18314,N_17599,N_15482);
or U18315 (N_18315,N_16084,N_15461);
nand U18316 (N_18316,N_15946,N_17937);
xnor U18317 (N_18317,N_17853,N_17802);
nand U18318 (N_18318,N_17534,N_16242);
nand U18319 (N_18319,N_16783,N_16898);
nand U18320 (N_18320,N_15105,N_17881);
nor U18321 (N_18321,N_16771,N_17211);
nand U18322 (N_18322,N_16656,N_15266);
nor U18323 (N_18323,N_15809,N_16355);
and U18324 (N_18324,N_17874,N_17645);
nor U18325 (N_18325,N_15272,N_15829);
nor U18326 (N_18326,N_16790,N_16239);
nand U18327 (N_18327,N_15143,N_16884);
nor U18328 (N_18328,N_16781,N_15972);
or U18329 (N_18329,N_17709,N_17413);
nor U18330 (N_18330,N_16107,N_17088);
xnor U18331 (N_18331,N_17745,N_16012);
and U18332 (N_18332,N_16729,N_16811);
xor U18333 (N_18333,N_17325,N_15360);
and U18334 (N_18334,N_17357,N_16497);
or U18335 (N_18335,N_16577,N_15260);
nor U18336 (N_18336,N_16645,N_15352);
xnor U18337 (N_18337,N_16769,N_16164);
or U18338 (N_18338,N_15097,N_15859);
nor U18339 (N_18339,N_16661,N_16881);
xor U18340 (N_18340,N_16527,N_16999);
nor U18341 (N_18341,N_15661,N_15781);
nor U18342 (N_18342,N_16131,N_17750);
nor U18343 (N_18343,N_17913,N_17856);
nand U18344 (N_18344,N_16274,N_16732);
or U18345 (N_18345,N_16763,N_17169);
nor U18346 (N_18346,N_15351,N_15182);
nand U18347 (N_18347,N_17798,N_17161);
or U18348 (N_18348,N_16672,N_15771);
and U18349 (N_18349,N_16377,N_16827);
nand U18350 (N_18350,N_15229,N_15736);
nor U18351 (N_18351,N_17722,N_15308);
nand U18352 (N_18352,N_16476,N_17200);
and U18353 (N_18353,N_16608,N_15407);
or U18354 (N_18354,N_16839,N_17285);
nor U18355 (N_18355,N_15566,N_16795);
nand U18356 (N_18356,N_15478,N_15693);
or U18357 (N_18357,N_16050,N_16322);
or U18358 (N_18358,N_16612,N_17974);
or U18359 (N_18359,N_15172,N_17141);
or U18360 (N_18360,N_17619,N_17277);
nand U18361 (N_18361,N_16345,N_15960);
nor U18362 (N_18362,N_15520,N_17019);
nand U18363 (N_18363,N_15665,N_15222);
and U18364 (N_18364,N_17867,N_16179);
xor U18365 (N_18365,N_15932,N_17862);
xor U18366 (N_18366,N_15321,N_15647);
xor U18367 (N_18367,N_17865,N_17265);
nand U18368 (N_18368,N_15279,N_16162);
xnor U18369 (N_18369,N_16885,N_17898);
or U18370 (N_18370,N_16332,N_17243);
xor U18371 (N_18371,N_17888,N_16334);
xor U18372 (N_18372,N_16985,N_17493);
nand U18373 (N_18373,N_15759,N_16472);
nand U18374 (N_18374,N_17317,N_17094);
nor U18375 (N_18375,N_17347,N_17973);
or U18376 (N_18376,N_16756,N_15952);
or U18377 (N_18377,N_15000,N_17159);
xnor U18378 (N_18378,N_15508,N_15363);
or U18379 (N_18379,N_15836,N_17398);
and U18380 (N_18380,N_17011,N_16658);
or U18381 (N_18381,N_17551,N_15135);
nor U18382 (N_18382,N_17370,N_17601);
or U18383 (N_18383,N_15707,N_17241);
xnor U18384 (N_18384,N_15903,N_17570);
or U18385 (N_18385,N_17060,N_16134);
xor U18386 (N_18386,N_17445,N_15637);
nor U18387 (N_18387,N_16630,N_15524);
xnor U18388 (N_18388,N_16535,N_17409);
and U18389 (N_18389,N_15185,N_15430);
or U18390 (N_18390,N_16583,N_16384);
nand U18391 (N_18391,N_15138,N_17015);
or U18392 (N_18392,N_17632,N_15685);
nor U18393 (N_18393,N_17659,N_15164);
xor U18394 (N_18394,N_16055,N_17566);
nor U18395 (N_18395,N_15486,N_15754);
or U18396 (N_18396,N_17521,N_16586);
and U18397 (N_18397,N_17465,N_16944);
xnor U18398 (N_18398,N_15244,N_16861);
nand U18399 (N_18399,N_16408,N_15536);
nor U18400 (N_18400,N_17379,N_15047);
nor U18401 (N_18401,N_17146,N_15334);
nand U18402 (N_18402,N_17079,N_16185);
xnor U18403 (N_18403,N_16523,N_15004);
and U18404 (N_18404,N_16320,N_15118);
nor U18405 (N_18405,N_16496,N_15090);
nand U18406 (N_18406,N_15618,N_17020);
nand U18407 (N_18407,N_17855,N_15828);
and U18408 (N_18408,N_17107,N_17334);
xnor U18409 (N_18409,N_16520,N_15455);
and U18410 (N_18410,N_17103,N_17351);
or U18411 (N_18411,N_17915,N_17882);
xor U18412 (N_18412,N_17501,N_15146);
xnor U18413 (N_18413,N_16062,N_16451);
and U18414 (N_18414,N_17920,N_15677);
or U18415 (N_18415,N_17212,N_15915);
and U18416 (N_18416,N_16801,N_17036);
xnor U18417 (N_18417,N_16449,N_16904);
nand U18418 (N_18418,N_17022,N_17373);
or U18419 (N_18419,N_16255,N_17272);
nor U18420 (N_18420,N_17528,N_16143);
and U18421 (N_18421,N_17082,N_16557);
xor U18422 (N_18422,N_16813,N_17304);
nand U18423 (N_18423,N_17366,N_15436);
xor U18424 (N_18424,N_15708,N_15703);
nor U18425 (N_18425,N_16717,N_15403);
nand U18426 (N_18426,N_17354,N_16680);
nand U18427 (N_18427,N_15951,N_15048);
or U18428 (N_18428,N_15626,N_15865);
and U18429 (N_18429,N_16678,N_17364);
and U18430 (N_18430,N_16391,N_15197);
or U18431 (N_18431,N_17852,N_15202);
or U18432 (N_18432,N_16465,N_15068);
or U18433 (N_18433,N_15832,N_17230);
nand U18434 (N_18434,N_16318,N_16951);
nor U18435 (N_18435,N_16774,N_15428);
nand U18436 (N_18436,N_17343,N_17028);
nand U18437 (N_18437,N_16300,N_16447);
or U18438 (N_18438,N_16514,N_15624);
nand U18439 (N_18439,N_16969,N_17007);
xnor U18440 (N_18440,N_17591,N_17583);
xnor U18441 (N_18441,N_17375,N_15978);
xnor U18442 (N_18442,N_15639,N_16980);
and U18443 (N_18443,N_15467,N_16880);
or U18444 (N_18444,N_17098,N_17854);
or U18445 (N_18445,N_16420,N_16715);
xor U18446 (N_18446,N_17013,N_16192);
and U18447 (N_18447,N_16267,N_15627);
and U18448 (N_18448,N_16406,N_15833);
nor U18449 (N_18449,N_17777,N_16924);
or U18450 (N_18450,N_16991,N_16887);
nand U18451 (N_18451,N_16541,N_16487);
and U18452 (N_18452,N_16960,N_15947);
xnor U18453 (N_18453,N_17637,N_15580);
nand U18454 (N_18454,N_16579,N_16826);
nor U18455 (N_18455,N_17542,N_16439);
nor U18456 (N_18456,N_16682,N_15929);
and U18457 (N_18457,N_16941,N_17655);
nand U18458 (N_18458,N_17844,N_17490);
and U18459 (N_18459,N_17868,N_17005);
nand U18460 (N_18460,N_15706,N_16537);
or U18461 (N_18461,N_17733,N_15356);
nand U18462 (N_18462,N_17199,N_15740);
nand U18463 (N_18463,N_16637,N_17545);
or U18464 (N_18464,N_17661,N_15556);
and U18465 (N_18465,N_15341,N_17556);
xor U18466 (N_18466,N_17361,N_15335);
or U18467 (N_18467,N_17990,N_16675);
or U18468 (N_18468,N_15030,N_17851);
nand U18469 (N_18469,N_17995,N_16014);
xor U18470 (N_18470,N_15995,N_15923);
nand U18471 (N_18471,N_16739,N_17768);
or U18472 (N_18472,N_15446,N_16066);
nor U18473 (N_18473,N_16988,N_17630);
and U18474 (N_18474,N_17807,N_15399);
xor U18475 (N_18475,N_17536,N_17677);
xnor U18476 (N_18476,N_17954,N_15554);
nor U18477 (N_18477,N_15236,N_16767);
or U18478 (N_18478,N_17563,N_16137);
nor U18479 (N_18479,N_15422,N_15492);
nor U18480 (N_18480,N_15663,N_17638);
xor U18481 (N_18481,N_16615,N_16222);
xor U18482 (N_18482,N_15379,N_16386);
nand U18483 (N_18483,N_16635,N_17008);
and U18484 (N_18484,N_16975,N_16958);
or U18485 (N_18485,N_16818,N_16534);
nand U18486 (N_18486,N_15982,N_15968);
and U18487 (N_18487,N_15541,N_16536);
and U18488 (N_18488,N_17506,N_17104);
nand U18489 (N_18489,N_15925,N_16652);
xor U18490 (N_18490,N_16664,N_17618);
nand U18491 (N_18491,N_16385,N_15458);
xnor U18492 (N_18492,N_17156,N_15668);
nor U18493 (N_18493,N_15199,N_17464);
nand U18494 (N_18494,N_16454,N_15999);
and U18495 (N_18495,N_15813,N_17620);
and U18496 (N_18496,N_16796,N_15970);
nand U18497 (N_18497,N_17573,N_16335);
nor U18498 (N_18498,N_16275,N_16631);
nand U18499 (N_18499,N_15209,N_16918);
and U18500 (N_18500,N_17492,N_15853);
xnor U18501 (N_18501,N_16110,N_15426);
or U18502 (N_18502,N_16329,N_17051);
xor U18503 (N_18503,N_16445,N_16961);
nor U18504 (N_18504,N_16530,N_17891);
xnor U18505 (N_18505,N_15307,N_16270);
xnor U18506 (N_18506,N_15476,N_17165);
xor U18507 (N_18507,N_15787,N_15847);
xor U18508 (N_18508,N_17823,N_16903);
and U18509 (N_18509,N_15041,N_16063);
nor U18510 (N_18510,N_15101,N_16401);
or U18511 (N_18511,N_15825,N_15208);
and U18512 (N_18512,N_15928,N_15504);
xnor U18513 (N_18513,N_15583,N_17623);
nand U18514 (N_18514,N_16906,N_17314);
or U18515 (N_18515,N_15645,N_17032);
nor U18516 (N_18516,N_17337,N_15263);
xnor U18517 (N_18517,N_16864,N_15728);
xor U18518 (N_18518,N_15881,N_16272);
xor U18519 (N_18519,N_16929,N_15827);
and U18520 (N_18520,N_15292,N_17070);
nor U18521 (N_18521,N_17656,N_17468);
or U18522 (N_18522,N_17989,N_17603);
and U18523 (N_18523,N_16295,N_15453);
and U18524 (N_18524,N_15945,N_15439);
nor U18525 (N_18525,N_15015,N_17925);
nor U18526 (N_18526,N_15894,N_16751);
and U18527 (N_18527,N_15033,N_16923);
or U18528 (N_18528,N_15336,N_16026);
xor U18529 (N_18529,N_16654,N_16712);
xnor U18530 (N_18530,N_17526,N_16606);
xor U18531 (N_18531,N_16422,N_16841);
and U18532 (N_18532,N_15249,N_17932);
and U18533 (N_18533,N_17071,N_17738);
nand U18534 (N_18534,N_17140,N_17473);
nand U18535 (N_18535,N_15318,N_15937);
nand U18536 (N_18536,N_17606,N_15270);
and U18537 (N_18537,N_17205,N_17095);
nor U18538 (N_18538,N_15391,N_16348);
xor U18539 (N_18539,N_15669,N_15924);
or U18540 (N_18540,N_16036,N_17557);
nand U18541 (N_18541,N_16138,N_15875);
and U18542 (N_18542,N_16659,N_17597);
or U18543 (N_18543,N_16375,N_15184);
or U18544 (N_18544,N_17516,N_15819);
nand U18545 (N_18545,N_17143,N_17533);
or U18546 (N_18546,N_15200,N_16909);
nand U18547 (N_18547,N_15542,N_16504);
xor U18548 (N_18548,N_16749,N_17588);
nand U18549 (N_18549,N_17754,N_15613);
or U18550 (N_18550,N_16667,N_17914);
nand U18551 (N_18551,N_15170,N_16364);
xnor U18552 (N_18552,N_15376,N_15917);
and U18553 (N_18553,N_16109,N_17001);
nor U18554 (N_18554,N_16916,N_17191);
or U18555 (N_18555,N_16494,N_17809);
nor U18556 (N_18556,N_17250,N_15802);
xor U18557 (N_18557,N_16025,N_16745);
and U18558 (N_18558,N_16488,N_17981);
and U18559 (N_18559,N_17726,N_15207);
nor U18560 (N_18560,N_17319,N_15163);
xor U18561 (N_18561,N_17721,N_16882);
and U18562 (N_18562,N_17349,N_15457);
or U18563 (N_18563,N_16040,N_16188);
xor U18564 (N_18564,N_17568,N_15895);
xnor U18565 (N_18565,N_15466,N_15572);
or U18566 (N_18566,N_15805,N_17017);
xor U18567 (N_18567,N_15907,N_16331);
and U18568 (N_18568,N_17735,N_16551);
or U18569 (N_18569,N_15044,N_17443);
xor U18570 (N_18570,N_15856,N_17828);
xnor U18571 (N_18571,N_15561,N_15948);
xor U18572 (N_18572,N_17206,N_16221);
and U18573 (N_18573,N_15559,N_17664);
xor U18574 (N_18574,N_17386,N_17024);
nand U18575 (N_18575,N_17286,N_15179);
xor U18576 (N_18576,N_15713,N_17598);
nor U18577 (N_18577,N_17266,N_17037);
or U18578 (N_18578,N_15650,N_15388);
xor U18579 (N_18579,N_16148,N_16254);
nand U18580 (N_18580,N_15839,N_17513);
xor U18581 (N_18581,N_16145,N_16676);
and U18582 (N_18582,N_15792,N_15821);
or U18583 (N_18583,N_17845,N_15413);
nand U18584 (N_18584,N_16831,N_15954);
nand U18585 (N_18585,N_16768,N_16836);
xnor U18586 (N_18586,N_15414,N_16064);
and U18587 (N_18587,N_16013,N_15695);
nor U18588 (N_18588,N_17510,N_16061);
xnor U18589 (N_18589,N_15887,N_16184);
or U18590 (N_18590,N_17951,N_16077);
xor U18591 (N_18591,N_15518,N_15145);
and U18592 (N_18592,N_15886,N_15198);
or U18593 (N_18593,N_15016,N_15250);
xnor U18594 (N_18594,N_15171,N_15600);
nand U18595 (N_18595,N_16886,N_15313);
and U18596 (N_18596,N_16321,N_17031);
nand U18597 (N_18597,N_16483,N_15850);
nand U18598 (N_18598,N_15380,N_17991);
and U18599 (N_18599,N_17249,N_15243);
nand U18600 (N_18600,N_15122,N_17411);
nand U18601 (N_18601,N_16319,N_16965);
xor U18602 (N_18602,N_16773,N_15798);
nor U18603 (N_18603,N_17822,N_17483);
nor U18604 (N_18604,N_15959,N_15225);
and U18605 (N_18605,N_17608,N_17461);
and U18606 (N_18606,N_16395,N_16176);
nor U18607 (N_18607,N_16227,N_16327);
nor U18608 (N_18608,N_15725,N_16462);
nand U18609 (N_18609,N_16891,N_15525);
xnor U18610 (N_18610,N_15408,N_15539);
or U18611 (N_18611,N_17734,N_15750);
and U18612 (N_18612,N_17174,N_17448);
nor U18613 (N_18613,N_17699,N_17058);
or U18614 (N_18614,N_16821,N_15681);
nor U18615 (N_18615,N_15994,N_15186);
xor U18616 (N_18616,N_17705,N_15555);
nor U18617 (N_18617,N_16413,N_17979);
and U18618 (N_18618,N_15919,N_16968);
nand U18619 (N_18619,N_15009,N_15855);
nor U18620 (N_18620,N_16132,N_17707);
xor U18621 (N_18621,N_17056,N_15816);
and U18622 (N_18622,N_15773,N_16627);
and U18623 (N_18623,N_16302,N_16142);
or U18624 (N_18624,N_17360,N_16039);
or U18625 (N_18625,N_15862,N_17430);
xnor U18626 (N_18626,N_15488,N_16901);
nor U18627 (N_18627,N_15395,N_17100);
nor U18628 (N_18628,N_16791,N_15206);
nand U18629 (N_18629,N_15123,N_17668);
and U18630 (N_18630,N_15957,N_17739);
or U18631 (N_18631,N_17916,N_17523);
and U18632 (N_18632,N_16939,N_17248);
and U18633 (N_18633,N_16601,N_16950);
nor U18634 (N_18634,N_17718,N_17106);
and U18635 (N_18635,N_15934,N_15538);
nor U18636 (N_18636,N_17909,N_15529);
nor U18637 (N_18637,N_16840,N_15752);
nand U18638 (N_18638,N_15527,N_15765);
or U18639 (N_18639,N_17899,N_17121);
nand U18640 (N_18640,N_17134,N_17969);
nand U18641 (N_18641,N_15053,N_17670);
nor U18642 (N_18642,N_17794,N_16370);
nand U18643 (N_18643,N_16911,N_15723);
nand U18644 (N_18644,N_15177,N_16544);
nor U18645 (N_18645,N_17220,N_16054);
nand U18646 (N_18646,N_16876,N_17399);
nand U18647 (N_18647,N_17450,N_17444);
nor U18648 (N_18648,N_16546,N_15070);
nor U18649 (N_18649,N_17442,N_16919);
nor U18650 (N_18650,N_15845,N_15470);
xnor U18651 (N_18651,N_16873,N_17090);
and U18652 (N_18652,N_17716,N_16456);
or U18653 (N_18653,N_16957,N_15045);
nor U18654 (N_18654,N_15666,N_16382);
or U18655 (N_18655,N_16058,N_15909);
and U18656 (N_18656,N_17820,N_17689);
xnor U18657 (N_18657,N_15291,N_15843);
nor U18658 (N_18658,N_17328,N_17760);
or U18659 (N_18659,N_15867,N_17857);
or U18660 (N_18660,N_16074,N_16210);
nor U18661 (N_18661,N_16807,N_17841);
nand U18662 (N_18662,N_17387,N_17945);
nor U18663 (N_18663,N_15974,N_17547);
xnor U18664 (N_18664,N_15742,N_16341);
and U18665 (N_18665,N_17894,N_15571);
nor U18666 (N_18666,N_15671,N_15797);
or U18667 (N_18667,N_15051,N_15073);
nand U18668 (N_18668,N_16639,N_15443);
nor U18669 (N_18669,N_16889,N_16430);
nand U18670 (N_18670,N_16311,N_17746);
and U18671 (N_18671,N_17066,N_15727);
and U18672 (N_18672,N_15148,N_17676);
or U18673 (N_18673,N_15775,N_15680);
and U18674 (N_18674,N_17429,N_16119);
nand U18675 (N_18675,N_17584,N_16298);
nor U18676 (N_18676,N_17876,N_16815);
xnor U18677 (N_18677,N_17672,N_16177);
xnor U18678 (N_18678,N_16981,N_17675);
or U18679 (N_18679,N_17785,N_17368);
nand U18680 (N_18680,N_17769,N_16046);
xor U18681 (N_18681,N_16421,N_15333);
and U18682 (N_18682,N_17340,N_17215);
or U18683 (N_18683,N_17596,N_16083);
nand U18684 (N_18684,N_15393,N_16622);
or U18685 (N_18685,N_16207,N_17296);
nand U18686 (N_18686,N_15120,N_16963);
or U18687 (N_18687,N_15694,N_17657);
or U18688 (N_18688,N_16035,N_16263);
nor U18689 (N_18689,N_15632,N_17748);
and U18690 (N_18690,N_16147,N_15872);
or U18691 (N_18691,N_16553,N_17482);
nor U18692 (N_18692,N_17209,N_15721);
or U18693 (N_18693,N_17420,N_15459);
or U18694 (N_18694,N_15468,N_16133);
xnor U18695 (N_18695,N_15770,N_15804);
nand U18696 (N_18696,N_15277,N_17475);
or U18697 (N_18697,N_17363,N_16043);
xor U18698 (N_18698,N_15018,N_16325);
nand U18699 (N_18699,N_15844,N_16765);
xnor U18700 (N_18700,N_15860,N_17072);
or U18701 (N_18701,N_17976,N_17166);
nor U18702 (N_18702,N_16307,N_16381);
nor U18703 (N_18703,N_16727,N_16709);
nor U18704 (N_18704,N_15089,N_16069);
or U18705 (N_18705,N_15955,N_17767);
xnor U18706 (N_18706,N_16940,N_15477);
and U18707 (N_18707,N_16027,N_15852);
xor U18708 (N_18708,N_15019,N_16097);
or U18709 (N_18709,N_16129,N_15830);
nand U18710 (N_18710,N_15072,N_16599);
xnor U18711 (N_18711,N_16087,N_15345);
nand U18712 (N_18712,N_16973,N_16113);
xnor U18713 (N_18713,N_16250,N_15265);
nand U18714 (N_18714,N_15676,N_17412);
xor U18715 (N_18715,N_17532,N_15176);
or U18716 (N_18716,N_16539,N_17688);
nor U18717 (N_18717,N_15790,N_16423);
xnor U18718 (N_18718,N_16784,N_15869);
xor U18719 (N_18719,N_17123,N_16044);
and U18720 (N_18720,N_15625,N_15672);
nand U18721 (N_18721,N_16860,N_15678);
nor U18722 (N_18722,N_15377,N_17269);
nand U18723 (N_18723,N_16616,N_16347);
or U18724 (N_18724,N_16436,N_17225);
and U18725 (N_18725,N_17023,N_16235);
or U18726 (N_18726,N_17609,N_15608);
xnor U18727 (N_18727,N_17310,N_16879);
nand U18728 (N_18728,N_16953,N_17600);
xor U18729 (N_18729,N_16584,N_17674);
xnor U18730 (N_18730,N_15140,N_16800);
xnor U18731 (N_18731,N_17247,N_16702);
nor U18732 (N_18732,N_15156,N_16197);
and U18733 (N_18733,N_15595,N_17110);
xor U18734 (N_18734,N_15169,N_15565);
xor U18735 (N_18735,N_17842,N_17797);
nor U18736 (N_18736,N_17255,N_17525);
or U18737 (N_18737,N_17546,N_17729);
nor U18738 (N_18738,N_15585,N_17312);
and U18739 (N_18739,N_15920,N_16766);
or U18740 (N_18740,N_17372,N_17271);
and U18741 (N_18741,N_16603,N_17763);
nand U18742 (N_18742,N_16144,N_17605);
or U18743 (N_18743,N_15757,N_17671);
nor U18744 (N_18744,N_16671,N_15800);
nor U18745 (N_18745,N_16024,N_17221);
and U18746 (N_18746,N_15481,N_16218);
nor U18747 (N_18747,N_17529,N_15149);
nor U18748 (N_18748,N_15662,N_16754);
or U18749 (N_18749,N_16477,N_16354);
and U18750 (N_18750,N_16338,N_17216);
nor U18751 (N_18751,N_16920,N_15751);
and U18752 (N_18752,N_15366,N_15649);
nor U18753 (N_18753,N_15085,N_16690);
or U18754 (N_18754,N_15897,N_17026);
or U18755 (N_18755,N_16428,N_17879);
and U18756 (N_18756,N_15648,N_17384);
and U18757 (N_18757,N_15515,N_15088);
xor U18758 (N_18758,N_17278,N_17669);
nor U18759 (N_18759,N_16045,N_16900);
nor U18760 (N_18760,N_15026,N_16820);
nand U18761 (N_18761,N_17030,N_15776);
or U18762 (N_18762,N_17004,N_15094);
or U18763 (N_18763,N_16072,N_17487);
nand U18764 (N_18764,N_15384,N_17803);
nand U18765 (N_18765,N_16871,N_15986);
nand U18766 (N_18766,N_17703,N_17604);
and U18767 (N_18767,N_17042,N_16700);
nand U18768 (N_18768,N_15715,N_15211);
xor U18769 (N_18769,N_15219,N_15949);
nand U18770 (N_18770,N_17239,N_17172);
nor U18771 (N_18771,N_17952,N_15027);
xor U18772 (N_18772,N_16506,N_16316);
and U18773 (N_18773,N_16565,N_15966);
nand U18774 (N_18774,N_17827,N_17625);
and U18775 (N_18775,N_15052,N_17982);
nor U18776 (N_18776,N_17396,N_17252);
nor U18777 (N_18777,N_17782,N_16198);
or U18778 (N_18778,N_17402,N_16387);
nor U18779 (N_18779,N_15421,N_16512);
and U18780 (N_18780,N_16685,N_16684);
or U18781 (N_18781,N_17824,N_15935);
nand U18782 (N_18782,N_17062,N_17985);
nand U18783 (N_18783,N_17538,N_16313);
or U18784 (N_18784,N_15590,N_15763);
nor U18785 (N_18785,N_17843,N_17918);
nand U18786 (N_18786,N_17713,N_15861);
xnor U18787 (N_18787,N_16760,N_16150);
nand U18788 (N_18788,N_17434,N_15500);
nand U18789 (N_18789,N_16647,N_17559);
nand U18790 (N_18790,N_16776,N_15930);
nor U18791 (N_18791,N_16037,N_16468);
nand U18792 (N_18792,N_15049,N_15434);
and U18793 (N_18793,N_17871,N_16178);
nor U18794 (N_18794,N_15106,N_15611);
or U18795 (N_18795,N_17391,N_17654);
nand U18796 (N_18796,N_15245,N_17667);
or U18797 (N_18797,N_17793,N_15823);
or U18798 (N_18798,N_15381,N_15490);
or U18799 (N_18799,N_17971,N_17704);
nand U18800 (N_18800,N_15387,N_15129);
and U18801 (N_18801,N_17829,N_15557);
xor U18802 (N_18802,N_15987,N_15294);
nand U18803 (N_18803,N_17788,N_15264);
or U18804 (N_18804,N_16798,N_16574);
nand U18805 (N_18805,N_17627,N_17069);
xnor U18806 (N_18806,N_17710,N_17186);
xnor U18807 (N_18807,N_15891,N_15548);
xor U18808 (N_18808,N_16556,N_16563);
nor U18809 (N_18809,N_17895,N_17150);
or U18810 (N_18810,N_15437,N_17045);
or U18811 (N_18811,N_17602,N_15042);
nand U18812 (N_18812,N_17491,N_16673);
xnor U18813 (N_18813,N_17953,N_15717);
nor U18814 (N_18814,N_16424,N_17999);
nor U18815 (N_18815,N_17408,N_16913);
xnor U18816 (N_18816,N_17992,N_17101);
nor U18817 (N_18817,N_15141,N_15331);
xor U18818 (N_18818,N_15332,N_16470);
nor U18819 (N_18819,N_16120,N_17980);
xnor U18820 (N_18820,N_16835,N_17068);
nor U18821 (N_18821,N_16333,N_15913);
xnor U18822 (N_18822,N_15546,N_15227);
xnor U18823 (N_18823,N_16892,N_15842);
and U18824 (N_18824,N_17778,N_15322);
or U18825 (N_18825,N_17404,N_15110);
nor U18826 (N_18826,N_17723,N_17222);
and U18827 (N_18827,N_15359,N_17063);
nor U18828 (N_18828,N_16993,N_16006);
or U18829 (N_18829,N_16378,N_15575);
and U18830 (N_18830,N_16759,N_15312);
nor U18831 (N_18831,N_16260,N_15874);
nand U18832 (N_18832,N_17846,N_15864);
and U18833 (N_18833,N_15675,N_15151);
nand U18834 (N_18834,N_15851,N_15193);
xnor U18835 (N_18835,N_16761,N_16611);
nand U18836 (N_18836,N_17816,N_17875);
or U18837 (N_18837,N_15730,N_17946);
nand U18838 (N_18838,N_15067,N_16337);
nor U18839 (N_18839,N_16236,N_15704);
and U18840 (N_18840,N_17163,N_16816);
or U18841 (N_18841,N_15732,N_17737);
nand U18842 (N_18842,N_17496,N_17291);
or U18843 (N_18843,N_17683,N_15096);
or U18844 (N_18844,N_16525,N_16517);
nand U18845 (N_18845,N_17811,N_16648);
or U18846 (N_18846,N_16269,N_17553);
xnor U18847 (N_18847,N_15337,N_15095);
or U18848 (N_18848,N_15065,N_15248);
and U18849 (N_18849,N_16617,N_17579);
or U18850 (N_18850,N_17477,N_17091);
and U18851 (N_18851,N_15339,N_16256);
nand U18852 (N_18852,N_15484,N_16594);
nor U18853 (N_18853,N_17880,N_16206);
nor U18854 (N_18854,N_17336,N_15810);
and U18855 (N_18855,N_15531,N_15442);
nor U18856 (N_18856,N_16634,N_16229);
nand U18857 (N_18857,N_16223,N_16559);
nand U18858 (N_18858,N_17612,N_17576);
nand U18859 (N_18859,N_15007,N_17073);
xnor U18860 (N_18860,N_15479,N_17861);
nand U18861 (N_18861,N_17345,N_15744);
nand U18862 (N_18862,N_16390,N_15902);
and U18863 (N_18863,N_17818,N_17590);
and U18864 (N_18864,N_15086,N_15116);
xor U18865 (N_18865,N_15168,N_17027);
or U18866 (N_18866,N_15679,N_17613);
or U18867 (N_18867,N_17940,N_15961);
nor U18868 (N_18868,N_17960,N_16533);
and U18869 (N_18869,N_15684,N_17639);
nor U18870 (N_18870,N_15160,N_17942);
xnor U18871 (N_18871,N_16214,N_17422);
or U18872 (N_18872,N_17297,N_16922);
xnor U18873 (N_18873,N_16088,N_17324);
xnor U18874 (N_18874,N_15389,N_16067);
and U18875 (N_18875,N_17235,N_15849);
xor U18876 (N_18876,N_16427,N_15196);
or U18877 (N_18877,N_15150,N_17866);
or U18878 (N_18878,N_16987,N_16293);
nand U18879 (N_18879,N_17757,N_16482);
xnor U18880 (N_18880,N_16020,N_15130);
nand U18881 (N_18881,N_17858,N_16914);
nor U18882 (N_18882,N_17087,N_16558);
nand U18883 (N_18883,N_16686,N_15252);
or U18884 (N_18884,N_15032,N_17292);
and U18885 (N_18885,N_17180,N_17658);
and U18886 (N_18886,N_15293,N_17930);
nand U18887 (N_18887,N_15262,N_16419);
nand U18888 (N_18888,N_15412,N_16358);
xnor U18889 (N_18889,N_16978,N_17923);
xnor U18890 (N_18890,N_17572,N_15038);
xor U18891 (N_18891,N_17644,N_17203);
and U18892 (N_18892,N_17059,N_15906);
nor U18893 (N_18893,N_17298,N_16967);
xnor U18894 (N_18894,N_17119,N_17416);
xor U18895 (N_18895,N_15441,N_15103);
nor U18896 (N_18896,N_17394,N_15091);
and U18897 (N_18897,N_15314,N_15401);
xnor U18898 (N_18898,N_15576,N_17614);
and U18899 (N_18899,N_15158,N_17571);
and U18900 (N_18900,N_15879,N_17238);
xnor U18901 (N_18901,N_16352,N_17791);
and U18902 (N_18902,N_15418,N_16444);
and U18903 (N_18903,N_16283,N_17395);
xor U18904 (N_18904,N_16130,N_15020);
or U18905 (N_18905,N_17167,N_15885);
or U18906 (N_18906,N_17835,N_15269);
or U18907 (N_18907,N_17451,N_16984);
or U18908 (N_18908,N_15784,N_16949);
or U18909 (N_18909,N_17322,N_16410);
and U18910 (N_18910,N_16194,N_15444);
or U18911 (N_18911,N_16992,N_16626);
xor U18912 (N_18912,N_16098,N_17418);
xor U18913 (N_18913,N_17752,N_15235);
and U18914 (N_18914,N_16003,N_17012);
or U18915 (N_18915,N_16587,N_17003);
xor U18916 (N_18916,N_16755,N_15316);
or U18917 (N_18917,N_17586,N_16265);
or U18918 (N_18918,N_15579,N_16857);
or U18919 (N_18919,N_16491,N_15513);
nand U18920 (N_18920,N_16078,N_17041);
nand U18921 (N_18921,N_15905,N_16505);
or U18922 (N_18922,N_16315,N_16662);
xnor U18923 (N_18923,N_16705,N_15487);
nand U18924 (N_18924,N_16572,N_16193);
nand U18925 (N_18925,N_16246,N_16021);
nor U18926 (N_18926,N_15782,N_16698);
nand U18927 (N_18927,N_15115,N_17695);
or U18928 (N_18928,N_16711,N_16722);
and U18929 (N_18929,N_16305,N_15003);
or U18930 (N_18930,N_15162,N_15098);
nand U18931 (N_18931,N_17628,N_16373);
nand U18932 (N_18932,N_16752,N_15826);
nor U18933 (N_18933,N_16251,N_16409);
xnor U18934 (N_18934,N_16808,N_16657);
and U18935 (N_18935,N_17838,N_17081);
xnor U18936 (N_18936,N_15876,N_15747);
and U18937 (N_18937,N_15013,N_17524);
or U18938 (N_18938,N_17237,N_17352);
nor U18939 (N_18939,N_16475,N_16296);
and U18940 (N_18940,N_15299,N_16507);
or U18941 (N_18941,N_15701,N_16665);
or U18942 (N_18942,N_17294,N_17000);
nand U18943 (N_18943,N_17488,N_17264);
or U18944 (N_18944,N_16699,N_17460);
nor U18945 (N_18945,N_16361,N_16708);
nor U18946 (N_18946,N_16403,N_16915);
and U18947 (N_18947,N_17469,N_16121);
or U18948 (N_18948,N_17906,N_15718);
nor U18949 (N_18949,N_16585,N_15008);
xnor U18950 (N_18950,N_16060,N_17724);
nor U18951 (N_18951,N_17057,N_16724);
xnor U18952 (N_18952,N_16866,N_16786);
nand U18953 (N_18953,N_17938,N_15709);
xnor U18954 (N_18954,N_17128,N_16059);
xor U18955 (N_18955,N_15069,N_17382);
nor U18956 (N_18956,N_16418,N_17311);
and U18957 (N_18957,N_16281,N_15355);
and U18958 (N_18958,N_15451,N_16604);
xnor U18959 (N_18959,N_17184,N_15788);
or U18960 (N_18960,N_17428,N_16070);
or U18961 (N_18961,N_15738,N_16312);
nand U18962 (N_18962,N_16694,N_16168);
or U18963 (N_18963,N_15155,N_16649);
or U18964 (N_18964,N_15233,N_16398);
xor U18965 (N_18965,N_15157,N_15558);
nor U18966 (N_18966,N_16522,N_16511);
nand U18967 (N_18967,N_16368,N_17233);
and U18968 (N_18968,N_15604,N_17780);
and U18969 (N_18969,N_16793,N_16552);
xnor U18970 (N_18970,N_16286,N_17175);
xor U18971 (N_18971,N_17776,N_17928);
and U18972 (N_18972,N_17074,N_16832);
xnor U18973 (N_18973,N_16838,N_15774);
xor U18974 (N_18974,N_17694,N_16076);
or U18975 (N_18975,N_17720,N_16056);
nand U18976 (N_18976,N_15495,N_16435);
or U18977 (N_18977,N_16498,N_16593);
or U18978 (N_18978,N_16189,N_17717);
and U18979 (N_18979,N_17162,N_15660);
nor U18980 (N_18980,N_17260,N_15108);
and U18981 (N_18981,N_17741,N_17381);
nor U18982 (N_18982,N_16582,N_17463);
and U18983 (N_18983,N_17641,N_15544);
xor U18984 (N_18984,N_17642,N_16948);
xnor U18985 (N_18985,N_17666,N_17333);
or U18986 (N_18986,N_17826,N_17770);
nor U18987 (N_18987,N_17792,N_17779);
xor U18988 (N_18988,N_15295,N_17176);
and U18989 (N_18989,N_15347,N_16529);
nor U18990 (N_18990,N_16547,N_17786);
xnor U18991 (N_18991,N_16417,N_16402);
nand U18992 (N_18992,N_16127,N_16628);
or U18993 (N_18993,N_17870,N_17697);
and U18994 (N_18994,N_17218,N_16216);
xor U18995 (N_18995,N_17457,N_17154);
xnor U18996 (N_18996,N_17151,N_15630);
nor U18997 (N_18997,N_17219,N_17262);
and U18998 (N_18998,N_15147,N_16897);
nor U18999 (N_18999,N_17629,N_16103);
nor U19000 (N_19000,N_17164,N_15963);
and U19001 (N_19001,N_16446,N_15659);
xnor U19002 (N_19002,N_17635,N_17055);
nand U19003 (N_19003,N_16643,N_16301);
nand U19004 (N_19004,N_17369,N_16367);
and U19005 (N_19005,N_16810,N_17997);
nand U19006 (N_19006,N_15911,N_17511);
or U19007 (N_19007,N_17839,N_17555);
nor U19008 (N_19008,N_16555,N_17273);
and U19009 (N_19009,N_17986,N_17742);
xor U19010 (N_19010,N_15409,N_16792);
nand U19011 (N_19011,N_16943,N_17043);
or U19012 (N_19012,N_16249,N_15657);
nand U19013 (N_19013,N_15620,N_15062);
and U19014 (N_19014,N_17240,N_15180);
nor U19015 (N_19015,N_17309,N_17499);
or U19016 (N_19016,N_16619,N_17787);
and U19017 (N_19017,N_15338,N_17652);
xnor U19018 (N_19018,N_15396,N_17283);
and U19019 (N_19019,N_16308,N_17831);
xnor U19020 (N_19020,N_16126,N_15329);
or U19021 (N_19021,N_17208,N_16230);
nand U19022 (N_19022,N_16245,N_17593);
nand U19023 (N_19023,N_16613,N_15532);
nand U19024 (N_19024,N_16641,N_15203);
nand U19025 (N_19025,N_17009,N_15741);
nand U19026 (N_19026,N_17132,N_17380);
xor U19027 (N_19027,N_16770,N_15040);
nand U19028 (N_19028,N_16017,N_17227);
nor U19029 (N_19029,N_15962,N_16159);
and U19030 (N_19030,N_16205,N_16856);
or U19031 (N_19031,N_16687,N_16405);
nand U19032 (N_19032,N_17173,N_15586);
nand U19033 (N_19033,N_15424,N_17244);
and U19034 (N_19034,N_16136,N_16314);
or U19035 (N_19035,N_16524,N_17712);
nor U19036 (N_19036,N_17500,N_17775);
nand U19037 (N_19037,N_15983,N_17626);
or U19038 (N_19038,N_16716,N_16287);
nor U19039 (N_19039,N_16357,N_17486);
or U19040 (N_19040,N_16629,N_15795);
nand U19041 (N_19041,N_17267,N_15132);
nor U19042 (N_19042,N_17708,N_17749);
and U19043 (N_19043,N_17860,N_16053);
or U19044 (N_19044,N_17771,N_17958);
xor U19045 (N_19045,N_15812,N_15888);
nand U19046 (N_19046,N_17254,N_16549);
nand U19047 (N_19047,N_15871,N_17047);
xor U19048 (N_19048,N_17410,N_15817);
xnor U19049 (N_19049,N_17371,N_16621);
xnor U19050 (N_19050,N_16031,N_17727);
or U19051 (N_19051,N_15834,N_15785);
and U19052 (N_19052,N_16650,N_15057);
nor U19053 (N_19053,N_15799,N_17455);
or U19054 (N_19054,N_15324,N_16706);
nand U19055 (N_19055,N_15942,N_15806);
or U19056 (N_19056,N_16268,N_17934);
xnor U19057 (N_19057,N_16730,N_17118);
or U19058 (N_19058,N_16186,N_17504);
nand U19059 (N_19059,N_17102,N_15764);
and U19060 (N_19060,N_17389,N_16847);
xor U19061 (N_19061,N_17470,N_16803);
xnor U19062 (N_19062,N_16493,N_17808);
or U19063 (N_19063,N_16473,N_15598);
nor U19064 (N_19064,N_17293,N_16467);
and U19065 (N_19065,N_15988,N_17907);
nand U19066 (N_19066,N_16868,N_15012);
or U19067 (N_19067,N_17801,N_16181);
xor U19068 (N_19068,N_17607,N_17756);
or U19069 (N_19069,N_17615,N_17796);
and U19070 (N_19070,N_15768,N_16560);
and U19071 (N_19071,N_16719,N_16365);
xor U19072 (N_19072,N_15344,N_15485);
nor U19073 (N_19073,N_15989,N_17053);
nand U19074 (N_19074,N_16735,N_16853);
and U19075 (N_19075,N_16733,N_15154);
and U19076 (N_19076,N_15139,N_17332);
or U19077 (N_19077,N_15521,N_16397);
xor U19078 (N_19078,N_17152,N_17949);
or U19079 (N_19079,N_15253,N_15178);
and U19080 (N_19080,N_16461,N_17592);
nor U19081 (N_19081,N_17268,N_17728);
and U19082 (N_19082,N_16674,N_16259);
nor U19083 (N_19083,N_15267,N_16797);
nand U19084 (N_19084,N_16812,N_17815);
xnor U19085 (N_19085,N_16721,N_15943);
or U19086 (N_19086,N_17093,N_16758);
xnor U19087 (N_19087,N_17821,N_17582);
or U19088 (N_19088,N_15240,N_15700);
nor U19089 (N_19089,N_16146,N_16257);
or U19090 (N_19090,N_16562,N_17275);
and U19091 (N_19091,N_17122,N_17790);
and U19092 (N_19092,N_15087,N_15113);
or U19093 (N_19093,N_15922,N_15317);
nand U19094 (N_19094,N_16016,N_17508);
or U19095 (N_19095,N_15820,N_17715);
nor U19096 (N_19096,N_16743,N_17964);
nand U19097 (N_19097,N_17245,N_16689);
nand U19098 (N_19098,N_16697,N_15079);
or U19099 (N_19099,N_16479,N_16474);
and U19100 (N_19100,N_15489,N_16515);
nand U19101 (N_19101,N_15731,N_15281);
nor U19102 (N_19102,N_17904,N_16004);
or U19103 (N_19103,N_16564,N_15689);
nand U19104 (N_19104,N_16501,N_17231);
or U19105 (N_19105,N_16495,N_17805);
nand U19106 (N_19106,N_17698,N_16997);
and U19107 (N_19107,N_17848,N_17929);
and U19108 (N_19108,N_15394,N_15014);
and U19109 (N_19109,N_16894,N_15285);
nand U19110 (N_19110,N_16371,N_17076);
and U19111 (N_19111,N_17157,N_15454);
or U19112 (N_19112,N_17299,N_17234);
and U19113 (N_19113,N_15433,N_17539);
and U19114 (N_19114,N_17968,N_16290);
xnor U19115 (N_19115,N_15699,N_17685);
and U19116 (N_19116,N_15438,N_17885);
nand U19117 (N_19117,N_17185,N_15493);
nor U19118 (N_19118,N_15256,N_15364);
nor U19119 (N_19119,N_15362,N_15111);
nand U19120 (N_19120,N_15142,N_16837);
nor U19121 (N_19121,N_17362,N_15815);
and U19122 (N_19122,N_15469,N_15644);
nor U19123 (N_19123,N_17994,N_15848);
xnor U19124 (N_19124,N_17113,N_17761);
nand U19125 (N_19125,N_16775,N_17956);
xnor U19126 (N_19126,N_17096,N_17595);
nor U19127 (N_19127,N_15803,N_15216);
nor U19128 (N_19128,N_17864,N_17339);
nand U19129 (N_19129,N_17884,N_16580);
nand U19130 (N_19130,N_16149,N_15152);
nor U19131 (N_19131,N_17996,N_15938);
or U19132 (N_19132,N_15537,N_15373);
xor U19133 (N_19133,N_17781,N_17415);
or U19134 (N_19134,N_17814,N_17436);
xor U19135 (N_19135,N_16292,N_16590);
or U19136 (N_19136,N_16930,N_17509);
nand U19137 (N_19137,N_15573,N_16094);
xnor U19138 (N_19138,N_17147,N_16091);
nand U19139 (N_19139,N_15780,N_15137);
nor U19140 (N_19140,N_16849,N_15214);
or U19141 (N_19141,N_15406,N_16575);
and U19142 (N_19142,N_15340,N_16183);
and U19143 (N_19143,N_15605,N_16878);
or U19144 (N_19144,N_17405,N_16469);
nor U19145 (N_19145,N_16480,N_17459);
and U19146 (N_19146,N_17259,N_15705);
nand U19147 (N_19147,N_16187,N_16464);
and U19148 (N_19148,N_16135,N_15035);
nor U19149 (N_19149,N_16100,N_15814);
or U19150 (N_19150,N_15733,N_15276);
or U19151 (N_19151,N_15601,N_16297);
nand U19152 (N_19152,N_15061,N_17307);
and U19153 (N_19153,N_16782,N_15921);
nor U19154 (N_19154,N_15480,N_16910);
or U19155 (N_19155,N_16431,N_16112);
nor U19156 (N_19156,N_16052,N_16519);
and U19157 (N_19157,N_16115,N_16833);
nand U19158 (N_19158,N_15967,N_16964);
and U19159 (N_19159,N_17892,N_16369);
xor U19160 (N_19160,N_17002,N_17975);
nor U19161 (N_19161,N_17965,N_16154);
and U19162 (N_19162,N_17901,N_16114);
or U19163 (N_19163,N_15242,N_16666);
or U19164 (N_19164,N_16592,N_15992);
xnor U19165 (N_19165,N_15641,N_15981);
xor U19166 (N_19166,N_15635,N_17124);
nor U19167 (N_19167,N_16095,N_16317);
nand U19168 (N_19168,N_15300,N_15976);
xnor U19169 (N_19169,N_15346,N_15519);
and U19170 (N_19170,N_17651,N_15369);
nor U19171 (N_19171,N_17424,N_15652);
or U19172 (N_19172,N_15501,N_17978);
nor U19173 (N_19173,N_17033,N_16632);
or U19174 (N_19174,N_17282,N_17338);
or U19175 (N_19175,N_15547,N_15112);
nor U19176 (N_19176,N_17507,N_17148);
xor U19177 (N_19177,N_15195,N_16068);
and U19178 (N_19178,N_16550,N_15884);
or U19179 (N_19179,N_15230,N_17040);
or U19180 (N_19180,N_16824,N_17514);
xnor U19181 (N_19181,N_17194,N_16393);
xnor U19182 (N_19182,N_17116,N_17419);
or U19183 (N_19183,N_15220,N_16231);
and U19184 (N_19184,N_17192,N_16640);
or U19185 (N_19185,N_16834,N_16166);
nand U19186 (N_19186,N_15353,N_16233);
xnor U19187 (N_19187,N_17549,N_17810);
and U19188 (N_19188,N_15698,N_17099);
xnor U19189 (N_19189,N_16463,N_17959);
xnor U19190 (N_19190,N_17963,N_15173);
or U19191 (N_19191,N_17680,N_15890);
and U19192 (N_19192,N_15969,N_15783);
nand U19193 (N_19193,N_16481,N_15507);
nor U19194 (N_19194,N_17774,N_17479);
and U19195 (N_19195,N_15232,N_17242);
xor U19196 (N_19196,N_17494,N_17589);
nand U19197 (N_19197,N_16033,N_17359);
and U19198 (N_19198,N_16339,N_16532);
xor U19199 (N_19199,N_17819,N_16389);
xnor U19200 (N_19200,N_15588,N_15683);
or U19201 (N_19201,N_16823,N_15687);
nor U19202 (N_19202,N_17168,N_17089);
nor U19203 (N_19203,N_15654,N_15899);
nor U19204 (N_19204,N_17730,N_15268);
nor U19205 (N_19205,N_17886,N_17764);
nand U19206 (N_19206,N_15753,N_15643);
xnor U19207 (N_19207,N_17665,N_15217);
nand U19208 (N_19208,N_17353,N_17049);
or U19209 (N_19209,N_15778,N_17565);
or U19210 (N_19210,N_15716,N_17515);
nor U19211 (N_19211,N_15996,N_15505);
or U19212 (N_19212,N_15686,N_17144);
or U19213 (N_19213,N_15255,N_16874);
and U19214 (N_19214,N_17355,N_17276);
and U19215 (N_19215,N_15194,N_17535);
or U19216 (N_19216,N_15646,N_17025);
and U19217 (N_19217,N_16971,N_17948);
and U19218 (N_19218,N_15462,N_15807);
nor U19219 (N_19219,N_15126,N_17288);
xnor U19220 (N_19220,N_16888,N_15287);
xor U19221 (N_19221,N_16955,N_15514);
or U19222 (N_19222,N_16000,N_15213);
nand U19223 (N_19223,N_16952,N_15127);
and U19224 (N_19224,N_15846,N_17725);
nand U19225 (N_19225,N_15472,N_16349);
and U19226 (N_19226,N_17050,N_15956);
xnor U19227 (N_19227,N_17029,N_16638);
and U19228 (N_19228,N_15349,N_17921);
or U19229 (N_19229,N_16741,N_15144);
or U19230 (N_19230,N_17517,N_16998);
or U19231 (N_19231,N_15769,N_17691);
xor U19232 (N_19232,N_17401,N_15416);
and U19233 (N_19233,N_16160,N_15025);
or U19234 (N_19234,N_17550,N_17274);
nand U19235 (N_19235,N_17377,N_15104);
and U19236 (N_19236,N_17966,N_16609);
or U19237 (N_19237,N_17433,N_16789);
or U19238 (N_19238,N_15029,N_17939);
and U19239 (N_19239,N_17649,N_16753);
xnor U19240 (N_19240,N_16174,N_16845);
xor U19241 (N_19241,N_17908,N_15361);
nor U19242 (N_19242,N_15348,N_15628);
or U19243 (N_19243,N_15328,N_16933);
xnor U19244 (N_19244,N_15499,N_16010);
nand U19245 (N_19245,N_16104,N_16830);
and U19246 (N_19246,N_17903,N_15077);
xnor U19247 (N_19247,N_16597,N_15251);
nor U19248 (N_19248,N_17983,N_15435);
xnor U19249 (N_19249,N_16032,N_17998);
nor U19250 (N_19250,N_17893,N_17611);
nor U19251 (N_19251,N_17126,N_15589);
xnor U19252 (N_19252,N_15372,N_16744);
or U19253 (N_19253,N_16877,N_16342);
and U19254 (N_19254,N_15404,N_15664);
nor U19255 (N_19255,N_16510,N_16976);
and U19256 (N_19256,N_16731,N_15793);
nand U19257 (N_19257,N_16452,N_17910);
xnor U19258 (N_19258,N_16232,N_16742);
nand U19259 (N_19259,N_16573,N_16400);
or U19260 (N_19260,N_15900,N_16692);
nand U19261 (N_19261,N_15602,N_16545);
xnor U19262 (N_19262,N_17092,N_15136);
nand U19263 (N_19263,N_16304,N_16124);
nand U19264 (N_19264,N_15081,N_17313);
and U19265 (N_19265,N_15656,N_15273);
xnor U19266 (N_19266,N_16344,N_16156);
and U19267 (N_19267,N_15552,N_16376);
xnor U19268 (N_19268,N_15183,N_16683);
or U19269 (N_19269,N_17086,N_17136);
nand U19270 (N_19270,N_17863,N_15165);
nand U19271 (N_19271,N_17034,N_16111);
and U19272 (N_19272,N_17594,N_15592);
nor U19273 (N_19273,N_16190,N_16548);
nor U19274 (N_19274,N_17358,N_16458);
or U19275 (N_19275,N_17127,N_16513);
nor U19276 (N_19276,N_16644,N_15284);
xnor U19277 (N_19277,N_16240,N_16757);
nor U19278 (N_19278,N_17569,N_16438);
and U19279 (N_19279,N_15564,N_15371);
nand U19280 (N_19280,N_16379,N_15692);
xor U19281 (N_19281,N_15617,N_17679);
or U19282 (N_19282,N_17170,N_15405);
xor U19283 (N_19283,N_17643,N_16937);
or U19284 (N_19284,N_15124,N_16209);
xor U19285 (N_19285,N_17616,N_15456);
nor U19286 (N_19286,N_15432,N_17423);
and U19287 (N_19287,N_17648,N_15714);
or U19288 (N_19288,N_15231,N_16440);
nand U19289 (N_19289,N_15254,N_16380);
or U19290 (N_19290,N_15483,N_15445);
nor U19291 (N_19291,N_17554,N_17114);
xnor U19292 (N_19292,N_17449,N_16346);
or U19293 (N_19293,N_16710,N_15325);
and U19294 (N_19294,N_17376,N_15167);
nor U19295 (N_19295,N_16163,N_15302);
xnor U19296 (N_19296,N_17217,N_17617);
and U19297 (N_19297,N_16822,N_17869);
nor U19298 (N_19298,N_15226,N_15638);
nand U19299 (N_19299,N_17933,N_15550);
and U19300 (N_19300,N_16038,N_16636);
or U19301 (N_19301,N_15985,N_15551);
nor U19302 (N_19302,N_16234,N_17197);
and U19303 (N_19303,N_15166,N_17452);
xor U19304 (N_19304,N_15901,N_16720);
or U19305 (N_19305,N_17481,N_16204);
nor U19306 (N_19306,N_17972,N_16029);
xor U19307 (N_19307,N_17977,N_16869);
nand U19308 (N_19308,N_16085,N_16153);
nor U19309 (N_19309,N_15908,N_15838);
or U19310 (N_19310,N_17783,N_15965);
and U19311 (N_19311,N_15258,N_15755);
xnor U19312 (N_19312,N_17993,N_17006);
nand U19313 (N_19313,N_17109,N_15074);
xnor U19314 (N_19314,N_16990,N_15189);
or U19315 (N_19315,N_16258,N_17061);
nand U19316 (N_19316,N_16867,N_15315);
and U19317 (N_19317,N_16663,N_16081);
nand U19318 (N_19318,N_16140,N_16170);
and U19319 (N_19319,N_15593,N_17743);
nor U19320 (N_19320,N_15581,N_15280);
or U19321 (N_19321,N_15274,N_17503);
xnor U19322 (N_19322,N_15697,N_16895);
nand U19323 (N_19323,N_17320,N_17108);
xnor U19324 (N_19324,N_15596,N_17789);
or U19325 (N_19325,N_17131,N_15837);
or U19326 (N_19326,N_17825,N_16139);
xor U19327 (N_19327,N_15460,N_16008);
or U19328 (N_19328,N_17917,N_17214);
and U19329 (N_19329,N_16099,N_15749);
nand U19330 (N_19330,N_17085,N_17077);
nand U19331 (N_19331,N_15621,N_15464);
or U19332 (N_19332,N_17472,N_17105);
and U19333 (N_19333,N_17437,N_16912);
nor U19334 (N_19334,N_16324,N_17558);
xnor U19335 (N_19335,N_15973,N_15024);
or U19336 (N_19336,N_16299,N_15534);
xnor U19337 (N_19337,N_15288,N_15224);
and U19338 (N_19338,N_16089,N_17224);
and U19339 (N_19339,N_17812,N_17681);
xor U19340 (N_19340,N_15350,N_16034);
and U19341 (N_19341,N_17344,N_17257);
and U19342 (N_19342,N_15612,N_15471);
xnor U19343 (N_19343,N_15526,N_15304);
nand U19344 (N_19344,N_15696,N_16509);
or U19345 (N_19345,N_16723,N_17474);
nand U19346 (N_19346,N_17766,N_17706);
or U19347 (N_19347,N_17097,N_17388);
or U19348 (N_19348,N_15218,N_15386);
nand U19349 (N_19349,N_16859,N_16740);
xnor U19350 (N_19350,N_16669,N_16679);
xor U19351 (N_19351,N_17476,N_16787);
xor U19352 (N_19352,N_16018,N_17497);
and U19353 (N_19353,N_17753,N_16028);
nor U19354 (N_19354,N_15201,N_15835);
nor U19355 (N_19355,N_16429,N_17125);
xor U19356 (N_19356,N_17229,N_16848);
nor U19357 (N_19357,N_15570,N_16934);
nor U19358 (N_19358,N_16182,N_15310);
nor U19359 (N_19359,N_16890,N_17417);
and U19360 (N_19360,N_15382,N_17520);
xnor U19361 (N_19361,N_17326,N_15502);
nor U19362 (N_19362,N_16485,N_17527);
xor U19363 (N_19363,N_15545,N_17765);
and U19364 (N_19364,N_16995,N_17544);
nor U19365 (N_19365,N_17232,N_16152);
nand U19366 (N_19366,N_17833,N_17327);
xnor U19367 (N_19367,N_16728,N_15779);
nor U19368 (N_19368,N_16695,N_16809);
xnor U19369 (N_19369,N_17155,N_17129);
xnor U19370 (N_19370,N_16521,N_16651);
xnor U19371 (N_19371,N_17970,N_17813);
or U19372 (N_19372,N_16323,N_15873);
nor U19373 (N_19373,N_17621,N_16598);
xor U19374 (N_19374,N_16970,N_17567);
xor U19375 (N_19375,N_15914,N_16080);
nor U19376 (N_19376,N_15046,N_17830);
xnor U19377 (N_19377,N_16105,N_15174);
or U19378 (N_19378,N_15616,N_16051);
nand U19379 (N_19379,N_16825,N_16736);
xnor U19380 (N_19380,N_16778,N_16554);
nor U19381 (N_19381,N_16578,N_17905);
and U19382 (N_19382,N_17478,N_15450);
xnor U19383 (N_19383,N_15039,N_15655);
nor U19384 (N_19384,N_15058,N_15640);
xor U19385 (N_19385,N_15841,N_16932);
nand U19386 (N_19386,N_15429,N_15610);
xnor U19387 (N_19387,N_15102,N_17799);
or U19388 (N_19388,N_15503,N_15023);
xnor U19389 (N_19389,N_16023,N_15607);
or U19390 (N_19390,N_15762,N_16954);
nand U19391 (N_19391,N_16625,N_17719);
nor U19392 (N_19392,N_17331,N_17195);
and U19393 (N_19393,N_15673,N_16219);
nor U19394 (N_19394,N_17318,N_15772);
or U19395 (N_19395,N_17236,N_16917);
and U19396 (N_19396,N_16977,N_17133);
or U19397 (N_19397,N_16175,N_15187);
nand U19398 (N_19398,N_16366,N_16248);
and U19399 (N_19399,N_17256,N_17466);
nor U19400 (N_19400,N_15991,N_15036);
nor U19401 (N_19401,N_15131,N_15383);
or U19402 (N_19402,N_15080,N_15283);
and U19403 (N_19403,N_15623,N_16220);
or U19404 (N_19404,N_16030,N_17518);
xnor U19405 (N_19405,N_15866,N_17522);
and U19406 (N_19406,N_16065,N_16646);
and U19407 (N_19407,N_17453,N_16846);
xnor U19408 (N_19408,N_16691,N_17253);
nand U19409 (N_19409,N_15275,N_16042);
or U19410 (N_19410,N_17662,N_16241);
and U19411 (N_19411,N_16956,N_15246);
or U19412 (N_19412,N_16655,N_17067);
xnor U19413 (N_19413,N_16125,N_17432);
nor U19414 (N_19414,N_17080,N_16086);
nor U19415 (N_19415,N_15497,N_17181);
nor U19416 (N_19416,N_17562,N_15609);
nor U19417 (N_19417,N_16982,N_16576);
nand U19418 (N_19418,N_17686,N_16141);
nand U19419 (N_19419,N_17039,N_15517);
and U19420 (N_19420,N_15528,N_15375);
nand U19421 (N_19421,N_16453,N_16007);
and U19422 (N_19422,N_17575,N_15615);
xnor U19423 (N_19423,N_17301,N_17640);
nor U19424 (N_19424,N_15290,N_15636);
nand U19425 (N_19425,N_16015,N_17889);
and U19426 (N_19426,N_17153,N_16264);
nand U19427 (N_19427,N_16392,N_17046);
and U19428 (N_19428,N_15099,N_15743);
nor U19429 (N_19429,N_17647,N_16096);
nand U19430 (N_19430,N_16199,N_15568);
nor U19431 (N_19431,N_15419,N_15427);
or U19432 (N_19432,N_17346,N_15622);
or U19433 (N_19433,N_17751,N_16896);
nor U19434 (N_19434,N_15653,N_17329);
and U19435 (N_19435,N_17279,N_17342);
or U19436 (N_19436,N_16806,N_17335);
nor U19437 (N_19437,N_17406,N_16383);
and U19438 (N_19438,N_15078,N_15582);
xor U19439 (N_19439,N_16276,N_15415);
and U19440 (N_19440,N_16571,N_17258);
nand U19441 (N_19441,N_15594,N_16005);
nor U19442 (N_19442,N_16854,N_17919);
and U19443 (N_19443,N_17984,N_17213);
nand U19444 (N_19444,N_17261,N_15926);
nor U19445 (N_19445,N_17290,N_15223);
and U19446 (N_19446,N_15574,N_16415);
or U19447 (N_19447,N_17400,N_16863);
nor U19448 (N_19448,N_16570,N_16865);
nand U19449 (N_19449,N_16228,N_15370);
nand U19450 (N_19450,N_17581,N_15975);
and U19451 (N_19451,N_17295,N_16284);
nand U19452 (N_19452,N_15107,N_17178);
nand U19453 (N_19453,N_16001,N_17228);
xnor U19454 (N_19454,N_15766,N_15378);
nor U19455 (N_19455,N_16471,N_15940);
xnor U19456 (N_19456,N_17393,N_15619);
xnor U19457 (N_19457,N_16668,N_16595);
nor U19458 (N_19458,N_16725,N_17300);
nor U19459 (N_19459,N_16489,N_17246);
or U19460 (N_19460,N_15882,N_15114);
nor U19461 (N_19461,N_17223,N_15449);
and U19462 (N_19462,N_17439,N_15614);
and U19463 (N_19463,N_15075,N_17817);
nand U19464 (N_19464,N_15261,N_15297);
nor U19465 (N_19465,N_15599,N_16225);
or U19466 (N_19466,N_15840,N_15133);
xnor U19467 (N_19467,N_15953,N_16200);
nand U19468 (N_19468,N_16011,N_17187);
and U19469 (N_19469,N_17927,N_17383);
and U19470 (N_19470,N_17836,N_15893);
or U19471 (N_19471,N_15711,N_17902);
nor U19472 (N_19472,N_15411,N_16670);
nand U19473 (N_19473,N_16893,N_15818);
nand U19474 (N_19474,N_16693,N_16374);
nand U19475 (N_19475,N_16108,N_16278);
nor U19476 (N_19476,N_16777,N_15737);
nand U19477 (N_19477,N_16983,N_16528);
nor U19478 (N_19478,N_17431,N_15670);
and U19479 (N_19479,N_17204,N_16543);
and U19480 (N_19480,N_16568,N_17263);
and U19481 (N_19481,N_17541,N_17859);
and U19482 (N_19482,N_15553,N_17044);
or U19483 (N_19483,N_17302,N_17512);
or U19484 (N_19484,N_17226,N_15870);
and U19485 (N_19485,N_17548,N_16623);
xor U19486 (N_19486,N_16151,N_15215);
nand U19487 (N_19487,N_17578,N_16441);
and U19488 (N_19488,N_15082,N_16161);
and U19489 (N_19489,N_15119,N_16048);
xnor U19490 (N_19490,N_15878,N_15323);
nor U19491 (N_19491,N_16931,N_17498);
or U19492 (N_19492,N_17631,N_16516);
nand U19493 (N_19493,N_16718,N_15491);
xnor U19494 (N_19494,N_17330,N_15117);
and U19495 (N_19495,N_17988,N_16569);
nand U19496 (N_19496,N_15789,N_16642);
nand U19497 (N_19497,N_15431,N_15175);
nand U19498 (N_19498,N_17048,N_15883);
nor U19499 (N_19499,N_16041,N_17543);
xor U19500 (N_19500,N_15604,N_15705);
and U19501 (N_19501,N_17071,N_15672);
nand U19502 (N_19502,N_16092,N_15708);
nand U19503 (N_19503,N_15307,N_15275);
xnor U19504 (N_19504,N_15630,N_15112);
or U19505 (N_19505,N_15891,N_15737);
and U19506 (N_19506,N_16233,N_15700);
xor U19507 (N_19507,N_16295,N_16682);
xor U19508 (N_19508,N_15719,N_15376);
nor U19509 (N_19509,N_16845,N_16822);
or U19510 (N_19510,N_17204,N_16398);
and U19511 (N_19511,N_17354,N_15192);
and U19512 (N_19512,N_15280,N_15495);
xor U19513 (N_19513,N_15386,N_15037);
nor U19514 (N_19514,N_15194,N_15827);
and U19515 (N_19515,N_17364,N_15032);
xnor U19516 (N_19516,N_16626,N_17195);
and U19517 (N_19517,N_15169,N_15356);
or U19518 (N_19518,N_17217,N_17830);
or U19519 (N_19519,N_15614,N_15733);
or U19520 (N_19520,N_17037,N_16359);
and U19521 (N_19521,N_16655,N_16522);
or U19522 (N_19522,N_17936,N_17580);
and U19523 (N_19523,N_15676,N_17285);
xnor U19524 (N_19524,N_15433,N_17950);
or U19525 (N_19525,N_15414,N_17889);
or U19526 (N_19526,N_16763,N_15412);
and U19527 (N_19527,N_15857,N_16396);
or U19528 (N_19528,N_17218,N_16370);
nand U19529 (N_19529,N_15963,N_16595);
and U19530 (N_19530,N_17595,N_15569);
nand U19531 (N_19531,N_17614,N_17701);
nand U19532 (N_19532,N_17844,N_15878);
nor U19533 (N_19533,N_16663,N_15178);
nor U19534 (N_19534,N_16693,N_17509);
nor U19535 (N_19535,N_17653,N_16394);
nor U19536 (N_19536,N_15939,N_17915);
nand U19537 (N_19537,N_17615,N_16977);
nand U19538 (N_19538,N_17055,N_17606);
and U19539 (N_19539,N_16732,N_17342);
nand U19540 (N_19540,N_17156,N_15639);
or U19541 (N_19541,N_15653,N_16927);
and U19542 (N_19542,N_16033,N_16684);
nand U19543 (N_19543,N_17128,N_15821);
or U19544 (N_19544,N_17775,N_17482);
nor U19545 (N_19545,N_16693,N_16071);
or U19546 (N_19546,N_17923,N_17072);
and U19547 (N_19547,N_17152,N_15011);
nor U19548 (N_19548,N_15579,N_15531);
or U19549 (N_19549,N_16185,N_15851);
nor U19550 (N_19550,N_15607,N_16862);
nand U19551 (N_19551,N_16090,N_16273);
nand U19552 (N_19552,N_15525,N_15750);
or U19553 (N_19553,N_15839,N_17709);
and U19554 (N_19554,N_16122,N_16895);
xnor U19555 (N_19555,N_15258,N_17903);
or U19556 (N_19556,N_17794,N_17260);
or U19557 (N_19557,N_16802,N_17082);
xnor U19558 (N_19558,N_15531,N_17961);
nor U19559 (N_19559,N_15686,N_15365);
nand U19560 (N_19560,N_16574,N_16409);
nand U19561 (N_19561,N_17397,N_15437);
nand U19562 (N_19562,N_17153,N_17796);
or U19563 (N_19563,N_16430,N_15707);
or U19564 (N_19564,N_17492,N_17766);
or U19565 (N_19565,N_16551,N_15031);
nor U19566 (N_19566,N_16920,N_15339);
xnor U19567 (N_19567,N_15857,N_15739);
nor U19568 (N_19568,N_16973,N_16192);
nand U19569 (N_19569,N_15641,N_15255);
and U19570 (N_19570,N_15757,N_16534);
nand U19571 (N_19571,N_17247,N_16113);
or U19572 (N_19572,N_17125,N_15093);
and U19573 (N_19573,N_15166,N_17246);
and U19574 (N_19574,N_16823,N_17476);
nor U19575 (N_19575,N_15618,N_16243);
nand U19576 (N_19576,N_15352,N_17846);
nor U19577 (N_19577,N_15526,N_15154);
nand U19578 (N_19578,N_17951,N_16893);
nor U19579 (N_19579,N_16129,N_17240);
or U19580 (N_19580,N_16640,N_15787);
or U19581 (N_19581,N_17958,N_15998);
nand U19582 (N_19582,N_16999,N_17002);
and U19583 (N_19583,N_15632,N_16432);
nor U19584 (N_19584,N_15493,N_16515);
xor U19585 (N_19585,N_15525,N_16804);
or U19586 (N_19586,N_15082,N_17768);
nor U19587 (N_19587,N_16664,N_17377);
nand U19588 (N_19588,N_15994,N_16399);
nor U19589 (N_19589,N_15986,N_16597);
nor U19590 (N_19590,N_17000,N_16437);
or U19591 (N_19591,N_15681,N_16101);
or U19592 (N_19592,N_16040,N_17089);
nor U19593 (N_19593,N_15551,N_16306);
and U19594 (N_19594,N_16550,N_16165);
nand U19595 (N_19595,N_17588,N_15311);
nor U19596 (N_19596,N_17504,N_16011);
and U19597 (N_19597,N_16477,N_17607);
nor U19598 (N_19598,N_17658,N_17833);
nand U19599 (N_19599,N_16665,N_15718);
or U19600 (N_19600,N_16160,N_17520);
nor U19601 (N_19601,N_16836,N_16618);
and U19602 (N_19602,N_17750,N_15478);
nand U19603 (N_19603,N_16730,N_17948);
nand U19604 (N_19604,N_17131,N_16225);
xnor U19605 (N_19605,N_16036,N_17190);
and U19606 (N_19606,N_17197,N_17158);
and U19607 (N_19607,N_16195,N_16702);
nand U19608 (N_19608,N_15053,N_16510);
nor U19609 (N_19609,N_17242,N_16015);
nand U19610 (N_19610,N_17749,N_16767);
xor U19611 (N_19611,N_15728,N_16228);
xnor U19612 (N_19612,N_15343,N_15027);
nor U19613 (N_19613,N_17272,N_15555);
or U19614 (N_19614,N_16284,N_17746);
nand U19615 (N_19615,N_16693,N_16144);
nor U19616 (N_19616,N_17213,N_15817);
nand U19617 (N_19617,N_16930,N_17222);
or U19618 (N_19618,N_17870,N_17745);
or U19619 (N_19619,N_15968,N_16996);
xnor U19620 (N_19620,N_17471,N_16039);
and U19621 (N_19621,N_15129,N_17778);
xor U19622 (N_19622,N_17453,N_15843);
xnor U19623 (N_19623,N_15219,N_15783);
and U19624 (N_19624,N_15122,N_15693);
or U19625 (N_19625,N_17806,N_17838);
xor U19626 (N_19626,N_16475,N_15557);
xnor U19627 (N_19627,N_15762,N_15279);
nand U19628 (N_19628,N_15954,N_17516);
or U19629 (N_19629,N_15150,N_15417);
nor U19630 (N_19630,N_15798,N_15626);
or U19631 (N_19631,N_17630,N_15491);
and U19632 (N_19632,N_16370,N_17063);
nand U19633 (N_19633,N_15676,N_15713);
nor U19634 (N_19634,N_17652,N_16508);
and U19635 (N_19635,N_17854,N_15411);
nor U19636 (N_19636,N_17280,N_15373);
xor U19637 (N_19637,N_16380,N_15551);
nand U19638 (N_19638,N_15415,N_15497);
or U19639 (N_19639,N_16474,N_16631);
nor U19640 (N_19640,N_17577,N_15464);
nor U19641 (N_19641,N_16921,N_15741);
and U19642 (N_19642,N_16220,N_15325);
xor U19643 (N_19643,N_16771,N_15743);
nor U19644 (N_19644,N_15586,N_16161);
and U19645 (N_19645,N_15686,N_17796);
and U19646 (N_19646,N_17626,N_15203);
or U19647 (N_19647,N_15753,N_15197);
nor U19648 (N_19648,N_15126,N_16060);
nor U19649 (N_19649,N_15857,N_15064);
nand U19650 (N_19650,N_15409,N_17668);
nor U19651 (N_19651,N_16359,N_17348);
xnor U19652 (N_19652,N_17981,N_15728);
nor U19653 (N_19653,N_15006,N_17762);
nor U19654 (N_19654,N_16583,N_15919);
nor U19655 (N_19655,N_17601,N_17351);
and U19656 (N_19656,N_17630,N_17000);
xnor U19657 (N_19657,N_16408,N_15431);
nand U19658 (N_19658,N_17762,N_17583);
nand U19659 (N_19659,N_15647,N_16971);
nand U19660 (N_19660,N_17132,N_17669);
nor U19661 (N_19661,N_16059,N_17630);
nand U19662 (N_19662,N_15090,N_15867);
nand U19663 (N_19663,N_16445,N_15667);
xor U19664 (N_19664,N_16189,N_15781);
or U19665 (N_19665,N_16076,N_16919);
and U19666 (N_19666,N_17343,N_17654);
and U19667 (N_19667,N_16357,N_16606);
and U19668 (N_19668,N_15514,N_15650);
xor U19669 (N_19669,N_17801,N_16856);
or U19670 (N_19670,N_16714,N_15052);
and U19671 (N_19671,N_16913,N_16425);
xnor U19672 (N_19672,N_16318,N_16087);
xor U19673 (N_19673,N_17299,N_15273);
or U19674 (N_19674,N_16014,N_16840);
nand U19675 (N_19675,N_16688,N_17424);
nand U19676 (N_19676,N_15833,N_16257);
and U19677 (N_19677,N_16837,N_16817);
nor U19678 (N_19678,N_15783,N_17299);
xnor U19679 (N_19679,N_17033,N_15602);
nand U19680 (N_19680,N_17259,N_15633);
nor U19681 (N_19681,N_16346,N_17533);
nor U19682 (N_19682,N_16912,N_16952);
nand U19683 (N_19683,N_16853,N_16975);
nand U19684 (N_19684,N_16856,N_15724);
and U19685 (N_19685,N_17140,N_15760);
nand U19686 (N_19686,N_16601,N_15251);
and U19687 (N_19687,N_17747,N_17523);
or U19688 (N_19688,N_16702,N_15616);
nand U19689 (N_19689,N_15673,N_15942);
xor U19690 (N_19690,N_15472,N_15999);
nand U19691 (N_19691,N_15898,N_17374);
and U19692 (N_19692,N_15961,N_15340);
nand U19693 (N_19693,N_15237,N_15721);
or U19694 (N_19694,N_17054,N_15306);
nor U19695 (N_19695,N_15852,N_16039);
or U19696 (N_19696,N_17232,N_16615);
or U19697 (N_19697,N_17630,N_16427);
nor U19698 (N_19698,N_16722,N_17637);
xnor U19699 (N_19699,N_17137,N_15682);
nor U19700 (N_19700,N_17586,N_16692);
and U19701 (N_19701,N_17491,N_15166);
or U19702 (N_19702,N_17548,N_17861);
nor U19703 (N_19703,N_17310,N_17522);
nor U19704 (N_19704,N_15705,N_17158);
xnor U19705 (N_19705,N_16906,N_16462);
and U19706 (N_19706,N_15645,N_16739);
nand U19707 (N_19707,N_16700,N_17848);
or U19708 (N_19708,N_15563,N_17239);
and U19709 (N_19709,N_17781,N_17394);
and U19710 (N_19710,N_16274,N_17428);
nand U19711 (N_19711,N_15623,N_17453);
nor U19712 (N_19712,N_15818,N_17753);
or U19713 (N_19713,N_17759,N_17794);
or U19714 (N_19714,N_16617,N_15607);
and U19715 (N_19715,N_16056,N_15498);
and U19716 (N_19716,N_17141,N_17906);
nor U19717 (N_19717,N_17490,N_16099);
and U19718 (N_19718,N_17057,N_17356);
nor U19719 (N_19719,N_17223,N_15158);
nand U19720 (N_19720,N_16863,N_16239);
and U19721 (N_19721,N_17324,N_17157);
nor U19722 (N_19722,N_16090,N_16874);
xnor U19723 (N_19723,N_17572,N_16801);
or U19724 (N_19724,N_15704,N_17048);
xor U19725 (N_19725,N_15969,N_16913);
xnor U19726 (N_19726,N_17529,N_16281);
nand U19727 (N_19727,N_16549,N_17901);
nand U19728 (N_19728,N_15348,N_17703);
and U19729 (N_19729,N_16408,N_16729);
nor U19730 (N_19730,N_15145,N_15293);
nand U19731 (N_19731,N_17737,N_16408);
and U19732 (N_19732,N_17027,N_16868);
nand U19733 (N_19733,N_17127,N_17911);
nand U19734 (N_19734,N_17847,N_15508);
and U19735 (N_19735,N_15389,N_16188);
nor U19736 (N_19736,N_16717,N_16281);
or U19737 (N_19737,N_17334,N_16416);
and U19738 (N_19738,N_17689,N_16141);
nor U19739 (N_19739,N_15149,N_16810);
xnor U19740 (N_19740,N_17747,N_15031);
and U19741 (N_19741,N_16177,N_15448);
and U19742 (N_19742,N_16777,N_16027);
xor U19743 (N_19743,N_17637,N_16355);
nor U19744 (N_19744,N_16747,N_17757);
xor U19745 (N_19745,N_17305,N_17715);
nor U19746 (N_19746,N_16709,N_16495);
nor U19747 (N_19747,N_16209,N_16461);
nand U19748 (N_19748,N_17751,N_16367);
and U19749 (N_19749,N_17119,N_16505);
nand U19750 (N_19750,N_16060,N_15885);
nor U19751 (N_19751,N_16637,N_15181);
or U19752 (N_19752,N_17597,N_17306);
xor U19753 (N_19753,N_17472,N_16126);
or U19754 (N_19754,N_15009,N_15853);
or U19755 (N_19755,N_16587,N_15960);
xor U19756 (N_19756,N_17689,N_15569);
and U19757 (N_19757,N_15862,N_17622);
nand U19758 (N_19758,N_15545,N_17960);
xor U19759 (N_19759,N_17216,N_15476);
or U19760 (N_19760,N_15352,N_15899);
and U19761 (N_19761,N_17825,N_15966);
or U19762 (N_19762,N_17378,N_17539);
or U19763 (N_19763,N_16493,N_16335);
nor U19764 (N_19764,N_17641,N_16579);
nor U19765 (N_19765,N_15951,N_17902);
and U19766 (N_19766,N_17718,N_17894);
xor U19767 (N_19767,N_16058,N_15823);
nor U19768 (N_19768,N_15661,N_16891);
and U19769 (N_19769,N_17886,N_17004);
xor U19770 (N_19770,N_17438,N_16157);
and U19771 (N_19771,N_16010,N_16833);
or U19772 (N_19772,N_17559,N_17469);
nor U19773 (N_19773,N_16506,N_15456);
nand U19774 (N_19774,N_17985,N_15961);
nand U19775 (N_19775,N_15377,N_16085);
nand U19776 (N_19776,N_17187,N_15666);
and U19777 (N_19777,N_17517,N_16218);
and U19778 (N_19778,N_16316,N_16852);
xor U19779 (N_19779,N_17088,N_17565);
nor U19780 (N_19780,N_17713,N_17267);
nor U19781 (N_19781,N_16975,N_16048);
xnor U19782 (N_19782,N_17671,N_17594);
nand U19783 (N_19783,N_16606,N_17629);
nand U19784 (N_19784,N_16728,N_15570);
nor U19785 (N_19785,N_16193,N_17208);
nor U19786 (N_19786,N_16497,N_16452);
and U19787 (N_19787,N_16327,N_17434);
nand U19788 (N_19788,N_17653,N_17183);
and U19789 (N_19789,N_17390,N_15409);
nor U19790 (N_19790,N_17533,N_15594);
and U19791 (N_19791,N_15655,N_16457);
and U19792 (N_19792,N_15596,N_16724);
nor U19793 (N_19793,N_15698,N_15794);
nor U19794 (N_19794,N_15596,N_16214);
nand U19795 (N_19795,N_17532,N_16162);
nand U19796 (N_19796,N_17007,N_17178);
xor U19797 (N_19797,N_15609,N_16561);
or U19798 (N_19798,N_17683,N_17694);
and U19799 (N_19799,N_17857,N_17737);
and U19800 (N_19800,N_15083,N_16110);
and U19801 (N_19801,N_15247,N_17164);
or U19802 (N_19802,N_17091,N_15288);
nand U19803 (N_19803,N_15110,N_15217);
xor U19804 (N_19804,N_16669,N_15269);
nor U19805 (N_19805,N_16437,N_15932);
and U19806 (N_19806,N_16149,N_15689);
nand U19807 (N_19807,N_15496,N_15810);
nor U19808 (N_19808,N_15097,N_16340);
and U19809 (N_19809,N_17013,N_17283);
nor U19810 (N_19810,N_16948,N_15437);
or U19811 (N_19811,N_15530,N_17416);
or U19812 (N_19812,N_17728,N_17474);
and U19813 (N_19813,N_15405,N_17254);
xor U19814 (N_19814,N_17952,N_17352);
and U19815 (N_19815,N_15279,N_15351);
nor U19816 (N_19816,N_16706,N_16340);
and U19817 (N_19817,N_15872,N_17521);
or U19818 (N_19818,N_15098,N_15727);
xnor U19819 (N_19819,N_16261,N_15788);
xnor U19820 (N_19820,N_16238,N_16006);
xnor U19821 (N_19821,N_17844,N_16360);
or U19822 (N_19822,N_16549,N_17140);
or U19823 (N_19823,N_17069,N_15345);
nand U19824 (N_19824,N_16957,N_15032);
xnor U19825 (N_19825,N_15553,N_15909);
nand U19826 (N_19826,N_17111,N_16170);
and U19827 (N_19827,N_16259,N_16244);
or U19828 (N_19828,N_15623,N_16605);
and U19829 (N_19829,N_16322,N_17708);
nand U19830 (N_19830,N_17810,N_17026);
nor U19831 (N_19831,N_17047,N_16556);
nand U19832 (N_19832,N_15622,N_17611);
nand U19833 (N_19833,N_15001,N_16863);
and U19834 (N_19834,N_15744,N_16228);
and U19835 (N_19835,N_17567,N_16252);
and U19836 (N_19836,N_17275,N_17415);
xnor U19837 (N_19837,N_15335,N_17595);
nor U19838 (N_19838,N_15342,N_16946);
nand U19839 (N_19839,N_16779,N_15046);
nor U19840 (N_19840,N_16601,N_17284);
or U19841 (N_19841,N_15573,N_17991);
and U19842 (N_19842,N_16449,N_15245);
and U19843 (N_19843,N_16968,N_15260);
xor U19844 (N_19844,N_16628,N_17730);
and U19845 (N_19845,N_15372,N_15153);
nor U19846 (N_19846,N_16129,N_16070);
and U19847 (N_19847,N_15433,N_17758);
and U19848 (N_19848,N_15883,N_16350);
nand U19849 (N_19849,N_15229,N_16783);
xor U19850 (N_19850,N_17394,N_16978);
or U19851 (N_19851,N_15280,N_17508);
or U19852 (N_19852,N_17943,N_17835);
or U19853 (N_19853,N_16575,N_15997);
nand U19854 (N_19854,N_17405,N_17591);
or U19855 (N_19855,N_16804,N_17968);
xor U19856 (N_19856,N_15779,N_17449);
or U19857 (N_19857,N_16132,N_15595);
nand U19858 (N_19858,N_15645,N_16713);
xor U19859 (N_19859,N_16061,N_16573);
nor U19860 (N_19860,N_15169,N_16315);
nor U19861 (N_19861,N_16455,N_16342);
and U19862 (N_19862,N_15521,N_17142);
and U19863 (N_19863,N_17122,N_17478);
nor U19864 (N_19864,N_17237,N_16657);
nand U19865 (N_19865,N_17459,N_17168);
and U19866 (N_19866,N_17987,N_16979);
nor U19867 (N_19867,N_16315,N_17676);
and U19868 (N_19868,N_17826,N_15803);
nor U19869 (N_19869,N_16925,N_16333);
or U19870 (N_19870,N_17305,N_17504);
or U19871 (N_19871,N_15340,N_15409);
nor U19872 (N_19872,N_15070,N_16280);
and U19873 (N_19873,N_15093,N_17238);
nand U19874 (N_19874,N_15701,N_15067);
or U19875 (N_19875,N_15037,N_17625);
xnor U19876 (N_19876,N_16600,N_17176);
nand U19877 (N_19877,N_15224,N_17660);
or U19878 (N_19878,N_15052,N_15640);
nor U19879 (N_19879,N_15348,N_17312);
xor U19880 (N_19880,N_17950,N_17468);
xor U19881 (N_19881,N_17821,N_17927);
or U19882 (N_19882,N_15683,N_15417);
xor U19883 (N_19883,N_15040,N_15969);
xor U19884 (N_19884,N_17365,N_17141);
nand U19885 (N_19885,N_15814,N_15138);
xnor U19886 (N_19886,N_17264,N_17687);
and U19887 (N_19887,N_16498,N_17047);
and U19888 (N_19888,N_15509,N_16613);
or U19889 (N_19889,N_17321,N_15849);
nand U19890 (N_19890,N_15329,N_16901);
or U19891 (N_19891,N_17805,N_16023);
and U19892 (N_19892,N_17470,N_16727);
and U19893 (N_19893,N_16002,N_17648);
nand U19894 (N_19894,N_17376,N_15072);
xnor U19895 (N_19895,N_15616,N_17717);
and U19896 (N_19896,N_17857,N_17602);
nand U19897 (N_19897,N_17689,N_16830);
xnor U19898 (N_19898,N_15897,N_15731);
and U19899 (N_19899,N_17813,N_16968);
or U19900 (N_19900,N_16144,N_17230);
nand U19901 (N_19901,N_17612,N_15540);
nor U19902 (N_19902,N_15449,N_17975);
xor U19903 (N_19903,N_16851,N_17390);
xor U19904 (N_19904,N_15501,N_17231);
and U19905 (N_19905,N_15823,N_15456);
nand U19906 (N_19906,N_16313,N_15420);
and U19907 (N_19907,N_16922,N_15085);
nor U19908 (N_19908,N_17369,N_15032);
or U19909 (N_19909,N_17203,N_15742);
nand U19910 (N_19910,N_15526,N_16183);
nand U19911 (N_19911,N_16141,N_16921);
or U19912 (N_19912,N_15542,N_16459);
nor U19913 (N_19913,N_16026,N_16373);
nor U19914 (N_19914,N_16516,N_16315);
and U19915 (N_19915,N_17532,N_15588);
nor U19916 (N_19916,N_17340,N_16715);
nor U19917 (N_19917,N_17592,N_17168);
xor U19918 (N_19918,N_16162,N_16946);
xnor U19919 (N_19919,N_15169,N_17043);
xnor U19920 (N_19920,N_15872,N_15216);
or U19921 (N_19921,N_16221,N_15054);
nor U19922 (N_19922,N_17726,N_17817);
xor U19923 (N_19923,N_15550,N_16662);
nor U19924 (N_19924,N_15465,N_15555);
nand U19925 (N_19925,N_17909,N_15296);
or U19926 (N_19926,N_15147,N_16970);
xor U19927 (N_19927,N_16435,N_16115);
nand U19928 (N_19928,N_16144,N_17234);
or U19929 (N_19929,N_15872,N_16512);
xnor U19930 (N_19930,N_17081,N_16900);
or U19931 (N_19931,N_15674,N_17491);
nor U19932 (N_19932,N_15369,N_15638);
and U19933 (N_19933,N_16021,N_17761);
nand U19934 (N_19934,N_17486,N_15959);
xor U19935 (N_19935,N_15278,N_16895);
nor U19936 (N_19936,N_17174,N_15032);
nand U19937 (N_19937,N_16755,N_15598);
or U19938 (N_19938,N_16588,N_17330);
xnor U19939 (N_19939,N_17408,N_17464);
nand U19940 (N_19940,N_16177,N_17816);
nand U19941 (N_19941,N_16964,N_15590);
xnor U19942 (N_19942,N_16966,N_16894);
and U19943 (N_19943,N_17069,N_17938);
nor U19944 (N_19944,N_17986,N_15530);
or U19945 (N_19945,N_17509,N_16382);
or U19946 (N_19946,N_16959,N_16394);
and U19947 (N_19947,N_17469,N_16848);
nor U19948 (N_19948,N_17076,N_17702);
nor U19949 (N_19949,N_15814,N_15464);
and U19950 (N_19950,N_16875,N_15444);
nand U19951 (N_19951,N_17160,N_16459);
nor U19952 (N_19952,N_17848,N_17291);
and U19953 (N_19953,N_15830,N_16957);
nand U19954 (N_19954,N_15507,N_16723);
or U19955 (N_19955,N_16972,N_15358);
or U19956 (N_19956,N_16464,N_15251);
xnor U19957 (N_19957,N_16190,N_17195);
or U19958 (N_19958,N_17237,N_17966);
or U19959 (N_19959,N_15491,N_16515);
xnor U19960 (N_19960,N_17976,N_15528);
or U19961 (N_19961,N_16768,N_17539);
or U19962 (N_19962,N_15655,N_15794);
and U19963 (N_19963,N_16972,N_15267);
xnor U19964 (N_19964,N_16361,N_17808);
and U19965 (N_19965,N_17430,N_16219);
nand U19966 (N_19966,N_15874,N_15574);
nor U19967 (N_19967,N_15422,N_17932);
or U19968 (N_19968,N_16240,N_16701);
nor U19969 (N_19969,N_17090,N_15660);
or U19970 (N_19970,N_16826,N_15690);
or U19971 (N_19971,N_16371,N_15017);
and U19972 (N_19972,N_16857,N_15935);
xor U19973 (N_19973,N_17290,N_15139);
nand U19974 (N_19974,N_17051,N_15180);
and U19975 (N_19975,N_17102,N_17151);
and U19976 (N_19976,N_15057,N_15130);
or U19977 (N_19977,N_17981,N_16631);
or U19978 (N_19978,N_16877,N_17917);
and U19979 (N_19979,N_15596,N_15820);
and U19980 (N_19980,N_15974,N_17217);
nor U19981 (N_19981,N_16065,N_17648);
and U19982 (N_19982,N_15102,N_16867);
and U19983 (N_19983,N_16979,N_17284);
or U19984 (N_19984,N_16418,N_17884);
nand U19985 (N_19985,N_15200,N_16465);
nor U19986 (N_19986,N_16965,N_17763);
nor U19987 (N_19987,N_17645,N_17281);
or U19988 (N_19988,N_17955,N_15611);
nand U19989 (N_19989,N_17446,N_17474);
xnor U19990 (N_19990,N_16940,N_17785);
nand U19991 (N_19991,N_17046,N_16774);
and U19992 (N_19992,N_15531,N_17970);
or U19993 (N_19993,N_17557,N_15563);
xor U19994 (N_19994,N_16901,N_16204);
nor U19995 (N_19995,N_16440,N_15745);
and U19996 (N_19996,N_17478,N_16545);
or U19997 (N_19997,N_17364,N_16867);
and U19998 (N_19998,N_17591,N_17355);
or U19999 (N_19999,N_15355,N_16431);
and U20000 (N_20000,N_15672,N_16681);
nand U20001 (N_20001,N_17992,N_17764);
or U20002 (N_20002,N_15755,N_17672);
nand U20003 (N_20003,N_16103,N_15181);
and U20004 (N_20004,N_16804,N_17493);
or U20005 (N_20005,N_16371,N_16883);
and U20006 (N_20006,N_15337,N_15018);
nand U20007 (N_20007,N_16837,N_15525);
nand U20008 (N_20008,N_16927,N_16867);
or U20009 (N_20009,N_15532,N_15147);
xor U20010 (N_20010,N_15533,N_17708);
xnor U20011 (N_20011,N_16558,N_17610);
or U20012 (N_20012,N_15841,N_16709);
and U20013 (N_20013,N_17848,N_16696);
xnor U20014 (N_20014,N_15676,N_17375);
nor U20015 (N_20015,N_15537,N_17518);
xor U20016 (N_20016,N_17227,N_15674);
or U20017 (N_20017,N_15335,N_16327);
or U20018 (N_20018,N_15960,N_16234);
or U20019 (N_20019,N_17462,N_15587);
or U20020 (N_20020,N_15106,N_17007);
nand U20021 (N_20021,N_16965,N_15602);
xor U20022 (N_20022,N_17196,N_17784);
and U20023 (N_20023,N_16544,N_16770);
or U20024 (N_20024,N_16894,N_15707);
nor U20025 (N_20025,N_15829,N_16916);
xor U20026 (N_20026,N_16791,N_16639);
nand U20027 (N_20027,N_17960,N_17993);
and U20028 (N_20028,N_15862,N_17700);
or U20029 (N_20029,N_15335,N_16161);
nand U20030 (N_20030,N_16482,N_17366);
nand U20031 (N_20031,N_16214,N_16160);
nand U20032 (N_20032,N_16461,N_16789);
nand U20033 (N_20033,N_16016,N_16470);
nor U20034 (N_20034,N_16690,N_16758);
nand U20035 (N_20035,N_16708,N_15407);
xor U20036 (N_20036,N_15074,N_16066);
nand U20037 (N_20037,N_16635,N_15150);
and U20038 (N_20038,N_17785,N_17502);
nand U20039 (N_20039,N_16582,N_15112);
nor U20040 (N_20040,N_15061,N_16565);
nand U20041 (N_20041,N_15221,N_17351);
nor U20042 (N_20042,N_17834,N_17709);
and U20043 (N_20043,N_15440,N_15251);
and U20044 (N_20044,N_15560,N_17545);
or U20045 (N_20045,N_17641,N_17354);
xor U20046 (N_20046,N_16087,N_15081);
nor U20047 (N_20047,N_16181,N_17595);
xor U20048 (N_20048,N_15388,N_16334);
or U20049 (N_20049,N_15355,N_17472);
nand U20050 (N_20050,N_17810,N_16890);
and U20051 (N_20051,N_17214,N_17971);
and U20052 (N_20052,N_16354,N_16877);
or U20053 (N_20053,N_17926,N_16456);
nand U20054 (N_20054,N_17936,N_15677);
nand U20055 (N_20055,N_15036,N_16069);
or U20056 (N_20056,N_16503,N_17477);
nand U20057 (N_20057,N_17474,N_17203);
or U20058 (N_20058,N_16229,N_16431);
nor U20059 (N_20059,N_15553,N_17706);
and U20060 (N_20060,N_16164,N_15568);
nand U20061 (N_20061,N_16559,N_16131);
nand U20062 (N_20062,N_17823,N_15831);
nor U20063 (N_20063,N_17569,N_15124);
nand U20064 (N_20064,N_16842,N_17192);
nand U20065 (N_20065,N_16407,N_17116);
xnor U20066 (N_20066,N_16440,N_16185);
and U20067 (N_20067,N_15398,N_15956);
and U20068 (N_20068,N_15894,N_17354);
nand U20069 (N_20069,N_16765,N_15101);
xor U20070 (N_20070,N_16758,N_17385);
xnor U20071 (N_20071,N_17875,N_17416);
nand U20072 (N_20072,N_16897,N_16389);
or U20073 (N_20073,N_15238,N_16858);
xnor U20074 (N_20074,N_16502,N_16744);
and U20075 (N_20075,N_17504,N_15298);
and U20076 (N_20076,N_17883,N_16160);
nor U20077 (N_20077,N_17700,N_16378);
and U20078 (N_20078,N_15569,N_16093);
xnor U20079 (N_20079,N_16650,N_16327);
nand U20080 (N_20080,N_17950,N_17659);
and U20081 (N_20081,N_16270,N_17350);
nor U20082 (N_20082,N_16162,N_16407);
xor U20083 (N_20083,N_16241,N_17975);
and U20084 (N_20084,N_16746,N_16497);
and U20085 (N_20085,N_15072,N_16702);
or U20086 (N_20086,N_15915,N_16412);
or U20087 (N_20087,N_16124,N_16440);
nand U20088 (N_20088,N_16718,N_16403);
and U20089 (N_20089,N_17797,N_15689);
nand U20090 (N_20090,N_15833,N_15911);
nand U20091 (N_20091,N_17369,N_15057);
or U20092 (N_20092,N_16088,N_16912);
xor U20093 (N_20093,N_15872,N_15193);
xnor U20094 (N_20094,N_15836,N_17228);
nor U20095 (N_20095,N_17545,N_16957);
or U20096 (N_20096,N_16828,N_15020);
and U20097 (N_20097,N_17876,N_17061);
xor U20098 (N_20098,N_16012,N_15323);
xor U20099 (N_20099,N_15253,N_17931);
and U20100 (N_20100,N_15515,N_15909);
nand U20101 (N_20101,N_17825,N_15749);
nand U20102 (N_20102,N_15406,N_17852);
nor U20103 (N_20103,N_17094,N_16861);
xnor U20104 (N_20104,N_16882,N_16603);
nor U20105 (N_20105,N_17089,N_17346);
xnor U20106 (N_20106,N_17379,N_15767);
or U20107 (N_20107,N_15029,N_16677);
nand U20108 (N_20108,N_15304,N_16782);
xor U20109 (N_20109,N_16438,N_17495);
xnor U20110 (N_20110,N_15511,N_16052);
nand U20111 (N_20111,N_17447,N_15367);
nor U20112 (N_20112,N_15239,N_16410);
xor U20113 (N_20113,N_17498,N_17352);
xor U20114 (N_20114,N_15959,N_16700);
nand U20115 (N_20115,N_16164,N_15396);
and U20116 (N_20116,N_16759,N_15544);
nor U20117 (N_20117,N_17210,N_15189);
nand U20118 (N_20118,N_17802,N_15246);
nor U20119 (N_20119,N_16661,N_17976);
nand U20120 (N_20120,N_16163,N_15769);
xnor U20121 (N_20121,N_16434,N_17807);
or U20122 (N_20122,N_17987,N_16252);
xor U20123 (N_20123,N_17952,N_15794);
nand U20124 (N_20124,N_15192,N_15022);
and U20125 (N_20125,N_16852,N_17998);
and U20126 (N_20126,N_16154,N_15604);
nand U20127 (N_20127,N_16769,N_16028);
nor U20128 (N_20128,N_15984,N_17599);
xnor U20129 (N_20129,N_16571,N_15573);
and U20130 (N_20130,N_16953,N_17239);
nand U20131 (N_20131,N_15390,N_17520);
and U20132 (N_20132,N_15651,N_16308);
or U20133 (N_20133,N_17239,N_17462);
xnor U20134 (N_20134,N_15941,N_16964);
nor U20135 (N_20135,N_15486,N_17892);
and U20136 (N_20136,N_16875,N_16596);
xor U20137 (N_20137,N_15477,N_15152);
or U20138 (N_20138,N_16023,N_16222);
xnor U20139 (N_20139,N_16814,N_17845);
nor U20140 (N_20140,N_16916,N_15011);
xor U20141 (N_20141,N_15458,N_15986);
nor U20142 (N_20142,N_16673,N_16736);
xnor U20143 (N_20143,N_16496,N_16600);
nor U20144 (N_20144,N_15986,N_16357);
or U20145 (N_20145,N_17878,N_15069);
nand U20146 (N_20146,N_17492,N_17097);
nor U20147 (N_20147,N_17409,N_17685);
xnor U20148 (N_20148,N_15856,N_15967);
xnor U20149 (N_20149,N_17469,N_17849);
and U20150 (N_20150,N_15842,N_15908);
nand U20151 (N_20151,N_15151,N_17343);
nand U20152 (N_20152,N_15454,N_16636);
or U20153 (N_20153,N_16421,N_17356);
nand U20154 (N_20154,N_16577,N_17160);
and U20155 (N_20155,N_15106,N_16768);
xnor U20156 (N_20156,N_17131,N_17919);
nand U20157 (N_20157,N_17965,N_16085);
xnor U20158 (N_20158,N_17715,N_17342);
or U20159 (N_20159,N_15568,N_15969);
nand U20160 (N_20160,N_15178,N_17589);
nor U20161 (N_20161,N_16363,N_17034);
nor U20162 (N_20162,N_16082,N_16111);
nand U20163 (N_20163,N_16160,N_17028);
nand U20164 (N_20164,N_17359,N_15901);
or U20165 (N_20165,N_15499,N_15874);
or U20166 (N_20166,N_17958,N_15903);
nand U20167 (N_20167,N_17235,N_15393);
or U20168 (N_20168,N_17746,N_17852);
nand U20169 (N_20169,N_15638,N_17234);
or U20170 (N_20170,N_16936,N_17241);
xor U20171 (N_20171,N_17771,N_15796);
xor U20172 (N_20172,N_15419,N_16606);
or U20173 (N_20173,N_15890,N_16167);
nand U20174 (N_20174,N_15314,N_15202);
nor U20175 (N_20175,N_15151,N_17180);
or U20176 (N_20176,N_15649,N_16953);
xor U20177 (N_20177,N_15408,N_16292);
and U20178 (N_20178,N_15471,N_17716);
and U20179 (N_20179,N_15879,N_16366);
xor U20180 (N_20180,N_15078,N_16082);
xnor U20181 (N_20181,N_15432,N_16950);
and U20182 (N_20182,N_17888,N_16728);
nand U20183 (N_20183,N_16482,N_16782);
nor U20184 (N_20184,N_17930,N_17248);
xnor U20185 (N_20185,N_17781,N_15929);
nand U20186 (N_20186,N_16175,N_17024);
and U20187 (N_20187,N_15040,N_16493);
or U20188 (N_20188,N_15196,N_16814);
nand U20189 (N_20189,N_17013,N_17002);
or U20190 (N_20190,N_16260,N_15671);
nor U20191 (N_20191,N_16904,N_17999);
xnor U20192 (N_20192,N_17267,N_17818);
xnor U20193 (N_20193,N_16161,N_15881);
and U20194 (N_20194,N_17514,N_17188);
and U20195 (N_20195,N_15298,N_16437);
xnor U20196 (N_20196,N_16596,N_16457);
nor U20197 (N_20197,N_15000,N_15740);
nand U20198 (N_20198,N_17939,N_17796);
nand U20199 (N_20199,N_17284,N_16198);
nand U20200 (N_20200,N_15171,N_15188);
xnor U20201 (N_20201,N_15063,N_15079);
xor U20202 (N_20202,N_17695,N_16460);
nor U20203 (N_20203,N_16463,N_15241);
nand U20204 (N_20204,N_17113,N_16923);
xnor U20205 (N_20205,N_17717,N_15151);
and U20206 (N_20206,N_17116,N_17886);
or U20207 (N_20207,N_15724,N_15250);
or U20208 (N_20208,N_15452,N_15740);
or U20209 (N_20209,N_16780,N_15200);
xnor U20210 (N_20210,N_16220,N_16204);
and U20211 (N_20211,N_17157,N_17276);
and U20212 (N_20212,N_17924,N_15504);
or U20213 (N_20213,N_16791,N_15354);
or U20214 (N_20214,N_16687,N_15831);
xnor U20215 (N_20215,N_17493,N_15864);
nor U20216 (N_20216,N_15064,N_17271);
nand U20217 (N_20217,N_15152,N_15569);
nor U20218 (N_20218,N_17152,N_17366);
and U20219 (N_20219,N_15574,N_15111);
xor U20220 (N_20220,N_17510,N_15251);
or U20221 (N_20221,N_17076,N_15091);
or U20222 (N_20222,N_17401,N_17717);
nor U20223 (N_20223,N_16459,N_16475);
nand U20224 (N_20224,N_17938,N_15949);
nor U20225 (N_20225,N_16067,N_17864);
xnor U20226 (N_20226,N_15102,N_16561);
or U20227 (N_20227,N_17310,N_15702);
xor U20228 (N_20228,N_17946,N_16979);
and U20229 (N_20229,N_17329,N_15580);
nor U20230 (N_20230,N_16554,N_17729);
and U20231 (N_20231,N_15732,N_17536);
xnor U20232 (N_20232,N_16024,N_16037);
and U20233 (N_20233,N_16062,N_17793);
xor U20234 (N_20234,N_17129,N_16827);
xor U20235 (N_20235,N_17956,N_16154);
and U20236 (N_20236,N_15607,N_15123);
xor U20237 (N_20237,N_16956,N_16192);
nand U20238 (N_20238,N_17861,N_16595);
or U20239 (N_20239,N_15522,N_15201);
and U20240 (N_20240,N_17618,N_16921);
nor U20241 (N_20241,N_17100,N_17210);
xor U20242 (N_20242,N_16213,N_16496);
nand U20243 (N_20243,N_16223,N_15441);
and U20244 (N_20244,N_17922,N_15022);
and U20245 (N_20245,N_15740,N_16940);
xnor U20246 (N_20246,N_16766,N_15313);
nand U20247 (N_20247,N_16645,N_15271);
or U20248 (N_20248,N_16275,N_15454);
and U20249 (N_20249,N_16531,N_15407);
nand U20250 (N_20250,N_16228,N_15098);
and U20251 (N_20251,N_15228,N_17379);
and U20252 (N_20252,N_15392,N_16263);
nor U20253 (N_20253,N_15237,N_17723);
and U20254 (N_20254,N_15846,N_15768);
nor U20255 (N_20255,N_16085,N_17228);
or U20256 (N_20256,N_17268,N_15780);
nor U20257 (N_20257,N_15381,N_16444);
and U20258 (N_20258,N_15242,N_17048);
and U20259 (N_20259,N_17817,N_16533);
or U20260 (N_20260,N_16010,N_17871);
or U20261 (N_20261,N_15647,N_15324);
nor U20262 (N_20262,N_15213,N_16964);
nand U20263 (N_20263,N_15190,N_17546);
or U20264 (N_20264,N_16086,N_17300);
or U20265 (N_20265,N_17494,N_17411);
xnor U20266 (N_20266,N_16398,N_17851);
nand U20267 (N_20267,N_16160,N_16361);
or U20268 (N_20268,N_15980,N_17805);
and U20269 (N_20269,N_15899,N_15249);
nand U20270 (N_20270,N_15376,N_16040);
and U20271 (N_20271,N_17992,N_15157);
or U20272 (N_20272,N_16468,N_17877);
or U20273 (N_20273,N_16736,N_16407);
nor U20274 (N_20274,N_15045,N_15433);
nand U20275 (N_20275,N_16543,N_17487);
nand U20276 (N_20276,N_16743,N_17504);
or U20277 (N_20277,N_16941,N_16114);
and U20278 (N_20278,N_15323,N_15124);
or U20279 (N_20279,N_16305,N_17483);
and U20280 (N_20280,N_17937,N_15630);
nor U20281 (N_20281,N_15313,N_16290);
or U20282 (N_20282,N_16385,N_16802);
xor U20283 (N_20283,N_16669,N_15611);
xor U20284 (N_20284,N_16970,N_16063);
nor U20285 (N_20285,N_17830,N_16130);
and U20286 (N_20286,N_17470,N_17887);
or U20287 (N_20287,N_17924,N_15614);
nor U20288 (N_20288,N_15794,N_15707);
nand U20289 (N_20289,N_15091,N_17779);
xor U20290 (N_20290,N_17778,N_16506);
nor U20291 (N_20291,N_15892,N_17491);
nor U20292 (N_20292,N_15378,N_15003);
nand U20293 (N_20293,N_17426,N_17339);
nor U20294 (N_20294,N_15174,N_15169);
nand U20295 (N_20295,N_17552,N_15607);
or U20296 (N_20296,N_16610,N_17368);
and U20297 (N_20297,N_15606,N_15682);
or U20298 (N_20298,N_17604,N_16097);
nor U20299 (N_20299,N_17164,N_15814);
or U20300 (N_20300,N_17960,N_17785);
and U20301 (N_20301,N_15649,N_16347);
nor U20302 (N_20302,N_16931,N_17730);
nand U20303 (N_20303,N_17576,N_16624);
nand U20304 (N_20304,N_16109,N_16511);
or U20305 (N_20305,N_16800,N_15832);
and U20306 (N_20306,N_15451,N_16194);
nand U20307 (N_20307,N_16096,N_15899);
and U20308 (N_20308,N_15619,N_17315);
or U20309 (N_20309,N_15725,N_15670);
or U20310 (N_20310,N_15912,N_16223);
or U20311 (N_20311,N_17136,N_17398);
nand U20312 (N_20312,N_16141,N_17010);
and U20313 (N_20313,N_17077,N_17840);
or U20314 (N_20314,N_15807,N_15625);
xor U20315 (N_20315,N_15637,N_17862);
nor U20316 (N_20316,N_15526,N_15375);
nand U20317 (N_20317,N_16441,N_17151);
or U20318 (N_20318,N_17328,N_16182);
and U20319 (N_20319,N_16439,N_15867);
and U20320 (N_20320,N_17075,N_15538);
or U20321 (N_20321,N_15958,N_17270);
nor U20322 (N_20322,N_15552,N_15627);
nor U20323 (N_20323,N_17298,N_17306);
nand U20324 (N_20324,N_15388,N_17211);
nor U20325 (N_20325,N_15387,N_16712);
nand U20326 (N_20326,N_17077,N_15837);
nand U20327 (N_20327,N_17088,N_16726);
xor U20328 (N_20328,N_16242,N_15123);
nor U20329 (N_20329,N_17409,N_17604);
nand U20330 (N_20330,N_17164,N_15418);
nand U20331 (N_20331,N_15359,N_17269);
nand U20332 (N_20332,N_15544,N_17497);
and U20333 (N_20333,N_16526,N_15311);
nand U20334 (N_20334,N_17730,N_15572);
or U20335 (N_20335,N_17834,N_15295);
or U20336 (N_20336,N_16467,N_16687);
nand U20337 (N_20337,N_16751,N_15778);
or U20338 (N_20338,N_17825,N_17499);
nor U20339 (N_20339,N_15883,N_15618);
nand U20340 (N_20340,N_17507,N_16839);
nand U20341 (N_20341,N_16909,N_16015);
and U20342 (N_20342,N_17270,N_16795);
and U20343 (N_20343,N_15763,N_15809);
or U20344 (N_20344,N_17252,N_17240);
xor U20345 (N_20345,N_17506,N_16163);
and U20346 (N_20346,N_17449,N_17279);
xor U20347 (N_20347,N_16515,N_15090);
nand U20348 (N_20348,N_16252,N_15516);
and U20349 (N_20349,N_17552,N_15990);
nor U20350 (N_20350,N_16576,N_17764);
or U20351 (N_20351,N_17417,N_15363);
and U20352 (N_20352,N_15612,N_17469);
and U20353 (N_20353,N_15766,N_16175);
xor U20354 (N_20354,N_16853,N_15141);
or U20355 (N_20355,N_16952,N_15722);
and U20356 (N_20356,N_16545,N_16847);
or U20357 (N_20357,N_17539,N_15655);
nor U20358 (N_20358,N_17655,N_16373);
nor U20359 (N_20359,N_15944,N_16127);
and U20360 (N_20360,N_15115,N_17754);
xor U20361 (N_20361,N_15175,N_15511);
or U20362 (N_20362,N_16214,N_15112);
nand U20363 (N_20363,N_15129,N_17671);
xor U20364 (N_20364,N_16403,N_16731);
and U20365 (N_20365,N_15231,N_17248);
nor U20366 (N_20366,N_16769,N_15626);
xnor U20367 (N_20367,N_17667,N_15740);
nand U20368 (N_20368,N_16178,N_17301);
or U20369 (N_20369,N_17724,N_17554);
xnor U20370 (N_20370,N_16856,N_16698);
xor U20371 (N_20371,N_17379,N_17639);
nand U20372 (N_20372,N_17696,N_17741);
or U20373 (N_20373,N_17775,N_17139);
or U20374 (N_20374,N_17218,N_17512);
and U20375 (N_20375,N_17838,N_17089);
and U20376 (N_20376,N_15766,N_17637);
or U20377 (N_20377,N_17152,N_17995);
or U20378 (N_20378,N_17832,N_15295);
and U20379 (N_20379,N_15778,N_16136);
xor U20380 (N_20380,N_17860,N_16391);
or U20381 (N_20381,N_16287,N_16647);
nand U20382 (N_20382,N_15019,N_17968);
nand U20383 (N_20383,N_15643,N_15122);
and U20384 (N_20384,N_17912,N_17587);
nor U20385 (N_20385,N_16352,N_17966);
or U20386 (N_20386,N_16731,N_17609);
xnor U20387 (N_20387,N_16861,N_15489);
or U20388 (N_20388,N_15934,N_15671);
nor U20389 (N_20389,N_15172,N_16255);
nor U20390 (N_20390,N_17704,N_15861);
and U20391 (N_20391,N_17327,N_15856);
nand U20392 (N_20392,N_15536,N_15193);
nand U20393 (N_20393,N_15619,N_17515);
nand U20394 (N_20394,N_17218,N_17555);
or U20395 (N_20395,N_16765,N_16307);
or U20396 (N_20396,N_16335,N_16545);
and U20397 (N_20397,N_17916,N_16826);
nor U20398 (N_20398,N_15789,N_17996);
xnor U20399 (N_20399,N_16336,N_17089);
nor U20400 (N_20400,N_17246,N_17335);
nor U20401 (N_20401,N_17776,N_16394);
and U20402 (N_20402,N_17071,N_16031);
nor U20403 (N_20403,N_17323,N_17676);
nor U20404 (N_20404,N_17789,N_16862);
xor U20405 (N_20405,N_15043,N_16465);
xnor U20406 (N_20406,N_15496,N_16222);
or U20407 (N_20407,N_15580,N_17979);
and U20408 (N_20408,N_15904,N_16838);
nand U20409 (N_20409,N_15951,N_15078);
nand U20410 (N_20410,N_15492,N_15251);
nor U20411 (N_20411,N_16717,N_15450);
nand U20412 (N_20412,N_16455,N_17669);
nor U20413 (N_20413,N_15885,N_15867);
and U20414 (N_20414,N_15983,N_17269);
xnor U20415 (N_20415,N_17239,N_16059);
xor U20416 (N_20416,N_15135,N_15844);
nor U20417 (N_20417,N_16954,N_15860);
nor U20418 (N_20418,N_16292,N_17658);
xnor U20419 (N_20419,N_15599,N_15996);
and U20420 (N_20420,N_17008,N_17254);
or U20421 (N_20421,N_16440,N_17381);
nand U20422 (N_20422,N_16657,N_15049);
xor U20423 (N_20423,N_15932,N_16709);
xor U20424 (N_20424,N_17257,N_15163);
xnor U20425 (N_20425,N_17699,N_16051);
nand U20426 (N_20426,N_15700,N_17469);
xor U20427 (N_20427,N_17845,N_16993);
and U20428 (N_20428,N_15464,N_17329);
nor U20429 (N_20429,N_16369,N_16466);
nand U20430 (N_20430,N_17378,N_15949);
nand U20431 (N_20431,N_16958,N_16269);
nor U20432 (N_20432,N_16600,N_15008);
xnor U20433 (N_20433,N_15067,N_17574);
nor U20434 (N_20434,N_15289,N_15377);
or U20435 (N_20435,N_15445,N_15852);
nor U20436 (N_20436,N_15723,N_16843);
nand U20437 (N_20437,N_17877,N_16947);
and U20438 (N_20438,N_16060,N_16309);
nor U20439 (N_20439,N_17800,N_17850);
xor U20440 (N_20440,N_17266,N_17671);
or U20441 (N_20441,N_15607,N_16209);
nor U20442 (N_20442,N_15427,N_16069);
and U20443 (N_20443,N_17335,N_15210);
nor U20444 (N_20444,N_17339,N_17206);
nor U20445 (N_20445,N_15211,N_16840);
xor U20446 (N_20446,N_15086,N_15584);
nor U20447 (N_20447,N_17221,N_15481);
or U20448 (N_20448,N_15926,N_17449);
and U20449 (N_20449,N_16462,N_16434);
xor U20450 (N_20450,N_15874,N_17172);
or U20451 (N_20451,N_16529,N_17594);
nand U20452 (N_20452,N_16252,N_15587);
xor U20453 (N_20453,N_15890,N_17914);
nor U20454 (N_20454,N_15813,N_17353);
nor U20455 (N_20455,N_17459,N_15323);
nand U20456 (N_20456,N_15419,N_17226);
xnor U20457 (N_20457,N_16531,N_15833);
or U20458 (N_20458,N_16508,N_17113);
or U20459 (N_20459,N_17156,N_17169);
and U20460 (N_20460,N_17283,N_16746);
nor U20461 (N_20461,N_15010,N_17255);
or U20462 (N_20462,N_17053,N_17333);
or U20463 (N_20463,N_16852,N_15706);
xnor U20464 (N_20464,N_15130,N_16516);
nand U20465 (N_20465,N_15801,N_16294);
nor U20466 (N_20466,N_17951,N_15512);
nand U20467 (N_20467,N_15807,N_15184);
nor U20468 (N_20468,N_15802,N_17180);
and U20469 (N_20469,N_16304,N_16909);
xor U20470 (N_20470,N_15301,N_16440);
nor U20471 (N_20471,N_15511,N_15810);
xor U20472 (N_20472,N_16406,N_17380);
nand U20473 (N_20473,N_15485,N_15617);
and U20474 (N_20474,N_17238,N_15955);
nand U20475 (N_20475,N_17381,N_15656);
nor U20476 (N_20476,N_17598,N_15101);
nand U20477 (N_20477,N_15807,N_17823);
and U20478 (N_20478,N_17420,N_15700);
xnor U20479 (N_20479,N_16133,N_17031);
nor U20480 (N_20480,N_17836,N_16762);
or U20481 (N_20481,N_15439,N_15062);
nand U20482 (N_20482,N_15230,N_15380);
xnor U20483 (N_20483,N_15257,N_17889);
nor U20484 (N_20484,N_17905,N_16744);
nor U20485 (N_20485,N_16550,N_17690);
or U20486 (N_20486,N_16675,N_16884);
nor U20487 (N_20487,N_17566,N_17059);
and U20488 (N_20488,N_15898,N_17720);
nand U20489 (N_20489,N_17112,N_15858);
and U20490 (N_20490,N_17170,N_16785);
nand U20491 (N_20491,N_15356,N_16710);
or U20492 (N_20492,N_15130,N_16898);
and U20493 (N_20493,N_16663,N_16648);
or U20494 (N_20494,N_15769,N_16676);
and U20495 (N_20495,N_15909,N_15248);
nand U20496 (N_20496,N_16412,N_16601);
xor U20497 (N_20497,N_17758,N_16710);
nand U20498 (N_20498,N_17336,N_17630);
or U20499 (N_20499,N_15774,N_16379);
nor U20500 (N_20500,N_16324,N_17854);
and U20501 (N_20501,N_17875,N_17519);
nor U20502 (N_20502,N_16366,N_17973);
xor U20503 (N_20503,N_16792,N_17314);
and U20504 (N_20504,N_17457,N_15323);
and U20505 (N_20505,N_17155,N_16596);
nand U20506 (N_20506,N_16744,N_17961);
and U20507 (N_20507,N_16314,N_16358);
nand U20508 (N_20508,N_15697,N_15894);
nor U20509 (N_20509,N_15628,N_15362);
or U20510 (N_20510,N_16843,N_15813);
or U20511 (N_20511,N_17345,N_15250);
and U20512 (N_20512,N_15729,N_17942);
nor U20513 (N_20513,N_16183,N_17984);
xor U20514 (N_20514,N_15578,N_17883);
nand U20515 (N_20515,N_17796,N_17770);
or U20516 (N_20516,N_17137,N_16491);
or U20517 (N_20517,N_17657,N_15454);
or U20518 (N_20518,N_16084,N_17459);
and U20519 (N_20519,N_16889,N_16227);
or U20520 (N_20520,N_17102,N_17773);
nand U20521 (N_20521,N_15201,N_15148);
and U20522 (N_20522,N_17388,N_17142);
xnor U20523 (N_20523,N_17196,N_17825);
nand U20524 (N_20524,N_16749,N_15549);
or U20525 (N_20525,N_17546,N_15290);
nand U20526 (N_20526,N_17746,N_16096);
nand U20527 (N_20527,N_16271,N_17347);
nor U20528 (N_20528,N_17133,N_15372);
or U20529 (N_20529,N_16342,N_16184);
or U20530 (N_20530,N_17718,N_16963);
nand U20531 (N_20531,N_17682,N_16936);
nor U20532 (N_20532,N_15075,N_17278);
xnor U20533 (N_20533,N_15228,N_16928);
or U20534 (N_20534,N_15201,N_17591);
nand U20535 (N_20535,N_16774,N_16541);
and U20536 (N_20536,N_15648,N_16252);
nand U20537 (N_20537,N_17518,N_16251);
xor U20538 (N_20538,N_16309,N_16646);
and U20539 (N_20539,N_15767,N_16083);
and U20540 (N_20540,N_17642,N_15153);
nand U20541 (N_20541,N_15390,N_16030);
and U20542 (N_20542,N_16569,N_17376);
nor U20543 (N_20543,N_16288,N_17440);
or U20544 (N_20544,N_15748,N_16908);
nand U20545 (N_20545,N_15402,N_17697);
nor U20546 (N_20546,N_15038,N_17178);
nand U20547 (N_20547,N_15661,N_16998);
nor U20548 (N_20548,N_17488,N_17561);
xnor U20549 (N_20549,N_16816,N_16911);
and U20550 (N_20550,N_15823,N_15409);
nor U20551 (N_20551,N_16968,N_15031);
and U20552 (N_20552,N_15327,N_16264);
nor U20553 (N_20553,N_16056,N_16408);
and U20554 (N_20554,N_17724,N_16357);
nand U20555 (N_20555,N_17669,N_16300);
or U20556 (N_20556,N_15889,N_17440);
xnor U20557 (N_20557,N_17858,N_15222);
xor U20558 (N_20558,N_17983,N_15155);
nor U20559 (N_20559,N_16941,N_15334);
or U20560 (N_20560,N_15923,N_15855);
and U20561 (N_20561,N_17806,N_17525);
or U20562 (N_20562,N_16435,N_16689);
or U20563 (N_20563,N_16337,N_17894);
xnor U20564 (N_20564,N_17516,N_16312);
and U20565 (N_20565,N_17321,N_17929);
xor U20566 (N_20566,N_15833,N_16486);
nand U20567 (N_20567,N_17325,N_15696);
or U20568 (N_20568,N_15268,N_15324);
and U20569 (N_20569,N_17291,N_15782);
nor U20570 (N_20570,N_15508,N_17134);
nor U20571 (N_20571,N_16647,N_17882);
nor U20572 (N_20572,N_15880,N_15362);
nor U20573 (N_20573,N_16267,N_15649);
nand U20574 (N_20574,N_15961,N_16008);
and U20575 (N_20575,N_15304,N_15257);
and U20576 (N_20576,N_15329,N_17808);
nor U20577 (N_20577,N_16815,N_15805);
nand U20578 (N_20578,N_15970,N_15725);
nand U20579 (N_20579,N_15175,N_17283);
nand U20580 (N_20580,N_17455,N_16620);
or U20581 (N_20581,N_17041,N_17649);
nand U20582 (N_20582,N_17595,N_16958);
nand U20583 (N_20583,N_17161,N_15881);
xnor U20584 (N_20584,N_17537,N_16469);
nor U20585 (N_20585,N_15349,N_16562);
xnor U20586 (N_20586,N_16235,N_17715);
xnor U20587 (N_20587,N_16064,N_16598);
or U20588 (N_20588,N_15256,N_16270);
or U20589 (N_20589,N_17183,N_16386);
and U20590 (N_20590,N_16157,N_16018);
xor U20591 (N_20591,N_15616,N_17335);
or U20592 (N_20592,N_15865,N_17784);
nand U20593 (N_20593,N_16707,N_17153);
nor U20594 (N_20594,N_16375,N_15016);
and U20595 (N_20595,N_17137,N_15371);
xnor U20596 (N_20596,N_17927,N_17708);
xnor U20597 (N_20597,N_17646,N_16178);
nor U20598 (N_20598,N_17291,N_15948);
or U20599 (N_20599,N_17110,N_15915);
or U20600 (N_20600,N_16541,N_15792);
and U20601 (N_20601,N_15351,N_16269);
nor U20602 (N_20602,N_17065,N_15599);
or U20603 (N_20603,N_16744,N_15982);
xnor U20604 (N_20604,N_15693,N_16666);
or U20605 (N_20605,N_16064,N_16230);
nor U20606 (N_20606,N_17140,N_15095);
or U20607 (N_20607,N_17091,N_17033);
or U20608 (N_20608,N_17300,N_15225);
nand U20609 (N_20609,N_15104,N_16504);
nor U20610 (N_20610,N_15509,N_16373);
xnor U20611 (N_20611,N_16433,N_16662);
or U20612 (N_20612,N_16972,N_17841);
nand U20613 (N_20613,N_16839,N_15317);
nor U20614 (N_20614,N_15343,N_17008);
nand U20615 (N_20615,N_15862,N_17352);
xor U20616 (N_20616,N_16599,N_17397);
nand U20617 (N_20617,N_17698,N_15839);
and U20618 (N_20618,N_15040,N_17422);
nand U20619 (N_20619,N_15214,N_15821);
nor U20620 (N_20620,N_16425,N_16566);
xnor U20621 (N_20621,N_16126,N_15770);
nand U20622 (N_20622,N_16136,N_15611);
and U20623 (N_20623,N_16219,N_17534);
or U20624 (N_20624,N_15536,N_15023);
xor U20625 (N_20625,N_17907,N_16416);
or U20626 (N_20626,N_16713,N_15379);
nand U20627 (N_20627,N_16519,N_17506);
nor U20628 (N_20628,N_17813,N_16222);
xor U20629 (N_20629,N_16263,N_16395);
or U20630 (N_20630,N_17286,N_15047);
nand U20631 (N_20631,N_16070,N_16883);
or U20632 (N_20632,N_15594,N_15928);
nor U20633 (N_20633,N_16251,N_15026);
and U20634 (N_20634,N_17706,N_16286);
xor U20635 (N_20635,N_16431,N_15535);
nand U20636 (N_20636,N_16095,N_17255);
nand U20637 (N_20637,N_16621,N_17845);
or U20638 (N_20638,N_16866,N_16573);
and U20639 (N_20639,N_16635,N_17199);
or U20640 (N_20640,N_17030,N_17913);
and U20641 (N_20641,N_17272,N_15840);
or U20642 (N_20642,N_16802,N_16872);
or U20643 (N_20643,N_15523,N_16477);
xnor U20644 (N_20644,N_15400,N_15803);
and U20645 (N_20645,N_16836,N_17875);
xor U20646 (N_20646,N_16377,N_16493);
nor U20647 (N_20647,N_15982,N_16248);
nor U20648 (N_20648,N_15094,N_17848);
nor U20649 (N_20649,N_15810,N_15199);
or U20650 (N_20650,N_16975,N_15364);
nand U20651 (N_20651,N_16536,N_16396);
and U20652 (N_20652,N_15412,N_17681);
xor U20653 (N_20653,N_16905,N_15567);
nand U20654 (N_20654,N_15871,N_17515);
xor U20655 (N_20655,N_17538,N_15308);
nor U20656 (N_20656,N_17564,N_15807);
nor U20657 (N_20657,N_16767,N_17889);
xnor U20658 (N_20658,N_17890,N_17888);
xnor U20659 (N_20659,N_17438,N_16664);
xnor U20660 (N_20660,N_17211,N_15389);
nand U20661 (N_20661,N_15608,N_17945);
and U20662 (N_20662,N_16675,N_16326);
xnor U20663 (N_20663,N_15239,N_16500);
nand U20664 (N_20664,N_15060,N_17481);
nor U20665 (N_20665,N_16870,N_16618);
nand U20666 (N_20666,N_15728,N_17693);
nor U20667 (N_20667,N_16607,N_15571);
xor U20668 (N_20668,N_16491,N_16709);
xor U20669 (N_20669,N_15293,N_17730);
or U20670 (N_20670,N_17211,N_15560);
xnor U20671 (N_20671,N_15322,N_16106);
nand U20672 (N_20672,N_17296,N_17858);
nor U20673 (N_20673,N_17263,N_17410);
or U20674 (N_20674,N_17358,N_15275);
and U20675 (N_20675,N_16794,N_16940);
nor U20676 (N_20676,N_15532,N_17630);
xnor U20677 (N_20677,N_15235,N_17689);
or U20678 (N_20678,N_17331,N_17586);
or U20679 (N_20679,N_17990,N_16934);
and U20680 (N_20680,N_15269,N_16945);
xor U20681 (N_20681,N_17179,N_17270);
or U20682 (N_20682,N_16230,N_15734);
nor U20683 (N_20683,N_15656,N_17242);
nor U20684 (N_20684,N_17405,N_16926);
and U20685 (N_20685,N_15692,N_17075);
xnor U20686 (N_20686,N_15301,N_16875);
nand U20687 (N_20687,N_15478,N_17105);
nand U20688 (N_20688,N_15297,N_17016);
nor U20689 (N_20689,N_15721,N_16401);
nor U20690 (N_20690,N_15778,N_17677);
nor U20691 (N_20691,N_15981,N_15788);
nor U20692 (N_20692,N_17772,N_16550);
xor U20693 (N_20693,N_17583,N_17444);
xnor U20694 (N_20694,N_15450,N_16416);
or U20695 (N_20695,N_16036,N_17051);
or U20696 (N_20696,N_17068,N_17830);
and U20697 (N_20697,N_17981,N_17218);
xnor U20698 (N_20698,N_16895,N_16776);
or U20699 (N_20699,N_15534,N_16298);
or U20700 (N_20700,N_15583,N_15144);
nor U20701 (N_20701,N_17599,N_17462);
nand U20702 (N_20702,N_16385,N_17851);
nand U20703 (N_20703,N_16412,N_16888);
xnor U20704 (N_20704,N_17550,N_16588);
and U20705 (N_20705,N_16520,N_15027);
nand U20706 (N_20706,N_16671,N_16992);
nor U20707 (N_20707,N_15826,N_17386);
or U20708 (N_20708,N_15020,N_17285);
or U20709 (N_20709,N_16563,N_17677);
xor U20710 (N_20710,N_17753,N_15454);
and U20711 (N_20711,N_17371,N_15252);
or U20712 (N_20712,N_15193,N_16948);
xor U20713 (N_20713,N_16485,N_15877);
nand U20714 (N_20714,N_15838,N_15225);
nand U20715 (N_20715,N_16639,N_16513);
or U20716 (N_20716,N_15330,N_17540);
or U20717 (N_20717,N_15938,N_17412);
and U20718 (N_20718,N_17321,N_16117);
nor U20719 (N_20719,N_15042,N_16187);
nor U20720 (N_20720,N_16460,N_17391);
xor U20721 (N_20721,N_16471,N_17603);
nor U20722 (N_20722,N_15838,N_15327);
xnor U20723 (N_20723,N_16947,N_16656);
nor U20724 (N_20724,N_15866,N_16385);
and U20725 (N_20725,N_17591,N_17819);
nand U20726 (N_20726,N_16781,N_17514);
xor U20727 (N_20727,N_17692,N_16233);
xor U20728 (N_20728,N_15877,N_15690);
nand U20729 (N_20729,N_15115,N_15261);
nand U20730 (N_20730,N_15067,N_15423);
xnor U20731 (N_20731,N_15609,N_17663);
xor U20732 (N_20732,N_16852,N_15254);
xnor U20733 (N_20733,N_15940,N_15787);
xnor U20734 (N_20734,N_17216,N_17634);
nor U20735 (N_20735,N_16039,N_17630);
xor U20736 (N_20736,N_16216,N_15379);
or U20737 (N_20737,N_16054,N_17644);
nor U20738 (N_20738,N_17940,N_17520);
nor U20739 (N_20739,N_15394,N_17641);
nand U20740 (N_20740,N_15406,N_17943);
and U20741 (N_20741,N_17303,N_16017);
and U20742 (N_20742,N_17576,N_16229);
and U20743 (N_20743,N_17277,N_16055);
xnor U20744 (N_20744,N_15634,N_15613);
or U20745 (N_20745,N_15450,N_16906);
and U20746 (N_20746,N_15627,N_15169);
nand U20747 (N_20747,N_17242,N_16932);
nand U20748 (N_20748,N_15229,N_16317);
nor U20749 (N_20749,N_17497,N_16560);
and U20750 (N_20750,N_15590,N_15128);
or U20751 (N_20751,N_16154,N_15975);
xnor U20752 (N_20752,N_16103,N_16173);
nand U20753 (N_20753,N_16740,N_17016);
or U20754 (N_20754,N_16405,N_16239);
nand U20755 (N_20755,N_17624,N_16820);
xor U20756 (N_20756,N_16708,N_16018);
nand U20757 (N_20757,N_16820,N_16903);
nor U20758 (N_20758,N_17581,N_16048);
and U20759 (N_20759,N_15587,N_16621);
and U20760 (N_20760,N_15813,N_16875);
nand U20761 (N_20761,N_17462,N_15224);
nor U20762 (N_20762,N_17721,N_16255);
and U20763 (N_20763,N_16024,N_16906);
nand U20764 (N_20764,N_17600,N_15049);
xnor U20765 (N_20765,N_15424,N_16799);
xnor U20766 (N_20766,N_17547,N_16662);
and U20767 (N_20767,N_17206,N_15905);
nor U20768 (N_20768,N_16159,N_17204);
or U20769 (N_20769,N_15460,N_16124);
nor U20770 (N_20770,N_16175,N_17753);
and U20771 (N_20771,N_17537,N_17206);
nand U20772 (N_20772,N_16354,N_16524);
xnor U20773 (N_20773,N_17660,N_17520);
xnor U20774 (N_20774,N_15374,N_15306);
or U20775 (N_20775,N_17245,N_16201);
and U20776 (N_20776,N_16918,N_15139);
xor U20777 (N_20777,N_17553,N_16032);
and U20778 (N_20778,N_16393,N_15797);
nor U20779 (N_20779,N_16529,N_17674);
or U20780 (N_20780,N_17137,N_15000);
or U20781 (N_20781,N_15360,N_16934);
nor U20782 (N_20782,N_16850,N_15417);
and U20783 (N_20783,N_16191,N_16264);
nand U20784 (N_20784,N_16294,N_15891);
nand U20785 (N_20785,N_17913,N_15949);
and U20786 (N_20786,N_15829,N_17567);
nand U20787 (N_20787,N_15821,N_15976);
xnor U20788 (N_20788,N_15294,N_17929);
xor U20789 (N_20789,N_16285,N_15683);
nor U20790 (N_20790,N_17598,N_17722);
and U20791 (N_20791,N_15672,N_15674);
and U20792 (N_20792,N_16759,N_15614);
nor U20793 (N_20793,N_17520,N_15795);
xnor U20794 (N_20794,N_16425,N_15263);
or U20795 (N_20795,N_17773,N_15975);
nand U20796 (N_20796,N_16998,N_17395);
nor U20797 (N_20797,N_15068,N_15625);
or U20798 (N_20798,N_16996,N_16366);
nor U20799 (N_20799,N_17752,N_17632);
and U20800 (N_20800,N_17901,N_15788);
or U20801 (N_20801,N_16987,N_15172);
and U20802 (N_20802,N_15308,N_15936);
nor U20803 (N_20803,N_17547,N_15727);
and U20804 (N_20804,N_16958,N_16132);
and U20805 (N_20805,N_17560,N_17328);
or U20806 (N_20806,N_17663,N_15440);
xnor U20807 (N_20807,N_15042,N_17930);
nand U20808 (N_20808,N_16945,N_15706);
nor U20809 (N_20809,N_17107,N_15490);
and U20810 (N_20810,N_16301,N_16453);
or U20811 (N_20811,N_17540,N_17609);
xnor U20812 (N_20812,N_16532,N_16440);
nor U20813 (N_20813,N_15626,N_15037);
nor U20814 (N_20814,N_16322,N_17724);
nor U20815 (N_20815,N_15213,N_15884);
or U20816 (N_20816,N_17600,N_17219);
nor U20817 (N_20817,N_16540,N_15716);
xor U20818 (N_20818,N_16461,N_15787);
xnor U20819 (N_20819,N_15142,N_17485);
nand U20820 (N_20820,N_16705,N_16228);
xnor U20821 (N_20821,N_17894,N_15072);
nand U20822 (N_20822,N_17417,N_15532);
and U20823 (N_20823,N_15194,N_16921);
or U20824 (N_20824,N_17373,N_17480);
nor U20825 (N_20825,N_16723,N_15903);
and U20826 (N_20826,N_15709,N_15621);
nand U20827 (N_20827,N_16858,N_15706);
and U20828 (N_20828,N_16804,N_15295);
nand U20829 (N_20829,N_17036,N_17338);
nand U20830 (N_20830,N_16153,N_15424);
nand U20831 (N_20831,N_16251,N_17920);
xnor U20832 (N_20832,N_16061,N_16356);
or U20833 (N_20833,N_15599,N_17982);
or U20834 (N_20834,N_16775,N_16258);
and U20835 (N_20835,N_15641,N_15224);
nor U20836 (N_20836,N_15500,N_17879);
nor U20837 (N_20837,N_15392,N_17807);
or U20838 (N_20838,N_17207,N_15393);
or U20839 (N_20839,N_17737,N_15430);
xor U20840 (N_20840,N_17173,N_17822);
and U20841 (N_20841,N_15632,N_16632);
nor U20842 (N_20842,N_15348,N_17377);
nand U20843 (N_20843,N_17988,N_17845);
xnor U20844 (N_20844,N_15694,N_17967);
and U20845 (N_20845,N_16037,N_16701);
and U20846 (N_20846,N_16986,N_16777);
and U20847 (N_20847,N_17216,N_16842);
nand U20848 (N_20848,N_17461,N_17026);
nor U20849 (N_20849,N_16511,N_17566);
or U20850 (N_20850,N_16620,N_17958);
or U20851 (N_20851,N_15891,N_15307);
and U20852 (N_20852,N_17560,N_16000);
nor U20853 (N_20853,N_16077,N_16070);
xnor U20854 (N_20854,N_17058,N_16547);
nor U20855 (N_20855,N_15094,N_15012);
and U20856 (N_20856,N_16850,N_15587);
or U20857 (N_20857,N_15303,N_15625);
nand U20858 (N_20858,N_17674,N_17959);
or U20859 (N_20859,N_15331,N_16925);
or U20860 (N_20860,N_17700,N_17320);
nor U20861 (N_20861,N_15880,N_17120);
nor U20862 (N_20862,N_16245,N_17895);
xnor U20863 (N_20863,N_16838,N_16252);
nand U20864 (N_20864,N_15065,N_15037);
xor U20865 (N_20865,N_16551,N_17551);
and U20866 (N_20866,N_17778,N_15975);
nor U20867 (N_20867,N_17820,N_17993);
xor U20868 (N_20868,N_17173,N_17539);
and U20869 (N_20869,N_16507,N_15277);
or U20870 (N_20870,N_17013,N_15428);
nand U20871 (N_20871,N_15953,N_16509);
nor U20872 (N_20872,N_15061,N_15185);
and U20873 (N_20873,N_15232,N_17371);
or U20874 (N_20874,N_17912,N_17814);
or U20875 (N_20875,N_17637,N_16278);
and U20876 (N_20876,N_17004,N_17416);
or U20877 (N_20877,N_15261,N_17569);
and U20878 (N_20878,N_16483,N_15551);
or U20879 (N_20879,N_16838,N_15329);
xor U20880 (N_20880,N_15265,N_17076);
and U20881 (N_20881,N_16984,N_15723);
and U20882 (N_20882,N_15066,N_17359);
and U20883 (N_20883,N_17597,N_15180);
nand U20884 (N_20884,N_16903,N_17838);
and U20885 (N_20885,N_17664,N_15152);
nor U20886 (N_20886,N_16886,N_16560);
nor U20887 (N_20887,N_16100,N_16293);
nand U20888 (N_20888,N_17650,N_16914);
or U20889 (N_20889,N_15141,N_16936);
or U20890 (N_20890,N_15900,N_17533);
nand U20891 (N_20891,N_16575,N_16612);
nor U20892 (N_20892,N_16834,N_16265);
nor U20893 (N_20893,N_15135,N_17500);
or U20894 (N_20894,N_15217,N_17322);
xnor U20895 (N_20895,N_15034,N_16691);
or U20896 (N_20896,N_15343,N_17607);
or U20897 (N_20897,N_16366,N_17232);
or U20898 (N_20898,N_15819,N_15612);
or U20899 (N_20899,N_15500,N_15394);
nor U20900 (N_20900,N_16147,N_15148);
xnor U20901 (N_20901,N_16013,N_16618);
nor U20902 (N_20902,N_16905,N_16142);
and U20903 (N_20903,N_17905,N_17292);
nand U20904 (N_20904,N_16799,N_15666);
and U20905 (N_20905,N_15767,N_17026);
xor U20906 (N_20906,N_16377,N_15670);
nor U20907 (N_20907,N_17499,N_17207);
nor U20908 (N_20908,N_16762,N_15089);
nor U20909 (N_20909,N_16220,N_17982);
xor U20910 (N_20910,N_17835,N_16697);
nand U20911 (N_20911,N_15557,N_15748);
nor U20912 (N_20912,N_17691,N_15531);
or U20913 (N_20913,N_16553,N_16512);
and U20914 (N_20914,N_16983,N_17002);
nor U20915 (N_20915,N_17175,N_16367);
xnor U20916 (N_20916,N_17179,N_15094);
xor U20917 (N_20917,N_17073,N_17491);
and U20918 (N_20918,N_17802,N_16517);
nor U20919 (N_20919,N_17931,N_16588);
and U20920 (N_20920,N_17072,N_17364);
or U20921 (N_20921,N_15810,N_16605);
or U20922 (N_20922,N_15461,N_16018);
xnor U20923 (N_20923,N_15602,N_17157);
or U20924 (N_20924,N_16452,N_17427);
xnor U20925 (N_20925,N_17558,N_15196);
or U20926 (N_20926,N_15876,N_16290);
and U20927 (N_20927,N_16282,N_16460);
xnor U20928 (N_20928,N_15934,N_17678);
and U20929 (N_20929,N_15984,N_17047);
xnor U20930 (N_20930,N_17859,N_15427);
and U20931 (N_20931,N_15169,N_16001);
nand U20932 (N_20932,N_15242,N_16572);
and U20933 (N_20933,N_15818,N_15236);
and U20934 (N_20934,N_16918,N_15224);
and U20935 (N_20935,N_17002,N_16411);
nand U20936 (N_20936,N_16941,N_16108);
xor U20937 (N_20937,N_15704,N_16869);
xor U20938 (N_20938,N_16249,N_15037);
or U20939 (N_20939,N_17507,N_16921);
nor U20940 (N_20940,N_16882,N_17093);
xor U20941 (N_20941,N_15597,N_17619);
or U20942 (N_20942,N_16250,N_16990);
and U20943 (N_20943,N_16190,N_15259);
and U20944 (N_20944,N_15271,N_17980);
and U20945 (N_20945,N_15336,N_17293);
nor U20946 (N_20946,N_17938,N_15540);
xnor U20947 (N_20947,N_16201,N_15425);
nor U20948 (N_20948,N_16543,N_16524);
nand U20949 (N_20949,N_17778,N_16330);
or U20950 (N_20950,N_16731,N_16525);
nand U20951 (N_20951,N_16220,N_15154);
nor U20952 (N_20952,N_17314,N_16598);
nor U20953 (N_20953,N_17967,N_17990);
and U20954 (N_20954,N_17703,N_15742);
nor U20955 (N_20955,N_16272,N_16629);
or U20956 (N_20956,N_16191,N_15840);
xnor U20957 (N_20957,N_15714,N_16801);
nor U20958 (N_20958,N_17445,N_16127);
and U20959 (N_20959,N_16718,N_15084);
and U20960 (N_20960,N_17422,N_16841);
xnor U20961 (N_20961,N_16310,N_16432);
nand U20962 (N_20962,N_16528,N_15633);
and U20963 (N_20963,N_16304,N_15636);
nand U20964 (N_20964,N_16541,N_17717);
nor U20965 (N_20965,N_15320,N_16886);
nand U20966 (N_20966,N_16953,N_15442);
and U20967 (N_20967,N_15831,N_15024);
xor U20968 (N_20968,N_16486,N_17715);
nand U20969 (N_20969,N_17532,N_17174);
xor U20970 (N_20970,N_17382,N_17803);
nand U20971 (N_20971,N_17943,N_16824);
and U20972 (N_20972,N_16770,N_16400);
and U20973 (N_20973,N_17247,N_16272);
nand U20974 (N_20974,N_16895,N_16162);
nor U20975 (N_20975,N_15037,N_17498);
or U20976 (N_20976,N_15134,N_16709);
xnor U20977 (N_20977,N_16840,N_15515);
and U20978 (N_20978,N_16152,N_15132);
nand U20979 (N_20979,N_17475,N_15323);
xor U20980 (N_20980,N_15969,N_16771);
and U20981 (N_20981,N_15345,N_16056);
and U20982 (N_20982,N_17978,N_17397);
and U20983 (N_20983,N_15654,N_16946);
or U20984 (N_20984,N_17332,N_15664);
and U20985 (N_20985,N_17667,N_15476);
and U20986 (N_20986,N_16557,N_16823);
nor U20987 (N_20987,N_17146,N_15799);
or U20988 (N_20988,N_15091,N_15298);
nand U20989 (N_20989,N_15857,N_16719);
and U20990 (N_20990,N_16048,N_16885);
xnor U20991 (N_20991,N_16786,N_17002);
nor U20992 (N_20992,N_15996,N_17539);
nor U20993 (N_20993,N_17704,N_15935);
xnor U20994 (N_20994,N_16909,N_17639);
nand U20995 (N_20995,N_17348,N_16460);
nand U20996 (N_20996,N_17538,N_17342);
or U20997 (N_20997,N_15925,N_17431);
or U20998 (N_20998,N_15954,N_17029);
nand U20999 (N_20999,N_16581,N_16024);
and U21000 (N_21000,N_20992,N_19858);
and U21001 (N_21001,N_20330,N_19358);
and U21002 (N_21002,N_19971,N_18823);
nor U21003 (N_21003,N_18311,N_20468);
or U21004 (N_21004,N_18180,N_18274);
and U21005 (N_21005,N_19616,N_19645);
xor U21006 (N_21006,N_20318,N_19700);
and U21007 (N_21007,N_19477,N_19376);
xnor U21008 (N_21008,N_20522,N_19984);
nor U21009 (N_21009,N_19032,N_18104);
or U21010 (N_21010,N_20551,N_18556);
or U21011 (N_21011,N_18866,N_18909);
nand U21012 (N_21012,N_19711,N_20579);
and U21013 (N_21013,N_18788,N_20740);
or U21014 (N_21014,N_18871,N_20609);
nand U21015 (N_21015,N_19588,N_19877);
nor U21016 (N_21016,N_18761,N_18613);
nand U21017 (N_21017,N_18949,N_20823);
nand U21018 (N_21018,N_18684,N_18365);
nand U21019 (N_21019,N_20366,N_18335);
or U21020 (N_21020,N_19391,N_18266);
nand U21021 (N_21021,N_19685,N_20126);
or U21022 (N_21022,N_18975,N_19139);
and U21023 (N_21023,N_18968,N_18345);
nor U21024 (N_21024,N_18994,N_20683);
nand U21025 (N_21025,N_20588,N_20103);
nand U21026 (N_21026,N_20674,N_18710);
xor U21027 (N_21027,N_20710,N_19874);
nand U21028 (N_21028,N_18867,N_18320);
or U21029 (N_21029,N_18955,N_19423);
nor U21030 (N_21030,N_20896,N_20585);
or U21031 (N_21031,N_19556,N_20036);
nor U21032 (N_21032,N_18562,N_18730);
or U21033 (N_21033,N_20263,N_19169);
or U21034 (N_21034,N_18037,N_20327);
or U21035 (N_21035,N_20183,N_19126);
or U21036 (N_21036,N_20933,N_20705);
nor U21037 (N_21037,N_18053,N_19405);
xor U21038 (N_21038,N_18649,N_18697);
and U21039 (N_21039,N_18681,N_18609);
and U21040 (N_21040,N_19441,N_19549);
nor U21041 (N_21041,N_19585,N_20688);
xor U21042 (N_21042,N_19676,N_20079);
nor U21043 (N_21043,N_18633,N_19909);
nand U21044 (N_21044,N_18476,N_19257);
nand U21045 (N_21045,N_20084,N_19418);
or U21046 (N_21046,N_18713,N_20008);
and U21047 (N_21047,N_20587,N_19193);
and U21048 (N_21048,N_20233,N_19394);
nor U21049 (N_21049,N_19857,N_20787);
nand U21050 (N_21050,N_19546,N_19946);
nand U21051 (N_21051,N_19173,N_18921);
xnor U21052 (N_21052,N_20730,N_19852);
xnor U21053 (N_21053,N_19657,N_19517);
nor U21054 (N_21054,N_19850,N_18386);
nor U21055 (N_21055,N_18007,N_18982);
nor U21056 (N_21056,N_20226,N_20068);
xnor U21057 (N_21057,N_20100,N_19849);
xnor U21058 (N_21058,N_18719,N_20241);
xnor U21059 (N_21059,N_19521,N_18227);
xor U21060 (N_21060,N_19188,N_19906);
or U21061 (N_21061,N_19410,N_19508);
nand U21062 (N_21062,N_20864,N_19045);
or U21063 (N_21063,N_18741,N_18243);
nor U21064 (N_21064,N_20876,N_20259);
and U21065 (N_21065,N_18069,N_20767);
and U21066 (N_21066,N_19213,N_18428);
xnor U21067 (N_21067,N_20108,N_18399);
nand U21068 (N_21068,N_19655,N_19631);
nor U21069 (N_21069,N_20088,N_20238);
or U21070 (N_21070,N_18256,N_18670);
and U21071 (N_21071,N_18603,N_19732);
and U21072 (N_21072,N_19002,N_19589);
and U21073 (N_21073,N_18144,N_19197);
nand U21074 (N_21074,N_20502,N_18917);
nand U21075 (N_21075,N_18686,N_20202);
and U21076 (N_21076,N_18179,N_20401);
nor U21077 (N_21077,N_18834,N_18152);
nor U21078 (N_21078,N_19966,N_18125);
or U21079 (N_21079,N_18403,N_20051);
nor U21080 (N_21080,N_18112,N_18291);
nor U21081 (N_21081,N_18383,N_19457);
and U21082 (N_21082,N_19958,N_20044);
and U21083 (N_21083,N_18624,N_20513);
or U21084 (N_21084,N_20148,N_20434);
nor U21085 (N_21085,N_18338,N_20707);
nand U21086 (N_21086,N_20806,N_19629);
nand U21087 (N_21087,N_20778,N_20793);
nor U21088 (N_21088,N_20632,N_18683);
nor U21089 (N_21089,N_19665,N_19342);
xor U21090 (N_21090,N_20696,N_18434);
nand U21091 (N_21091,N_19261,N_20189);
xnor U21092 (N_21092,N_18465,N_19602);
or U21093 (N_21093,N_20494,N_20299);
xnor U21094 (N_21094,N_19949,N_20016);
and U21095 (N_21095,N_18087,N_18279);
and U21096 (N_21096,N_19901,N_20005);
xor U21097 (N_21097,N_20677,N_19789);
and U21098 (N_21098,N_19177,N_20638);
nor U21099 (N_21099,N_20724,N_20165);
and U21100 (N_21100,N_20466,N_19472);
xor U21101 (N_21101,N_19619,N_19361);
nor U21102 (N_21102,N_20708,N_19747);
nand U21103 (N_21103,N_18899,N_18828);
nand U21104 (N_21104,N_20755,N_20412);
or U21105 (N_21105,N_18824,N_20244);
nor U21106 (N_21106,N_18288,N_20033);
and U21107 (N_21107,N_20023,N_20083);
nor U21108 (N_21108,N_19317,N_19401);
nand U21109 (N_21109,N_19708,N_19600);
or U21110 (N_21110,N_20130,N_18540);
nand U21111 (N_21111,N_19338,N_20795);
or U21112 (N_21112,N_18971,N_18737);
or U21113 (N_21113,N_19910,N_20133);
or U21114 (N_21114,N_20162,N_18767);
or U21115 (N_21115,N_19201,N_18582);
and U21116 (N_21116,N_20568,N_20610);
nor U21117 (N_21117,N_19328,N_18988);
nor U21118 (N_21118,N_18416,N_20996);
xor U21119 (N_21119,N_20671,N_19962);
nand U21120 (N_21120,N_20745,N_19027);
and U21121 (N_21121,N_18889,N_19437);
nand U21122 (N_21122,N_20704,N_18711);
nand U21123 (N_21123,N_20622,N_19968);
and U21124 (N_21124,N_18964,N_20865);
xor U21125 (N_21125,N_19648,N_19044);
nand U21126 (N_21126,N_18922,N_18211);
and U21127 (N_21127,N_19840,N_19351);
xnor U21128 (N_21128,N_20644,N_19478);
nand U21129 (N_21129,N_18723,N_18758);
nor U21130 (N_21130,N_18950,N_18046);
xor U21131 (N_21131,N_20075,N_20961);
nor U21132 (N_21132,N_18640,N_20972);
nand U21133 (N_21133,N_20628,N_19512);
and U21134 (N_21134,N_18090,N_19337);
or U21135 (N_21135,N_18530,N_19876);
nor U21136 (N_21136,N_19604,N_18265);
nand U21137 (N_21137,N_20091,N_20910);
nand U21138 (N_21138,N_19977,N_19621);
xor U21139 (N_21139,N_20209,N_18778);
nor U21140 (N_21140,N_18573,N_20408);
nor U21141 (N_21141,N_19241,N_19471);
nor U21142 (N_21142,N_19753,N_19015);
or U21143 (N_21143,N_20985,N_18371);
xor U21144 (N_21144,N_18825,N_18490);
and U21145 (N_21145,N_19729,N_19297);
nor U21146 (N_21146,N_20277,N_19536);
nand U21147 (N_21147,N_20321,N_19520);
nand U21148 (N_21148,N_18570,N_20890);
nand U21149 (N_21149,N_19101,N_20676);
and U21150 (N_21150,N_20111,N_19356);
and U21151 (N_21151,N_20934,N_18198);
or U21152 (N_21152,N_20930,N_19305);
nand U21153 (N_21153,N_19218,N_20403);
nand U21154 (N_21154,N_19454,N_20218);
nor U21155 (N_21155,N_19825,N_18143);
xnor U21156 (N_21156,N_20457,N_20771);
or U21157 (N_21157,N_20557,N_19581);
and U21158 (N_21158,N_20030,N_19097);
or U21159 (N_21159,N_18690,N_19082);
and U21160 (N_21160,N_19761,N_18716);
nor U21161 (N_21161,N_18468,N_19945);
or U21162 (N_21162,N_20558,N_18354);
xnor U21163 (N_21163,N_18580,N_18843);
xor U21164 (N_21164,N_18821,N_18896);
nand U21165 (N_21165,N_18021,N_20124);
nor U21166 (N_21166,N_20067,N_20645);
xor U21167 (N_21167,N_20143,N_19243);
xnor U21168 (N_21168,N_18389,N_18408);
and U21169 (N_21169,N_20839,N_20310);
nand U21170 (N_21170,N_19773,N_18261);
nand U21171 (N_21171,N_19499,N_20580);
and U21172 (N_21172,N_20820,N_20515);
and U21173 (N_21173,N_20946,N_19851);
nor U21174 (N_21174,N_20352,N_20990);
nor U21175 (N_21175,N_19598,N_19592);
xor U21176 (N_21176,N_19155,N_19688);
and U21177 (N_21177,N_20156,N_19274);
and U21178 (N_21178,N_20650,N_19768);
nor U21179 (N_21179,N_20373,N_18654);
and U21180 (N_21180,N_18248,N_20651);
xnor U21181 (N_21181,N_18531,N_19092);
or U21182 (N_21182,N_19004,N_20596);
xnor U21183 (N_21183,N_19972,N_18221);
nor U21184 (N_21184,N_19164,N_19555);
or U21185 (N_21185,N_18210,N_19653);
and U21186 (N_21186,N_18663,N_19845);
xnor U21187 (N_21187,N_19103,N_18860);
and U21188 (N_21188,N_19380,N_19625);
nor U21189 (N_21189,N_20922,N_19794);
xor U21190 (N_21190,N_20142,N_18606);
xnor U21191 (N_21191,N_18804,N_20526);
nor U21192 (N_21192,N_20102,N_18477);
and U21193 (N_21193,N_19883,N_18142);
nand U21194 (N_21194,N_18839,N_19231);
and U21195 (N_21195,N_20831,N_20007);
or U21196 (N_21196,N_20766,N_20739);
xnor U21197 (N_21197,N_19083,N_19371);
and U21198 (N_21198,N_18561,N_19805);
and U21199 (N_21199,N_19301,N_18067);
and U21200 (N_21200,N_19149,N_18492);
nor U21201 (N_21201,N_19759,N_18214);
nor U21202 (N_21202,N_18470,N_18138);
and U21203 (N_21203,N_20534,N_18308);
xnor U21204 (N_21204,N_19630,N_20355);
nor U21205 (N_21205,N_20786,N_19205);
nand U21206 (N_21206,N_19704,N_18615);
nand U21207 (N_21207,N_20128,N_19310);
or U21208 (N_21208,N_19063,N_19673);
or U21209 (N_21209,N_20022,N_20542);
or U21210 (N_21210,N_20032,N_20014);
nor U21211 (N_21211,N_18299,N_20278);
nor U21212 (N_21212,N_19220,N_19746);
or U21213 (N_21213,N_20019,N_20763);
nor U21214 (N_21214,N_20532,N_19727);
xnor U21215 (N_21215,N_19827,N_20090);
xnor U21216 (N_21216,N_18699,N_18424);
nor U21217 (N_21217,N_20061,N_18602);
and U21218 (N_21218,N_19889,N_18190);
and U21219 (N_21219,N_20120,N_20584);
nor U21220 (N_21220,N_18159,N_18727);
or U21221 (N_21221,N_18709,N_20488);
nor U21222 (N_21222,N_19530,N_19095);
nand U21223 (N_21223,N_20877,N_20448);
nand U21224 (N_21224,N_19160,N_20347);
nand U21225 (N_21225,N_20358,N_18344);
nand U21226 (N_21226,N_19576,N_20407);
and U21227 (N_21227,N_20040,N_18471);
nor U21228 (N_21228,N_18213,N_20811);
nor U21229 (N_21229,N_19465,N_19190);
xnor U21230 (N_21230,N_18063,N_20747);
nand U21231 (N_21231,N_20909,N_20926);
nor U21232 (N_21232,N_20641,N_19025);
xor U21233 (N_21233,N_20472,N_18966);
and U21234 (N_21234,N_20861,N_18521);
nor U21235 (N_21235,N_20335,N_20255);
xor U21236 (N_21236,N_20668,N_20132);
nor U21237 (N_21237,N_19677,N_20243);
nand U21238 (N_21238,N_18822,N_18870);
nand U21239 (N_21239,N_18297,N_19728);
or U21240 (N_21240,N_18194,N_19099);
or U21241 (N_21241,N_20733,N_20479);
xnor U21242 (N_21242,N_18566,N_20809);
nand U21243 (N_21243,N_19105,N_20665);
nor U21244 (N_21244,N_20283,N_20944);
xor U21245 (N_21245,N_18546,N_19931);
and U21246 (N_21246,N_18427,N_20734);
or U21247 (N_21247,N_20997,N_19395);
nor U21248 (N_21248,N_20198,N_18002);
and U21249 (N_21249,N_19841,N_19107);
and U21250 (N_21250,N_19667,N_19726);
xor U21251 (N_21251,N_19493,N_20791);
xnor U21252 (N_21252,N_20476,N_19771);
or U21253 (N_21253,N_19515,N_19758);
nor U21254 (N_21254,N_18293,N_18040);
or U21255 (N_21255,N_20147,N_19836);
xor U21256 (N_21256,N_18370,N_19679);
or U21257 (N_21257,N_18281,N_19007);
xnor U21258 (N_21258,N_19622,N_18442);
nand U21259 (N_21259,N_19871,N_19802);
and U21260 (N_21260,N_20919,N_18061);
xnor U21261 (N_21261,N_18278,N_18555);
nor U21262 (N_21262,N_20058,N_18880);
xnor U21263 (N_21263,N_19607,N_18722);
and U21264 (N_21264,N_20978,N_19223);
or U21265 (N_21265,N_19253,N_18548);
or U21266 (N_21266,N_19869,N_19661);
nand U21267 (N_21267,N_19703,N_19470);
nand U21268 (N_21268,N_19790,N_18932);
xnor U21269 (N_21269,N_20034,N_18268);
nand U21270 (N_21270,N_18323,N_19096);
nand U21271 (N_21271,N_19070,N_18844);
or U21272 (N_21272,N_20868,N_19683);
or U21273 (N_21273,N_19374,N_18944);
nand U21274 (N_21274,N_18739,N_18358);
nor U21275 (N_21275,N_20426,N_18850);
nand U21276 (N_21276,N_20372,N_20938);
and U21277 (N_21277,N_19541,N_19762);
xor U21278 (N_21278,N_20294,N_20658);
xnor U21279 (N_21279,N_18625,N_20582);
and U21280 (N_21280,N_20054,N_20554);
nor U21281 (N_21281,N_18914,N_19184);
and U21282 (N_21282,N_18036,N_19313);
or U21283 (N_21283,N_19449,N_18280);
nor U21284 (N_21284,N_19786,N_20150);
xor U21285 (N_21285,N_20474,N_18749);
or U21286 (N_21286,N_19343,N_20810);
nor U21287 (N_21287,N_20234,N_19999);
nand U21288 (N_21288,N_20105,N_18195);
nor U21289 (N_21289,N_19720,N_18042);
nand U21290 (N_21290,N_19228,N_19826);
or U21291 (N_21291,N_19719,N_19324);
nor U21292 (N_21292,N_19591,N_19733);
and U21293 (N_21293,N_20953,N_19506);
nor U21294 (N_21294,N_19050,N_18901);
and U21295 (N_21295,N_19658,N_20981);
and U21296 (N_21296,N_19800,N_19263);
nand U21297 (N_21297,N_20866,N_20043);
or U21298 (N_21298,N_20463,N_20828);
xnor U21299 (N_21299,N_18991,N_18894);
and U21300 (N_21300,N_20388,N_18564);
xor U21301 (N_21301,N_19247,N_20171);
and U21302 (N_21302,N_19964,N_18451);
xor U21303 (N_21303,N_20342,N_20576);
and U21304 (N_21304,N_18588,N_20237);
xnor U21305 (N_21305,N_18431,N_18970);
nor U21306 (N_21306,N_18551,N_18475);
or U21307 (N_21307,N_18731,N_20415);
nand U21308 (N_21308,N_19487,N_20959);
and U21309 (N_21309,N_20672,N_19976);
and U21310 (N_21310,N_19366,N_20287);
xnor U21311 (N_21311,N_18666,N_19141);
xor U21312 (N_21312,N_20550,N_18397);
or U21313 (N_21313,N_19666,N_19518);
nand U21314 (N_21314,N_18887,N_18908);
nand U21315 (N_21315,N_18937,N_18216);
or U21316 (N_21316,N_18237,N_20499);
nand U21317 (N_21317,N_18608,N_19340);
and U21318 (N_21318,N_18992,N_20138);
xnor U21319 (N_21319,N_18836,N_20948);
nand U21320 (N_21320,N_20569,N_20246);
xnor U21321 (N_21321,N_20304,N_18407);
nand U21322 (N_21322,N_20871,N_18435);
or U21323 (N_21323,N_20857,N_20652);
xor U21324 (N_21324,N_20444,N_18132);
nor U21325 (N_21325,N_20439,N_20637);
nor U21326 (N_21326,N_20935,N_19034);
and U21327 (N_21327,N_19059,N_19398);
nand U21328 (N_21328,N_19260,N_19567);
nand U21329 (N_21329,N_18811,N_18220);
or U21330 (N_21330,N_19792,N_20965);
or U21331 (N_21331,N_19076,N_19458);
or U21332 (N_21332,N_19387,N_19519);
xnor U21333 (N_21333,N_19580,N_19386);
nor U21334 (N_21334,N_18651,N_19156);
and U21335 (N_21335,N_20056,N_19887);
and U21336 (N_21336,N_19494,N_20521);
or U21337 (N_21337,N_19244,N_20958);
or U21338 (N_21338,N_20510,N_19364);
xor U21339 (N_21339,N_18618,N_20776);
nand U21340 (N_21340,N_20885,N_19068);
and U21341 (N_21341,N_18513,N_20364);
nand U21342 (N_21342,N_18322,N_18107);
nand U21343 (N_21343,N_19040,N_18498);
nor U21344 (N_21344,N_18733,N_18756);
or U21345 (N_21345,N_18328,N_20242);
nand U21346 (N_21346,N_20493,N_19230);
and U21347 (N_21347,N_20538,N_19955);
nor U21348 (N_21348,N_18361,N_20383);
xnor U21349 (N_21349,N_18100,N_19583);
and U21350 (N_21350,N_19372,N_18276);
nand U21351 (N_21351,N_19656,N_18604);
xor U21352 (N_21352,N_18306,N_19303);
or U21353 (N_21353,N_18832,N_20604);
nand U21354 (N_21354,N_20850,N_19250);
and U21355 (N_21355,N_20702,N_20615);
nand U21356 (N_21356,N_18350,N_18559);
nor U21357 (N_21357,N_19229,N_19293);
or U21358 (N_21358,N_20302,N_20594);
and U21359 (N_21359,N_18136,N_20492);
xor U21360 (N_21360,N_20451,N_18952);
xor U21361 (N_21361,N_19690,N_19533);
xor U21362 (N_21362,N_19705,N_20545);
or U21363 (N_21363,N_19060,N_18205);
and U21364 (N_21364,N_20858,N_18495);
nand U21365 (N_21365,N_20769,N_19785);
or U21366 (N_21366,N_20681,N_19782);
xor U21367 (N_21367,N_19818,N_19486);
nor U21368 (N_21368,N_19528,N_19145);
nor U21369 (N_21369,N_20331,N_19885);
and U21370 (N_21370,N_19638,N_19843);
and U21371 (N_21371,N_20151,N_18724);
nand U21372 (N_21372,N_19578,N_18990);
and U21373 (N_21373,N_18203,N_19422);
or U21374 (N_21374,N_18406,N_18869);
nand U21375 (N_21375,N_19172,N_20653);
or U21376 (N_21376,N_19256,N_18351);
and U21377 (N_21377,N_20146,N_20842);
or U21378 (N_21378,N_19837,N_19130);
and U21379 (N_21379,N_20561,N_20800);
nor U21380 (N_21380,N_18349,N_18652);
nand U21381 (N_21381,N_18907,N_20107);
and U21382 (N_21382,N_20574,N_18418);
nor U21383 (N_21383,N_18842,N_20350);
nor U21384 (N_21384,N_20158,N_19316);
or U21385 (N_21385,N_19686,N_18010);
and U21386 (N_21386,N_20437,N_20916);
and U21387 (N_21387,N_20410,N_20154);
xor U21388 (N_21388,N_19288,N_20853);
and U21389 (N_21389,N_18300,N_18440);
and U21390 (N_21390,N_20026,N_18634);
nor U21391 (N_21391,N_20085,N_19384);
nor U21392 (N_21392,N_20306,N_18172);
and U21393 (N_21393,N_19579,N_18044);
nor U21394 (N_21394,N_20619,N_18725);
nand U21395 (N_21395,N_20214,N_18425);
or U21396 (N_21396,N_18433,N_20344);
nor U21397 (N_21397,N_20441,N_19023);
or U21398 (N_21398,N_18135,N_20537);
and U21399 (N_21399,N_18368,N_19649);
xor U21400 (N_21400,N_18996,N_18089);
xor U21401 (N_21401,N_20633,N_20157);
or U21402 (N_21402,N_20779,N_19626);
and U21403 (N_21403,N_20496,N_19428);
xor U21404 (N_21404,N_19388,N_20325);
nor U21405 (N_21405,N_18786,N_19087);
xnor U21406 (N_21406,N_20602,N_18182);
xor U21407 (N_21407,N_20177,N_19886);
nand U21408 (N_21408,N_19382,N_20540);
nor U21409 (N_21409,N_19012,N_19772);
xor U21410 (N_21410,N_19776,N_18485);
nand U21411 (N_21411,N_19276,N_19717);
xor U21412 (N_21412,N_19969,N_20911);
or U21413 (N_21413,N_19524,N_18167);
or U21414 (N_21414,N_19842,N_19459);
xor U21415 (N_21415,N_19525,N_18919);
or U21416 (N_21416,N_20837,N_20379);
nand U21417 (N_21417,N_19222,N_18396);
or U21418 (N_21418,N_18953,N_20312);
xnor U21419 (N_21419,N_20436,N_20393);
nand U21420 (N_21420,N_20541,N_18805);
xnor U21421 (N_21421,N_19135,N_19959);
xor U21422 (N_21422,N_18494,N_18765);
or U21423 (N_21423,N_19136,N_20888);
and U21424 (N_21424,N_18395,N_20236);
nand U21425 (N_21425,N_18174,N_19994);
or U21426 (N_21426,N_20149,N_19041);
xor U21427 (N_21427,N_19928,N_19284);
and U21428 (N_21428,N_20685,N_20334);
nand U21429 (N_21429,N_20994,N_20519);
nor U21430 (N_21430,N_19752,N_20881);
or U21431 (N_21431,N_19026,N_18018);
nor U21432 (N_21432,N_19482,N_20382);
nor U21433 (N_21433,N_18382,N_20924);
and U21434 (N_21434,N_18385,N_19980);
and U21435 (N_21435,N_18126,N_18450);
or U21436 (N_21436,N_19609,N_20332);
and U21437 (N_21437,N_20768,N_19242);
nor U21438 (N_21438,N_19204,N_18339);
and U21439 (N_21439,N_20931,N_19559);
xnor U21440 (N_21440,N_18432,N_20761);
and U21441 (N_21441,N_18675,N_18232);
nand U21442 (N_21442,N_19174,N_18974);
or U21443 (N_21443,N_19991,N_19119);
and U21444 (N_21444,N_18827,N_20908);
nor U21445 (N_21445,N_20135,N_20046);
xor U21446 (N_21446,N_18881,N_19856);
and U21447 (N_21447,N_20416,N_20790);
or U21448 (N_21448,N_19051,N_20846);
xor U21449 (N_21449,N_20117,N_20282);
nor U21450 (N_21450,N_19755,N_20004);
xor U21451 (N_21451,N_19754,N_19397);
nor U21452 (N_21452,N_19643,N_20071);
or U21453 (N_21453,N_20741,N_18391);
xnor U21454 (N_21454,N_18148,N_19618);
xnor U21455 (N_21455,N_20082,N_18830);
and U21456 (N_21456,N_18655,N_20631);
nor U21457 (N_21457,N_20792,N_20893);
nand U21458 (N_21458,N_20969,N_18664);
or U21459 (N_21459,N_20251,N_19957);
and U21460 (N_21460,N_19820,N_19049);
xnor U21461 (N_21461,N_20169,N_20988);
nand U21462 (N_21462,N_19283,N_19817);
nor U21463 (N_21463,N_18499,N_20446);
nor U21464 (N_21464,N_20957,N_20447);
nor U21465 (N_21465,N_19175,N_19924);
xor U21466 (N_21466,N_19272,N_20386);
xnor U21467 (N_21467,N_20190,N_18092);
nor U21468 (N_21468,N_20785,N_18736);
nor U21469 (N_21469,N_19271,N_20726);
xnor U21470 (N_21470,N_18622,N_20660);
or U21471 (N_21471,N_19474,N_20544);
nand U21472 (N_21472,N_20315,N_18983);
and U21473 (N_21473,N_19133,N_18454);
and U21474 (N_21474,N_20200,N_19322);
nor U21475 (N_21475,N_18253,N_20455);
or U21476 (N_21476,N_18377,N_20297);
or U21477 (N_21477,N_19286,N_18581);
and U21478 (N_21478,N_18882,N_19937);
or U21479 (N_21479,N_19651,N_18627);
xnor U21480 (N_21480,N_18533,N_19640);
xor U21481 (N_21481,N_19947,N_20581);
and U21482 (N_21482,N_20673,N_19075);
nor U21483 (N_21483,N_18110,N_19346);
or U21484 (N_21484,N_18815,N_20706);
nor U21485 (N_21485,N_20453,N_20686);
nor U21486 (N_21486,N_18305,N_20359);
or U21487 (N_21487,N_18462,N_18457);
or U21488 (N_21488,N_20855,N_20491);
and U21489 (N_21489,N_20649,N_19724);
nor U21490 (N_21490,N_18507,N_18552);
xor U21491 (N_21491,N_18005,N_19150);
or U21492 (N_21492,N_19212,N_18636);
nor U21493 (N_21493,N_18001,N_18809);
xnor U21494 (N_21494,N_18892,N_20752);
or U21495 (N_21495,N_18113,N_18302);
or U21496 (N_21496,N_18333,N_19278);
xnor U21497 (N_21497,N_18706,N_19017);
xnor U21498 (N_21498,N_20074,N_19509);
xnor U21499 (N_21499,N_18364,N_19684);
or U21500 (N_21500,N_19217,N_18712);
nand U21501 (N_21501,N_18249,N_20497);
xnor U21502 (N_21502,N_18885,N_18998);
nand U21503 (N_21503,N_20798,N_18156);
nor U21504 (N_21504,N_19617,N_19961);
nand U21505 (N_21505,N_18043,N_20089);
or U21506 (N_21506,N_20818,N_19121);
and U21507 (N_21507,N_19331,N_20387);
or U21508 (N_21508,N_20607,N_19791);
xor U21509 (N_21509,N_20470,N_18977);
or U21510 (N_21510,N_19514,N_20119);
xnor U21511 (N_21511,N_18959,N_20122);
nor U21512 (N_21512,N_19614,N_20072);
xnor U21513 (N_21513,N_19233,N_20194);
nand U21514 (N_21514,N_20514,N_19844);
xnor U21515 (N_21515,N_19813,N_20249);
xnor U21516 (N_21516,N_19033,N_18029);
or U21517 (N_21517,N_20967,N_20047);
nor U21518 (N_21518,N_20593,N_18554);
xor U21519 (N_21519,N_20732,N_20886);
or U21520 (N_21520,N_20062,N_18517);
and U21521 (N_21521,N_18486,N_19613);
nor U21522 (N_21522,N_20833,N_19353);
nand U21523 (N_21523,N_18411,N_18330);
nand U21524 (N_21524,N_18209,N_18831);
and U21525 (N_21525,N_19801,N_20152);
and U21526 (N_21526,N_20182,N_19848);
xor U21527 (N_21527,N_20163,N_18592);
nor U21528 (N_21528,N_18234,N_19446);
and U21529 (N_21529,N_18074,N_19760);
nor U21530 (N_21530,N_18667,N_19290);
nand U21531 (N_21531,N_20483,N_19210);
nor U21532 (N_21532,N_18904,N_18597);
nor U21533 (N_21533,N_20808,N_20720);
nor U21534 (N_21534,N_18076,N_20252);
nand U21535 (N_21535,N_18114,N_20824);
or U21536 (N_21536,N_18242,N_19867);
or U21537 (N_21537,N_19511,N_18818);
xnor U21538 (N_21538,N_20319,N_20353);
nand U21539 (N_21539,N_20356,N_20348);
xor U21540 (N_21540,N_20737,N_20101);
xor U21541 (N_21541,N_19185,N_18164);
xor U21542 (N_21542,N_19262,N_20336);
and U21543 (N_21543,N_20374,N_20655);
xor U21544 (N_21544,N_18587,N_19833);
nand U21545 (N_21545,N_20052,N_18933);
xnor U21546 (N_21546,N_18659,N_20093);
nand U21547 (N_21547,N_18091,N_20895);
or U21548 (N_21548,N_20114,N_18876);
nand U21549 (N_21549,N_19416,N_18394);
and U21550 (N_21550,N_19381,N_20181);
xnor U21551 (N_21551,N_18678,N_18474);
nor U21552 (N_21552,N_19744,N_18591);
nor U21553 (N_21553,N_18341,N_20848);
or U21554 (N_21554,N_18926,N_20210);
or U21555 (N_21555,N_19970,N_20433);
nor U21556 (N_21556,N_19796,N_19880);
nor U21557 (N_21557,N_18726,N_18458);
or U21558 (N_21558,N_19106,N_20636);
nor U21559 (N_21559,N_20698,N_19563);
and U21560 (N_21560,N_18414,N_18764);
and U21561 (N_21561,N_19325,N_19192);
xnor U21562 (N_21562,N_19730,N_19429);
or U21563 (N_21563,N_19569,N_19855);
nand U21564 (N_21564,N_18057,N_20875);
nand U21565 (N_21565,N_20774,N_18147);
nand U21566 (N_21566,N_18472,N_19385);
and U21567 (N_21567,N_18309,N_20498);
nor U21568 (N_21568,N_18436,N_18630);
nand U21569 (N_21569,N_18599,N_18791);
and U21570 (N_21570,N_18589,N_20367);
and U21571 (N_21571,N_19333,N_19419);
xnor U21572 (N_21572,N_18117,N_20844);
xnor U21573 (N_21573,N_20803,N_18673);
nand U21574 (N_21574,N_18460,N_18463);
or U21575 (N_21575,N_18070,N_20137);
or U21576 (N_21576,N_19227,N_18660);
or U21577 (N_21577,N_19623,N_20914);
and U21578 (N_21578,N_18073,N_18859);
xor U21579 (N_21579,N_20873,N_18426);
nand U21580 (N_21580,N_19120,N_19152);
or U21581 (N_21581,N_19929,N_20756);
xnor U21582 (N_21582,N_19902,N_18181);
and U21583 (N_21583,N_18593,N_20399);
or U21584 (N_21584,N_20835,N_19862);
or U21585 (N_21585,N_18366,N_19501);
nand U21586 (N_21586,N_18168,N_18296);
nor U21587 (N_21587,N_18157,N_18793);
or U21588 (N_21588,N_20620,N_20031);
or U21589 (N_21589,N_18004,N_20878);
or U21590 (N_21590,N_19393,N_18837);
nand U21591 (N_21591,N_20504,N_18151);
xnor U21592 (N_21592,N_20419,N_18863);
and U21593 (N_21593,N_19151,N_20572);
xnor U21594 (N_21594,N_19125,N_18497);
and U21595 (N_21595,N_19345,N_18400);
or U21596 (N_21596,N_20646,N_19042);
and U21597 (N_21597,N_20361,N_18995);
and U21598 (N_21598,N_18550,N_19571);
or U21599 (N_21599,N_19200,N_18421);
and U21600 (N_21600,N_20413,N_19161);
nand U21601 (N_21601,N_20339,N_18845);
nand U21602 (N_21602,N_19000,N_20450);
and U21603 (N_21603,N_20095,N_18705);
nor U21604 (N_21604,N_20381,N_18694);
or U21605 (N_21605,N_20900,N_19865);
nand U21606 (N_21606,N_20634,N_19529);
xnor U21607 (N_21607,N_20845,N_18772);
and U21608 (N_21608,N_19178,N_18648);
or U21609 (N_21609,N_20001,N_19979);
or U21610 (N_21610,N_20300,N_20635);
or U21611 (N_21611,N_18097,N_18437);
nand U21612 (N_21612,N_20743,N_18957);
nand U21613 (N_21613,N_20565,N_19716);
xnor U21614 (N_21614,N_20856,N_20758);
nand U21615 (N_21615,N_20925,N_20060);
or U21616 (N_21616,N_20375,N_20341);
nor U21617 (N_21617,N_20639,N_19180);
nand U21618 (N_21618,N_20316,N_18572);
nor U21619 (N_21619,N_19779,N_20814);
nor U21620 (N_21620,N_19072,N_18617);
or U21621 (N_21621,N_18331,N_20929);
and U21622 (N_21622,N_20106,N_20357);
xor U21623 (N_21623,N_18453,N_19707);
nor U21624 (N_21624,N_20153,N_19829);
nor U21625 (N_21625,N_18217,N_19564);
xnor U21626 (N_21626,N_20041,N_19504);
xnor U21627 (N_21627,N_19987,N_19895);
nor U21628 (N_21628,N_19903,N_18204);
or U21629 (N_21629,N_20495,N_18115);
and U21630 (N_21630,N_19295,N_19507);
or U21631 (N_21631,N_18222,N_19312);
or U21632 (N_21632,N_20424,N_18487);
nand U21633 (N_21633,N_18861,N_20208);
and U21634 (N_21634,N_18347,N_20642);
or U21635 (N_21635,N_18567,N_18569);
nand U21636 (N_21636,N_19383,N_20883);
nor U21637 (N_21637,N_18121,N_18956);
and U21638 (N_21638,N_19627,N_20417);
xnor U21639 (N_21639,N_20960,N_18077);
nand U21640 (N_21640,N_18638,N_18353);
and U21641 (N_21641,N_18623,N_20420);
or U21642 (N_21642,N_20289,N_19214);
and U21643 (N_21643,N_18972,N_19208);
nand U21644 (N_21644,N_19403,N_20293);
nand U21645 (N_21645,N_19535,N_19940);
and U21646 (N_21646,N_18807,N_19456);
and U21647 (N_21647,N_18619,N_18698);
nand U21648 (N_21648,N_18083,N_20854);
nor U21649 (N_21649,N_19897,N_19327);
or U21650 (N_21650,N_19995,N_18819);
or U21651 (N_21651,N_18401,N_18833);
nor U21652 (N_21652,N_19234,N_20505);
nor U21653 (N_21653,N_20445,N_19432);
and U21654 (N_21654,N_18255,N_20484);
and U21655 (N_21655,N_18641,N_20178);
and U21656 (N_21656,N_18668,N_20397);
and U21657 (N_21657,N_19756,N_18938);
nand U21658 (N_21658,N_18522,N_20729);
and U21659 (N_21659,N_20281,N_20024);
nor U21660 (N_21660,N_18410,N_19258);
nand U21661 (N_21661,N_19142,N_18025);
xor U21662 (N_21662,N_20385,N_20715);
nand U21663 (N_21663,N_19442,N_18160);
and U21664 (N_21664,N_20722,N_20966);
nand U21665 (N_21665,N_18372,N_19859);
or U21666 (N_21666,N_20991,N_19795);
and U21667 (N_21667,N_19011,N_19144);
nand U21668 (N_21668,N_18639,N_18542);
nor U21669 (N_21669,N_18378,N_18420);
and U21670 (N_21670,N_18696,N_20764);
nor U21671 (N_21671,N_20245,N_20780);
nand U21672 (N_21672,N_18916,N_20597);
nand U21673 (N_21673,N_18653,N_19531);
xor U21674 (N_21674,N_20184,N_18084);
nand U21675 (N_21675,N_20207,N_20535);
and U21676 (N_21676,N_18140,N_18049);
or U21677 (N_21677,N_20109,N_19122);
nor U21678 (N_21678,N_18590,N_20028);
xnor U21679 (N_21679,N_19207,N_20943);
or U21680 (N_21680,N_20765,N_18802);
or U21681 (N_21681,N_18506,N_19159);
or U21682 (N_21682,N_18212,N_19539);
xor U21683 (N_21683,N_18218,N_20971);
xor U21684 (N_21684,N_19469,N_19430);
or U21685 (N_21685,N_18402,N_18961);
or U21686 (N_21686,N_19128,N_20723);
and U21687 (N_21687,N_20254,N_19282);
xor U21688 (N_21688,N_18423,N_18379);
and U21689 (N_21689,N_20175,N_18877);
and U21690 (N_21690,N_18680,N_20168);
or U21691 (N_21691,N_18689,N_20920);
xnor U21692 (N_21692,N_20849,N_20678);
and U21693 (N_21693,N_20187,N_19373);
nor U21694 (N_21694,N_19176,N_19357);
xor U21695 (N_21695,N_20013,N_19030);
or U21696 (N_21696,N_19675,N_20257);
or U21697 (N_21697,N_19485,N_18228);
nor U21698 (N_21698,N_18976,N_19367);
and U21699 (N_21699,N_19237,N_20219);
nand U21700 (N_21700,N_18958,N_20338);
xnor U21701 (N_21701,N_18523,N_19320);
xor U21702 (N_21702,N_19674,N_18801);
xor U21703 (N_21703,N_18984,N_20402);
nor U21704 (N_21704,N_19311,N_18473);
or U21705 (N_21705,N_19490,N_19248);
nand U21706 (N_21706,N_18332,N_19584);
nand U21707 (N_21707,N_18388,N_20936);
or U21708 (N_21708,N_19919,N_18695);
nor U21709 (N_21709,N_19913,N_18898);
nand U21710 (N_21710,N_19816,N_19407);
or U21711 (N_21711,N_20539,N_20092);
nor U21712 (N_21712,N_18047,N_20529);
and U21713 (N_21713,N_19365,N_18874);
nor U21714 (N_21714,N_19455,N_18444);
or U21715 (N_21715,N_19934,N_18883);
nand U21716 (N_21716,N_19078,N_18728);
and U21717 (N_21717,N_18224,N_18913);
or U21718 (N_21718,N_19809,N_20391);
nand U21719 (N_21719,N_20369,N_18019);
nor U21720 (N_21720,N_18795,N_20188);
or U21721 (N_21721,N_18853,N_18176);
nor U21722 (N_21722,N_20998,N_20204);
nor U21723 (N_21723,N_19094,N_19832);
or U21724 (N_21724,N_19694,N_20220);
nor U21725 (N_21725,N_18128,N_18745);
or U21726 (N_21726,N_18771,N_18387);
or U21727 (N_21727,N_18817,N_19548);
nor U21728 (N_21728,N_20716,N_19834);
nor U21729 (N_21729,N_20368,N_19468);
nand U21730 (N_21730,N_18940,N_18015);
nor U21731 (N_21731,N_18229,N_19412);
or U21732 (N_21732,N_20731,N_19839);
nor U21733 (N_21733,N_18191,N_20384);
nor U21734 (N_21734,N_20976,N_20552);
and U21735 (N_21735,N_20295,N_20819);
and U21736 (N_21736,N_19100,N_19055);
and U21737 (N_21737,N_19907,N_19399);
nor U21738 (N_21738,N_20827,N_20066);
nand U21739 (N_21739,N_19047,N_19341);
or U21740 (N_21740,N_19404,N_20927);
or U21741 (N_21741,N_18509,N_20889);
nand U21742 (N_21742,N_18312,N_18480);
and U21743 (N_21743,N_20603,N_18202);
nor U21744 (N_21744,N_19988,N_19189);
or U21745 (N_21745,N_18873,N_20173);
nand U21746 (N_21746,N_19066,N_19888);
and U21747 (N_21747,N_19725,N_19495);
nor U21748 (N_21748,N_18911,N_18244);
or U21749 (N_21749,N_20482,N_19005);
nand U21750 (N_21750,N_19035,N_20486);
or U21751 (N_21751,N_18544,N_19672);
or U21752 (N_21752,N_18035,N_18951);
xnor U21753 (N_21753,N_18665,N_20662);
and U21754 (N_21754,N_18319,N_18455);
nand U21755 (N_21755,N_18360,N_18783);
xnor U21756 (N_21756,N_20805,N_18865);
nand U21757 (N_21757,N_18075,N_19641);
or U21758 (N_21758,N_18456,N_19080);
nand U21759 (N_21759,N_20377,N_19091);
nor U21760 (N_21760,N_18008,N_20759);
xnor U21761 (N_21761,N_19935,N_19370);
and U21762 (N_21762,N_18482,N_19973);
and U21763 (N_21763,N_20465,N_18915);
nor U21764 (N_21764,N_20675,N_19596);
and U21765 (N_21765,N_19226,N_18744);
and U21766 (N_21766,N_20754,N_18163);
and U21767 (N_21767,N_19203,N_18527);
nor U21768 (N_21768,N_18718,N_18806);
nand U21769 (N_21769,N_18565,N_19003);
nor U21770 (N_21770,N_20394,N_20852);
and U21771 (N_21771,N_19634,N_18026);
xor U21772 (N_21772,N_18153,N_18131);
or U21773 (N_21773,N_18539,N_18146);
nor U21774 (N_21774,N_18607,N_20421);
and U21775 (N_21775,N_18247,N_20456);
nand U21776 (N_21776,N_20423,N_18999);
and U21777 (N_21777,N_20964,N_18054);
nor U21778 (N_21778,N_18674,N_18321);
nor U21779 (N_21779,N_20240,N_19183);
or U21780 (N_21780,N_19323,N_20974);
nand U21781 (N_21781,N_19721,N_20021);
xor U21782 (N_21782,N_19489,N_19582);
nand U21783 (N_21783,N_20270,N_19289);
xor U21784 (N_21784,N_20110,N_20970);
or U21785 (N_21785,N_20134,N_18441);
and U21786 (N_21786,N_18848,N_18993);
and U21787 (N_21787,N_20400,N_18285);
nor U21788 (N_21788,N_19179,N_19315);
or U21789 (N_21789,N_20428,N_18906);
xnor U21790 (N_21790,N_20872,N_18166);
nor U21791 (N_21791,N_18616,N_18356);
xor U21792 (N_21792,N_19239,N_20081);
nor U21793 (N_21793,N_19492,N_18415);
nor U21794 (N_21794,N_19251,N_18626);
nand U21795 (N_21795,N_19861,N_19712);
xnor U21796 (N_21796,N_18079,N_19847);
nand U21797 (N_21797,N_19028,N_18362);
nand U21798 (N_21798,N_19157,N_18936);
and U21799 (N_21799,N_18596,N_19221);
nand U21800 (N_21800,N_20172,N_18119);
nand U21801 (N_21801,N_19206,N_18858);
nor U21802 (N_21802,N_19497,N_18986);
or U21803 (N_21803,N_20224,N_18536);
xnor U21804 (N_21804,N_19930,N_20422);
nand U21805 (N_21805,N_20216,N_20223);
nor U21806 (N_21806,N_18841,N_20921);
xnor U21807 (N_21807,N_19194,N_20727);
nor U21808 (N_21808,N_18315,N_19332);
nor U21809 (N_21809,N_20140,N_19330);
and U21810 (N_21810,N_18488,N_19590);
nor U21811 (N_21811,N_18838,N_19777);
nor U21812 (N_21812,N_18943,N_18282);
nand U21813 (N_21813,N_18732,N_18612);
nand U21814 (N_21814,N_20038,N_19314);
nor U21815 (N_21815,N_19039,N_20983);
and U21816 (N_21816,N_18000,N_18286);
xor U21817 (N_21817,N_18851,N_18835);
and U21818 (N_21818,N_18510,N_19797);
nand U21819 (N_21819,N_19573,N_19046);
nor U21820 (N_21820,N_20599,N_20987);
xor U21821 (N_21821,N_20562,N_20796);
nor U21822 (N_21822,N_18629,N_19024);
xnor U21823 (N_21823,N_19196,N_20042);
xor U21824 (N_21824,N_20950,N_20692);
nand U21825 (N_21825,N_18594,N_20395);
nand U21826 (N_21826,N_20324,N_20176);
nand U21827 (N_21827,N_19769,N_19014);
or U21828 (N_21828,N_18500,N_20232);
and U21829 (N_21829,N_18826,N_20753);
and U21830 (N_21830,N_19513,N_18236);
nor U21831 (N_21831,N_20530,N_19784);
xor U21832 (N_21832,N_18154,N_20583);
nand U21833 (N_21833,N_20454,N_18729);
nor U21834 (N_21834,N_18071,N_18504);
and U21835 (N_21835,N_20564,N_20449);
or U21836 (N_21836,N_20945,N_20309);
nor U21837 (N_21837,N_18225,N_20902);
or U21838 (N_21838,N_20076,N_18183);
xor U21839 (N_21839,N_19309,N_19925);
and U21840 (N_21840,N_19846,N_18575);
and U21841 (N_21841,N_19823,N_18635);
and U21842 (N_21842,N_19985,N_19359);
nor U21843 (N_21843,N_19757,N_19021);
or U21844 (N_21844,N_20029,N_18481);
or U21845 (N_21845,N_19182,N_18048);
and U21846 (N_21846,N_19875,N_18796);
or U21847 (N_21847,N_20018,N_19787);
nor U21848 (N_21848,N_20360,N_18177);
and U21849 (N_21849,N_19163,N_18095);
xor U21850 (N_21850,N_18052,N_18294);
or U21851 (N_21851,N_20601,N_19445);
and U21852 (N_21852,N_20196,N_20104);
or U21853 (N_21853,N_18103,N_20264);
xor U21854 (N_21854,N_19687,N_20378);
nor U21855 (N_21855,N_19932,N_19606);
xor U21856 (N_21856,N_19864,N_20782);
or U21857 (N_21857,N_18750,N_18145);
and U21858 (N_21858,N_19551,N_19997);
and U21859 (N_21859,N_18491,N_20509);
nor U21860 (N_21860,N_19879,N_19038);
xor U21861 (N_21861,N_20939,N_18413);
nor U21862 (N_21862,N_19350,N_20520);
or U21863 (N_21863,N_20904,N_18030);
or U21864 (N_21864,N_18645,N_18980);
or U21865 (N_21865,N_19636,N_19209);
nand U21866 (N_21866,N_20313,N_18557);
and U21867 (N_21867,N_19195,N_19741);
nor U21868 (N_21868,N_18405,N_20265);
nor U21869 (N_21869,N_20308,N_19088);
nor U21870 (N_21870,N_20039,N_20113);
or U21871 (N_21871,N_18316,N_20458);
or U21872 (N_21872,N_20314,N_20231);
and U21873 (N_21873,N_19803,N_18927);
nand U21874 (N_21874,N_19111,N_20918);
nor U21875 (N_21875,N_18301,N_19240);
xnor U21876 (N_21876,N_18133,N_20789);
or U21877 (N_21877,N_20629,N_20979);
xnor U21878 (N_21878,N_19498,N_18197);
nand U21879 (N_21879,N_19434,N_19644);
nor U21880 (N_21880,N_18985,N_19168);
nor U21881 (N_21881,N_19936,N_19926);
nand U21882 (N_21882,N_18782,N_19146);
nor U21883 (N_21883,N_19824,N_19090);
nand U21884 (N_21884,N_20328,N_20003);
or U21885 (N_21885,N_19425,N_20000);
nor U21886 (N_21886,N_20624,N_20680);
nor U21887 (N_21887,N_20784,N_18545);
xor U21888 (N_21888,N_18620,N_19369);
and U21889 (N_21889,N_18346,N_20429);
nand U21890 (N_21890,N_18676,N_19948);
xor U21891 (N_21891,N_19917,N_20349);
nor U21892 (N_21892,N_19368,N_20317);
or U21893 (N_21893,N_19822,N_19998);
nor U21894 (N_21894,N_18417,N_18610);
or U21895 (N_21895,N_20567,N_20989);
nor U21896 (N_21896,N_18122,N_18656);
nor U21897 (N_21897,N_20371,N_20906);
xor U21898 (N_21898,N_19304,N_19778);
xor U21899 (N_21899,N_20700,N_19774);
nor U21900 (N_21900,N_20398,N_19678);
or U21901 (N_21901,N_18262,N_20010);
nor U21902 (N_21902,N_19806,N_19920);
xnor U21903 (N_21903,N_20099,N_19287);
and U21904 (N_21904,N_19054,N_20073);
or U21905 (N_21905,N_18310,N_18799);
and U21906 (N_21906,N_20518,N_20380);
nor U21907 (N_21907,N_20913,N_18558);
or U21908 (N_21908,N_18857,N_20701);
or U21909 (N_21909,N_19808,N_19073);
nand U21910 (N_21910,N_19292,N_18479);
xor U21911 (N_21911,N_20477,N_18313);
and U21912 (N_21912,N_19993,N_20621);
nor U21913 (N_21913,N_20907,N_18250);
nor U21914 (N_21914,N_18020,N_18158);
or U21915 (N_21915,N_18577,N_19043);
nor U21916 (N_21916,N_18502,N_19735);
nand U21917 (N_21917,N_18856,N_18829);
xnor U21918 (N_21918,N_20507,N_19697);
and U21919 (N_21919,N_20670,N_18810);
xnor U21920 (N_21920,N_19466,N_18740);
nand U21921 (N_21921,N_19526,N_20442);
nor U21922 (N_21922,N_18171,N_20746);
and U21923 (N_21923,N_20508,N_20389);
and U21924 (N_21924,N_19347,N_20719);
and U21925 (N_21925,N_19433,N_19577);
or U21926 (N_21926,N_19911,N_19894);
nor U21927 (N_21927,N_20870,N_19540);
xor U21928 (N_21928,N_20697,N_20221);
or U21929 (N_21929,N_20627,N_18704);
nand U21930 (N_21930,N_18459,N_18967);
xnor U21931 (N_21931,N_19069,N_20063);
xor U21932 (N_21932,N_19440,N_18700);
xnor U21933 (N_21933,N_19134,N_20064);
nand U21934 (N_21934,N_19647,N_18289);
nor U21935 (N_21935,N_19873,N_20199);
or U21936 (N_21936,N_19224,N_19689);
nor U21937 (N_21937,N_20461,N_18518);
and U21938 (N_21938,N_18679,N_19691);
or U21939 (N_21939,N_20116,N_20816);
xnor U21940 (N_21940,N_18948,N_19408);
and U21941 (N_21941,N_19944,N_20690);
nor U21942 (N_21942,N_19561,N_18928);
and U21943 (N_21943,N_18287,N_18685);
nor U21944 (N_21944,N_19307,N_19996);
and U21945 (N_21945,N_20301,N_19318);
xor U21946 (N_21946,N_18130,N_19914);
or U21947 (N_21947,N_18263,N_19268);
nor U21948 (N_21948,N_20693,N_18798);
or U21949 (N_21949,N_19245,N_20815);
nand U21950 (N_21950,N_20630,N_19952);
nor U21951 (N_21951,N_19019,N_20213);
nand U21952 (N_21952,N_18094,N_20305);
nand U21953 (N_21953,N_20115,N_19783);
or U21954 (N_21954,N_19400,N_18585);
xnor U21955 (N_21955,N_19642,N_18329);
nand U21956 (N_21956,N_20942,N_20559);
nand U21957 (N_21957,N_18283,N_20346);
xnor U21958 (N_21958,N_20666,N_19693);
or U21959 (N_21959,N_18787,N_20772);
nor U21960 (N_21960,N_20516,N_19603);
and U21961 (N_21961,N_18931,N_18098);
nor U21962 (N_21962,N_18081,N_20563);
nor U21963 (N_21963,N_20751,N_19319);
nand U21964 (N_21964,N_18780,N_19277);
or U21965 (N_21965,N_20748,N_20193);
nand U21966 (N_21966,N_20197,N_20239);
nor U21967 (N_21967,N_19375,N_20262);
nand U21968 (N_21968,N_20699,N_19633);
and U21969 (N_21969,N_19978,N_20480);
nand U21970 (N_21970,N_19020,N_18340);
nor U21971 (N_21971,N_20123,N_18803);
and U21972 (N_21972,N_19550,N_19236);
xnor U21973 (N_21973,N_20139,N_20267);
xor U21974 (N_21974,N_18511,N_20460);
nand U21975 (N_21975,N_18032,N_18065);
xor U21976 (N_21976,N_20131,N_19545);
or U21977 (N_21977,N_19715,N_18814);
xnor U21978 (N_21978,N_19951,N_18272);
and U21979 (N_21979,N_19943,N_20370);
nor U21980 (N_21980,N_19635,N_18954);
xnor U21981 (N_21981,N_20956,N_18039);
nor U21982 (N_21982,N_18118,N_18979);
and U21983 (N_21983,N_19632,N_18129);
nor U21984 (N_21984,N_19575,N_18947);
or U21985 (N_21985,N_18096,N_18794);
xnor U21986 (N_21986,N_18538,N_20869);
nor U21987 (N_21987,N_19748,N_18945);
xor U21988 (N_21988,N_20573,N_18124);
and U21989 (N_21989,N_18520,N_18547);
nor U21990 (N_21990,N_20648,N_20141);
nand U21991 (N_21991,N_20425,N_20543);
nor U21992 (N_21992,N_18342,N_18254);
or U21993 (N_21993,N_20859,N_18187);
and U21994 (N_21994,N_20404,N_20217);
nor U21995 (N_21995,N_20838,N_20817);
nor U21996 (N_21996,N_18006,N_18535);
or U21997 (N_21997,N_18050,N_19927);
nand U21998 (N_21998,N_19922,N_19148);
or U21999 (N_21999,N_19706,N_18483);
nor U22000 (N_22000,N_18934,N_18139);
nor U22001 (N_22001,N_19431,N_20225);
or U22002 (N_22002,N_19306,N_18336);
or U22003 (N_22003,N_19334,N_19898);
xor U22004 (N_22004,N_19056,N_19158);
or U22005 (N_22005,N_19452,N_19587);
xnor U22006 (N_22006,N_19699,N_18467);
and U22007 (N_22007,N_18584,N_19279);
nor U22008 (N_22008,N_18064,N_20887);
xnor U22009 (N_22009,N_20840,N_19597);
xnor U22010 (N_22010,N_18820,N_19908);
or U22011 (N_22011,N_18969,N_19639);
xnor U22012 (N_22012,N_19086,N_20980);
nand U22013 (N_22013,N_18326,N_20206);
or U22014 (N_22014,N_20414,N_18170);
or U22015 (N_22015,N_19981,N_19269);
xor U22016 (N_22016,N_20363,N_19574);
nand U22017 (N_22017,N_18503,N_19390);
or U22018 (N_22018,N_20329,N_18946);
nor U22019 (N_22019,N_20303,N_20757);
and U22020 (N_22020,N_19942,N_19547);
nand U22021 (N_22021,N_19965,N_20211);
and U22022 (N_22022,N_19464,N_18149);
nand U22023 (N_22023,N_20999,N_20689);
or U22024 (N_22024,N_18162,N_20851);
and U22025 (N_22025,N_19001,N_18307);
nand U22026 (N_22026,N_19064,N_18605);
nand U22027 (N_22027,N_18614,N_20762);
xor U22028 (N_22028,N_19505,N_18099);
or U22029 (N_22029,N_19171,N_19281);
nand U22030 (N_22030,N_19013,N_18925);
xnor U22031 (N_22031,N_19360,N_20531);
or U22032 (N_22032,N_19671,N_18942);
nand U22033 (N_22033,N_18238,N_18058);
nor U22034 (N_22034,N_18404,N_18563);
nand U22035 (N_22035,N_19167,N_19131);
xnor U22036 (N_22036,N_19481,N_18430);
xnor U22037 (N_22037,N_18800,N_20298);
xnor U22038 (N_22038,N_19389,N_20749);
and U22039 (N_22039,N_18251,N_20794);
or U22040 (N_22040,N_18496,N_20343);
xnor U22041 (N_22041,N_19542,N_20777);
nand U22042 (N_22042,N_20897,N_20269);
xor U22043 (N_22043,N_20166,N_18864);
nand U22044 (N_22044,N_18534,N_20951);
nand U22045 (N_22045,N_18769,N_19451);
nor U22046 (N_22046,N_18017,N_19537);
nor U22047 (N_22047,N_19285,N_20272);
or U22048 (N_22048,N_19165,N_18165);
nor U22049 (N_22049,N_18348,N_19129);
nor U22050 (N_22050,N_19467,N_19812);
or U22051 (N_22051,N_20506,N_19298);
nor U22052 (N_22052,N_18359,N_18918);
nand U22053 (N_22053,N_19896,N_18893);
xnor U22054 (N_22054,N_20144,N_18524);
and U22055 (N_22055,N_19799,N_18381);
or U22056 (N_22056,N_19941,N_19308);
or U22057 (N_22057,N_20788,N_20192);
or U22058 (N_22058,N_20928,N_20735);
nand U22059 (N_22059,N_19444,N_19702);
nand U22060 (N_22060,N_20825,N_18169);
nor U22061 (N_22061,N_19764,N_19335);
xor U22062 (N_22062,N_18621,N_20874);
xor U22063 (N_22063,N_20822,N_20070);
or U22064 (N_22064,N_18009,N_18773);
or U22065 (N_22065,N_19899,N_19299);
or U22066 (N_22066,N_20781,N_20230);
nor U22067 (N_22067,N_20053,N_19254);
nor U22068 (N_22068,N_18241,N_19275);
nand U22069 (N_22069,N_19362,N_20320);
nor U22070 (N_22070,N_19939,N_18448);
and U22071 (N_22071,N_19669,N_19831);
nor U22072 (N_22072,N_19058,N_18746);
nor U22073 (N_22073,N_19814,N_19807);
and U22074 (N_22074,N_18260,N_20440);
nor U22075 (N_22075,N_20045,N_20009);
nor U22076 (N_22076,N_20025,N_18571);
xnor U22077 (N_22077,N_20340,N_18516);
xnor U22078 (N_22078,N_20011,N_20711);
nor U22079 (N_22079,N_19104,N_20523);
nor U22080 (N_22080,N_20078,N_20525);
xor U22081 (N_22081,N_19116,N_18753);
xnor U22082 (N_22082,N_19488,N_19414);
or U22083 (N_22083,N_20640,N_19491);
xor U22084 (N_22084,N_19714,N_20365);
xor U22085 (N_22085,N_19186,N_18568);
or U22086 (N_22086,N_20867,N_20112);
nand U22087 (N_22087,N_19181,N_19435);
xor U22088 (N_22088,N_19085,N_20248);
nand U22089 (N_22089,N_20687,N_20713);
nor U22090 (N_22090,N_18196,N_18671);
nand U22091 (N_22091,N_20566,N_20485);
and U22092 (N_22092,N_18813,N_18647);
nand U22093 (N_22093,N_19396,N_18337);
or U22094 (N_22094,N_20963,N_19267);
nor U22095 (N_22095,N_20284,N_20501);
xor U22096 (N_22096,N_18137,N_18452);
and U22097 (N_22097,N_18284,N_19956);
xnor U22098 (N_22098,N_19933,N_18997);
and U22099 (N_22099,N_18586,N_19484);
or U22100 (N_22100,N_18363,N_20968);
xor U22101 (N_22101,N_19663,N_20326);
or U22102 (N_22102,N_19067,N_20847);
nor U22103 (N_22103,N_18840,N_18235);
or U22104 (N_22104,N_20578,N_18766);
or U22105 (N_22105,N_20118,N_20086);
or U22106 (N_22106,N_18369,N_19532);
xor U22107 (N_22107,N_20984,N_18779);
or U22108 (N_22108,N_20598,N_19191);
xnor U22109 (N_22109,N_18789,N_20703);
or U22110 (N_22110,N_20268,N_18747);
nor U22111 (N_22111,N_19112,N_18240);
or U22112 (N_22112,N_19349,N_19552);
or U22113 (N_22113,N_20291,N_19071);
xnor U22114 (N_22114,N_20280,N_18175);
nor U22115 (N_22115,N_19815,N_18016);
and U22116 (N_22116,N_20773,N_18161);
and U22117 (N_22117,N_19560,N_20478);
xnor U22118 (N_22118,N_19698,N_18259);
nand U22119 (N_22119,N_19696,N_20669);
nor U22120 (N_22120,N_20489,N_19117);
and U22121 (N_22121,N_20993,N_19187);
xor U22122 (N_22122,N_19534,N_18277);
nand U22123 (N_22123,N_18601,N_18033);
and U22124 (N_22124,N_19915,N_18409);
and U22125 (N_22125,N_19745,N_18939);
nor U22126 (N_22126,N_20553,N_19127);
and U22127 (N_22127,N_19775,N_19974);
nand U22128 (N_22128,N_20901,N_18012);
nor U22129 (N_22129,N_18443,N_18657);
or U22130 (N_22130,N_20125,N_18658);
or U22131 (N_22131,N_18743,N_20879);
xnor U22132 (N_22132,N_19763,N_19650);
nor U22133 (N_22133,N_18231,N_19967);
or U22134 (N_22134,N_18334,N_19605);
and U22135 (N_22135,N_20643,N_19264);
or U22136 (N_22136,N_19954,N_20884);
or U22137 (N_22137,N_18192,N_20898);
xnor U22138 (N_22138,N_20167,N_20547);
and U22139 (N_22139,N_18270,N_18755);
nor U22140 (N_22140,N_20986,N_19219);
and U22141 (N_22141,N_20843,N_19061);
or U22142 (N_22142,N_19162,N_20503);
nand U22143 (N_22143,N_18355,N_19426);
nor U22144 (N_22144,N_18735,N_18045);
and U22145 (N_22145,N_20899,N_18515);
nand U22146 (N_22146,N_19881,N_18398);
nor U22147 (N_22147,N_19736,N_20589);
or U22148 (N_22148,N_19392,N_18784);
nand U22149 (N_22149,N_18357,N_18380);
nand U22150 (N_22150,N_19225,N_18989);
and U22151 (N_22151,N_20555,N_18528);
nand U22152 (N_22152,N_20617,N_18068);
nand U22153 (N_22153,N_20435,N_19053);
and U22154 (N_22154,N_19216,N_19102);
or U22155 (N_22155,N_20279,N_19461);
nand U22156 (N_22156,N_18219,N_18186);
nor U22157 (N_22157,N_20799,N_18682);
nor U22158 (N_22158,N_20258,N_20015);
nand U22159 (N_22159,N_19670,N_18962);
nor U22160 (N_22160,N_20659,N_18056);
or U22161 (N_22161,N_18066,N_19863);
xnor U22162 (N_22162,N_20682,N_19904);
xnor U22163 (N_22163,N_18895,N_18770);
nand U22164 (N_22164,N_19652,N_20783);
nand U22165 (N_22165,N_19891,N_19916);
xnor U22166 (N_22166,N_19562,N_18478);
and U22167 (N_22167,N_19065,N_20892);
nor U22168 (N_22168,N_20027,N_18252);
and U22169 (N_22169,N_19500,N_18038);
and U22170 (N_22170,N_18532,N_18702);
or U22171 (N_22171,N_20323,N_20260);
or U22172 (N_22172,N_18902,N_18290);
or U22173 (N_22173,N_20829,N_19654);
and U22174 (N_22174,N_18579,N_20185);
nor U22175 (N_22175,N_18466,N_18127);
xnor U22176 (N_22176,N_19302,N_18264);
or U22177 (N_22177,N_20657,N_19734);
nand U22178 (N_22178,N_20292,N_20717);
nand U22179 (N_22179,N_19037,N_18489);
xor U22180 (N_22180,N_20571,N_20452);
xnor U22181 (N_22181,N_19198,N_20473);
nand U22182 (N_22182,N_18464,N_19646);
or U22183 (N_22183,N_20409,N_18193);
and U22184 (N_22184,N_19770,N_19615);
nand U22185 (N_22185,N_20459,N_20253);
and U22186 (N_22186,N_20500,N_18392);
and U22187 (N_22187,N_20736,N_18847);
and U22188 (N_22188,N_18246,N_19124);
or U22189 (N_22189,N_18875,N_19723);
nand U22190 (N_22190,N_20612,N_18714);
xor U22191 (N_22191,N_20427,N_20834);
nand U22192 (N_22192,N_20684,N_20546);
nor U22193 (N_22193,N_20623,N_18541);
nand U22194 (N_22194,N_18650,N_18897);
nor U22195 (N_22195,N_19170,N_18512);
nand U22196 (N_22196,N_18930,N_18200);
or U22197 (N_22197,N_20975,N_18298);
and U22198 (N_22198,N_19923,N_18960);
nand U22199 (N_22199,N_18484,N_19415);
xor U22200 (N_22200,N_20430,N_18543);
nor U22201 (N_22201,N_19438,N_19273);
xnor U22202 (N_22202,N_18295,N_19781);
or U22203 (N_22203,N_19232,N_20059);
nor U22204 (N_22204,N_19767,N_19211);
nand U22205 (N_22205,N_19872,N_19008);
xnor U22206 (N_22206,N_20750,N_18141);
nand U22207 (N_22207,N_19611,N_19659);
nor U22208 (N_22208,N_19870,N_18792);
xnor U22209 (N_22209,N_18185,N_19522);
or U22210 (N_22210,N_19344,N_18762);
nor U22211 (N_22211,N_18207,N_19595);
or U22212 (N_22212,N_20973,N_19938);
and U22213 (N_22213,N_18429,N_20613);
or U22214 (N_22214,N_20738,N_20712);
nand U22215 (N_22215,N_18703,N_19612);
nand U22216 (N_22216,N_19259,N_20006);
xor U22217 (N_22217,N_19853,N_19062);
and U22218 (N_22218,N_19108,N_19637);
nor U22219 (N_22219,N_20351,N_20212);
nor U22220 (N_22220,N_20937,N_20679);
or U22221 (N_22221,N_19402,N_18108);
nand U22222 (N_22222,N_20661,N_18720);
nand U22223 (N_22223,N_18230,N_18223);
nor U22224 (N_22224,N_20591,N_19523);
xnor U22225 (N_22225,N_18105,N_20592);
or U22226 (N_22226,N_18900,N_19114);
xor U22227 (N_22227,N_19113,N_20663);
nor U22228 (N_22228,N_18269,N_18693);
nor U22229 (N_22229,N_18903,N_20801);
nand U22230 (N_22230,N_18422,N_20307);
and U22231 (N_22231,N_20017,N_18560);
xor U22232 (N_22232,N_18751,N_18886);
xor U22233 (N_22233,N_19354,N_19479);
and U22234 (N_22234,N_20804,N_18669);
xnor U22235 (N_22235,N_19352,N_20860);
and U22236 (N_22236,N_20616,N_18120);
xor U22237 (N_22237,N_18757,N_18672);
nor U22238 (N_22238,N_18576,N_20286);
nor U22239 (N_22239,N_20057,N_19713);
or U22240 (N_22240,N_19417,N_20311);
xor U22241 (N_22241,N_18111,N_20560);
or U22242 (N_22242,N_20097,N_19628);
nor U22243 (N_22243,N_19554,N_19378);
xnor U22244 (N_22244,N_20276,N_18812);
nor U22245 (N_22245,N_19544,N_19480);
and U22246 (N_22246,N_20590,N_19593);
nand U22247 (N_22247,N_19246,N_18325);
or U22248 (N_22248,N_18245,N_20432);
xor U22249 (N_22249,N_18884,N_19447);
nor U22250 (N_22250,N_20608,N_19427);
and U22251 (N_22251,N_18924,N_18501);
nor U22252 (N_22252,N_19624,N_18790);
nand U22253 (N_22253,N_19620,N_20203);
nand U22254 (N_22254,N_19029,N_20077);
or U22255 (N_22255,N_18691,N_18085);
nor U22256 (N_22256,N_20392,N_19265);
xor U22257 (N_22257,N_18888,N_20080);
nor U22258 (N_22258,N_20285,N_18677);
nor U22259 (N_22259,N_20577,N_18549);
and U22260 (N_22260,N_18027,N_19963);
and U22261 (N_22261,N_20094,N_20273);
or U22262 (N_22262,N_19079,N_19793);
nand U22263 (N_22263,N_19766,N_20714);
nand U22264 (N_22264,N_18852,N_19300);
and U22265 (N_22265,N_18643,N_20275);
nor U22266 (N_22266,N_20982,N_20467);
and U22267 (N_22267,N_18583,N_18846);
or U22268 (N_22268,N_20709,N_20667);
or U22269 (N_22269,N_19804,N_19118);
nand U22270 (N_22270,N_18257,N_19266);
nor U22271 (N_22271,N_19765,N_19599);
nor U22272 (N_22272,N_20977,N_20917);
and U22273 (N_22273,N_19166,N_20274);
or U22274 (N_22274,N_18505,N_20862);
nand U22275 (N_22275,N_20012,N_20290);
nand U22276 (N_22276,N_19199,N_20647);
and U22277 (N_22277,N_19557,N_18178);
or U22278 (N_22278,N_18072,N_18314);
nand U22279 (N_22279,N_19409,N_19838);
and U22280 (N_22280,N_19018,N_19249);
nand U22281 (N_22281,N_18024,N_18393);
and U22282 (N_22282,N_20905,N_18352);
nor U22283 (N_22283,N_18754,N_19749);
xor U22284 (N_22284,N_20512,N_18734);
or U22285 (N_22285,N_20121,N_20826);
xor U22286 (N_22286,N_18637,N_18978);
nand U22287 (N_22287,N_20949,N_20940);
and U22288 (N_22288,N_20694,N_19296);
or U22289 (N_22289,N_18226,N_19664);
nor U22290 (N_22290,N_20345,N_18082);
xnor U22291 (N_22291,N_19348,N_18508);
or U22292 (N_22292,N_19031,N_19439);
nor U22293 (N_22293,N_19294,N_20728);
or U22294 (N_22294,N_19695,N_18101);
nor U22295 (N_22295,N_18023,N_19443);
xor U22296 (N_22296,N_18275,N_19084);
xnor U22297 (N_22297,N_19594,N_18519);
or U22298 (N_22298,N_19990,N_20201);
xnor U22299 (N_22299,N_19565,N_18447);
and U22300 (N_22300,N_18374,N_20618);
and U22301 (N_22301,N_19983,N_18258);
nand U22302 (N_22302,N_19570,N_18595);
xor U22303 (N_22303,N_19238,N_19462);
nor U22304 (N_22304,N_20127,N_19215);
and U22305 (N_22305,N_19010,N_20841);
xnor U22306 (N_22306,N_19738,N_19830);
nor U22307 (N_22307,N_18661,N_19921);
and U22308 (N_22308,N_18632,N_18317);
nand U22309 (N_22309,N_19036,N_18318);
or U22310 (N_22310,N_20475,N_20250);
xnor U22311 (N_22311,N_20882,N_18384);
nand U22312 (N_22312,N_18763,N_18031);
or U22313 (N_22313,N_18376,N_19137);
nor U22314 (N_22314,N_20288,N_19339);
and U22315 (N_22315,N_20721,N_18327);
nor U22316 (N_22316,N_19077,N_19321);
and U22317 (N_22317,N_19510,N_20469);
nor U22318 (N_22318,N_19740,N_19868);
xnor U22319 (N_22319,N_20333,N_19202);
nand U22320 (N_22320,N_20995,N_18905);
nor U22321 (N_22321,N_18662,N_19553);
nand U22322 (N_22322,N_19109,N_20155);
or U22323 (N_22323,N_20055,N_19601);
and U22324 (N_22324,N_20418,N_20222);
xor U22325 (N_22325,N_18738,N_19912);
or U22326 (N_22326,N_19115,N_20161);
nor U22327 (N_22327,N_20912,N_20227);
xnor U22328 (N_22328,N_19132,N_19821);
nand U22329 (N_22329,N_19878,N_18134);
xor U22330 (N_22330,N_18059,N_18760);
and U22331 (N_22331,N_20903,N_20049);
nand U22332 (N_22332,N_20362,N_20626);
nor U22333 (N_22333,N_18055,N_20807);
nor U22334 (N_22334,N_18060,N_20812);
nor U22335 (N_22335,N_18303,N_20191);
and U22336 (N_22336,N_20271,N_18106);
and U22337 (N_22337,N_19989,N_19892);
nor U22338 (N_22338,N_18816,N_20186);
xor U22339 (N_22339,N_20894,N_19138);
or U22340 (N_22340,N_19052,N_18116);
xor U22341 (N_22341,N_19074,N_18923);
or U22342 (N_22342,N_20164,N_19377);
and U22343 (N_22343,N_19448,N_18776);
or U22344 (N_22344,N_19692,N_20775);
xnor U22345 (N_22345,N_20863,N_20813);
nor U22346 (N_22346,N_19992,N_18646);
or U22347 (N_22347,N_18373,N_20524);
and U22348 (N_22348,N_19953,N_20595);
nor U22349 (N_22349,N_20179,N_18449);
or U22350 (N_22350,N_18692,N_19860);
nor U22351 (N_22351,N_19718,N_20797);
nor U22352 (N_22352,N_18375,N_20431);
nor U22353 (N_22353,N_20725,N_20836);
and U22354 (N_22354,N_19280,N_19476);
nand U22355 (N_22355,N_20955,N_19048);
nor U22356 (N_22356,N_19255,N_20880);
xnor U22357 (N_22357,N_18188,N_18367);
xor U22358 (N_22358,N_20941,N_18878);
nor U22359 (N_22359,N_20002,N_19355);
xnor U22360 (N_22360,N_20575,N_18777);
nor U22361 (N_22361,N_18935,N_19866);
or U22362 (N_22362,N_19081,N_19143);
xnor U22363 (N_22363,N_18742,N_18529);
or U22364 (N_22364,N_18708,N_19884);
or U22365 (N_22365,N_18849,N_19900);
or U22366 (N_22366,N_20256,N_18721);
or U22367 (N_22367,N_19751,N_20611);
or U22368 (N_22368,N_19291,N_20145);
and U22369 (N_22369,N_18717,N_20954);
or U22370 (N_22370,N_19436,N_19140);
or U22371 (N_22371,N_18461,N_20228);
nor U22372 (N_22372,N_18781,N_19123);
nand U22373 (N_22373,N_19798,N_20664);
and U22374 (N_22374,N_20549,N_20411);
nand U22375 (N_22375,N_19709,N_18123);
and U22376 (N_22376,N_20932,N_19572);
xnor U22377 (N_22377,N_18701,N_18150);
or U22378 (N_22378,N_18941,N_18304);
nor U22379 (N_22379,N_19982,N_20556);
nand U22380 (N_22380,N_18324,N_18014);
and U22381 (N_22381,N_20915,N_18273);
nor U22382 (N_22382,N_20035,N_19662);
nor U22383 (N_22383,N_19680,N_20438);
and U22384 (N_22384,N_20528,N_20891);
xor U22385 (N_22385,N_19110,N_18525);
nand U22386 (N_22386,N_20548,N_20376);
nor U22387 (N_22387,N_19986,N_20517);
or U22388 (N_22388,N_20096,N_19022);
or U22389 (N_22389,N_19098,N_19743);
nand U22390 (N_22390,N_20511,N_19722);
xor U22391 (N_22391,N_18526,N_18872);
nand U22392 (N_22392,N_19475,N_20695);
nand U22393 (N_22393,N_20744,N_19089);
and U22394 (N_22394,N_20605,N_20322);
xor U22395 (N_22395,N_19566,N_18292);
nand U22396 (N_22396,N_20235,N_19701);
nand U22397 (N_22397,N_20048,N_18086);
nand U22398 (N_22398,N_18574,N_18233);
nor U22399 (N_22399,N_19975,N_20354);
xnor U22400 (N_22400,N_20098,N_19527);
and U22401 (N_22401,N_19731,N_18051);
and U22402 (N_22402,N_19516,N_19363);
nor U22403 (N_22403,N_20205,N_19608);
nand U22404 (N_22404,N_18644,N_19336);
or U22405 (N_22405,N_18155,N_18445);
xnor U22406 (N_22406,N_18439,N_18267);
xor U22407 (N_22407,N_19093,N_19153);
xor U22408 (N_22408,N_19681,N_19568);
xor U22409 (N_22409,N_20471,N_20625);
nor U22410 (N_22410,N_19854,N_20065);
and U22411 (N_22411,N_20337,N_18173);
xnor U22412 (N_22412,N_20832,N_19810);
or U22413 (N_22413,N_18785,N_20923);
nand U22414 (N_22414,N_19742,N_18600);
and U22415 (N_22415,N_18774,N_20405);
and U22416 (N_22416,N_18199,N_18929);
nand U22417 (N_22417,N_20487,N_18688);
nand U22418 (N_22418,N_20069,N_19502);
or U22419 (N_22419,N_20266,N_20396);
xor U22420 (N_22420,N_20180,N_19421);
or U22421 (N_22421,N_20606,N_19057);
nor U22422 (N_22422,N_18206,N_20443);
or U22423 (N_22423,N_19893,N_19788);
xnor U22424 (N_22424,N_19543,N_19006);
or U22425 (N_22425,N_18215,N_20952);
nor U22426 (N_22426,N_19739,N_20050);
and U22427 (N_22427,N_20760,N_18013);
or U22428 (N_22428,N_19660,N_20802);
and U22429 (N_22429,N_19668,N_19890);
nand U22430 (N_22430,N_19586,N_18390);
nand U22431 (N_22431,N_18687,N_19835);
and U22432 (N_22432,N_18890,N_18912);
or U22433 (N_22433,N_18963,N_18537);
nor U22434 (N_22434,N_19737,N_18768);
nor U22435 (N_22435,N_19411,N_18184);
nand U22436 (N_22436,N_18514,N_20770);
and U22437 (N_22437,N_19413,N_20160);
xnor U22438 (N_22438,N_20136,N_18752);
or U22439 (N_22439,N_19503,N_19905);
nand U22440 (N_22440,N_20481,N_19154);
nand U22441 (N_22441,N_18011,N_20570);
or U22442 (N_22442,N_18868,N_18062);
nand U22443 (N_22443,N_18343,N_20037);
xor U22444 (N_22444,N_20947,N_18271);
or U22445 (N_22445,N_19424,N_20962);
or U22446 (N_22446,N_18891,N_20654);
nand U22447 (N_22447,N_19960,N_19496);
nor U22448 (N_22448,N_18879,N_20261);
nor U22449 (N_22449,N_19483,N_20742);
xor U22450 (N_22450,N_20020,N_20390);
or U22451 (N_22451,N_18987,N_20600);
nor U22452 (N_22452,N_19235,N_20195);
and U22453 (N_22453,N_19270,N_20247);
nor U22454 (N_22454,N_18109,N_18208);
nand U22455 (N_22455,N_19460,N_19558);
xnor U22456 (N_22456,N_18088,N_19147);
or U22457 (N_22457,N_18707,N_20170);
xor U22458 (N_22458,N_18003,N_18759);
and U22459 (N_22459,N_20159,N_20614);
xnor U22460 (N_22460,N_18965,N_20406);
nand U22461 (N_22461,N_18553,N_19009);
nand U22462 (N_22462,N_18854,N_18910);
and U22463 (N_22463,N_20586,N_20821);
or U22464 (N_22464,N_19780,N_18611);
xnor U22465 (N_22465,N_19473,N_19252);
or U22466 (N_22466,N_19329,N_18855);
nor U22467 (N_22467,N_20490,N_19016);
nand U22468 (N_22468,N_20296,N_18973);
nand U22469 (N_22469,N_19450,N_20215);
nor U22470 (N_22470,N_19379,N_19463);
xnor U22471 (N_22471,N_18598,N_18493);
and U22472 (N_22472,N_19420,N_19710);
nor U22473 (N_22473,N_19950,N_18080);
or U22474 (N_22474,N_18078,N_18093);
or U22475 (N_22475,N_20691,N_20229);
or U22476 (N_22476,N_20464,N_18189);
xnor U22477 (N_22477,N_19453,N_20087);
xnor U22478 (N_22478,N_18412,N_20718);
or U22479 (N_22479,N_19750,N_18797);
or U22480 (N_22480,N_20129,N_18578);
nor U22481 (N_22481,N_18446,N_19682);
nand U22482 (N_22482,N_18642,N_19610);
nor U22483 (N_22483,N_18981,N_20533);
nand U22484 (N_22484,N_19326,N_18631);
nand U22485 (N_22485,N_20527,N_18808);
xnor U22486 (N_22486,N_19882,N_20656);
xnor U22487 (N_22487,N_18201,N_18419);
nand U22488 (N_22488,N_20174,N_18239);
nor U22489 (N_22489,N_18041,N_18102);
nand U22490 (N_22490,N_18748,N_20536);
nor U22491 (N_22491,N_18469,N_18438);
xnor U22492 (N_22492,N_18034,N_20830);
or U22493 (N_22493,N_19538,N_19918);
or U22494 (N_22494,N_20462,N_18028);
xnor U22495 (N_22495,N_18628,N_19828);
nand U22496 (N_22496,N_18920,N_18775);
xnor U22497 (N_22497,N_19811,N_18862);
nand U22498 (N_22498,N_18022,N_18715);
or U22499 (N_22499,N_19406,N_19819);
nor U22500 (N_22500,N_18243,N_18977);
nor U22501 (N_22501,N_20880,N_19877);
nor U22502 (N_22502,N_18558,N_20297);
and U22503 (N_22503,N_19512,N_20354);
or U22504 (N_22504,N_20518,N_18927);
and U22505 (N_22505,N_19910,N_20455);
xor U22506 (N_22506,N_18714,N_20857);
nand U22507 (N_22507,N_19181,N_18157);
nor U22508 (N_22508,N_19105,N_19122);
nor U22509 (N_22509,N_19199,N_18625);
or U22510 (N_22510,N_19118,N_20829);
and U22511 (N_22511,N_20622,N_18246);
or U22512 (N_22512,N_19273,N_19337);
nand U22513 (N_22513,N_20815,N_19040);
and U22514 (N_22514,N_20483,N_19295);
or U22515 (N_22515,N_20537,N_20612);
nor U22516 (N_22516,N_19457,N_19734);
and U22517 (N_22517,N_19399,N_20616);
xor U22518 (N_22518,N_20299,N_20469);
and U22519 (N_22519,N_20043,N_19657);
nand U22520 (N_22520,N_19656,N_19181);
or U22521 (N_22521,N_20109,N_20396);
and U22522 (N_22522,N_19632,N_19320);
xnor U22523 (N_22523,N_19520,N_18993);
nand U22524 (N_22524,N_19444,N_20032);
nor U22525 (N_22525,N_20383,N_20334);
xnor U22526 (N_22526,N_19312,N_19834);
nor U22527 (N_22527,N_19898,N_20924);
or U22528 (N_22528,N_20872,N_18306);
nand U22529 (N_22529,N_20966,N_18048);
nand U22530 (N_22530,N_19081,N_18983);
xor U22531 (N_22531,N_18724,N_20615);
xnor U22532 (N_22532,N_19110,N_20572);
and U22533 (N_22533,N_20853,N_18345);
and U22534 (N_22534,N_20211,N_18002);
nand U22535 (N_22535,N_19746,N_20344);
xor U22536 (N_22536,N_18718,N_20818);
xor U22537 (N_22537,N_19838,N_18298);
nor U22538 (N_22538,N_19197,N_18639);
nor U22539 (N_22539,N_19972,N_19883);
nand U22540 (N_22540,N_19283,N_20540);
nor U22541 (N_22541,N_18402,N_18876);
or U22542 (N_22542,N_20855,N_20607);
nor U22543 (N_22543,N_18587,N_19305);
nor U22544 (N_22544,N_19434,N_20795);
and U22545 (N_22545,N_20184,N_20704);
or U22546 (N_22546,N_18227,N_20393);
xor U22547 (N_22547,N_19680,N_19158);
nand U22548 (N_22548,N_18105,N_19782);
nor U22549 (N_22549,N_19285,N_20020);
xor U22550 (N_22550,N_20444,N_18172);
xnor U22551 (N_22551,N_19563,N_18258);
or U22552 (N_22552,N_20868,N_20061);
and U22553 (N_22553,N_20266,N_20942);
nor U22554 (N_22554,N_19903,N_20001);
or U22555 (N_22555,N_20672,N_20144);
or U22556 (N_22556,N_20681,N_19968);
nor U22557 (N_22557,N_20053,N_18175);
nand U22558 (N_22558,N_20688,N_19933);
or U22559 (N_22559,N_18135,N_20999);
nand U22560 (N_22560,N_19569,N_18142);
nand U22561 (N_22561,N_18695,N_20517);
nor U22562 (N_22562,N_19508,N_18392);
nand U22563 (N_22563,N_20899,N_20977);
nand U22564 (N_22564,N_18286,N_18753);
xnor U22565 (N_22565,N_18399,N_18030);
xnor U22566 (N_22566,N_19176,N_20529);
xor U22567 (N_22567,N_18570,N_18329);
and U22568 (N_22568,N_19797,N_19020);
nor U22569 (N_22569,N_19729,N_18481);
xor U22570 (N_22570,N_18568,N_18522);
nor U22571 (N_22571,N_19067,N_20425);
xor U22572 (N_22572,N_18193,N_19633);
or U22573 (N_22573,N_18320,N_18802);
nor U22574 (N_22574,N_19029,N_20260);
or U22575 (N_22575,N_18769,N_18696);
nor U22576 (N_22576,N_18441,N_19226);
and U22577 (N_22577,N_20677,N_18298);
nand U22578 (N_22578,N_20142,N_19913);
xor U22579 (N_22579,N_18797,N_20955);
and U22580 (N_22580,N_20054,N_20092);
and U22581 (N_22581,N_19349,N_18925);
nor U22582 (N_22582,N_19407,N_20295);
and U22583 (N_22583,N_18008,N_18955);
nand U22584 (N_22584,N_19995,N_19977);
nand U22585 (N_22585,N_18685,N_18709);
and U22586 (N_22586,N_18235,N_20539);
or U22587 (N_22587,N_20018,N_19370);
xnor U22588 (N_22588,N_20150,N_18851);
nand U22589 (N_22589,N_18878,N_20045);
xor U22590 (N_22590,N_20945,N_20476);
and U22591 (N_22591,N_19935,N_19647);
nor U22592 (N_22592,N_20069,N_19211);
or U22593 (N_22593,N_19345,N_18282);
nand U22594 (N_22594,N_20294,N_20990);
and U22595 (N_22595,N_18213,N_18386);
or U22596 (N_22596,N_18457,N_19527);
or U22597 (N_22597,N_19724,N_19574);
xnor U22598 (N_22598,N_18457,N_20001);
nor U22599 (N_22599,N_19052,N_19282);
or U22600 (N_22600,N_20070,N_18453);
and U22601 (N_22601,N_18319,N_20233);
nor U22602 (N_22602,N_18128,N_18497);
or U22603 (N_22603,N_19584,N_18467);
nand U22604 (N_22604,N_19147,N_20174);
nand U22605 (N_22605,N_19529,N_19115);
nor U22606 (N_22606,N_18778,N_20053);
nand U22607 (N_22607,N_18043,N_18936);
xor U22608 (N_22608,N_18866,N_18578);
and U22609 (N_22609,N_19179,N_20742);
and U22610 (N_22610,N_18539,N_19605);
and U22611 (N_22611,N_19279,N_19209);
nor U22612 (N_22612,N_18077,N_18662);
and U22613 (N_22613,N_20243,N_20701);
nor U22614 (N_22614,N_19083,N_19837);
nor U22615 (N_22615,N_19998,N_20525);
and U22616 (N_22616,N_19583,N_20251);
or U22617 (N_22617,N_20871,N_19541);
nand U22618 (N_22618,N_18265,N_18993);
nor U22619 (N_22619,N_18126,N_19503);
xnor U22620 (N_22620,N_20337,N_18814);
nand U22621 (N_22621,N_20346,N_20531);
nor U22622 (N_22622,N_19389,N_20319);
and U22623 (N_22623,N_19600,N_19480);
and U22624 (N_22624,N_19641,N_19398);
xnor U22625 (N_22625,N_18608,N_20163);
or U22626 (N_22626,N_20285,N_18935);
xnor U22627 (N_22627,N_19156,N_20302);
or U22628 (N_22628,N_19541,N_19275);
nor U22629 (N_22629,N_19766,N_18553);
nor U22630 (N_22630,N_20697,N_19040);
or U22631 (N_22631,N_20879,N_18383);
and U22632 (N_22632,N_18159,N_19866);
or U22633 (N_22633,N_20498,N_20536);
nand U22634 (N_22634,N_19013,N_18742);
nand U22635 (N_22635,N_18493,N_20615);
nand U22636 (N_22636,N_19374,N_19297);
xor U22637 (N_22637,N_20633,N_20308);
nand U22638 (N_22638,N_20407,N_19484);
and U22639 (N_22639,N_20790,N_20804);
nor U22640 (N_22640,N_19922,N_19876);
and U22641 (N_22641,N_18012,N_18828);
or U22642 (N_22642,N_20557,N_19010);
and U22643 (N_22643,N_20051,N_19239);
or U22644 (N_22644,N_20905,N_18834);
nand U22645 (N_22645,N_18275,N_18562);
or U22646 (N_22646,N_19150,N_18252);
xor U22647 (N_22647,N_18363,N_19542);
or U22648 (N_22648,N_18974,N_18931);
and U22649 (N_22649,N_20962,N_19705);
nor U22650 (N_22650,N_18778,N_19772);
xor U22651 (N_22651,N_20139,N_18569);
nor U22652 (N_22652,N_20836,N_18544);
xnor U22653 (N_22653,N_20525,N_20383);
nor U22654 (N_22654,N_20752,N_19906);
nor U22655 (N_22655,N_19430,N_20222);
or U22656 (N_22656,N_20997,N_18069);
and U22657 (N_22657,N_19966,N_18334);
nand U22658 (N_22658,N_18317,N_20588);
nand U22659 (N_22659,N_19629,N_20868);
and U22660 (N_22660,N_18958,N_20080);
nand U22661 (N_22661,N_18703,N_19472);
or U22662 (N_22662,N_20858,N_19159);
nand U22663 (N_22663,N_19937,N_20644);
nor U22664 (N_22664,N_20233,N_20833);
xnor U22665 (N_22665,N_18524,N_19666);
or U22666 (N_22666,N_19520,N_19060);
nand U22667 (N_22667,N_18488,N_18557);
nand U22668 (N_22668,N_18001,N_20375);
or U22669 (N_22669,N_18759,N_20402);
and U22670 (N_22670,N_19893,N_20642);
and U22671 (N_22671,N_18374,N_19868);
nand U22672 (N_22672,N_20606,N_20580);
and U22673 (N_22673,N_18957,N_18054);
nand U22674 (N_22674,N_18131,N_20841);
nand U22675 (N_22675,N_19582,N_18313);
and U22676 (N_22676,N_20100,N_20692);
xor U22677 (N_22677,N_20778,N_19421);
nor U22678 (N_22678,N_20616,N_19058);
and U22679 (N_22679,N_20294,N_18075);
nor U22680 (N_22680,N_20780,N_20195);
xor U22681 (N_22681,N_20722,N_18322);
nand U22682 (N_22682,N_18603,N_20791);
xnor U22683 (N_22683,N_20286,N_18504);
nand U22684 (N_22684,N_18461,N_18603);
or U22685 (N_22685,N_18449,N_18249);
and U22686 (N_22686,N_18860,N_20027);
and U22687 (N_22687,N_19476,N_18864);
nand U22688 (N_22688,N_18673,N_20501);
and U22689 (N_22689,N_19909,N_19579);
nor U22690 (N_22690,N_20395,N_18870);
xnor U22691 (N_22691,N_19996,N_18762);
or U22692 (N_22692,N_19886,N_20644);
nor U22693 (N_22693,N_19435,N_18562);
and U22694 (N_22694,N_19383,N_19815);
nand U22695 (N_22695,N_20925,N_20917);
nor U22696 (N_22696,N_19754,N_18864);
and U22697 (N_22697,N_19601,N_20520);
nor U22698 (N_22698,N_18582,N_19763);
xor U22699 (N_22699,N_18467,N_20481);
and U22700 (N_22700,N_18597,N_18569);
or U22701 (N_22701,N_18047,N_19480);
xnor U22702 (N_22702,N_18319,N_20998);
or U22703 (N_22703,N_19124,N_20093);
nor U22704 (N_22704,N_20405,N_20048);
nand U22705 (N_22705,N_18261,N_18718);
and U22706 (N_22706,N_19407,N_20802);
nor U22707 (N_22707,N_19006,N_20709);
or U22708 (N_22708,N_20629,N_20958);
and U22709 (N_22709,N_19282,N_19620);
nor U22710 (N_22710,N_19109,N_19210);
or U22711 (N_22711,N_20894,N_19305);
nor U22712 (N_22712,N_19445,N_19308);
and U22713 (N_22713,N_20432,N_20733);
nor U22714 (N_22714,N_18556,N_20402);
and U22715 (N_22715,N_18234,N_18200);
xor U22716 (N_22716,N_19668,N_18181);
nand U22717 (N_22717,N_19634,N_20718);
nand U22718 (N_22718,N_18144,N_20495);
or U22719 (N_22719,N_20703,N_20877);
xnor U22720 (N_22720,N_20779,N_20571);
xnor U22721 (N_22721,N_19033,N_19878);
and U22722 (N_22722,N_20230,N_19536);
xor U22723 (N_22723,N_18306,N_18440);
nand U22724 (N_22724,N_20453,N_19682);
xor U22725 (N_22725,N_19789,N_20410);
nor U22726 (N_22726,N_18330,N_19705);
nor U22727 (N_22727,N_20508,N_18931);
or U22728 (N_22728,N_19815,N_20837);
xor U22729 (N_22729,N_19930,N_20379);
nand U22730 (N_22730,N_20842,N_18687);
xor U22731 (N_22731,N_20273,N_18753);
and U22732 (N_22732,N_19857,N_20023);
xor U22733 (N_22733,N_18855,N_19977);
xnor U22734 (N_22734,N_20381,N_19139);
and U22735 (N_22735,N_20779,N_18522);
xnor U22736 (N_22736,N_20329,N_19038);
xnor U22737 (N_22737,N_19482,N_20723);
or U22738 (N_22738,N_20398,N_20963);
or U22739 (N_22739,N_19750,N_19610);
or U22740 (N_22740,N_19541,N_18144);
and U22741 (N_22741,N_18182,N_20917);
nand U22742 (N_22742,N_19362,N_18247);
or U22743 (N_22743,N_20434,N_18392);
nor U22744 (N_22744,N_18536,N_20809);
nor U22745 (N_22745,N_18295,N_19203);
and U22746 (N_22746,N_19925,N_20546);
nor U22747 (N_22747,N_18783,N_20822);
or U22748 (N_22748,N_18031,N_19412);
nand U22749 (N_22749,N_20864,N_20184);
and U22750 (N_22750,N_19871,N_19452);
nand U22751 (N_22751,N_18588,N_18853);
nand U22752 (N_22752,N_18614,N_18172);
nand U22753 (N_22753,N_18546,N_20469);
and U22754 (N_22754,N_20309,N_18774);
or U22755 (N_22755,N_18344,N_19883);
nand U22756 (N_22756,N_18421,N_20388);
or U22757 (N_22757,N_18344,N_19045);
xor U22758 (N_22758,N_19462,N_18374);
or U22759 (N_22759,N_19774,N_20759);
and U22760 (N_22760,N_19617,N_18100);
nor U22761 (N_22761,N_20011,N_19647);
and U22762 (N_22762,N_18190,N_19519);
and U22763 (N_22763,N_18051,N_20555);
or U22764 (N_22764,N_19092,N_18576);
nor U22765 (N_22765,N_20717,N_19492);
or U22766 (N_22766,N_20676,N_19614);
or U22767 (N_22767,N_20120,N_19795);
nand U22768 (N_22768,N_18972,N_20723);
xnor U22769 (N_22769,N_18989,N_18005);
nor U22770 (N_22770,N_18738,N_20960);
or U22771 (N_22771,N_18494,N_19536);
nor U22772 (N_22772,N_18267,N_20056);
nand U22773 (N_22773,N_20958,N_20094);
xnor U22774 (N_22774,N_19296,N_20672);
nand U22775 (N_22775,N_20113,N_19567);
and U22776 (N_22776,N_18212,N_20301);
or U22777 (N_22777,N_18964,N_19086);
and U22778 (N_22778,N_19107,N_19465);
xnor U22779 (N_22779,N_19918,N_19719);
nor U22780 (N_22780,N_19610,N_20696);
nand U22781 (N_22781,N_20174,N_19748);
or U22782 (N_22782,N_18110,N_18672);
and U22783 (N_22783,N_18849,N_19090);
nand U22784 (N_22784,N_18109,N_20987);
nor U22785 (N_22785,N_18949,N_20329);
or U22786 (N_22786,N_18082,N_19214);
or U22787 (N_22787,N_20439,N_20768);
and U22788 (N_22788,N_20832,N_19878);
and U22789 (N_22789,N_19278,N_20471);
xor U22790 (N_22790,N_20148,N_18227);
and U22791 (N_22791,N_19192,N_18678);
nor U22792 (N_22792,N_20137,N_18569);
nor U22793 (N_22793,N_20476,N_18734);
or U22794 (N_22794,N_19705,N_20228);
or U22795 (N_22795,N_19774,N_19437);
nand U22796 (N_22796,N_18759,N_19129);
nor U22797 (N_22797,N_19372,N_19947);
or U22798 (N_22798,N_20453,N_20813);
xor U22799 (N_22799,N_19578,N_20625);
nand U22800 (N_22800,N_19653,N_19163);
or U22801 (N_22801,N_18635,N_18759);
nand U22802 (N_22802,N_18525,N_19759);
xor U22803 (N_22803,N_18190,N_20505);
nor U22804 (N_22804,N_18361,N_18185);
nor U22805 (N_22805,N_20429,N_19413);
nand U22806 (N_22806,N_20749,N_20368);
or U22807 (N_22807,N_19694,N_20773);
nand U22808 (N_22808,N_20553,N_18484);
nand U22809 (N_22809,N_19375,N_20349);
nand U22810 (N_22810,N_20357,N_19234);
and U22811 (N_22811,N_20499,N_18026);
and U22812 (N_22812,N_20318,N_20870);
nand U22813 (N_22813,N_19917,N_19646);
xor U22814 (N_22814,N_20239,N_18140);
and U22815 (N_22815,N_20127,N_20926);
nand U22816 (N_22816,N_19829,N_19828);
or U22817 (N_22817,N_18955,N_18204);
and U22818 (N_22818,N_18733,N_19577);
xor U22819 (N_22819,N_18825,N_18580);
or U22820 (N_22820,N_19719,N_18666);
or U22821 (N_22821,N_20846,N_18711);
and U22822 (N_22822,N_20224,N_20756);
or U22823 (N_22823,N_20481,N_19237);
xor U22824 (N_22824,N_18581,N_19716);
nor U22825 (N_22825,N_19977,N_19984);
or U22826 (N_22826,N_18374,N_19694);
nor U22827 (N_22827,N_19160,N_19814);
nor U22828 (N_22828,N_19228,N_20189);
or U22829 (N_22829,N_20471,N_19143);
nor U22830 (N_22830,N_19163,N_19845);
xor U22831 (N_22831,N_20111,N_20244);
nor U22832 (N_22832,N_18734,N_20272);
or U22833 (N_22833,N_20764,N_19836);
nor U22834 (N_22834,N_19040,N_18679);
or U22835 (N_22835,N_19870,N_20289);
and U22836 (N_22836,N_20724,N_18774);
and U22837 (N_22837,N_20030,N_19864);
and U22838 (N_22838,N_20675,N_18630);
nand U22839 (N_22839,N_18252,N_19464);
nand U22840 (N_22840,N_20009,N_19531);
xor U22841 (N_22841,N_19240,N_20594);
nor U22842 (N_22842,N_19012,N_19951);
nand U22843 (N_22843,N_18607,N_19127);
nor U22844 (N_22844,N_20420,N_18163);
and U22845 (N_22845,N_18997,N_19721);
and U22846 (N_22846,N_20046,N_18936);
nand U22847 (N_22847,N_20527,N_18279);
nor U22848 (N_22848,N_20602,N_19983);
xor U22849 (N_22849,N_18136,N_18016);
nand U22850 (N_22850,N_20889,N_19302);
and U22851 (N_22851,N_20102,N_18465);
xor U22852 (N_22852,N_20106,N_20703);
nor U22853 (N_22853,N_20693,N_18359);
nand U22854 (N_22854,N_18395,N_19263);
or U22855 (N_22855,N_20885,N_19324);
xnor U22856 (N_22856,N_18774,N_20008);
nor U22857 (N_22857,N_19210,N_20231);
xor U22858 (N_22858,N_19840,N_20409);
or U22859 (N_22859,N_20632,N_19888);
or U22860 (N_22860,N_18238,N_20061);
or U22861 (N_22861,N_18336,N_20730);
nand U22862 (N_22862,N_20365,N_20403);
nor U22863 (N_22863,N_18555,N_18648);
and U22864 (N_22864,N_20980,N_18226);
and U22865 (N_22865,N_20137,N_20601);
nand U22866 (N_22866,N_20991,N_18257);
nor U22867 (N_22867,N_19452,N_19409);
or U22868 (N_22868,N_18026,N_19558);
or U22869 (N_22869,N_19955,N_18294);
nor U22870 (N_22870,N_19444,N_19835);
nand U22871 (N_22871,N_19636,N_18877);
nand U22872 (N_22872,N_20390,N_19596);
nor U22873 (N_22873,N_20185,N_20621);
and U22874 (N_22874,N_20589,N_19128);
and U22875 (N_22875,N_18157,N_18680);
xnor U22876 (N_22876,N_19738,N_19221);
xnor U22877 (N_22877,N_18707,N_20609);
xnor U22878 (N_22878,N_20373,N_20039);
nor U22879 (N_22879,N_19377,N_18367);
nand U22880 (N_22880,N_18070,N_20583);
nand U22881 (N_22881,N_19877,N_18307);
and U22882 (N_22882,N_19372,N_19016);
and U22883 (N_22883,N_18568,N_19520);
nor U22884 (N_22884,N_19179,N_19067);
xor U22885 (N_22885,N_20813,N_18548);
nor U22886 (N_22886,N_18004,N_19952);
nand U22887 (N_22887,N_19244,N_19746);
and U22888 (N_22888,N_20675,N_18636);
or U22889 (N_22889,N_18473,N_18061);
nand U22890 (N_22890,N_18228,N_20448);
nor U22891 (N_22891,N_19614,N_19920);
nand U22892 (N_22892,N_18545,N_19782);
nand U22893 (N_22893,N_20919,N_20054);
nand U22894 (N_22894,N_18215,N_20997);
xor U22895 (N_22895,N_20251,N_20818);
or U22896 (N_22896,N_20542,N_18011);
nor U22897 (N_22897,N_20180,N_20726);
nand U22898 (N_22898,N_19073,N_18492);
and U22899 (N_22899,N_18565,N_19586);
nor U22900 (N_22900,N_18917,N_18439);
xnor U22901 (N_22901,N_20566,N_19690);
nand U22902 (N_22902,N_18689,N_18990);
xor U22903 (N_22903,N_20862,N_18297);
xnor U22904 (N_22904,N_19384,N_19498);
xnor U22905 (N_22905,N_18480,N_19244);
or U22906 (N_22906,N_18256,N_18703);
or U22907 (N_22907,N_18820,N_20208);
and U22908 (N_22908,N_20505,N_19766);
nor U22909 (N_22909,N_20825,N_20286);
nor U22910 (N_22910,N_19131,N_18490);
or U22911 (N_22911,N_19920,N_18992);
nor U22912 (N_22912,N_19615,N_18722);
nand U22913 (N_22913,N_20544,N_18002);
nand U22914 (N_22914,N_19800,N_19778);
or U22915 (N_22915,N_18636,N_20472);
nand U22916 (N_22916,N_18254,N_18481);
nand U22917 (N_22917,N_19423,N_20350);
xor U22918 (N_22918,N_18782,N_18839);
xnor U22919 (N_22919,N_18155,N_20822);
nor U22920 (N_22920,N_20600,N_19841);
nor U22921 (N_22921,N_18295,N_19057);
nor U22922 (N_22922,N_19198,N_19637);
nor U22923 (N_22923,N_18127,N_19335);
nor U22924 (N_22924,N_19652,N_19232);
xnor U22925 (N_22925,N_19684,N_18235);
xor U22926 (N_22926,N_18498,N_18843);
and U22927 (N_22927,N_19955,N_20482);
xor U22928 (N_22928,N_20519,N_19637);
xnor U22929 (N_22929,N_19216,N_18817);
nand U22930 (N_22930,N_18934,N_20437);
or U22931 (N_22931,N_20944,N_20421);
xor U22932 (N_22932,N_19892,N_20151);
and U22933 (N_22933,N_19156,N_20807);
xnor U22934 (N_22934,N_20462,N_19971);
nand U22935 (N_22935,N_19862,N_18599);
nand U22936 (N_22936,N_18253,N_20477);
or U22937 (N_22937,N_18052,N_19995);
or U22938 (N_22938,N_19121,N_18907);
xnor U22939 (N_22939,N_19021,N_19833);
or U22940 (N_22940,N_20557,N_18183);
nand U22941 (N_22941,N_19428,N_20367);
nor U22942 (N_22942,N_19385,N_18798);
xnor U22943 (N_22943,N_18875,N_19297);
nor U22944 (N_22944,N_19164,N_18892);
nand U22945 (N_22945,N_20742,N_19225);
nand U22946 (N_22946,N_20778,N_20110);
nor U22947 (N_22947,N_19255,N_20393);
xor U22948 (N_22948,N_19795,N_18134);
nand U22949 (N_22949,N_19951,N_18142);
and U22950 (N_22950,N_20183,N_18743);
xnor U22951 (N_22951,N_18675,N_18674);
or U22952 (N_22952,N_20908,N_20337);
xor U22953 (N_22953,N_18287,N_18835);
or U22954 (N_22954,N_20454,N_20036);
and U22955 (N_22955,N_20323,N_18281);
or U22956 (N_22956,N_20099,N_19162);
nand U22957 (N_22957,N_20284,N_20998);
xor U22958 (N_22958,N_18878,N_19877);
and U22959 (N_22959,N_19146,N_18435);
or U22960 (N_22960,N_18914,N_18803);
or U22961 (N_22961,N_20337,N_18131);
nand U22962 (N_22962,N_19222,N_19207);
or U22963 (N_22963,N_20330,N_19252);
nand U22964 (N_22964,N_19134,N_19171);
or U22965 (N_22965,N_19872,N_19157);
or U22966 (N_22966,N_20020,N_18401);
nand U22967 (N_22967,N_18326,N_20786);
and U22968 (N_22968,N_20927,N_18945);
and U22969 (N_22969,N_19630,N_19762);
or U22970 (N_22970,N_18456,N_19613);
xor U22971 (N_22971,N_20555,N_20112);
xor U22972 (N_22972,N_19424,N_19785);
nor U22973 (N_22973,N_18427,N_18990);
nand U22974 (N_22974,N_18232,N_18627);
nor U22975 (N_22975,N_18036,N_20606);
nor U22976 (N_22976,N_19406,N_19718);
nand U22977 (N_22977,N_20885,N_20781);
and U22978 (N_22978,N_19441,N_20332);
xor U22979 (N_22979,N_20924,N_18665);
nor U22980 (N_22980,N_20780,N_18006);
nand U22981 (N_22981,N_20078,N_19857);
nor U22982 (N_22982,N_20036,N_20533);
xnor U22983 (N_22983,N_18485,N_20666);
nand U22984 (N_22984,N_18654,N_19062);
nor U22985 (N_22985,N_19049,N_20320);
nand U22986 (N_22986,N_19999,N_19043);
nand U22987 (N_22987,N_19380,N_18400);
xnor U22988 (N_22988,N_20212,N_19567);
or U22989 (N_22989,N_18974,N_20012);
xor U22990 (N_22990,N_18430,N_18562);
and U22991 (N_22991,N_18372,N_18410);
nor U22992 (N_22992,N_18712,N_19509);
xor U22993 (N_22993,N_19270,N_18044);
and U22994 (N_22994,N_19296,N_19114);
or U22995 (N_22995,N_18684,N_18569);
nand U22996 (N_22996,N_19264,N_18519);
or U22997 (N_22997,N_18574,N_19039);
xor U22998 (N_22998,N_19372,N_19620);
or U22999 (N_22999,N_19633,N_19437);
nand U23000 (N_23000,N_20782,N_20156);
or U23001 (N_23001,N_20916,N_18494);
nand U23002 (N_23002,N_18647,N_20823);
and U23003 (N_23003,N_20192,N_19045);
or U23004 (N_23004,N_20956,N_19089);
nor U23005 (N_23005,N_19850,N_19200);
or U23006 (N_23006,N_20478,N_20423);
and U23007 (N_23007,N_18880,N_18479);
or U23008 (N_23008,N_20548,N_19607);
and U23009 (N_23009,N_19273,N_18718);
nor U23010 (N_23010,N_20815,N_20366);
nor U23011 (N_23011,N_18735,N_19697);
nand U23012 (N_23012,N_20860,N_19842);
or U23013 (N_23013,N_19798,N_18210);
xnor U23014 (N_23014,N_18253,N_20768);
nand U23015 (N_23015,N_19587,N_19519);
nor U23016 (N_23016,N_19081,N_19839);
nand U23017 (N_23017,N_19584,N_20736);
and U23018 (N_23018,N_20754,N_18120);
xnor U23019 (N_23019,N_18801,N_20568);
nor U23020 (N_23020,N_20034,N_20586);
nand U23021 (N_23021,N_18102,N_19749);
and U23022 (N_23022,N_18892,N_20872);
or U23023 (N_23023,N_18895,N_18083);
or U23024 (N_23024,N_18101,N_18291);
and U23025 (N_23025,N_19806,N_19444);
nand U23026 (N_23026,N_18482,N_19470);
and U23027 (N_23027,N_19683,N_19216);
nor U23028 (N_23028,N_18697,N_20834);
xor U23029 (N_23029,N_19624,N_20581);
or U23030 (N_23030,N_20945,N_20537);
xor U23031 (N_23031,N_20423,N_19404);
nand U23032 (N_23032,N_18117,N_19025);
or U23033 (N_23033,N_20169,N_18226);
xor U23034 (N_23034,N_19536,N_18826);
nand U23035 (N_23035,N_19344,N_18287);
nor U23036 (N_23036,N_18352,N_19047);
and U23037 (N_23037,N_18517,N_19958);
and U23038 (N_23038,N_20094,N_18025);
xnor U23039 (N_23039,N_19416,N_20809);
nor U23040 (N_23040,N_20588,N_18661);
or U23041 (N_23041,N_20449,N_19978);
nand U23042 (N_23042,N_19766,N_19323);
xnor U23043 (N_23043,N_19409,N_20953);
and U23044 (N_23044,N_19078,N_19145);
and U23045 (N_23045,N_18155,N_20677);
xnor U23046 (N_23046,N_18087,N_19360);
or U23047 (N_23047,N_20879,N_18343);
nor U23048 (N_23048,N_20827,N_20015);
or U23049 (N_23049,N_20501,N_18478);
nor U23050 (N_23050,N_20841,N_19171);
and U23051 (N_23051,N_20867,N_19583);
and U23052 (N_23052,N_19313,N_20518);
and U23053 (N_23053,N_20126,N_18141);
and U23054 (N_23054,N_18830,N_19826);
nor U23055 (N_23055,N_18904,N_20749);
and U23056 (N_23056,N_20729,N_20787);
xor U23057 (N_23057,N_20916,N_19598);
nor U23058 (N_23058,N_20276,N_20079);
and U23059 (N_23059,N_18354,N_19047);
nor U23060 (N_23060,N_18735,N_18247);
nand U23061 (N_23061,N_20269,N_19707);
nand U23062 (N_23062,N_18001,N_18518);
xor U23063 (N_23063,N_19335,N_18744);
and U23064 (N_23064,N_19499,N_20548);
xor U23065 (N_23065,N_19023,N_18072);
nor U23066 (N_23066,N_20647,N_19191);
or U23067 (N_23067,N_18800,N_18301);
xor U23068 (N_23068,N_18861,N_18359);
nand U23069 (N_23069,N_20336,N_20361);
or U23070 (N_23070,N_19569,N_18847);
nor U23071 (N_23071,N_19256,N_20077);
and U23072 (N_23072,N_19598,N_20941);
nand U23073 (N_23073,N_18790,N_20816);
xor U23074 (N_23074,N_18606,N_19879);
xor U23075 (N_23075,N_18032,N_19661);
nor U23076 (N_23076,N_18396,N_19726);
or U23077 (N_23077,N_18497,N_20878);
and U23078 (N_23078,N_19548,N_18720);
and U23079 (N_23079,N_18246,N_19905);
or U23080 (N_23080,N_19611,N_18928);
xor U23081 (N_23081,N_19743,N_18397);
or U23082 (N_23082,N_19549,N_18932);
and U23083 (N_23083,N_19714,N_19258);
xor U23084 (N_23084,N_19235,N_18107);
and U23085 (N_23085,N_18501,N_20586);
xnor U23086 (N_23086,N_18510,N_18969);
nand U23087 (N_23087,N_20473,N_20652);
nand U23088 (N_23088,N_20475,N_18339);
and U23089 (N_23089,N_20152,N_19066);
xor U23090 (N_23090,N_19374,N_20496);
nand U23091 (N_23091,N_19419,N_19819);
and U23092 (N_23092,N_20347,N_18565);
or U23093 (N_23093,N_19033,N_20614);
and U23094 (N_23094,N_19037,N_19011);
nand U23095 (N_23095,N_20771,N_18585);
nand U23096 (N_23096,N_20998,N_18316);
and U23097 (N_23097,N_20258,N_18220);
nand U23098 (N_23098,N_18095,N_19130);
nor U23099 (N_23099,N_18050,N_19810);
or U23100 (N_23100,N_19947,N_20166);
nor U23101 (N_23101,N_20725,N_18385);
or U23102 (N_23102,N_18425,N_18374);
nand U23103 (N_23103,N_18985,N_18145);
nor U23104 (N_23104,N_18511,N_19475);
and U23105 (N_23105,N_18870,N_19580);
nor U23106 (N_23106,N_18130,N_19331);
nor U23107 (N_23107,N_18092,N_20405);
or U23108 (N_23108,N_19403,N_19600);
nor U23109 (N_23109,N_19547,N_20861);
nand U23110 (N_23110,N_18367,N_19380);
and U23111 (N_23111,N_18277,N_19409);
xor U23112 (N_23112,N_20260,N_20379);
or U23113 (N_23113,N_20495,N_20252);
and U23114 (N_23114,N_18494,N_19621);
or U23115 (N_23115,N_18790,N_18218);
and U23116 (N_23116,N_20915,N_19397);
nand U23117 (N_23117,N_18125,N_19090);
or U23118 (N_23118,N_20101,N_20986);
nor U23119 (N_23119,N_20903,N_20807);
and U23120 (N_23120,N_20280,N_19302);
or U23121 (N_23121,N_18053,N_20634);
and U23122 (N_23122,N_20976,N_19172);
xnor U23123 (N_23123,N_20508,N_18527);
or U23124 (N_23124,N_18406,N_18505);
and U23125 (N_23125,N_20372,N_20244);
and U23126 (N_23126,N_18570,N_19090);
nand U23127 (N_23127,N_19895,N_19149);
or U23128 (N_23128,N_19001,N_20420);
nand U23129 (N_23129,N_18888,N_18277);
nor U23130 (N_23130,N_18150,N_20101);
nor U23131 (N_23131,N_20404,N_19331);
or U23132 (N_23132,N_20093,N_19654);
nand U23133 (N_23133,N_20797,N_20899);
and U23134 (N_23134,N_20385,N_20367);
and U23135 (N_23135,N_20488,N_18556);
nor U23136 (N_23136,N_19966,N_20221);
xnor U23137 (N_23137,N_20763,N_20931);
xnor U23138 (N_23138,N_20295,N_18533);
and U23139 (N_23139,N_18805,N_20201);
or U23140 (N_23140,N_20612,N_19031);
or U23141 (N_23141,N_18205,N_18973);
nor U23142 (N_23142,N_20325,N_20808);
nor U23143 (N_23143,N_19215,N_20277);
and U23144 (N_23144,N_18601,N_18584);
and U23145 (N_23145,N_20992,N_19412);
nand U23146 (N_23146,N_18546,N_20612);
nand U23147 (N_23147,N_18749,N_18005);
and U23148 (N_23148,N_20386,N_20153);
xor U23149 (N_23149,N_20285,N_19459);
nand U23150 (N_23150,N_19334,N_20964);
and U23151 (N_23151,N_18849,N_20148);
nor U23152 (N_23152,N_18700,N_19875);
and U23153 (N_23153,N_20378,N_20820);
and U23154 (N_23154,N_18796,N_18476);
nand U23155 (N_23155,N_19204,N_19717);
or U23156 (N_23156,N_18001,N_20866);
and U23157 (N_23157,N_20090,N_19624);
xor U23158 (N_23158,N_19974,N_20742);
nand U23159 (N_23159,N_18032,N_19166);
or U23160 (N_23160,N_19382,N_20716);
or U23161 (N_23161,N_18951,N_18619);
and U23162 (N_23162,N_19655,N_20422);
or U23163 (N_23163,N_18536,N_19962);
nand U23164 (N_23164,N_20813,N_20977);
xor U23165 (N_23165,N_20670,N_20654);
xnor U23166 (N_23166,N_18710,N_19495);
nor U23167 (N_23167,N_19790,N_20866);
and U23168 (N_23168,N_19341,N_18766);
nor U23169 (N_23169,N_19334,N_19273);
or U23170 (N_23170,N_19815,N_19166);
or U23171 (N_23171,N_18430,N_19896);
nand U23172 (N_23172,N_19897,N_20166);
or U23173 (N_23173,N_20160,N_19357);
or U23174 (N_23174,N_18050,N_18637);
xor U23175 (N_23175,N_20062,N_19627);
and U23176 (N_23176,N_19641,N_18842);
or U23177 (N_23177,N_18028,N_18848);
or U23178 (N_23178,N_20636,N_18562);
and U23179 (N_23179,N_19939,N_18710);
nor U23180 (N_23180,N_20472,N_20458);
or U23181 (N_23181,N_20310,N_18394);
nand U23182 (N_23182,N_20125,N_19339);
and U23183 (N_23183,N_20672,N_19041);
and U23184 (N_23184,N_19774,N_18912);
xor U23185 (N_23185,N_19195,N_18740);
xor U23186 (N_23186,N_19301,N_18203);
or U23187 (N_23187,N_19875,N_19076);
or U23188 (N_23188,N_20211,N_19837);
and U23189 (N_23189,N_18738,N_19418);
nand U23190 (N_23190,N_19899,N_19407);
nor U23191 (N_23191,N_18173,N_20291);
nor U23192 (N_23192,N_20336,N_20915);
nand U23193 (N_23193,N_19590,N_19563);
or U23194 (N_23194,N_19956,N_19140);
xnor U23195 (N_23195,N_19196,N_19685);
nor U23196 (N_23196,N_20667,N_18599);
nand U23197 (N_23197,N_18390,N_18705);
nand U23198 (N_23198,N_20071,N_19077);
xnor U23199 (N_23199,N_18698,N_18502);
xnor U23200 (N_23200,N_19899,N_18031);
nor U23201 (N_23201,N_19911,N_19635);
nand U23202 (N_23202,N_18137,N_18287);
and U23203 (N_23203,N_18622,N_18628);
xor U23204 (N_23204,N_19135,N_20060);
xnor U23205 (N_23205,N_18859,N_20881);
nor U23206 (N_23206,N_20585,N_18415);
nand U23207 (N_23207,N_18552,N_18638);
or U23208 (N_23208,N_19724,N_18159);
xnor U23209 (N_23209,N_19790,N_20744);
xor U23210 (N_23210,N_19423,N_19108);
and U23211 (N_23211,N_20064,N_20470);
or U23212 (N_23212,N_19028,N_18488);
and U23213 (N_23213,N_20611,N_19212);
xor U23214 (N_23214,N_19644,N_18883);
nand U23215 (N_23215,N_18208,N_19973);
or U23216 (N_23216,N_18936,N_20977);
xor U23217 (N_23217,N_18247,N_18570);
nand U23218 (N_23218,N_19376,N_20836);
xnor U23219 (N_23219,N_20777,N_19774);
and U23220 (N_23220,N_18020,N_19902);
or U23221 (N_23221,N_18773,N_20700);
or U23222 (N_23222,N_19784,N_19568);
or U23223 (N_23223,N_20317,N_19369);
and U23224 (N_23224,N_18191,N_20696);
or U23225 (N_23225,N_19790,N_18408);
and U23226 (N_23226,N_20127,N_19727);
or U23227 (N_23227,N_19872,N_18394);
nand U23228 (N_23228,N_20859,N_18382);
xor U23229 (N_23229,N_20386,N_19973);
nand U23230 (N_23230,N_20763,N_18889);
nand U23231 (N_23231,N_18708,N_19108);
and U23232 (N_23232,N_19781,N_18262);
nor U23233 (N_23233,N_20462,N_18555);
xnor U23234 (N_23234,N_20344,N_20487);
nand U23235 (N_23235,N_19201,N_19195);
nor U23236 (N_23236,N_20219,N_18388);
nand U23237 (N_23237,N_20268,N_18313);
nand U23238 (N_23238,N_19146,N_18995);
xor U23239 (N_23239,N_18645,N_18906);
and U23240 (N_23240,N_19902,N_18102);
nand U23241 (N_23241,N_18954,N_18039);
or U23242 (N_23242,N_18148,N_19677);
or U23243 (N_23243,N_20350,N_20430);
or U23244 (N_23244,N_19397,N_20851);
xor U23245 (N_23245,N_20368,N_20010);
and U23246 (N_23246,N_19913,N_18306);
or U23247 (N_23247,N_18163,N_19946);
nand U23248 (N_23248,N_19674,N_20864);
nor U23249 (N_23249,N_18756,N_18781);
and U23250 (N_23250,N_19939,N_18311);
nand U23251 (N_23251,N_19059,N_19169);
and U23252 (N_23252,N_20108,N_20818);
and U23253 (N_23253,N_19106,N_19427);
xor U23254 (N_23254,N_18864,N_20737);
and U23255 (N_23255,N_18312,N_19381);
nor U23256 (N_23256,N_18995,N_19420);
and U23257 (N_23257,N_19853,N_18317);
nand U23258 (N_23258,N_18747,N_18436);
xnor U23259 (N_23259,N_20481,N_20005);
and U23260 (N_23260,N_20109,N_20231);
or U23261 (N_23261,N_19133,N_20523);
nor U23262 (N_23262,N_20351,N_20973);
nor U23263 (N_23263,N_20366,N_19395);
nand U23264 (N_23264,N_18179,N_20164);
nor U23265 (N_23265,N_18439,N_18981);
and U23266 (N_23266,N_18372,N_19983);
or U23267 (N_23267,N_19479,N_20008);
nor U23268 (N_23268,N_20675,N_18038);
or U23269 (N_23269,N_19441,N_18832);
nand U23270 (N_23270,N_19547,N_18937);
or U23271 (N_23271,N_19010,N_20078);
and U23272 (N_23272,N_20097,N_20600);
xor U23273 (N_23273,N_20614,N_19514);
nor U23274 (N_23274,N_20661,N_19615);
xor U23275 (N_23275,N_20868,N_18749);
xnor U23276 (N_23276,N_18314,N_18839);
and U23277 (N_23277,N_20837,N_19773);
and U23278 (N_23278,N_18590,N_18491);
nor U23279 (N_23279,N_18706,N_19758);
or U23280 (N_23280,N_20180,N_19553);
xnor U23281 (N_23281,N_18137,N_19413);
nand U23282 (N_23282,N_19562,N_20206);
nand U23283 (N_23283,N_19804,N_18787);
and U23284 (N_23284,N_19052,N_18947);
nor U23285 (N_23285,N_19880,N_18032);
nand U23286 (N_23286,N_18592,N_19651);
nor U23287 (N_23287,N_19997,N_19454);
xor U23288 (N_23288,N_20922,N_19165);
nor U23289 (N_23289,N_19309,N_19391);
or U23290 (N_23290,N_19306,N_19315);
and U23291 (N_23291,N_19870,N_18027);
nor U23292 (N_23292,N_20210,N_18602);
and U23293 (N_23293,N_19660,N_20931);
nand U23294 (N_23294,N_18433,N_19478);
or U23295 (N_23295,N_20578,N_20807);
nand U23296 (N_23296,N_19703,N_19882);
xnor U23297 (N_23297,N_20518,N_19986);
xnor U23298 (N_23298,N_20917,N_19108);
nor U23299 (N_23299,N_19257,N_19545);
nor U23300 (N_23300,N_18166,N_20050);
xnor U23301 (N_23301,N_18097,N_20956);
and U23302 (N_23302,N_20394,N_20305);
xnor U23303 (N_23303,N_19454,N_18893);
and U23304 (N_23304,N_19983,N_18560);
or U23305 (N_23305,N_20964,N_19209);
or U23306 (N_23306,N_20221,N_20869);
xor U23307 (N_23307,N_19457,N_19088);
nor U23308 (N_23308,N_19107,N_19836);
and U23309 (N_23309,N_19900,N_18386);
nand U23310 (N_23310,N_19797,N_19923);
xnor U23311 (N_23311,N_20459,N_19750);
nor U23312 (N_23312,N_19654,N_20103);
nor U23313 (N_23313,N_19226,N_18166);
nor U23314 (N_23314,N_20146,N_19111);
nand U23315 (N_23315,N_18067,N_18353);
nand U23316 (N_23316,N_18594,N_18738);
nand U23317 (N_23317,N_18850,N_19623);
or U23318 (N_23318,N_19474,N_18391);
or U23319 (N_23319,N_20522,N_20667);
nor U23320 (N_23320,N_19597,N_19516);
xnor U23321 (N_23321,N_20647,N_18774);
nand U23322 (N_23322,N_19833,N_20544);
xor U23323 (N_23323,N_18925,N_20005);
nor U23324 (N_23324,N_20710,N_19302);
nand U23325 (N_23325,N_18075,N_20478);
and U23326 (N_23326,N_20423,N_18597);
xor U23327 (N_23327,N_20345,N_18864);
nand U23328 (N_23328,N_18148,N_20629);
nand U23329 (N_23329,N_20626,N_19570);
or U23330 (N_23330,N_19111,N_18861);
or U23331 (N_23331,N_18520,N_20374);
nand U23332 (N_23332,N_18687,N_19021);
nor U23333 (N_23333,N_20589,N_19093);
nor U23334 (N_23334,N_19805,N_19904);
and U23335 (N_23335,N_20170,N_20837);
nand U23336 (N_23336,N_19751,N_20583);
and U23337 (N_23337,N_18969,N_20029);
nor U23338 (N_23338,N_20513,N_20277);
nand U23339 (N_23339,N_19176,N_19715);
and U23340 (N_23340,N_18625,N_19695);
or U23341 (N_23341,N_20514,N_18895);
nor U23342 (N_23342,N_19064,N_20937);
nor U23343 (N_23343,N_18587,N_18632);
and U23344 (N_23344,N_18096,N_19366);
xnor U23345 (N_23345,N_18912,N_19124);
nand U23346 (N_23346,N_20437,N_19881);
nand U23347 (N_23347,N_20478,N_20779);
or U23348 (N_23348,N_18187,N_19536);
xnor U23349 (N_23349,N_18365,N_18481);
nand U23350 (N_23350,N_20198,N_20606);
nand U23351 (N_23351,N_20977,N_18338);
nor U23352 (N_23352,N_18916,N_20947);
xnor U23353 (N_23353,N_18437,N_19504);
xor U23354 (N_23354,N_18457,N_19673);
xnor U23355 (N_23355,N_18401,N_19626);
nand U23356 (N_23356,N_18177,N_18137);
nor U23357 (N_23357,N_19616,N_18235);
and U23358 (N_23358,N_19368,N_19887);
and U23359 (N_23359,N_20570,N_18755);
xor U23360 (N_23360,N_18705,N_20882);
nor U23361 (N_23361,N_18080,N_19539);
xnor U23362 (N_23362,N_19091,N_20758);
or U23363 (N_23363,N_19786,N_19991);
xor U23364 (N_23364,N_20427,N_18414);
and U23365 (N_23365,N_19653,N_18929);
nor U23366 (N_23366,N_19339,N_19269);
or U23367 (N_23367,N_18596,N_18316);
nand U23368 (N_23368,N_18142,N_20527);
and U23369 (N_23369,N_20837,N_18991);
xnor U23370 (N_23370,N_19494,N_19483);
or U23371 (N_23371,N_20261,N_19981);
nand U23372 (N_23372,N_20362,N_18153);
xnor U23373 (N_23373,N_20111,N_20106);
nor U23374 (N_23374,N_18934,N_20058);
nand U23375 (N_23375,N_20130,N_19647);
nor U23376 (N_23376,N_18911,N_18608);
nor U23377 (N_23377,N_18681,N_20653);
and U23378 (N_23378,N_19452,N_20179);
and U23379 (N_23379,N_20551,N_18178);
and U23380 (N_23380,N_19856,N_18397);
nand U23381 (N_23381,N_18753,N_19319);
or U23382 (N_23382,N_20738,N_18657);
nor U23383 (N_23383,N_18842,N_18016);
nand U23384 (N_23384,N_18942,N_20927);
nand U23385 (N_23385,N_20965,N_18868);
nor U23386 (N_23386,N_20500,N_20529);
and U23387 (N_23387,N_20117,N_19598);
and U23388 (N_23388,N_20842,N_20568);
nand U23389 (N_23389,N_20259,N_19527);
nand U23390 (N_23390,N_18146,N_18965);
and U23391 (N_23391,N_19941,N_19088);
nand U23392 (N_23392,N_19980,N_18879);
nor U23393 (N_23393,N_19732,N_18092);
nand U23394 (N_23394,N_20276,N_19234);
nor U23395 (N_23395,N_20016,N_20301);
or U23396 (N_23396,N_18612,N_20875);
xnor U23397 (N_23397,N_20903,N_20779);
or U23398 (N_23398,N_19398,N_20956);
and U23399 (N_23399,N_20597,N_19409);
or U23400 (N_23400,N_20226,N_18133);
and U23401 (N_23401,N_19458,N_19270);
xnor U23402 (N_23402,N_20864,N_18218);
or U23403 (N_23403,N_20728,N_19159);
and U23404 (N_23404,N_20440,N_18587);
nor U23405 (N_23405,N_20191,N_19667);
nor U23406 (N_23406,N_18168,N_20515);
nand U23407 (N_23407,N_19703,N_20342);
xor U23408 (N_23408,N_18921,N_19683);
or U23409 (N_23409,N_18189,N_20289);
nor U23410 (N_23410,N_20272,N_18241);
and U23411 (N_23411,N_18061,N_20782);
or U23412 (N_23412,N_18336,N_19938);
or U23413 (N_23413,N_18780,N_20795);
xor U23414 (N_23414,N_19765,N_19739);
nand U23415 (N_23415,N_20870,N_18905);
nor U23416 (N_23416,N_19247,N_18215);
nor U23417 (N_23417,N_20128,N_20927);
nand U23418 (N_23418,N_19315,N_20143);
nor U23419 (N_23419,N_18855,N_18752);
xor U23420 (N_23420,N_20592,N_20875);
xnor U23421 (N_23421,N_19089,N_18559);
or U23422 (N_23422,N_18260,N_19012);
nand U23423 (N_23423,N_19676,N_19859);
xnor U23424 (N_23424,N_20967,N_20911);
and U23425 (N_23425,N_18081,N_19371);
nor U23426 (N_23426,N_20485,N_20295);
nor U23427 (N_23427,N_18199,N_18669);
nor U23428 (N_23428,N_18223,N_20654);
or U23429 (N_23429,N_20193,N_18509);
xor U23430 (N_23430,N_19248,N_18642);
xnor U23431 (N_23431,N_19029,N_19459);
or U23432 (N_23432,N_18838,N_18898);
or U23433 (N_23433,N_19788,N_19777);
nor U23434 (N_23434,N_18838,N_19414);
nor U23435 (N_23435,N_20098,N_19006);
nor U23436 (N_23436,N_18305,N_18324);
nor U23437 (N_23437,N_20999,N_18725);
nor U23438 (N_23438,N_20272,N_18931);
or U23439 (N_23439,N_19622,N_19075);
nor U23440 (N_23440,N_18156,N_18397);
nor U23441 (N_23441,N_20525,N_20730);
or U23442 (N_23442,N_19319,N_18674);
nand U23443 (N_23443,N_20261,N_18287);
nand U23444 (N_23444,N_19009,N_20927);
nand U23445 (N_23445,N_20529,N_18458);
or U23446 (N_23446,N_19029,N_18079);
and U23447 (N_23447,N_18023,N_20098);
nand U23448 (N_23448,N_19257,N_19560);
nor U23449 (N_23449,N_20872,N_20808);
nand U23450 (N_23450,N_19165,N_19279);
xnor U23451 (N_23451,N_19364,N_18846);
nand U23452 (N_23452,N_19098,N_19236);
and U23453 (N_23453,N_19966,N_19991);
nor U23454 (N_23454,N_18382,N_19656);
xor U23455 (N_23455,N_19586,N_19277);
nand U23456 (N_23456,N_20893,N_19518);
and U23457 (N_23457,N_20472,N_19423);
nand U23458 (N_23458,N_20840,N_19531);
xor U23459 (N_23459,N_20499,N_19480);
nor U23460 (N_23460,N_18436,N_20749);
and U23461 (N_23461,N_20107,N_19590);
nand U23462 (N_23462,N_19025,N_20937);
nand U23463 (N_23463,N_18099,N_20035);
xnor U23464 (N_23464,N_18328,N_19061);
nand U23465 (N_23465,N_19041,N_18980);
or U23466 (N_23466,N_20196,N_20601);
and U23467 (N_23467,N_20081,N_18371);
or U23468 (N_23468,N_19478,N_20808);
or U23469 (N_23469,N_19621,N_19681);
xor U23470 (N_23470,N_20039,N_19606);
nor U23471 (N_23471,N_20114,N_19099);
nand U23472 (N_23472,N_20761,N_20665);
nand U23473 (N_23473,N_20700,N_19011);
nor U23474 (N_23474,N_18207,N_20823);
xor U23475 (N_23475,N_19495,N_18902);
nor U23476 (N_23476,N_18333,N_20976);
xor U23477 (N_23477,N_19501,N_18670);
nor U23478 (N_23478,N_18330,N_18116);
nand U23479 (N_23479,N_19890,N_20628);
nor U23480 (N_23480,N_18852,N_20469);
xnor U23481 (N_23481,N_18158,N_19807);
nand U23482 (N_23482,N_18493,N_20201);
xnor U23483 (N_23483,N_20932,N_20717);
and U23484 (N_23484,N_19113,N_20854);
nor U23485 (N_23485,N_18309,N_18779);
or U23486 (N_23486,N_19080,N_18420);
or U23487 (N_23487,N_20344,N_18591);
or U23488 (N_23488,N_19973,N_20541);
nor U23489 (N_23489,N_20927,N_20114);
or U23490 (N_23490,N_19975,N_20267);
nor U23491 (N_23491,N_20363,N_19762);
and U23492 (N_23492,N_18032,N_20883);
nor U23493 (N_23493,N_18509,N_18404);
nand U23494 (N_23494,N_18555,N_18085);
nor U23495 (N_23495,N_20239,N_19568);
nand U23496 (N_23496,N_18723,N_19999);
or U23497 (N_23497,N_20645,N_20963);
xnor U23498 (N_23498,N_19517,N_20794);
xor U23499 (N_23499,N_20694,N_18983);
xor U23500 (N_23500,N_18183,N_18869);
nor U23501 (N_23501,N_19119,N_18716);
nand U23502 (N_23502,N_19176,N_20749);
nor U23503 (N_23503,N_20215,N_18610);
and U23504 (N_23504,N_18773,N_19436);
or U23505 (N_23505,N_18273,N_18406);
nor U23506 (N_23506,N_20323,N_18152);
nand U23507 (N_23507,N_19717,N_19157);
nor U23508 (N_23508,N_18521,N_20401);
and U23509 (N_23509,N_19793,N_19354);
nor U23510 (N_23510,N_18555,N_20356);
xnor U23511 (N_23511,N_19843,N_19274);
or U23512 (N_23512,N_18440,N_20335);
and U23513 (N_23513,N_20423,N_20583);
xnor U23514 (N_23514,N_18224,N_20799);
nor U23515 (N_23515,N_20710,N_18983);
and U23516 (N_23516,N_19080,N_19807);
and U23517 (N_23517,N_19996,N_20429);
and U23518 (N_23518,N_19491,N_20442);
and U23519 (N_23519,N_20318,N_20742);
nor U23520 (N_23520,N_18445,N_20351);
nand U23521 (N_23521,N_20187,N_18100);
xor U23522 (N_23522,N_19899,N_18076);
or U23523 (N_23523,N_20170,N_19723);
or U23524 (N_23524,N_20991,N_19777);
nand U23525 (N_23525,N_19798,N_20779);
or U23526 (N_23526,N_18061,N_19238);
and U23527 (N_23527,N_18087,N_20080);
nand U23528 (N_23528,N_18910,N_18408);
xor U23529 (N_23529,N_20134,N_19680);
or U23530 (N_23530,N_19029,N_19071);
or U23531 (N_23531,N_18784,N_18976);
nor U23532 (N_23532,N_18645,N_18899);
nor U23533 (N_23533,N_20333,N_20437);
or U23534 (N_23534,N_19322,N_18005);
nor U23535 (N_23535,N_20437,N_18725);
or U23536 (N_23536,N_19744,N_19271);
xnor U23537 (N_23537,N_20966,N_19828);
nor U23538 (N_23538,N_19773,N_20144);
or U23539 (N_23539,N_20184,N_18349);
nor U23540 (N_23540,N_19380,N_19737);
and U23541 (N_23541,N_18832,N_19370);
nand U23542 (N_23542,N_19928,N_18993);
nor U23543 (N_23543,N_19784,N_19127);
or U23544 (N_23544,N_18186,N_18669);
and U23545 (N_23545,N_20686,N_18168);
and U23546 (N_23546,N_20334,N_18556);
xnor U23547 (N_23547,N_20042,N_18599);
and U23548 (N_23548,N_20082,N_19270);
or U23549 (N_23549,N_18767,N_19906);
xnor U23550 (N_23550,N_19124,N_20794);
or U23551 (N_23551,N_19577,N_18336);
nand U23552 (N_23552,N_19028,N_18168);
nand U23553 (N_23553,N_18113,N_18791);
nor U23554 (N_23554,N_19873,N_18820);
and U23555 (N_23555,N_20531,N_20012);
or U23556 (N_23556,N_19315,N_20476);
nor U23557 (N_23557,N_18109,N_19953);
nand U23558 (N_23558,N_18990,N_18756);
or U23559 (N_23559,N_20740,N_18217);
xor U23560 (N_23560,N_19106,N_19478);
xnor U23561 (N_23561,N_19255,N_20421);
and U23562 (N_23562,N_19244,N_19157);
and U23563 (N_23563,N_19576,N_19669);
nand U23564 (N_23564,N_19781,N_20291);
nand U23565 (N_23565,N_18632,N_18433);
nand U23566 (N_23566,N_19389,N_18083);
nor U23567 (N_23567,N_20784,N_20228);
or U23568 (N_23568,N_19710,N_19626);
xor U23569 (N_23569,N_20742,N_18973);
nand U23570 (N_23570,N_19071,N_18218);
and U23571 (N_23571,N_20618,N_19208);
nand U23572 (N_23572,N_18855,N_18417);
nor U23573 (N_23573,N_20262,N_18670);
nand U23574 (N_23574,N_19369,N_20758);
nand U23575 (N_23575,N_19012,N_19417);
nor U23576 (N_23576,N_20935,N_18904);
nand U23577 (N_23577,N_18796,N_18770);
nor U23578 (N_23578,N_18104,N_18120);
nand U23579 (N_23579,N_20646,N_18701);
nand U23580 (N_23580,N_20996,N_18568);
xor U23581 (N_23581,N_18583,N_20947);
and U23582 (N_23582,N_18343,N_20607);
nor U23583 (N_23583,N_19650,N_19384);
nor U23584 (N_23584,N_18166,N_20993);
or U23585 (N_23585,N_18166,N_19872);
nand U23586 (N_23586,N_20449,N_18575);
nand U23587 (N_23587,N_19225,N_19977);
and U23588 (N_23588,N_19921,N_19400);
xor U23589 (N_23589,N_18171,N_19748);
nor U23590 (N_23590,N_20576,N_19393);
nor U23591 (N_23591,N_18093,N_20143);
nor U23592 (N_23592,N_18251,N_18269);
nand U23593 (N_23593,N_19123,N_18531);
nand U23594 (N_23594,N_18145,N_18324);
xor U23595 (N_23595,N_18755,N_18896);
xor U23596 (N_23596,N_20280,N_19690);
nor U23597 (N_23597,N_18999,N_20828);
or U23598 (N_23598,N_18606,N_20468);
and U23599 (N_23599,N_19693,N_20324);
nand U23600 (N_23600,N_19859,N_20426);
and U23601 (N_23601,N_18773,N_20715);
nand U23602 (N_23602,N_19197,N_18759);
nand U23603 (N_23603,N_20982,N_18230);
and U23604 (N_23604,N_18614,N_19593);
nand U23605 (N_23605,N_18452,N_19878);
nand U23606 (N_23606,N_19916,N_19715);
nand U23607 (N_23607,N_18034,N_20918);
nor U23608 (N_23608,N_20521,N_18395);
xor U23609 (N_23609,N_19269,N_20303);
nand U23610 (N_23610,N_18894,N_19796);
nor U23611 (N_23611,N_19432,N_19983);
nand U23612 (N_23612,N_18303,N_19623);
and U23613 (N_23613,N_18420,N_18275);
and U23614 (N_23614,N_20166,N_18440);
nand U23615 (N_23615,N_20485,N_19209);
or U23616 (N_23616,N_19691,N_20654);
nor U23617 (N_23617,N_20896,N_20027);
and U23618 (N_23618,N_18251,N_18291);
nor U23619 (N_23619,N_20964,N_18745);
and U23620 (N_23620,N_20297,N_19469);
xnor U23621 (N_23621,N_19036,N_20903);
and U23622 (N_23622,N_20154,N_20512);
nand U23623 (N_23623,N_18852,N_18893);
or U23624 (N_23624,N_18316,N_19686);
and U23625 (N_23625,N_18907,N_19182);
nor U23626 (N_23626,N_19650,N_19994);
or U23627 (N_23627,N_18528,N_20093);
or U23628 (N_23628,N_20809,N_18391);
and U23629 (N_23629,N_18190,N_20829);
or U23630 (N_23630,N_20681,N_20107);
and U23631 (N_23631,N_20546,N_19403);
xnor U23632 (N_23632,N_19027,N_18319);
xnor U23633 (N_23633,N_20972,N_20351);
xor U23634 (N_23634,N_19635,N_20505);
xor U23635 (N_23635,N_19851,N_20240);
or U23636 (N_23636,N_19091,N_19239);
nand U23637 (N_23637,N_19712,N_20843);
xnor U23638 (N_23638,N_18251,N_19484);
nor U23639 (N_23639,N_18836,N_19744);
nor U23640 (N_23640,N_20156,N_19251);
xor U23641 (N_23641,N_19109,N_19583);
and U23642 (N_23642,N_20498,N_18942);
nand U23643 (N_23643,N_18514,N_20229);
xor U23644 (N_23644,N_20941,N_18545);
and U23645 (N_23645,N_19074,N_20033);
nand U23646 (N_23646,N_20635,N_18512);
and U23647 (N_23647,N_20305,N_20472);
and U23648 (N_23648,N_19032,N_18618);
xnor U23649 (N_23649,N_20625,N_18218);
nand U23650 (N_23650,N_20280,N_18639);
or U23651 (N_23651,N_20942,N_19279);
nand U23652 (N_23652,N_20397,N_19571);
xor U23653 (N_23653,N_19711,N_20019);
nand U23654 (N_23654,N_19877,N_18122);
xnor U23655 (N_23655,N_18177,N_19013);
xnor U23656 (N_23656,N_18866,N_18961);
xor U23657 (N_23657,N_18009,N_19165);
or U23658 (N_23658,N_19172,N_18147);
xor U23659 (N_23659,N_19793,N_20156);
and U23660 (N_23660,N_18400,N_20267);
nand U23661 (N_23661,N_20772,N_18970);
xnor U23662 (N_23662,N_19452,N_18069);
xor U23663 (N_23663,N_18262,N_19120);
nor U23664 (N_23664,N_19091,N_18827);
and U23665 (N_23665,N_19042,N_18745);
xnor U23666 (N_23666,N_20312,N_18301);
and U23667 (N_23667,N_18760,N_19606);
and U23668 (N_23668,N_18932,N_19604);
or U23669 (N_23669,N_19810,N_20667);
xor U23670 (N_23670,N_19284,N_20358);
or U23671 (N_23671,N_20828,N_19298);
or U23672 (N_23672,N_20511,N_18415);
nor U23673 (N_23673,N_18397,N_19679);
and U23674 (N_23674,N_20768,N_18953);
xor U23675 (N_23675,N_18064,N_19540);
or U23676 (N_23676,N_20924,N_18929);
and U23677 (N_23677,N_19506,N_19210);
or U23678 (N_23678,N_20581,N_19681);
nand U23679 (N_23679,N_18855,N_20646);
nor U23680 (N_23680,N_18014,N_18358);
nand U23681 (N_23681,N_19987,N_20532);
xnor U23682 (N_23682,N_18113,N_19084);
or U23683 (N_23683,N_18309,N_18125);
and U23684 (N_23684,N_20701,N_18888);
nor U23685 (N_23685,N_18928,N_20818);
and U23686 (N_23686,N_19504,N_18323);
and U23687 (N_23687,N_20657,N_20637);
nand U23688 (N_23688,N_20419,N_20303);
nor U23689 (N_23689,N_19677,N_18477);
nand U23690 (N_23690,N_20940,N_20545);
and U23691 (N_23691,N_19643,N_18373);
nor U23692 (N_23692,N_18375,N_18469);
nor U23693 (N_23693,N_19159,N_19964);
nor U23694 (N_23694,N_20355,N_20753);
xor U23695 (N_23695,N_20125,N_18204);
or U23696 (N_23696,N_19635,N_18486);
or U23697 (N_23697,N_20743,N_19879);
nand U23698 (N_23698,N_18038,N_19560);
or U23699 (N_23699,N_20615,N_19609);
and U23700 (N_23700,N_19604,N_20682);
nand U23701 (N_23701,N_19194,N_18912);
or U23702 (N_23702,N_19035,N_18349);
or U23703 (N_23703,N_18356,N_19089);
nand U23704 (N_23704,N_20894,N_19041);
xnor U23705 (N_23705,N_18993,N_18573);
and U23706 (N_23706,N_20170,N_20500);
xor U23707 (N_23707,N_19269,N_20026);
xnor U23708 (N_23708,N_18373,N_18739);
xor U23709 (N_23709,N_18926,N_18426);
or U23710 (N_23710,N_18873,N_18428);
nand U23711 (N_23711,N_20312,N_19281);
xnor U23712 (N_23712,N_20061,N_19810);
nand U23713 (N_23713,N_20428,N_20580);
nor U23714 (N_23714,N_19172,N_20753);
nor U23715 (N_23715,N_20343,N_18575);
and U23716 (N_23716,N_20204,N_19668);
and U23717 (N_23717,N_18385,N_19924);
or U23718 (N_23718,N_20890,N_18179);
or U23719 (N_23719,N_20250,N_19980);
nand U23720 (N_23720,N_19190,N_20863);
nand U23721 (N_23721,N_18930,N_20169);
xnor U23722 (N_23722,N_20234,N_19428);
xor U23723 (N_23723,N_19542,N_20419);
nand U23724 (N_23724,N_19863,N_18868);
nand U23725 (N_23725,N_19612,N_20299);
and U23726 (N_23726,N_19408,N_18305);
or U23727 (N_23727,N_19329,N_19855);
xor U23728 (N_23728,N_19870,N_18827);
nand U23729 (N_23729,N_18492,N_20853);
or U23730 (N_23730,N_18976,N_20747);
nor U23731 (N_23731,N_19072,N_20602);
nor U23732 (N_23732,N_20640,N_19887);
and U23733 (N_23733,N_19269,N_19971);
nor U23734 (N_23734,N_18606,N_18840);
nand U23735 (N_23735,N_18859,N_18823);
xnor U23736 (N_23736,N_19711,N_18313);
or U23737 (N_23737,N_18861,N_20116);
and U23738 (N_23738,N_19828,N_18766);
or U23739 (N_23739,N_19046,N_18801);
nor U23740 (N_23740,N_19307,N_20192);
nor U23741 (N_23741,N_19245,N_19370);
and U23742 (N_23742,N_19560,N_20784);
nand U23743 (N_23743,N_19241,N_18899);
nand U23744 (N_23744,N_18011,N_19361);
and U23745 (N_23745,N_20237,N_19304);
and U23746 (N_23746,N_18656,N_19235);
nor U23747 (N_23747,N_19000,N_20488);
nand U23748 (N_23748,N_19900,N_19990);
and U23749 (N_23749,N_20213,N_19388);
or U23750 (N_23750,N_18620,N_20858);
xor U23751 (N_23751,N_20272,N_19698);
nor U23752 (N_23752,N_20574,N_18743);
and U23753 (N_23753,N_19431,N_18129);
nor U23754 (N_23754,N_20655,N_19563);
or U23755 (N_23755,N_18456,N_19650);
and U23756 (N_23756,N_19006,N_18410);
xnor U23757 (N_23757,N_18690,N_20691);
nor U23758 (N_23758,N_20063,N_18628);
xor U23759 (N_23759,N_20948,N_20864);
xnor U23760 (N_23760,N_20230,N_20338);
xnor U23761 (N_23761,N_19818,N_18478);
nor U23762 (N_23762,N_19799,N_20765);
nor U23763 (N_23763,N_20176,N_18794);
or U23764 (N_23764,N_19974,N_18388);
or U23765 (N_23765,N_19497,N_20744);
xnor U23766 (N_23766,N_19543,N_19003);
nand U23767 (N_23767,N_20280,N_20971);
nand U23768 (N_23768,N_19046,N_18816);
or U23769 (N_23769,N_18278,N_19129);
and U23770 (N_23770,N_19468,N_18876);
or U23771 (N_23771,N_19913,N_19095);
nand U23772 (N_23772,N_18848,N_20091);
or U23773 (N_23773,N_20010,N_20575);
xnor U23774 (N_23774,N_18538,N_18761);
xor U23775 (N_23775,N_18092,N_19067);
nand U23776 (N_23776,N_18286,N_18610);
nand U23777 (N_23777,N_19945,N_18436);
or U23778 (N_23778,N_19414,N_20395);
and U23779 (N_23779,N_18105,N_18640);
or U23780 (N_23780,N_19618,N_18192);
nor U23781 (N_23781,N_19369,N_19111);
nor U23782 (N_23782,N_18938,N_20447);
nand U23783 (N_23783,N_19632,N_19298);
nor U23784 (N_23784,N_18309,N_19828);
and U23785 (N_23785,N_20224,N_20906);
nand U23786 (N_23786,N_19576,N_19120);
nand U23787 (N_23787,N_19670,N_18729);
xnor U23788 (N_23788,N_18878,N_18368);
xor U23789 (N_23789,N_19896,N_18972);
xnor U23790 (N_23790,N_18224,N_19827);
nor U23791 (N_23791,N_20829,N_20601);
or U23792 (N_23792,N_18472,N_20376);
nand U23793 (N_23793,N_18932,N_19715);
nand U23794 (N_23794,N_19798,N_18095);
or U23795 (N_23795,N_18916,N_20760);
or U23796 (N_23796,N_20221,N_20972);
and U23797 (N_23797,N_18116,N_19695);
and U23798 (N_23798,N_19060,N_18079);
or U23799 (N_23799,N_19744,N_18924);
nand U23800 (N_23800,N_19521,N_18715);
nor U23801 (N_23801,N_18831,N_19265);
or U23802 (N_23802,N_18792,N_18468);
and U23803 (N_23803,N_20546,N_19636);
nor U23804 (N_23804,N_18552,N_19123);
nor U23805 (N_23805,N_18593,N_19908);
nand U23806 (N_23806,N_18367,N_20992);
and U23807 (N_23807,N_18584,N_18045);
nor U23808 (N_23808,N_18351,N_18785);
nand U23809 (N_23809,N_19399,N_18106);
nor U23810 (N_23810,N_18971,N_20657);
xnor U23811 (N_23811,N_20192,N_19902);
xnor U23812 (N_23812,N_19249,N_20557);
nor U23813 (N_23813,N_19509,N_18007);
and U23814 (N_23814,N_20425,N_20770);
or U23815 (N_23815,N_19254,N_19188);
or U23816 (N_23816,N_18789,N_19016);
or U23817 (N_23817,N_19817,N_20127);
nand U23818 (N_23818,N_19796,N_20388);
or U23819 (N_23819,N_19435,N_18324);
or U23820 (N_23820,N_18419,N_20560);
and U23821 (N_23821,N_19318,N_19956);
and U23822 (N_23822,N_18226,N_19849);
nand U23823 (N_23823,N_20095,N_19412);
xnor U23824 (N_23824,N_20760,N_20971);
nand U23825 (N_23825,N_18610,N_18935);
or U23826 (N_23826,N_18114,N_20338);
xor U23827 (N_23827,N_19230,N_19758);
nand U23828 (N_23828,N_20014,N_19436);
and U23829 (N_23829,N_20625,N_19048);
xor U23830 (N_23830,N_20348,N_18351);
and U23831 (N_23831,N_18082,N_19913);
or U23832 (N_23832,N_18804,N_20797);
nand U23833 (N_23833,N_19422,N_18281);
xnor U23834 (N_23834,N_19614,N_19488);
or U23835 (N_23835,N_18736,N_19596);
and U23836 (N_23836,N_20559,N_19413);
nor U23837 (N_23837,N_18418,N_20331);
xor U23838 (N_23838,N_20879,N_20179);
xor U23839 (N_23839,N_18660,N_19649);
or U23840 (N_23840,N_18934,N_20923);
or U23841 (N_23841,N_18479,N_20907);
nand U23842 (N_23842,N_19673,N_18705);
nand U23843 (N_23843,N_20870,N_20211);
and U23844 (N_23844,N_20038,N_20365);
nor U23845 (N_23845,N_18845,N_18116);
nor U23846 (N_23846,N_18138,N_18715);
xor U23847 (N_23847,N_20699,N_18069);
or U23848 (N_23848,N_19941,N_18366);
and U23849 (N_23849,N_18784,N_18931);
nor U23850 (N_23850,N_19394,N_18938);
xnor U23851 (N_23851,N_19311,N_18189);
or U23852 (N_23852,N_18655,N_20483);
xnor U23853 (N_23853,N_18626,N_18922);
or U23854 (N_23854,N_18004,N_18357);
nor U23855 (N_23855,N_18496,N_20246);
and U23856 (N_23856,N_20210,N_20104);
and U23857 (N_23857,N_18226,N_19421);
or U23858 (N_23858,N_18661,N_19914);
xnor U23859 (N_23859,N_20405,N_18200);
nand U23860 (N_23860,N_20115,N_19277);
or U23861 (N_23861,N_19917,N_18875);
nor U23862 (N_23862,N_18887,N_18036);
or U23863 (N_23863,N_20278,N_19842);
or U23864 (N_23864,N_20663,N_20179);
xor U23865 (N_23865,N_20643,N_19524);
nor U23866 (N_23866,N_20627,N_19797);
nand U23867 (N_23867,N_18141,N_18635);
nand U23868 (N_23868,N_20154,N_19666);
nor U23869 (N_23869,N_20741,N_20765);
xor U23870 (N_23870,N_18114,N_19331);
and U23871 (N_23871,N_19769,N_20446);
or U23872 (N_23872,N_19028,N_20707);
nor U23873 (N_23873,N_20450,N_20559);
or U23874 (N_23874,N_20681,N_18665);
nor U23875 (N_23875,N_19193,N_20240);
xor U23876 (N_23876,N_19717,N_19665);
nand U23877 (N_23877,N_18104,N_19013);
xnor U23878 (N_23878,N_19868,N_19687);
xor U23879 (N_23879,N_19837,N_20968);
and U23880 (N_23880,N_20899,N_18280);
or U23881 (N_23881,N_18974,N_20245);
xnor U23882 (N_23882,N_18789,N_20265);
xnor U23883 (N_23883,N_20117,N_18730);
xor U23884 (N_23884,N_19440,N_19812);
nor U23885 (N_23885,N_19237,N_19198);
nand U23886 (N_23886,N_20397,N_20658);
or U23887 (N_23887,N_18712,N_19180);
xor U23888 (N_23888,N_19425,N_18470);
xor U23889 (N_23889,N_19535,N_19621);
xor U23890 (N_23890,N_18553,N_19780);
nand U23891 (N_23891,N_20871,N_19421);
or U23892 (N_23892,N_20707,N_20508);
nor U23893 (N_23893,N_18450,N_20588);
or U23894 (N_23894,N_19044,N_19157);
nand U23895 (N_23895,N_18546,N_18389);
nor U23896 (N_23896,N_20217,N_20158);
or U23897 (N_23897,N_20030,N_19783);
and U23898 (N_23898,N_18228,N_18696);
and U23899 (N_23899,N_18086,N_18078);
nand U23900 (N_23900,N_18391,N_19144);
nand U23901 (N_23901,N_18277,N_20308);
and U23902 (N_23902,N_18345,N_18369);
or U23903 (N_23903,N_19820,N_20097);
and U23904 (N_23904,N_18022,N_20184);
xor U23905 (N_23905,N_18530,N_20004);
nand U23906 (N_23906,N_18837,N_18628);
or U23907 (N_23907,N_20063,N_20155);
or U23908 (N_23908,N_20176,N_19363);
and U23909 (N_23909,N_20306,N_18664);
xnor U23910 (N_23910,N_20138,N_19752);
or U23911 (N_23911,N_18941,N_19270);
nand U23912 (N_23912,N_18259,N_20008);
nand U23913 (N_23913,N_20686,N_18415);
nor U23914 (N_23914,N_18261,N_18107);
or U23915 (N_23915,N_18841,N_20669);
nand U23916 (N_23916,N_18682,N_20692);
nor U23917 (N_23917,N_20188,N_19912);
xor U23918 (N_23918,N_18024,N_20768);
and U23919 (N_23919,N_20666,N_20186);
nand U23920 (N_23920,N_20511,N_18049);
and U23921 (N_23921,N_20654,N_18545);
or U23922 (N_23922,N_19646,N_20157);
nand U23923 (N_23923,N_18859,N_19201);
and U23924 (N_23924,N_20989,N_20736);
nor U23925 (N_23925,N_20770,N_20547);
xnor U23926 (N_23926,N_18426,N_20222);
nor U23927 (N_23927,N_18434,N_18055);
xnor U23928 (N_23928,N_19617,N_18363);
or U23929 (N_23929,N_18229,N_18939);
nor U23930 (N_23930,N_20376,N_18709);
xnor U23931 (N_23931,N_18702,N_18623);
nand U23932 (N_23932,N_20505,N_19902);
or U23933 (N_23933,N_19829,N_20332);
or U23934 (N_23934,N_20669,N_18534);
and U23935 (N_23935,N_19760,N_19977);
and U23936 (N_23936,N_18083,N_18422);
or U23937 (N_23937,N_19473,N_19040);
nor U23938 (N_23938,N_18381,N_18130);
and U23939 (N_23939,N_20612,N_18837);
and U23940 (N_23940,N_20767,N_18156);
nand U23941 (N_23941,N_19218,N_18666);
and U23942 (N_23942,N_18305,N_20925);
nor U23943 (N_23943,N_20661,N_19521);
xnor U23944 (N_23944,N_19746,N_19025);
nand U23945 (N_23945,N_19028,N_19232);
xor U23946 (N_23946,N_19272,N_19316);
nand U23947 (N_23947,N_18526,N_19360);
and U23948 (N_23948,N_20171,N_19508);
xor U23949 (N_23949,N_18162,N_18740);
and U23950 (N_23950,N_18349,N_18691);
nand U23951 (N_23951,N_18415,N_19877);
and U23952 (N_23952,N_19481,N_19834);
nor U23953 (N_23953,N_19790,N_20635);
and U23954 (N_23954,N_18176,N_20101);
xor U23955 (N_23955,N_19628,N_18436);
and U23956 (N_23956,N_19477,N_20066);
nand U23957 (N_23957,N_19301,N_18848);
nand U23958 (N_23958,N_20775,N_19129);
and U23959 (N_23959,N_20331,N_19703);
nor U23960 (N_23960,N_20490,N_18634);
nand U23961 (N_23961,N_20145,N_18935);
nand U23962 (N_23962,N_18106,N_18758);
or U23963 (N_23963,N_19704,N_20868);
or U23964 (N_23964,N_19549,N_19688);
or U23965 (N_23965,N_19807,N_18468);
nor U23966 (N_23966,N_19360,N_20142);
nand U23967 (N_23967,N_20223,N_19273);
nand U23968 (N_23968,N_18366,N_20689);
and U23969 (N_23969,N_18047,N_20647);
nor U23970 (N_23970,N_19428,N_20169);
nor U23971 (N_23971,N_18893,N_20550);
and U23972 (N_23972,N_19507,N_20727);
or U23973 (N_23973,N_19336,N_19872);
nand U23974 (N_23974,N_19046,N_20633);
nand U23975 (N_23975,N_18278,N_19772);
nor U23976 (N_23976,N_18024,N_20076);
and U23977 (N_23977,N_18673,N_20675);
and U23978 (N_23978,N_20003,N_19172);
and U23979 (N_23979,N_19672,N_20112);
or U23980 (N_23980,N_20450,N_19419);
or U23981 (N_23981,N_19075,N_18486);
and U23982 (N_23982,N_20126,N_19400);
and U23983 (N_23983,N_19005,N_19705);
or U23984 (N_23984,N_18862,N_19648);
or U23985 (N_23985,N_18236,N_20566);
nand U23986 (N_23986,N_18632,N_18061);
or U23987 (N_23987,N_19341,N_18020);
nand U23988 (N_23988,N_20369,N_20662);
and U23989 (N_23989,N_18730,N_19815);
xnor U23990 (N_23990,N_18247,N_19528);
nand U23991 (N_23991,N_19036,N_19874);
or U23992 (N_23992,N_20020,N_18442);
nor U23993 (N_23993,N_20160,N_18100);
or U23994 (N_23994,N_20767,N_19649);
nor U23995 (N_23995,N_18121,N_19802);
nand U23996 (N_23996,N_18232,N_20883);
or U23997 (N_23997,N_20864,N_18772);
or U23998 (N_23998,N_20681,N_18814);
xnor U23999 (N_23999,N_18200,N_18460);
xnor U24000 (N_24000,N_22766,N_23606);
or U24001 (N_24001,N_22984,N_23519);
and U24002 (N_24002,N_21840,N_23354);
or U24003 (N_24003,N_22645,N_23236);
xor U24004 (N_24004,N_23243,N_23635);
nor U24005 (N_24005,N_21693,N_22596);
or U24006 (N_24006,N_22430,N_23316);
nand U24007 (N_24007,N_22918,N_23920);
or U24008 (N_24008,N_22529,N_21828);
and U24009 (N_24009,N_22203,N_23416);
nand U24010 (N_24010,N_23535,N_21820);
xnor U24011 (N_24011,N_23493,N_23851);
xnor U24012 (N_24012,N_22665,N_23867);
nand U24013 (N_24013,N_22157,N_21149);
nand U24014 (N_24014,N_21649,N_23835);
and U24015 (N_24015,N_23751,N_23222);
and U24016 (N_24016,N_21801,N_22934);
xor U24017 (N_24017,N_21882,N_23165);
xnor U24018 (N_24018,N_23198,N_21762);
or U24019 (N_24019,N_21119,N_22653);
xor U24020 (N_24020,N_23647,N_23177);
nor U24021 (N_24021,N_22813,N_21296);
nor U24022 (N_24022,N_21896,N_23224);
nand U24023 (N_24023,N_21277,N_23050);
and U24024 (N_24024,N_23853,N_23529);
nand U24025 (N_24025,N_22874,N_22499);
nand U24026 (N_24026,N_23710,N_23526);
and U24027 (N_24027,N_22524,N_23210);
or U24028 (N_24028,N_22117,N_23139);
nand U24029 (N_24029,N_21130,N_23722);
nor U24030 (N_24030,N_22176,N_22990);
and U24031 (N_24031,N_23207,N_23332);
and U24032 (N_24032,N_23330,N_23731);
and U24033 (N_24033,N_22457,N_21609);
xor U24034 (N_24034,N_22268,N_22843);
nor U24035 (N_24035,N_21124,N_23926);
nor U24036 (N_24036,N_21421,N_23217);
nor U24037 (N_24037,N_21646,N_23321);
and U24038 (N_24038,N_22301,N_21702);
or U24039 (N_24039,N_21629,N_21495);
or U24040 (N_24040,N_23840,N_22396);
and U24041 (N_24041,N_21053,N_21613);
nand U24042 (N_24042,N_23323,N_23600);
xnor U24043 (N_24043,N_23318,N_23547);
or U24044 (N_24044,N_23730,N_22635);
or U24045 (N_24045,N_23972,N_23464);
nand U24046 (N_24046,N_21689,N_22664);
xnor U24047 (N_24047,N_21071,N_23087);
and U24048 (N_24048,N_22633,N_22121);
nor U24049 (N_24049,N_21981,N_21926);
nand U24050 (N_24050,N_22437,N_21739);
and U24051 (N_24051,N_21110,N_21829);
nor U24052 (N_24052,N_21152,N_21144);
nand U24053 (N_24053,N_21187,N_23718);
and U24054 (N_24054,N_22274,N_21169);
nand U24055 (N_24055,N_21331,N_23447);
nor U24056 (N_24056,N_22903,N_23041);
nand U24057 (N_24057,N_23197,N_22646);
or U24058 (N_24058,N_22381,N_23513);
and U24059 (N_24059,N_21092,N_23508);
and U24060 (N_24060,N_21447,N_21979);
nand U24061 (N_24061,N_21938,N_22383);
or U24062 (N_24062,N_23775,N_23062);
or U24063 (N_24063,N_23393,N_21462);
or U24064 (N_24064,N_21579,N_22746);
nand U24065 (N_24065,N_21150,N_21474);
nand U24066 (N_24066,N_21089,N_21639);
or U24067 (N_24067,N_23051,N_21767);
or U24068 (N_24068,N_22788,N_22395);
nor U24069 (N_24069,N_21575,N_23620);
nor U24070 (N_24070,N_23875,N_23812);
or U24071 (N_24071,N_23175,N_21723);
and U24072 (N_24072,N_23172,N_21589);
nand U24073 (N_24073,N_21271,N_21472);
nor U24074 (N_24074,N_22745,N_22679);
nand U24075 (N_24075,N_22644,N_22111);
xor U24076 (N_24076,N_23530,N_22331);
xnor U24077 (N_24077,N_21791,N_22423);
and U24078 (N_24078,N_21626,N_21788);
nor U24079 (N_24079,N_21714,N_23297);
and U24080 (N_24080,N_21991,N_22300);
or U24081 (N_24081,N_21466,N_23490);
nor U24082 (N_24082,N_23040,N_23525);
or U24083 (N_24083,N_21257,N_21996);
xnor U24084 (N_24084,N_23199,N_21832);
xnor U24085 (N_24085,N_21258,N_23151);
xnor U24086 (N_24086,N_23415,N_21163);
nor U24087 (N_24087,N_23860,N_22087);
nor U24088 (N_24088,N_23260,N_23049);
or U24089 (N_24089,N_22774,N_23232);
or U24090 (N_24090,N_21814,N_21846);
nor U24091 (N_24091,N_23675,N_21232);
xnor U24092 (N_24092,N_21240,N_22211);
and U24093 (N_24093,N_22483,N_23994);
nor U24094 (N_24094,N_22888,N_23810);
or U24095 (N_24095,N_23263,N_22458);
and U24096 (N_24096,N_21743,N_22494);
and U24097 (N_24097,N_21024,N_23191);
xor U24098 (N_24098,N_23322,N_21803);
or U24099 (N_24099,N_21494,N_21334);
nor U24100 (N_24100,N_22075,N_22053);
or U24101 (N_24101,N_22208,N_22463);
or U24102 (N_24102,N_22558,N_23220);
or U24103 (N_24103,N_22915,N_22591);
nand U24104 (N_24104,N_22527,N_21279);
or U24105 (N_24105,N_23697,N_21284);
nor U24106 (N_24106,N_23690,N_21823);
nand U24107 (N_24107,N_22357,N_22961);
nor U24108 (N_24108,N_22827,N_21233);
nand U24109 (N_24109,N_22974,N_23023);
and U24110 (N_24110,N_22092,N_22019);
and U24111 (N_24111,N_23757,N_23476);
xor U24112 (N_24112,N_23708,N_23967);
xnor U24113 (N_24113,N_22674,N_23616);
or U24114 (N_24114,N_22787,N_23090);
nand U24115 (N_24115,N_23029,N_21108);
or U24116 (N_24116,N_22728,N_21622);
and U24117 (N_24117,N_21899,N_23787);
and U24118 (N_24118,N_23400,N_22384);
nand U24119 (N_24119,N_23132,N_23195);
or U24120 (N_24120,N_22126,N_21405);
nand U24121 (N_24121,N_23239,N_21865);
nor U24122 (N_24122,N_22701,N_21485);
xnor U24123 (N_24123,N_22688,N_23194);
nand U24124 (N_24124,N_23358,N_22749);
nor U24125 (N_24125,N_23178,N_22509);
and U24126 (N_24126,N_22882,N_22251);
or U24127 (N_24127,N_23923,N_22505);
and U24128 (N_24128,N_22611,N_22639);
xnor U24129 (N_24129,N_22508,N_23341);
nor U24130 (N_24130,N_22060,N_23017);
xor U24131 (N_24131,N_23497,N_22163);
xor U24132 (N_24132,N_22227,N_23912);
xor U24133 (N_24133,N_22660,N_23219);
and U24134 (N_24134,N_21912,N_22077);
nor U24135 (N_24135,N_22120,N_21434);
and U24136 (N_24136,N_23597,N_21855);
and U24137 (N_24137,N_21311,N_23861);
nor U24138 (N_24138,N_21033,N_22538);
nor U24139 (N_24139,N_22663,N_21999);
xnor U24140 (N_24140,N_23668,N_23906);
or U24141 (N_24141,N_23752,N_23968);
xor U24142 (N_24142,N_23326,N_22206);
xnor U24143 (N_24143,N_23723,N_22319);
or U24144 (N_24144,N_21709,N_21054);
nand U24145 (N_24145,N_21404,N_21994);
nor U24146 (N_24146,N_22577,N_21628);
nand U24147 (N_24147,N_21191,N_23998);
or U24148 (N_24148,N_21733,N_21562);
and U24149 (N_24149,N_21891,N_22333);
nand U24150 (N_24150,N_22860,N_23784);
and U24151 (N_24151,N_22617,N_22118);
xor U24152 (N_24152,N_23881,N_22299);
nor U24153 (N_24153,N_22104,N_22175);
or U24154 (N_24154,N_22562,N_21977);
nor U24155 (N_24155,N_23543,N_21555);
nand U24156 (N_24156,N_23975,N_23011);
and U24157 (N_24157,N_23266,N_21862);
nor U24158 (N_24158,N_21660,N_21195);
nand U24159 (N_24159,N_22154,N_21278);
xnor U24160 (N_24160,N_23782,N_22794);
xor U24161 (N_24161,N_23460,N_21262);
and U24162 (N_24162,N_21193,N_22631);
and U24163 (N_24163,N_23943,N_23003);
nor U24164 (N_24164,N_21724,N_23225);
or U24165 (N_24165,N_21207,N_23873);
nand U24166 (N_24166,N_23976,N_22654);
nand U24167 (N_24167,N_21413,N_23855);
nor U24168 (N_24168,N_21378,N_23268);
nand U24169 (N_24169,N_21515,N_22359);
or U24170 (N_24170,N_22977,N_22295);
and U24171 (N_24171,N_21225,N_23420);
or U24172 (N_24172,N_21787,N_21112);
xor U24173 (N_24173,N_22440,N_22899);
nor U24174 (N_24174,N_21269,N_22199);
and U24175 (N_24175,N_23201,N_22532);
or U24176 (N_24176,N_21155,N_23442);
xnor U24177 (N_24177,N_21664,N_21857);
nor U24178 (N_24178,N_22128,N_22346);
nor U24179 (N_24179,N_22021,N_22699);
and U24180 (N_24180,N_22986,N_23160);
nor U24181 (N_24181,N_21872,N_21498);
nor U24182 (N_24182,N_23807,N_23694);
nor U24183 (N_24183,N_22759,N_21394);
nor U24184 (N_24184,N_22824,N_21403);
or U24185 (N_24185,N_21154,N_21230);
and U24186 (N_24186,N_23780,N_23455);
xor U24187 (N_24187,N_22939,N_22724);
and U24188 (N_24188,N_21077,N_23568);
nand U24189 (N_24189,N_22139,N_22488);
and U24190 (N_24190,N_23063,N_21604);
nand U24191 (N_24191,N_21997,N_22360);
nand U24192 (N_24192,N_23838,N_22545);
nand U24193 (N_24193,N_22369,N_23370);
and U24194 (N_24194,N_21081,N_23031);
and U24195 (N_24195,N_23559,N_23544);
nand U24196 (N_24196,N_22707,N_23858);
nand U24197 (N_24197,N_21076,N_23938);
nor U24198 (N_24198,N_21605,N_21314);
xor U24199 (N_24199,N_22246,N_21487);
or U24200 (N_24200,N_22443,N_22168);
nand U24201 (N_24201,N_23091,N_22957);
nand U24202 (N_24202,N_22005,N_21510);
and U24203 (N_24203,N_21643,N_21493);
or U24204 (N_24204,N_21048,N_23149);
nor U24205 (N_24205,N_23134,N_22838);
or U24206 (N_24206,N_21878,N_21780);
and U24207 (N_24207,N_22328,N_22071);
or U24208 (N_24208,N_22050,N_22234);
and U24209 (N_24209,N_21352,N_23472);
xor U24210 (N_24210,N_22011,N_22242);
nor U24211 (N_24211,N_22044,N_21615);
or U24212 (N_24212,N_21858,N_23507);
xor U24213 (N_24213,N_23671,N_21095);
and U24214 (N_24214,N_23421,N_22810);
xor U24215 (N_24215,N_21557,N_23148);
xnor U24216 (N_24216,N_21672,N_21252);
xor U24217 (N_24217,N_23557,N_22221);
and U24218 (N_24218,N_22834,N_22637);
nor U24219 (N_24219,N_23699,N_21023);
xnor U24220 (N_24220,N_22244,N_21580);
nor U24221 (N_24221,N_22720,N_22626);
or U24222 (N_24222,N_21795,N_22432);
nand U24223 (N_24223,N_23735,N_22051);
and U24224 (N_24224,N_23566,N_22090);
or U24225 (N_24225,N_21669,N_21167);
or U24226 (N_24226,N_22641,N_21638);
and U24227 (N_24227,N_22835,N_23742);
xnor U24228 (N_24228,N_21684,N_21354);
xor U24229 (N_24229,N_21236,N_22945);
or U24230 (N_24230,N_23395,N_21758);
nand U24231 (N_24231,N_21159,N_21574);
nand U24232 (N_24232,N_22238,N_22754);
or U24233 (N_24233,N_22785,N_22703);
and U24234 (N_24234,N_23588,N_23363);
nor U24235 (N_24235,N_23066,N_21074);
nand U24236 (N_24236,N_23590,N_22800);
nand U24237 (N_24237,N_23785,N_23186);
xor U24238 (N_24238,N_23902,N_22535);
xnor U24239 (N_24239,N_22110,N_23852);
or U24240 (N_24240,N_21824,N_23964);
nor U24241 (N_24241,N_22141,N_23836);
nand U24242 (N_24242,N_22279,N_22738);
xnor U24243 (N_24243,N_21889,N_23504);
nor U24244 (N_24244,N_22192,N_23383);
or U24245 (N_24245,N_23261,N_23646);
and U24246 (N_24246,N_21424,N_22039);
and U24247 (N_24247,N_22544,N_23633);
xnor U24248 (N_24248,N_23577,N_21449);
and U24249 (N_24249,N_23848,N_22479);
nand U24250 (N_24250,N_21968,N_23607);
nand U24251 (N_24251,N_21573,N_22893);
or U24252 (N_24252,N_23461,N_22144);
and U24253 (N_24253,N_23367,N_21002);
and U24254 (N_24254,N_21319,N_22937);
nand U24255 (N_24255,N_22065,N_23686);
and U24256 (N_24256,N_23039,N_22407);
or U24257 (N_24257,N_22303,N_22287);
nand U24258 (N_24258,N_23102,N_21879);
nor U24259 (N_24259,N_22938,N_22883);
nor U24260 (N_24260,N_23038,N_23407);
nor U24261 (N_24261,N_22704,N_21798);
or U24262 (N_24262,N_21897,N_21822);
nand U24263 (N_24263,N_21239,N_22656);
nand U24264 (N_24264,N_23154,N_21584);
or U24265 (N_24265,N_23494,N_21630);
nand U24266 (N_24266,N_22892,N_21633);
nand U24267 (N_24267,N_21942,N_23313);
xnor U24268 (N_24268,N_21886,N_21381);
or U24269 (N_24269,N_22702,N_23247);
nor U24270 (N_24270,N_23350,N_22022);
and U24271 (N_24271,N_21375,N_22477);
and U24272 (N_24272,N_21520,N_21126);
nor U24273 (N_24273,N_23680,N_21307);
nor U24274 (N_24274,N_21482,N_23248);
nor U24275 (N_24275,N_22811,N_21402);
xnor U24276 (N_24276,N_23006,N_22612);
and U24277 (N_24277,N_23463,N_23745);
and U24278 (N_24278,N_23546,N_21710);
and U24279 (N_24279,N_21224,N_21379);
xnor U24280 (N_24280,N_22447,N_23479);
and U24281 (N_24281,N_23891,N_21080);
and U24282 (N_24282,N_23892,N_22233);
xor U24283 (N_24283,N_23079,N_23966);
xor U24284 (N_24284,N_21025,N_21980);
or U24285 (N_24285,N_23803,N_21545);
nor U24286 (N_24286,N_21754,N_21836);
nor U24287 (N_24287,N_22158,N_22292);
and U24288 (N_24288,N_23850,N_21172);
xnor U24289 (N_24289,N_22207,N_21250);
nor U24290 (N_24290,N_21342,N_21755);
and U24291 (N_24291,N_22456,N_22278);
xnor U24292 (N_24292,N_23021,N_22958);
nand U24293 (N_24293,N_22793,N_22764);
or U24294 (N_24294,N_23603,N_22431);
nor U24295 (N_24295,N_21567,N_23503);
or U24296 (N_24296,N_22404,N_21948);
or U24297 (N_24297,N_21200,N_21433);
or U24298 (N_24298,N_21175,N_23314);
xor U24299 (N_24299,N_23271,N_22978);
and U24300 (N_24300,N_23740,N_22107);
nand U24301 (N_24301,N_21995,N_22991);
xor U24302 (N_24302,N_23369,N_21044);
and U24303 (N_24303,N_22010,N_21779);
nor U24304 (N_24304,N_23874,N_22084);
nand U24305 (N_24305,N_22992,N_22582);
nand U24306 (N_24306,N_21655,N_22136);
or U24307 (N_24307,N_23424,N_21376);
nand U24308 (N_24308,N_23798,N_23484);
and U24309 (N_24309,N_22831,N_23679);
or U24310 (N_24310,N_23099,N_21949);
nor U24311 (N_24311,N_23763,N_22137);
nand U24312 (N_24312,N_22027,N_23138);
nor U24313 (N_24313,N_22445,N_22729);
nor U24314 (N_24314,N_22782,N_21827);
xor U24315 (N_24315,N_21241,N_21201);
xor U24316 (N_24316,N_22083,N_21294);
nand U24317 (N_24317,N_22392,N_21676);
nor U24318 (N_24318,N_22894,N_23653);
nor U24319 (N_24319,N_23007,N_22969);
nor U24320 (N_24320,N_23080,N_21599);
and U24321 (N_24321,N_23258,N_22105);
nor U24322 (N_24322,N_21728,N_21255);
and U24323 (N_24323,N_21715,N_21321);
or U24324 (N_24324,N_21476,N_22362);
and U24325 (N_24325,N_22507,N_22519);
nand U24326 (N_24326,N_21223,N_23602);
nand U24327 (N_24327,N_23346,N_21060);
nor U24328 (N_24328,N_22775,N_21037);
xor U24329 (N_24329,N_21812,N_22563);
and U24330 (N_24330,N_23375,N_21543);
and U24331 (N_24331,N_23884,N_23127);
or U24332 (N_24332,N_22798,N_21473);
xnor U24333 (N_24333,N_22349,N_23897);
and U24334 (N_24334,N_22040,N_21677);
or U24335 (N_24335,N_23534,N_21004);
and U24336 (N_24336,N_21559,N_22734);
nand U24337 (N_24337,N_22815,N_23016);
or U24338 (N_24338,N_21777,N_21070);
and U24339 (N_24339,N_22391,N_22671);
xnor U24340 (N_24340,N_21393,N_21888);
xnor U24341 (N_24341,N_22337,N_22224);
nand U24342 (N_24342,N_21934,N_22284);
nand U24343 (N_24343,N_23522,N_23556);
nor U24344 (N_24344,N_23684,N_23233);
nand U24345 (N_24345,N_21870,N_23841);
and U24346 (N_24346,N_22747,N_21075);
or U24347 (N_24347,N_21299,N_21310);
nand U24348 (N_24348,N_22898,N_23769);
nand U24349 (N_24349,N_22293,N_23914);
xnor U24350 (N_24350,N_22905,N_23610);
or U24351 (N_24351,N_23311,N_22881);
xor U24352 (N_24352,N_22896,N_22455);
and U24353 (N_24353,N_23660,N_22901);
xor U24354 (N_24354,N_21137,N_23755);
xor U24355 (N_24355,N_22576,N_23744);
or U24356 (N_24356,N_21067,N_22259);
and U24357 (N_24357,N_22210,N_21332);
nor U24358 (N_24358,N_23648,N_23084);
and U24359 (N_24359,N_21701,N_22159);
xor U24360 (N_24360,N_21174,N_23100);
nor U24361 (N_24361,N_21385,N_22363);
nand U24362 (N_24362,N_23046,N_23302);
xor U24363 (N_24363,N_23364,N_23280);
nor U24364 (N_24364,N_21517,N_21783);
and U24365 (N_24365,N_21800,N_23008);
nor U24366 (N_24366,N_23622,N_23857);
or U24367 (N_24367,N_21313,N_22965);
and U24368 (N_24368,N_22062,N_23935);
nand U24369 (N_24369,N_21446,N_23528);
xor U24370 (N_24370,N_23842,N_22318);
or U24371 (N_24371,N_21205,N_22814);
nor U24372 (N_24372,N_23044,N_21212);
nor U24373 (N_24373,N_21963,N_23324);
or U24374 (N_24374,N_22897,N_22552);
xnor U24375 (N_24375,N_21302,N_21259);
or U24376 (N_24376,N_23473,N_21884);
nor U24377 (N_24377,N_21102,N_23987);
and U24378 (N_24378,N_21962,N_21478);
or U24379 (N_24379,N_21349,N_23262);
xnor U24380 (N_24380,N_21500,N_23562);
xor U24381 (N_24381,N_23249,N_22498);
nand U24382 (N_24382,N_23012,N_21536);
or U24383 (N_24383,N_21055,N_23520);
nand U24384 (N_24384,N_21887,N_22967);
nand U24385 (N_24385,N_23643,N_23918);
nand U24386 (N_24386,N_22756,N_23811);
and U24387 (N_24387,N_23078,N_22496);
nand U24388 (N_24388,N_22116,N_23707);
and U24389 (N_24389,N_22099,N_21885);
and U24390 (N_24390,N_21450,N_22481);
and U24391 (N_24391,N_23283,N_23862);
and U24392 (N_24392,N_23737,N_22780);
xnor U24393 (N_24393,N_23783,N_23491);
or U24394 (N_24394,N_22988,N_22334);
xnor U24395 (N_24395,N_22540,N_22776);
and U24396 (N_24396,N_23917,N_21451);
and U24397 (N_24397,N_21362,N_22033);
and U24398 (N_24398,N_23250,N_21909);
xor U24399 (N_24399,N_22602,N_22045);
nor U24400 (N_24400,N_23876,N_23541);
or U24401 (N_24401,N_23894,N_23813);
nor U24402 (N_24402,N_21436,N_23721);
xor U24403 (N_24403,N_21338,N_21524);
or U24404 (N_24404,N_22112,N_22161);
nand U24405 (N_24405,N_21353,N_21595);
nand U24406 (N_24406,N_22615,N_21550);
nor U24407 (N_24407,N_22253,N_22147);
or U24408 (N_24408,N_21084,N_22891);
and U24409 (N_24409,N_23093,N_22678);
and U24410 (N_24410,N_21964,N_23781);
nor U24411 (N_24411,N_22066,N_22721);
or U24412 (N_24412,N_21087,N_22917);
nor U24413 (N_24413,N_23361,N_23765);
nor U24414 (N_24414,N_23042,N_23366);
nand U24415 (N_24415,N_21637,N_22366);
nand U24416 (N_24416,N_23440,N_21837);
or U24417 (N_24417,N_22580,N_21566);
and U24418 (N_24418,N_22439,N_22108);
xnor U24419 (N_24419,N_22655,N_23152);
nand U24420 (N_24420,N_22658,N_22020);
nor U24421 (N_24421,N_21959,N_23453);
or U24422 (N_24422,N_22711,N_21691);
and U24423 (N_24423,N_23770,N_22941);
and U24424 (N_24424,N_23432,N_22348);
or U24425 (N_24425,N_23058,N_22845);
nor U24426 (N_24426,N_22871,N_21392);
or U24427 (N_24427,N_23772,N_23898);
xor U24428 (N_24428,N_21467,N_21531);
or U24429 (N_24429,N_23337,N_23736);
nor U24430 (N_24430,N_23517,N_23703);
xor U24431 (N_24431,N_23119,N_23057);
xor U24432 (N_24432,N_23073,N_22604);
xnor U24433 (N_24433,N_22046,N_22098);
and U24434 (N_24434,N_21014,N_22832);
and U24435 (N_24435,N_22980,N_23114);
nand U24436 (N_24436,N_21317,N_21292);
or U24437 (N_24437,N_22907,N_22353);
nand U24438 (N_24438,N_23980,N_21211);
and U24439 (N_24439,N_23483,N_22593);
nand U24440 (N_24440,N_22607,N_21158);
nand U24441 (N_24441,N_22398,N_21142);
nand U24442 (N_24442,N_21969,N_22770);
or U24443 (N_24443,N_21966,N_23804);
or U24444 (N_24444,N_21086,N_21143);
nor U24445 (N_24445,N_23663,N_21497);
nand U24446 (N_24446,N_23909,N_21782);
nor U24447 (N_24447,N_21898,N_21490);
xnor U24448 (N_24448,N_21128,N_21202);
nand U24449 (N_24449,N_22741,N_22869);
and U24450 (N_24450,N_22610,N_23101);
or U24451 (N_24451,N_23069,N_22146);
xnor U24452 (N_24452,N_21797,N_21985);
nand U24453 (N_24453,N_21073,N_23287);
nor U24454 (N_24454,N_23509,N_23325);
xor U24455 (N_24455,N_21597,N_21592);
xnor U24456 (N_24456,N_22296,N_21558);
xnor U24457 (N_24457,N_22204,N_21178);
or U24458 (N_24458,N_21748,N_22531);
xnor U24459 (N_24459,N_22063,N_22243);
nand U24460 (N_24460,N_21505,N_22429);
and U24461 (N_24461,N_21644,N_23372);
xnor U24462 (N_24462,N_22125,N_22568);
nor U24463 (N_24463,N_22232,N_23617);
xor U24464 (N_24464,N_23578,N_21192);
and U24465 (N_24465,N_23594,N_21363);
nor U24466 (N_24466,N_23028,N_23571);
or U24467 (N_24467,N_21096,N_23060);
xnor U24468 (N_24468,N_23124,N_22737);
nor U24469 (N_24469,N_22426,N_22068);
nor U24470 (N_24470,N_23551,N_21869);
nand U24471 (N_24471,N_22599,N_23071);
and U24472 (N_24472,N_21513,N_22474);
and U24473 (N_24473,N_22692,N_23709);
xnor U24474 (N_24474,N_22584,N_21244);
nor U24475 (N_24475,N_21203,N_21345);
and U24476 (N_24476,N_23117,N_23936);
xnor U24477 (N_24477,N_21547,N_23642);
and U24478 (N_24478,N_23893,N_22501);
xor U24479 (N_24479,N_22515,N_21213);
nand U24480 (N_24480,N_23104,N_21571);
nor U24481 (N_24481,N_21518,N_22317);
nor U24482 (N_24482,N_21526,N_23128);
nor U24483 (N_24483,N_22718,N_21861);
nor U24484 (N_24484,N_21343,N_21667);
or U24485 (N_24485,N_21412,N_21350);
or U24486 (N_24486,N_22997,N_23171);
nand U24487 (N_24487,N_21841,N_22371);
xor U24488 (N_24488,N_23385,N_21246);
and U24489 (N_24489,N_23129,N_22167);
and U24490 (N_24490,N_22739,N_21382);
or U24491 (N_24491,N_21064,N_22380);
xnor U24492 (N_24492,N_23885,N_22884);
or U24493 (N_24493,N_23462,N_21383);
and U24494 (N_24494,N_21136,N_22281);
xor U24495 (N_24495,N_23844,N_23767);
or U24496 (N_24496,N_21227,N_22876);
nand U24497 (N_24497,N_23627,N_21113);
and U24498 (N_24498,N_21411,N_22628);
and U24499 (N_24499,N_21906,N_23317);
nor U24500 (N_24500,N_21365,N_21859);
nor U24501 (N_24501,N_22821,N_21698);
and U24502 (N_24502,N_22247,N_22783);
or U24503 (N_24503,N_22927,N_21355);
nor U24504 (N_24504,N_23118,N_23570);
xnor U24505 (N_24505,N_22130,N_22943);
nor U24506 (N_24506,N_22989,N_21789);
and U24507 (N_24507,N_23125,N_21162);
xor U24508 (N_24508,N_23147,N_22638);
nor U24509 (N_24509,N_23871,N_21951);
or U24510 (N_24510,N_21032,N_23439);
or U24511 (N_24511,N_22179,N_21528);
nand U24512 (N_24512,N_21471,N_22581);
or U24513 (N_24513,N_22057,N_23634);
and U24514 (N_24514,N_21958,N_21683);
and U24515 (N_24515,N_21457,N_21123);
or U24516 (N_24516,N_21645,N_21688);
xor U24517 (N_24517,N_23817,N_23941);
and U24518 (N_24518,N_21160,N_21548);
nand U24519 (N_24519,N_21650,N_23009);
or U24520 (N_24520,N_23146,N_22142);
nor U24521 (N_24521,N_22082,N_21591);
xnor U24522 (N_24522,N_23428,N_23110);
and U24523 (N_24523,N_21017,N_22323);
nor U24524 (N_24524,N_21161,N_22231);
nand U24525 (N_24525,N_23065,N_23215);
nand U24526 (N_24526,N_21456,N_21716);
nand U24527 (N_24527,N_22670,N_22839);
nor U24528 (N_24528,N_22786,N_23315);
and U24529 (N_24529,N_22236,N_21093);
or U24530 (N_24530,N_22795,N_21972);
nand U24531 (N_24531,N_21692,N_22960);
nand U24532 (N_24532,N_23673,N_21750);
nand U24533 (N_24533,N_21180,N_23505);
xor U24534 (N_24534,N_23150,N_23379);
or U24535 (N_24535,N_21329,N_22372);
nor U24536 (N_24536,N_22261,N_23845);
nand U24537 (N_24537,N_22223,N_22351);
nor U24538 (N_24538,N_22209,N_22352);
xnor U24539 (N_24539,N_23037,N_23061);
nand U24540 (N_24540,N_23523,N_23814);
nor U24541 (N_24541,N_22885,N_21565);
or U24542 (N_24542,N_22572,N_23320);
and U24543 (N_24543,N_21936,N_21168);
nand U24544 (N_24544,N_23458,N_22996);
nand U24545 (N_24545,N_21138,N_23214);
nor U24546 (N_24546,N_22288,N_21374);
or U24547 (N_24547,N_21881,N_22954);
nand U24548 (N_24548,N_23678,N_22712);
or U24549 (N_24549,N_22690,N_21204);
nand U24550 (N_24550,N_23589,N_21632);
nand U24551 (N_24551,N_23308,N_22940);
or U24552 (N_24552,N_21026,N_23698);
nand U24553 (N_24553,N_22636,N_23856);
or U24554 (N_24554,N_22408,N_22187);
nor U24555 (N_24555,N_23024,N_21785);
nand U24556 (N_24556,N_23575,N_21720);
or U24557 (N_24557,N_23286,N_22000);
nor U24558 (N_24558,N_23982,N_23401);
xnor U24559 (N_24559,N_21868,N_22361);
nor U24560 (N_24560,N_21031,N_21298);
xor U24561 (N_24561,N_21892,N_23467);
and U24562 (N_24562,N_23700,N_21747);
xnor U24563 (N_24563,N_22661,N_22450);
nand U24564 (N_24564,N_23688,N_21725);
nor U24565 (N_24565,N_23300,N_21441);
or U24566 (N_24566,N_21078,N_21873);
nand U24567 (N_24567,N_21512,N_22812);
xnor U24568 (N_24568,N_21809,N_22064);
and U24569 (N_24569,N_21593,N_23211);
nand U24570 (N_24570,N_23984,N_21611);
nor U24571 (N_24571,N_23339,N_21953);
xnor U24572 (N_24572,N_21327,N_21367);
and U24573 (N_24573,N_21663,N_23624);
nand U24574 (N_24574,N_22342,N_22487);
or U24575 (N_24575,N_23580,N_23689);
nand U24576 (N_24576,N_21431,N_23636);
nand U24577 (N_24577,N_23934,N_22557);
or U24578 (N_24578,N_23711,N_21749);
or U24579 (N_24579,N_23045,N_21094);
nor U24580 (N_24580,N_21978,N_21852);
or U24581 (N_24581,N_21553,N_21662);
nor U24582 (N_24582,N_21551,N_22422);
or U24583 (N_24583,N_22276,N_22922);
and U24584 (N_24584,N_21121,N_22131);
nand U24585 (N_24585,N_23854,N_22560);
and U24586 (N_24586,N_22526,N_23625);
or U24587 (N_24587,N_23754,N_23928);
nand U24588 (N_24588,N_23106,N_23651);
xor U24589 (N_24589,N_21753,N_22416);
nor U24590 (N_24590,N_23345,N_23750);
or U24591 (N_24591,N_21333,N_21905);
xnor U24592 (N_24592,N_22595,N_21468);
xnor U24593 (N_24593,N_22180,N_21856);
and U24594 (N_24594,N_23806,N_22826);
nor U24595 (N_24595,N_23900,N_21293);
nand U24596 (N_24596,N_23116,N_23123);
nor U24597 (N_24597,N_21900,N_21083);
xor U24598 (N_24598,N_22514,N_23552);
and U24599 (N_24599,N_23184,N_23229);
or U24600 (N_24600,N_22201,N_22076);
nand U24601 (N_24601,N_21955,N_21602);
or U24602 (N_24602,N_21320,N_23574);
nand U24603 (N_24603,N_22908,N_22662);
and U24604 (N_24604,N_22235,N_22282);
xnor U24605 (N_24605,N_22009,N_21486);
and U24606 (N_24606,N_21699,N_21652);
xor U24607 (N_24607,N_22668,N_21871);
and U24608 (N_24608,N_23135,N_21903);
nand U24609 (N_24609,N_22446,N_22553);
xnor U24610 (N_24610,N_23921,N_22727);
xor U24611 (N_24611,N_22473,N_22657);
nor U24612 (N_24612,N_21006,N_22564);
nand U24613 (N_24613,N_23329,N_21740);
nor U24614 (N_24614,N_22072,N_23296);
nor U24615 (N_24615,N_22579,N_22034);
and U24616 (N_24616,N_21848,N_23418);
or U24617 (N_24617,N_22340,N_23377);
nor U24618 (N_24618,N_23758,N_21297);
nand U24619 (N_24619,N_23410,N_23020);
and U24620 (N_24620,N_22589,N_22588);
nor U24621 (N_24621,N_21097,N_21335);
nor U24622 (N_24622,N_21880,N_22036);
or U24623 (N_24623,N_23961,N_22561);
nand U24624 (N_24624,N_21902,N_21254);
nand U24625 (N_24625,N_22936,N_22388);
nor U24626 (N_24626,N_23939,N_21727);
nor U24627 (N_24627,N_23153,N_23985);
and U24628 (N_24628,N_23880,N_23614);
xor U24629 (N_24629,N_21415,N_22921);
and U24630 (N_24630,N_22983,N_22280);
and U24631 (N_24631,N_22855,N_22401);
nand U24632 (N_24632,N_22804,N_23142);
nor U24633 (N_24633,N_22262,N_23554);
and U24634 (N_24634,N_22829,N_22405);
or U24635 (N_24635,N_22387,N_21647);
xor U24636 (N_24636,N_23759,N_22982);
or U24637 (N_24637,N_21826,N_22889);
xor U24638 (N_24638,N_23404,N_23168);
and U24639 (N_24639,N_22609,N_22433);
xnor U24640 (N_24640,N_23202,N_21577);
xnor U24641 (N_24641,N_22620,N_22616);
and U24642 (N_24642,N_21998,N_23362);
nand U24643 (N_24643,N_22925,N_21035);
nor U24644 (N_24644,N_21546,N_22283);
or U24645 (N_24645,N_22002,N_22402);
and U24646 (N_24646,N_21464,N_23542);
nand U24647 (N_24647,N_21802,N_22442);
nand U24648 (N_24648,N_23396,N_22748);
or U24649 (N_24649,N_22364,N_23212);
or U24650 (N_24650,N_21019,N_23081);
xnor U24651 (N_24651,N_21268,N_21640);
and U24652 (N_24652,N_22987,N_22651);
nand U24653 (N_24653,N_23581,N_23877);
nand U24654 (N_24654,N_21917,N_22302);
nor U24655 (N_24655,N_23705,N_22390);
nor U24656 (N_24656,N_22495,N_23109);
nor U24657 (N_24657,N_23993,N_22042);
xor U24658 (N_24658,N_23829,N_21290);
and U24659 (N_24659,N_23299,N_21675);
or U24660 (N_24660,N_21001,N_23488);
nor U24661 (N_24661,N_21007,N_21051);
or U24662 (N_24662,N_21830,N_22170);
nand U24663 (N_24663,N_21818,N_22947);
xor U24664 (N_24664,N_21000,N_22484);
nor U24665 (N_24665,N_22263,N_23425);
nor U24666 (N_24666,N_23822,N_21616);
nor U24667 (N_24667,N_22218,N_22648);
nand U24668 (N_24668,N_21439,N_23847);
nor U24669 (N_24669,N_21181,N_23036);
nor U24670 (N_24670,N_23357,N_23301);
nand U24671 (N_24671,N_23766,N_21085);
nand U24672 (N_24672,N_22256,N_21043);
xnor U24673 (N_24673,N_22149,N_21406);
and U24674 (N_24674,N_22830,N_21115);
nor U24675 (N_24675,N_22751,N_23724);
nor U24676 (N_24676,N_21435,N_21484);
nand U24677 (N_24677,N_23349,N_23792);
nand U24678 (N_24678,N_21134,N_21717);
xnor U24679 (N_24679,N_21924,N_21696);
nor U24680 (N_24680,N_22106,N_21588);
and U24681 (N_24681,N_22928,N_22124);
nor U24682 (N_24682,N_22614,N_23572);
nor U24683 (N_24683,N_22669,N_22503);
nand U24684 (N_24684,N_22550,N_21771);
xnor U24685 (N_24685,N_22480,N_23365);
nor U24686 (N_24686,N_21731,N_22627);
or U24687 (N_24687,N_21578,N_22842);
and U24688 (N_24688,N_21282,N_22666);
nand U24689 (N_24689,N_22325,N_21417);
nor U24690 (N_24690,N_23384,N_23793);
or U24691 (N_24691,N_22530,N_23259);
nor U24692 (N_24692,N_23951,N_23919);
xor U24693 (N_24693,N_22710,N_22041);
and U24694 (N_24694,N_23816,N_22054);
and U24695 (N_24695,N_21146,N_23913);
xor U24696 (N_24696,N_21661,N_22877);
or U24697 (N_24697,N_21220,N_23108);
xnor U24698 (N_24698,N_22367,N_23701);
nor U24699 (N_24699,N_21606,N_22763);
and U24700 (N_24700,N_21988,N_23392);
or U24701 (N_24701,N_22249,N_23957);
xnor U24702 (N_24702,N_22102,N_22590);
or U24703 (N_24703,N_22089,N_22948);
xnor U24704 (N_24704,N_21625,N_22758);
nor U24705 (N_24705,N_23693,N_23965);
or U24706 (N_24706,N_21678,N_23818);
or U24707 (N_24707,N_23799,N_23833);
nor U24708 (N_24708,N_22166,N_21430);
and U24709 (N_24709,N_21954,N_23514);
xnor U24710 (N_24710,N_22285,N_23824);
nor U24711 (N_24711,N_22080,N_22056);
nand U24712 (N_24712,N_23502,N_21184);
nand U24713 (N_24713,N_22188,N_23555);
and U24714 (N_24714,N_21539,N_22730);
nor U24715 (N_24715,N_23355,N_23417);
xor U24716 (N_24716,N_22547,N_22023);
nand U24717 (N_24717,N_22448,N_22846);
nand U24718 (N_24718,N_23959,N_21491);
nand U24719 (N_24719,N_22081,N_23294);
nand U24720 (N_24720,N_23082,N_21423);
xor U24721 (N_24721,N_21530,N_21380);
or U24722 (N_24722,N_23468,N_23601);
nor U24723 (N_24723,N_23216,N_22861);
xor U24724 (N_24724,N_22373,N_22613);
or U24725 (N_24725,N_22078,N_23105);
nor U24726 (N_24726,N_21839,N_22828);
xnor U24727 (N_24727,N_23727,N_21011);
xor U24728 (N_24728,N_21300,N_23786);
nand U24729 (N_24729,N_23143,N_21883);
xor U24730 (N_24730,N_21849,N_23681);
nand U24731 (N_24731,N_23591,N_22240);
or U24732 (N_24732,N_23741,N_22271);
nor U24733 (N_24733,N_22878,N_22566);
nor U24734 (N_24734,N_21961,N_23482);
xnor U24735 (N_24735,N_23837,N_21389);
xor U24736 (N_24736,N_23336,N_21100);
nand U24737 (N_24737,N_23070,N_21617);
and U24738 (N_24738,N_22672,N_23406);
xnor U24739 (N_24739,N_22725,N_23915);
or U24740 (N_24740,N_22975,N_22968);
xnor U24741 (N_24741,N_23569,N_23956);
nor U24742 (N_24742,N_21330,N_22859);
xnor U24743 (N_24743,N_22621,N_23743);
nor U24744 (N_24744,N_21272,N_21177);
nand U24745 (N_24745,N_22413,N_23470);
and U24746 (N_24746,N_23661,N_21425);
or U24747 (N_24747,N_23306,N_22858);
or U24748 (N_24748,N_21005,N_21266);
nor U24749 (N_24749,N_23878,N_21732);
and U24750 (N_24750,N_21318,N_23952);
nor U24751 (N_24751,N_22909,N_22376);
xnor U24752 (N_24752,N_22230,N_22949);
nand U24753 (N_24753,N_21316,N_22732);
nor U24754 (N_24754,N_23846,N_21104);
or U24755 (N_24755,N_22461,N_21141);
nor U24756 (N_24756,N_21315,N_22971);
nand U24757 (N_24757,N_22435,N_22478);
and U24758 (N_24758,N_22245,N_23279);
nor U24759 (N_24759,N_23903,N_23889);
nor U24760 (N_24760,N_21974,N_23052);
and U24761 (N_24761,N_23427,N_22286);
nor U24762 (N_24762,N_23550,N_21989);
and U24763 (N_24763,N_21741,N_21488);
or U24764 (N_24764,N_22119,N_22652);
or U24765 (N_24765,N_23120,N_21930);
xor U24766 (N_24766,N_23685,N_23756);
nand U24767 (N_24767,N_22875,N_23382);
or U24768 (N_24768,N_23398,N_22421);
xor U24769 (N_24769,N_23805,N_21766);
nor U24770 (N_24770,N_22008,N_21122);
nor U24771 (N_24771,N_23540,N_23911);
nor U24772 (N_24772,N_21635,N_22906);
xor U24773 (N_24773,N_22771,N_22942);
nor U24774 (N_24774,N_23328,N_23537);
nor U24775 (N_24775,N_22031,N_22914);
xor U24776 (N_24776,N_22549,N_23669);
nand U24777 (N_24777,N_21796,N_23506);
or U24778 (N_24778,N_23196,N_23312);
nand U24779 (N_24779,N_22470,N_22802);
nand U24780 (N_24780,N_21621,N_23048);
or U24781 (N_24781,N_22966,N_23989);
xnor U24782 (N_24782,N_21370,N_21147);
and U24783 (N_24783,N_21623,N_23790);
nand U24784 (N_24784,N_22976,N_22964);
or U24785 (N_24785,N_21916,N_22320);
xnor U24786 (N_24786,N_22870,N_22177);
and U24787 (N_24787,N_23524,N_22059);
xnor U24788 (N_24788,N_23726,N_23823);
nor U24789 (N_24789,N_22229,N_23843);
nand U24790 (N_24790,N_21066,N_21477);
and U24791 (N_24791,N_22930,N_21807);
and U24792 (N_24792,N_23677,N_21793);
and U24793 (N_24793,N_21120,N_23564);
or U24794 (N_24794,N_23137,N_22833);
nand U24795 (N_24795,N_23035,N_21967);
nand U24796 (N_24796,N_22886,N_23213);
or U24797 (N_24797,N_23068,N_21874);
xor U24798 (N_24798,N_22241,N_22541);
or U24799 (N_24799,N_21819,N_23429);
or U24800 (N_24800,N_21950,N_21058);
nand U24801 (N_24801,N_23916,N_22308);
nor U24802 (N_24802,N_23826,N_22140);
nor U24803 (N_24803,N_21992,N_23870);
nor U24804 (N_24804,N_22805,N_23553);
nand U24805 (N_24805,N_22160,N_21016);
nand U24806 (N_24806,N_23596,N_23158);
xnor U24807 (N_24807,N_21570,N_21556);
xor U24808 (N_24808,N_22578,N_22397);
and U24809 (N_24809,N_23162,N_23027);
and U24810 (N_24810,N_21784,N_23820);
or U24811 (N_24811,N_21041,N_22848);
nand U24812 (N_24812,N_22512,N_22255);
nand U24813 (N_24813,N_23715,N_21893);
xnor U24814 (N_24814,N_21229,N_21427);
and U24815 (N_24815,N_23788,N_23285);
and U24816 (N_24816,N_22185,N_22569);
or U24817 (N_24817,N_22156,N_21534);
xor U24818 (N_24818,N_22873,N_23288);
nand U24819 (N_24819,N_21774,N_23276);
or U24820 (N_24820,N_23953,N_22822);
or U24821 (N_24821,N_22935,N_22471);
xnor U24822 (N_24822,N_23459,N_21943);
or U24823 (N_24823,N_21922,N_22809);
and U24824 (N_24824,N_22272,N_23628);
xnor U24825 (N_24825,N_21907,N_22091);
nand U24826 (N_24826,N_21508,N_22571);
and U24827 (N_24827,N_21915,N_21853);
and U24828 (N_24828,N_21222,N_22733);
xor U24829 (N_24829,N_21176,N_22451);
nand U24830 (N_24830,N_22150,N_23644);
and U24831 (N_24831,N_23430,N_21651);
and U24832 (N_24832,N_23639,N_21189);
xor U24833 (N_24833,N_22929,N_22355);
nand U24834 (N_24834,N_22536,N_22803);
nand U24835 (N_24835,N_23549,N_21153);
nor U24836 (N_24836,N_23777,N_23932);
and U24837 (N_24837,N_23971,N_22517);
xnor U24838 (N_24838,N_21521,N_22409);
nor U24839 (N_24839,N_22597,N_23333);
and U24840 (N_24840,N_23097,N_22801);
nand U24841 (N_24841,N_21769,N_21712);
nand U24842 (N_24842,N_22632,N_23032);
nor U24843 (N_24843,N_21773,N_23933);
or U24844 (N_24844,N_22095,N_23521);
or U24845 (N_24845,N_23335,N_21384);
nor U24846 (N_24846,N_21281,N_23631);
and U24847 (N_24847,N_21444,N_21685);
nand U24848 (N_24848,N_23613,N_22680);
nand U24849 (N_24849,N_22681,N_21634);
xor U24850 (N_24850,N_22750,N_21418);
or U24851 (N_24851,N_22113,N_23729);
nor U24852 (N_24852,N_23391,N_22684);
nand U24853 (N_24853,N_22038,N_21947);
nand U24854 (N_24854,N_23492,N_23981);
nor U24855 (N_24855,N_23431,N_22345);
nand U24856 (N_24856,N_21082,N_23378);
nand U24857 (N_24857,N_21360,N_23327);
nor U24858 (N_24858,N_21718,N_21658);
xnor U24859 (N_24859,N_23725,N_21323);
xnor U24860 (N_24860,N_23075,N_22277);
xor U24861 (N_24861,N_21460,N_23156);
nand U24862 (N_24862,N_21761,N_23533);
nand U24863 (N_24863,N_23477,N_21369);
xor U24864 (N_24864,N_23353,N_21834);
xnor U24865 (N_24865,N_23254,N_23227);
nand U24866 (N_24866,N_23072,N_22389);
and U24867 (N_24867,N_22004,N_21618);
nor U24868 (N_24868,N_22151,N_21346);
nand U24869 (N_24869,N_23849,N_23284);
and U24870 (N_24870,N_21582,N_23748);
xnor U24871 (N_24871,N_22260,N_22467);
nand U24872 (N_24872,N_23929,N_23776);
and U24873 (N_24873,N_23465,N_23802);
nor U24874 (N_24874,N_22305,N_23791);
xor U24875 (N_24875,N_21218,N_22411);
and U24876 (N_24876,N_23373,N_23426);
xor U24877 (N_24877,N_23014,N_21079);
and U24878 (N_24878,N_21361,N_21756);
nor U24879 (N_24879,N_21746,N_21186);
nand U24880 (N_24880,N_21831,N_21697);
or U24881 (N_24881,N_22379,N_22001);
or U24882 (N_24882,N_22425,N_21039);
xor U24883 (N_24883,N_23304,N_21535);
xor U24884 (N_24884,N_22689,N_22214);
nand U24885 (N_24885,N_21458,N_21285);
or U24886 (N_24886,N_21116,N_21695);
or U24887 (N_24887,N_22239,N_22250);
and U24888 (N_24888,N_22191,N_22264);
nand U24889 (N_24889,N_21012,N_23618);
nand U24890 (N_24890,N_23638,N_23830);
nand U24891 (N_24891,N_23827,N_22994);
nor U24892 (N_24892,N_21432,N_22777);
xor U24893 (N_24893,N_22386,N_21631);
and U24894 (N_24894,N_23319,N_23872);
nor U24895 (N_24895,N_21671,N_22606);
xor U24896 (N_24896,N_23632,N_21851);
xnor U24897 (N_24897,N_21726,N_22520);
and U24898 (N_24898,N_21799,N_22594);
xnor U24899 (N_24899,N_21921,N_21806);
nand U24900 (N_24900,N_23059,N_21713);
or U24901 (N_24901,N_23434,N_23656);
nor U24902 (N_24902,N_22500,N_21603);
nor U24903 (N_24903,N_21764,N_23695);
xor U24904 (N_24904,N_21933,N_22546);
and U24905 (N_24905,N_22713,N_22841);
or U24906 (N_24906,N_22109,N_21388);
nor U24907 (N_24907,N_23277,N_21514);
nand U24908 (N_24908,N_23221,N_21911);
nand U24909 (N_24909,N_22998,N_22510);
nand U24910 (N_24910,N_23237,N_21428);
xnor U24911 (N_24911,N_23281,N_22145);
nor U24912 (N_24912,N_22012,N_23376);
xnor U24913 (N_24913,N_23974,N_21306);
xor U24914 (N_24914,N_22592,N_21939);
xor U24915 (N_24915,N_21173,N_21790);
xor U24916 (N_24916,N_22735,N_21757);
or U24917 (N_24917,N_22043,N_21422);
nand U24918 (N_24918,N_21410,N_21503);
xnor U24919 (N_24919,N_22539,N_23088);
nand U24920 (N_24920,N_23501,N_23558);
nand U24921 (N_24921,N_21504,N_22472);
xnor U24922 (N_24922,N_21875,N_23176);
nor U24923 (N_24923,N_21438,N_21804);
and U24924 (N_24924,N_21525,N_21303);
or U24925 (N_24925,N_21983,N_22368);
nand U24926 (N_24926,N_22258,N_22779);
nor U24927 (N_24927,N_21492,N_23203);
or U24928 (N_24928,N_21587,N_23389);
xnor U24929 (N_24929,N_21280,N_23586);
or U24930 (N_24930,N_22073,N_21341);
nand U24931 (N_24931,N_21607,N_22951);
nor U24932 (N_24932,N_23821,N_23413);
nor U24933 (N_24933,N_23868,N_22521);
and U24934 (N_24934,N_21021,N_23103);
nor U24935 (N_24935,N_22138,N_23655);
or U24936 (N_24936,N_22676,N_22172);
and U24937 (N_24937,N_21682,N_21908);
and U24938 (N_24938,N_22356,N_22502);
xor U24939 (N_24939,N_21068,N_21564);
or U24940 (N_24940,N_23185,N_21208);
nor U24941 (N_24941,N_23657,N_23466);
nand U24942 (N_24942,N_21975,N_21527);
nor U24943 (N_24943,N_21656,N_21443);
and U24944 (N_24944,N_21131,N_21391);
nor U24945 (N_24945,N_23992,N_21324);
nor U24946 (N_24946,N_21700,N_23979);
or U24947 (N_24947,N_22476,N_22573);
xor U24948 (N_24948,N_22959,N_21040);
or U24949 (N_24949,N_22630,N_23583);
and U24950 (N_24950,N_22736,N_22322);
or U24951 (N_24951,N_22420,N_22061);
or U24952 (N_24952,N_21261,N_21705);
nor U24953 (N_24953,N_21171,N_23863);
nor U24954 (N_24954,N_22316,N_21228);
xnor U24955 (N_24955,N_21059,N_23025);
and U24956 (N_24956,N_22691,N_22452);
and U24957 (N_24957,N_22466,N_22486);
xnor U24958 (N_24958,N_22806,N_23940);
nor U24959 (N_24959,N_23005,N_23561);
nand U24960 (N_24960,N_23717,N_22944);
nor U24961 (N_24961,N_23536,N_21304);
and U24962 (N_24962,N_21594,N_23592);
and U24963 (N_24963,N_21665,N_22981);
or U24964 (N_24964,N_23654,N_22438);
nand U24965 (N_24965,N_22953,N_22096);
xnor U24966 (N_24966,N_22849,N_22772);
nor U24967 (N_24967,N_21091,N_21253);
nand U24968 (N_24968,N_21805,N_22887);
or U24969 (N_24969,N_21359,N_23226);
nor U24970 (N_24970,N_22695,N_22344);
and U24971 (N_24971,N_23356,N_23691);
nand U24972 (N_24972,N_21833,N_21151);
and U24973 (N_24973,N_21653,N_22335);
or U24974 (N_24974,N_22753,N_22625);
or U24975 (N_24975,N_22074,N_22879);
nor U24976 (N_24976,N_23815,N_21711);
nor U24977 (N_24977,N_21850,N_21072);
nand U24978 (N_24978,N_21679,N_23696);
nand U24979 (N_24979,N_22273,N_21305);
or U24980 (N_24980,N_23443,N_23115);
and U24981 (N_24981,N_22490,N_21775);
or U24982 (N_24982,N_21583,N_22910);
or U24983 (N_24983,N_21455,N_22731);
and U24984 (N_24984,N_21737,N_22014);
xnor U24985 (N_24985,N_22270,N_23768);
or U24986 (N_24986,N_22339,N_22624);
or U24987 (N_24987,N_21301,N_22864);
xor U24988 (N_24988,N_22485,N_23133);
xnor U24989 (N_24989,N_22248,N_22762);
nor U24990 (N_24990,N_21781,N_23419);
or U24991 (N_24991,N_23747,N_21744);
nand U24992 (N_24992,N_22924,N_21251);
nand U24993 (N_24993,N_23422,N_21326);
and U24994 (N_24994,N_22673,N_21322);
xor U24995 (N_24995,N_21502,N_22313);
xor U24996 (N_24996,N_22037,N_23761);
xnor U24997 (N_24997,N_22100,N_23746);
xnor U24998 (N_24998,N_23907,N_23265);
nor U24999 (N_24999,N_23995,N_21586);
xnor U25000 (N_25000,N_21736,N_23342);
or U25001 (N_25001,N_21877,N_23665);
nor U25002 (N_25002,N_23192,N_21516);
xnor U25003 (N_25003,N_21941,N_23733);
or U25004 (N_25004,N_22493,N_23794);
nor U25005 (N_25005,N_21165,N_22923);
xor U25006 (N_25006,N_21022,N_21090);
and U25007 (N_25007,N_21276,N_23368);
nand U25008 (N_25008,N_23182,N_23585);
nor U25009 (N_25009,N_23098,N_23344);
and U25010 (N_25010,N_21047,N_22200);
xnor U25011 (N_25011,N_22634,N_23942);
and U25012 (N_25012,N_23054,N_23205);
xnor U25013 (N_25013,N_21815,N_22697);
nand U25014 (N_25014,N_22768,N_22365);
nor U25015 (N_25015,N_23352,N_23452);
and U25016 (N_25016,N_23883,N_23394);
and U25017 (N_25017,N_22797,N_22086);
nand U25018 (N_25018,N_21768,N_21103);
nor U25019 (N_25019,N_22694,N_21794);
and U25020 (N_25020,N_21863,N_22744);
and U25021 (N_25021,N_22778,N_22598);
and U25022 (N_25022,N_22693,N_23587);
xnor U25023 (N_25023,N_21918,N_21283);
nor U25024 (N_25024,N_23548,N_23937);
nand U25025 (N_25025,N_21274,N_22257);
nor U25026 (N_25026,N_23640,N_23340);
nor U25027 (N_25027,N_21063,N_21132);
nor U25028 (N_25028,N_21585,N_23706);
or U25029 (N_25029,N_23086,N_21409);
and U25030 (N_25030,N_22796,N_22377);
and U25031 (N_25031,N_23714,N_21465);
xnor U25032 (N_25032,N_22298,N_21420);
or U25033 (N_25033,N_22799,N_21442);
xnor U25034 (N_25034,N_22003,N_21448);
nor U25035 (N_25035,N_22851,N_23828);
or U25036 (N_25036,N_21400,N_22226);
or U25037 (N_25037,N_22122,N_21560);
xnor U25038 (N_25038,N_21289,N_21519);
xnor U25039 (N_25039,N_22132,N_22311);
nor U25040 (N_25040,N_21982,N_22006);
nand U25041 (N_25041,N_23471,N_23033);
nor U25042 (N_25042,N_21666,N_22719);
xor U25043 (N_25043,N_23130,N_22765);
nor U25044 (N_25044,N_23043,N_23010);
and U25045 (N_25045,N_23945,N_21312);
nand U25046 (N_25046,N_22275,N_23970);
nand U25047 (N_25047,N_23567,N_21867);
nor U25048 (N_25048,N_22865,N_22601);
and U25049 (N_25049,N_23511,N_23474);
or U25050 (N_25050,N_22706,N_21927);
xor U25051 (N_25051,N_22133,N_21440);
or U25052 (N_25052,N_23886,N_23437);
nand U25053 (N_25053,N_23292,N_21845);
nor U25054 (N_25054,N_22304,N_22030);
and U25055 (N_25055,N_23950,N_22932);
xor U25056 (N_25056,N_23235,N_22341);
xnor U25057 (N_25057,N_22844,N_23609);
xor U25058 (N_25058,N_23866,N_22169);
nand U25059 (N_25059,N_23584,N_22819);
nand U25060 (N_25060,N_22194,N_21088);
xor U25061 (N_25061,N_23180,N_23002);
xnor U25062 (N_25062,N_22216,N_22329);
nor U25063 (N_25063,N_22880,N_21340);
xnor U25064 (N_25064,N_21013,N_23962);
nand U25065 (N_25065,N_21366,N_23113);
nor U25066 (N_25066,N_23649,N_22551);
nand U25067 (N_25067,N_22709,N_23228);
nor U25068 (N_25068,N_21734,N_21356);
or U25069 (N_25069,N_22162,N_21164);
nand U25070 (N_25070,N_23579,N_23760);
nand U25071 (N_25071,N_21844,N_23869);
and U25072 (N_25072,N_21437,N_21533);
nor U25073 (N_25073,N_21601,N_23664);
nand U25074 (N_25074,N_22215,N_22726);
and U25075 (N_25075,N_23001,N_23441);
xor U25076 (N_25076,N_22070,N_22586);
nor U25077 (N_25077,N_21690,N_23107);
nor U25078 (N_25078,N_22513,N_23977);
nor U25079 (N_25079,N_23789,N_22700);
nor U25080 (N_25080,N_22350,N_22542);
and U25081 (N_25081,N_22528,N_21419);
or U25082 (N_25082,N_23295,N_23289);
nand U25083 (N_25083,N_22913,N_21760);
nand U25084 (N_25084,N_23157,N_22129);
or U25085 (N_25085,N_22035,N_21009);
nor U25086 (N_25086,N_23022,N_21377);
nor U25087 (N_25087,N_21541,N_22952);
and U25088 (N_25088,N_23896,N_22556);
and U25089 (N_25089,N_22600,N_22338);
xnor U25090 (N_25090,N_21772,N_22181);
or U25091 (N_25091,N_23960,N_21034);
or U25092 (N_25092,N_21348,N_23659);
and U25093 (N_25093,N_21932,N_23595);
nand U25094 (N_25094,N_21452,N_22784);
nor U25095 (N_25095,N_22946,N_21453);
xor U25096 (N_25096,N_23480,N_21408);
and U25097 (N_25097,N_21946,N_22291);
and U25098 (N_25098,N_21620,N_22619);
and U25099 (N_25099,N_22444,N_22326);
or U25100 (N_25100,N_22385,N_23095);
nand U25101 (N_25101,N_23208,N_22904);
nor U25102 (N_25102,N_22312,N_22374);
nor U25103 (N_25103,N_23444,N_22618);
nor U25104 (N_25104,N_23371,N_22400);
nor U25105 (N_25105,N_21339,N_23004);
nand U25106 (N_25106,N_23749,N_23307);
nor U25107 (N_25107,N_21459,N_23047);
nor U25108 (N_25108,N_21049,N_21894);
and U25109 (N_25109,N_21216,N_21608);
nor U25110 (N_25110,N_23516,N_22649);
nor U25111 (N_25111,N_23650,N_23988);
or U25112 (N_25112,N_21641,N_21295);
or U25113 (N_25113,N_23720,N_21763);
nor U25114 (N_25114,N_22013,N_22029);
or U25115 (N_25115,N_21273,N_22454);
nor U25116 (N_25116,N_21198,N_21337);
nor U25117 (N_25117,N_21109,N_22847);
and U25118 (N_25118,N_23563,N_21576);
nor U25119 (N_25119,N_23865,N_22382);
and U25120 (N_25120,N_21125,N_21183);
xor U25121 (N_25121,N_22862,N_23448);
and U25122 (N_25122,N_22543,N_23053);
or U25123 (N_25123,N_23963,N_21730);
xor U25124 (N_25124,N_23055,N_23170);
or U25125 (N_25125,N_23034,N_21199);
nand U25126 (N_25126,N_22228,N_21042);
nand U25127 (N_25127,N_21901,N_22853);
or U25128 (N_25128,N_23495,N_22310);
nor U25129 (N_25129,N_22252,N_23076);
xor U25130 (N_25130,N_22868,N_23719);
xnor U25131 (N_25131,N_22225,N_23347);
or U25132 (N_25132,N_23739,N_21694);
xnor U25133 (N_25133,N_22213,N_23253);
nand U25134 (N_25134,N_22534,N_23255);
and U25135 (N_25135,N_21563,N_21401);
and U25136 (N_25136,N_22453,N_23190);
nand U25137 (N_25137,N_22127,N_23126);
xnor U25138 (N_25138,N_22773,N_23246);
nor U25139 (N_25139,N_22781,N_23670);
nand U25140 (N_25140,N_23611,N_21572);
nand U25141 (N_25141,N_23969,N_21015);
nand U25142 (N_25142,N_21373,N_21038);
xor U25143 (N_25143,N_21735,N_22265);
nand U25144 (N_25144,N_22370,N_22007);
and U25145 (N_25145,N_23166,N_21904);
xnor U25146 (N_25146,N_23200,N_23188);
nand U25147 (N_25147,N_23629,N_21956);
xor U25148 (N_25148,N_22079,N_22314);
xnor U25149 (N_25149,N_22995,N_21569);
nand U25150 (N_25150,N_22424,N_22963);
or U25151 (N_25151,N_23825,N_23890);
and U25152 (N_25152,N_23272,N_23986);
nor U25153 (N_25153,N_22205,N_22920);
xor U25154 (N_25154,N_23155,N_21721);
xnor U25155 (N_25155,N_21759,N_21215);
and U25156 (N_25156,N_21111,N_21778);
or U25157 (N_25157,N_22427,N_23796);
xor U25158 (N_25158,N_23122,N_23257);
nor U25159 (N_25159,N_21398,N_22993);
or U25160 (N_25160,N_21196,N_22103);
nor U25161 (N_25161,N_23161,N_22434);
and U25162 (N_25162,N_22752,N_23582);
or U25163 (N_25163,N_22173,N_23996);
xor U25164 (N_25164,N_22973,N_21358);
nor U25165 (N_25165,N_21937,N_22419);
nor U25166 (N_25166,N_21046,N_21707);
xor U25167 (N_25167,N_21719,N_23187);
or U25168 (N_25168,N_23223,N_21368);
nor U25169 (N_25169,N_23682,N_22807);
and U25170 (N_25170,N_22441,N_21910);
nand U25171 (N_25171,N_21854,N_23949);
nor U25172 (N_25172,N_21291,N_22816);
nand U25173 (N_25173,N_23206,N_22321);
nor U25174 (N_25174,N_22489,N_22565);
nand U25175 (N_25175,N_22412,N_23832);
nor U25176 (N_25176,N_23604,N_21061);
or U25177 (N_25177,N_23438,N_22643);
xor U25178 (N_25178,N_23026,N_21590);
nand U25179 (N_25179,N_22165,N_22155);
xnor U25180 (N_25180,N_21129,N_21654);
nand U25181 (N_25181,N_22152,N_22715);
xor U25182 (N_25182,N_21786,N_21540);
nand U25183 (N_25183,N_22585,N_23230);
and U25184 (N_25184,N_23374,N_21984);
nor U25185 (N_25185,N_22916,N_21928);
nand U25186 (N_25186,N_21843,N_21287);
nor U25187 (N_25187,N_21673,N_21135);
and U25188 (N_25188,N_21357,N_22016);
or U25189 (N_25189,N_22047,N_23531);
or U25190 (N_25190,N_22332,N_21496);
xnor U25191 (N_25191,N_22955,N_22237);
xnor U25192 (N_25192,N_23240,N_23879);
nand U25193 (N_25193,N_22686,N_21231);
or U25194 (N_25194,N_22516,N_23489);
nor U25195 (N_25195,N_23500,N_23955);
or U25196 (N_25196,N_23888,N_23899);
and U25197 (N_25197,N_23282,N_21973);
or U25198 (N_25198,N_21479,N_22999);
or U25199 (N_25199,N_21598,N_21935);
nand U25200 (N_25200,N_21309,N_21636);
and U25201 (N_25201,N_22183,N_22190);
xor U25202 (N_25202,N_22682,N_22414);
nor U25203 (N_25203,N_23887,N_22315);
nor U25204 (N_25204,N_21461,N_21018);
nor U25205 (N_25205,N_23290,N_22171);
and U25206 (N_25206,N_21971,N_22823);
and U25207 (N_25207,N_21065,N_23515);
and U25208 (N_25208,N_21145,N_23067);
xor U25209 (N_25209,N_21140,N_21770);
or U25210 (N_25210,N_23774,N_21957);
nand U25211 (N_25211,N_22189,N_22825);
xor U25212 (N_25212,N_21923,N_22403);
xor U25213 (N_25213,N_22267,N_23839);
xor U25214 (N_25214,N_22330,N_23209);
or U25215 (N_25215,N_21703,N_21036);
nand U25216 (N_25216,N_21687,N_23245);
nor U25217 (N_25217,N_21816,N_23560);
nor U25218 (N_25218,N_23449,N_22254);
nor U25219 (N_25219,N_21351,N_23141);
nand U25220 (N_25220,N_21166,N_21426);
nor U25221 (N_25221,N_23456,N_23423);
xor U25222 (N_25222,N_23083,N_23702);
and U25223 (N_25223,N_23931,N_22574);
or U25224 (N_25224,N_22717,N_23408);
nor U25225 (N_25225,N_22394,N_23013);
nor U25226 (N_25226,N_21050,N_21107);
nand U25227 (N_25227,N_21407,N_22743);
nor U25228 (N_25228,N_22085,N_21552);
nor U25229 (N_25229,N_22297,N_21542);
xnor U25230 (N_25230,N_21612,N_22895);
and U25231 (N_25231,N_22143,N_21817);
or U25232 (N_25232,N_23674,N_23267);
nand U25233 (N_25233,N_23797,N_22164);
nand U25234 (N_25234,N_23131,N_23351);
nor U25235 (N_25235,N_21234,N_21847);
or U25236 (N_25236,N_22931,N_21127);
xnor U25237 (N_25237,N_23527,N_23510);
nor U25238 (N_25238,N_23475,N_21581);
nand U25239 (N_25239,N_22555,N_22623);
xor U25240 (N_25240,N_22866,N_22025);
and U25241 (N_25241,N_21529,N_22418);
or U25242 (N_25242,N_23734,N_22506);
or U25243 (N_25243,N_22742,N_21976);
and U25244 (N_25244,N_23274,N_21920);
nor U25245 (N_25245,N_21245,N_22024);
xor U25246 (N_25246,N_21069,N_23598);
nor U25247 (N_25247,N_22115,N_21027);
nand U25248 (N_25248,N_22761,N_21940);
nor U25249 (N_25249,N_23380,N_23411);
nor U25250 (N_25250,N_22399,N_23599);
nor U25251 (N_25251,N_23800,N_21221);
or U25252 (N_25252,N_22269,N_22015);
and U25253 (N_25253,N_23983,N_22970);
or U25254 (N_25254,N_23334,N_21099);
or U25255 (N_25255,N_23136,N_22926);
or U25256 (N_25256,N_21445,N_22760);
and U25257 (N_25257,N_23238,N_22548);
xnor U25258 (N_25258,N_23539,N_22058);
nand U25259 (N_25259,N_21117,N_22642);
and U25260 (N_25260,N_22469,N_22222);
xnor U25261 (N_25261,N_23454,N_23762);
nand U25262 (N_25262,N_21838,N_21264);
nand U25263 (N_25263,N_22629,N_21020);
and U25264 (N_25264,N_21537,N_21792);
and U25265 (N_25265,N_21249,N_22950);
xor U25266 (N_25266,N_22055,N_21399);
nand U25267 (N_25267,N_21680,N_21929);
nand U25268 (N_25268,N_23925,N_23140);
nor U25269 (N_25269,N_21397,N_21509);
nand U25270 (N_25270,N_22465,N_23498);
xnor U25271 (N_25271,N_21568,N_23496);
and U25272 (N_25272,N_22962,N_23269);
nand U25273 (N_25273,N_22212,N_21260);
nand U25274 (N_25274,N_22028,N_22186);
xnor U25275 (N_25275,N_23771,N_21235);
xor U25276 (N_25276,N_23645,N_23015);
nand U25277 (N_25277,N_23947,N_22640);
nor U25278 (N_25278,N_23630,N_21808);
nor U25279 (N_25279,N_22347,N_23728);
nand U25280 (N_25280,N_22820,N_22428);
nand U25281 (N_25281,N_22307,N_23908);
nand U25282 (N_25282,N_21209,N_23946);
nand U25283 (N_25283,N_23958,N_21148);
nor U25284 (N_25284,N_23612,N_23692);
and U25285 (N_25285,N_23387,N_22791);
xnor U25286 (N_25286,N_23605,N_21098);
nand U25287 (N_25287,N_21738,N_22217);
nor U25288 (N_25288,N_21706,N_23167);
or U25289 (N_25289,N_23809,N_22049);
or U25290 (N_25290,N_21708,N_23795);
xor U25291 (N_25291,N_22052,N_23922);
or U25292 (N_25292,N_21157,N_22511);
and U25293 (N_25293,N_23204,N_22705);
nand U25294 (N_25294,N_21396,N_21197);
or U25295 (N_25295,N_22504,N_21106);
or U25296 (N_25296,N_21561,N_22863);
or U25297 (N_25297,N_23270,N_22972);
and U25298 (N_25298,N_22378,N_22497);
or U25299 (N_25299,N_22097,N_22698);
nor U25300 (N_25300,N_23687,N_22587);
nor U25301 (N_25301,N_23652,N_21105);
nor U25302 (N_25302,N_22327,N_21336);
xnor U25303 (N_25303,N_22818,N_23573);
and U25304 (N_25304,N_23412,N_22872);
and U25305 (N_25305,N_22525,N_23111);
nor U25306 (N_25306,N_22714,N_22343);
xnor U25307 (N_25307,N_21416,N_23808);
or U25308 (N_25308,N_22570,N_23662);
nor U25309 (N_25309,N_22567,N_23637);
xnor U25310 (N_25310,N_23778,N_23973);
and U25311 (N_25311,N_21776,N_21139);
or U25312 (N_25312,N_21475,N_21931);
or U25313 (N_25313,N_23077,N_22358);
nand U25314 (N_25314,N_21970,N_21028);
nand U25315 (N_25315,N_21668,N_22789);
nor U25316 (N_25316,N_21045,N_23121);
nand U25317 (N_25317,N_22460,N_22716);
or U25318 (N_25318,N_23278,N_21538);
nand U25319 (N_25319,N_22767,N_23641);
and U25320 (N_25320,N_21347,N_21729);
xor U25321 (N_25321,N_22290,N_22854);
nor U25322 (N_25322,N_23990,N_21242);
or U25323 (N_25323,N_22219,N_22491);
and U25324 (N_25324,N_21210,N_22482);
nand U25325 (N_25325,N_21194,N_23331);
and U25326 (N_25326,N_22324,N_23402);
xnor U25327 (N_25327,N_21188,N_21190);
nor U25328 (N_25328,N_23451,N_23565);
nand U25329 (N_25329,N_23381,N_23738);
xor U25330 (N_25330,N_23164,N_21263);
xnor U25331 (N_25331,N_21866,N_23273);
nor U25332 (N_25332,N_22492,N_21010);
nand U25333 (N_25333,N_23242,N_21483);
and U25334 (N_25334,N_21275,N_21214);
nand U25335 (N_25335,N_23310,N_23450);
nor U25336 (N_25336,N_23713,N_21554);
nor U25337 (N_25337,N_23291,N_23089);
xnor U25338 (N_25338,N_21267,N_23576);
xor U25339 (N_25339,N_23732,N_22902);
nand U25340 (N_25340,N_23779,N_21914);
nor U25341 (N_25341,N_22309,N_23716);
and U25342 (N_25342,N_21544,N_22740);
and U25343 (N_25343,N_23218,N_21648);
or U25344 (N_25344,N_22306,N_23954);
or U25345 (N_25345,N_23676,N_23608);
and U25346 (N_25346,N_23905,N_23309);
nand U25347 (N_25347,N_22468,N_23619);
xor U25348 (N_25348,N_23436,N_22101);
nand U25349 (N_25349,N_21549,N_22184);
xnor U25350 (N_25350,N_21288,N_23469);
nand U25351 (N_25351,N_21371,N_22336);
and U25352 (N_25352,N_21325,N_21217);
nor U25353 (N_25353,N_22153,N_23181);
or U25354 (N_25354,N_23486,N_23252);
and U25355 (N_25355,N_23615,N_23174);
nand U25356 (N_25356,N_23360,N_22195);
nor U25357 (N_25357,N_23303,N_23144);
xor U25358 (N_25358,N_23244,N_21286);
nor U25359 (N_25359,N_22266,N_22933);
xor U25360 (N_25360,N_23512,N_23910);
nand U25361 (N_25361,N_23927,N_22836);
nor U25362 (N_25362,N_21722,N_22406);
nand U25363 (N_25363,N_23112,N_23405);
xnor U25364 (N_25364,N_21372,N_22537);
nand U25365 (N_25365,N_21945,N_21185);
nor U25366 (N_25366,N_22659,N_21243);
xnor U25367 (N_25367,N_21876,N_21990);
nand U25368 (N_25368,N_21657,N_23414);
or U25369 (N_25369,N_23397,N_23895);
or U25370 (N_25370,N_22790,N_23305);
nor U25371 (N_25371,N_23275,N_22667);
nor U25372 (N_25372,N_22459,N_21835);
nor U25373 (N_25373,N_23538,N_23882);
nand U25374 (N_25374,N_22808,N_21270);
nand U25375 (N_25375,N_23390,N_22603);
nor U25376 (N_25376,N_21062,N_23904);
nand U25377 (N_25377,N_21745,N_21960);
and U25378 (N_25378,N_22583,N_21596);
xor U25379 (N_25379,N_22533,N_23403);
nand U25380 (N_25380,N_21101,N_22018);
nand U25381 (N_25381,N_22837,N_21256);
and U25382 (N_25382,N_23924,N_23487);
nand U25383 (N_25383,N_21810,N_22650);
nand U25384 (N_25384,N_22375,N_22048);
nor U25385 (N_25385,N_21454,N_23056);
nand U25386 (N_25386,N_22289,N_23094);
or U25387 (N_25387,N_21811,N_21328);
nor U25388 (N_25388,N_22518,N_21825);
nor U25389 (N_25389,N_23000,N_23864);
and U25390 (N_25390,N_21642,N_22410);
nor U25391 (N_25391,N_22069,N_23231);
and U25392 (N_25392,N_21501,N_22032);
nor U25393 (N_25393,N_21523,N_22134);
xor U25394 (N_25394,N_23683,N_23948);
nand U25395 (N_25395,N_22135,N_21237);
nor U25396 (N_25396,N_21030,N_22449);
nand U25397 (N_25397,N_23819,N_21506);
and U25398 (N_25398,N_22687,N_22393);
or U25399 (N_25399,N_22850,N_23189);
nand U25400 (N_25400,N_23944,N_22182);
nor U25401 (N_25401,N_23623,N_21133);
nor U25402 (N_25402,N_21686,N_22197);
nor U25403 (N_25403,N_23532,N_21206);
or U25404 (N_25404,N_21265,N_21890);
nor U25405 (N_25405,N_23831,N_22840);
nand U25406 (N_25406,N_21860,N_23445);
and U25407 (N_25407,N_22193,N_22708);
and U25408 (N_25408,N_21919,N_23930);
and U25409 (N_25409,N_23834,N_23173);
nor U25410 (N_25410,N_22856,N_23145);
nor U25411 (N_25411,N_23193,N_23901);
or U25412 (N_25412,N_22462,N_22417);
nand U25413 (N_25413,N_22415,N_22093);
or U25414 (N_25414,N_22792,N_21742);
xnor U25415 (N_25415,N_22026,N_23626);
and U25416 (N_25416,N_21390,N_23801);
xor U25417 (N_25417,N_21842,N_21864);
xnor U25418 (N_25418,N_23658,N_21619);
and U25419 (N_25419,N_22890,N_21386);
xor U25420 (N_25420,N_23667,N_22475);
nand U25421 (N_25421,N_21925,N_23163);
xnor U25422 (N_25422,N_22685,N_23074);
or U25423 (N_25423,N_22900,N_22354);
and U25424 (N_25424,N_21056,N_21247);
xnor U25425 (N_25425,N_23433,N_22769);
nand U25426 (N_25426,N_22956,N_23264);
or U25427 (N_25427,N_23666,N_23159);
nor U25428 (N_25428,N_21429,N_21480);
nor U25429 (N_25429,N_23773,N_22696);
xnor U25430 (N_25430,N_22174,N_22198);
and U25431 (N_25431,N_23183,N_23518);
nor U25432 (N_25432,N_21179,N_21944);
nor U25433 (N_25433,N_22757,N_23019);
nand U25434 (N_25434,N_23298,N_23859);
and U25435 (N_25435,N_22723,N_22622);
xor U25436 (N_25436,N_23169,N_23409);
xor U25437 (N_25437,N_21114,N_21913);
nand U25438 (N_25438,N_23481,N_23179);
and U25439 (N_25439,N_21674,N_22178);
xor U25440 (N_25440,N_21993,N_21395);
nor U25441 (N_25441,N_21226,N_22857);
nand U25442 (N_25442,N_22912,N_23991);
or U25443 (N_25443,N_23388,N_23018);
xor U25444 (N_25444,N_22559,N_23704);
xor U25445 (N_25445,N_22817,N_21610);
nor U25446 (N_25446,N_22202,N_22067);
and U25447 (N_25447,N_23234,N_21170);
nor U25448 (N_25448,N_23030,N_22123);
nor U25449 (N_25449,N_22094,N_22114);
nor U25450 (N_25450,N_21008,N_22148);
or U25451 (N_25451,N_21614,N_21052);
xnor U25452 (N_25452,N_22911,N_21387);
nor U25453 (N_25453,N_22294,N_23085);
or U25454 (N_25454,N_22522,N_23621);
and U25455 (N_25455,N_21965,N_22464);
or U25456 (N_25456,N_21765,N_21463);
nor U25457 (N_25457,N_21751,N_23997);
or U25458 (N_25458,N_21470,N_21952);
nand U25459 (N_25459,N_21156,N_22979);
nor U25460 (N_25460,N_21182,N_23256);
xor U25461 (N_25461,N_21986,N_23386);
nand U25462 (N_25462,N_22605,N_23712);
nor U25463 (N_25463,N_23499,N_21987);
nand U25464 (N_25464,N_21364,N_22919);
and U25465 (N_25465,N_21600,N_22220);
nor U25466 (N_25466,N_23764,N_22683);
and U25467 (N_25467,N_21344,N_21248);
xnor U25468 (N_25468,N_23999,N_22755);
and U25469 (N_25469,N_22608,N_22677);
xor U25470 (N_25470,N_21627,N_21532);
and U25471 (N_25471,N_21308,N_21029);
nor U25472 (N_25472,N_23251,N_21489);
xnor U25473 (N_25473,N_23478,N_22675);
nor U25474 (N_25474,N_21681,N_22722);
and U25475 (N_25475,N_21821,N_22196);
nor U25476 (N_25476,N_21057,N_21414);
xor U25477 (N_25477,N_23092,N_23593);
or U25478 (N_25478,N_22436,N_23338);
xnor U25479 (N_25479,N_21481,N_22575);
nor U25480 (N_25480,N_22867,N_23753);
or U25481 (N_25481,N_21219,N_22017);
and U25482 (N_25482,N_21670,N_23545);
xor U25483 (N_25483,N_21511,N_21752);
or U25484 (N_25484,N_23399,N_22088);
or U25485 (N_25485,N_23343,N_21522);
or U25486 (N_25486,N_21813,N_21003);
xor U25487 (N_25487,N_23457,N_23348);
and U25488 (N_25488,N_22523,N_23485);
xnor U25489 (N_25489,N_22554,N_21704);
nand U25490 (N_25490,N_23096,N_23241);
xnor U25491 (N_25491,N_23978,N_22852);
nand U25492 (N_25492,N_23293,N_23435);
and U25493 (N_25493,N_23672,N_21499);
or U25494 (N_25494,N_21895,N_21238);
or U25495 (N_25495,N_22647,N_22985);
nor U25496 (N_25496,N_21659,N_21624);
xnor U25497 (N_25497,N_21507,N_21469);
nand U25498 (N_25498,N_21118,N_23064);
nand U25499 (N_25499,N_23446,N_23359);
and U25500 (N_25500,N_23853,N_21631);
nand U25501 (N_25501,N_21822,N_22407);
or U25502 (N_25502,N_22450,N_21946);
nand U25503 (N_25503,N_23283,N_23417);
nand U25504 (N_25504,N_21666,N_23635);
or U25505 (N_25505,N_23010,N_22174);
or U25506 (N_25506,N_22378,N_21678);
nand U25507 (N_25507,N_22048,N_21289);
nand U25508 (N_25508,N_22024,N_23138);
xor U25509 (N_25509,N_23334,N_23549);
or U25510 (N_25510,N_22101,N_23488);
xor U25511 (N_25511,N_23556,N_21385);
nand U25512 (N_25512,N_22448,N_21579);
nand U25513 (N_25513,N_22434,N_22752);
nor U25514 (N_25514,N_23810,N_23262);
nand U25515 (N_25515,N_22185,N_21650);
and U25516 (N_25516,N_23105,N_23865);
xnor U25517 (N_25517,N_21114,N_21222);
and U25518 (N_25518,N_21877,N_22957);
xor U25519 (N_25519,N_21549,N_21444);
nand U25520 (N_25520,N_21910,N_23888);
nor U25521 (N_25521,N_23193,N_21335);
or U25522 (N_25522,N_22625,N_22784);
nor U25523 (N_25523,N_21922,N_23589);
and U25524 (N_25524,N_21304,N_22233);
and U25525 (N_25525,N_22386,N_21497);
nor U25526 (N_25526,N_22561,N_21855);
nor U25527 (N_25527,N_23074,N_23601);
and U25528 (N_25528,N_21866,N_22354);
xor U25529 (N_25529,N_21210,N_21632);
xor U25530 (N_25530,N_21082,N_21118);
nor U25531 (N_25531,N_21467,N_21253);
nand U25532 (N_25532,N_21629,N_23427);
nand U25533 (N_25533,N_22880,N_22064);
nor U25534 (N_25534,N_22341,N_22391);
nor U25535 (N_25535,N_22791,N_22810);
or U25536 (N_25536,N_22385,N_21212);
xor U25537 (N_25537,N_23198,N_22333);
nor U25538 (N_25538,N_22248,N_22442);
nor U25539 (N_25539,N_22958,N_21443);
and U25540 (N_25540,N_21370,N_23717);
nand U25541 (N_25541,N_21766,N_21062);
nand U25542 (N_25542,N_22232,N_23677);
nor U25543 (N_25543,N_22598,N_22379);
nor U25544 (N_25544,N_23080,N_23192);
xnor U25545 (N_25545,N_21471,N_21556);
nor U25546 (N_25546,N_22046,N_22090);
or U25547 (N_25547,N_23170,N_23571);
nand U25548 (N_25548,N_23817,N_22518);
nor U25549 (N_25549,N_23481,N_23207);
nor U25550 (N_25550,N_21091,N_23157);
xnor U25551 (N_25551,N_23219,N_21302);
and U25552 (N_25552,N_23043,N_23907);
nor U25553 (N_25553,N_23450,N_23720);
or U25554 (N_25554,N_21119,N_22196);
xnor U25555 (N_25555,N_21376,N_21531);
xor U25556 (N_25556,N_22496,N_23050);
or U25557 (N_25557,N_22672,N_22998);
nor U25558 (N_25558,N_22743,N_21871);
xnor U25559 (N_25559,N_23896,N_22244);
nand U25560 (N_25560,N_23795,N_23072);
or U25561 (N_25561,N_22082,N_21735);
xor U25562 (N_25562,N_21190,N_23058);
nand U25563 (N_25563,N_22476,N_23846);
xnor U25564 (N_25564,N_22793,N_23031);
nand U25565 (N_25565,N_23144,N_23899);
and U25566 (N_25566,N_22069,N_22639);
nand U25567 (N_25567,N_23119,N_23635);
or U25568 (N_25568,N_23208,N_21597);
nor U25569 (N_25569,N_22064,N_21379);
nor U25570 (N_25570,N_22776,N_22506);
or U25571 (N_25571,N_23776,N_23093);
or U25572 (N_25572,N_22016,N_21111);
or U25573 (N_25573,N_23593,N_22646);
or U25574 (N_25574,N_23261,N_22570);
nor U25575 (N_25575,N_21923,N_21694);
xnor U25576 (N_25576,N_23634,N_21764);
or U25577 (N_25577,N_21769,N_23192);
nor U25578 (N_25578,N_21335,N_23680);
or U25579 (N_25579,N_23748,N_21386);
and U25580 (N_25580,N_22920,N_23229);
xnor U25581 (N_25581,N_23056,N_23275);
xor U25582 (N_25582,N_23435,N_22233);
nor U25583 (N_25583,N_22444,N_22753);
nor U25584 (N_25584,N_21180,N_22916);
xnor U25585 (N_25585,N_23976,N_22158);
nand U25586 (N_25586,N_21179,N_23843);
nand U25587 (N_25587,N_23723,N_22749);
and U25588 (N_25588,N_22586,N_23899);
xnor U25589 (N_25589,N_23844,N_21987);
or U25590 (N_25590,N_22232,N_22081);
xnor U25591 (N_25591,N_21344,N_23077);
or U25592 (N_25592,N_22430,N_23915);
nand U25593 (N_25593,N_23297,N_21558);
nand U25594 (N_25594,N_23155,N_21502);
nor U25595 (N_25595,N_22023,N_22292);
nand U25596 (N_25596,N_22082,N_22770);
or U25597 (N_25597,N_23476,N_22249);
or U25598 (N_25598,N_22690,N_22887);
xor U25599 (N_25599,N_21724,N_22110);
nor U25600 (N_25600,N_21029,N_23074);
nand U25601 (N_25601,N_21722,N_22490);
and U25602 (N_25602,N_21569,N_21717);
nand U25603 (N_25603,N_23348,N_21454);
nand U25604 (N_25604,N_22609,N_22289);
or U25605 (N_25605,N_23270,N_23131);
nand U25606 (N_25606,N_22265,N_22726);
xor U25607 (N_25607,N_23171,N_22734);
nand U25608 (N_25608,N_23844,N_23131);
xor U25609 (N_25609,N_23365,N_23821);
nor U25610 (N_25610,N_21734,N_23747);
nand U25611 (N_25611,N_22566,N_22572);
or U25612 (N_25612,N_22740,N_21459);
nor U25613 (N_25613,N_22930,N_21371);
or U25614 (N_25614,N_23322,N_22981);
or U25615 (N_25615,N_23679,N_21076);
or U25616 (N_25616,N_23297,N_21148);
nor U25617 (N_25617,N_23136,N_22859);
nand U25618 (N_25618,N_23661,N_21223);
nor U25619 (N_25619,N_23987,N_21927);
xor U25620 (N_25620,N_23359,N_22718);
or U25621 (N_25621,N_22065,N_23569);
nand U25622 (N_25622,N_23994,N_23076);
nand U25623 (N_25623,N_23998,N_21051);
nand U25624 (N_25624,N_21622,N_21113);
and U25625 (N_25625,N_22202,N_23433);
nor U25626 (N_25626,N_22631,N_21647);
nand U25627 (N_25627,N_22442,N_22679);
or U25628 (N_25628,N_22100,N_22925);
xnor U25629 (N_25629,N_23875,N_23504);
and U25630 (N_25630,N_23863,N_23480);
nand U25631 (N_25631,N_22887,N_23395);
nor U25632 (N_25632,N_22873,N_23683);
or U25633 (N_25633,N_23465,N_23845);
or U25634 (N_25634,N_23880,N_21987);
or U25635 (N_25635,N_22611,N_21110);
nor U25636 (N_25636,N_23309,N_22119);
nand U25637 (N_25637,N_22216,N_22743);
nand U25638 (N_25638,N_23684,N_23120);
xor U25639 (N_25639,N_22875,N_22619);
nor U25640 (N_25640,N_21805,N_22126);
xor U25641 (N_25641,N_22836,N_22458);
nand U25642 (N_25642,N_21454,N_23506);
nand U25643 (N_25643,N_23322,N_21094);
nor U25644 (N_25644,N_22754,N_23771);
nand U25645 (N_25645,N_21151,N_21228);
or U25646 (N_25646,N_21484,N_21755);
xor U25647 (N_25647,N_23201,N_23043);
nor U25648 (N_25648,N_21401,N_21067);
nor U25649 (N_25649,N_23059,N_23201);
or U25650 (N_25650,N_22141,N_23919);
nand U25651 (N_25651,N_23076,N_22632);
and U25652 (N_25652,N_22474,N_22468);
or U25653 (N_25653,N_22998,N_22478);
and U25654 (N_25654,N_21350,N_23633);
xnor U25655 (N_25655,N_22253,N_21338);
nand U25656 (N_25656,N_22391,N_21672);
xnor U25657 (N_25657,N_23384,N_22432);
nand U25658 (N_25658,N_21913,N_23499);
and U25659 (N_25659,N_22341,N_21079);
xnor U25660 (N_25660,N_23539,N_22664);
or U25661 (N_25661,N_22728,N_21364);
or U25662 (N_25662,N_21220,N_23688);
or U25663 (N_25663,N_23101,N_21015);
xnor U25664 (N_25664,N_22410,N_22986);
nor U25665 (N_25665,N_22701,N_22912);
nand U25666 (N_25666,N_21211,N_23079);
nand U25667 (N_25667,N_21302,N_22479);
and U25668 (N_25668,N_23949,N_23290);
xnor U25669 (N_25669,N_23461,N_22882);
or U25670 (N_25670,N_23417,N_23528);
nand U25671 (N_25671,N_22606,N_23211);
nand U25672 (N_25672,N_21474,N_22891);
xnor U25673 (N_25673,N_23609,N_22124);
nand U25674 (N_25674,N_22910,N_21674);
nor U25675 (N_25675,N_23355,N_21814);
or U25676 (N_25676,N_21883,N_22275);
nand U25677 (N_25677,N_23203,N_21162);
xnor U25678 (N_25678,N_23495,N_21009);
or U25679 (N_25679,N_21237,N_23977);
nand U25680 (N_25680,N_23556,N_23957);
nand U25681 (N_25681,N_23475,N_23075);
nor U25682 (N_25682,N_21980,N_23078);
xor U25683 (N_25683,N_21475,N_22437);
or U25684 (N_25684,N_22453,N_23950);
xor U25685 (N_25685,N_22380,N_23158);
nor U25686 (N_25686,N_21003,N_22912);
xnor U25687 (N_25687,N_22990,N_21368);
nor U25688 (N_25688,N_23051,N_21368);
or U25689 (N_25689,N_22039,N_22806);
or U25690 (N_25690,N_21339,N_22253);
xor U25691 (N_25691,N_23036,N_23432);
nor U25692 (N_25692,N_22755,N_22920);
and U25693 (N_25693,N_23742,N_23434);
nand U25694 (N_25694,N_22248,N_21922);
nand U25695 (N_25695,N_21185,N_21390);
and U25696 (N_25696,N_22393,N_23370);
and U25697 (N_25697,N_23620,N_23406);
nor U25698 (N_25698,N_22800,N_23272);
nor U25699 (N_25699,N_23416,N_21882);
nand U25700 (N_25700,N_22688,N_21576);
or U25701 (N_25701,N_22191,N_21447);
xnor U25702 (N_25702,N_22275,N_21361);
or U25703 (N_25703,N_21919,N_21400);
and U25704 (N_25704,N_22580,N_22972);
and U25705 (N_25705,N_23250,N_21772);
nand U25706 (N_25706,N_21431,N_21873);
xnor U25707 (N_25707,N_22072,N_21747);
or U25708 (N_25708,N_22595,N_23453);
xor U25709 (N_25709,N_23586,N_22192);
and U25710 (N_25710,N_21446,N_22540);
nand U25711 (N_25711,N_23598,N_23220);
nand U25712 (N_25712,N_23021,N_21951);
xnor U25713 (N_25713,N_21946,N_21739);
nor U25714 (N_25714,N_22332,N_21057);
nor U25715 (N_25715,N_21890,N_23158);
xor U25716 (N_25716,N_21088,N_21237);
and U25717 (N_25717,N_23823,N_21645);
nand U25718 (N_25718,N_22727,N_22431);
and U25719 (N_25719,N_21036,N_22605);
or U25720 (N_25720,N_21269,N_21383);
xor U25721 (N_25721,N_21254,N_23436);
or U25722 (N_25722,N_21077,N_23500);
xnor U25723 (N_25723,N_22392,N_22789);
nand U25724 (N_25724,N_23818,N_23824);
and U25725 (N_25725,N_23262,N_23745);
xor U25726 (N_25726,N_23939,N_23927);
and U25727 (N_25727,N_22993,N_22169);
xnor U25728 (N_25728,N_21584,N_22784);
nand U25729 (N_25729,N_23311,N_22199);
nand U25730 (N_25730,N_21918,N_22834);
nand U25731 (N_25731,N_23492,N_22772);
nand U25732 (N_25732,N_22566,N_21521);
and U25733 (N_25733,N_21743,N_22102);
or U25734 (N_25734,N_22191,N_21522);
nand U25735 (N_25735,N_23135,N_22395);
xor U25736 (N_25736,N_21242,N_23582);
nand U25737 (N_25737,N_22121,N_23820);
nor U25738 (N_25738,N_23140,N_23349);
or U25739 (N_25739,N_23648,N_23944);
and U25740 (N_25740,N_23601,N_21994);
and U25741 (N_25741,N_21107,N_23248);
nand U25742 (N_25742,N_21121,N_22829);
and U25743 (N_25743,N_23957,N_23237);
or U25744 (N_25744,N_22834,N_21728);
xor U25745 (N_25745,N_22308,N_22180);
nor U25746 (N_25746,N_23538,N_21547);
or U25747 (N_25747,N_22068,N_21509);
or U25748 (N_25748,N_21256,N_22901);
nor U25749 (N_25749,N_23372,N_22335);
and U25750 (N_25750,N_22977,N_23544);
nor U25751 (N_25751,N_22754,N_22574);
xor U25752 (N_25752,N_23994,N_23609);
and U25753 (N_25753,N_23748,N_23110);
or U25754 (N_25754,N_23037,N_21187);
and U25755 (N_25755,N_21820,N_22872);
nor U25756 (N_25756,N_21003,N_22462);
and U25757 (N_25757,N_22158,N_22446);
and U25758 (N_25758,N_21178,N_23227);
nor U25759 (N_25759,N_21582,N_22488);
nor U25760 (N_25760,N_22425,N_21558);
nor U25761 (N_25761,N_21148,N_23126);
nor U25762 (N_25762,N_22449,N_22035);
xor U25763 (N_25763,N_22375,N_22320);
nand U25764 (N_25764,N_23502,N_22961);
and U25765 (N_25765,N_23023,N_23829);
and U25766 (N_25766,N_22676,N_21995);
nor U25767 (N_25767,N_23362,N_21796);
nand U25768 (N_25768,N_21086,N_21912);
and U25769 (N_25769,N_23350,N_23979);
nand U25770 (N_25770,N_21086,N_23839);
xor U25771 (N_25771,N_21504,N_23765);
and U25772 (N_25772,N_23377,N_23456);
xnor U25773 (N_25773,N_22087,N_21148);
xor U25774 (N_25774,N_22635,N_23527);
nor U25775 (N_25775,N_22945,N_21637);
and U25776 (N_25776,N_22310,N_21262);
xor U25777 (N_25777,N_22949,N_22985);
nor U25778 (N_25778,N_21907,N_23600);
nand U25779 (N_25779,N_23615,N_21807);
xnor U25780 (N_25780,N_23197,N_23541);
and U25781 (N_25781,N_22453,N_21153);
nor U25782 (N_25782,N_21459,N_22612);
nor U25783 (N_25783,N_21062,N_22390);
nor U25784 (N_25784,N_22152,N_23954);
xor U25785 (N_25785,N_22280,N_21816);
xor U25786 (N_25786,N_22815,N_23446);
and U25787 (N_25787,N_23710,N_23740);
nor U25788 (N_25788,N_21978,N_23580);
or U25789 (N_25789,N_23974,N_23102);
and U25790 (N_25790,N_21741,N_21279);
or U25791 (N_25791,N_23166,N_21439);
nand U25792 (N_25792,N_21270,N_22260);
nand U25793 (N_25793,N_22523,N_22746);
and U25794 (N_25794,N_23732,N_21055);
nor U25795 (N_25795,N_23365,N_21018);
xnor U25796 (N_25796,N_23690,N_21587);
and U25797 (N_25797,N_21572,N_23028);
nor U25798 (N_25798,N_23793,N_23846);
xor U25799 (N_25799,N_23706,N_23331);
or U25800 (N_25800,N_21326,N_22505);
nand U25801 (N_25801,N_22081,N_23911);
or U25802 (N_25802,N_21576,N_22380);
and U25803 (N_25803,N_21878,N_21792);
and U25804 (N_25804,N_23980,N_23664);
nor U25805 (N_25805,N_22678,N_23142);
nand U25806 (N_25806,N_21038,N_21388);
or U25807 (N_25807,N_23756,N_22903);
and U25808 (N_25808,N_23385,N_21545);
or U25809 (N_25809,N_21616,N_21988);
and U25810 (N_25810,N_23849,N_22990);
and U25811 (N_25811,N_23589,N_23501);
nand U25812 (N_25812,N_22376,N_23213);
or U25813 (N_25813,N_22614,N_23914);
xor U25814 (N_25814,N_22639,N_23777);
nand U25815 (N_25815,N_22873,N_21014);
and U25816 (N_25816,N_22311,N_23248);
nor U25817 (N_25817,N_22952,N_21418);
nor U25818 (N_25818,N_22851,N_21878);
and U25819 (N_25819,N_22973,N_23104);
nor U25820 (N_25820,N_23302,N_23036);
nand U25821 (N_25821,N_23906,N_23818);
and U25822 (N_25822,N_22131,N_21838);
nor U25823 (N_25823,N_23776,N_23500);
nand U25824 (N_25824,N_22329,N_22809);
nor U25825 (N_25825,N_21072,N_23981);
nand U25826 (N_25826,N_23668,N_22437);
xor U25827 (N_25827,N_22235,N_21127);
and U25828 (N_25828,N_23353,N_21875);
and U25829 (N_25829,N_22699,N_22483);
nor U25830 (N_25830,N_21092,N_21554);
nand U25831 (N_25831,N_21871,N_21762);
xor U25832 (N_25832,N_22234,N_21979);
and U25833 (N_25833,N_22286,N_23725);
nand U25834 (N_25834,N_21524,N_21719);
nor U25835 (N_25835,N_21397,N_21818);
and U25836 (N_25836,N_23307,N_22943);
or U25837 (N_25837,N_22956,N_21993);
nor U25838 (N_25838,N_21236,N_21525);
xor U25839 (N_25839,N_22101,N_21865);
and U25840 (N_25840,N_21093,N_22458);
or U25841 (N_25841,N_22295,N_21168);
nor U25842 (N_25842,N_21430,N_22864);
or U25843 (N_25843,N_21123,N_21890);
xor U25844 (N_25844,N_23636,N_21683);
xor U25845 (N_25845,N_23096,N_23923);
nand U25846 (N_25846,N_22250,N_22409);
nor U25847 (N_25847,N_23402,N_22048);
nand U25848 (N_25848,N_22541,N_23019);
nor U25849 (N_25849,N_21309,N_22958);
nor U25850 (N_25850,N_23019,N_22179);
nor U25851 (N_25851,N_22591,N_21794);
nor U25852 (N_25852,N_23486,N_23012);
and U25853 (N_25853,N_22189,N_22663);
and U25854 (N_25854,N_23650,N_22146);
or U25855 (N_25855,N_23055,N_21447);
and U25856 (N_25856,N_21382,N_21025);
or U25857 (N_25857,N_21001,N_23297);
and U25858 (N_25858,N_22397,N_23493);
or U25859 (N_25859,N_21582,N_21354);
xor U25860 (N_25860,N_23047,N_22127);
xor U25861 (N_25861,N_22845,N_23937);
and U25862 (N_25862,N_23163,N_22244);
or U25863 (N_25863,N_22249,N_21780);
or U25864 (N_25864,N_21266,N_22098);
nor U25865 (N_25865,N_23371,N_22128);
nand U25866 (N_25866,N_21528,N_22450);
xnor U25867 (N_25867,N_21501,N_22235);
nor U25868 (N_25868,N_21008,N_22211);
and U25869 (N_25869,N_22297,N_23865);
and U25870 (N_25870,N_23109,N_23325);
nand U25871 (N_25871,N_22263,N_22462);
nor U25872 (N_25872,N_23610,N_22858);
xnor U25873 (N_25873,N_22404,N_23481);
nand U25874 (N_25874,N_21842,N_22128);
or U25875 (N_25875,N_21087,N_21261);
and U25876 (N_25876,N_23287,N_21308);
nand U25877 (N_25877,N_22454,N_23101);
xor U25878 (N_25878,N_22725,N_21389);
nor U25879 (N_25879,N_21244,N_21548);
xnor U25880 (N_25880,N_23115,N_22921);
nand U25881 (N_25881,N_22355,N_21403);
xor U25882 (N_25882,N_23803,N_21061);
xnor U25883 (N_25883,N_21170,N_22492);
and U25884 (N_25884,N_21745,N_22855);
nor U25885 (N_25885,N_22166,N_23481);
or U25886 (N_25886,N_22909,N_22107);
nand U25887 (N_25887,N_21948,N_21525);
or U25888 (N_25888,N_22299,N_23171);
and U25889 (N_25889,N_21066,N_21636);
nor U25890 (N_25890,N_22911,N_23658);
nor U25891 (N_25891,N_22983,N_21409);
nor U25892 (N_25892,N_21503,N_23550);
or U25893 (N_25893,N_23695,N_23027);
and U25894 (N_25894,N_23779,N_23214);
or U25895 (N_25895,N_23615,N_23797);
nand U25896 (N_25896,N_23245,N_21528);
xnor U25897 (N_25897,N_23424,N_21707);
or U25898 (N_25898,N_21338,N_23006);
nor U25899 (N_25899,N_23564,N_23193);
or U25900 (N_25900,N_22906,N_21938);
xnor U25901 (N_25901,N_21957,N_21172);
nor U25902 (N_25902,N_23839,N_22961);
xor U25903 (N_25903,N_21581,N_22714);
nand U25904 (N_25904,N_21978,N_23509);
xor U25905 (N_25905,N_23233,N_21633);
xnor U25906 (N_25906,N_22873,N_22644);
nor U25907 (N_25907,N_22995,N_23861);
and U25908 (N_25908,N_23312,N_22072);
nor U25909 (N_25909,N_21909,N_21528);
or U25910 (N_25910,N_23561,N_22145);
or U25911 (N_25911,N_22734,N_22572);
nand U25912 (N_25912,N_23631,N_21019);
nand U25913 (N_25913,N_23176,N_21987);
xnor U25914 (N_25914,N_21177,N_23857);
nor U25915 (N_25915,N_21753,N_21276);
or U25916 (N_25916,N_22251,N_21375);
nor U25917 (N_25917,N_21819,N_21468);
nand U25918 (N_25918,N_21561,N_23106);
nand U25919 (N_25919,N_23157,N_21134);
and U25920 (N_25920,N_23186,N_22722);
xnor U25921 (N_25921,N_22289,N_21161);
and U25922 (N_25922,N_22765,N_23166);
and U25923 (N_25923,N_23990,N_22892);
and U25924 (N_25924,N_22132,N_23459);
xor U25925 (N_25925,N_21765,N_21651);
and U25926 (N_25926,N_21591,N_21643);
xnor U25927 (N_25927,N_23911,N_21203);
xnor U25928 (N_25928,N_23263,N_22510);
nor U25929 (N_25929,N_21468,N_21829);
or U25930 (N_25930,N_22092,N_22669);
or U25931 (N_25931,N_23647,N_23456);
xnor U25932 (N_25932,N_21374,N_21110);
nor U25933 (N_25933,N_23680,N_22706);
and U25934 (N_25934,N_23869,N_23314);
nor U25935 (N_25935,N_22841,N_23540);
and U25936 (N_25936,N_22340,N_23618);
and U25937 (N_25937,N_21483,N_22774);
nor U25938 (N_25938,N_22586,N_22621);
nand U25939 (N_25939,N_21909,N_21449);
or U25940 (N_25940,N_23488,N_23126);
xnor U25941 (N_25941,N_21467,N_21294);
or U25942 (N_25942,N_23389,N_23977);
or U25943 (N_25943,N_21903,N_21070);
nand U25944 (N_25944,N_21474,N_22513);
or U25945 (N_25945,N_21539,N_22418);
nand U25946 (N_25946,N_21063,N_22463);
nand U25947 (N_25947,N_23810,N_22584);
or U25948 (N_25948,N_22953,N_21425);
and U25949 (N_25949,N_23895,N_21968);
or U25950 (N_25950,N_22122,N_23440);
xor U25951 (N_25951,N_23475,N_21198);
nor U25952 (N_25952,N_22756,N_23017);
nand U25953 (N_25953,N_21592,N_22411);
and U25954 (N_25954,N_23362,N_22691);
or U25955 (N_25955,N_23698,N_22839);
or U25956 (N_25956,N_23322,N_23796);
nor U25957 (N_25957,N_23060,N_21956);
and U25958 (N_25958,N_23709,N_22270);
and U25959 (N_25959,N_23476,N_21226);
nand U25960 (N_25960,N_21572,N_23481);
nor U25961 (N_25961,N_21164,N_21852);
and U25962 (N_25962,N_23219,N_21381);
xnor U25963 (N_25963,N_21657,N_21470);
xor U25964 (N_25964,N_23015,N_21507);
xnor U25965 (N_25965,N_21227,N_21982);
nand U25966 (N_25966,N_22921,N_21538);
xor U25967 (N_25967,N_21156,N_22333);
nor U25968 (N_25968,N_22154,N_21957);
nand U25969 (N_25969,N_23867,N_21272);
xor U25970 (N_25970,N_21708,N_23778);
and U25971 (N_25971,N_21346,N_23650);
or U25972 (N_25972,N_23822,N_22172);
nor U25973 (N_25973,N_21463,N_21564);
and U25974 (N_25974,N_23310,N_22613);
and U25975 (N_25975,N_22576,N_22996);
xnor U25976 (N_25976,N_21710,N_23096);
nor U25977 (N_25977,N_21201,N_21678);
and U25978 (N_25978,N_22954,N_21760);
nor U25979 (N_25979,N_23826,N_21174);
nor U25980 (N_25980,N_21763,N_22012);
nand U25981 (N_25981,N_23553,N_22287);
nor U25982 (N_25982,N_21545,N_23084);
xnor U25983 (N_25983,N_23166,N_21849);
xor U25984 (N_25984,N_21296,N_23825);
nor U25985 (N_25985,N_21315,N_23604);
nor U25986 (N_25986,N_22750,N_23090);
xnor U25987 (N_25987,N_21923,N_23443);
nor U25988 (N_25988,N_21350,N_21729);
and U25989 (N_25989,N_22491,N_22156);
nand U25990 (N_25990,N_23344,N_21927);
nand U25991 (N_25991,N_23074,N_22962);
nor U25992 (N_25992,N_23798,N_23760);
and U25993 (N_25993,N_23494,N_21663);
xor U25994 (N_25994,N_22897,N_23788);
nand U25995 (N_25995,N_23386,N_21873);
nand U25996 (N_25996,N_22294,N_21374);
nor U25997 (N_25997,N_21111,N_22026);
xnor U25998 (N_25998,N_23393,N_23459);
or U25999 (N_25999,N_22251,N_21599);
nand U26000 (N_26000,N_22306,N_23183);
or U26001 (N_26001,N_22065,N_21351);
xor U26002 (N_26002,N_23858,N_22757);
and U26003 (N_26003,N_23797,N_21298);
or U26004 (N_26004,N_22905,N_23889);
xnor U26005 (N_26005,N_23953,N_21360);
or U26006 (N_26006,N_22185,N_22616);
or U26007 (N_26007,N_22856,N_22820);
and U26008 (N_26008,N_21693,N_23021);
xnor U26009 (N_26009,N_21968,N_22274);
and U26010 (N_26010,N_22173,N_21372);
or U26011 (N_26011,N_23712,N_23353);
and U26012 (N_26012,N_22648,N_22560);
xnor U26013 (N_26013,N_22808,N_23640);
nand U26014 (N_26014,N_22736,N_23569);
or U26015 (N_26015,N_23958,N_21132);
nor U26016 (N_26016,N_23479,N_21274);
or U26017 (N_26017,N_22232,N_21102);
nor U26018 (N_26018,N_22329,N_21266);
xnor U26019 (N_26019,N_21547,N_22134);
nand U26020 (N_26020,N_21712,N_23494);
nor U26021 (N_26021,N_21105,N_23947);
or U26022 (N_26022,N_23064,N_21310);
xor U26023 (N_26023,N_23534,N_21838);
nand U26024 (N_26024,N_21626,N_21274);
or U26025 (N_26025,N_21833,N_22463);
nor U26026 (N_26026,N_22871,N_21662);
xor U26027 (N_26027,N_22738,N_23192);
nor U26028 (N_26028,N_23327,N_21455);
or U26029 (N_26029,N_21580,N_22985);
nor U26030 (N_26030,N_21582,N_21476);
xnor U26031 (N_26031,N_22287,N_23875);
nor U26032 (N_26032,N_23840,N_23944);
nor U26033 (N_26033,N_23015,N_23798);
and U26034 (N_26034,N_22459,N_22522);
or U26035 (N_26035,N_23647,N_22600);
and U26036 (N_26036,N_21165,N_21868);
or U26037 (N_26037,N_23494,N_22793);
xor U26038 (N_26038,N_23057,N_21109);
xor U26039 (N_26039,N_21537,N_21192);
and U26040 (N_26040,N_22083,N_23341);
nand U26041 (N_26041,N_23400,N_21394);
nand U26042 (N_26042,N_21792,N_22816);
and U26043 (N_26043,N_23138,N_23809);
nor U26044 (N_26044,N_21027,N_22183);
nor U26045 (N_26045,N_23836,N_23146);
nor U26046 (N_26046,N_22936,N_23755);
and U26047 (N_26047,N_21370,N_21407);
nor U26048 (N_26048,N_23065,N_22987);
xor U26049 (N_26049,N_23035,N_23905);
and U26050 (N_26050,N_21914,N_23252);
or U26051 (N_26051,N_23274,N_23400);
or U26052 (N_26052,N_23549,N_23386);
nor U26053 (N_26053,N_21830,N_21407);
nor U26054 (N_26054,N_23355,N_23332);
or U26055 (N_26055,N_22417,N_21750);
nor U26056 (N_26056,N_22323,N_22601);
nand U26057 (N_26057,N_21107,N_22177);
xnor U26058 (N_26058,N_22752,N_23799);
nand U26059 (N_26059,N_23804,N_22647);
xnor U26060 (N_26060,N_21244,N_21740);
or U26061 (N_26061,N_23914,N_21729);
xor U26062 (N_26062,N_23062,N_21365);
and U26063 (N_26063,N_21501,N_23913);
xnor U26064 (N_26064,N_23521,N_21037);
nor U26065 (N_26065,N_23362,N_23332);
xnor U26066 (N_26066,N_22948,N_23729);
and U26067 (N_26067,N_21127,N_23133);
and U26068 (N_26068,N_21846,N_21947);
xnor U26069 (N_26069,N_21190,N_22263);
or U26070 (N_26070,N_21028,N_21994);
xnor U26071 (N_26071,N_21280,N_23322);
or U26072 (N_26072,N_21646,N_22471);
xnor U26073 (N_26073,N_22307,N_21775);
nor U26074 (N_26074,N_21248,N_22718);
and U26075 (N_26075,N_22144,N_22435);
and U26076 (N_26076,N_22199,N_23508);
and U26077 (N_26077,N_21929,N_21903);
nand U26078 (N_26078,N_21293,N_23968);
nand U26079 (N_26079,N_23153,N_21392);
nand U26080 (N_26080,N_23479,N_21162);
xnor U26081 (N_26081,N_21936,N_23173);
and U26082 (N_26082,N_23278,N_21124);
or U26083 (N_26083,N_21789,N_22852);
xor U26084 (N_26084,N_21457,N_21347);
and U26085 (N_26085,N_21889,N_22872);
or U26086 (N_26086,N_23741,N_22514);
or U26087 (N_26087,N_21715,N_22283);
xor U26088 (N_26088,N_21171,N_23903);
nor U26089 (N_26089,N_21235,N_22090);
or U26090 (N_26090,N_22682,N_21208);
nand U26091 (N_26091,N_23952,N_21473);
nor U26092 (N_26092,N_21760,N_22512);
xor U26093 (N_26093,N_21057,N_21996);
nor U26094 (N_26094,N_23715,N_21890);
or U26095 (N_26095,N_21807,N_22956);
xor U26096 (N_26096,N_21577,N_21799);
xor U26097 (N_26097,N_23313,N_23641);
nand U26098 (N_26098,N_22659,N_21787);
or U26099 (N_26099,N_22826,N_21748);
xnor U26100 (N_26100,N_23943,N_22333);
xor U26101 (N_26101,N_21197,N_22350);
or U26102 (N_26102,N_21474,N_22188);
and U26103 (N_26103,N_21352,N_21477);
and U26104 (N_26104,N_21519,N_22235);
and U26105 (N_26105,N_21688,N_22966);
xnor U26106 (N_26106,N_22505,N_22267);
nand U26107 (N_26107,N_22884,N_21871);
or U26108 (N_26108,N_23576,N_22933);
nand U26109 (N_26109,N_21201,N_23643);
and U26110 (N_26110,N_21984,N_23660);
and U26111 (N_26111,N_22126,N_23501);
nor U26112 (N_26112,N_23805,N_23538);
xor U26113 (N_26113,N_21040,N_23113);
and U26114 (N_26114,N_23570,N_23432);
or U26115 (N_26115,N_22932,N_21067);
nand U26116 (N_26116,N_22439,N_23352);
or U26117 (N_26117,N_21626,N_23337);
nand U26118 (N_26118,N_23148,N_23645);
nor U26119 (N_26119,N_23175,N_23736);
or U26120 (N_26120,N_21098,N_23420);
and U26121 (N_26121,N_22984,N_22819);
and U26122 (N_26122,N_23182,N_21770);
and U26123 (N_26123,N_22161,N_23933);
xnor U26124 (N_26124,N_22353,N_21624);
nand U26125 (N_26125,N_21804,N_22821);
nand U26126 (N_26126,N_21191,N_22275);
nor U26127 (N_26127,N_22692,N_22842);
or U26128 (N_26128,N_23129,N_22001);
nand U26129 (N_26129,N_21270,N_21172);
nor U26130 (N_26130,N_23939,N_23305);
and U26131 (N_26131,N_23635,N_21656);
and U26132 (N_26132,N_23653,N_21341);
and U26133 (N_26133,N_22336,N_21189);
or U26134 (N_26134,N_22388,N_22448);
xor U26135 (N_26135,N_21147,N_21067);
nand U26136 (N_26136,N_21427,N_21271);
nand U26137 (N_26137,N_23804,N_22886);
nor U26138 (N_26138,N_22221,N_23515);
or U26139 (N_26139,N_23242,N_23800);
or U26140 (N_26140,N_23121,N_23303);
or U26141 (N_26141,N_23222,N_21866);
xor U26142 (N_26142,N_21548,N_21361);
nor U26143 (N_26143,N_21046,N_21182);
nand U26144 (N_26144,N_21046,N_22561);
and U26145 (N_26145,N_21279,N_23796);
nand U26146 (N_26146,N_21526,N_21726);
nand U26147 (N_26147,N_21705,N_21912);
nand U26148 (N_26148,N_22376,N_22549);
or U26149 (N_26149,N_21016,N_21957);
nand U26150 (N_26150,N_21285,N_21183);
and U26151 (N_26151,N_23735,N_23600);
nand U26152 (N_26152,N_22621,N_23486);
and U26153 (N_26153,N_23762,N_21930);
and U26154 (N_26154,N_22350,N_23355);
nor U26155 (N_26155,N_23692,N_22225);
nor U26156 (N_26156,N_21470,N_21131);
nand U26157 (N_26157,N_22530,N_22639);
or U26158 (N_26158,N_22861,N_21909);
nor U26159 (N_26159,N_23377,N_23230);
nor U26160 (N_26160,N_22862,N_21411);
or U26161 (N_26161,N_21534,N_22102);
xor U26162 (N_26162,N_21145,N_23459);
nor U26163 (N_26163,N_21574,N_21945);
nand U26164 (N_26164,N_22042,N_22402);
nand U26165 (N_26165,N_22556,N_22618);
or U26166 (N_26166,N_21232,N_22818);
and U26167 (N_26167,N_21164,N_21239);
nand U26168 (N_26168,N_23306,N_22668);
xnor U26169 (N_26169,N_22831,N_21546);
nor U26170 (N_26170,N_23525,N_21400);
nor U26171 (N_26171,N_21974,N_23528);
and U26172 (N_26172,N_22520,N_21548);
and U26173 (N_26173,N_23390,N_22559);
xor U26174 (N_26174,N_21796,N_23311);
nand U26175 (N_26175,N_23891,N_21052);
nor U26176 (N_26176,N_21525,N_21453);
nand U26177 (N_26177,N_21441,N_22102);
nand U26178 (N_26178,N_21024,N_23285);
nand U26179 (N_26179,N_22418,N_21938);
and U26180 (N_26180,N_21765,N_21365);
xor U26181 (N_26181,N_23038,N_23541);
and U26182 (N_26182,N_22402,N_23737);
xor U26183 (N_26183,N_22845,N_22244);
or U26184 (N_26184,N_21018,N_21760);
and U26185 (N_26185,N_22615,N_23483);
and U26186 (N_26186,N_22345,N_21459);
nand U26187 (N_26187,N_22910,N_21157);
xnor U26188 (N_26188,N_23409,N_22705);
nand U26189 (N_26189,N_21269,N_23827);
nor U26190 (N_26190,N_23508,N_22263);
nand U26191 (N_26191,N_21503,N_22940);
or U26192 (N_26192,N_23565,N_23729);
nor U26193 (N_26193,N_22907,N_23004);
xor U26194 (N_26194,N_23221,N_23978);
xnor U26195 (N_26195,N_21933,N_23969);
nor U26196 (N_26196,N_23822,N_23180);
nor U26197 (N_26197,N_23257,N_23234);
or U26198 (N_26198,N_23127,N_22616);
xnor U26199 (N_26199,N_22941,N_23418);
nand U26200 (N_26200,N_22706,N_23244);
nand U26201 (N_26201,N_22273,N_21505);
xor U26202 (N_26202,N_23674,N_23969);
or U26203 (N_26203,N_21834,N_22777);
or U26204 (N_26204,N_23222,N_23960);
nor U26205 (N_26205,N_22803,N_21873);
and U26206 (N_26206,N_22346,N_21499);
or U26207 (N_26207,N_22186,N_21175);
and U26208 (N_26208,N_21975,N_23978);
and U26209 (N_26209,N_22141,N_23613);
nor U26210 (N_26210,N_23925,N_22499);
and U26211 (N_26211,N_23948,N_22792);
xnor U26212 (N_26212,N_21705,N_22219);
or U26213 (N_26213,N_22386,N_22928);
nand U26214 (N_26214,N_23612,N_23275);
or U26215 (N_26215,N_22102,N_23109);
xnor U26216 (N_26216,N_22704,N_21379);
nor U26217 (N_26217,N_22399,N_22708);
or U26218 (N_26218,N_21925,N_21591);
nand U26219 (N_26219,N_22977,N_21236);
or U26220 (N_26220,N_21628,N_22895);
or U26221 (N_26221,N_22965,N_23160);
nor U26222 (N_26222,N_21214,N_21958);
xnor U26223 (N_26223,N_22912,N_21465);
nor U26224 (N_26224,N_21189,N_23174);
and U26225 (N_26225,N_22606,N_23575);
or U26226 (N_26226,N_21259,N_21576);
xor U26227 (N_26227,N_23513,N_23113);
nand U26228 (N_26228,N_21805,N_21884);
xnor U26229 (N_26229,N_23252,N_22264);
nor U26230 (N_26230,N_23066,N_21538);
nand U26231 (N_26231,N_22554,N_22962);
xnor U26232 (N_26232,N_23039,N_22156);
xnor U26233 (N_26233,N_21108,N_21210);
and U26234 (N_26234,N_22296,N_21916);
nand U26235 (N_26235,N_23975,N_23594);
nor U26236 (N_26236,N_22870,N_22845);
or U26237 (N_26237,N_23485,N_23933);
and U26238 (N_26238,N_22226,N_21969);
nor U26239 (N_26239,N_23998,N_23727);
nand U26240 (N_26240,N_21722,N_22616);
or U26241 (N_26241,N_22923,N_21829);
or U26242 (N_26242,N_22885,N_22033);
and U26243 (N_26243,N_21300,N_21554);
nand U26244 (N_26244,N_23159,N_23949);
or U26245 (N_26245,N_21376,N_21238);
nand U26246 (N_26246,N_22423,N_21584);
or U26247 (N_26247,N_22793,N_22465);
and U26248 (N_26248,N_22228,N_23875);
and U26249 (N_26249,N_21721,N_22654);
xnor U26250 (N_26250,N_23267,N_23144);
and U26251 (N_26251,N_22457,N_23702);
nor U26252 (N_26252,N_23410,N_21630);
and U26253 (N_26253,N_21770,N_23000);
nor U26254 (N_26254,N_23315,N_23724);
or U26255 (N_26255,N_21074,N_23298);
nand U26256 (N_26256,N_22367,N_23610);
or U26257 (N_26257,N_23244,N_22335);
or U26258 (N_26258,N_23136,N_21112);
nand U26259 (N_26259,N_22738,N_21133);
xnor U26260 (N_26260,N_22675,N_21373);
or U26261 (N_26261,N_21591,N_21889);
xor U26262 (N_26262,N_22700,N_22872);
nor U26263 (N_26263,N_23313,N_23949);
nand U26264 (N_26264,N_23232,N_23435);
or U26265 (N_26265,N_23446,N_22968);
nand U26266 (N_26266,N_22293,N_21548);
and U26267 (N_26267,N_23369,N_22378);
and U26268 (N_26268,N_22642,N_21848);
nor U26269 (N_26269,N_22318,N_22796);
nor U26270 (N_26270,N_22492,N_23363);
and U26271 (N_26271,N_21194,N_23450);
xor U26272 (N_26272,N_23535,N_23385);
nand U26273 (N_26273,N_22313,N_22468);
nand U26274 (N_26274,N_22416,N_22966);
nor U26275 (N_26275,N_23664,N_23089);
or U26276 (N_26276,N_22069,N_23028);
nor U26277 (N_26277,N_22818,N_22051);
nand U26278 (N_26278,N_23810,N_23356);
xor U26279 (N_26279,N_23167,N_22001);
and U26280 (N_26280,N_23137,N_22103);
or U26281 (N_26281,N_23284,N_21502);
nand U26282 (N_26282,N_23586,N_23642);
nand U26283 (N_26283,N_22692,N_23685);
xnor U26284 (N_26284,N_23510,N_21964);
nor U26285 (N_26285,N_21120,N_22392);
and U26286 (N_26286,N_23469,N_21472);
or U26287 (N_26287,N_23390,N_22974);
and U26288 (N_26288,N_22008,N_21301);
nand U26289 (N_26289,N_21327,N_22553);
xor U26290 (N_26290,N_23165,N_23124);
or U26291 (N_26291,N_21148,N_21895);
xor U26292 (N_26292,N_23958,N_23910);
and U26293 (N_26293,N_23418,N_22724);
nor U26294 (N_26294,N_21499,N_23663);
nor U26295 (N_26295,N_23041,N_21692);
xor U26296 (N_26296,N_22551,N_22783);
nor U26297 (N_26297,N_21265,N_23570);
or U26298 (N_26298,N_23416,N_22536);
and U26299 (N_26299,N_23818,N_22353);
nand U26300 (N_26300,N_23818,N_21708);
xnor U26301 (N_26301,N_22612,N_22216);
nor U26302 (N_26302,N_22473,N_21983);
or U26303 (N_26303,N_21855,N_23109);
xnor U26304 (N_26304,N_23470,N_23569);
nand U26305 (N_26305,N_23049,N_22179);
nor U26306 (N_26306,N_21709,N_23834);
nor U26307 (N_26307,N_21005,N_21577);
and U26308 (N_26308,N_23826,N_22007);
and U26309 (N_26309,N_22541,N_21678);
nand U26310 (N_26310,N_23547,N_23426);
nand U26311 (N_26311,N_21274,N_21081);
nand U26312 (N_26312,N_21363,N_23237);
or U26313 (N_26313,N_23842,N_23677);
xnor U26314 (N_26314,N_21182,N_22044);
nand U26315 (N_26315,N_21691,N_23441);
xor U26316 (N_26316,N_21275,N_23087);
and U26317 (N_26317,N_21590,N_21436);
and U26318 (N_26318,N_22156,N_23309);
and U26319 (N_26319,N_23782,N_23170);
nand U26320 (N_26320,N_23134,N_21103);
xor U26321 (N_26321,N_23843,N_22954);
and U26322 (N_26322,N_23548,N_22642);
and U26323 (N_26323,N_23780,N_22718);
nor U26324 (N_26324,N_21092,N_21249);
nor U26325 (N_26325,N_21978,N_23040);
nor U26326 (N_26326,N_22099,N_21497);
xnor U26327 (N_26327,N_22911,N_23969);
nor U26328 (N_26328,N_22733,N_21695);
nand U26329 (N_26329,N_23109,N_22971);
nor U26330 (N_26330,N_22943,N_23123);
nand U26331 (N_26331,N_21157,N_22740);
or U26332 (N_26332,N_23720,N_22539);
or U26333 (N_26333,N_21271,N_21650);
xor U26334 (N_26334,N_23439,N_23593);
xnor U26335 (N_26335,N_21438,N_23160);
xnor U26336 (N_26336,N_21291,N_22190);
xor U26337 (N_26337,N_23455,N_22823);
xor U26338 (N_26338,N_23826,N_23793);
nor U26339 (N_26339,N_21848,N_23312);
nor U26340 (N_26340,N_23445,N_23289);
nand U26341 (N_26341,N_21247,N_22537);
xor U26342 (N_26342,N_22250,N_22910);
nor U26343 (N_26343,N_23472,N_23017);
nand U26344 (N_26344,N_21130,N_23818);
xor U26345 (N_26345,N_21337,N_21820);
and U26346 (N_26346,N_23789,N_23790);
nand U26347 (N_26347,N_21211,N_21099);
nor U26348 (N_26348,N_21586,N_23113);
nand U26349 (N_26349,N_21320,N_22716);
nand U26350 (N_26350,N_22728,N_23751);
nor U26351 (N_26351,N_22368,N_21198);
or U26352 (N_26352,N_22368,N_22990);
xnor U26353 (N_26353,N_21386,N_21143);
xor U26354 (N_26354,N_23758,N_23905);
nor U26355 (N_26355,N_23305,N_21018);
nand U26356 (N_26356,N_22326,N_21387);
nand U26357 (N_26357,N_23498,N_22204);
or U26358 (N_26358,N_23534,N_22759);
nand U26359 (N_26359,N_21803,N_23221);
nor U26360 (N_26360,N_22703,N_22913);
xnor U26361 (N_26361,N_23399,N_22497);
or U26362 (N_26362,N_22086,N_22478);
or U26363 (N_26363,N_21906,N_21452);
or U26364 (N_26364,N_23672,N_23921);
nor U26365 (N_26365,N_21140,N_21107);
and U26366 (N_26366,N_21065,N_21192);
and U26367 (N_26367,N_21524,N_21860);
or U26368 (N_26368,N_22903,N_23258);
or U26369 (N_26369,N_22888,N_22407);
xnor U26370 (N_26370,N_21774,N_22717);
nand U26371 (N_26371,N_23993,N_22239);
nor U26372 (N_26372,N_21918,N_22707);
and U26373 (N_26373,N_23701,N_21635);
nor U26374 (N_26374,N_21257,N_23609);
and U26375 (N_26375,N_23898,N_23287);
and U26376 (N_26376,N_23023,N_21898);
nor U26377 (N_26377,N_21343,N_21050);
nor U26378 (N_26378,N_21593,N_22610);
xnor U26379 (N_26379,N_21247,N_21136);
xor U26380 (N_26380,N_21821,N_22705);
or U26381 (N_26381,N_21490,N_22581);
nand U26382 (N_26382,N_21343,N_21411);
xnor U26383 (N_26383,N_21303,N_21674);
xor U26384 (N_26384,N_23520,N_23820);
nor U26385 (N_26385,N_22802,N_21627);
xor U26386 (N_26386,N_21327,N_21333);
nand U26387 (N_26387,N_22835,N_21017);
nand U26388 (N_26388,N_22299,N_23810);
xor U26389 (N_26389,N_22474,N_22197);
nor U26390 (N_26390,N_21388,N_21681);
nand U26391 (N_26391,N_23585,N_21644);
nand U26392 (N_26392,N_23746,N_22480);
nor U26393 (N_26393,N_21123,N_23040);
or U26394 (N_26394,N_22157,N_22821);
or U26395 (N_26395,N_23080,N_23431);
or U26396 (N_26396,N_23834,N_23032);
and U26397 (N_26397,N_21366,N_23540);
xnor U26398 (N_26398,N_22341,N_23827);
or U26399 (N_26399,N_21962,N_23548);
nor U26400 (N_26400,N_23778,N_23603);
nand U26401 (N_26401,N_22329,N_21395);
xor U26402 (N_26402,N_21685,N_21450);
and U26403 (N_26403,N_22152,N_23749);
and U26404 (N_26404,N_21825,N_21175);
xnor U26405 (N_26405,N_22921,N_23788);
nand U26406 (N_26406,N_23113,N_22319);
and U26407 (N_26407,N_23822,N_21971);
xor U26408 (N_26408,N_23601,N_22530);
xnor U26409 (N_26409,N_22841,N_22215);
nand U26410 (N_26410,N_23374,N_21414);
or U26411 (N_26411,N_23090,N_21211);
or U26412 (N_26412,N_22540,N_22679);
xor U26413 (N_26413,N_23673,N_23846);
and U26414 (N_26414,N_22267,N_23557);
and U26415 (N_26415,N_23602,N_22164);
xnor U26416 (N_26416,N_22054,N_21715);
and U26417 (N_26417,N_23863,N_22345);
and U26418 (N_26418,N_23574,N_21931);
nand U26419 (N_26419,N_21226,N_21764);
nor U26420 (N_26420,N_23656,N_22103);
xnor U26421 (N_26421,N_23669,N_21916);
or U26422 (N_26422,N_22895,N_23261);
or U26423 (N_26423,N_23323,N_23644);
or U26424 (N_26424,N_22124,N_22117);
xnor U26425 (N_26425,N_21725,N_23804);
nor U26426 (N_26426,N_22328,N_21837);
and U26427 (N_26427,N_21260,N_22070);
xor U26428 (N_26428,N_23050,N_23342);
and U26429 (N_26429,N_23702,N_21354);
xnor U26430 (N_26430,N_22114,N_23160);
or U26431 (N_26431,N_22426,N_23086);
nor U26432 (N_26432,N_23982,N_22458);
xor U26433 (N_26433,N_22685,N_23642);
xnor U26434 (N_26434,N_23840,N_23811);
nand U26435 (N_26435,N_22570,N_23151);
xnor U26436 (N_26436,N_23464,N_22391);
nor U26437 (N_26437,N_21673,N_21148);
nand U26438 (N_26438,N_23962,N_22615);
nor U26439 (N_26439,N_22657,N_22108);
nand U26440 (N_26440,N_21891,N_21223);
and U26441 (N_26441,N_23280,N_22071);
nor U26442 (N_26442,N_23228,N_23914);
nand U26443 (N_26443,N_22945,N_23817);
xor U26444 (N_26444,N_21579,N_23460);
nand U26445 (N_26445,N_23178,N_23369);
or U26446 (N_26446,N_21201,N_23175);
and U26447 (N_26447,N_22891,N_21052);
nor U26448 (N_26448,N_22322,N_22599);
and U26449 (N_26449,N_21875,N_23484);
xor U26450 (N_26450,N_22422,N_21472);
nand U26451 (N_26451,N_23160,N_21618);
nand U26452 (N_26452,N_21262,N_21681);
xor U26453 (N_26453,N_21225,N_21670);
and U26454 (N_26454,N_22918,N_21168);
and U26455 (N_26455,N_23998,N_23916);
xnor U26456 (N_26456,N_22376,N_23183);
or U26457 (N_26457,N_21603,N_23329);
nand U26458 (N_26458,N_23299,N_22003);
xnor U26459 (N_26459,N_22111,N_22814);
nand U26460 (N_26460,N_23737,N_22577);
or U26461 (N_26461,N_22506,N_21071);
and U26462 (N_26462,N_23861,N_22936);
or U26463 (N_26463,N_22118,N_21731);
and U26464 (N_26464,N_22270,N_21294);
and U26465 (N_26465,N_21815,N_22662);
and U26466 (N_26466,N_23642,N_23975);
xor U26467 (N_26467,N_23121,N_21919);
and U26468 (N_26468,N_21610,N_23216);
or U26469 (N_26469,N_23900,N_23174);
xnor U26470 (N_26470,N_23544,N_22698);
xnor U26471 (N_26471,N_23971,N_22626);
xnor U26472 (N_26472,N_23201,N_22228);
or U26473 (N_26473,N_23571,N_23389);
or U26474 (N_26474,N_23540,N_22688);
nand U26475 (N_26475,N_22479,N_22807);
nand U26476 (N_26476,N_21980,N_21828);
nand U26477 (N_26477,N_23798,N_22221);
nor U26478 (N_26478,N_23218,N_21898);
nand U26479 (N_26479,N_21072,N_21420);
nand U26480 (N_26480,N_23824,N_23420);
and U26481 (N_26481,N_21591,N_22685);
and U26482 (N_26482,N_23116,N_23638);
or U26483 (N_26483,N_21689,N_22709);
and U26484 (N_26484,N_22290,N_23587);
nand U26485 (N_26485,N_22501,N_22790);
nor U26486 (N_26486,N_22175,N_21085);
xnor U26487 (N_26487,N_21381,N_23429);
xnor U26488 (N_26488,N_23831,N_23688);
and U26489 (N_26489,N_22523,N_22286);
xnor U26490 (N_26490,N_22252,N_22210);
nor U26491 (N_26491,N_23313,N_21609);
or U26492 (N_26492,N_22283,N_23153);
nand U26493 (N_26493,N_22498,N_23047);
xnor U26494 (N_26494,N_21289,N_23523);
and U26495 (N_26495,N_22121,N_23100);
nand U26496 (N_26496,N_23963,N_21159);
nor U26497 (N_26497,N_22007,N_21810);
or U26498 (N_26498,N_22086,N_23462);
xnor U26499 (N_26499,N_22949,N_23525);
and U26500 (N_26500,N_22548,N_21914);
xnor U26501 (N_26501,N_22745,N_21969);
and U26502 (N_26502,N_22118,N_22358);
or U26503 (N_26503,N_23290,N_22190);
nand U26504 (N_26504,N_23685,N_23867);
and U26505 (N_26505,N_22778,N_22668);
xor U26506 (N_26506,N_21533,N_23096);
or U26507 (N_26507,N_23284,N_23651);
and U26508 (N_26508,N_23754,N_23035);
xnor U26509 (N_26509,N_23693,N_21898);
and U26510 (N_26510,N_23663,N_23100);
or U26511 (N_26511,N_23837,N_22932);
nor U26512 (N_26512,N_23241,N_22748);
nor U26513 (N_26513,N_23505,N_23389);
or U26514 (N_26514,N_23828,N_23144);
nand U26515 (N_26515,N_21383,N_22361);
nand U26516 (N_26516,N_22438,N_22830);
nand U26517 (N_26517,N_23517,N_22801);
or U26518 (N_26518,N_23035,N_22986);
nor U26519 (N_26519,N_22831,N_21762);
or U26520 (N_26520,N_22030,N_21126);
xor U26521 (N_26521,N_21095,N_21618);
nor U26522 (N_26522,N_21852,N_22521);
or U26523 (N_26523,N_23885,N_21580);
xnor U26524 (N_26524,N_23063,N_23226);
or U26525 (N_26525,N_23980,N_22337);
xor U26526 (N_26526,N_23390,N_23359);
and U26527 (N_26527,N_23819,N_21121);
nand U26528 (N_26528,N_23311,N_21210);
nand U26529 (N_26529,N_21162,N_23474);
and U26530 (N_26530,N_21826,N_22229);
nor U26531 (N_26531,N_22479,N_22501);
or U26532 (N_26532,N_22618,N_22288);
nand U26533 (N_26533,N_23413,N_22387);
and U26534 (N_26534,N_22532,N_21004);
or U26535 (N_26535,N_21435,N_22664);
and U26536 (N_26536,N_22557,N_23497);
nor U26537 (N_26537,N_22736,N_21506);
and U26538 (N_26538,N_21148,N_22098);
nand U26539 (N_26539,N_23119,N_21293);
nand U26540 (N_26540,N_23869,N_22763);
nor U26541 (N_26541,N_21544,N_21286);
nand U26542 (N_26542,N_21494,N_22689);
nor U26543 (N_26543,N_23764,N_22013);
and U26544 (N_26544,N_21795,N_22203);
xnor U26545 (N_26545,N_21384,N_22193);
xnor U26546 (N_26546,N_21674,N_21244);
nor U26547 (N_26547,N_21091,N_21090);
and U26548 (N_26548,N_22774,N_22674);
xnor U26549 (N_26549,N_21342,N_22356);
or U26550 (N_26550,N_21087,N_23386);
and U26551 (N_26551,N_22652,N_23039);
xnor U26552 (N_26552,N_21953,N_22798);
nand U26553 (N_26553,N_22162,N_22605);
nand U26554 (N_26554,N_21738,N_23064);
nor U26555 (N_26555,N_21814,N_22309);
nand U26556 (N_26556,N_23036,N_22518);
nand U26557 (N_26557,N_21717,N_23946);
and U26558 (N_26558,N_22471,N_23523);
or U26559 (N_26559,N_23564,N_22758);
and U26560 (N_26560,N_23349,N_23382);
nand U26561 (N_26561,N_22182,N_23024);
xnor U26562 (N_26562,N_21552,N_22505);
xnor U26563 (N_26563,N_23499,N_21403);
and U26564 (N_26564,N_22523,N_21849);
nand U26565 (N_26565,N_22798,N_21193);
nand U26566 (N_26566,N_22749,N_22970);
or U26567 (N_26567,N_23955,N_23624);
xnor U26568 (N_26568,N_23454,N_22967);
or U26569 (N_26569,N_21485,N_21118);
nor U26570 (N_26570,N_22609,N_22371);
xnor U26571 (N_26571,N_21130,N_22968);
and U26572 (N_26572,N_22702,N_22703);
and U26573 (N_26573,N_23948,N_21733);
xnor U26574 (N_26574,N_21102,N_23896);
and U26575 (N_26575,N_21864,N_23406);
and U26576 (N_26576,N_23045,N_21062);
and U26577 (N_26577,N_21752,N_22291);
xnor U26578 (N_26578,N_21013,N_22803);
and U26579 (N_26579,N_21368,N_23476);
or U26580 (N_26580,N_23380,N_21173);
xor U26581 (N_26581,N_23263,N_23660);
or U26582 (N_26582,N_23148,N_21961);
and U26583 (N_26583,N_23928,N_21541);
xor U26584 (N_26584,N_21277,N_21858);
nor U26585 (N_26585,N_21896,N_23801);
nand U26586 (N_26586,N_21795,N_21229);
xnor U26587 (N_26587,N_21280,N_22051);
nand U26588 (N_26588,N_23599,N_23349);
or U26589 (N_26589,N_21878,N_21644);
nor U26590 (N_26590,N_23740,N_22198);
nor U26591 (N_26591,N_21669,N_22540);
nand U26592 (N_26592,N_21733,N_21287);
and U26593 (N_26593,N_23616,N_22126);
xor U26594 (N_26594,N_22916,N_23103);
and U26595 (N_26595,N_21778,N_21386);
and U26596 (N_26596,N_22205,N_22519);
nor U26597 (N_26597,N_22722,N_21094);
or U26598 (N_26598,N_21380,N_21545);
and U26599 (N_26599,N_21630,N_23713);
nor U26600 (N_26600,N_22546,N_22462);
xor U26601 (N_26601,N_21978,N_21908);
and U26602 (N_26602,N_23827,N_22497);
xnor U26603 (N_26603,N_23033,N_21532);
nor U26604 (N_26604,N_23286,N_22127);
xnor U26605 (N_26605,N_23367,N_23137);
nand U26606 (N_26606,N_23750,N_23951);
xnor U26607 (N_26607,N_22142,N_22244);
and U26608 (N_26608,N_23685,N_22383);
nor U26609 (N_26609,N_22135,N_23414);
nand U26610 (N_26610,N_23289,N_22185);
and U26611 (N_26611,N_21538,N_22487);
xnor U26612 (N_26612,N_22123,N_21257);
and U26613 (N_26613,N_22638,N_22524);
and U26614 (N_26614,N_22289,N_22812);
xor U26615 (N_26615,N_21085,N_23067);
and U26616 (N_26616,N_22897,N_21220);
nor U26617 (N_26617,N_23133,N_21822);
xnor U26618 (N_26618,N_22768,N_21670);
and U26619 (N_26619,N_22876,N_23394);
nor U26620 (N_26620,N_21634,N_23388);
xnor U26621 (N_26621,N_22814,N_23261);
xor U26622 (N_26622,N_21660,N_23126);
nand U26623 (N_26623,N_21255,N_21067);
xor U26624 (N_26624,N_21443,N_23960);
nand U26625 (N_26625,N_21284,N_21212);
nand U26626 (N_26626,N_23536,N_21753);
nor U26627 (N_26627,N_21781,N_21101);
nand U26628 (N_26628,N_21593,N_21411);
xor U26629 (N_26629,N_22216,N_23127);
or U26630 (N_26630,N_23625,N_21863);
nor U26631 (N_26631,N_23087,N_22738);
nor U26632 (N_26632,N_22341,N_21741);
nand U26633 (N_26633,N_23144,N_22466);
and U26634 (N_26634,N_21069,N_23873);
nor U26635 (N_26635,N_21789,N_21647);
nor U26636 (N_26636,N_22654,N_22369);
or U26637 (N_26637,N_21198,N_21861);
nor U26638 (N_26638,N_22154,N_21832);
xnor U26639 (N_26639,N_23458,N_22885);
nand U26640 (N_26640,N_22036,N_22945);
nor U26641 (N_26641,N_21073,N_21100);
xnor U26642 (N_26642,N_22712,N_22897);
or U26643 (N_26643,N_23903,N_22236);
nand U26644 (N_26644,N_23004,N_23461);
nand U26645 (N_26645,N_21837,N_21657);
nand U26646 (N_26646,N_23269,N_22433);
nand U26647 (N_26647,N_23579,N_22280);
xor U26648 (N_26648,N_22047,N_22604);
nor U26649 (N_26649,N_21049,N_22917);
or U26650 (N_26650,N_22705,N_21299);
nand U26651 (N_26651,N_22512,N_21485);
nor U26652 (N_26652,N_23942,N_21699);
nand U26653 (N_26653,N_21740,N_23159);
nor U26654 (N_26654,N_22801,N_23502);
and U26655 (N_26655,N_22928,N_21902);
and U26656 (N_26656,N_22621,N_21061);
or U26657 (N_26657,N_23956,N_22528);
and U26658 (N_26658,N_22743,N_23469);
or U26659 (N_26659,N_22197,N_22660);
or U26660 (N_26660,N_21246,N_22938);
xor U26661 (N_26661,N_23379,N_22176);
and U26662 (N_26662,N_22030,N_23636);
and U26663 (N_26663,N_21395,N_22556);
xnor U26664 (N_26664,N_21150,N_21570);
nor U26665 (N_26665,N_21462,N_22149);
or U26666 (N_26666,N_21651,N_21294);
nor U26667 (N_26667,N_22242,N_22022);
or U26668 (N_26668,N_22510,N_21314);
nand U26669 (N_26669,N_21085,N_22999);
nand U26670 (N_26670,N_21257,N_21072);
xnor U26671 (N_26671,N_22011,N_22281);
xor U26672 (N_26672,N_21982,N_21942);
nand U26673 (N_26673,N_21450,N_22981);
nand U26674 (N_26674,N_22758,N_21950);
or U26675 (N_26675,N_22502,N_21998);
nor U26676 (N_26676,N_21707,N_22447);
nor U26677 (N_26677,N_22534,N_21414);
and U26678 (N_26678,N_23263,N_21704);
nor U26679 (N_26679,N_21330,N_22328);
nand U26680 (N_26680,N_22471,N_21565);
or U26681 (N_26681,N_22451,N_21969);
xor U26682 (N_26682,N_21539,N_23357);
and U26683 (N_26683,N_21719,N_22025);
nand U26684 (N_26684,N_23032,N_23474);
xnor U26685 (N_26685,N_22619,N_22179);
and U26686 (N_26686,N_21156,N_21269);
xnor U26687 (N_26687,N_23461,N_22693);
xnor U26688 (N_26688,N_23140,N_23400);
or U26689 (N_26689,N_23376,N_21320);
xnor U26690 (N_26690,N_23179,N_23446);
xor U26691 (N_26691,N_21162,N_22423);
nand U26692 (N_26692,N_21443,N_23706);
and U26693 (N_26693,N_23369,N_22209);
xor U26694 (N_26694,N_23815,N_21508);
or U26695 (N_26695,N_22856,N_21782);
or U26696 (N_26696,N_23315,N_21186);
nand U26697 (N_26697,N_21576,N_23409);
nor U26698 (N_26698,N_21616,N_23749);
xor U26699 (N_26699,N_21106,N_22602);
or U26700 (N_26700,N_21194,N_23995);
or U26701 (N_26701,N_21972,N_23504);
and U26702 (N_26702,N_22608,N_21346);
xor U26703 (N_26703,N_22842,N_22650);
xor U26704 (N_26704,N_21747,N_23778);
xor U26705 (N_26705,N_21920,N_22398);
xnor U26706 (N_26706,N_22043,N_21694);
xnor U26707 (N_26707,N_21850,N_22101);
nor U26708 (N_26708,N_22190,N_23784);
nor U26709 (N_26709,N_23222,N_22108);
nand U26710 (N_26710,N_21273,N_23351);
nand U26711 (N_26711,N_22424,N_23443);
and U26712 (N_26712,N_21976,N_22019);
or U26713 (N_26713,N_23846,N_23865);
or U26714 (N_26714,N_22021,N_23832);
nand U26715 (N_26715,N_23394,N_22071);
and U26716 (N_26716,N_23169,N_23632);
nand U26717 (N_26717,N_22144,N_21506);
nand U26718 (N_26718,N_22542,N_23329);
and U26719 (N_26719,N_21322,N_22116);
nand U26720 (N_26720,N_21236,N_21515);
or U26721 (N_26721,N_22602,N_21361);
xnor U26722 (N_26722,N_21742,N_22755);
and U26723 (N_26723,N_23560,N_22230);
nand U26724 (N_26724,N_23482,N_22043);
nand U26725 (N_26725,N_23884,N_21606);
xor U26726 (N_26726,N_21342,N_23074);
and U26727 (N_26727,N_21429,N_22056);
nor U26728 (N_26728,N_22601,N_21572);
and U26729 (N_26729,N_22718,N_21815);
xor U26730 (N_26730,N_22158,N_23744);
or U26731 (N_26731,N_22639,N_23941);
nor U26732 (N_26732,N_23963,N_21758);
and U26733 (N_26733,N_21548,N_21140);
xor U26734 (N_26734,N_22005,N_23207);
nand U26735 (N_26735,N_23952,N_21375);
nand U26736 (N_26736,N_21657,N_22690);
and U26737 (N_26737,N_21061,N_21173);
xor U26738 (N_26738,N_23014,N_23594);
xnor U26739 (N_26739,N_22391,N_21404);
nor U26740 (N_26740,N_23438,N_22107);
nand U26741 (N_26741,N_23261,N_23509);
xor U26742 (N_26742,N_21604,N_22086);
nand U26743 (N_26743,N_21453,N_21835);
or U26744 (N_26744,N_21029,N_23453);
nand U26745 (N_26745,N_21704,N_23056);
xnor U26746 (N_26746,N_23148,N_23608);
xor U26747 (N_26747,N_21933,N_23215);
nor U26748 (N_26748,N_22824,N_23550);
nor U26749 (N_26749,N_21072,N_22197);
nor U26750 (N_26750,N_22266,N_23121);
or U26751 (N_26751,N_21652,N_22585);
or U26752 (N_26752,N_22676,N_23833);
or U26753 (N_26753,N_22132,N_22138);
or U26754 (N_26754,N_21443,N_22775);
and U26755 (N_26755,N_21010,N_23585);
xnor U26756 (N_26756,N_23661,N_21479);
nand U26757 (N_26757,N_23215,N_22720);
or U26758 (N_26758,N_22736,N_22896);
and U26759 (N_26759,N_21713,N_21647);
xnor U26760 (N_26760,N_23849,N_23664);
nor U26761 (N_26761,N_23572,N_22796);
or U26762 (N_26762,N_21178,N_23415);
nand U26763 (N_26763,N_21536,N_23150);
nand U26764 (N_26764,N_23825,N_23230);
nor U26765 (N_26765,N_21900,N_22703);
or U26766 (N_26766,N_23071,N_23945);
or U26767 (N_26767,N_22649,N_23440);
nand U26768 (N_26768,N_22920,N_22434);
nand U26769 (N_26769,N_21741,N_22550);
nand U26770 (N_26770,N_21014,N_23907);
nand U26771 (N_26771,N_23482,N_21573);
xor U26772 (N_26772,N_23843,N_23079);
and U26773 (N_26773,N_22374,N_22509);
nand U26774 (N_26774,N_22951,N_23039);
nand U26775 (N_26775,N_21044,N_22908);
and U26776 (N_26776,N_23481,N_23996);
and U26777 (N_26777,N_22208,N_21700);
nor U26778 (N_26778,N_21343,N_21627);
nand U26779 (N_26779,N_23426,N_22535);
xnor U26780 (N_26780,N_22611,N_23126);
and U26781 (N_26781,N_21490,N_21909);
nor U26782 (N_26782,N_23821,N_23776);
nor U26783 (N_26783,N_23183,N_23379);
and U26784 (N_26784,N_22165,N_22651);
nand U26785 (N_26785,N_22441,N_22368);
or U26786 (N_26786,N_23344,N_21371);
xor U26787 (N_26787,N_23797,N_21388);
and U26788 (N_26788,N_23461,N_22885);
nor U26789 (N_26789,N_21577,N_22223);
or U26790 (N_26790,N_23684,N_21052);
xnor U26791 (N_26791,N_21199,N_21425);
xnor U26792 (N_26792,N_22895,N_22041);
or U26793 (N_26793,N_22229,N_21669);
or U26794 (N_26794,N_23375,N_23819);
and U26795 (N_26795,N_22659,N_22645);
or U26796 (N_26796,N_23599,N_23950);
nand U26797 (N_26797,N_22969,N_23990);
or U26798 (N_26798,N_21270,N_21260);
xor U26799 (N_26799,N_22792,N_23038);
nand U26800 (N_26800,N_23677,N_23538);
or U26801 (N_26801,N_21154,N_22618);
nand U26802 (N_26802,N_22997,N_21956);
xnor U26803 (N_26803,N_21225,N_23334);
nor U26804 (N_26804,N_22218,N_21696);
nand U26805 (N_26805,N_23299,N_22060);
and U26806 (N_26806,N_22639,N_22978);
and U26807 (N_26807,N_21758,N_23181);
and U26808 (N_26808,N_23282,N_23215);
and U26809 (N_26809,N_23741,N_23497);
or U26810 (N_26810,N_22104,N_23323);
or U26811 (N_26811,N_23570,N_21244);
xnor U26812 (N_26812,N_23688,N_21202);
nand U26813 (N_26813,N_22435,N_23428);
nor U26814 (N_26814,N_23807,N_21486);
and U26815 (N_26815,N_22680,N_21121);
nor U26816 (N_26816,N_21331,N_21423);
nand U26817 (N_26817,N_22299,N_22843);
nand U26818 (N_26818,N_22710,N_23697);
nand U26819 (N_26819,N_23936,N_22882);
nor U26820 (N_26820,N_21766,N_21635);
nand U26821 (N_26821,N_21746,N_22963);
or U26822 (N_26822,N_23643,N_23260);
nand U26823 (N_26823,N_23331,N_23220);
xor U26824 (N_26824,N_21409,N_23948);
nor U26825 (N_26825,N_23517,N_21947);
nand U26826 (N_26826,N_21771,N_21968);
or U26827 (N_26827,N_21923,N_23107);
nor U26828 (N_26828,N_22498,N_22087);
xnor U26829 (N_26829,N_23776,N_23031);
and U26830 (N_26830,N_23467,N_21116);
and U26831 (N_26831,N_21116,N_22692);
or U26832 (N_26832,N_22442,N_23481);
and U26833 (N_26833,N_23457,N_23729);
nor U26834 (N_26834,N_23352,N_23920);
xnor U26835 (N_26835,N_21659,N_21039);
xnor U26836 (N_26836,N_21535,N_21484);
and U26837 (N_26837,N_23125,N_23822);
and U26838 (N_26838,N_21634,N_21268);
nor U26839 (N_26839,N_23860,N_22974);
and U26840 (N_26840,N_21923,N_21980);
nand U26841 (N_26841,N_23897,N_22848);
and U26842 (N_26842,N_22121,N_21268);
xnor U26843 (N_26843,N_23696,N_23985);
xor U26844 (N_26844,N_22009,N_23390);
or U26845 (N_26845,N_21069,N_23378);
or U26846 (N_26846,N_21876,N_23344);
nand U26847 (N_26847,N_22642,N_23469);
nand U26848 (N_26848,N_23526,N_22036);
or U26849 (N_26849,N_23921,N_22980);
xor U26850 (N_26850,N_21313,N_22101);
nand U26851 (N_26851,N_23150,N_23396);
nor U26852 (N_26852,N_22141,N_22115);
or U26853 (N_26853,N_22194,N_21859);
xor U26854 (N_26854,N_22625,N_21851);
or U26855 (N_26855,N_23913,N_23385);
or U26856 (N_26856,N_23737,N_22568);
nand U26857 (N_26857,N_23374,N_21999);
nor U26858 (N_26858,N_23340,N_22674);
and U26859 (N_26859,N_23716,N_23939);
and U26860 (N_26860,N_23638,N_23412);
xnor U26861 (N_26861,N_23580,N_21344);
nand U26862 (N_26862,N_23174,N_22928);
xnor U26863 (N_26863,N_23916,N_22282);
nor U26864 (N_26864,N_23825,N_22282);
or U26865 (N_26865,N_22550,N_21501);
nor U26866 (N_26866,N_22624,N_21761);
nor U26867 (N_26867,N_21704,N_22018);
nand U26868 (N_26868,N_22189,N_23459);
and U26869 (N_26869,N_23269,N_22451);
nand U26870 (N_26870,N_22514,N_23648);
and U26871 (N_26871,N_22672,N_23338);
nor U26872 (N_26872,N_23160,N_22176);
nand U26873 (N_26873,N_23829,N_23111);
nor U26874 (N_26874,N_21952,N_22162);
nor U26875 (N_26875,N_23555,N_23511);
and U26876 (N_26876,N_23456,N_21212);
or U26877 (N_26877,N_22841,N_23723);
nor U26878 (N_26878,N_21018,N_21361);
and U26879 (N_26879,N_23901,N_21649);
nor U26880 (N_26880,N_23863,N_21708);
xnor U26881 (N_26881,N_23726,N_23099);
and U26882 (N_26882,N_21746,N_21349);
xor U26883 (N_26883,N_23039,N_21756);
and U26884 (N_26884,N_21835,N_21868);
or U26885 (N_26885,N_22128,N_21839);
and U26886 (N_26886,N_22709,N_22245);
xor U26887 (N_26887,N_23235,N_21945);
nand U26888 (N_26888,N_22175,N_21962);
or U26889 (N_26889,N_21294,N_22409);
nor U26890 (N_26890,N_21593,N_21128);
xnor U26891 (N_26891,N_22739,N_21675);
and U26892 (N_26892,N_22815,N_21817);
and U26893 (N_26893,N_23080,N_23202);
xnor U26894 (N_26894,N_21166,N_23995);
nor U26895 (N_26895,N_21960,N_22656);
or U26896 (N_26896,N_21139,N_23461);
nor U26897 (N_26897,N_23715,N_23990);
and U26898 (N_26898,N_23928,N_23816);
nor U26899 (N_26899,N_21307,N_21703);
nor U26900 (N_26900,N_23483,N_23150);
xnor U26901 (N_26901,N_23914,N_23012);
nor U26902 (N_26902,N_23990,N_21270);
and U26903 (N_26903,N_21087,N_22950);
and U26904 (N_26904,N_22046,N_22558);
or U26905 (N_26905,N_23824,N_23073);
xnor U26906 (N_26906,N_22588,N_21626);
or U26907 (N_26907,N_22465,N_21042);
nor U26908 (N_26908,N_21421,N_23748);
and U26909 (N_26909,N_22305,N_22587);
nor U26910 (N_26910,N_22024,N_21172);
nor U26911 (N_26911,N_23153,N_21652);
or U26912 (N_26912,N_22303,N_22045);
nor U26913 (N_26913,N_21404,N_23234);
nor U26914 (N_26914,N_22100,N_22365);
xnor U26915 (N_26915,N_21076,N_22895);
nand U26916 (N_26916,N_21880,N_22348);
xor U26917 (N_26917,N_23660,N_22471);
xnor U26918 (N_26918,N_21906,N_21493);
nor U26919 (N_26919,N_22262,N_21913);
or U26920 (N_26920,N_21338,N_22023);
nand U26921 (N_26921,N_23942,N_23218);
nand U26922 (N_26922,N_21175,N_22887);
or U26923 (N_26923,N_23160,N_21459);
xor U26924 (N_26924,N_22000,N_23931);
or U26925 (N_26925,N_23377,N_23412);
and U26926 (N_26926,N_23702,N_23807);
or U26927 (N_26927,N_22220,N_22862);
nor U26928 (N_26928,N_21595,N_21209);
xor U26929 (N_26929,N_22175,N_21807);
nor U26930 (N_26930,N_23193,N_23669);
or U26931 (N_26931,N_22153,N_23025);
nand U26932 (N_26932,N_23370,N_23375);
nor U26933 (N_26933,N_23326,N_23837);
or U26934 (N_26934,N_21866,N_23981);
nand U26935 (N_26935,N_21841,N_21867);
xnor U26936 (N_26936,N_22005,N_23775);
or U26937 (N_26937,N_21357,N_21609);
xnor U26938 (N_26938,N_23359,N_23647);
nand U26939 (N_26939,N_22247,N_21494);
and U26940 (N_26940,N_21940,N_22667);
and U26941 (N_26941,N_21570,N_22958);
xnor U26942 (N_26942,N_22093,N_22527);
xor U26943 (N_26943,N_22948,N_22807);
nor U26944 (N_26944,N_21726,N_21170);
nor U26945 (N_26945,N_23395,N_21325);
or U26946 (N_26946,N_22123,N_21361);
nand U26947 (N_26947,N_21134,N_21529);
xnor U26948 (N_26948,N_22033,N_21003);
and U26949 (N_26949,N_21395,N_21777);
or U26950 (N_26950,N_22195,N_22153);
nor U26951 (N_26951,N_22704,N_21952);
or U26952 (N_26952,N_22529,N_21204);
and U26953 (N_26953,N_22075,N_23550);
xor U26954 (N_26954,N_23627,N_21396);
or U26955 (N_26955,N_23036,N_21637);
and U26956 (N_26956,N_21436,N_23916);
and U26957 (N_26957,N_23535,N_22342);
and U26958 (N_26958,N_23322,N_21775);
or U26959 (N_26959,N_22186,N_21001);
xor U26960 (N_26960,N_22886,N_22671);
and U26961 (N_26961,N_21410,N_21461);
or U26962 (N_26962,N_23975,N_22699);
or U26963 (N_26963,N_22720,N_22924);
nand U26964 (N_26964,N_23627,N_21969);
xor U26965 (N_26965,N_23212,N_23455);
or U26966 (N_26966,N_23599,N_23793);
or U26967 (N_26967,N_22760,N_21227);
nor U26968 (N_26968,N_22455,N_22180);
nor U26969 (N_26969,N_21340,N_23760);
xnor U26970 (N_26970,N_23890,N_21862);
and U26971 (N_26971,N_22660,N_21382);
nor U26972 (N_26972,N_21021,N_22871);
or U26973 (N_26973,N_23583,N_23853);
nor U26974 (N_26974,N_21115,N_22047);
nor U26975 (N_26975,N_22634,N_22369);
nor U26976 (N_26976,N_21053,N_22479);
and U26977 (N_26977,N_23646,N_21148);
nand U26978 (N_26978,N_21132,N_23913);
nor U26979 (N_26979,N_21078,N_21930);
or U26980 (N_26980,N_23599,N_22787);
nand U26981 (N_26981,N_23735,N_21480);
or U26982 (N_26982,N_21509,N_21268);
and U26983 (N_26983,N_21682,N_23181);
nand U26984 (N_26984,N_21985,N_22052);
or U26985 (N_26985,N_22637,N_22517);
xor U26986 (N_26986,N_21816,N_23349);
nor U26987 (N_26987,N_22410,N_23832);
and U26988 (N_26988,N_21492,N_23031);
nor U26989 (N_26989,N_21661,N_22798);
xor U26990 (N_26990,N_22638,N_22126);
nor U26991 (N_26991,N_23082,N_21637);
nand U26992 (N_26992,N_22373,N_21448);
and U26993 (N_26993,N_22105,N_23500);
nand U26994 (N_26994,N_21582,N_23776);
xnor U26995 (N_26995,N_21587,N_21435);
nand U26996 (N_26996,N_23287,N_22034);
nor U26997 (N_26997,N_22991,N_22891);
or U26998 (N_26998,N_22740,N_23536);
or U26999 (N_26999,N_22848,N_21214);
or U27000 (N_27000,N_25495,N_24265);
or U27001 (N_27001,N_26482,N_25979);
xnor U27002 (N_27002,N_25890,N_26726);
and U27003 (N_27003,N_26879,N_24079);
nand U27004 (N_27004,N_25068,N_24012);
nand U27005 (N_27005,N_24056,N_26074);
or U27006 (N_27006,N_25598,N_26258);
nand U27007 (N_27007,N_26041,N_26572);
nand U27008 (N_27008,N_25444,N_26913);
and U27009 (N_27009,N_26903,N_25707);
xor U27010 (N_27010,N_26861,N_26246);
nor U27011 (N_27011,N_25583,N_24368);
or U27012 (N_27012,N_25347,N_24468);
or U27013 (N_27013,N_26198,N_24699);
or U27014 (N_27014,N_26576,N_26354);
or U27015 (N_27015,N_24868,N_25298);
or U27016 (N_27016,N_24382,N_24075);
nand U27017 (N_27017,N_25006,N_24181);
xor U27018 (N_27018,N_24131,N_24034);
xor U27019 (N_27019,N_24830,N_25261);
or U27020 (N_27020,N_26128,N_25763);
xnor U27021 (N_27021,N_24527,N_25791);
nand U27022 (N_27022,N_25287,N_25742);
or U27023 (N_27023,N_26611,N_26029);
nand U27024 (N_27024,N_25722,N_25281);
or U27025 (N_27025,N_24543,N_26118);
xor U27026 (N_27026,N_26713,N_26057);
xnor U27027 (N_27027,N_24727,N_25810);
nor U27028 (N_27028,N_26729,N_26515);
and U27029 (N_27029,N_24748,N_24348);
xnor U27030 (N_27030,N_25839,N_26504);
nand U27031 (N_27031,N_25361,N_26011);
or U27032 (N_27032,N_26626,N_26380);
and U27033 (N_27033,N_26648,N_25512);
or U27034 (N_27034,N_25228,N_25842);
and U27035 (N_27035,N_26831,N_25715);
and U27036 (N_27036,N_24182,N_26667);
nor U27037 (N_27037,N_26015,N_24927);
and U27038 (N_27038,N_26534,N_24253);
nor U27039 (N_27039,N_26071,N_26953);
xnor U27040 (N_27040,N_26502,N_24163);
and U27041 (N_27041,N_25573,N_26428);
nor U27042 (N_27042,N_25808,N_26523);
xor U27043 (N_27043,N_24807,N_24299);
and U27044 (N_27044,N_26881,N_24824);
nor U27045 (N_27045,N_24027,N_25067);
xnor U27046 (N_27046,N_24551,N_26890);
and U27047 (N_27047,N_24890,N_26250);
or U27048 (N_27048,N_24135,N_26751);
or U27049 (N_27049,N_25792,N_24115);
xnor U27050 (N_27050,N_24975,N_24808);
nand U27051 (N_27051,N_25472,N_26708);
and U27052 (N_27052,N_26538,N_26429);
or U27053 (N_27053,N_26349,N_26750);
nand U27054 (N_27054,N_26860,N_25295);
and U27055 (N_27055,N_24255,N_24710);
nand U27056 (N_27056,N_24719,N_26093);
and U27057 (N_27057,N_24603,N_24610);
nor U27058 (N_27058,N_26760,N_24838);
xor U27059 (N_27059,N_25857,N_26477);
xor U27060 (N_27060,N_24871,N_26937);
xnor U27061 (N_27061,N_24567,N_26604);
nor U27062 (N_27062,N_24682,N_26674);
and U27063 (N_27063,N_24070,N_25299);
xnor U27064 (N_27064,N_25334,N_26253);
and U27065 (N_27065,N_24134,N_24385);
nor U27066 (N_27066,N_25868,N_25343);
and U27067 (N_27067,N_25003,N_24829);
xnor U27068 (N_27068,N_24498,N_24978);
nand U27069 (N_27069,N_25827,N_25273);
xnor U27070 (N_27070,N_26509,N_25059);
nor U27071 (N_27071,N_24519,N_24338);
and U27072 (N_27072,N_24760,N_24203);
or U27073 (N_27073,N_24640,N_25655);
and U27074 (N_27074,N_26863,N_24129);
xor U27075 (N_27075,N_24305,N_24965);
nor U27076 (N_27076,N_26302,N_25706);
nand U27077 (N_27077,N_26641,N_26783);
nand U27078 (N_27078,N_24678,N_24683);
nor U27079 (N_27079,N_25734,N_25383);
and U27080 (N_27080,N_25253,N_24314);
and U27081 (N_27081,N_24806,N_25449);
xnor U27082 (N_27082,N_24423,N_26470);
nand U27083 (N_27083,N_26615,N_25740);
xnor U27084 (N_27084,N_25889,N_26151);
and U27085 (N_27085,N_25112,N_25367);
nor U27086 (N_27086,N_26837,N_26418);
nand U27087 (N_27087,N_25799,N_26653);
nand U27088 (N_27088,N_26218,N_26711);
nor U27089 (N_27089,N_25242,N_25524);
xnor U27090 (N_27090,N_26787,N_24251);
and U27091 (N_27091,N_26035,N_25082);
xnor U27092 (N_27092,N_24502,N_25352);
xnor U27093 (N_27093,N_24529,N_26695);
nor U27094 (N_27094,N_25030,N_25038);
nand U27095 (N_27095,N_24096,N_25263);
nor U27096 (N_27096,N_24036,N_24189);
xor U27097 (N_27097,N_25834,N_26191);
nor U27098 (N_27098,N_24483,N_24749);
nand U27099 (N_27099,N_26951,N_25507);
xor U27100 (N_27100,N_25438,N_24404);
and U27101 (N_27101,N_24509,N_25234);
xor U27102 (N_27102,N_25131,N_24648);
nor U27103 (N_27103,N_25618,N_26047);
nand U27104 (N_27104,N_26257,N_24414);
nor U27105 (N_27105,N_26716,N_26275);
nor U27106 (N_27106,N_24615,N_24173);
and U27107 (N_27107,N_25136,N_25167);
or U27108 (N_27108,N_24174,N_26053);
or U27109 (N_27109,N_25206,N_26402);
or U27110 (N_27110,N_26875,N_24779);
xor U27111 (N_27111,N_25117,N_24153);
or U27112 (N_27112,N_25757,N_25159);
xnor U27113 (N_27113,N_24508,N_25798);
and U27114 (N_27114,N_24371,N_26663);
nand U27115 (N_27115,N_25019,N_25670);
xor U27116 (N_27116,N_25677,N_24039);
or U27117 (N_27117,N_25671,N_24478);
nand U27118 (N_27118,N_25650,N_24561);
or U27119 (N_27119,N_25959,N_26812);
xnor U27120 (N_27120,N_26274,N_25044);
nand U27121 (N_27121,N_24815,N_26201);
nor U27122 (N_27122,N_25966,N_26019);
xnor U27123 (N_27123,N_25851,N_25571);
nand U27124 (N_27124,N_25313,N_26807);
xnor U27125 (N_27125,N_25812,N_24292);
and U27126 (N_27126,N_26025,N_26455);
and U27127 (N_27127,N_25364,N_26329);
or U27128 (N_27128,N_25631,N_25619);
nor U27129 (N_27129,N_25328,N_26487);
nand U27130 (N_27130,N_24624,N_25991);
xnor U27131 (N_27131,N_26578,N_24452);
or U27132 (N_27132,N_26671,N_24739);
nor U27133 (N_27133,N_26795,N_24982);
and U27134 (N_27134,N_26055,N_26008);
nand U27135 (N_27135,N_25119,N_25271);
and U27136 (N_27136,N_26271,N_24457);
nor U27137 (N_27137,N_26330,N_25908);
nand U27138 (N_27138,N_25770,N_26901);
and U27139 (N_27139,N_26227,N_24381);
or U27140 (N_27140,N_26410,N_26654);
nand U27141 (N_27141,N_25559,N_24121);
or U27142 (N_27142,N_26762,N_26683);
and U27143 (N_27143,N_24187,N_25245);
xor U27144 (N_27144,N_24392,N_26232);
or U27145 (N_27145,N_25033,N_25621);
nand U27146 (N_27146,N_26252,N_25374);
or U27147 (N_27147,N_26338,N_25375);
xor U27148 (N_27148,N_24107,N_25874);
nor U27149 (N_27149,N_24432,N_26318);
nor U27150 (N_27150,N_26507,N_26844);
nand U27151 (N_27151,N_24102,N_24016);
and U27152 (N_27152,N_25041,N_25321);
nand U27153 (N_27153,N_24471,N_24198);
nand U27154 (N_27154,N_26520,N_24104);
or U27155 (N_27155,N_24084,N_26981);
or U27156 (N_27156,N_25589,N_26183);
xnor U27157 (N_27157,N_24332,N_25310);
and U27158 (N_27158,N_24114,N_24233);
nand U27159 (N_27159,N_25915,N_24585);
and U27160 (N_27160,N_24670,N_26173);
or U27161 (N_27161,N_26585,N_24903);
nand U27162 (N_27162,N_25013,N_26289);
xor U27163 (N_27163,N_26744,N_25341);
xnor U27164 (N_27164,N_26174,N_26301);
nor U27165 (N_27165,N_24178,N_25630);
nand U27166 (N_27166,N_25828,N_25262);
xor U27167 (N_27167,N_26423,N_26249);
or U27168 (N_27168,N_24499,N_24440);
nor U27169 (N_27169,N_25846,N_24883);
nand U27170 (N_27170,N_26606,N_25468);
nand U27171 (N_27171,N_25578,N_25932);
nand U27172 (N_27172,N_26133,N_26188);
or U27173 (N_27173,N_24594,N_24261);
and U27174 (N_27174,N_24571,N_24298);
and U27175 (N_27175,N_24325,N_24554);
nand U27176 (N_27176,N_26153,N_26833);
nand U27177 (N_27177,N_26521,N_24335);
or U27178 (N_27178,N_26152,N_25405);
or U27179 (N_27179,N_25668,N_26048);
xor U27180 (N_27180,N_26925,N_25554);
nor U27181 (N_27181,N_26313,N_24535);
or U27182 (N_27182,N_26669,N_25066);
xnor U27183 (N_27183,N_25888,N_25777);
xor U27184 (N_27184,N_25442,N_26493);
and U27185 (N_27185,N_24977,N_26541);
nand U27186 (N_27186,N_25431,N_24281);
and U27187 (N_27187,N_25325,N_25489);
and U27188 (N_27188,N_25535,N_24328);
and U27189 (N_27189,N_25930,N_26827);
nand U27190 (N_27190,N_25766,N_26239);
xnor U27191 (N_27191,N_26316,N_25698);
xnor U27192 (N_27192,N_25771,N_24168);
xor U27193 (N_27193,N_26290,N_24304);
nand U27194 (N_27194,N_26341,N_26333);
xnor U27195 (N_27195,N_24773,N_26122);
xor U27196 (N_27196,N_25071,N_24176);
nor U27197 (N_27197,N_24028,N_24329);
or U27198 (N_27198,N_25543,N_25940);
nand U27199 (N_27199,N_24920,N_26524);
and U27200 (N_27200,N_26883,N_24844);
nor U27201 (N_27201,N_24800,N_25807);
nor U27202 (N_27202,N_25413,N_25396);
or U27203 (N_27203,N_24525,N_24949);
or U27204 (N_27204,N_25390,N_24081);
nand U27205 (N_27205,N_26510,N_26506);
and U27206 (N_27206,N_25258,N_25362);
and U27207 (N_27207,N_24043,N_26596);
xor U27208 (N_27208,N_26426,N_24132);
and U27209 (N_27209,N_24149,N_24072);
or U27210 (N_27210,N_26649,N_25606);
xnor U27211 (N_27211,N_26251,N_26207);
or U27212 (N_27212,N_24130,N_24848);
xor U27213 (N_27213,N_24677,N_24395);
nor U27214 (N_27214,N_26893,N_25899);
xor U27215 (N_27215,N_24767,N_24405);
and U27216 (N_27216,N_24972,N_26052);
nor U27217 (N_27217,N_26868,N_25199);
or U27218 (N_27218,N_26453,N_25229);
or U27219 (N_27219,N_26384,N_25982);
xnor U27220 (N_27220,N_24256,N_26836);
xor U27221 (N_27221,N_25613,N_26365);
or U27222 (N_27222,N_26556,N_25469);
xnor U27223 (N_27223,N_26392,N_25661);
xnor U27224 (N_27224,N_24127,N_24490);
and U27225 (N_27225,N_25702,N_24315);
xor U27226 (N_27226,N_25214,N_24518);
nand U27227 (N_27227,N_26554,N_26832);
nor U27228 (N_27228,N_25793,N_24420);
or U27229 (N_27229,N_25765,N_26593);
and U27230 (N_27230,N_24960,N_26573);
xnor U27231 (N_27231,N_24961,N_26226);
nor U27232 (N_27232,N_26267,N_25829);
nor U27233 (N_27233,N_26344,N_25703);
or U27234 (N_27234,N_24901,N_24796);
and U27235 (N_27235,N_26033,N_25759);
and U27236 (N_27236,N_25337,N_26007);
nand U27237 (N_27237,N_25219,N_24629);
xor U27238 (N_27238,N_24186,N_26871);
nor U27239 (N_27239,N_26602,N_26517);
nor U27240 (N_27240,N_25173,N_26772);
and U27241 (N_27241,N_26739,N_25737);
nor U27242 (N_27242,N_24126,N_24996);
and U27243 (N_27243,N_26437,N_25290);
or U27244 (N_27244,N_26874,N_26245);
nand U27245 (N_27245,N_25461,N_24723);
and U27246 (N_27246,N_25397,N_25539);
and U27247 (N_27247,N_26206,N_24826);
nor U27248 (N_27248,N_24358,N_24513);
or U27249 (N_27249,N_25609,N_26377);
or U27250 (N_27250,N_26081,N_24409);
xor U27251 (N_27251,N_26968,N_25804);
nand U27252 (N_27252,N_24985,N_25678);
nand U27253 (N_27253,N_26622,N_25045);
nand U27254 (N_27254,N_26414,N_25443);
nand U27255 (N_27255,N_25756,N_26818);
and U27256 (N_27256,N_26105,N_25648);
and U27257 (N_27257,N_26297,N_25917);
and U27258 (N_27258,N_26389,N_25533);
nor U27259 (N_27259,N_24696,N_24363);
or U27260 (N_27260,N_26940,N_25014);
xor U27261 (N_27261,N_25855,N_26401);
and U27262 (N_27262,N_26679,N_26457);
and U27263 (N_27263,N_24387,N_24744);
or U27264 (N_27264,N_24042,N_26955);
nand U27265 (N_27265,N_25028,N_24133);
and U27266 (N_27266,N_25949,N_26415);
nand U27267 (N_27267,N_25815,N_24974);
or U27268 (N_27268,N_25169,N_26677);
xnor U27269 (N_27269,N_26830,N_26490);
nand U27270 (N_27270,N_25976,N_26031);
nand U27271 (N_27271,N_26963,N_25046);
nand U27272 (N_27272,N_24501,N_24422);
or U27273 (N_27273,N_25197,N_26793);
xnor U27274 (N_27274,N_26138,N_25717);
xnor U27275 (N_27275,N_24263,N_24419);
xnor U27276 (N_27276,N_25089,N_26001);
xnor U27277 (N_27277,N_24538,N_26018);
nand U27278 (N_27278,N_24896,N_25754);
nor U27279 (N_27279,N_24520,N_26568);
or U27280 (N_27280,N_24865,N_24879);
xnor U27281 (N_27281,N_24786,N_26975);
nor U27282 (N_27282,N_24221,N_25723);
and U27283 (N_27283,N_26806,N_25638);
and U27284 (N_27284,N_25674,N_25731);
and U27285 (N_27285,N_25526,N_24078);
or U27286 (N_27286,N_25482,N_26042);
xnor U27287 (N_27287,N_25651,N_24763);
and U27288 (N_27288,N_26355,N_26110);
nand U27289 (N_27289,N_26966,N_26984);
and U27290 (N_27290,N_25213,N_25433);
and U27291 (N_27291,N_26592,N_26906);
xnor U27292 (N_27292,N_26148,N_24033);
nor U27293 (N_27293,N_26815,N_24526);
nor U27294 (N_27294,N_26030,N_24546);
nor U27295 (N_27295,N_26911,N_25988);
and U27296 (N_27296,N_25487,N_26443);
nand U27297 (N_27297,N_26723,N_25530);
nor U27298 (N_27298,N_24522,N_24536);
nor U27299 (N_27299,N_26104,N_24946);
nand U27300 (N_27300,N_26575,N_24435);
or U27301 (N_27301,N_24475,N_25087);
nor U27302 (N_27302,N_24784,N_24447);
xor U27303 (N_27303,N_26814,N_24616);
or U27304 (N_27304,N_26917,N_25106);
nand U27305 (N_27305,N_24429,N_24852);
nand U27306 (N_27306,N_26303,N_25975);
and U27307 (N_27307,N_26876,N_24403);
and U27308 (N_27308,N_25574,N_26235);
nor U27309 (N_27309,N_25065,N_24792);
nand U27310 (N_27310,N_24714,N_26887);
and U27311 (N_27311,N_26977,N_24738);
or U27312 (N_27312,N_25994,N_24321);
or U27313 (N_27313,N_24354,N_24040);
nor U27314 (N_27314,N_26092,N_25615);
nor U27315 (N_27315,N_26186,N_26168);
nand U27316 (N_27316,N_26741,N_26149);
and U27317 (N_27317,N_24038,N_26096);
or U27318 (N_27318,N_24679,N_24228);
nand U27319 (N_27319,N_24359,N_25653);
and U27320 (N_27320,N_24365,N_24811);
and U27321 (N_27321,N_26731,N_24476);
nor U27322 (N_27322,N_24416,N_24512);
nor U27323 (N_27323,N_26195,N_25816);
nor U27324 (N_27324,N_26135,N_24971);
nor U27325 (N_27325,N_26439,N_24572);
or U27326 (N_27326,N_24924,N_26948);
and U27327 (N_27327,N_26113,N_25686);
nand U27328 (N_27328,N_24391,N_24524);
nor U27329 (N_27329,N_25556,N_26532);
nand U27330 (N_27330,N_25254,N_26801);
xnor U27331 (N_27331,N_26869,N_26283);
and U27332 (N_27332,N_24817,N_24073);
xor U27333 (N_27333,N_25177,N_26175);
xnor U27334 (N_27334,N_25641,N_26537);
nor U27335 (N_27335,N_26447,N_24492);
nor U27336 (N_27336,N_25241,N_26411);
nor U27337 (N_27337,N_24477,N_25185);
xor U27338 (N_27338,N_25788,N_24148);
and U27339 (N_27339,N_25212,N_26407);
nor U27340 (N_27340,N_25342,N_25523);
nand U27341 (N_27341,N_24407,N_26928);
nor U27342 (N_27342,N_24374,N_24230);
or U27343 (N_27343,N_24649,N_24421);
nand U27344 (N_27344,N_25264,N_24367);
nand U27345 (N_27345,N_26114,N_25555);
nand U27346 (N_27346,N_25531,N_25938);
or U27347 (N_27347,N_24757,N_25164);
xnor U27348 (N_27348,N_25905,N_26758);
and U27349 (N_27349,N_26381,N_25399);
or U27350 (N_27350,N_25079,N_25121);
nand U27351 (N_27351,N_24532,N_26422);
nor U27352 (N_27352,N_25259,N_24962);
or U27353 (N_27353,N_25503,N_24582);
or U27354 (N_27354,N_24689,N_24847);
nor U27355 (N_27355,N_25680,N_24915);
and U27356 (N_27356,N_26970,N_26637);
nand U27357 (N_27357,N_25595,N_25860);
and U27358 (N_27358,N_26542,N_26165);
or U27359 (N_27359,N_24930,N_25639);
nand U27360 (N_27360,N_26260,N_24346);
xor U27361 (N_27361,N_26369,N_25200);
nor U27362 (N_27362,N_26942,N_25158);
xor U27363 (N_27363,N_25201,N_26560);
nor U27364 (N_27364,N_25467,N_25353);
or U27365 (N_27365,N_26718,N_24283);
xor U27366 (N_27366,N_24711,N_24236);
xor U27367 (N_27367,N_26205,N_24243);
xnor U27368 (N_27368,N_24832,N_26213);
nand U27369 (N_27369,N_25062,N_24528);
or U27370 (N_27370,N_26296,N_25351);
nor U27371 (N_27371,N_24030,N_24663);
xor U27372 (N_27372,N_24644,N_25646);
nor U27373 (N_27373,N_26090,N_24495);
or U27374 (N_27374,N_24287,N_26681);
or U27375 (N_27375,N_25499,N_24294);
nor U27376 (N_27376,N_25711,N_24336);
or U27377 (N_27377,N_24445,N_25752);
nand U27378 (N_27378,N_25802,N_25775);
nand U27379 (N_27379,N_25492,N_25780);
xor U27380 (N_27380,N_25854,N_26310);
or U27381 (N_27381,N_25502,N_24545);
nand U27382 (N_27382,N_26347,N_25563);
and U27383 (N_27383,N_24768,N_24057);
nor U27384 (N_27384,N_24692,N_25830);
or U27385 (N_27385,N_26036,N_25505);
nand U27386 (N_27386,N_25773,N_24631);
nor U27387 (N_27387,N_26676,N_25863);
and U27388 (N_27388,N_26220,N_26494);
or U27389 (N_27389,N_25001,N_26489);
xnor U27390 (N_27390,N_26027,N_24238);
and U27391 (N_27391,N_24245,N_26706);
and U27392 (N_27392,N_25251,N_25260);
xnor U27393 (N_27393,N_24100,N_24618);
nor U27394 (N_27394,N_24280,N_25268);
and U27395 (N_27395,N_25144,N_25948);
or U27396 (N_27396,N_26129,N_24825);
and U27397 (N_27397,N_25952,N_24608);
or U27398 (N_27398,N_25382,N_26550);
nand U27399 (N_27399,N_25542,N_26399);
nand U27400 (N_27400,N_24850,N_24693);
nand U27401 (N_27401,N_26752,N_25823);
and U27402 (N_27402,N_26281,N_26583);
nand U27403 (N_27403,N_26864,N_26800);
nand U27404 (N_27404,N_26343,N_24576);
and U27405 (N_27405,N_25017,N_24145);
nor U27406 (N_27406,N_25963,N_25644);
or U27407 (N_27407,N_25772,N_24482);
xor U27408 (N_27408,N_26819,N_26900);
nor U27409 (N_27409,N_24741,N_24019);
nor U27410 (N_27410,N_26337,N_25822);
nor U27411 (N_27411,N_26761,N_24171);
nor U27412 (N_27412,N_24555,N_24886);
or U27413 (N_27413,N_26780,N_25824);
nor U27414 (N_27414,N_24899,N_24065);
or U27415 (N_27415,N_24088,N_25925);
xnor U27416 (N_27416,N_24958,N_24339);
nor U27417 (N_27417,N_26350,N_26046);
xnor U27418 (N_27418,N_24667,N_25695);
and U27419 (N_27419,N_25285,N_26432);
nand U27420 (N_27420,N_26999,N_25034);
nor U27421 (N_27421,N_24559,N_24870);
nor U27422 (N_27422,N_24241,N_26087);
nand U27423 (N_27423,N_24352,N_25729);
xor U27424 (N_27424,N_26370,N_25256);
xor U27425 (N_27425,N_24776,N_25247);
or U27426 (N_27426,N_25728,N_25162);
nand U27427 (N_27427,N_26088,N_26228);
and U27428 (N_27428,N_24970,N_25377);
and U27429 (N_27429,N_26024,N_26987);
or U27430 (N_27430,N_24681,N_25995);
and U27431 (N_27431,N_25048,N_26768);
or U27432 (N_27432,N_24628,N_25453);
nand U27433 (N_27433,N_25782,N_26898);
or U27434 (N_27434,N_24595,N_26063);
nand U27435 (N_27435,N_24976,N_24231);
xnor U27436 (N_27436,N_26775,N_24751);
or U27437 (N_27437,N_25480,N_25047);
or U27438 (N_27438,N_24276,N_26277);
xor U27439 (N_27439,N_26485,N_25231);
or U27440 (N_27440,N_26180,N_25694);
nand U27441 (N_27441,N_25446,N_24853);
xor U27442 (N_27442,N_24914,N_25712);
or U27443 (N_27443,N_25008,N_26878);
or U27444 (N_27444,N_24152,N_24783);
nand U27445 (N_27445,N_25867,N_24735);
xnor U27446 (N_27446,N_25393,N_25277);
and U27447 (N_27447,N_25588,N_26748);
nand U27448 (N_27448,N_25244,N_25887);
nor U27449 (N_27449,N_25274,N_24918);
xnor U27450 (N_27450,N_24099,N_24717);
nor U27451 (N_27451,N_26625,N_25276);
and U27452 (N_27452,N_25416,N_26311);
xnor U27453 (N_27453,N_24606,N_25898);
xnor U27454 (N_27454,N_26460,N_26295);
or U27455 (N_27455,N_24156,N_25525);
and U27456 (N_27456,N_25768,N_26442);
nor U27457 (N_27457,N_24657,N_25983);
and U27458 (N_27458,N_25474,N_25660);
or U27459 (N_27459,N_25818,N_24882);
or U27460 (N_27460,N_25892,N_24647);
or U27461 (N_27461,N_26581,N_26644);
xor U27462 (N_27462,N_25497,N_24664);
nor U27463 (N_27463,N_25123,N_26373);
or U27464 (N_27464,N_25369,N_25881);
and U27465 (N_27465,N_24810,N_26111);
or U27466 (N_27466,N_24400,N_26687);
nor U27467 (N_27467,N_26705,N_24630);
xor U27468 (N_27468,N_25430,N_26777);
xor U27469 (N_27469,N_24531,N_26853);
nor U27470 (N_27470,N_26527,N_24269);
nand U27471 (N_27471,N_24973,N_26382);
xor U27472 (N_27472,N_24398,N_24802);
nand U27473 (N_27473,N_24345,N_25738);
or U27474 (N_27474,N_26569,N_25378);
nor U27475 (N_27475,N_25488,N_24430);
or U27476 (N_27476,N_24257,N_26476);
nor U27477 (N_27477,N_26935,N_25186);
nor U27478 (N_27478,N_26745,N_26995);
and U27479 (N_27479,N_26454,N_26371);
or U27480 (N_27480,N_25819,N_24399);
or U27481 (N_27481,N_24983,N_26244);
nand U27482 (N_27482,N_24089,N_24922);
xnor U27483 (N_27483,N_24705,N_25157);
nand U27484 (N_27484,N_25811,N_25004);
and U27485 (N_27485,N_25088,N_25408);
and U27486 (N_27486,N_25324,N_26077);
nor U27487 (N_27487,N_25882,N_25081);
nand U27488 (N_27488,N_24845,N_24885);
nand U27489 (N_27489,N_26620,N_26279);
and U27490 (N_27490,N_24061,N_26997);
and U27491 (N_27491,N_25189,N_24260);
and U27492 (N_27492,N_25292,N_25955);
nor U27493 (N_27493,N_25180,N_26693);
xnor U27494 (N_27494,N_24963,N_25101);
and U27495 (N_27495,N_26689,N_25758);
xnor U27496 (N_27496,N_25312,N_26192);
nand U27497 (N_27497,N_24942,N_25871);
nor U27498 (N_27498,N_26501,N_25165);
nand U27499 (N_27499,N_26967,N_26664);
and U27500 (N_27500,N_24436,N_25091);
xor U27501 (N_27501,N_25308,N_24840);
xor U27502 (N_27502,N_25813,N_25070);
or U27503 (N_27503,N_24510,N_25891);
xnor U27504 (N_27504,N_25724,N_24362);
nor U27505 (N_27505,N_25211,N_25900);
nand U27506 (N_27506,N_25072,N_26699);
xor U27507 (N_27507,N_24376,N_25597);
or U27508 (N_27508,N_25509,N_25400);
nand U27509 (N_27509,N_24434,N_26466);
nand U27510 (N_27510,N_25585,N_26431);
and U27511 (N_27511,N_26385,N_25005);
nand U27512 (N_27512,N_25175,N_25942);
and U27513 (N_27513,N_25354,N_24085);
nand U27514 (N_27514,N_25370,N_24316);
and U27515 (N_27515,N_24864,N_25465);
nand U27516 (N_27516,N_24583,N_25429);
xor U27517 (N_27517,N_25395,N_26945);
nor U27518 (N_27518,N_25849,N_25269);
nor U27519 (N_27519,N_26789,N_26850);
nor U27520 (N_27520,N_25187,N_26496);
and U27521 (N_27521,N_26714,N_25879);
and U27522 (N_27522,N_24787,N_25055);
nor U27523 (N_27523,N_26769,N_26471);
xor U27524 (N_27524,N_26960,N_24433);
nor U27525 (N_27525,N_26662,N_24122);
or U27526 (N_27526,N_26609,N_26395);
nor U27527 (N_27527,N_25394,N_24721);
or U27528 (N_27528,N_24921,N_25669);
nand U27529 (N_27529,N_25074,N_26811);
and U27530 (N_27530,N_26998,N_24394);
xnor U27531 (N_27531,N_24195,N_24003);
nor U27532 (N_27532,N_26949,N_25239);
or U27533 (N_27533,N_25856,N_26266);
nor U27534 (N_27534,N_26782,N_24732);
nor U27535 (N_27535,N_24201,N_25331);
or U27536 (N_27536,N_26287,N_26242);
and U27537 (N_27537,N_25098,N_26131);
and U27538 (N_27538,N_24209,N_26388);
nor U27539 (N_27539,N_25108,N_24402);
and U27540 (N_27540,N_26557,N_24312);
nand U27541 (N_27541,N_24504,N_25697);
or U27542 (N_27542,N_24239,N_25454);
nand U27543 (N_27543,N_26808,N_26552);
or U27544 (N_27544,N_26056,N_26764);
xnor U27545 (N_27545,N_25414,N_26383);
and U27546 (N_27546,N_24226,N_26372);
and U27547 (N_27547,N_25944,N_26529);
nand U27548 (N_27548,N_25985,N_25913);
or U27549 (N_27549,N_24855,N_25594);
or U27550 (N_27550,N_26736,N_26545);
xor U27551 (N_27551,N_26276,N_24074);
or U27552 (N_27552,N_24472,N_25387);
nor U27553 (N_27553,N_24247,N_25886);
xor U27554 (N_27554,N_26364,N_26095);
xnor U27555 (N_27555,N_25225,N_26100);
or U27556 (N_27556,N_25974,N_26091);
and U27557 (N_27557,N_24698,N_25684);
nand U27558 (N_27558,N_26512,N_24293);
and U27559 (N_27559,N_25419,N_26680);
nor U27560 (N_27560,N_25778,N_24736);
and U27561 (N_27561,N_25478,N_26003);
and U27562 (N_27562,N_24386,N_26156);
nor U27563 (N_27563,N_26044,N_24289);
nand U27564 (N_27564,N_26479,N_25872);
nor U27565 (N_27565,N_26934,N_26743);
nand U27566 (N_27566,N_25923,N_26375);
nand U27567 (N_27567,N_26441,N_24925);
xnor U27568 (N_27568,N_25491,N_26712);
and U27569 (N_27569,N_26264,N_24484);
nand U27570 (N_27570,N_26895,N_26914);
nor U27571 (N_27571,N_25667,N_24177);
nand U27572 (N_27572,N_24047,N_25859);
nand U27573 (N_27573,N_25208,N_26254);
or U27574 (N_27574,N_24892,N_25953);
xor U27575 (N_27575,N_26992,N_24302);
xor U27576 (N_27576,N_25662,N_24789);
and U27577 (N_27577,N_26394,N_24138);
nand U27578 (N_27578,N_26553,N_25386);
and U27579 (N_27579,N_25226,N_25205);
xor U27580 (N_27580,N_26954,N_26786);
and U27581 (N_27581,N_26624,N_26549);
and U27582 (N_27582,N_24474,N_25876);
nor U27583 (N_27583,N_26952,N_26503);
nand U27584 (N_27584,N_25163,N_25010);
nand U27585 (N_27585,N_26217,N_26941);
xnor U27586 (N_27586,N_26639,N_25023);
or U27587 (N_27587,N_25184,N_26846);
nor U27588 (N_27588,N_24599,N_25753);
nand U27589 (N_27589,N_25602,N_25977);
xor U27590 (N_27590,N_24712,N_25906);
or U27591 (N_27591,N_25306,N_25025);
xor U27592 (N_27592,N_26614,N_26378);
nor U27593 (N_27593,N_26673,N_24311);
nor U27594 (N_27594,N_24388,N_26256);
or U27595 (N_27595,N_26690,N_26498);
nand U27596 (N_27596,N_25452,N_25116);
nand U27597 (N_27597,N_24939,N_24425);
or U27598 (N_27598,N_25848,N_25250);
nand U27599 (N_27599,N_24116,N_26158);
or U27600 (N_27600,N_25565,N_25666);
nor U27601 (N_27601,N_26005,N_26017);
nand U27602 (N_27602,N_25035,N_24022);
or U27603 (N_27603,N_26884,N_24745);
xor U27604 (N_27604,N_25086,N_25633);
xnor U27605 (N_27605,N_24756,N_24093);
xor U27606 (N_27606,N_24690,N_26064);
and U27607 (N_27607,N_24645,N_25562);
and U27608 (N_27608,N_25950,N_26229);
xor U27609 (N_27609,N_25767,N_25659);
nor U27610 (N_27610,N_26406,N_25645);
xnor U27611 (N_27611,N_26665,N_25152);
and U27612 (N_27612,N_25100,N_24103);
nor U27613 (N_27613,N_24912,N_26514);
nor U27614 (N_27614,N_26894,N_26076);
nand U27615 (N_27615,N_26763,N_25128);
or U27616 (N_27616,N_24700,N_24212);
nor U27617 (N_27617,N_26464,N_24951);
nand U27618 (N_27618,N_25139,N_26317);
nand U27619 (N_27619,N_24244,N_26838);
or U27620 (N_27620,N_25385,N_26766);
nand U27621 (N_27621,N_24091,N_24943);
nor U27622 (N_27622,N_24916,N_25636);
nand U27623 (N_27623,N_24708,N_25805);
or U27624 (N_27624,N_26109,N_25368);
nand U27625 (N_27625,N_24734,N_25730);
xnor U27626 (N_27626,N_25240,N_24324);
xnor U27627 (N_27627,N_24688,N_25705);
nor U27628 (N_27628,N_26721,N_26136);
nor U27629 (N_27629,N_26284,N_24765);
nand U27630 (N_27630,N_24713,N_26430);
or U27631 (N_27631,N_25359,N_26616);
or U27632 (N_27632,N_26075,N_26140);
and U27633 (N_27633,N_26589,N_25996);
nand U27634 (N_27634,N_24884,N_25227);
nor U27635 (N_27635,N_24048,N_26822);
xor U27636 (N_27636,N_26849,N_26182);
nor U27637 (N_27637,N_26724,N_26518);
nand U27638 (N_27638,N_25617,N_26405);
nand U27639 (N_27639,N_26166,N_25693);
xor U27640 (N_27640,N_25713,N_26702);
or U27641 (N_27641,N_26886,N_26638);
nor U27642 (N_27642,N_25864,N_25785);
xor U27643 (N_27643,N_24507,N_24966);
xor U27644 (N_27644,N_24486,N_24308);
xor U27645 (N_27645,N_25420,N_24213);
nor U27646 (N_27646,N_24846,N_26234);
nor U27647 (N_27647,N_24701,N_26185);
and U27648 (N_27648,N_24533,N_24650);
and U27649 (N_27649,N_24347,N_26026);
nor U27650 (N_27650,N_24068,N_25806);
xnor U27651 (N_27651,N_24809,N_25870);
or U27652 (N_27652,N_24408,N_24364);
or U27653 (N_27653,N_24202,N_25110);
nor U27654 (N_27654,N_24790,N_26060);
and U27655 (N_27655,N_26916,N_24515);
nand U27656 (N_27656,N_25536,N_26920);
or U27657 (N_27657,N_24340,N_24503);
xor U27658 (N_27658,N_26255,N_24570);
nand U27659 (N_27659,N_24553,N_24170);
nand U27660 (N_27660,N_25147,N_26902);
nand U27661 (N_27661,N_26440,N_24858);
nand U27662 (N_27662,N_26603,N_25224);
nor U27663 (N_27663,N_26632,N_26661);
nand U27664 (N_27664,N_26134,N_24453);
nor U27665 (N_27665,N_24059,N_24550);
xor U27666 (N_27666,N_26610,N_24987);
and U27667 (N_27667,N_24199,N_25549);
nand U27668 (N_27668,N_25564,N_26468);
nand U27669 (N_27669,N_25097,N_25115);
or U27670 (N_27670,N_25275,N_26738);
xor U27671 (N_27671,N_26225,N_26320);
nand U27672 (N_27672,N_24207,N_26597);
and U27673 (N_27673,N_25538,N_25861);
nor U27674 (N_27674,N_25971,N_24083);
nor U27675 (N_27675,N_24706,N_24485);
and U27676 (N_27676,N_26709,N_24586);
or U27677 (N_27677,N_25140,N_26484);
nor U27678 (N_27678,N_24473,N_25789);
nand U27679 (N_27679,N_26334,N_24449);
xor U27680 (N_27680,N_26288,N_25056);
nand U27681 (N_27681,N_25349,N_25198);
or U27682 (N_27682,N_24632,N_25193);
or U27683 (N_27683,N_26599,N_25441);
xor U27684 (N_27684,N_25243,N_25457);
and U27685 (N_27685,N_26732,N_25357);
xor U27686 (N_27686,N_24589,N_24843);
xor U27687 (N_27687,N_26757,N_24834);
xnor U27688 (N_27688,N_26564,N_25272);
nor U27689 (N_27689,N_24569,N_24227);
nor U27690 (N_27690,N_25553,N_26571);
xor U27691 (N_27691,N_25418,N_25346);
nor U27692 (N_27692,N_25690,N_24197);
or U27693 (N_27693,N_24379,N_24095);
nor U27694 (N_27694,N_24052,N_26016);
and U27695 (N_27695,N_26269,N_26374);
nand U27696 (N_27696,N_26101,N_25462);
and U27697 (N_27697,N_25040,N_26642);
xor U27698 (N_27698,N_25150,N_25672);
xor U27699 (N_27699,N_24775,N_25914);
or U27700 (N_27700,N_24344,N_26474);
xor U27701 (N_27701,N_26700,N_25166);
and U27702 (N_27702,N_25642,N_24307);
nor U27703 (N_27703,N_26162,N_24248);
xnor U27704 (N_27704,N_24192,N_25043);
and U27705 (N_27705,N_25841,N_25125);
nand U27706 (N_27706,N_24990,N_26607);
and U27707 (N_27707,N_24087,N_24778);
nor U27708 (N_27708,N_26219,N_24439);
xnor U27709 (N_27709,N_26896,N_24493);
or U27710 (N_27710,N_25455,N_25363);
nor U27711 (N_27711,N_24355,N_25579);
nor U27712 (N_27712,N_26450,N_24300);
xnor U27713 (N_27713,N_24590,N_25154);
or U27714 (N_27714,N_26660,N_26522);
nor U27715 (N_27715,N_26839,N_25022);
nor U27716 (N_27716,N_24082,N_25335);
xor U27717 (N_27717,N_26929,N_24821);
nor U27718 (N_27718,N_26820,N_25989);
or U27719 (N_27719,N_25883,N_24933);
xnor U27720 (N_27720,N_25909,N_25391);
nand U27721 (N_27721,N_24557,N_26944);
or U27722 (N_27722,N_24098,N_26858);
or U27723 (N_27723,N_25451,N_24448);
nor U27724 (N_27724,N_24671,N_26691);
nor U27725 (N_27725,N_25632,N_26368);
nand U27726 (N_27726,N_25987,N_26433);
xnor U27727 (N_27727,N_26049,N_24639);
nor U27728 (N_27728,N_24356,N_24229);
nor U27729 (N_27729,N_26262,N_26958);
or U27730 (N_27730,N_24743,N_26636);
and U27731 (N_27731,N_25493,N_25837);
or U27732 (N_27732,N_26897,N_25787);
nor U27733 (N_27733,N_26852,N_26804);
nand U27734 (N_27734,N_26434,N_24957);
nand U27735 (N_27735,N_26448,N_25783);
or U27736 (N_27736,N_24271,N_25138);
nor U27737 (N_27737,N_24979,N_25540);
nor U27738 (N_27738,N_25009,N_26240);
nand U27739 (N_27739,N_26167,N_24905);
nand U27740 (N_27740,N_24902,N_26686);
nor U27741 (N_27741,N_26880,N_25440);
or U27742 (N_27742,N_26054,N_25278);
nor U27743 (N_27743,N_24794,N_26452);
or U27744 (N_27744,N_24175,N_26427);
nor U27745 (N_27745,N_25727,N_26835);
or U27746 (N_27746,N_25779,N_26196);
xnor U27747 (N_27747,N_25604,N_26212);
and U27748 (N_27748,N_24157,N_25450);
and U27749 (N_27749,N_26802,N_25485);
and U27750 (N_27750,N_24218,N_24437);
xor U27751 (N_27751,N_24428,N_26034);
nand U27752 (N_27752,N_24264,N_26986);
nor U27753 (N_27753,N_25118,N_24219);
nand U27754 (N_27754,N_24716,N_25736);
and U27755 (N_27755,N_24319,N_25939);
xor U27756 (N_27756,N_24579,N_24279);
and U27757 (N_27757,N_24101,N_25520);
xor U27758 (N_27758,N_24934,N_24383);
or U27759 (N_27759,N_24161,N_24270);
and U27760 (N_27760,N_26039,N_26678);
or U27761 (N_27761,N_24835,N_26177);
or U27762 (N_27762,N_24993,N_25345);
xnor U27763 (N_27763,N_25340,N_24242);
and U27764 (N_27764,N_24866,N_26103);
nand U27765 (N_27765,N_26386,N_26247);
xnor U27766 (N_27766,N_24333,N_25835);
xor U27767 (N_27767,N_26722,N_26753);
or U27768 (N_27768,N_24050,N_26877);
xnor U27769 (N_27769,N_26068,N_26009);
nor U27770 (N_27770,N_24537,N_25652);
nand U27771 (N_27771,N_26927,N_24764);
nor U27772 (N_27772,N_26323,N_25288);
and U27773 (N_27773,N_24998,N_25054);
nand U27774 (N_27774,N_26630,N_25714);
xnor U27775 (N_27775,N_24881,N_24146);
nor U27776 (N_27776,N_25284,N_24593);
or U27777 (N_27777,N_25701,N_26548);
nor U27778 (N_27778,N_26684,N_25172);
nor U27779 (N_27779,N_26692,N_24718);
nor U27780 (N_27780,N_24286,N_25132);
nor U27781 (N_27781,N_26544,N_24046);
xor U27782 (N_27782,N_24859,N_24144);
nand U27783 (N_27783,N_25929,N_26742);
and U27784 (N_27784,N_26321,N_24220);
or U27785 (N_27785,N_24266,N_26872);
nand U27786 (N_27786,N_24413,N_24206);
nor U27787 (N_27787,N_26688,N_26969);
and U27788 (N_27788,N_24588,N_24724);
nor U27789 (N_27789,N_25873,N_25073);
nand U27790 (N_27790,N_24568,N_24923);
or U27791 (N_27791,N_25687,N_25582);
nand U27792 (N_27792,N_26843,N_25230);
and U27793 (N_27793,N_24155,N_26892);
xnor U27794 (N_27794,N_25380,N_24444);
or U27795 (N_27795,N_26826,N_25176);
nor U27796 (N_27796,N_25997,N_25183);
nor U27797 (N_27797,N_26360,N_26265);
xor U27798 (N_27798,N_26322,N_25605);
nand U27799 (N_27799,N_26790,N_24063);
nand U27800 (N_27800,N_25845,N_25447);
nand U27801 (N_27801,N_25528,N_24697);
nand U27802 (N_27802,N_26307,N_24124);
or U27803 (N_27803,N_24791,N_25155);
xnor U27804 (N_27804,N_25570,N_24458);
nand U27805 (N_27805,N_26300,N_26282);
xnor U27806 (N_27806,N_25372,N_24044);
nor U27807 (N_27807,N_24465,N_26889);
or U27808 (N_27808,N_26991,N_24500);
or U27809 (N_27809,N_26587,N_26792);
xor U27810 (N_27810,N_25320,N_25475);
nand U27811 (N_27811,N_25196,N_24442);
xor U27812 (N_27812,N_24297,N_24653);
and U27813 (N_27813,N_25221,N_25327);
nand U27814 (N_27814,N_25926,N_25102);
and U27815 (N_27815,N_25847,N_24814);
and U27816 (N_27816,N_26083,N_26659);
nand U27817 (N_27817,N_24360,N_25494);
nand U27818 (N_27818,N_24895,N_24393);
xor U27819 (N_27819,N_25078,N_25649);
nand U27820 (N_27820,N_26623,N_25133);
or U27821 (N_27821,N_26108,N_24625);
nor U27822 (N_27822,N_24819,N_24730);
nand U27823 (N_27823,N_26263,N_26921);
nor U27824 (N_27824,N_25057,N_26734);
nand U27825 (N_27825,N_24480,N_26089);
nand U27826 (N_27826,N_24798,N_25683);
xor U27827 (N_27827,N_24636,N_26559);
nor U27828 (N_27828,N_26285,N_24267);
xor U27829 (N_27829,N_26582,N_26910);
and U27830 (N_27830,N_24799,N_26345);
and U27831 (N_27831,N_26891,N_24323);
nor U27832 (N_27832,N_24740,N_26308);
nor U27833 (N_27833,N_26696,N_24277);
xnor U27834 (N_27834,N_25458,N_26065);
and U27835 (N_27835,N_24051,N_25776);
and U27836 (N_27836,N_25466,N_26481);
or U27837 (N_27837,N_26098,N_24296);
or U27838 (N_27838,N_25307,N_25675);
and U27839 (N_27839,N_25060,N_24349);
nor U27840 (N_27840,N_25122,N_24816);
or U27841 (N_27841,N_26137,N_24438);
and U27842 (N_27842,N_26059,N_24469);
and U27843 (N_27843,N_26657,N_24769);
or U27844 (N_27844,N_26356,N_25406);
xnor U27845 (N_27845,N_25236,N_26397);
nor U27846 (N_27846,N_24643,N_24861);
nor U27847 (N_27847,N_24854,N_24801);
and U27848 (N_27848,N_24935,N_24989);
and U27849 (N_27849,N_26972,N_26784);
or U27850 (N_27850,N_24054,N_25760);
nor U27851 (N_27851,N_26467,N_24194);
nand U27852 (N_27852,N_24675,N_26720);
nand U27853 (N_27853,N_25075,N_26608);
nand U27854 (N_27854,N_26730,N_25194);
nor U27855 (N_27855,N_24511,N_26650);
or U27856 (N_27856,N_26327,N_24772);
nand U27857 (N_27857,N_25749,N_25411);
nand U27858 (N_27858,N_25689,N_26907);
and U27859 (N_27859,N_25797,N_24411);
or U27860 (N_27860,N_25114,N_24232);
nand U27861 (N_27861,N_26668,N_25896);
nor U27862 (N_27862,N_24326,N_26856);
and U27863 (N_27863,N_25350,N_26781);
nand U27864 (N_27864,N_26417,N_24224);
or U27865 (N_27865,N_25521,N_24872);
and U27866 (N_27866,N_26420,N_26749);
or U27867 (N_27867,N_26171,N_25627);
or U27868 (N_27868,N_24090,N_25592);
or U27869 (N_27869,N_25527,N_25360);
xnor U27870 (N_27870,N_24762,N_24412);
xnor U27871 (N_27871,N_26184,N_24183);
or U27872 (N_27872,N_25238,N_24611);
nand U27873 (N_27873,N_26037,N_25425);
nand U27874 (N_27874,N_25880,N_24208);
nand U27875 (N_27875,N_24431,N_26824);
nor U27876 (N_27876,N_24523,N_26424);
nor U27877 (N_27877,N_25207,N_26862);
nand U27878 (N_27878,N_25969,N_25266);
and U27879 (N_27879,N_25960,N_25459);
nor U27880 (N_27880,N_24534,N_25704);
xor U27881 (N_27881,N_26159,N_25255);
or U27882 (N_27882,N_24780,N_26272);
nand U27883 (N_27883,N_25304,N_26965);
nand U27884 (N_27884,N_24932,N_26621);
xnor U27885 (N_27885,N_26915,N_25676);
nand U27886 (N_27886,N_25398,N_24666);
and U27887 (N_27887,N_26223,N_24900);
or U27888 (N_27888,N_25252,N_25981);
or U27889 (N_27889,N_26444,N_24944);
or U27890 (N_27890,N_26146,N_26102);
xor U27891 (N_27891,N_25587,N_25113);
nand U27892 (N_27892,N_26233,N_26794);
or U27893 (N_27893,N_25297,N_24008);
or U27894 (N_27894,N_25215,N_25718);
xor U27895 (N_27895,N_26396,N_25510);
xnor U27896 (N_27896,N_26613,N_24427);
nand U27897 (N_27897,N_25984,N_24577);
or U27898 (N_27898,N_24023,N_24113);
nor U27899 (N_27899,N_25129,N_24626);
nand U27900 (N_27900,N_24986,N_25832);
nor U27901 (N_27901,N_24904,N_25316);
nor U27902 (N_27902,N_24162,N_24397);
xnor U27903 (N_27903,N_26324,N_26859);
nor U27904 (N_27904,N_25967,N_24337);
xnor U27905 (N_27905,N_25216,N_25744);
nand U27906 (N_27906,N_25748,N_26643);
nor U27907 (N_27907,N_24731,N_26335);
nand U27908 (N_27908,N_26002,N_24357);
and U27909 (N_27909,N_24659,N_26094);
nand U27910 (N_27910,N_24761,N_24396);
and U27911 (N_27911,N_25560,N_24373);
nor U27912 (N_27912,N_24426,N_24953);
or U27913 (N_27913,N_25576,N_24622);
nand U27914 (N_27914,N_24919,N_24273);
or U27915 (N_27915,N_25188,N_26446);
and U27916 (N_27916,N_26873,N_26204);
and U27917 (N_27917,N_26605,N_26885);
and U27918 (N_27918,N_25149,N_26957);
xor U27919 (N_27919,N_26456,N_25336);
nand U27920 (N_27920,N_24860,N_24123);
nand U27921 (N_27921,N_25436,N_24733);
nand U27922 (N_27922,N_24827,N_24390);
and U27923 (N_27923,N_25069,N_24010);
and U27924 (N_27924,N_26346,N_24137);
nor U27925 (N_27925,N_26580,N_26038);
or U27926 (N_27926,N_26505,N_24968);
nor U27927 (N_27927,N_25293,N_24301);
and U27928 (N_27928,N_24464,N_25878);
nor U27929 (N_27929,N_24211,N_24911);
nor U27930 (N_27930,N_25192,N_25257);
and U27931 (N_27931,N_26899,N_26904);
or U27932 (N_27932,N_25591,N_24831);
xnor U27933 (N_27933,N_26325,N_25844);
and U27934 (N_27934,N_25099,N_24015);
and U27935 (N_27935,N_24216,N_24282);
and U27936 (N_27936,N_25586,N_24873);
nand U27937 (N_27937,N_25596,N_25315);
nand U27938 (N_27938,N_26006,N_25220);
or U27939 (N_27939,N_25992,N_25755);
and U27940 (N_27940,N_25912,N_26558);
and U27941 (N_27941,N_25142,N_25223);
xnor U27942 (N_27942,N_26348,N_24530);
nor U27943 (N_27943,N_24818,N_26315);
or U27944 (N_27944,N_26500,N_25784);
nand U27945 (N_27945,N_26363,N_25700);
nor U27946 (N_27946,N_25170,N_24862);
and U27947 (N_27947,N_24686,N_26293);
and U27948 (N_27948,N_24725,N_25515);
nand U27949 (N_27949,N_26070,N_25761);
or U27950 (N_27950,N_24234,N_25814);
nor U27951 (N_27951,N_25514,N_25986);
or U27952 (N_27952,N_24295,N_26144);
xnor U27953 (N_27953,N_24119,N_26771);
or U27954 (N_27954,N_24204,N_24378);
nor U27955 (N_27955,N_25235,N_26200);
xor U27956 (N_27956,N_25739,N_24120);
and U27957 (N_27957,N_25096,N_25637);
or U27958 (N_27958,N_24563,N_26672);
xnor U27959 (N_27959,N_26163,N_25519);
nor U27960 (N_27960,N_26194,N_26409);
nand U27961 (N_27961,N_26043,N_26342);
or U27962 (N_27962,N_24071,N_24805);
nand U27963 (N_27963,N_26150,N_25012);
xor U27964 (N_27964,N_25858,N_24154);
xnor U27965 (N_27965,N_26685,N_25608);
nand U27966 (N_27966,N_25296,N_24954);
or U27967 (N_27967,N_24926,N_24797);
nor U27968 (N_27968,N_26066,N_25569);
and U27969 (N_27969,N_25545,N_24812);
and U27970 (N_27970,N_24077,N_24343);
or U27971 (N_27971,N_25972,N_24353);
and U27972 (N_27972,N_26776,N_25501);
nand U27973 (N_27973,N_26203,N_24109);
or U27974 (N_27974,N_26419,N_24450);
and U27975 (N_27975,N_24956,N_26241);
and U27976 (N_27976,N_25379,N_24694);
or U27977 (N_27977,N_24317,N_24268);
or U27978 (N_27978,N_26413,N_24097);
xnor U27979 (N_27979,N_24907,N_24788);
nor U27980 (N_27980,N_24285,N_25076);
nand U27981 (N_27981,N_25427,N_26472);
xnor U27982 (N_27982,N_24372,N_24169);
nor U27983 (N_27983,N_24552,N_25232);
or U27984 (N_27984,N_24547,N_25504);
xor U27985 (N_27985,N_25332,N_25473);
xnor U27986 (N_27986,N_26021,N_26511);
xnor U27987 (N_27987,N_26717,N_26099);
or U27988 (N_27988,N_24782,N_24111);
nor U27989 (N_27989,N_25735,N_25862);
and U27990 (N_27990,N_25498,N_26535);
nor U27991 (N_27991,N_25922,N_26357);
or U27992 (N_27992,N_24823,N_25486);
and U27993 (N_27993,N_24166,N_26362);
xnor U27994 (N_27994,N_24185,N_25000);
nand U27995 (N_27995,N_24999,N_25161);
or U27996 (N_27996,N_26366,N_25795);
xnor U27997 (N_27997,N_24619,N_25937);
nand U27998 (N_27998,N_26051,N_26588);
nand U27999 (N_27999,N_25721,N_25148);
nor U28000 (N_28000,N_25558,N_25840);
and U28001 (N_28001,N_26618,N_24249);
or U28002 (N_28002,N_24581,N_25935);
nor U28003 (N_28003,N_25145,N_26164);
nand U28004 (N_28004,N_25428,N_25663);
or U28005 (N_28005,N_24820,N_25439);
nor U28006 (N_28006,N_24995,N_25921);
nand U28007 (N_28007,N_25376,N_26516);
xor U28008 (N_28008,N_25409,N_25820);
nand U28009 (N_28009,N_26976,N_26189);
or U28010 (N_28010,N_26286,N_25007);
nand U28011 (N_28011,N_26072,N_26215);
or U28012 (N_28012,N_24891,N_25135);
nand U28013 (N_28013,N_26740,N_24331);
or U28014 (N_28014,N_24521,N_26682);
nand U28015 (N_28015,N_24443,N_26004);
or U28016 (N_28016,N_25720,N_26010);
nand U28017 (N_28017,N_26980,N_26598);
or U28018 (N_28018,N_26546,N_24539);
and U28019 (N_28019,N_24674,N_26798);
or U28020 (N_28020,N_26926,N_24105);
or U28021 (N_28021,N_24497,N_25866);
nor U28022 (N_28022,N_26746,N_25877);
nand U28023 (N_28023,N_26309,N_25696);
xor U28024 (N_28024,N_26222,N_25283);
and U28025 (N_28025,N_25567,N_24196);
xor U28026 (N_28026,N_24602,N_26658);
nand U28027 (N_28027,N_24310,N_25904);
xor U28028 (N_28028,N_24151,N_25647);
and U28029 (N_28029,N_24002,N_26469);
nand U28030 (N_28030,N_26273,N_24952);
nor U28031 (N_28031,N_26756,N_24804);
or U28032 (N_28032,N_25111,N_24031);
xor U28033 (N_28033,N_26393,N_26142);
xor U28034 (N_28034,N_24676,N_24680);
and U28035 (N_28035,N_24049,N_24184);
nor U28036 (N_28036,N_24032,N_26478);
and U28037 (N_28037,N_26112,N_24737);
or U28038 (N_28038,N_26810,N_26817);
or U28039 (N_28039,N_24106,N_25931);
and U28040 (N_28040,N_24836,N_25174);
nand U28041 (N_28041,N_25624,N_26491);
nand U28042 (N_28042,N_25534,N_25092);
nand U28043 (N_28043,N_24575,N_25581);
nor U28044 (N_28044,N_24897,N_24375);
xor U28045 (N_28045,N_26962,N_24180);
nand U28046 (N_28046,N_25572,N_26187);
nand U28047 (N_28047,N_26214,N_24246);
nor U28048 (N_28048,N_24290,N_24125);
nand U28049 (N_28049,N_25291,N_24112);
and U28050 (N_28050,N_26528,N_26176);
and U28051 (N_28051,N_26555,N_24179);
nand U28052 (N_28052,N_26231,N_26788);
nor U28053 (N_28053,N_25237,N_25203);
nand U28054 (N_28054,N_26106,N_24660);
and U28055 (N_28055,N_26936,N_24600);
or U28056 (N_28056,N_25990,N_26331);
xnor U28057 (N_28057,N_25490,N_25051);
nor U28058 (N_28058,N_25402,N_25050);
and U28059 (N_28059,N_25178,N_24128);
nor U28060 (N_28060,N_25685,N_25168);
xor U28061 (N_28061,N_24803,N_24754);
nand U28062 (N_28062,N_26473,N_26499);
and U28063 (N_28063,N_25301,N_24948);
xor U28064 (N_28064,N_25544,N_25120);
and U28065 (N_28065,N_26259,N_24612);
nor U28066 (N_28066,N_24190,N_25943);
and U28067 (N_28067,N_24841,N_24318);
nor U28068 (N_28068,N_25933,N_24158);
nor U28069 (N_28069,N_26845,N_24542);
nor U28070 (N_28070,N_24781,N_26996);
and U28071 (N_28071,N_26882,N_25090);
and U28072 (N_28072,N_25517,N_26627);
nor U28073 (N_28073,N_25105,N_26461);
nor U28074 (N_28074,N_24759,N_25421);
nor U28075 (N_28075,N_26540,N_25970);
or U28076 (N_28076,N_24320,N_25836);
and U28077 (N_28077,N_25222,N_25080);
nand U28078 (N_28078,N_26238,N_25024);
and U28079 (N_28079,N_26652,N_26728);
and U28080 (N_28080,N_25611,N_24598);
nor U28081 (N_28081,N_26577,N_26465);
or U28082 (N_28082,N_24758,N_24638);
nor U28083 (N_28083,N_24147,N_26797);
nor U28084 (N_28084,N_25317,N_26508);
xor U28085 (N_28085,N_26994,N_24722);
and U28086 (N_28086,N_26492,N_25884);
and U28087 (N_28087,N_25483,N_26169);
nand U28088 (N_28088,N_26710,N_26463);
and U28089 (N_28089,N_25747,N_24969);
nand U28090 (N_28090,N_26120,N_26379);
or U28091 (N_28091,N_25557,N_25190);
xnor U28092 (N_28092,N_24322,N_24029);
xor U28093 (N_28093,N_25688,N_26278);
and U28094 (N_28094,N_26584,N_26125);
nand U28095 (N_28095,N_25634,N_25961);
and U28096 (N_28096,N_25973,N_26747);
xnor U28097 (N_28097,N_24406,N_25920);
xnor U28098 (N_28098,N_24947,N_24454);
xnor U28099 (N_28099,N_24945,N_25620);
and U28100 (N_28100,N_24560,N_25625);
or U28101 (N_28101,N_26298,N_25319);
nand U28102 (N_28102,N_25016,N_24938);
or U28103 (N_28103,N_24876,N_26340);
nor U28104 (N_28104,N_25885,N_25934);
nor U28105 (N_28105,N_25434,N_24851);
xor U28106 (N_28106,N_24058,N_25305);
nor U28107 (N_28107,N_24828,N_24869);
or U28108 (N_28108,N_24709,N_24941);
and U28109 (N_28109,N_24351,N_24441);
and U28110 (N_28110,N_25803,N_24668);
and U28111 (N_28111,N_24278,N_26594);
nor U28112 (N_28112,N_26172,N_25628);
and U28113 (N_28113,N_25726,N_26211);
xnor U28114 (N_28114,N_25053,N_26261);
nand U28115 (N_28115,N_26990,N_24172);
nor U28116 (N_28116,N_26436,N_24259);
nor U28117 (N_28117,N_25338,N_24288);
nand U28118 (N_28118,N_25941,N_26855);
or U28119 (N_28119,N_25424,N_26670);
xnor U28120 (N_28120,N_25910,N_26121);
nand U28121 (N_28121,N_26040,N_25456);
nand U28122 (N_28122,N_26985,N_26312);
and U28123 (N_28123,N_26707,N_24635);
or U28124 (N_28124,N_25084,N_24601);
nand U28125 (N_28125,N_25601,N_24813);
nor U28126 (N_28126,N_25160,N_24770);
nand U28127 (N_28127,N_26796,N_26533);
nor U28128 (N_28128,N_24931,N_24466);
or U28129 (N_28129,N_26412,N_25432);
nand U28130 (N_28130,N_26268,N_24591);
nand U28131 (N_28131,N_24908,N_24596);
nand U28132 (N_28132,N_26939,N_26759);
nand U28133 (N_28133,N_26656,N_26851);
nor U28134 (N_28134,N_24894,N_26947);
and U28135 (N_28135,N_25796,N_26117);
and U28136 (N_28136,N_24041,N_26640);
or U28137 (N_28137,N_25426,N_26028);
nor U28138 (N_28138,N_25064,N_25435);
xor U28139 (N_28139,N_26767,N_24637);
and U28140 (N_28140,N_26236,N_26619);
xor U28141 (N_28141,N_26459,N_25181);
nand U28142 (N_28142,N_26774,N_26634);
nand U28143 (N_28143,N_26909,N_26770);
xor U28144 (N_28144,N_24303,N_25945);
nand U28145 (N_28145,N_26069,N_24771);
and U28146 (N_28146,N_26351,N_25769);
and U28147 (N_28147,N_25445,N_26943);
or U28148 (N_28148,N_24200,N_25309);
or U28149 (N_28149,N_26574,N_25801);
and U28150 (N_28150,N_26526,N_24898);
nor U28151 (N_28151,N_26773,N_24729);
nor U28152 (N_28152,N_25957,N_26950);
and U28153 (N_28153,N_25918,N_25825);
nand U28154 (N_28154,N_25575,N_25809);
or U28155 (N_28155,N_24014,N_25954);
nor U28156 (N_28156,N_26326,N_24191);
or U28157 (N_28157,N_24210,N_26974);
xnor U28158 (N_28158,N_24940,N_24004);
nor U28159 (N_28159,N_25300,N_26635);
or U28160 (N_28160,N_25318,N_26097);
nor U28161 (N_28161,N_26139,N_25865);
nand U28162 (N_28162,N_24462,N_26933);
or U28163 (N_28163,N_24750,N_25577);
or U28164 (N_28164,N_25294,N_24877);
nor U28165 (N_28165,N_26912,N_25679);
nor U28166 (N_28166,N_24005,N_26842);
and U28167 (N_28167,N_26847,N_25629);
nand U28168 (N_28168,N_26181,N_24370);
or U28169 (N_28169,N_25999,N_24018);
and U28170 (N_28170,N_24496,N_26922);
nor U28171 (N_28171,N_26563,N_26989);
xor U28172 (N_28172,N_24118,N_26561);
or U28173 (N_28173,N_25020,N_26000);
xor U28174 (N_28174,N_25437,N_24467);
or U28175 (N_28175,N_26210,N_24742);
nand U28176 (N_28176,N_25460,N_25373);
nor U28177 (N_28177,N_25063,N_25130);
or U28178 (N_28178,N_24341,N_24424);
nand U28179 (N_28179,N_26586,N_25833);
or U28180 (N_28180,N_26115,N_24455);
xor U28181 (N_28181,N_25202,N_24291);
xor U28182 (N_28182,N_26971,N_24587);
or U28183 (N_28183,N_25998,N_24839);
nand U28184 (N_28184,N_26022,N_26237);
xor U28185 (N_28185,N_24597,N_24017);
xnor U28186 (N_28186,N_25853,N_25042);
and U28187 (N_28187,N_26170,N_26084);
or U28188 (N_28188,N_25339,N_26857);
and U28189 (N_28189,N_25103,N_24967);
nor U28190 (N_28190,N_26292,N_25725);
xnor U28191 (N_28191,N_25267,N_26631);
nor U28192 (N_28192,N_25964,N_26130);
nand U28193 (N_28193,N_24641,N_25599);
xnor U28194 (N_28194,N_24489,N_26959);
xnor U28195 (N_28195,N_24446,N_24837);
or U28196 (N_28196,N_25403,N_26924);
nor U28197 (N_28197,N_24007,N_25826);
nor U28198 (N_28198,N_26400,N_26932);
or U28199 (N_28199,N_25980,N_26821);
xnor U28200 (N_28200,N_26905,N_24274);
and U28201 (N_28201,N_26141,N_25600);
or U28202 (N_28202,N_26918,N_25603);
and U28203 (N_28203,N_24350,N_25852);
nor U28204 (N_28204,N_24880,N_24992);
xor U28205 (N_28205,N_25058,N_25484);
xor U28206 (N_28206,N_24517,N_24562);
and U28207 (N_28207,N_25794,N_26143);
nor U28208 (N_28208,N_26421,N_25993);
and U28209 (N_28209,N_26361,N_25762);
or U28210 (N_28210,N_25195,N_26628);
nor U28211 (N_28211,N_26280,N_26458);
nor U28212 (N_28212,N_26404,N_25282);
xnor U28213 (N_28213,N_25781,N_25477);
xor U28214 (N_28214,N_24867,N_24055);
or U28215 (N_28215,N_25052,N_24913);
nor U28216 (N_28216,N_26698,N_26061);
or U28217 (N_28217,N_26304,N_24936);
nand U28218 (N_28218,N_25481,N_26701);
and U28219 (N_28219,N_26202,N_25330);
and U28220 (N_28220,N_24774,N_25248);
nand U28221 (N_28221,N_26291,N_26828);
or U28222 (N_28222,N_26840,N_25919);
nor U28223 (N_28223,N_24959,N_26147);
xnor U28224 (N_28224,N_24045,N_26161);
or U28225 (N_28225,N_26328,N_24139);
and U28226 (N_28226,N_24929,N_25664);
and U28227 (N_28227,N_25817,N_24024);
nor U28228 (N_28228,N_26570,N_25179);
nor U28229 (N_28229,N_25348,N_25552);
xor U28230 (N_28230,N_25018,N_25741);
nand U28231 (N_28231,N_26449,N_25204);
nor U28232 (N_28232,N_25958,N_26179);
xor U28233 (N_28233,N_25743,N_26813);
and U28234 (N_28234,N_26591,N_25786);
and U28235 (N_28235,N_24272,N_26704);
or U28236 (N_28236,N_24633,N_25532);
or U28237 (N_28237,N_26157,N_25965);
nor U28238 (N_28238,N_25745,N_26946);
nor U28239 (N_28239,N_24143,N_25831);
and U28240 (N_28240,N_24252,N_25392);
nor U28241 (N_28241,N_26408,N_26155);
nor U28242 (N_28242,N_25962,N_25513);
and U28243 (N_28243,N_24067,N_24418);
or U28244 (N_28244,N_25323,N_26190);
or U28245 (N_28245,N_25156,N_26080);
xor U28246 (N_28246,N_25656,N_24691);
xor U28247 (N_28247,N_25143,N_25895);
and U28248 (N_28248,N_25279,N_26755);
nand U28249 (N_28249,N_25422,N_25371);
xnor U28250 (N_28250,N_25049,N_25516);
xnor U28251 (N_28251,N_24655,N_24254);
nor U28252 (N_28252,N_24863,N_25423);
nand U28253 (N_28253,N_24707,N_26866);
xor U28254 (N_28254,N_26600,N_24069);
or U28255 (N_28255,N_24235,N_26336);
nand U28256 (N_28256,N_26647,N_25107);
nor U28257 (N_28257,N_25191,N_26012);
nor U28258 (N_28258,N_24025,N_26809);
or U28259 (N_28259,N_25709,N_24240);
xnor U28260 (N_28260,N_24658,N_26216);
or U28261 (N_28261,N_24607,N_25901);
or U28262 (N_28262,N_24887,N_24313);
xor U28263 (N_28263,N_24013,N_24459);
nor U28264 (N_28264,N_25541,N_24487);
xnor U28265 (N_28265,N_25774,N_25869);
and U28266 (N_28266,N_24793,N_25821);
nand U28267 (N_28267,N_25326,N_26629);
and U28268 (N_28268,N_25537,N_26982);
nand U28269 (N_28269,N_26961,N_24980);
xor U28270 (N_28270,N_24558,N_26124);
nand U28271 (N_28271,N_25506,N_24702);
or U28272 (N_28272,N_26539,N_25002);
or U28273 (N_28273,N_25302,N_25401);
or U28274 (N_28274,N_24327,N_25182);
nand U28275 (N_28275,N_26956,N_25126);
nand U28276 (N_28276,N_26050,N_25547);
nor U28277 (N_28277,N_24580,N_24609);
and U28278 (N_28278,N_25654,N_26483);
and U28279 (N_28279,N_24092,N_26531);
and U28280 (N_28280,N_26923,N_26358);
xnor U28281 (N_28281,N_26938,N_24214);
or U28282 (N_28282,N_24614,N_25407);
nand U28283 (N_28283,N_26107,N_26209);
nand U28284 (N_28284,N_26888,N_25903);
or U28285 (N_28285,N_25303,N_26243);
nand U28286 (N_28286,N_24110,N_25916);
or U28287 (N_28287,N_25061,N_24167);
and U28288 (N_28288,N_26497,N_24369);
nor U28289 (N_28289,N_24795,N_25518);
or U28290 (N_28290,N_24642,N_24284);
and U28291 (N_28291,N_25471,N_24874);
or U28292 (N_28292,N_24950,N_24893);
nand U28293 (N_28293,N_25508,N_24164);
xnor U28294 (N_28294,N_26633,N_26445);
or U28295 (N_28295,N_25289,N_25607);
nand U28296 (N_28296,N_26082,N_24505);
or U28297 (N_28297,N_25463,N_25665);
xor U28298 (N_28298,N_26979,N_25077);
and U28299 (N_28299,N_26645,N_26854);
nand U28300 (N_28300,N_24634,N_25246);
and U28301 (N_28301,N_26565,N_26305);
or U28302 (N_28302,N_24703,N_24565);
nand U28303 (N_28303,N_26480,N_24909);
or U28304 (N_28304,N_25716,N_24094);
nand U28305 (N_28305,N_25153,N_24623);
and U28306 (N_28306,N_24140,N_26566);
xnor U28307 (N_28307,N_26352,N_24704);
and U28308 (N_28308,N_25031,N_25746);
and U28309 (N_28309,N_24906,N_26931);
nor U28310 (N_28310,N_24460,N_24159);
or U28311 (N_28311,N_24415,N_26451);
nand U28312 (N_28312,N_24661,N_26579);
or U28313 (N_28313,N_25404,N_25356);
xor U28314 (N_28314,N_26525,N_25355);
or U28315 (N_28315,N_26655,N_24652);
nand U28316 (N_28316,N_24009,N_26435);
xnor U28317 (N_28317,N_24514,N_26438);
nand U28318 (N_28318,N_24672,N_24964);
or U28319 (N_28319,N_24549,N_25590);
xor U28320 (N_28320,N_25314,N_25464);
nor U28321 (N_28321,N_24237,N_24470);
nor U28322 (N_28322,N_26495,N_24026);
nand U28323 (N_28323,N_25479,N_24053);
nor U28324 (N_28324,N_26086,N_25270);
nor U28325 (N_28325,N_25616,N_24401);
and U28326 (N_28326,N_25658,N_25838);
nor U28327 (N_28327,N_24604,N_24451);
nand U28328 (N_28328,N_24020,N_25095);
xor U28329 (N_28329,N_24250,N_25946);
xnor U28330 (N_28330,N_25691,N_25085);
nor U28331 (N_28331,N_25015,N_26160);
or U28332 (N_28332,N_26543,N_24141);
and U28333 (N_28333,N_24687,N_26725);
nand U28334 (N_28334,N_24086,N_26765);
or U28335 (N_28335,N_26908,N_25029);
nor U28336 (N_28336,N_26078,N_26547);
xor U28337 (N_28337,N_24621,N_24062);
xor U28338 (N_28338,N_24225,N_25476);
and U28339 (N_28339,N_26964,N_26779);
xor U28340 (N_28340,N_26601,N_24728);
xor U28341 (N_28341,N_25614,N_24984);
and U28342 (N_28342,N_24011,N_26754);
nand U28343 (N_28343,N_25897,N_26376);
xor U28344 (N_28344,N_25551,N_26085);
xnor U28345 (N_28345,N_24117,N_25311);
nand U28346 (N_28346,N_24064,N_24566);
nand U28347 (N_28347,N_25093,N_24888);
or U28348 (N_28348,N_24417,N_26848);
or U28349 (N_28349,N_26488,N_24937);
and U28350 (N_28350,N_24613,N_24857);
nand U28351 (N_28351,N_26595,N_25366);
nor U28352 (N_28352,N_25036,N_25417);
and U28353 (N_28353,N_24463,N_26079);
nand U28354 (N_28354,N_26230,N_24108);
xor U28355 (N_28355,N_24578,N_26675);
and U28356 (N_28356,N_26403,N_26930);
and U28357 (N_28357,N_25021,N_24669);
or U28358 (N_28358,N_24275,N_25568);
xnor U28359 (N_28359,N_25381,N_25127);
nor U28360 (N_28360,N_24380,N_24309);
nand U28361 (N_28361,N_26666,N_26988);
xor U28362 (N_28362,N_26612,N_25094);
xor U28363 (N_28363,N_25511,N_25610);
and U28364 (N_28364,N_25751,N_25673);
and U28365 (N_28365,N_25546,N_24917);
and U28366 (N_28366,N_24656,N_25548);
nor U28367 (N_28367,N_26735,N_24205);
nor U28368 (N_28368,N_24540,N_24910);
xor U28369 (N_28369,N_26867,N_24456);
nand U28370 (N_28370,N_26530,N_25233);
or U28371 (N_28371,N_26513,N_26799);
or U28372 (N_28372,N_24384,N_24715);
xor U28373 (N_28373,N_25850,N_24627);
and U28374 (N_28374,N_24410,N_26126);
or U28375 (N_28375,N_26208,N_26193);
nand U28376 (N_28376,N_24223,N_25104);
and U28377 (N_28377,N_26314,N_26248);
and U28378 (N_28378,N_24479,N_25622);
and U28379 (N_28379,N_26398,N_26791);
nand U28380 (N_28380,N_24481,N_24136);
nand U28381 (N_28381,N_24150,N_26221);
or U28382 (N_28382,N_26299,N_24548);
nand U28383 (N_28383,N_24060,N_24258);
and U28384 (N_28384,N_24997,N_24994);
or U28385 (N_28385,N_24494,N_24080);
or U28386 (N_28386,N_24160,N_26803);
xnor U28387 (N_28387,N_24662,N_24752);
nand U28388 (N_28388,N_26154,N_25790);
xor U28389 (N_28389,N_26993,N_25928);
xnor U28390 (N_28390,N_25217,N_25719);
nor U28391 (N_28391,N_25843,N_24556);
and U28392 (N_28392,N_25561,N_26727);
nor U28393 (N_28393,N_25496,N_25612);
xor U28394 (N_28394,N_24306,N_25124);
xnor U28395 (N_28395,N_25732,N_26733);
xnor U28396 (N_28396,N_26719,N_25956);
and U28397 (N_28397,N_24755,N_26132);
nor U28398 (N_28398,N_25470,N_24334);
nand U28399 (N_28399,N_25584,N_26829);
nor U28400 (N_28400,N_24584,N_25218);
and U28401 (N_28401,N_26224,N_24564);
nand U28402 (N_28402,N_24654,N_26425);
nor U28403 (N_28403,N_25907,N_26270);
nand U28404 (N_28404,N_25682,N_26123);
nand U28405 (N_28405,N_26823,N_24366);
and U28406 (N_28406,N_24006,N_25911);
and U28407 (N_28407,N_26339,N_24875);
nor U28408 (N_28408,N_26567,N_25529);
nor U28409 (N_28409,N_26805,N_25265);
nand U28410 (N_28410,N_25893,N_25692);
and U28411 (N_28411,N_24673,N_25640);
nand U28412 (N_28412,N_25384,N_24617);
nor U28413 (N_28413,N_26023,N_26703);
xor U28414 (N_28414,N_24747,N_26694);
or U28415 (N_28415,N_26032,N_26462);
and U28416 (N_28416,N_24928,N_26119);
nor U28417 (N_28417,N_24620,N_26697);
and U28418 (N_28418,N_24573,N_26737);
nand U28419 (N_28419,N_25643,N_26367);
xor U28420 (N_28420,N_25936,N_24506);
nor U28421 (N_28421,N_25032,N_25500);
nor U28422 (N_28422,N_26617,N_24188);
xor U28423 (N_28423,N_25580,N_24217);
and U28424 (N_28424,N_25333,N_26416);
xor U28425 (N_28425,N_24785,N_25389);
nor U28426 (N_28426,N_24021,N_26816);
or U28427 (N_28427,N_24165,N_25027);
xor U28428 (N_28428,N_25412,N_25286);
nand U28429 (N_28429,N_25039,N_26294);
xnor U28430 (N_28430,N_25657,N_26062);
nand U28431 (N_28431,N_25388,N_24991);
xnor U28432 (N_28432,N_25141,N_24037);
nor U28433 (N_28433,N_25083,N_26519);
or U28434 (N_28434,N_26045,N_26536);
nand U28435 (N_28435,N_26486,N_24491);
or U28436 (N_28436,N_24076,N_26127);
or U28437 (N_28437,N_25109,N_24461);
or U28438 (N_28438,N_24035,N_26590);
or U28439 (N_28439,N_26646,N_26785);
and U28440 (N_28440,N_25699,N_24389);
or U28441 (N_28441,N_24889,N_26778);
nand U28442 (N_28442,N_25322,N_25522);
nor U28443 (N_28443,N_24001,N_26390);
nor U28444 (N_28444,N_24000,N_25210);
nor U28445 (N_28445,N_25902,N_26058);
and U28446 (N_28446,N_24685,N_26715);
nand U28447 (N_28447,N_24066,N_25365);
nand U28448 (N_28448,N_25550,N_24766);
or U28449 (N_28449,N_24746,N_25875);
nand U28450 (N_28450,N_24665,N_25924);
xor U28451 (N_28451,N_25626,N_24574);
nand U28452 (N_28452,N_26475,N_24377);
xnor U28453 (N_28453,N_25894,N_25026);
or U28454 (N_28454,N_24142,N_25249);
nand U28455 (N_28455,N_26841,N_26013);
nand U28456 (N_28456,N_26973,N_24684);
nor U28457 (N_28457,N_25344,N_24726);
xnor U28458 (N_28458,N_25764,N_24842);
xor U28459 (N_28459,N_25968,N_26014);
nor U28460 (N_28460,N_25011,N_26978);
nand U28461 (N_28461,N_26306,N_24516);
nor U28462 (N_28462,N_26651,N_25710);
nand U28463 (N_28463,N_24955,N_25750);
nor U28464 (N_28464,N_25037,N_25733);
nand U28465 (N_28465,N_25146,N_26551);
nor U28466 (N_28466,N_26391,N_25566);
xor U28467 (N_28467,N_26332,N_24222);
nand U28468 (N_28468,N_25681,N_25927);
and U28469 (N_28469,N_24878,N_24361);
and U28470 (N_28470,N_24342,N_25593);
xnor U28471 (N_28471,N_26919,N_26983);
nand U28472 (N_28472,N_24215,N_25947);
and U28473 (N_28473,N_26145,N_26825);
nor U28474 (N_28474,N_25151,N_24541);
or U28475 (N_28475,N_26116,N_24592);
nand U28476 (N_28476,N_25623,N_25329);
or U28477 (N_28477,N_24651,N_26562);
nor U28478 (N_28478,N_26073,N_24753);
and U28479 (N_28479,N_24330,N_24988);
or U28480 (N_28480,N_24695,N_25635);
or U28481 (N_28481,N_26020,N_24605);
and U28482 (N_28482,N_24833,N_24822);
nor U28483 (N_28483,N_24262,N_26870);
xnor U28484 (N_28484,N_24849,N_24981);
nand U28485 (N_28485,N_25137,N_24856);
nor U28486 (N_28486,N_25951,N_25800);
or U28487 (N_28487,N_26834,N_24488);
and U28488 (N_28488,N_25358,N_25134);
or U28489 (N_28489,N_26067,N_25708);
xor U28490 (N_28490,N_26319,N_24646);
xor U28491 (N_28491,N_25280,N_25448);
or U28492 (N_28492,N_26197,N_26199);
nor U28493 (N_28493,N_24544,N_25171);
or U28494 (N_28494,N_25978,N_25415);
nand U28495 (N_28495,N_26387,N_25209);
or U28496 (N_28496,N_24193,N_24777);
nor U28497 (N_28497,N_26178,N_26353);
or U28498 (N_28498,N_25410,N_24720);
or U28499 (N_28499,N_26359,N_26865);
and U28500 (N_28500,N_26164,N_24878);
nand U28501 (N_28501,N_26803,N_26001);
or U28502 (N_28502,N_25605,N_24238);
and U28503 (N_28503,N_25328,N_26348);
nand U28504 (N_28504,N_26199,N_26054);
or U28505 (N_28505,N_26069,N_26378);
nor U28506 (N_28506,N_24086,N_24855);
or U28507 (N_28507,N_24161,N_25002);
nor U28508 (N_28508,N_26024,N_25860);
xnor U28509 (N_28509,N_25284,N_24321);
nand U28510 (N_28510,N_25323,N_26368);
and U28511 (N_28511,N_24204,N_24314);
nand U28512 (N_28512,N_25811,N_25831);
nor U28513 (N_28513,N_25845,N_26324);
xnor U28514 (N_28514,N_26939,N_24744);
nand U28515 (N_28515,N_25359,N_25980);
or U28516 (N_28516,N_25880,N_24110);
nor U28517 (N_28517,N_26305,N_25933);
nand U28518 (N_28518,N_26316,N_24651);
xor U28519 (N_28519,N_26202,N_24265);
nor U28520 (N_28520,N_24479,N_26194);
nor U28521 (N_28521,N_26106,N_26345);
xor U28522 (N_28522,N_24373,N_24413);
xor U28523 (N_28523,N_25029,N_24114);
nor U28524 (N_28524,N_24042,N_24041);
nor U28525 (N_28525,N_24835,N_26361);
and U28526 (N_28526,N_24477,N_26678);
nor U28527 (N_28527,N_24066,N_25723);
nor U28528 (N_28528,N_24930,N_24769);
or U28529 (N_28529,N_26800,N_24875);
nand U28530 (N_28530,N_24798,N_24919);
nand U28531 (N_28531,N_25607,N_25889);
nand U28532 (N_28532,N_26622,N_24335);
nand U28533 (N_28533,N_25363,N_26492);
nor U28534 (N_28534,N_26529,N_26558);
or U28535 (N_28535,N_25951,N_26767);
nor U28536 (N_28536,N_24595,N_24384);
nor U28537 (N_28537,N_26293,N_25748);
nand U28538 (N_28538,N_24104,N_26083);
or U28539 (N_28539,N_26869,N_24890);
or U28540 (N_28540,N_25839,N_24190);
nor U28541 (N_28541,N_25558,N_24252);
nand U28542 (N_28542,N_24292,N_24224);
nor U28543 (N_28543,N_24257,N_26590);
and U28544 (N_28544,N_26706,N_25245);
and U28545 (N_28545,N_25917,N_25337);
xor U28546 (N_28546,N_24451,N_25868);
nor U28547 (N_28547,N_25597,N_24522);
or U28548 (N_28548,N_24278,N_24682);
xnor U28549 (N_28549,N_25804,N_25981);
nand U28550 (N_28550,N_26385,N_26463);
nor U28551 (N_28551,N_25736,N_24570);
or U28552 (N_28552,N_24109,N_26224);
nand U28553 (N_28553,N_25318,N_25044);
nor U28554 (N_28554,N_25592,N_25013);
xnor U28555 (N_28555,N_26342,N_24208);
and U28556 (N_28556,N_25119,N_24489);
and U28557 (N_28557,N_26452,N_25586);
nand U28558 (N_28558,N_25553,N_25927);
and U28559 (N_28559,N_24752,N_25584);
nor U28560 (N_28560,N_24687,N_25947);
nor U28561 (N_28561,N_25018,N_25736);
and U28562 (N_28562,N_26485,N_26322);
nor U28563 (N_28563,N_24116,N_26319);
nor U28564 (N_28564,N_26126,N_26469);
or U28565 (N_28565,N_25899,N_26251);
nand U28566 (N_28566,N_25056,N_24389);
or U28567 (N_28567,N_25013,N_26616);
nor U28568 (N_28568,N_26233,N_26942);
xnor U28569 (N_28569,N_24732,N_24850);
nor U28570 (N_28570,N_26507,N_26533);
xor U28571 (N_28571,N_26713,N_25099);
and U28572 (N_28572,N_25682,N_26984);
and U28573 (N_28573,N_25613,N_25979);
or U28574 (N_28574,N_24781,N_26324);
xor U28575 (N_28575,N_24660,N_26653);
or U28576 (N_28576,N_24073,N_24767);
xnor U28577 (N_28577,N_24870,N_24189);
nor U28578 (N_28578,N_24238,N_25039);
or U28579 (N_28579,N_26625,N_26706);
xor U28580 (N_28580,N_25620,N_26432);
and U28581 (N_28581,N_26590,N_26380);
xnor U28582 (N_28582,N_24607,N_25387);
and U28583 (N_28583,N_25668,N_26308);
and U28584 (N_28584,N_24175,N_26713);
or U28585 (N_28585,N_26418,N_24613);
and U28586 (N_28586,N_25355,N_26129);
nor U28587 (N_28587,N_25510,N_26669);
xor U28588 (N_28588,N_25699,N_24704);
nand U28589 (N_28589,N_26239,N_26960);
nand U28590 (N_28590,N_24716,N_24347);
nor U28591 (N_28591,N_25476,N_24550);
and U28592 (N_28592,N_26382,N_25738);
and U28593 (N_28593,N_24716,N_26753);
xnor U28594 (N_28594,N_26212,N_24347);
or U28595 (N_28595,N_24404,N_24584);
nor U28596 (N_28596,N_25954,N_24198);
or U28597 (N_28597,N_25011,N_24769);
or U28598 (N_28598,N_26106,N_24952);
nor U28599 (N_28599,N_25408,N_26471);
nand U28600 (N_28600,N_25628,N_26535);
and U28601 (N_28601,N_25542,N_26689);
xor U28602 (N_28602,N_24781,N_24670);
and U28603 (N_28603,N_25793,N_25027);
nand U28604 (N_28604,N_25225,N_24784);
and U28605 (N_28605,N_26570,N_25136);
nand U28606 (N_28606,N_25658,N_25466);
and U28607 (N_28607,N_25772,N_24142);
or U28608 (N_28608,N_26635,N_24799);
or U28609 (N_28609,N_25701,N_25371);
nand U28610 (N_28610,N_26609,N_25215);
and U28611 (N_28611,N_25455,N_25628);
or U28612 (N_28612,N_24561,N_26479);
nor U28613 (N_28613,N_26639,N_26830);
nor U28614 (N_28614,N_26104,N_25861);
nor U28615 (N_28615,N_25794,N_24434);
or U28616 (N_28616,N_24759,N_24238);
xnor U28617 (N_28617,N_25383,N_24437);
nor U28618 (N_28618,N_24717,N_26840);
or U28619 (N_28619,N_24452,N_24090);
and U28620 (N_28620,N_26586,N_26024);
nand U28621 (N_28621,N_25814,N_25604);
xor U28622 (N_28622,N_24850,N_24383);
xor U28623 (N_28623,N_25569,N_26475);
nand U28624 (N_28624,N_24861,N_26266);
and U28625 (N_28625,N_24175,N_25244);
xnor U28626 (N_28626,N_25225,N_26029);
nor U28627 (N_28627,N_24690,N_25917);
and U28628 (N_28628,N_26228,N_25214);
xor U28629 (N_28629,N_25066,N_26664);
nor U28630 (N_28630,N_25771,N_26138);
xor U28631 (N_28631,N_26791,N_24621);
nand U28632 (N_28632,N_26305,N_24692);
or U28633 (N_28633,N_26558,N_24405);
or U28634 (N_28634,N_25834,N_24335);
nand U28635 (N_28635,N_24137,N_24637);
nand U28636 (N_28636,N_26842,N_24878);
xnor U28637 (N_28637,N_24059,N_24430);
nor U28638 (N_28638,N_25189,N_26496);
xor U28639 (N_28639,N_25230,N_26021);
nand U28640 (N_28640,N_26947,N_26813);
nand U28641 (N_28641,N_24651,N_26373);
nand U28642 (N_28642,N_24572,N_24435);
and U28643 (N_28643,N_24183,N_24258);
and U28644 (N_28644,N_24615,N_25101);
nor U28645 (N_28645,N_26500,N_24428);
and U28646 (N_28646,N_24853,N_24469);
xnor U28647 (N_28647,N_25694,N_26090);
nor U28648 (N_28648,N_26247,N_26725);
or U28649 (N_28649,N_26593,N_24582);
or U28650 (N_28650,N_26319,N_26176);
and U28651 (N_28651,N_25501,N_25690);
or U28652 (N_28652,N_26505,N_24404);
xnor U28653 (N_28653,N_24700,N_24798);
xor U28654 (N_28654,N_26358,N_25197);
nor U28655 (N_28655,N_26496,N_26876);
or U28656 (N_28656,N_25049,N_25201);
and U28657 (N_28657,N_25333,N_25586);
xor U28658 (N_28658,N_25365,N_26917);
nor U28659 (N_28659,N_26928,N_26128);
nand U28660 (N_28660,N_25638,N_24500);
nand U28661 (N_28661,N_26079,N_24015);
and U28662 (N_28662,N_25878,N_26595);
xnor U28663 (N_28663,N_25598,N_25091);
xor U28664 (N_28664,N_26277,N_24639);
xnor U28665 (N_28665,N_24876,N_25369);
nor U28666 (N_28666,N_26204,N_26348);
nor U28667 (N_28667,N_25337,N_24607);
nand U28668 (N_28668,N_26079,N_25402);
and U28669 (N_28669,N_26728,N_24271);
nor U28670 (N_28670,N_24037,N_26562);
or U28671 (N_28671,N_26980,N_26566);
xor U28672 (N_28672,N_26193,N_25805);
or U28673 (N_28673,N_26266,N_26855);
or U28674 (N_28674,N_24880,N_25757);
xnor U28675 (N_28675,N_26965,N_25233);
nor U28676 (N_28676,N_24252,N_24649);
or U28677 (N_28677,N_26100,N_25282);
and U28678 (N_28678,N_25109,N_25576);
nor U28679 (N_28679,N_24562,N_25274);
nor U28680 (N_28680,N_24505,N_26867);
nor U28681 (N_28681,N_24705,N_24396);
nand U28682 (N_28682,N_25309,N_26879);
or U28683 (N_28683,N_25322,N_26562);
or U28684 (N_28684,N_24171,N_26736);
and U28685 (N_28685,N_26127,N_24979);
and U28686 (N_28686,N_26849,N_24005);
and U28687 (N_28687,N_25531,N_24499);
nand U28688 (N_28688,N_26797,N_25756);
nand U28689 (N_28689,N_25777,N_25214);
nand U28690 (N_28690,N_24037,N_26237);
and U28691 (N_28691,N_24460,N_24894);
xnor U28692 (N_28692,N_24248,N_24544);
nor U28693 (N_28693,N_24521,N_25761);
or U28694 (N_28694,N_26035,N_26570);
or U28695 (N_28695,N_26254,N_24731);
xor U28696 (N_28696,N_24879,N_25702);
nor U28697 (N_28697,N_26311,N_25857);
nor U28698 (N_28698,N_26345,N_26620);
xnor U28699 (N_28699,N_24264,N_24135);
or U28700 (N_28700,N_25518,N_24264);
nor U28701 (N_28701,N_24256,N_25033);
nor U28702 (N_28702,N_26408,N_25505);
or U28703 (N_28703,N_24941,N_26634);
or U28704 (N_28704,N_24794,N_25507);
nor U28705 (N_28705,N_24031,N_24667);
xnor U28706 (N_28706,N_24295,N_26535);
nor U28707 (N_28707,N_24485,N_25555);
xnor U28708 (N_28708,N_24434,N_25239);
nand U28709 (N_28709,N_24314,N_25161);
nand U28710 (N_28710,N_26621,N_26410);
or U28711 (N_28711,N_25232,N_24936);
xor U28712 (N_28712,N_24203,N_24595);
nand U28713 (N_28713,N_26166,N_26751);
or U28714 (N_28714,N_25102,N_25492);
nand U28715 (N_28715,N_24132,N_26128);
and U28716 (N_28716,N_26326,N_25279);
xor U28717 (N_28717,N_24764,N_24439);
and U28718 (N_28718,N_26354,N_24795);
or U28719 (N_28719,N_25835,N_24269);
nor U28720 (N_28720,N_25506,N_26937);
or U28721 (N_28721,N_25268,N_26281);
nor U28722 (N_28722,N_25607,N_25092);
and U28723 (N_28723,N_25634,N_25264);
nor U28724 (N_28724,N_24689,N_26485);
or U28725 (N_28725,N_24741,N_24787);
xor U28726 (N_28726,N_24739,N_26631);
nand U28727 (N_28727,N_26845,N_25118);
and U28728 (N_28728,N_25323,N_24148);
nor U28729 (N_28729,N_25103,N_25666);
or U28730 (N_28730,N_24279,N_25310);
nand U28731 (N_28731,N_24253,N_25265);
xnor U28732 (N_28732,N_25950,N_24222);
xnor U28733 (N_28733,N_24204,N_25201);
nor U28734 (N_28734,N_24996,N_25245);
or U28735 (N_28735,N_25620,N_26108);
nor U28736 (N_28736,N_26424,N_24182);
and U28737 (N_28737,N_24810,N_26538);
or U28738 (N_28738,N_26510,N_24846);
xor U28739 (N_28739,N_26742,N_24466);
nand U28740 (N_28740,N_24014,N_25819);
nor U28741 (N_28741,N_26610,N_25926);
or U28742 (N_28742,N_24074,N_25999);
or U28743 (N_28743,N_26300,N_24381);
and U28744 (N_28744,N_24052,N_25753);
nand U28745 (N_28745,N_26933,N_26462);
nand U28746 (N_28746,N_25737,N_26873);
nand U28747 (N_28747,N_24410,N_26929);
or U28748 (N_28748,N_24882,N_25097);
or U28749 (N_28749,N_25977,N_26382);
and U28750 (N_28750,N_25975,N_24503);
or U28751 (N_28751,N_26215,N_26633);
or U28752 (N_28752,N_24369,N_24842);
nor U28753 (N_28753,N_26781,N_24306);
or U28754 (N_28754,N_26956,N_25612);
or U28755 (N_28755,N_24149,N_24202);
nor U28756 (N_28756,N_25443,N_24957);
nand U28757 (N_28757,N_26710,N_26179);
xnor U28758 (N_28758,N_24004,N_24894);
xor U28759 (N_28759,N_24525,N_25144);
and U28760 (N_28760,N_26116,N_26369);
nand U28761 (N_28761,N_25194,N_24277);
and U28762 (N_28762,N_26971,N_25680);
nor U28763 (N_28763,N_24928,N_25257);
and U28764 (N_28764,N_26696,N_24286);
nand U28765 (N_28765,N_25159,N_24289);
or U28766 (N_28766,N_24140,N_24435);
xor U28767 (N_28767,N_24814,N_26267);
nor U28768 (N_28768,N_26205,N_26151);
nor U28769 (N_28769,N_24609,N_24488);
and U28770 (N_28770,N_26033,N_24684);
nor U28771 (N_28771,N_25824,N_25686);
nor U28772 (N_28772,N_24231,N_24180);
nor U28773 (N_28773,N_26947,N_25798);
and U28774 (N_28774,N_26653,N_25831);
or U28775 (N_28775,N_26003,N_25705);
or U28776 (N_28776,N_24538,N_24451);
and U28777 (N_28777,N_26015,N_24800);
or U28778 (N_28778,N_24897,N_25315);
nand U28779 (N_28779,N_26225,N_26437);
and U28780 (N_28780,N_24044,N_24819);
or U28781 (N_28781,N_25076,N_26300);
or U28782 (N_28782,N_25072,N_24286);
or U28783 (N_28783,N_24297,N_25757);
or U28784 (N_28784,N_24895,N_25452);
and U28785 (N_28785,N_24134,N_24115);
nor U28786 (N_28786,N_24000,N_24254);
and U28787 (N_28787,N_25959,N_24571);
xor U28788 (N_28788,N_26530,N_25670);
and U28789 (N_28789,N_24672,N_24853);
or U28790 (N_28790,N_25610,N_24157);
nand U28791 (N_28791,N_26320,N_26510);
and U28792 (N_28792,N_25252,N_26861);
nor U28793 (N_28793,N_26458,N_26571);
nor U28794 (N_28794,N_24534,N_25495);
xnor U28795 (N_28795,N_26605,N_24075);
xnor U28796 (N_28796,N_24232,N_25012);
or U28797 (N_28797,N_25185,N_25239);
xnor U28798 (N_28798,N_26791,N_24121);
or U28799 (N_28799,N_25295,N_25453);
nor U28800 (N_28800,N_26548,N_26352);
nor U28801 (N_28801,N_24515,N_26273);
and U28802 (N_28802,N_26970,N_24638);
xor U28803 (N_28803,N_25025,N_25796);
nand U28804 (N_28804,N_26788,N_25817);
nor U28805 (N_28805,N_25439,N_24251);
nand U28806 (N_28806,N_24717,N_24102);
nor U28807 (N_28807,N_25767,N_25228);
xor U28808 (N_28808,N_24251,N_25406);
or U28809 (N_28809,N_24588,N_25129);
nand U28810 (N_28810,N_25428,N_25763);
nand U28811 (N_28811,N_24217,N_25456);
nor U28812 (N_28812,N_26411,N_26787);
xor U28813 (N_28813,N_24241,N_25779);
xnor U28814 (N_28814,N_25448,N_26820);
xor U28815 (N_28815,N_26009,N_25284);
and U28816 (N_28816,N_25927,N_25996);
nor U28817 (N_28817,N_24763,N_26723);
or U28818 (N_28818,N_24522,N_24564);
nand U28819 (N_28819,N_24471,N_24722);
nor U28820 (N_28820,N_26931,N_25379);
nor U28821 (N_28821,N_26351,N_24898);
nor U28822 (N_28822,N_25988,N_26199);
nor U28823 (N_28823,N_26603,N_25744);
nor U28824 (N_28824,N_24523,N_24163);
nor U28825 (N_28825,N_24512,N_26026);
or U28826 (N_28826,N_24122,N_25534);
nor U28827 (N_28827,N_26476,N_26295);
xnor U28828 (N_28828,N_26845,N_25020);
nor U28829 (N_28829,N_24221,N_25159);
nand U28830 (N_28830,N_26595,N_24827);
nor U28831 (N_28831,N_25203,N_25929);
nor U28832 (N_28832,N_24533,N_24567);
nor U28833 (N_28833,N_24979,N_24721);
or U28834 (N_28834,N_26331,N_26068);
nand U28835 (N_28835,N_26023,N_26045);
nand U28836 (N_28836,N_25877,N_26531);
nand U28837 (N_28837,N_24166,N_24440);
xnor U28838 (N_28838,N_24391,N_26733);
and U28839 (N_28839,N_25930,N_24571);
or U28840 (N_28840,N_25940,N_26445);
and U28841 (N_28841,N_25218,N_24778);
and U28842 (N_28842,N_26593,N_24549);
xor U28843 (N_28843,N_24613,N_24333);
xor U28844 (N_28844,N_24441,N_25072);
nand U28845 (N_28845,N_26274,N_24291);
xor U28846 (N_28846,N_25905,N_24085);
and U28847 (N_28847,N_26308,N_25490);
and U28848 (N_28848,N_26869,N_24501);
nand U28849 (N_28849,N_26591,N_26436);
or U28850 (N_28850,N_24938,N_26435);
nor U28851 (N_28851,N_26603,N_24227);
nor U28852 (N_28852,N_26975,N_25956);
nor U28853 (N_28853,N_24431,N_25545);
nand U28854 (N_28854,N_26829,N_24589);
nor U28855 (N_28855,N_24248,N_26291);
xor U28856 (N_28856,N_24560,N_26765);
and U28857 (N_28857,N_26072,N_26396);
nor U28858 (N_28858,N_26315,N_24089);
nor U28859 (N_28859,N_24464,N_25188);
nand U28860 (N_28860,N_25791,N_25395);
nor U28861 (N_28861,N_26695,N_26999);
nor U28862 (N_28862,N_24038,N_26868);
or U28863 (N_28863,N_25015,N_26055);
nor U28864 (N_28864,N_25390,N_24070);
nor U28865 (N_28865,N_26997,N_26336);
or U28866 (N_28866,N_24099,N_24497);
xor U28867 (N_28867,N_24009,N_24112);
or U28868 (N_28868,N_24982,N_25880);
nand U28869 (N_28869,N_24863,N_24734);
nor U28870 (N_28870,N_26019,N_24547);
and U28871 (N_28871,N_24428,N_24857);
nand U28872 (N_28872,N_24230,N_25771);
nand U28873 (N_28873,N_25780,N_26880);
nand U28874 (N_28874,N_26442,N_25375);
and U28875 (N_28875,N_24781,N_26289);
xor U28876 (N_28876,N_24288,N_26948);
xor U28877 (N_28877,N_25974,N_25103);
and U28878 (N_28878,N_25490,N_24459);
xnor U28879 (N_28879,N_25403,N_25931);
nand U28880 (N_28880,N_25550,N_24642);
nor U28881 (N_28881,N_24753,N_26266);
xnor U28882 (N_28882,N_26644,N_25277);
xnor U28883 (N_28883,N_26807,N_24063);
nand U28884 (N_28884,N_24670,N_26149);
and U28885 (N_28885,N_26691,N_24317);
nand U28886 (N_28886,N_24952,N_26550);
xor U28887 (N_28887,N_24558,N_25997);
nand U28888 (N_28888,N_25865,N_25499);
xor U28889 (N_28889,N_26579,N_25611);
nand U28890 (N_28890,N_24316,N_24134);
nand U28891 (N_28891,N_26134,N_24751);
or U28892 (N_28892,N_25372,N_24723);
xnor U28893 (N_28893,N_25288,N_26827);
xnor U28894 (N_28894,N_26625,N_25176);
xor U28895 (N_28895,N_24710,N_26958);
and U28896 (N_28896,N_24319,N_26399);
and U28897 (N_28897,N_24960,N_26879);
nand U28898 (N_28898,N_24534,N_25205);
nand U28899 (N_28899,N_25435,N_25221);
or U28900 (N_28900,N_25897,N_26250);
or U28901 (N_28901,N_24428,N_26047);
nand U28902 (N_28902,N_24821,N_24387);
nand U28903 (N_28903,N_24275,N_24674);
xor U28904 (N_28904,N_25584,N_25039);
xnor U28905 (N_28905,N_26975,N_25289);
nand U28906 (N_28906,N_24219,N_25167);
nand U28907 (N_28907,N_24523,N_25400);
xor U28908 (N_28908,N_26734,N_26524);
xor U28909 (N_28909,N_25633,N_25172);
and U28910 (N_28910,N_26534,N_25460);
and U28911 (N_28911,N_25089,N_26256);
and U28912 (N_28912,N_25479,N_26053);
nand U28913 (N_28913,N_25171,N_25415);
xnor U28914 (N_28914,N_26866,N_26149);
and U28915 (N_28915,N_24574,N_24795);
and U28916 (N_28916,N_25706,N_24034);
nor U28917 (N_28917,N_25995,N_24640);
and U28918 (N_28918,N_26486,N_25600);
or U28919 (N_28919,N_26908,N_26777);
xor U28920 (N_28920,N_26448,N_26089);
nor U28921 (N_28921,N_25188,N_24106);
or U28922 (N_28922,N_25352,N_25865);
nand U28923 (N_28923,N_26288,N_25576);
or U28924 (N_28924,N_26583,N_26870);
or U28925 (N_28925,N_26467,N_24524);
and U28926 (N_28926,N_24250,N_24769);
xnor U28927 (N_28927,N_25787,N_24717);
nor U28928 (N_28928,N_25629,N_24692);
xor U28929 (N_28929,N_25004,N_25631);
xor U28930 (N_28930,N_24734,N_24048);
nor U28931 (N_28931,N_25459,N_25643);
nand U28932 (N_28932,N_26347,N_25426);
nand U28933 (N_28933,N_26148,N_25166);
nor U28934 (N_28934,N_24317,N_24336);
nand U28935 (N_28935,N_25328,N_26786);
nand U28936 (N_28936,N_25763,N_24549);
or U28937 (N_28937,N_25115,N_24645);
and U28938 (N_28938,N_25530,N_24257);
or U28939 (N_28939,N_26428,N_25608);
and U28940 (N_28940,N_24174,N_25229);
nor U28941 (N_28941,N_26143,N_25489);
and U28942 (N_28942,N_26497,N_26379);
or U28943 (N_28943,N_26333,N_24230);
and U28944 (N_28944,N_24582,N_25965);
nand U28945 (N_28945,N_26042,N_24897);
and U28946 (N_28946,N_25678,N_24898);
or U28947 (N_28947,N_26024,N_24603);
and U28948 (N_28948,N_25603,N_24352);
xnor U28949 (N_28949,N_25067,N_24511);
or U28950 (N_28950,N_26773,N_25797);
and U28951 (N_28951,N_24552,N_26867);
xor U28952 (N_28952,N_26857,N_26916);
nand U28953 (N_28953,N_24173,N_25152);
or U28954 (N_28954,N_26920,N_24305);
or U28955 (N_28955,N_24942,N_24946);
and U28956 (N_28956,N_26033,N_26035);
nor U28957 (N_28957,N_25109,N_24519);
nor U28958 (N_28958,N_25951,N_25526);
nor U28959 (N_28959,N_25126,N_25653);
xnor U28960 (N_28960,N_24807,N_26423);
xnor U28961 (N_28961,N_26582,N_24142);
xor U28962 (N_28962,N_26964,N_24999);
xnor U28963 (N_28963,N_25376,N_25950);
xnor U28964 (N_28964,N_26839,N_24047);
or U28965 (N_28965,N_25196,N_25667);
nor U28966 (N_28966,N_24801,N_26112);
and U28967 (N_28967,N_25014,N_25575);
xnor U28968 (N_28968,N_26892,N_25686);
nand U28969 (N_28969,N_25548,N_26806);
and U28970 (N_28970,N_24328,N_24474);
nand U28971 (N_28971,N_24323,N_26247);
nand U28972 (N_28972,N_25968,N_26744);
and U28973 (N_28973,N_25644,N_25646);
and U28974 (N_28974,N_24691,N_25196);
nor U28975 (N_28975,N_24396,N_24084);
nand U28976 (N_28976,N_26993,N_25839);
and U28977 (N_28977,N_24197,N_26125);
nand U28978 (N_28978,N_25094,N_24462);
or U28979 (N_28979,N_24501,N_24886);
nand U28980 (N_28980,N_24460,N_25934);
nor U28981 (N_28981,N_25943,N_26864);
nand U28982 (N_28982,N_24315,N_25406);
or U28983 (N_28983,N_25026,N_26885);
nand U28984 (N_28984,N_24806,N_26898);
xnor U28985 (N_28985,N_25429,N_25473);
and U28986 (N_28986,N_24602,N_24084);
or U28987 (N_28987,N_26376,N_24776);
nand U28988 (N_28988,N_26542,N_24207);
nor U28989 (N_28989,N_26639,N_24928);
nor U28990 (N_28990,N_26047,N_25721);
and U28991 (N_28991,N_25564,N_24336);
nand U28992 (N_28992,N_24339,N_24752);
xnor U28993 (N_28993,N_24182,N_24063);
nand U28994 (N_28994,N_24587,N_25168);
nor U28995 (N_28995,N_25584,N_24645);
nor U28996 (N_28996,N_24813,N_25530);
nor U28997 (N_28997,N_25225,N_26280);
nand U28998 (N_28998,N_25476,N_24185);
or U28999 (N_28999,N_26000,N_24315);
nand U29000 (N_29000,N_25545,N_26717);
nor U29001 (N_29001,N_25642,N_24777);
nor U29002 (N_29002,N_26348,N_24754);
nor U29003 (N_29003,N_24558,N_25508);
nand U29004 (N_29004,N_25385,N_26643);
or U29005 (N_29005,N_24788,N_26843);
nand U29006 (N_29006,N_25531,N_26836);
xnor U29007 (N_29007,N_25598,N_26868);
nor U29008 (N_29008,N_26518,N_25296);
xnor U29009 (N_29009,N_24100,N_25770);
or U29010 (N_29010,N_26669,N_25889);
nand U29011 (N_29011,N_24867,N_25756);
xnor U29012 (N_29012,N_24489,N_26152);
and U29013 (N_29013,N_24370,N_24348);
nor U29014 (N_29014,N_26276,N_24967);
or U29015 (N_29015,N_24229,N_25040);
and U29016 (N_29016,N_24240,N_26191);
nand U29017 (N_29017,N_26608,N_24009);
nand U29018 (N_29018,N_26998,N_26596);
and U29019 (N_29019,N_25402,N_24241);
and U29020 (N_29020,N_25388,N_26420);
nand U29021 (N_29021,N_26904,N_25899);
or U29022 (N_29022,N_25219,N_25405);
or U29023 (N_29023,N_25863,N_25918);
nand U29024 (N_29024,N_26922,N_25261);
nor U29025 (N_29025,N_26281,N_25932);
and U29026 (N_29026,N_26198,N_25457);
nor U29027 (N_29027,N_24840,N_26333);
nand U29028 (N_29028,N_26685,N_24391);
and U29029 (N_29029,N_25846,N_25583);
nand U29030 (N_29030,N_24727,N_26646);
nand U29031 (N_29031,N_26405,N_24005);
nor U29032 (N_29032,N_25105,N_24507);
nor U29033 (N_29033,N_25501,N_26115);
or U29034 (N_29034,N_26574,N_25561);
and U29035 (N_29035,N_24690,N_26475);
nor U29036 (N_29036,N_25706,N_24995);
and U29037 (N_29037,N_26617,N_26124);
xnor U29038 (N_29038,N_25728,N_26893);
xor U29039 (N_29039,N_25231,N_24073);
nand U29040 (N_29040,N_25575,N_26470);
nor U29041 (N_29041,N_24694,N_24693);
and U29042 (N_29042,N_25999,N_25019);
and U29043 (N_29043,N_25023,N_24611);
and U29044 (N_29044,N_25394,N_26727);
xnor U29045 (N_29045,N_24548,N_24438);
xnor U29046 (N_29046,N_25552,N_26816);
nor U29047 (N_29047,N_24428,N_25281);
nand U29048 (N_29048,N_25726,N_24100);
xnor U29049 (N_29049,N_25201,N_24199);
or U29050 (N_29050,N_26510,N_26249);
and U29051 (N_29051,N_24962,N_26876);
xnor U29052 (N_29052,N_25274,N_26354);
or U29053 (N_29053,N_26738,N_24305);
nor U29054 (N_29054,N_26618,N_24798);
nand U29055 (N_29055,N_25847,N_24946);
or U29056 (N_29056,N_26716,N_26237);
and U29057 (N_29057,N_24599,N_24868);
xor U29058 (N_29058,N_24925,N_24671);
and U29059 (N_29059,N_25677,N_24294);
nor U29060 (N_29060,N_24860,N_26794);
xnor U29061 (N_29061,N_24609,N_26577);
nor U29062 (N_29062,N_26214,N_26844);
or U29063 (N_29063,N_24327,N_24404);
and U29064 (N_29064,N_26655,N_25029);
and U29065 (N_29065,N_24523,N_25218);
nand U29066 (N_29066,N_26476,N_25712);
and U29067 (N_29067,N_25594,N_26885);
nor U29068 (N_29068,N_25196,N_25724);
and U29069 (N_29069,N_26051,N_25682);
or U29070 (N_29070,N_25819,N_25349);
or U29071 (N_29071,N_26885,N_25729);
nand U29072 (N_29072,N_24908,N_26954);
and U29073 (N_29073,N_25196,N_24443);
nand U29074 (N_29074,N_24372,N_25476);
xnor U29075 (N_29075,N_25455,N_25764);
or U29076 (N_29076,N_26762,N_25082);
xnor U29077 (N_29077,N_26365,N_26437);
and U29078 (N_29078,N_25186,N_26706);
nor U29079 (N_29079,N_24830,N_26672);
xor U29080 (N_29080,N_24365,N_24844);
nand U29081 (N_29081,N_24217,N_24879);
nand U29082 (N_29082,N_26838,N_24098);
or U29083 (N_29083,N_24864,N_24418);
nand U29084 (N_29084,N_25385,N_24350);
nand U29085 (N_29085,N_24766,N_25211);
or U29086 (N_29086,N_26778,N_25294);
or U29087 (N_29087,N_26790,N_26338);
xor U29088 (N_29088,N_26888,N_26445);
and U29089 (N_29089,N_25254,N_25414);
and U29090 (N_29090,N_26419,N_25531);
and U29091 (N_29091,N_26020,N_26146);
and U29092 (N_29092,N_25273,N_25574);
or U29093 (N_29093,N_24707,N_24526);
xnor U29094 (N_29094,N_24846,N_25515);
nor U29095 (N_29095,N_25594,N_24201);
and U29096 (N_29096,N_24905,N_25117);
or U29097 (N_29097,N_24846,N_24019);
and U29098 (N_29098,N_24515,N_25812);
nand U29099 (N_29099,N_25746,N_26498);
and U29100 (N_29100,N_26119,N_26190);
nor U29101 (N_29101,N_26670,N_24903);
nor U29102 (N_29102,N_24040,N_24274);
nand U29103 (N_29103,N_25024,N_25308);
xor U29104 (N_29104,N_25345,N_25778);
and U29105 (N_29105,N_24467,N_25945);
nor U29106 (N_29106,N_25108,N_25251);
xnor U29107 (N_29107,N_26896,N_24397);
nand U29108 (N_29108,N_24851,N_26300);
xor U29109 (N_29109,N_26429,N_24953);
nand U29110 (N_29110,N_25943,N_24822);
nand U29111 (N_29111,N_24853,N_24629);
xor U29112 (N_29112,N_26986,N_26442);
or U29113 (N_29113,N_25491,N_26609);
or U29114 (N_29114,N_26152,N_25391);
nor U29115 (N_29115,N_26395,N_26725);
or U29116 (N_29116,N_25807,N_26008);
nor U29117 (N_29117,N_25308,N_25137);
or U29118 (N_29118,N_24040,N_25368);
or U29119 (N_29119,N_26264,N_25485);
nor U29120 (N_29120,N_24742,N_24895);
xnor U29121 (N_29121,N_26011,N_24732);
and U29122 (N_29122,N_24941,N_24237);
or U29123 (N_29123,N_26012,N_25586);
and U29124 (N_29124,N_25242,N_24300);
and U29125 (N_29125,N_24785,N_25959);
nand U29126 (N_29126,N_26604,N_24786);
or U29127 (N_29127,N_24893,N_24800);
or U29128 (N_29128,N_24107,N_24633);
nor U29129 (N_29129,N_25001,N_26941);
nor U29130 (N_29130,N_24127,N_26629);
and U29131 (N_29131,N_24946,N_26988);
nor U29132 (N_29132,N_26394,N_24925);
xnor U29133 (N_29133,N_24363,N_26868);
and U29134 (N_29134,N_26621,N_26251);
nand U29135 (N_29135,N_25346,N_25907);
nand U29136 (N_29136,N_25267,N_24462);
or U29137 (N_29137,N_26373,N_25795);
or U29138 (N_29138,N_26160,N_24777);
nor U29139 (N_29139,N_24140,N_26890);
and U29140 (N_29140,N_24975,N_24475);
nand U29141 (N_29141,N_25681,N_24730);
and U29142 (N_29142,N_26189,N_26393);
and U29143 (N_29143,N_24493,N_25085);
or U29144 (N_29144,N_24047,N_24255);
xor U29145 (N_29145,N_25375,N_26484);
and U29146 (N_29146,N_25496,N_25629);
or U29147 (N_29147,N_25995,N_26407);
or U29148 (N_29148,N_25783,N_25069);
nand U29149 (N_29149,N_26077,N_25194);
nor U29150 (N_29150,N_26230,N_26008);
xnor U29151 (N_29151,N_25782,N_26597);
xnor U29152 (N_29152,N_25125,N_26121);
and U29153 (N_29153,N_26168,N_24012);
nor U29154 (N_29154,N_24273,N_26723);
nor U29155 (N_29155,N_25532,N_26350);
xor U29156 (N_29156,N_26212,N_25590);
or U29157 (N_29157,N_26504,N_24144);
and U29158 (N_29158,N_26275,N_24390);
nor U29159 (N_29159,N_25432,N_26803);
nand U29160 (N_29160,N_26276,N_25271);
or U29161 (N_29161,N_24082,N_26478);
nand U29162 (N_29162,N_26731,N_26237);
nor U29163 (N_29163,N_26879,N_25451);
nand U29164 (N_29164,N_26081,N_25598);
and U29165 (N_29165,N_25328,N_24795);
or U29166 (N_29166,N_24977,N_24025);
xnor U29167 (N_29167,N_24318,N_26085);
nand U29168 (N_29168,N_26267,N_26872);
nor U29169 (N_29169,N_26194,N_24374);
nand U29170 (N_29170,N_26496,N_24046);
or U29171 (N_29171,N_25452,N_24575);
or U29172 (N_29172,N_25293,N_26876);
and U29173 (N_29173,N_24886,N_26686);
or U29174 (N_29174,N_26401,N_25646);
or U29175 (N_29175,N_26387,N_25161);
or U29176 (N_29176,N_26590,N_26925);
xor U29177 (N_29177,N_24845,N_25031);
nor U29178 (N_29178,N_26983,N_25642);
xnor U29179 (N_29179,N_25763,N_25178);
nand U29180 (N_29180,N_25170,N_25856);
nand U29181 (N_29181,N_24415,N_24804);
nand U29182 (N_29182,N_24473,N_24613);
or U29183 (N_29183,N_25135,N_24080);
xnor U29184 (N_29184,N_25736,N_25335);
nand U29185 (N_29185,N_24428,N_24107);
nor U29186 (N_29186,N_25668,N_26926);
or U29187 (N_29187,N_26754,N_25773);
or U29188 (N_29188,N_25520,N_25702);
and U29189 (N_29189,N_26151,N_24734);
nor U29190 (N_29190,N_24841,N_24243);
nor U29191 (N_29191,N_25503,N_26588);
and U29192 (N_29192,N_26061,N_26267);
xnor U29193 (N_29193,N_25305,N_25377);
or U29194 (N_29194,N_24658,N_26668);
nor U29195 (N_29195,N_24229,N_24292);
nand U29196 (N_29196,N_25543,N_24271);
xor U29197 (N_29197,N_25173,N_26968);
xnor U29198 (N_29198,N_25959,N_24582);
xnor U29199 (N_29199,N_26011,N_26379);
nand U29200 (N_29200,N_24154,N_26870);
nor U29201 (N_29201,N_26560,N_26493);
nor U29202 (N_29202,N_25787,N_25275);
nor U29203 (N_29203,N_25728,N_24427);
or U29204 (N_29204,N_24907,N_24451);
or U29205 (N_29205,N_26481,N_24622);
nor U29206 (N_29206,N_24426,N_25600);
nor U29207 (N_29207,N_25320,N_24827);
nor U29208 (N_29208,N_25983,N_25144);
xnor U29209 (N_29209,N_26910,N_25229);
and U29210 (N_29210,N_24269,N_24713);
nor U29211 (N_29211,N_24114,N_24307);
nor U29212 (N_29212,N_25344,N_24173);
and U29213 (N_29213,N_25758,N_26574);
or U29214 (N_29214,N_26256,N_24245);
xor U29215 (N_29215,N_25482,N_25960);
xnor U29216 (N_29216,N_24881,N_24945);
nor U29217 (N_29217,N_26439,N_25308);
or U29218 (N_29218,N_25953,N_24511);
nor U29219 (N_29219,N_25568,N_25578);
nand U29220 (N_29220,N_24272,N_26469);
nand U29221 (N_29221,N_26200,N_24833);
and U29222 (N_29222,N_24398,N_26298);
or U29223 (N_29223,N_24147,N_25606);
nand U29224 (N_29224,N_26156,N_24541);
or U29225 (N_29225,N_24694,N_26168);
and U29226 (N_29226,N_24357,N_25854);
xor U29227 (N_29227,N_24165,N_26446);
xnor U29228 (N_29228,N_25223,N_24711);
nand U29229 (N_29229,N_26600,N_25966);
nor U29230 (N_29230,N_26437,N_25024);
nand U29231 (N_29231,N_25320,N_24566);
xnor U29232 (N_29232,N_26008,N_24203);
nor U29233 (N_29233,N_26634,N_26576);
xnor U29234 (N_29234,N_26731,N_26784);
xor U29235 (N_29235,N_25547,N_26152);
or U29236 (N_29236,N_24240,N_26043);
nand U29237 (N_29237,N_25148,N_25311);
nand U29238 (N_29238,N_24742,N_24721);
nor U29239 (N_29239,N_25914,N_26626);
nor U29240 (N_29240,N_26213,N_26980);
nor U29241 (N_29241,N_25119,N_25479);
xnor U29242 (N_29242,N_25016,N_26220);
or U29243 (N_29243,N_26066,N_24631);
and U29244 (N_29244,N_25893,N_24133);
nand U29245 (N_29245,N_26470,N_26947);
xor U29246 (N_29246,N_24618,N_26537);
nand U29247 (N_29247,N_26356,N_24722);
nand U29248 (N_29248,N_26710,N_25840);
xnor U29249 (N_29249,N_24496,N_24276);
or U29250 (N_29250,N_26804,N_25854);
nor U29251 (N_29251,N_25419,N_24316);
and U29252 (N_29252,N_26631,N_25757);
nor U29253 (N_29253,N_25833,N_24843);
xnor U29254 (N_29254,N_26363,N_24716);
and U29255 (N_29255,N_25567,N_25145);
or U29256 (N_29256,N_24316,N_26225);
xnor U29257 (N_29257,N_25986,N_26948);
or U29258 (N_29258,N_25982,N_24691);
xnor U29259 (N_29259,N_25284,N_26273);
nand U29260 (N_29260,N_24506,N_26774);
nor U29261 (N_29261,N_25112,N_24592);
nor U29262 (N_29262,N_26563,N_26630);
nand U29263 (N_29263,N_25067,N_25006);
nand U29264 (N_29264,N_24836,N_26360);
or U29265 (N_29265,N_24612,N_26101);
and U29266 (N_29266,N_24151,N_26953);
nand U29267 (N_29267,N_25829,N_24912);
or U29268 (N_29268,N_26286,N_24332);
and U29269 (N_29269,N_24183,N_26614);
xor U29270 (N_29270,N_25686,N_26150);
nor U29271 (N_29271,N_26184,N_25303);
and U29272 (N_29272,N_25485,N_24812);
nand U29273 (N_29273,N_24035,N_26964);
or U29274 (N_29274,N_25444,N_26226);
xnor U29275 (N_29275,N_25893,N_25226);
nor U29276 (N_29276,N_24376,N_24393);
or U29277 (N_29277,N_26949,N_24681);
or U29278 (N_29278,N_24634,N_26400);
xor U29279 (N_29279,N_25954,N_24459);
xnor U29280 (N_29280,N_24562,N_24147);
xnor U29281 (N_29281,N_24712,N_24276);
xor U29282 (N_29282,N_24427,N_24946);
and U29283 (N_29283,N_25962,N_25609);
xnor U29284 (N_29284,N_26267,N_25468);
nand U29285 (N_29285,N_26390,N_26289);
or U29286 (N_29286,N_26382,N_24968);
and U29287 (N_29287,N_26653,N_25508);
and U29288 (N_29288,N_26658,N_26015);
or U29289 (N_29289,N_25123,N_26024);
nor U29290 (N_29290,N_25116,N_26247);
nand U29291 (N_29291,N_25908,N_24818);
nand U29292 (N_29292,N_25377,N_26620);
nor U29293 (N_29293,N_24260,N_25872);
nand U29294 (N_29294,N_26323,N_25730);
xor U29295 (N_29295,N_24590,N_25064);
and U29296 (N_29296,N_24427,N_25315);
or U29297 (N_29297,N_24460,N_24459);
or U29298 (N_29298,N_26958,N_24796);
and U29299 (N_29299,N_25087,N_24255);
nor U29300 (N_29300,N_25644,N_25072);
nand U29301 (N_29301,N_25124,N_24875);
xor U29302 (N_29302,N_25515,N_24879);
nand U29303 (N_29303,N_24037,N_25389);
nand U29304 (N_29304,N_26722,N_25449);
nor U29305 (N_29305,N_24124,N_24018);
and U29306 (N_29306,N_26006,N_24156);
or U29307 (N_29307,N_24747,N_24697);
nor U29308 (N_29308,N_26952,N_26037);
nand U29309 (N_29309,N_24269,N_24615);
nor U29310 (N_29310,N_25341,N_24475);
nor U29311 (N_29311,N_25920,N_26545);
or U29312 (N_29312,N_24668,N_25020);
xnor U29313 (N_29313,N_26351,N_26093);
nand U29314 (N_29314,N_24712,N_24314);
or U29315 (N_29315,N_26901,N_26985);
nor U29316 (N_29316,N_25307,N_26701);
xor U29317 (N_29317,N_26501,N_26418);
or U29318 (N_29318,N_24067,N_26315);
and U29319 (N_29319,N_25204,N_25507);
nor U29320 (N_29320,N_25957,N_24727);
xor U29321 (N_29321,N_25458,N_26128);
or U29322 (N_29322,N_25320,N_26236);
and U29323 (N_29323,N_26191,N_26247);
nor U29324 (N_29324,N_25562,N_24013);
and U29325 (N_29325,N_25271,N_24254);
xor U29326 (N_29326,N_24055,N_25230);
xor U29327 (N_29327,N_24501,N_25775);
nor U29328 (N_29328,N_25457,N_24805);
xnor U29329 (N_29329,N_26376,N_26544);
nor U29330 (N_29330,N_25409,N_24008);
nand U29331 (N_29331,N_26639,N_25173);
nand U29332 (N_29332,N_24372,N_25585);
and U29333 (N_29333,N_24192,N_26704);
nand U29334 (N_29334,N_25046,N_24365);
xnor U29335 (N_29335,N_26695,N_24052);
and U29336 (N_29336,N_24254,N_26052);
nand U29337 (N_29337,N_25828,N_25577);
xor U29338 (N_29338,N_25180,N_26533);
or U29339 (N_29339,N_26530,N_24595);
or U29340 (N_29340,N_24496,N_25916);
nand U29341 (N_29341,N_24972,N_26021);
or U29342 (N_29342,N_26893,N_24204);
xnor U29343 (N_29343,N_25452,N_26170);
nor U29344 (N_29344,N_26837,N_26931);
nor U29345 (N_29345,N_25573,N_26395);
and U29346 (N_29346,N_25115,N_25449);
nor U29347 (N_29347,N_24193,N_24680);
or U29348 (N_29348,N_26869,N_25654);
nor U29349 (N_29349,N_24564,N_26875);
nor U29350 (N_29350,N_26925,N_26692);
or U29351 (N_29351,N_26988,N_25928);
or U29352 (N_29352,N_24760,N_24709);
nand U29353 (N_29353,N_24806,N_24551);
or U29354 (N_29354,N_24993,N_24286);
xor U29355 (N_29355,N_25482,N_25651);
nand U29356 (N_29356,N_26920,N_26114);
nor U29357 (N_29357,N_25929,N_24956);
nand U29358 (N_29358,N_26223,N_24917);
or U29359 (N_29359,N_26439,N_24996);
or U29360 (N_29360,N_25994,N_26003);
xor U29361 (N_29361,N_24728,N_25607);
xnor U29362 (N_29362,N_24868,N_25656);
xnor U29363 (N_29363,N_25215,N_24272);
xnor U29364 (N_29364,N_24072,N_24313);
nor U29365 (N_29365,N_26442,N_25028);
or U29366 (N_29366,N_24037,N_25183);
xor U29367 (N_29367,N_24101,N_24195);
or U29368 (N_29368,N_24889,N_26876);
xnor U29369 (N_29369,N_25700,N_24048);
and U29370 (N_29370,N_25003,N_26167);
xnor U29371 (N_29371,N_25788,N_24298);
or U29372 (N_29372,N_25045,N_26454);
nand U29373 (N_29373,N_26225,N_24289);
and U29374 (N_29374,N_25062,N_25633);
or U29375 (N_29375,N_25437,N_26149);
nor U29376 (N_29376,N_26781,N_26174);
nand U29377 (N_29377,N_25734,N_24565);
and U29378 (N_29378,N_24737,N_24231);
and U29379 (N_29379,N_26532,N_24345);
xnor U29380 (N_29380,N_26242,N_24286);
or U29381 (N_29381,N_24721,N_24105);
nand U29382 (N_29382,N_25762,N_25500);
xor U29383 (N_29383,N_25586,N_26895);
and U29384 (N_29384,N_26268,N_26731);
nor U29385 (N_29385,N_26310,N_25954);
and U29386 (N_29386,N_25372,N_25874);
xnor U29387 (N_29387,N_24207,N_25381);
nand U29388 (N_29388,N_24108,N_26823);
nor U29389 (N_29389,N_26306,N_24561);
nor U29390 (N_29390,N_24858,N_26226);
and U29391 (N_29391,N_25058,N_25496);
nor U29392 (N_29392,N_25982,N_24428);
or U29393 (N_29393,N_25471,N_24236);
nor U29394 (N_29394,N_26472,N_25496);
and U29395 (N_29395,N_25956,N_26863);
nand U29396 (N_29396,N_25278,N_24932);
and U29397 (N_29397,N_25289,N_25106);
and U29398 (N_29398,N_25272,N_25539);
or U29399 (N_29399,N_26967,N_25036);
or U29400 (N_29400,N_26064,N_26651);
and U29401 (N_29401,N_26790,N_24013);
or U29402 (N_29402,N_24589,N_24939);
nand U29403 (N_29403,N_24365,N_24405);
xnor U29404 (N_29404,N_24214,N_24671);
or U29405 (N_29405,N_25638,N_26207);
nand U29406 (N_29406,N_25836,N_26755);
and U29407 (N_29407,N_25934,N_24181);
nand U29408 (N_29408,N_24938,N_26420);
or U29409 (N_29409,N_25612,N_24344);
xor U29410 (N_29410,N_24968,N_24822);
xnor U29411 (N_29411,N_26969,N_24664);
xnor U29412 (N_29412,N_25849,N_26059);
nor U29413 (N_29413,N_26817,N_25442);
xor U29414 (N_29414,N_25000,N_25242);
and U29415 (N_29415,N_25205,N_24719);
nor U29416 (N_29416,N_25013,N_25340);
nand U29417 (N_29417,N_26581,N_26611);
and U29418 (N_29418,N_24998,N_25164);
nor U29419 (N_29419,N_25060,N_25665);
and U29420 (N_29420,N_25805,N_24726);
or U29421 (N_29421,N_26784,N_26366);
nand U29422 (N_29422,N_25535,N_24066);
nand U29423 (N_29423,N_25706,N_25844);
or U29424 (N_29424,N_26357,N_24844);
xor U29425 (N_29425,N_24487,N_26265);
nand U29426 (N_29426,N_26717,N_26496);
and U29427 (N_29427,N_26364,N_24956);
nor U29428 (N_29428,N_24814,N_25112);
nand U29429 (N_29429,N_24519,N_24594);
nor U29430 (N_29430,N_26307,N_26972);
xor U29431 (N_29431,N_26052,N_24957);
xor U29432 (N_29432,N_25009,N_25108);
xnor U29433 (N_29433,N_25733,N_25703);
xor U29434 (N_29434,N_24163,N_26266);
xor U29435 (N_29435,N_26048,N_24979);
xor U29436 (N_29436,N_24817,N_26047);
or U29437 (N_29437,N_25782,N_24253);
nor U29438 (N_29438,N_24121,N_24013);
or U29439 (N_29439,N_26200,N_26011);
or U29440 (N_29440,N_24615,N_24335);
or U29441 (N_29441,N_25837,N_24431);
xnor U29442 (N_29442,N_25512,N_26596);
and U29443 (N_29443,N_24484,N_25044);
xor U29444 (N_29444,N_25577,N_24161);
nand U29445 (N_29445,N_25913,N_26342);
nand U29446 (N_29446,N_24934,N_25521);
nand U29447 (N_29447,N_26580,N_24625);
nand U29448 (N_29448,N_25209,N_25645);
or U29449 (N_29449,N_25180,N_26435);
nand U29450 (N_29450,N_26526,N_26760);
or U29451 (N_29451,N_25357,N_24428);
nor U29452 (N_29452,N_25003,N_24124);
or U29453 (N_29453,N_26025,N_25076);
or U29454 (N_29454,N_24520,N_24082);
nand U29455 (N_29455,N_24058,N_24374);
nand U29456 (N_29456,N_26883,N_26386);
xor U29457 (N_29457,N_26655,N_24831);
or U29458 (N_29458,N_26416,N_25595);
xor U29459 (N_29459,N_24110,N_24958);
xor U29460 (N_29460,N_26183,N_24033);
or U29461 (N_29461,N_25164,N_26303);
nor U29462 (N_29462,N_24334,N_24804);
nor U29463 (N_29463,N_25911,N_26830);
xnor U29464 (N_29464,N_25981,N_26216);
nor U29465 (N_29465,N_24882,N_24186);
nand U29466 (N_29466,N_26482,N_25623);
nand U29467 (N_29467,N_24401,N_24067);
or U29468 (N_29468,N_24681,N_25098);
or U29469 (N_29469,N_24800,N_26157);
xnor U29470 (N_29470,N_24397,N_24064);
nor U29471 (N_29471,N_26272,N_26491);
and U29472 (N_29472,N_26356,N_26502);
nand U29473 (N_29473,N_25258,N_24826);
and U29474 (N_29474,N_24248,N_26979);
or U29475 (N_29475,N_26117,N_24370);
nor U29476 (N_29476,N_24098,N_26745);
and U29477 (N_29477,N_26698,N_24116);
or U29478 (N_29478,N_25430,N_24959);
and U29479 (N_29479,N_26926,N_25466);
xor U29480 (N_29480,N_24993,N_24868);
or U29481 (N_29481,N_25590,N_24188);
xnor U29482 (N_29482,N_26724,N_25519);
xnor U29483 (N_29483,N_25626,N_26054);
xnor U29484 (N_29484,N_26089,N_26953);
xor U29485 (N_29485,N_24524,N_25083);
nor U29486 (N_29486,N_25478,N_25323);
nor U29487 (N_29487,N_24160,N_26052);
and U29488 (N_29488,N_26526,N_25994);
and U29489 (N_29489,N_25153,N_25355);
or U29490 (N_29490,N_25775,N_24558);
or U29491 (N_29491,N_25106,N_25059);
and U29492 (N_29492,N_26091,N_25354);
and U29493 (N_29493,N_25071,N_26569);
nand U29494 (N_29494,N_26881,N_24912);
and U29495 (N_29495,N_24836,N_26368);
nor U29496 (N_29496,N_24297,N_24808);
nand U29497 (N_29497,N_26626,N_26089);
xnor U29498 (N_29498,N_24528,N_24070);
xnor U29499 (N_29499,N_25867,N_26662);
nand U29500 (N_29500,N_26512,N_25462);
or U29501 (N_29501,N_24684,N_26940);
nor U29502 (N_29502,N_25333,N_25258);
and U29503 (N_29503,N_24319,N_25840);
or U29504 (N_29504,N_26012,N_25159);
and U29505 (N_29505,N_25920,N_25175);
or U29506 (N_29506,N_25225,N_26747);
nand U29507 (N_29507,N_24077,N_25511);
xor U29508 (N_29508,N_24745,N_24441);
or U29509 (N_29509,N_25889,N_24948);
and U29510 (N_29510,N_25864,N_26567);
nand U29511 (N_29511,N_24305,N_24718);
and U29512 (N_29512,N_26137,N_24326);
nand U29513 (N_29513,N_24591,N_24304);
xnor U29514 (N_29514,N_25146,N_26321);
or U29515 (N_29515,N_25544,N_26429);
and U29516 (N_29516,N_24712,N_26306);
and U29517 (N_29517,N_26105,N_25080);
nand U29518 (N_29518,N_24600,N_25976);
xor U29519 (N_29519,N_26966,N_24540);
or U29520 (N_29520,N_24362,N_24285);
nand U29521 (N_29521,N_26452,N_25438);
xor U29522 (N_29522,N_24302,N_26976);
and U29523 (N_29523,N_25659,N_25665);
or U29524 (N_29524,N_26521,N_24966);
or U29525 (N_29525,N_24539,N_26776);
and U29526 (N_29526,N_26117,N_25151);
nand U29527 (N_29527,N_24726,N_24453);
and U29528 (N_29528,N_26950,N_24655);
nand U29529 (N_29529,N_25222,N_24481);
xnor U29530 (N_29530,N_24668,N_25555);
nor U29531 (N_29531,N_26824,N_26834);
or U29532 (N_29532,N_26259,N_25688);
nand U29533 (N_29533,N_26221,N_26779);
nor U29534 (N_29534,N_24896,N_24330);
nand U29535 (N_29535,N_25923,N_26579);
or U29536 (N_29536,N_26818,N_26971);
and U29537 (N_29537,N_26047,N_24809);
and U29538 (N_29538,N_24428,N_24968);
or U29539 (N_29539,N_26210,N_25358);
and U29540 (N_29540,N_26234,N_24803);
nor U29541 (N_29541,N_25100,N_24029);
or U29542 (N_29542,N_26606,N_25947);
xnor U29543 (N_29543,N_25697,N_25199);
nor U29544 (N_29544,N_25697,N_25479);
and U29545 (N_29545,N_24271,N_24584);
and U29546 (N_29546,N_26354,N_24767);
xor U29547 (N_29547,N_25642,N_25335);
or U29548 (N_29548,N_25459,N_25587);
or U29549 (N_29549,N_26308,N_25213);
or U29550 (N_29550,N_26201,N_24797);
nor U29551 (N_29551,N_25436,N_26310);
nor U29552 (N_29552,N_25375,N_25684);
nand U29553 (N_29553,N_25473,N_26847);
nor U29554 (N_29554,N_24706,N_26843);
and U29555 (N_29555,N_26325,N_25681);
xor U29556 (N_29556,N_26326,N_24944);
and U29557 (N_29557,N_24173,N_25019);
nand U29558 (N_29558,N_24588,N_26617);
xor U29559 (N_29559,N_24168,N_24550);
and U29560 (N_29560,N_25573,N_24169);
and U29561 (N_29561,N_24857,N_24196);
nand U29562 (N_29562,N_25642,N_25757);
and U29563 (N_29563,N_25953,N_25520);
and U29564 (N_29564,N_26522,N_26532);
xnor U29565 (N_29565,N_26232,N_24788);
or U29566 (N_29566,N_26341,N_25066);
nor U29567 (N_29567,N_26789,N_24726);
nor U29568 (N_29568,N_26492,N_25325);
and U29569 (N_29569,N_25210,N_24797);
and U29570 (N_29570,N_26028,N_24802);
xor U29571 (N_29571,N_25631,N_24829);
nand U29572 (N_29572,N_25917,N_24807);
nor U29573 (N_29573,N_24810,N_24146);
nor U29574 (N_29574,N_24410,N_26793);
xor U29575 (N_29575,N_26135,N_24530);
or U29576 (N_29576,N_26320,N_25932);
and U29577 (N_29577,N_24302,N_25862);
nand U29578 (N_29578,N_24822,N_26232);
xor U29579 (N_29579,N_24257,N_26350);
nand U29580 (N_29580,N_24035,N_26832);
and U29581 (N_29581,N_26447,N_26788);
nor U29582 (N_29582,N_25120,N_24678);
or U29583 (N_29583,N_25810,N_25948);
nand U29584 (N_29584,N_26629,N_26189);
xnor U29585 (N_29585,N_24385,N_26490);
xor U29586 (N_29586,N_24970,N_24912);
xor U29587 (N_29587,N_25630,N_24315);
nand U29588 (N_29588,N_26778,N_26918);
and U29589 (N_29589,N_26491,N_26428);
or U29590 (N_29590,N_25135,N_25309);
and U29591 (N_29591,N_25428,N_26686);
nand U29592 (N_29592,N_24199,N_26600);
and U29593 (N_29593,N_25744,N_25298);
xnor U29594 (N_29594,N_25481,N_24740);
xnor U29595 (N_29595,N_26746,N_25174);
xor U29596 (N_29596,N_26601,N_25779);
xor U29597 (N_29597,N_24831,N_25280);
or U29598 (N_29598,N_25432,N_26843);
nand U29599 (N_29599,N_25582,N_24480);
and U29600 (N_29600,N_26895,N_25302);
or U29601 (N_29601,N_26426,N_25974);
and U29602 (N_29602,N_25567,N_24153);
or U29603 (N_29603,N_25882,N_26582);
nor U29604 (N_29604,N_26670,N_24278);
nand U29605 (N_29605,N_25218,N_26521);
and U29606 (N_29606,N_24304,N_24037);
or U29607 (N_29607,N_25217,N_26146);
and U29608 (N_29608,N_26678,N_25212);
xnor U29609 (N_29609,N_24295,N_24608);
xor U29610 (N_29610,N_25424,N_26178);
or U29611 (N_29611,N_24382,N_24921);
xnor U29612 (N_29612,N_26886,N_25673);
nor U29613 (N_29613,N_24776,N_26113);
nand U29614 (N_29614,N_24086,N_26831);
or U29615 (N_29615,N_25439,N_25293);
and U29616 (N_29616,N_25579,N_26680);
or U29617 (N_29617,N_25325,N_26676);
and U29618 (N_29618,N_26617,N_25646);
xnor U29619 (N_29619,N_26416,N_24107);
xor U29620 (N_29620,N_25622,N_24696);
nand U29621 (N_29621,N_25563,N_25934);
or U29622 (N_29622,N_24993,N_26790);
nor U29623 (N_29623,N_25175,N_24972);
xnor U29624 (N_29624,N_24950,N_24238);
and U29625 (N_29625,N_25311,N_26267);
nand U29626 (N_29626,N_26482,N_26411);
or U29627 (N_29627,N_24126,N_24047);
and U29628 (N_29628,N_25948,N_25789);
and U29629 (N_29629,N_24977,N_26576);
nor U29630 (N_29630,N_24788,N_25972);
nor U29631 (N_29631,N_26893,N_25690);
or U29632 (N_29632,N_25562,N_26071);
nor U29633 (N_29633,N_26773,N_24775);
nand U29634 (N_29634,N_26627,N_25488);
nand U29635 (N_29635,N_26584,N_25048);
xnor U29636 (N_29636,N_26086,N_24555);
nor U29637 (N_29637,N_26108,N_25895);
nor U29638 (N_29638,N_26055,N_26197);
nand U29639 (N_29639,N_25036,N_24092);
nor U29640 (N_29640,N_26139,N_26264);
nand U29641 (N_29641,N_24034,N_25892);
nor U29642 (N_29642,N_26140,N_24282);
nand U29643 (N_29643,N_26158,N_25069);
nor U29644 (N_29644,N_25220,N_24783);
or U29645 (N_29645,N_26647,N_26363);
nand U29646 (N_29646,N_25668,N_26552);
and U29647 (N_29647,N_26091,N_25997);
nor U29648 (N_29648,N_24741,N_24444);
or U29649 (N_29649,N_26875,N_26836);
or U29650 (N_29650,N_26759,N_25765);
nor U29651 (N_29651,N_25271,N_24752);
nor U29652 (N_29652,N_25826,N_24674);
nand U29653 (N_29653,N_25341,N_25866);
nor U29654 (N_29654,N_26999,N_25288);
or U29655 (N_29655,N_24650,N_25052);
nand U29656 (N_29656,N_26675,N_26744);
or U29657 (N_29657,N_26723,N_25435);
nor U29658 (N_29658,N_25387,N_26853);
or U29659 (N_29659,N_26294,N_24504);
nor U29660 (N_29660,N_25417,N_24129);
nand U29661 (N_29661,N_26813,N_24836);
and U29662 (N_29662,N_24435,N_24563);
xor U29663 (N_29663,N_24201,N_25025);
nand U29664 (N_29664,N_24545,N_26303);
or U29665 (N_29665,N_25988,N_26782);
or U29666 (N_29666,N_25126,N_26107);
and U29667 (N_29667,N_26075,N_24213);
nand U29668 (N_29668,N_26141,N_26017);
nor U29669 (N_29669,N_24519,N_25583);
nor U29670 (N_29670,N_25848,N_25433);
or U29671 (N_29671,N_26355,N_26172);
nand U29672 (N_29672,N_24980,N_24728);
xor U29673 (N_29673,N_24434,N_26188);
nor U29674 (N_29674,N_26035,N_25174);
nand U29675 (N_29675,N_24450,N_25911);
xnor U29676 (N_29676,N_24354,N_26644);
and U29677 (N_29677,N_25505,N_26713);
nand U29678 (N_29678,N_25777,N_26441);
or U29679 (N_29679,N_24750,N_25824);
xor U29680 (N_29680,N_25682,N_24859);
nand U29681 (N_29681,N_25680,N_25894);
nand U29682 (N_29682,N_26213,N_25202);
and U29683 (N_29683,N_25756,N_26968);
nand U29684 (N_29684,N_26891,N_24801);
or U29685 (N_29685,N_25648,N_24969);
and U29686 (N_29686,N_25396,N_24244);
nor U29687 (N_29687,N_26484,N_26075);
nand U29688 (N_29688,N_26551,N_25249);
nand U29689 (N_29689,N_25031,N_24803);
nand U29690 (N_29690,N_26327,N_25972);
and U29691 (N_29691,N_26522,N_25074);
nor U29692 (N_29692,N_26625,N_24437);
or U29693 (N_29693,N_24019,N_26387);
and U29694 (N_29694,N_24900,N_26876);
xnor U29695 (N_29695,N_26694,N_26460);
nor U29696 (N_29696,N_25580,N_24840);
or U29697 (N_29697,N_25986,N_26994);
nor U29698 (N_29698,N_26715,N_24242);
and U29699 (N_29699,N_24338,N_26098);
nand U29700 (N_29700,N_25427,N_25388);
nand U29701 (N_29701,N_26379,N_25819);
nand U29702 (N_29702,N_25497,N_26269);
nand U29703 (N_29703,N_26324,N_25009);
xor U29704 (N_29704,N_25841,N_24159);
xor U29705 (N_29705,N_26704,N_24417);
and U29706 (N_29706,N_25834,N_24946);
nor U29707 (N_29707,N_26601,N_24528);
xnor U29708 (N_29708,N_24307,N_26829);
nand U29709 (N_29709,N_26870,N_26957);
and U29710 (N_29710,N_26168,N_24925);
xor U29711 (N_29711,N_25836,N_24270);
and U29712 (N_29712,N_25102,N_24833);
nor U29713 (N_29713,N_24275,N_24801);
and U29714 (N_29714,N_26437,N_26000);
or U29715 (N_29715,N_24563,N_25942);
and U29716 (N_29716,N_25580,N_25828);
xnor U29717 (N_29717,N_25979,N_24790);
nand U29718 (N_29718,N_25095,N_26736);
and U29719 (N_29719,N_25989,N_24909);
and U29720 (N_29720,N_24302,N_25615);
or U29721 (N_29721,N_24707,N_26436);
nand U29722 (N_29722,N_24156,N_26031);
and U29723 (N_29723,N_26650,N_25097);
nor U29724 (N_29724,N_24351,N_24396);
xnor U29725 (N_29725,N_26122,N_26280);
xnor U29726 (N_29726,N_25233,N_26853);
and U29727 (N_29727,N_26712,N_24390);
xor U29728 (N_29728,N_25272,N_25339);
and U29729 (N_29729,N_24834,N_24711);
xnor U29730 (N_29730,N_25341,N_24262);
xor U29731 (N_29731,N_25118,N_25432);
nor U29732 (N_29732,N_24170,N_24442);
nand U29733 (N_29733,N_25381,N_26836);
xor U29734 (N_29734,N_25138,N_26810);
nor U29735 (N_29735,N_26929,N_26398);
nand U29736 (N_29736,N_24289,N_26245);
and U29737 (N_29737,N_26126,N_26659);
xnor U29738 (N_29738,N_24616,N_26616);
or U29739 (N_29739,N_26179,N_24791);
and U29740 (N_29740,N_24913,N_26710);
nand U29741 (N_29741,N_24154,N_25138);
nor U29742 (N_29742,N_24511,N_24345);
and U29743 (N_29743,N_25174,N_26428);
nor U29744 (N_29744,N_26086,N_24897);
and U29745 (N_29745,N_26287,N_25297);
nand U29746 (N_29746,N_25896,N_26018);
and U29747 (N_29747,N_24070,N_26151);
and U29748 (N_29748,N_25729,N_26740);
or U29749 (N_29749,N_26267,N_26225);
or U29750 (N_29750,N_24141,N_25596);
nand U29751 (N_29751,N_24054,N_25779);
nor U29752 (N_29752,N_25353,N_24496);
and U29753 (N_29753,N_26260,N_24683);
and U29754 (N_29754,N_26810,N_25254);
nor U29755 (N_29755,N_26974,N_24946);
nand U29756 (N_29756,N_25820,N_26613);
and U29757 (N_29757,N_26147,N_24656);
xor U29758 (N_29758,N_24454,N_24571);
and U29759 (N_29759,N_25664,N_24622);
or U29760 (N_29760,N_26602,N_26522);
or U29761 (N_29761,N_26286,N_26626);
nand U29762 (N_29762,N_26837,N_25651);
nand U29763 (N_29763,N_24686,N_25068);
nor U29764 (N_29764,N_25707,N_26018);
and U29765 (N_29765,N_26355,N_26401);
nand U29766 (N_29766,N_25546,N_26210);
nor U29767 (N_29767,N_25005,N_25702);
nor U29768 (N_29768,N_26090,N_25161);
and U29769 (N_29769,N_25391,N_26078);
and U29770 (N_29770,N_24844,N_25449);
nor U29771 (N_29771,N_25990,N_26903);
nor U29772 (N_29772,N_26501,N_26129);
nand U29773 (N_29773,N_26585,N_26304);
and U29774 (N_29774,N_24607,N_26602);
and U29775 (N_29775,N_26762,N_25163);
and U29776 (N_29776,N_24933,N_24495);
nor U29777 (N_29777,N_24249,N_25877);
or U29778 (N_29778,N_24390,N_24860);
or U29779 (N_29779,N_24037,N_26498);
and U29780 (N_29780,N_24552,N_26904);
nand U29781 (N_29781,N_26876,N_24281);
nand U29782 (N_29782,N_26899,N_24256);
and U29783 (N_29783,N_24874,N_26129);
and U29784 (N_29784,N_24316,N_26979);
xor U29785 (N_29785,N_26677,N_26240);
xnor U29786 (N_29786,N_25568,N_26292);
or U29787 (N_29787,N_24595,N_24049);
and U29788 (N_29788,N_25891,N_24683);
nor U29789 (N_29789,N_24044,N_24161);
or U29790 (N_29790,N_24041,N_25378);
and U29791 (N_29791,N_24254,N_26987);
xor U29792 (N_29792,N_26044,N_26423);
xor U29793 (N_29793,N_26329,N_24328);
nand U29794 (N_29794,N_24869,N_26388);
or U29795 (N_29795,N_26002,N_24987);
nand U29796 (N_29796,N_24092,N_25548);
nor U29797 (N_29797,N_24638,N_26335);
xor U29798 (N_29798,N_26915,N_26373);
nand U29799 (N_29799,N_26291,N_25100);
or U29800 (N_29800,N_26285,N_25594);
and U29801 (N_29801,N_25205,N_26316);
or U29802 (N_29802,N_26304,N_26401);
and U29803 (N_29803,N_24608,N_26152);
nand U29804 (N_29804,N_24953,N_26664);
and U29805 (N_29805,N_25342,N_25240);
and U29806 (N_29806,N_25985,N_25154);
xnor U29807 (N_29807,N_25355,N_24967);
or U29808 (N_29808,N_24548,N_26993);
nor U29809 (N_29809,N_24743,N_26397);
or U29810 (N_29810,N_24136,N_24671);
nand U29811 (N_29811,N_26970,N_24931);
nand U29812 (N_29812,N_25542,N_25088);
or U29813 (N_29813,N_25827,N_24511);
nand U29814 (N_29814,N_25102,N_26772);
xor U29815 (N_29815,N_26179,N_26754);
nor U29816 (N_29816,N_24812,N_24744);
or U29817 (N_29817,N_24940,N_24701);
and U29818 (N_29818,N_25626,N_26012);
nand U29819 (N_29819,N_24501,N_25476);
or U29820 (N_29820,N_24988,N_25563);
nand U29821 (N_29821,N_24088,N_26974);
xnor U29822 (N_29822,N_25384,N_24973);
and U29823 (N_29823,N_26074,N_26520);
or U29824 (N_29824,N_24728,N_26060);
xor U29825 (N_29825,N_25996,N_24761);
nand U29826 (N_29826,N_26191,N_24777);
and U29827 (N_29827,N_24196,N_25313);
nor U29828 (N_29828,N_26065,N_26434);
and U29829 (N_29829,N_26007,N_25995);
and U29830 (N_29830,N_25928,N_25898);
and U29831 (N_29831,N_26503,N_24470);
or U29832 (N_29832,N_24610,N_25749);
xnor U29833 (N_29833,N_25078,N_24223);
xor U29834 (N_29834,N_26534,N_25475);
xnor U29835 (N_29835,N_24625,N_24318);
or U29836 (N_29836,N_24227,N_25540);
and U29837 (N_29837,N_26374,N_26713);
nor U29838 (N_29838,N_26958,N_26547);
nor U29839 (N_29839,N_26241,N_26732);
nand U29840 (N_29840,N_26773,N_24700);
nor U29841 (N_29841,N_24284,N_26523);
and U29842 (N_29842,N_26042,N_26137);
nand U29843 (N_29843,N_26549,N_25992);
xor U29844 (N_29844,N_25861,N_26790);
or U29845 (N_29845,N_25020,N_26792);
or U29846 (N_29846,N_24787,N_25252);
xnor U29847 (N_29847,N_24187,N_24290);
nor U29848 (N_29848,N_25889,N_25012);
nand U29849 (N_29849,N_24566,N_25912);
and U29850 (N_29850,N_26511,N_26717);
and U29851 (N_29851,N_24772,N_24873);
and U29852 (N_29852,N_25120,N_24744);
nand U29853 (N_29853,N_25693,N_25889);
nor U29854 (N_29854,N_25736,N_24328);
or U29855 (N_29855,N_25008,N_25537);
and U29856 (N_29856,N_25120,N_25279);
xor U29857 (N_29857,N_25129,N_26747);
xor U29858 (N_29858,N_26917,N_26674);
and U29859 (N_29859,N_26070,N_25983);
and U29860 (N_29860,N_24949,N_26961);
or U29861 (N_29861,N_24155,N_25092);
nor U29862 (N_29862,N_24364,N_26324);
nor U29863 (N_29863,N_26834,N_25250);
nor U29864 (N_29864,N_26051,N_26210);
xor U29865 (N_29865,N_26024,N_24299);
xor U29866 (N_29866,N_26335,N_24852);
nand U29867 (N_29867,N_25371,N_24543);
nand U29868 (N_29868,N_24964,N_25008);
nand U29869 (N_29869,N_26792,N_25814);
nor U29870 (N_29870,N_25740,N_25627);
or U29871 (N_29871,N_24202,N_25618);
nand U29872 (N_29872,N_26994,N_26305);
or U29873 (N_29873,N_24544,N_25102);
nand U29874 (N_29874,N_25109,N_26019);
nand U29875 (N_29875,N_25548,N_26312);
or U29876 (N_29876,N_24181,N_24324);
or U29877 (N_29877,N_25859,N_26491);
nor U29878 (N_29878,N_24424,N_25023);
or U29879 (N_29879,N_26543,N_25724);
xnor U29880 (N_29880,N_24137,N_25391);
or U29881 (N_29881,N_26713,N_26751);
xnor U29882 (N_29882,N_24644,N_26789);
xor U29883 (N_29883,N_26394,N_25302);
xnor U29884 (N_29884,N_24155,N_25130);
nor U29885 (N_29885,N_25888,N_24792);
xnor U29886 (N_29886,N_26125,N_25343);
and U29887 (N_29887,N_25563,N_26440);
or U29888 (N_29888,N_24683,N_25064);
nand U29889 (N_29889,N_26033,N_26194);
and U29890 (N_29890,N_25600,N_24350);
nor U29891 (N_29891,N_26634,N_25232);
and U29892 (N_29892,N_24680,N_26061);
and U29893 (N_29893,N_25730,N_24059);
nand U29894 (N_29894,N_25643,N_24468);
nand U29895 (N_29895,N_25624,N_24625);
or U29896 (N_29896,N_24736,N_25554);
xor U29897 (N_29897,N_26119,N_26738);
nand U29898 (N_29898,N_25925,N_25421);
and U29899 (N_29899,N_25022,N_25377);
xnor U29900 (N_29900,N_24914,N_26686);
nor U29901 (N_29901,N_25426,N_25423);
nor U29902 (N_29902,N_24703,N_25738);
nor U29903 (N_29903,N_24047,N_24964);
nand U29904 (N_29904,N_26289,N_26091);
xnor U29905 (N_29905,N_25038,N_24850);
or U29906 (N_29906,N_26811,N_25252);
nor U29907 (N_29907,N_24772,N_24666);
xor U29908 (N_29908,N_25948,N_25527);
xor U29909 (N_29909,N_25215,N_24483);
nor U29910 (N_29910,N_24324,N_25124);
xor U29911 (N_29911,N_25358,N_24397);
and U29912 (N_29912,N_24011,N_25146);
nand U29913 (N_29913,N_26528,N_24308);
nor U29914 (N_29914,N_24561,N_25027);
and U29915 (N_29915,N_26025,N_25758);
and U29916 (N_29916,N_24637,N_26309);
nand U29917 (N_29917,N_24698,N_25343);
nor U29918 (N_29918,N_25795,N_24952);
or U29919 (N_29919,N_25298,N_24231);
nor U29920 (N_29920,N_24650,N_26730);
or U29921 (N_29921,N_24404,N_25350);
and U29922 (N_29922,N_26740,N_24867);
or U29923 (N_29923,N_24320,N_25807);
and U29924 (N_29924,N_24326,N_26806);
nand U29925 (N_29925,N_26042,N_25105);
and U29926 (N_29926,N_25262,N_26286);
and U29927 (N_29927,N_25803,N_24187);
or U29928 (N_29928,N_25760,N_26595);
nor U29929 (N_29929,N_25225,N_26257);
nand U29930 (N_29930,N_25788,N_24688);
and U29931 (N_29931,N_24047,N_26571);
nand U29932 (N_29932,N_24896,N_26890);
and U29933 (N_29933,N_25546,N_26712);
xnor U29934 (N_29934,N_25010,N_24210);
or U29935 (N_29935,N_25088,N_24392);
and U29936 (N_29936,N_26704,N_26727);
nor U29937 (N_29937,N_26275,N_25995);
nand U29938 (N_29938,N_24923,N_26199);
xnor U29939 (N_29939,N_26863,N_26490);
and U29940 (N_29940,N_26598,N_25060);
nand U29941 (N_29941,N_26665,N_24550);
nor U29942 (N_29942,N_26100,N_24633);
nor U29943 (N_29943,N_26705,N_26237);
or U29944 (N_29944,N_24114,N_25892);
nand U29945 (N_29945,N_24842,N_26861);
or U29946 (N_29946,N_25757,N_25960);
or U29947 (N_29947,N_24665,N_24102);
and U29948 (N_29948,N_26872,N_26932);
nor U29949 (N_29949,N_24307,N_24406);
nand U29950 (N_29950,N_24641,N_24775);
xnor U29951 (N_29951,N_24133,N_26982);
xnor U29952 (N_29952,N_25562,N_24351);
nor U29953 (N_29953,N_25391,N_24074);
nand U29954 (N_29954,N_25240,N_26238);
or U29955 (N_29955,N_24589,N_26259);
nand U29956 (N_29956,N_26537,N_25029);
xor U29957 (N_29957,N_26376,N_24288);
and U29958 (N_29958,N_26245,N_26925);
nand U29959 (N_29959,N_24166,N_26473);
xnor U29960 (N_29960,N_24468,N_25581);
nor U29961 (N_29961,N_24754,N_26347);
nor U29962 (N_29962,N_24297,N_24775);
xor U29963 (N_29963,N_26038,N_25385);
nand U29964 (N_29964,N_24101,N_24033);
and U29965 (N_29965,N_26856,N_26566);
xnor U29966 (N_29966,N_24413,N_26680);
and U29967 (N_29967,N_26417,N_26875);
nor U29968 (N_29968,N_25892,N_24970);
nand U29969 (N_29969,N_24030,N_26732);
or U29970 (N_29970,N_25813,N_26030);
and U29971 (N_29971,N_24709,N_24410);
nand U29972 (N_29972,N_26720,N_26070);
or U29973 (N_29973,N_26025,N_24047);
nand U29974 (N_29974,N_26654,N_24428);
or U29975 (N_29975,N_24735,N_25533);
nor U29976 (N_29976,N_26152,N_25135);
xor U29977 (N_29977,N_26740,N_24838);
nand U29978 (N_29978,N_24076,N_24463);
and U29979 (N_29979,N_25364,N_25865);
xnor U29980 (N_29980,N_26201,N_24925);
nand U29981 (N_29981,N_26331,N_24194);
nor U29982 (N_29982,N_24138,N_26773);
xor U29983 (N_29983,N_25397,N_24911);
or U29984 (N_29984,N_26774,N_25436);
nand U29985 (N_29985,N_25745,N_26373);
and U29986 (N_29986,N_25458,N_26900);
or U29987 (N_29987,N_24470,N_26773);
nand U29988 (N_29988,N_25866,N_25218);
xnor U29989 (N_29989,N_25723,N_25716);
or U29990 (N_29990,N_26318,N_25292);
nor U29991 (N_29991,N_25040,N_24350);
nor U29992 (N_29992,N_25946,N_25441);
nor U29993 (N_29993,N_26768,N_24294);
and U29994 (N_29994,N_26623,N_26890);
and U29995 (N_29995,N_24984,N_25725);
and U29996 (N_29996,N_26201,N_25623);
xnor U29997 (N_29997,N_26107,N_26702);
xnor U29998 (N_29998,N_24126,N_26613);
xor U29999 (N_29999,N_25914,N_24802);
xor UO_0 (O_0,N_29179,N_29656);
and UO_1 (O_1,N_28412,N_27011);
or UO_2 (O_2,N_29251,N_27458);
and UO_3 (O_3,N_27617,N_27057);
nand UO_4 (O_4,N_28280,N_29643);
and UO_5 (O_5,N_29159,N_27392);
nand UO_6 (O_6,N_29239,N_27743);
or UO_7 (O_7,N_27729,N_27940);
xor UO_8 (O_8,N_27097,N_27911);
nand UO_9 (O_9,N_29531,N_27843);
xnor UO_10 (O_10,N_28388,N_27518);
nand UO_11 (O_11,N_28530,N_29313);
or UO_12 (O_12,N_29190,N_29861);
or UO_13 (O_13,N_27820,N_27908);
or UO_14 (O_14,N_27204,N_28724);
and UO_15 (O_15,N_28274,N_27888);
or UO_16 (O_16,N_29495,N_29778);
and UO_17 (O_17,N_29538,N_29007);
nor UO_18 (O_18,N_27497,N_29259);
nor UO_19 (O_19,N_28376,N_27174);
or UO_20 (O_20,N_29205,N_28720);
nor UO_21 (O_21,N_29961,N_29636);
or UO_22 (O_22,N_29601,N_27399);
and UO_23 (O_23,N_29930,N_28362);
or UO_24 (O_24,N_29958,N_29960);
and UO_25 (O_25,N_28754,N_29068);
and UO_26 (O_26,N_27469,N_27074);
and UO_27 (O_27,N_27736,N_28746);
nand UO_28 (O_28,N_29837,N_28888);
nand UO_29 (O_29,N_28606,N_28011);
nor UO_30 (O_30,N_28884,N_27781);
nand UO_31 (O_31,N_29921,N_27079);
and UO_32 (O_32,N_27784,N_27506);
and UO_33 (O_33,N_27724,N_28428);
nor UO_34 (O_34,N_29234,N_27535);
nand UO_35 (O_35,N_27633,N_28215);
nand UO_36 (O_36,N_28069,N_29868);
or UO_37 (O_37,N_27866,N_29722);
or UO_38 (O_38,N_28802,N_27301);
or UO_39 (O_39,N_27587,N_29945);
nor UO_40 (O_40,N_28400,N_27500);
or UO_41 (O_41,N_28704,N_28080);
nand UO_42 (O_42,N_29955,N_27612);
nand UO_43 (O_43,N_28217,N_28903);
nand UO_44 (O_44,N_28482,N_27734);
xor UO_45 (O_45,N_29415,N_27412);
nand UO_46 (O_46,N_28022,N_29064);
nor UO_47 (O_47,N_27995,N_27693);
or UO_48 (O_48,N_28378,N_27658);
xor UO_49 (O_49,N_29646,N_29265);
and UO_50 (O_50,N_28355,N_29249);
nand UO_51 (O_51,N_29248,N_28869);
nor UO_52 (O_52,N_27765,N_29588);
nand UO_53 (O_53,N_27006,N_28491);
nand UO_54 (O_54,N_27672,N_27698);
nand UO_55 (O_55,N_27049,N_29836);
and UO_56 (O_56,N_27905,N_28387);
nor UO_57 (O_57,N_28978,N_27267);
or UO_58 (O_58,N_27524,N_27433);
nand UO_59 (O_59,N_29390,N_28375);
xnor UO_60 (O_60,N_27046,N_27952);
and UO_61 (O_61,N_29027,N_27692);
and UO_62 (O_62,N_27434,N_27815);
or UO_63 (O_63,N_28590,N_29221);
xor UO_64 (O_64,N_29031,N_29474);
xor UO_65 (O_65,N_27769,N_28909);
nor UO_66 (O_66,N_27117,N_28706);
nor UO_67 (O_67,N_29139,N_28543);
xor UO_68 (O_68,N_29499,N_28092);
nand UO_69 (O_69,N_27884,N_29908);
nand UO_70 (O_70,N_29148,N_29286);
xnor UO_71 (O_71,N_29619,N_28921);
and UO_72 (O_72,N_28453,N_27146);
or UO_73 (O_73,N_28858,N_27984);
or UO_74 (O_74,N_28402,N_28140);
and UO_75 (O_75,N_29212,N_28605);
nor UO_76 (O_76,N_28851,N_28913);
nand UO_77 (O_77,N_29553,N_29336);
xor UO_78 (O_78,N_28301,N_27833);
nand UO_79 (O_79,N_27033,N_27013);
nor UO_80 (O_80,N_27741,N_27935);
nand UO_81 (O_81,N_28928,N_29931);
nor UO_82 (O_82,N_28121,N_27848);
or UO_83 (O_83,N_29845,N_27192);
nor UO_84 (O_84,N_29215,N_28054);
nor UO_85 (O_85,N_27598,N_27607);
or UO_86 (O_86,N_27716,N_27746);
nand UO_87 (O_87,N_29476,N_28283);
nand UO_88 (O_88,N_28573,N_29462);
and UO_89 (O_89,N_28962,N_28498);
and UO_90 (O_90,N_28193,N_28075);
nor UO_91 (O_91,N_29006,N_28827);
or UO_92 (O_92,N_27590,N_27705);
and UO_93 (O_93,N_28617,N_29564);
and UO_94 (O_94,N_29719,N_28915);
xnor UO_95 (O_95,N_27648,N_29302);
xnor UO_96 (O_96,N_29400,N_28423);
nor UO_97 (O_97,N_27227,N_28919);
nor UO_98 (O_98,N_29078,N_28105);
and UO_99 (O_99,N_28684,N_27160);
nand UO_100 (O_100,N_29356,N_28566);
nand UO_101 (O_101,N_27066,N_28821);
xnor UO_102 (O_102,N_27676,N_27346);
or UO_103 (O_103,N_27774,N_29144);
xnor UO_104 (O_104,N_28448,N_27120);
nand UO_105 (O_105,N_27557,N_29555);
or UO_106 (O_106,N_29918,N_27675);
nor UO_107 (O_107,N_29678,N_28697);
or UO_108 (O_108,N_28023,N_28649);
or UO_109 (O_109,N_29453,N_29922);
or UO_110 (O_110,N_27463,N_29291);
xnor UO_111 (O_111,N_28271,N_28451);
and UO_112 (O_112,N_29098,N_29261);
nand UO_113 (O_113,N_28956,N_28894);
and UO_114 (O_114,N_29459,N_29393);
nand UO_115 (O_115,N_27112,N_28158);
nor UO_116 (O_116,N_29335,N_28088);
or UO_117 (O_117,N_27320,N_29762);
nor UO_118 (O_118,N_27667,N_27094);
and UO_119 (O_119,N_27449,N_29645);
xor UO_120 (O_120,N_28325,N_27345);
and UO_121 (O_121,N_27404,N_27730);
and UO_122 (O_122,N_29652,N_28805);
xor UO_123 (O_123,N_29408,N_27153);
and UO_124 (O_124,N_28296,N_29074);
and UO_125 (O_125,N_28418,N_27534);
xnor UO_126 (O_126,N_29230,N_27946);
nand UO_127 (O_127,N_28184,N_27542);
nor UO_128 (O_128,N_27517,N_27789);
nor UO_129 (O_129,N_29477,N_28346);
and UO_130 (O_130,N_27187,N_27055);
nand UO_131 (O_131,N_27181,N_28582);
nor UO_132 (O_132,N_27466,N_28990);
xnor UO_133 (O_133,N_29649,N_28523);
nand UO_134 (O_134,N_28776,N_28863);
or UO_135 (O_135,N_27699,N_27180);
or UO_136 (O_136,N_28644,N_28469);
or UO_137 (O_137,N_29515,N_29565);
or UO_138 (O_138,N_29297,N_27154);
or UO_139 (O_139,N_29520,N_27727);
nand UO_140 (O_140,N_29013,N_27488);
nand UO_141 (O_141,N_29511,N_28791);
and UO_142 (O_142,N_28598,N_29222);
or UO_143 (O_143,N_27374,N_28016);
or UO_144 (O_144,N_29432,N_29754);
or UO_145 (O_145,N_28855,N_29153);
and UO_146 (O_146,N_29079,N_29829);
nand UO_147 (O_147,N_29414,N_27673);
and UO_148 (O_148,N_29238,N_29445);
or UO_149 (O_149,N_27615,N_28799);
or UO_150 (O_150,N_29391,N_29717);
and UO_151 (O_151,N_27137,N_29653);
nand UO_152 (O_152,N_29568,N_27683);
and UO_153 (O_153,N_27514,N_28258);
xnor UO_154 (O_154,N_27552,N_27415);
nor UO_155 (O_155,N_28098,N_28436);
or UO_156 (O_156,N_27168,N_28584);
and UO_157 (O_157,N_27318,N_29549);
nor UO_158 (O_158,N_28082,N_27568);
or UO_159 (O_159,N_28291,N_29493);
nor UO_160 (O_160,N_27785,N_28624);
nand UO_161 (O_161,N_28675,N_27974);
nand UO_162 (O_162,N_29523,N_29723);
or UO_163 (O_163,N_28793,N_27442);
nor UO_164 (O_164,N_28638,N_29536);
and UO_165 (O_165,N_29244,N_29933);
nand UO_166 (O_166,N_28429,N_27677);
and UO_167 (O_167,N_27430,N_28288);
and UO_168 (O_168,N_29864,N_27255);
or UO_169 (O_169,N_29949,N_28896);
and UO_170 (O_170,N_27232,N_27242);
or UO_171 (O_171,N_28439,N_27519);
and UO_172 (O_172,N_29800,N_28930);
and UO_173 (O_173,N_29529,N_28440);
nor UO_174 (O_174,N_28289,N_29644);
nor UO_175 (O_175,N_28957,N_28923);
nand UO_176 (O_176,N_28232,N_28323);
nor UO_177 (O_177,N_27619,N_29578);
nor UO_178 (O_178,N_28731,N_28848);
or UO_179 (O_179,N_29688,N_27830);
xor UO_180 (O_180,N_28281,N_29434);
xnor UO_181 (O_181,N_29566,N_28090);
xnor UO_182 (O_182,N_27476,N_28838);
nand UO_183 (O_183,N_28500,N_28238);
nor UO_184 (O_184,N_27982,N_29990);
xnor UO_185 (O_185,N_27377,N_27173);
xor UO_186 (O_186,N_27681,N_27801);
nand UO_187 (O_187,N_29420,N_29301);
nand UO_188 (O_188,N_27080,N_29269);
nand UO_189 (O_189,N_29347,N_28991);
nand UO_190 (O_190,N_27357,N_27694);
xor UO_191 (O_191,N_27048,N_27106);
nor UO_192 (O_192,N_28172,N_28654);
and UO_193 (O_193,N_29739,N_29494);
nand UO_194 (O_194,N_29062,N_27445);
nand UO_195 (O_195,N_28862,N_29607);
nand UO_196 (O_196,N_29785,N_28256);
xor UO_197 (O_197,N_27788,N_28342);
nor UO_198 (O_198,N_28305,N_28782);
and UO_199 (O_199,N_27498,N_28028);
nand UO_200 (O_200,N_27897,N_27157);
xnor UO_201 (O_201,N_27269,N_29976);
and UO_202 (O_202,N_27319,N_28550);
or UO_203 (O_203,N_28349,N_29740);
xnor UO_204 (O_204,N_28309,N_28872);
nand UO_205 (O_205,N_29797,N_28327);
and UO_206 (O_206,N_27281,N_29579);
xor UO_207 (O_207,N_29895,N_29295);
nor UO_208 (O_208,N_29699,N_28564);
and UO_209 (O_209,N_28488,N_27014);
and UO_210 (O_210,N_28842,N_29614);
or UO_211 (O_211,N_27611,N_29326);
nor UO_212 (O_212,N_29987,N_28828);
xor UO_213 (O_213,N_29630,N_29506);
and UO_214 (O_214,N_28815,N_28065);
nor UO_215 (O_215,N_27031,N_28020);
or UO_216 (O_216,N_28614,N_29072);
or UO_217 (O_217,N_28417,N_29428);
xnor UO_218 (O_218,N_27898,N_27855);
xnor UO_219 (O_219,N_29809,N_28314);
or UO_220 (O_220,N_29032,N_29663);
and UO_221 (O_221,N_27042,N_27240);
and UO_222 (O_222,N_27359,N_27712);
or UO_223 (O_223,N_27203,N_28463);
or UO_224 (O_224,N_29368,N_27058);
and UO_225 (O_225,N_28895,N_29551);
nor UO_226 (O_226,N_29721,N_27997);
nor UO_227 (O_227,N_27100,N_28977);
nor UO_228 (O_228,N_29469,N_29528);
xor UO_229 (O_229,N_29189,N_29272);
nand UO_230 (O_230,N_29448,N_29070);
nor UO_231 (O_231,N_29957,N_29254);
nand UO_232 (O_232,N_28655,N_28181);
or UO_233 (O_233,N_28634,N_29804);
nand UO_234 (O_234,N_29177,N_28611);
nor UO_235 (O_235,N_29917,N_29631);
and UO_236 (O_236,N_28150,N_27142);
xnor UO_237 (O_237,N_29787,N_28292);
xor UO_238 (O_238,N_28535,N_27367);
or UO_239 (O_239,N_28473,N_29805);
or UO_240 (O_240,N_27287,N_27628);
and UO_241 (O_241,N_27777,N_29436);
xor UO_242 (O_242,N_27914,N_29132);
xor UO_243 (O_243,N_28047,N_29855);
nand UO_244 (O_244,N_27300,N_29142);
nor UO_245 (O_245,N_29701,N_27207);
or UO_246 (O_246,N_28653,N_29262);
nor UO_247 (O_247,N_27069,N_29143);
xnor UO_248 (O_248,N_29540,N_27728);
and UO_249 (O_249,N_28240,N_28180);
and UO_250 (O_250,N_27902,N_29417);
nor UO_251 (O_251,N_29424,N_28540);
and UO_252 (O_252,N_27128,N_29231);
or UO_253 (O_253,N_28825,N_29478);
and UO_254 (O_254,N_29939,N_27719);
nand UO_255 (O_255,N_27516,N_28242);
xor UO_256 (O_256,N_29083,N_28286);
xor UO_257 (O_257,N_27523,N_29289);
or UO_258 (O_258,N_29831,N_27877);
nor UO_259 (O_259,N_28361,N_28339);
xor UO_260 (O_260,N_27448,N_28067);
xor UO_261 (O_261,N_29396,N_29869);
and UO_262 (O_262,N_29751,N_27717);
and UO_263 (O_263,N_28148,N_29123);
xnor UO_264 (O_264,N_28911,N_28259);
or UO_265 (O_265,N_27505,N_28003);
or UO_266 (O_266,N_27233,N_28156);
nand UO_267 (O_267,N_29314,N_28413);
nand UO_268 (O_268,N_27022,N_29042);
nand UO_269 (O_269,N_29294,N_29541);
nor UO_270 (O_270,N_28886,N_28421);
nor UO_271 (O_271,N_29734,N_28639);
or UO_272 (O_272,N_28132,N_29217);
or UO_273 (O_273,N_27018,N_29902);
and UO_274 (O_274,N_27572,N_27299);
and UO_275 (O_275,N_29983,N_29874);
and UO_276 (O_276,N_27403,N_29461);
and UO_277 (O_277,N_29627,N_27937);
and UO_278 (O_278,N_29321,N_27229);
xor UO_279 (O_279,N_29967,N_29219);
nand UO_280 (O_280,N_28447,N_27322);
nor UO_281 (O_281,N_27393,N_27674);
or UO_282 (O_282,N_27970,N_29211);
or UO_283 (O_283,N_28685,N_27001);
xor UO_284 (O_284,N_27875,N_28068);
and UO_285 (O_285,N_29300,N_27155);
nand UO_286 (O_286,N_27793,N_28489);
or UO_287 (O_287,N_27446,N_29546);
xor UO_288 (O_288,N_28513,N_28719);
nor UO_289 (O_289,N_27533,N_29532);
and UO_290 (O_290,N_28477,N_27917);
or UO_291 (O_291,N_29613,N_28700);
nand UO_292 (O_292,N_28954,N_28931);
nand UO_293 (O_293,N_29076,N_28580);
or UO_294 (O_294,N_28622,N_28998);
nand UO_295 (O_295,N_27973,N_28632);
and UO_296 (O_296,N_28087,N_29073);
nor UO_297 (O_297,N_28307,N_27496);
or UO_298 (O_298,N_29772,N_29946);
nand UO_299 (O_299,N_29709,N_27162);
and UO_300 (O_300,N_29556,N_27803);
xnor UO_301 (O_301,N_27444,N_27679);
nor UO_302 (O_302,N_29882,N_27807);
and UO_303 (O_303,N_27259,N_27314);
and UO_304 (O_304,N_29371,N_27230);
nand UO_305 (O_305,N_28845,N_28608);
xor UO_306 (O_306,N_29992,N_28265);
nand UO_307 (O_307,N_28427,N_27870);
or UO_308 (O_308,N_29747,N_28204);
and UO_309 (O_309,N_27328,N_29150);
nor UO_310 (O_310,N_27825,N_27596);
or UO_311 (O_311,N_29165,N_28974);
xor UO_312 (O_312,N_27994,N_27208);
nor UO_313 (O_313,N_28446,N_29322);
nand UO_314 (O_314,N_27682,N_28357);
and UO_315 (O_315,N_29599,N_27686);
nor UO_316 (O_316,N_29102,N_29329);
and UO_317 (O_317,N_28982,N_27526);
nand UO_318 (O_318,N_28328,N_27355);
or UO_319 (O_319,N_27718,N_29250);
or UO_320 (O_320,N_27333,N_27759);
and UO_321 (O_321,N_27313,N_27749);
nor UO_322 (O_322,N_29484,N_29849);
and UO_323 (O_323,N_28248,N_28391);
or UO_324 (O_324,N_27130,N_28358);
xor UO_325 (O_325,N_28424,N_28175);
xnor UO_326 (O_326,N_29667,N_28381);
nor UO_327 (O_327,N_27249,N_28006);
nor UO_328 (O_328,N_29163,N_27198);
nor UO_329 (O_329,N_28330,N_29071);
nand UO_330 (O_330,N_27456,N_28501);
nand UO_331 (O_331,N_28433,N_29750);
xor UO_332 (O_332,N_27571,N_27271);
xor UO_333 (O_333,N_29256,N_27577);
xnor UO_334 (O_334,N_27244,N_27060);
or UO_335 (O_335,N_29317,N_29047);
nand UO_336 (O_336,N_29969,N_29736);
or UO_337 (O_337,N_29374,N_28662);
or UO_338 (O_338,N_28899,N_29664);
nand UO_339 (O_339,N_29051,N_29848);
or UO_340 (O_340,N_27297,N_29035);
nor UO_341 (O_341,N_29896,N_27510);
nor UO_342 (O_342,N_27356,N_27655);
or UO_343 (O_343,N_27817,N_29905);
xor UO_344 (O_344,N_28251,N_27169);
nor UO_345 (O_345,N_28640,N_28134);
or UO_346 (O_346,N_29629,N_27512);
or UO_347 (O_347,N_28942,N_28876);
and UO_348 (O_348,N_28127,N_27113);
nand UO_349 (O_349,N_29524,N_28359);
and UO_350 (O_350,N_28396,N_27307);
nor UO_351 (O_351,N_27580,N_27981);
xnor UO_352 (O_352,N_28004,N_28567);
and UO_353 (O_353,N_29067,N_28732);
or UO_354 (O_354,N_29765,N_29623);
or UO_355 (O_355,N_28290,N_29640);
nand UO_356 (O_356,N_28519,N_29381);
and UO_357 (O_357,N_28694,N_27707);
nor UO_358 (O_358,N_27840,N_29048);
and UO_359 (O_359,N_27382,N_28091);
xor UO_360 (O_360,N_29367,N_27179);
nand UO_361 (O_361,N_27538,N_27625);
or UO_362 (O_362,N_29973,N_28889);
nand UO_363 (O_363,N_29331,N_28315);
and UO_364 (O_364,N_29991,N_28390);
and UO_365 (O_365,N_29161,N_27141);
or UO_366 (O_366,N_29503,N_29028);
and UO_367 (O_367,N_28239,N_27814);
xnor UO_368 (O_368,N_29609,N_28494);
or UO_369 (O_369,N_29573,N_28951);
or UO_370 (O_370,N_28514,N_29686);
xnor UO_371 (O_371,N_27105,N_28021);
nor UO_372 (O_372,N_28182,N_28460);
and UO_373 (O_373,N_27899,N_28379);
xor UO_374 (O_374,N_27447,N_27738);
nand UO_375 (O_375,N_27939,N_27284);
or UO_376 (O_376,N_28744,N_28596);
and UO_377 (O_377,N_27652,N_29433);
or UO_378 (O_378,N_29698,N_27723);
nor UO_379 (O_379,N_27929,N_28595);
nand UO_380 (O_380,N_28508,N_28343);
or UO_381 (O_381,N_29220,N_29943);
or UO_382 (O_382,N_28667,N_29009);
nand UO_383 (O_383,N_29604,N_29953);
and UO_384 (O_384,N_29792,N_27603);
nand UO_385 (O_385,N_28437,N_28225);
nand UO_386 (O_386,N_27083,N_28681);
nor UO_387 (O_387,N_27629,N_28351);
nand UO_388 (O_388,N_29611,N_29866);
and UO_389 (O_389,N_27821,N_27161);
or UO_390 (O_390,N_27104,N_27035);
xnor UO_391 (O_391,N_29543,N_28260);
nand UO_392 (O_392,N_27753,N_27184);
or UO_393 (O_393,N_29235,N_29004);
xor UO_394 (O_394,N_28057,N_29888);
nand UO_395 (O_395,N_29731,N_27706);
and UO_396 (O_396,N_27000,N_27760);
or UO_397 (O_397,N_28633,N_29544);
or UO_398 (O_398,N_28814,N_28136);
nor UO_399 (O_399,N_28118,N_28701);
and UO_400 (O_400,N_28282,N_28865);
nand UO_401 (O_401,N_29403,N_29187);
nand UO_402 (O_402,N_29635,N_28490);
xnor UO_403 (O_403,N_28813,N_28364);
xor UO_404 (O_404,N_27165,N_29971);
xor UO_405 (O_405,N_28972,N_29878);
nor UO_406 (O_406,N_27487,N_27582);
xor UO_407 (O_407,N_27964,N_28244);
and UO_408 (O_408,N_29483,N_29054);
nor UO_409 (O_409,N_27998,N_27129);
nand UO_410 (O_410,N_27258,N_28620);
or UO_411 (O_411,N_28918,N_28946);
xnor UO_412 (O_412,N_28032,N_27387);
nand UO_413 (O_413,N_27934,N_28431);
or UO_414 (O_414,N_28665,N_27023);
or UO_415 (O_415,N_28920,N_28784);
and UO_416 (O_416,N_29581,N_28496);
xnor UO_417 (O_417,N_29121,N_28013);
xor UO_418 (O_418,N_28602,N_29775);
xor UO_419 (O_419,N_27747,N_27930);
xnor UO_420 (O_420,N_28306,N_27660);
xor UO_421 (O_421,N_29392,N_28541);
or UO_422 (O_422,N_28616,N_29385);
xnor UO_423 (O_423,N_29275,N_28571);
and UO_424 (O_424,N_28973,N_27077);
nor UO_425 (O_425,N_27780,N_29174);
or UO_426 (O_426,N_29811,N_29303);
or UO_427 (O_427,N_28228,N_27455);
nor UO_428 (O_428,N_27334,N_29312);
nor UO_429 (O_429,N_28304,N_27918);
xor UO_430 (O_430,N_27581,N_27892);
nor UO_431 (O_431,N_29351,N_27098);
xnor UO_432 (O_432,N_27796,N_27967);
nand UO_433 (O_433,N_27391,N_27171);
and UO_434 (O_434,N_28707,N_28109);
nand UO_435 (O_435,N_29464,N_28333);
xor UO_436 (O_436,N_27122,N_27241);
xor UO_437 (O_437,N_29372,N_29061);
and UO_438 (O_438,N_29038,N_29936);
nor UO_439 (O_439,N_27321,N_29449);
xor UO_440 (O_440,N_29398,N_29674);
nand UO_441 (O_441,N_28046,N_28370);
nand UO_442 (O_442,N_29180,N_28853);
nand UO_443 (O_443,N_27896,N_28669);
nor UO_444 (O_444,N_28812,N_28777);
nor UO_445 (O_445,N_27933,N_29340);
or UO_446 (O_446,N_28659,N_29853);
xnor UO_447 (O_447,N_27178,N_27782);
and UO_448 (O_448,N_28741,N_27744);
xor UO_449 (O_449,N_28334,N_28760);
nor UO_450 (O_450,N_27024,N_27566);
or UO_451 (O_451,N_27402,N_28416);
xor UO_452 (O_452,N_28775,N_29842);
nor UO_453 (O_453,N_28867,N_27624);
or UO_454 (O_454,N_28161,N_29875);
nor UO_455 (O_455,N_28808,N_29082);
or UO_456 (O_456,N_29164,N_29271);
xor UO_457 (O_457,N_27344,N_28648);
or UO_458 (O_458,N_29624,N_28045);
nand UO_459 (O_459,N_27850,N_28495);
xor UO_460 (O_460,N_28176,N_29703);
or UO_461 (O_461,N_27324,N_27539);
or UO_462 (O_462,N_29608,N_27613);
nand UO_463 (O_463,N_29802,N_29606);
nor UO_464 (O_464,N_27969,N_29407);
nor UO_465 (O_465,N_29692,N_27653);
and UO_466 (O_466,N_29847,N_27992);
or UO_467 (O_467,N_28717,N_29018);
nand UO_468 (O_468,N_29610,N_29569);
nand UO_469 (O_469,N_29716,N_29117);
and UO_470 (O_470,N_28594,N_28578);
nor UO_471 (O_471,N_27621,N_27697);
nor UO_472 (O_472,N_28729,N_27254);
xnor UO_473 (O_473,N_29060,N_28967);
nor UO_474 (O_474,N_28832,N_29362);
or UO_475 (O_475,N_29111,N_27150);
xnor UO_476 (O_476,N_28167,N_27152);
and UO_477 (O_477,N_28205,N_28179);
or UO_478 (O_478,N_27501,N_27051);
or UO_479 (O_479,N_27966,N_29937);
nor UO_480 (O_480,N_28017,N_28154);
or UO_481 (O_481,N_29560,N_29416);
nor UO_482 (O_482,N_27108,N_27725);
or UO_483 (O_483,N_29363,N_29146);
nor UO_484 (O_484,N_27750,N_28506);
nand UO_485 (O_485,N_29252,N_27604);
or UO_486 (O_486,N_27405,N_29388);
or UO_487 (O_487,N_28189,N_28103);
and UO_488 (O_488,N_27177,N_27742);
xor UO_489 (O_489,N_29602,N_28104);
and UO_490 (O_490,N_27589,N_29545);
and UO_491 (O_491,N_28859,N_27980);
and UO_492 (O_492,N_28243,N_28615);
nor UO_493 (O_493,N_27925,N_27585);
xor UO_494 (O_494,N_28432,N_27560);
and UO_495 (O_495,N_29258,N_29769);
xnor UO_496 (O_496,N_28916,N_28397);
or UO_497 (O_497,N_28861,N_27191);
nor UO_498 (O_498,N_27823,N_28561);
nand UO_499 (O_499,N_27547,N_28925);
and UO_500 (O_500,N_28849,N_29753);
nand UO_501 (O_501,N_29181,N_29049);
nor UO_502 (O_502,N_27722,N_28976);
and UO_503 (O_503,N_29683,N_29263);
and UO_504 (O_504,N_27339,N_27839);
xnor UO_505 (O_505,N_29577,N_27068);
xnor UO_506 (O_506,N_27038,N_28941);
nand UO_507 (O_507,N_28806,N_29087);
or UO_508 (O_508,N_28471,N_29223);
xnor UO_509 (O_509,N_28094,N_29170);
nand UO_510 (O_510,N_27954,N_27745);
nor UO_511 (O_511,N_28478,N_27428);
and UO_512 (O_512,N_29395,N_28001);
or UO_513 (O_513,N_29225,N_28171);
xnor UO_514 (O_514,N_29757,N_27927);
or UO_515 (O_515,N_27895,N_29830);
nor UO_516 (O_516,N_28143,N_28630);
and UO_517 (O_517,N_28768,N_28079);
nand UO_518 (O_518,N_28173,N_28618);
and UO_519 (O_519,N_27390,N_29594);
nand UO_520 (O_520,N_29486,N_27236);
and UO_521 (O_521,N_28353,N_27827);
xor UO_522 (O_522,N_29745,N_27030);
and UO_523 (O_523,N_27443,N_27503);
nand UO_524 (O_524,N_29152,N_28019);
xnor UO_525 (O_525,N_27138,N_28117);
or UO_526 (O_526,N_27665,N_29518);
and UO_527 (O_527,N_28263,N_28367);
or UO_528 (O_528,N_29708,N_27989);
xor UO_529 (O_529,N_29912,N_29015);
nand UO_530 (O_530,N_27687,N_27869);
nor UO_531 (O_531,N_28880,N_28545);
xnor UO_532 (O_532,N_28209,N_27306);
nor UO_533 (O_533,N_29412,N_29232);
or UO_534 (O_534,N_27265,N_27824);
or UO_535 (O_535,N_29526,N_28671);
and UO_536 (O_536,N_28317,N_28038);
nand UO_537 (O_537,N_27620,N_29517);
xnor UO_538 (O_538,N_29525,N_29213);
xor UO_539 (O_539,N_28264,N_29788);
and UO_540 (O_540,N_28613,N_29923);
and UO_541 (O_541,N_29097,N_29670);
nand UO_542 (O_542,N_29793,N_27252);
and UO_543 (O_543,N_28874,N_29352);
and UO_544 (O_544,N_28932,N_29030);
nand UO_545 (O_545,N_29380,N_28690);
or UO_546 (O_546,N_28955,N_27007);
xnor UO_547 (O_547,N_29425,N_29767);
nand UO_548 (O_548,N_29046,N_28177);
and UO_549 (O_549,N_29979,N_28186);
or UO_550 (O_550,N_27912,N_27485);
and UO_551 (O_551,N_28987,N_28986);
or UO_552 (O_552,N_28981,N_29729);
or UO_553 (O_553,N_27757,N_28005);
xor UO_554 (O_554,N_27894,N_29404);
nor UO_555 (O_555,N_28338,N_27545);
and UO_556 (O_556,N_27493,N_29088);
nand UO_557 (O_557,N_29178,N_28619);
and UO_558 (O_558,N_27555,N_28831);
xor UO_559 (O_559,N_28686,N_27668);
nor UO_560 (O_560,N_28610,N_27436);
nand UO_561 (O_561,N_28503,N_28472);
nand UO_562 (O_562,N_27091,N_28668);
and UO_563 (O_563,N_29561,N_29050);
nor UO_564 (O_564,N_27431,N_28547);
nor UO_565 (O_565,N_28350,N_29475);
nand UO_566 (O_566,N_29344,N_29125);
nand UO_567 (O_567,N_28324,N_29118);
or UO_568 (O_568,N_27862,N_28823);
nor UO_569 (O_569,N_29101,N_28159);
and UO_570 (O_570,N_28174,N_29266);
xor UO_571 (O_571,N_28787,N_29509);
xnor UO_572 (O_572,N_27295,N_29737);
or UO_573 (O_573,N_28230,N_29514);
or UO_574 (O_574,N_29676,N_28692);
or UO_575 (O_575,N_29268,N_29828);
xnor UO_576 (O_576,N_27114,N_28036);
and UO_577 (O_577,N_29867,N_29122);
xor UO_578 (O_578,N_29548,N_27845);
xor UO_579 (O_579,N_28072,N_29846);
and UO_580 (O_580,N_27158,N_27957);
and UO_581 (O_581,N_27972,N_29537);
or UO_582 (O_582,N_27635,N_29278);
xnor UO_583 (O_583,N_27372,N_28442);
nor UO_584 (O_584,N_27770,N_28377);
or UO_585 (O_585,N_27502,N_28052);
nor UO_586 (O_586,N_27525,N_28927);
nor UO_587 (O_587,N_28457,N_27642);
nand UO_588 (O_588,N_27323,N_28406);
xnor UO_589 (O_589,N_28102,N_29012);
nand UO_590 (O_590,N_29157,N_27189);
nand UO_591 (O_591,N_29468,N_29816);
nor UO_592 (O_592,N_28940,N_28246);
and UO_593 (O_593,N_28245,N_29777);
xor UO_594 (O_594,N_27308,N_29240);
nand UO_595 (O_595,N_28185,N_28847);
xor UO_596 (O_596,N_27958,N_28456);
nand UO_597 (O_597,N_28002,N_27132);
xor UO_598 (O_598,N_27816,N_27977);
or UO_599 (O_599,N_27605,N_29338);
nand UO_600 (O_600,N_29901,N_27085);
and UO_601 (O_601,N_27872,N_28476);
nand UO_602 (O_602,N_29827,N_27071);
xor UO_603 (O_603,N_27231,N_27421);
nand UO_604 (O_604,N_27025,N_29657);
and UO_605 (O_605,N_28601,N_27423);
or UO_606 (O_606,N_28629,N_29799);
and UO_607 (O_607,N_27579,N_27923);
and UO_608 (O_608,N_28018,N_28835);
or UO_609 (O_609,N_28319,N_29784);
nand UO_610 (O_610,N_28818,N_28664);
nand UO_611 (O_611,N_29724,N_28949);
nand UO_612 (O_612,N_28947,N_29521);
nand UO_613 (O_613,N_27826,N_27838);
nor UO_614 (O_614,N_27294,N_29648);
nor UO_615 (O_615,N_29204,N_29039);
nand UO_616 (O_616,N_29637,N_29916);
nor UO_617 (O_617,N_27397,N_27928);
nand UO_618 (O_618,N_28549,N_28426);
xor UO_619 (O_619,N_27167,N_28645);
nand UO_620 (O_620,N_28910,N_29859);
or UO_621 (O_621,N_29790,N_29197);
nor UO_622 (O_622,N_28833,N_28860);
and UO_623 (O_623,N_28577,N_28781);
nand UO_624 (O_624,N_28537,N_28557);
nand UO_625 (O_625,N_27127,N_27887);
and UO_626 (O_626,N_28252,N_28468);
xor UO_627 (O_627,N_29685,N_28666);
or UO_628 (O_628,N_29660,N_28214);
nor UO_629 (O_629,N_29357,N_29172);
or UO_630 (O_630,N_28623,N_28516);
and UO_631 (O_631,N_28202,N_28129);
and UO_632 (O_632,N_27479,N_29200);
xor UO_633 (O_633,N_29010,N_28738);
or UO_634 (O_634,N_27987,N_28199);
nand UO_635 (O_635,N_28555,N_27197);
nor UO_636 (O_636,N_27309,N_27832);
or UO_637 (O_637,N_29768,N_28348);
and UO_638 (O_638,N_28336,N_29423);
and UO_639 (O_639,N_28830,N_27133);
xor UO_640 (O_640,N_29033,N_29654);
or UO_641 (O_641,N_29003,N_28191);
nor UO_642 (O_642,N_29169,N_29993);
xor UO_643 (O_643,N_27864,N_27695);
nand UO_644 (O_644,N_27956,N_27330);
and UO_645 (O_645,N_27076,N_27664);
nor UO_646 (O_646,N_27016,N_27429);
nand UO_647 (O_647,N_27851,N_29280);
xor UO_648 (O_648,N_29669,N_27504);
nand UO_649 (O_649,N_28677,N_29890);
nand UO_650 (O_650,N_29409,N_27944);
xnor UO_651 (O_651,N_27861,N_29690);
and UO_652 (O_652,N_27225,N_28438);
or UO_653 (O_653,N_27809,N_29377);
or UO_654 (O_654,N_28755,N_28445);
xor UO_655 (O_655,N_28807,N_29974);
and UO_656 (O_656,N_29639,N_29584);
xnor UO_657 (O_657,N_29008,N_28120);
xor UO_658 (O_658,N_27491,N_29612);
nor UO_659 (O_659,N_27550,N_28201);
nor UO_660 (O_660,N_27139,N_28492);
and UO_661 (O_661,N_29539,N_28646);
or UO_662 (O_662,N_27867,N_27690);
nand UO_663 (O_663,N_29191,N_27623);
and UO_664 (O_664,N_29596,N_28532);
and UO_665 (O_665,N_28108,N_28026);
nor UO_666 (O_666,N_28740,N_28316);
or UO_667 (O_667,N_29066,N_29292);
nor UO_668 (O_668,N_29998,N_29485);
and UO_669 (O_669,N_27291,N_29628);
xor UO_670 (O_670,N_27732,N_27818);
nor UO_671 (O_671,N_28769,N_28546);
nand UO_672 (O_672,N_27947,N_29091);
or UO_673 (O_673,N_28834,N_28365);
nor UO_674 (O_674,N_27420,N_27708);
nand UO_675 (O_675,N_27544,N_29095);
nor UO_676 (O_676,N_27103,N_28394);
or UO_677 (O_677,N_28914,N_29794);
and UO_678 (O_678,N_29934,N_29634);
nand UO_679 (O_679,N_28055,N_29705);
or UO_680 (O_680,N_27711,N_27806);
and UO_681 (O_681,N_29752,N_28678);
nand UO_682 (O_682,N_27900,N_27546);
xor UO_683 (O_683,N_28059,N_27052);
nand UO_684 (O_684,N_28892,N_29376);
xor UO_685 (O_685,N_28563,N_29950);
nor UO_686 (O_686,N_27841,N_28035);
nor UO_687 (O_687,N_27779,N_28255);
and UO_688 (O_688,N_29386,N_28691);
xnor UO_689 (O_689,N_29910,N_29706);
nand UO_690 (O_690,N_27288,N_29870);
nor UO_691 (O_691,N_29002,N_27311);
nor UO_692 (O_692,N_27661,N_29668);
xor UO_693 (O_693,N_28133,N_27156);
or UO_694 (O_694,N_28213,N_28454);
xor UO_695 (O_695,N_28086,N_28081);
nand UO_696 (O_696,N_27962,N_29576);
nand UO_697 (O_697,N_29501,N_28037);
and UO_698 (O_698,N_27941,N_27685);
or UO_699 (O_699,N_29452,N_28221);
and UO_700 (O_700,N_28409,N_27410);
or UO_701 (O_701,N_27593,N_27578);
xnor UO_702 (O_702,N_28278,N_28757);
xnor UO_703 (O_703,N_28992,N_29430);
nand UO_704 (O_704,N_28352,N_29903);
xor UO_705 (O_705,N_29481,N_27145);
or UO_706 (O_706,N_28761,N_28558);
xnor UO_707 (O_707,N_27651,N_29997);
and UO_708 (O_708,N_29605,N_29497);
and UO_709 (O_709,N_27805,N_29129);
nor UO_710 (O_710,N_28313,N_28077);
nand UO_711 (O_711,N_29839,N_28285);
or UO_712 (O_712,N_28642,N_29763);
nor UO_713 (O_713,N_28229,N_27657);
nand UO_714 (O_714,N_27121,N_28562);
xor UO_715 (O_715,N_27226,N_28907);
xnor UO_716 (O_716,N_27985,N_29463);
and UO_717 (O_717,N_27406,N_28560);
and UO_718 (O_718,N_29715,N_27880);
nor UO_719 (O_719,N_27243,N_29382);
xor UO_720 (O_720,N_28637,N_27509);
and UO_721 (O_721,N_27045,N_27247);
and UO_722 (O_722,N_29887,N_28950);
and UO_723 (O_723,N_29176,N_29137);
and UO_724 (O_724,N_27282,N_27285);
nor UO_725 (O_725,N_27758,N_29052);
nand UO_726 (O_726,N_29037,N_28997);
nor UO_727 (O_727,N_28208,N_29858);
and UO_728 (O_728,N_28093,N_29673);
xnor UO_729 (O_729,N_27131,N_27715);
nor UO_730 (O_730,N_28881,N_28603);
nand UO_731 (O_731,N_29704,N_27527);
and UO_732 (O_732,N_27111,N_29782);
nand UO_733 (O_733,N_29622,N_28841);
or UO_734 (O_734,N_27264,N_27595);
nand UO_735 (O_735,N_28771,N_29410);
or UO_736 (O_736,N_28486,N_29632);
xnor UO_737 (O_737,N_29041,N_27860);
nand UO_738 (O_738,N_29977,N_28795);
nand UO_739 (O_739,N_29766,N_27248);
nor UO_740 (O_740,N_28162,N_27351);
xor UO_741 (O_741,N_29516,N_28948);
nand UO_742 (O_742,N_27124,N_29311);
or UO_743 (O_743,N_28458,N_27647);
or UO_744 (O_744,N_28099,N_29527);
nor UO_745 (O_745,N_27089,N_28206);
xnor UO_746 (O_746,N_29963,N_29496);
or UO_747 (O_747,N_28125,N_28042);
or UO_748 (O_748,N_29185,N_29865);
nor UO_749 (O_749,N_29952,N_27521);
and UO_750 (O_750,N_28009,N_29439);
nand UO_751 (O_751,N_29909,N_27065);
nand UO_752 (O_752,N_28247,N_29746);
or UO_753 (O_753,N_29671,N_27388);
or UO_754 (O_754,N_28960,N_29077);
nand UO_755 (O_755,N_28063,N_29810);
and UO_756 (O_756,N_28058,N_29354);
or UO_757 (O_757,N_27812,N_28890);
and UO_758 (O_758,N_29755,N_28879);
nand UO_759 (O_759,N_29642,N_27795);
xnor UO_760 (O_760,N_28368,N_28674);
and UO_761 (O_761,N_29591,N_27804);
or UO_762 (O_762,N_28898,N_27986);
nand UO_763 (O_763,N_29358,N_29133);
nand UO_764 (O_764,N_27609,N_29615);
nand UO_765 (O_765,N_29519,N_29298);
and UO_766 (O_766,N_27650,N_28583);
and UO_767 (O_767,N_29808,N_27163);
nor UO_768 (O_768,N_29020,N_28111);
or UO_769 (O_769,N_28465,N_28138);
xor UO_770 (O_770,N_27714,N_29884);
or UO_771 (O_771,N_29720,N_27853);
xnor UO_772 (O_772,N_29898,N_27889);
nor UO_773 (O_773,N_27426,N_27764);
or UO_774 (O_774,N_29105,N_29821);
nor UO_775 (O_775,N_29399,N_28538);
nand UO_776 (O_776,N_29552,N_29926);
nor UO_777 (O_777,N_28483,N_27125);
nand UO_778 (O_778,N_27553,N_28656);
and UO_779 (O_779,N_27384,N_27400);
or UO_780 (O_780,N_28170,N_27961);
xnor UO_781 (O_781,N_29589,N_28906);
or UO_782 (O_782,N_29488,N_27289);
and UO_783 (O_783,N_28718,N_27411);
and UO_784 (O_784,N_28178,N_28525);
nor UO_785 (O_785,N_28322,N_27432);
nor UO_786 (O_786,N_29780,N_27453);
xor UO_787 (O_787,N_29360,N_27999);
or UO_788 (O_788,N_29019,N_27822);
nand UO_789 (O_789,N_29089,N_28123);
nand UO_790 (O_790,N_27136,N_28399);
nand UO_791 (O_791,N_27159,N_29996);
nand UO_792 (O_792,N_29277,N_28548);
or UO_793 (O_793,N_29981,N_28078);
and UO_794 (O_794,N_27800,N_27050);
nand UO_795 (O_795,N_28236,N_29188);
or UO_796 (O_796,N_27976,N_29951);
xnor UO_797 (O_797,N_27205,N_29938);
nand UO_798 (O_798,N_27062,N_27486);
xor UO_799 (O_799,N_27365,N_29687);
nor UO_800 (O_800,N_28912,N_28369);
and UO_801 (O_801,N_29840,N_27965);
xor UO_802 (O_802,N_29201,N_28066);
xnor UO_803 (O_803,N_27883,N_29247);
xnor UO_804 (O_804,N_28166,N_28303);
or UO_805 (O_805,N_29460,N_28984);
and UO_806 (O_806,N_28794,N_28857);
xor UO_807 (O_807,N_28484,N_29110);
nand UO_808 (O_808,N_27148,N_27015);
nor UO_809 (O_809,N_28124,N_27858);
nand UO_810 (O_810,N_28822,N_29279);
and UO_811 (O_811,N_27088,N_27831);
xnor UO_812 (O_812,N_28559,N_28188);
and UO_813 (O_813,N_27235,N_28676);
nand UO_814 (O_814,N_27327,N_28395);
nor UO_815 (O_815,N_28575,N_27451);
nand UO_816 (O_816,N_27854,N_28536);
or UO_817 (O_817,N_27634,N_27082);
nand UO_818 (O_818,N_29978,N_29679);
nor UO_819 (O_819,N_28050,N_28461);
xnor UO_820 (O_820,N_27915,N_28015);
and UO_821 (O_821,N_28621,N_27275);
nand UO_822 (O_822,N_29440,N_27070);
nor UO_823 (O_823,N_29965,N_28266);
and UO_824 (O_824,N_28836,N_29756);
nand UO_825 (O_825,N_28689,N_29894);
nor UO_826 (O_826,N_27748,N_27201);
xnor UO_827 (O_827,N_27008,N_29025);
nand UO_828 (O_828,N_29284,N_28147);
or UO_829 (O_829,N_29838,N_28734);
nor UO_830 (O_830,N_27360,N_29554);
nor UO_831 (O_831,N_29237,N_27960);
or UO_832 (O_832,N_29534,N_29216);
or UO_833 (O_833,N_29092,N_27959);
nand UO_834 (O_834,N_28145,N_27280);
nor UO_835 (O_835,N_28027,N_28040);
nor UO_836 (O_836,N_29138,N_29455);
xnor UO_837 (O_837,N_29168,N_28041);
nor UO_838 (O_838,N_28965,N_27370);
xnor UO_839 (O_839,N_29173,N_27010);
and UO_840 (O_840,N_29287,N_27040);
or UO_841 (O_841,N_27268,N_28031);
nand UO_842 (O_842,N_28415,N_29288);
and UO_843 (O_843,N_27041,N_29491);
nand UO_844 (O_844,N_27188,N_27101);
xnor UO_845 (O_845,N_29798,N_29999);
nor UO_846 (O_846,N_28101,N_27090);
or UO_847 (O_847,N_27700,N_28939);
and UO_848 (O_848,N_29959,N_28728);
or UO_849 (O_849,N_28820,N_28122);
nor UO_850 (O_850,N_27353,N_28137);
nand UO_851 (O_851,N_28295,N_28599);
xor UO_852 (O_852,N_28298,N_28135);
xor UO_853 (O_853,N_28254,N_29574);
nand UO_854 (O_854,N_29886,N_29135);
nand UO_855 (O_855,N_27594,N_27775);
and UO_856 (O_856,N_27564,N_28609);
nor UO_857 (O_857,N_28785,N_28574);
nor UO_858 (O_858,N_28151,N_29112);
or UO_859 (O_859,N_27766,N_28995);
and UO_860 (O_860,N_28360,N_27262);
or UO_861 (O_861,N_28533,N_29021);
nor UO_862 (O_862,N_28341,N_29625);
and UO_863 (O_863,N_29131,N_29964);
and UO_864 (O_864,N_29005,N_29228);
nor UO_865 (O_865,N_29333,N_27522);
and UO_866 (O_866,N_29891,N_28531);
xor UO_867 (O_867,N_28539,N_27978);
xnor UO_868 (O_868,N_29956,N_29233);
or UO_869 (O_869,N_28475,N_28131);
nor UO_870 (O_870,N_27175,N_27868);
nand UO_871 (O_871,N_27678,N_29571);
xnor UO_872 (O_872,N_29427,N_28764);
nand UO_873 (O_873,N_27643,N_28008);
or UO_874 (O_874,N_28824,N_28553);
xnor UO_875 (O_875,N_27636,N_29130);
nor UO_876 (O_876,N_28854,N_29726);
xor UO_877 (O_877,N_28499,N_27483);
nand UO_878 (O_878,N_29728,N_28153);
nand UO_879 (O_879,N_27263,N_28223);
and UO_880 (O_880,N_28866,N_28552);
and UO_881 (O_881,N_29346,N_27645);
nor UO_882 (O_882,N_29318,N_28725);
xnor UO_883 (O_883,N_27790,N_28169);
xnor UO_884 (O_884,N_29127,N_29236);
nor UO_885 (O_885,N_29108,N_28868);
nor UO_886 (O_886,N_27565,N_28710);
xor UO_887 (O_887,N_27740,N_29786);
nand UO_888 (O_888,N_28250,N_28612);
or UO_889 (O_889,N_29700,N_28407);
nor UO_890 (O_890,N_27398,N_29113);
nand UO_891 (O_891,N_27118,N_29968);
nor UO_892 (O_892,N_29270,N_28844);
nand UO_893 (O_893,N_27292,N_29330);
and UO_894 (O_894,N_29043,N_27835);
and UO_895 (O_895,N_27043,N_28030);
xor UO_896 (O_896,N_29795,N_27293);
or UO_897 (O_897,N_28773,N_29447);
xnor UO_898 (O_898,N_28643,N_28311);
nand UO_899 (O_899,N_28512,N_27786);
nor UO_900 (O_900,N_29282,N_27761);
nor UO_901 (O_901,N_29590,N_29283);
xor UO_902 (O_902,N_27874,N_29682);
nand UO_903 (O_903,N_27844,N_28670);
nand UO_904 (O_904,N_27279,N_29832);
xor UO_905 (O_905,N_27644,N_29081);
xor UO_906 (O_906,N_27515,N_29458);
and UO_907 (O_907,N_27639,N_28073);
and UO_908 (O_908,N_29733,N_29198);
nor UO_909 (O_909,N_27622,N_28222);
xnor UO_910 (O_910,N_27435,N_29770);
nand UO_911 (O_911,N_28800,N_27037);
xor UO_912 (O_912,N_28262,N_28130);
nor UO_913 (O_913,N_27425,N_27343);
or UO_914 (O_914,N_29158,N_28945);
or UO_915 (O_915,N_28788,N_28347);
nand UO_916 (O_916,N_29970,N_29879);
or UO_917 (O_917,N_27762,N_27591);
xnor UO_918 (O_918,N_28975,N_27290);
or UO_919 (O_919,N_27332,N_29273);
and UO_920 (O_920,N_28372,N_28658);
xnor UO_921 (O_921,N_29319,N_28366);
xor UO_922 (O_922,N_29175,N_28139);
nor UO_923 (O_923,N_28587,N_28048);
nand UO_924 (O_924,N_27438,N_28902);
xnor UO_925 (O_925,N_28856,N_28227);
nand UO_926 (O_926,N_27439,N_27910);
or UO_927 (O_927,N_29014,N_29411);
or UO_928 (O_928,N_28389,N_28320);
nand UO_929 (O_929,N_27666,N_29817);
nand UO_930 (O_930,N_27702,N_29877);
or UO_931 (O_931,N_29954,N_29086);
xnor UO_932 (O_932,N_29325,N_29100);
nand UO_933 (O_933,N_29444,N_27419);
nand UO_934 (O_934,N_27859,N_29776);
nor UO_935 (O_935,N_27756,N_27846);
nor UO_936 (O_936,N_27696,N_27849);
nand UO_937 (O_937,N_28627,N_27312);
or UO_938 (O_938,N_29229,N_27379);
xor UO_939 (O_939,N_28505,N_29774);
nand UO_940 (O_940,N_28126,N_27228);
and UO_941 (O_941,N_27110,N_29140);
and UO_942 (O_942,N_29920,N_27441);
nor UO_943 (O_943,N_27331,N_29986);
or UO_944 (O_944,N_29580,N_28970);
nor UO_945 (O_945,N_29489,N_28968);
and UO_946 (O_946,N_29149,N_29145);
and UO_947 (O_947,N_29210,N_29862);
nand UO_948 (O_948,N_27341,N_29822);
nor UO_949 (O_949,N_27559,N_28414);
and UO_950 (O_950,N_29162,N_27608);
or UO_951 (O_951,N_28726,N_27886);
xnor UO_952 (O_952,N_28107,N_29693);
nand UO_953 (O_953,N_27464,N_27296);
and UO_954 (O_954,N_27484,N_28544);
nor UO_955 (O_955,N_27993,N_27414);
or UO_956 (O_956,N_29582,N_28384);
nor UO_957 (O_957,N_28589,N_29136);
nand UO_958 (O_958,N_29530,N_29761);
xnor UO_959 (O_959,N_28792,N_28287);
or UO_960 (O_960,N_29711,N_28572);
nor UO_961 (O_961,N_27401,N_28207);
or UO_962 (O_962,N_28679,N_27215);
or UO_963 (O_963,N_27219,N_27054);
and UO_964 (O_964,N_27116,N_29812);
nand UO_965 (O_965,N_27975,N_27520);
or UO_966 (O_966,N_27873,N_28517);
or UO_967 (O_967,N_29310,N_28518);
nand UO_968 (O_968,N_28759,N_27626);
nand UO_969 (O_969,N_29479,N_29557);
and UO_970 (O_970,N_28344,N_28935);
nand UO_971 (O_971,N_29470,N_28959);
xor UO_972 (O_972,N_27654,N_28450);
xor UO_973 (O_973,N_29471,N_27214);
xnor UO_974 (O_974,N_27950,N_27631);
nor UO_975 (O_975,N_27885,N_27720);
or UO_976 (O_976,N_28029,N_28231);
and UO_977 (O_977,N_28750,N_28592);
nand UO_978 (O_978,N_27427,N_28722);
xnor UO_979 (O_979,N_29296,N_28628);
or UO_980 (O_980,N_29713,N_28084);
xnor UO_981 (O_981,N_27329,N_27123);
nand UO_982 (O_982,N_29807,N_27407);
or UO_983 (O_983,N_29932,N_27270);
and UO_984 (O_984,N_29029,N_29227);
nor UO_985 (O_985,N_27988,N_28294);
or UO_986 (O_986,N_27971,N_29480);
and UO_987 (O_987,N_27395,N_27490);
and UO_988 (O_988,N_27026,N_29450);
and UO_989 (O_989,N_27472,N_28695);
nor UO_990 (O_990,N_29988,N_27238);
and UO_991 (O_991,N_28748,N_28934);
and UO_992 (O_992,N_29119,N_27701);
nand UO_993 (O_993,N_29764,N_27381);
xor UO_994 (O_994,N_29267,N_29402);
nand UO_995 (O_995,N_27363,N_28321);
and UO_996 (O_996,N_27863,N_28211);
nor UO_997 (O_997,N_29323,N_27551);
and UO_998 (O_998,N_27691,N_28160);
xor UO_999 (O_999,N_27837,N_27576);
nand UO_1000 (O_1000,N_28374,N_29339);
xor UO_1001 (O_1001,N_27422,N_27791);
or UO_1002 (O_1002,N_29307,N_27570);
and UO_1003 (O_1003,N_28816,N_28569);
nand UO_1004 (O_1004,N_29507,N_29925);
or UO_1005 (O_1005,N_27342,N_28593);
and UO_1006 (O_1006,N_29633,N_29421);
and UO_1007 (O_1007,N_27836,N_27276);
xnor UO_1008 (O_1008,N_29718,N_27004);
and UO_1009 (O_1009,N_27368,N_29995);
nor UO_1010 (O_1010,N_29844,N_28708);
or UO_1011 (O_1011,N_29490,N_29207);
and UO_1012 (O_1012,N_27283,N_29141);
nor UO_1013 (O_1013,N_28083,N_27588);
and UO_1014 (O_1014,N_27627,N_27549);
and UO_1015 (O_1015,N_28864,N_27931);
nor UO_1016 (O_1016,N_29114,N_28702);
and UO_1017 (O_1017,N_27480,N_28996);
and UO_1018 (O_1018,N_28393,N_29422);
xor UO_1019 (O_1019,N_28386,N_29835);
xnor UO_1020 (O_1020,N_27317,N_27808);
or UO_1021 (O_1021,N_28875,N_28234);
or UO_1022 (O_1022,N_29985,N_28786);
nor UO_1023 (O_1023,N_28647,N_27495);
xor UO_1024 (O_1024,N_29508,N_29675);
and UO_1025 (O_1025,N_27670,N_27073);
nand UO_1026 (O_1026,N_27039,N_27278);
xor UO_1027 (O_1027,N_28758,N_27176);
xnor UO_1028 (O_1028,N_28443,N_27471);
nand UO_1029 (O_1029,N_27135,N_28279);
nor UO_1030 (O_1030,N_29120,N_28502);
xor UO_1031 (O_1031,N_28766,N_28999);
and UO_1032 (O_1032,N_29348,N_29876);
or UO_1033 (O_1033,N_29104,N_28014);
xnor UO_1034 (O_1034,N_29435,N_27890);
nand UO_1035 (O_1035,N_27017,N_27021);
nand UO_1036 (O_1036,N_29666,N_28749);
and UO_1037 (O_1037,N_29492,N_29929);
nand UO_1038 (O_1038,N_29316,N_28752);
or UO_1039 (O_1039,N_28522,N_28196);
nor UO_1040 (O_1040,N_28723,N_27310);
xor UO_1041 (O_1041,N_29919,N_28272);
and UO_1042 (O_1042,N_28837,N_28579);
nor UO_1043 (O_1043,N_29084,N_28200);
or UO_1044 (O_1044,N_29824,N_27473);
xnor UO_1045 (O_1045,N_29603,N_28843);
nor UO_1046 (O_1046,N_28164,N_29320);
nor UO_1047 (O_1047,N_27369,N_28779);
nor UO_1048 (O_1048,N_29860,N_28509);
or UO_1049 (O_1049,N_27616,N_27876);
and UO_1050 (O_1050,N_28883,N_28470);
nor UO_1051 (O_1051,N_29823,N_27072);
nor UO_1052 (O_1052,N_28554,N_28411);
and UO_1053 (O_1053,N_27482,N_28085);
nand UO_1054 (O_1054,N_27834,N_28404);
xor UO_1055 (O_1055,N_29059,N_29242);
nor UO_1056 (O_1056,N_29016,N_29334);
xnor UO_1057 (O_1057,N_29467,N_27528);
or UO_1058 (O_1058,N_29871,N_29134);
and UO_1059 (O_1059,N_29820,N_28345);
or UO_1060 (O_1060,N_29397,N_28168);
nand UO_1061 (O_1061,N_27373,N_28657);
and UO_1062 (O_1062,N_29913,N_29182);
xnor UO_1063 (O_1063,N_27286,N_29349);
nor UO_1064 (O_1064,N_27389,N_27460);
nor UO_1065 (O_1065,N_28885,N_27086);
and UO_1066 (O_1066,N_29547,N_27477);
nand UO_1067 (O_1067,N_28113,N_29749);
and UO_1068 (O_1068,N_28000,N_27813);
nand UO_1069 (O_1069,N_28354,N_27710);
nand UO_1070 (O_1070,N_29852,N_29758);
xnor UO_1071 (O_1071,N_28789,N_28607);
nor UO_1072 (O_1072,N_27272,N_29732);
xnor UO_1073 (O_1073,N_29023,N_28270);
and UO_1074 (O_1074,N_29948,N_28591);
xnor UO_1075 (O_1075,N_27903,N_29378);
and UO_1076 (O_1076,N_27773,N_29661);
nor UO_1077 (O_1077,N_27592,N_29055);
xor UO_1078 (O_1078,N_28224,N_27217);
nor UO_1079 (O_1079,N_28811,N_27783);
nor UO_1080 (O_1080,N_29364,N_27573);
nand UO_1081 (O_1081,N_28373,N_27029);
or UO_1082 (O_1082,N_28025,N_28529);
xnor UO_1083 (O_1083,N_27754,N_27424);
nand UO_1084 (O_1084,N_29924,N_29702);
nor UO_1085 (O_1085,N_29899,N_29454);
xor UO_1086 (O_1086,N_28422,N_28459);
nor UO_1087 (O_1087,N_27562,N_27092);
nand UO_1088 (O_1088,N_28661,N_29472);
xnor UO_1089 (O_1089,N_28565,N_28146);
or UO_1090 (O_1090,N_27739,N_29880);
or UO_1091 (O_1091,N_29833,N_29813);
or UO_1092 (O_1092,N_27277,N_29106);
and UO_1093 (O_1093,N_29406,N_29691);
and UO_1094 (O_1094,N_29982,N_28452);
nand UO_1095 (O_1095,N_28273,N_27216);
and UO_1096 (O_1096,N_27440,N_29504);
or UO_1097 (O_1097,N_27376,N_27494);
nand UO_1098 (O_1098,N_27926,N_29826);
or UO_1099 (O_1099,N_29984,N_29156);
xnor UO_1100 (O_1100,N_28908,N_29246);
and UO_1101 (O_1101,N_29617,N_29681);
nand UO_1102 (O_1102,N_27170,N_27614);
xor UO_1103 (O_1103,N_28891,N_27671);
or UO_1104 (O_1104,N_29658,N_27916);
nor UO_1105 (O_1105,N_27979,N_29011);
or UO_1106 (O_1106,N_28839,N_29022);
and UO_1107 (O_1107,N_27078,N_27646);
xor UO_1108 (O_1108,N_27470,N_27475);
nor UO_1109 (O_1109,N_28774,N_28819);
or UO_1110 (O_1110,N_28114,N_27532);
or UO_1111 (O_1111,N_27347,N_28269);
and UO_1112 (O_1112,N_27099,N_29080);
nor UO_1113 (O_1113,N_27413,N_29856);
nand UO_1114 (O_1114,N_27943,N_29915);
or UO_1115 (O_1115,N_28310,N_29742);
and UO_1116 (O_1116,N_29806,N_29456);
or UO_1117 (O_1117,N_29697,N_27340);
nor UO_1118 (O_1118,N_28356,N_28276);
or UO_1119 (O_1119,N_28071,N_28299);
nand UO_1120 (O_1120,N_29575,N_27543);
or UO_1121 (O_1121,N_28983,N_29650);
nand UO_1122 (O_1122,N_27919,N_27583);
and UO_1123 (O_1123,N_27335,N_27417);
and UO_1124 (O_1124,N_29281,N_29069);
xnor UO_1125 (O_1125,N_29315,N_28703);
or UO_1126 (O_1126,N_28926,N_28284);
xnor UO_1127 (O_1127,N_27810,N_27942);
and UO_1128 (O_1128,N_28631,N_27009);
nor UO_1129 (O_1129,N_28652,N_29783);
nand UO_1130 (O_1130,N_28142,N_27771);
xor UO_1131 (O_1131,N_29116,N_29741);
nor UO_1132 (O_1132,N_29680,N_27358);
or UO_1133 (O_1133,N_28985,N_27951);
or UO_1134 (O_1134,N_29446,N_28257);
and UO_1135 (O_1135,N_28061,N_27418);
and UO_1136 (O_1136,N_29208,N_27462);
nor UO_1137 (O_1137,N_28551,N_28698);
xor UO_1138 (O_1138,N_28297,N_28772);
nand UO_1139 (O_1139,N_28804,N_29451);
and UO_1140 (O_1140,N_28798,N_29550);
nand UO_1141 (O_1141,N_28534,N_29942);
nor UO_1142 (O_1142,N_27767,N_28119);
or UO_1143 (O_1143,N_29944,N_29466);
nor UO_1144 (O_1144,N_28871,N_28419);
nand UO_1145 (O_1145,N_29199,N_28625);
and UO_1146 (O_1146,N_27968,N_29857);
nand UO_1147 (O_1147,N_28380,N_29094);
xor UO_1148 (O_1148,N_29620,N_28964);
and UO_1149 (O_1149,N_28332,N_27663);
and UO_1150 (O_1150,N_28335,N_28852);
or UO_1151 (O_1151,N_28778,N_28237);
nor UO_1152 (O_1152,N_29585,N_27193);
and UO_1153 (O_1153,N_27084,N_28747);
xnor UO_1154 (O_1154,N_29195,N_28783);
nand UO_1155 (O_1155,N_28568,N_27361);
xor UO_1156 (O_1156,N_29361,N_28753);
nand UO_1157 (O_1157,N_27260,N_28056);
and UO_1158 (O_1158,N_28487,N_29738);
nand UO_1159 (O_1159,N_28989,N_27563);
or UO_1160 (O_1160,N_28917,N_28203);
xor UO_1161 (O_1161,N_29226,N_28218);
xor UO_1162 (O_1162,N_28074,N_28106);
or UO_1163 (O_1163,N_29160,N_29940);
xnor UO_1164 (O_1164,N_28878,N_29542);
nor UO_1165 (O_1165,N_27064,N_27751);
nor UO_1166 (O_1166,N_28024,N_27246);
and UO_1167 (O_1167,N_28680,N_27182);
nand UO_1168 (O_1168,N_28846,N_27558);
nand UO_1169 (O_1169,N_29593,N_27450);
and UO_1170 (O_1170,N_28597,N_29202);
nand UO_1171 (O_1171,N_27618,N_29324);
nand UO_1172 (O_1172,N_27202,N_27778);
and UO_1173 (O_1173,N_29401,N_28095);
xnor UO_1174 (O_1174,N_28195,N_28988);
nand UO_1175 (O_1175,N_29789,N_29171);
xnor UO_1176 (O_1176,N_27102,N_28900);
or UO_1177 (O_1177,N_28873,N_29851);
and UO_1178 (O_1178,N_28253,N_27164);
or UO_1179 (O_1179,N_28687,N_27452);
or UO_1180 (O_1180,N_28051,N_27298);
or UO_1181 (O_1181,N_27185,N_27948);
nand UO_1182 (O_1182,N_27437,N_27047);
and UO_1183 (O_1183,N_27755,N_28474);
xor UO_1184 (O_1184,N_28100,N_28979);
xor UO_1185 (O_1185,N_27183,N_27224);
nor UO_1186 (O_1186,N_27250,N_29563);
xnor UO_1187 (O_1187,N_28980,N_28521);
nand UO_1188 (O_1188,N_27366,N_28922);
xnor UO_1189 (O_1189,N_29203,N_28929);
nand UO_1190 (O_1190,N_27865,N_29911);
and UO_1191 (O_1191,N_28542,N_28641);
and UO_1192 (O_1192,N_28576,N_28405);
nand UO_1193 (O_1193,N_29218,N_27063);
nand UO_1194 (O_1194,N_29843,N_28904);
and UO_1195 (O_1195,N_28220,N_28527);
or UO_1196 (O_1196,N_29255,N_28520);
nand UO_1197 (O_1197,N_27003,N_27223);
nand UO_1198 (O_1198,N_27640,N_27680);
nand UO_1199 (O_1199,N_29253,N_27303);
nor UO_1200 (O_1200,N_27326,N_29337);
nor UO_1201 (O_1201,N_28756,N_29241);
or UO_1202 (O_1202,N_27752,N_27731);
nand UO_1203 (O_1203,N_27206,N_27222);
and UO_1204 (O_1204,N_28850,N_28441);
nor UO_1205 (O_1205,N_27878,N_28721);
nor UO_1206 (O_1206,N_27656,N_27195);
xnor UO_1207 (O_1207,N_28526,N_27662);
nand UO_1208 (O_1208,N_28034,N_29341);
nand UO_1209 (O_1209,N_27304,N_28801);
or UO_1210 (O_1210,N_27140,N_27036);
xor UO_1211 (O_1211,N_28765,N_28745);
and UO_1212 (O_1212,N_28715,N_28958);
nor UO_1213 (O_1213,N_28060,N_27220);
nor UO_1214 (O_1214,N_29442,N_27348);
or UO_1215 (O_1215,N_27218,N_28302);
nand UO_1216 (O_1216,N_29109,N_27274);
and UO_1217 (O_1217,N_29850,N_27336);
or UO_1218 (O_1218,N_27842,N_28585);
xnor UO_1219 (O_1219,N_27983,N_28331);
or UO_1220 (O_1220,N_27245,N_29405);
or UO_1221 (O_1221,N_29276,N_27186);
xnor UO_1222 (O_1222,N_29989,N_28210);
and UO_1223 (O_1223,N_28963,N_29641);
and UO_1224 (O_1224,N_27963,N_29274);
nor UO_1225 (O_1225,N_29883,N_28212);
nor UO_1226 (O_1226,N_27337,N_29587);
or UO_1227 (O_1227,N_29186,N_29192);
and UO_1228 (O_1228,N_29000,N_27095);
xnor UO_1229 (O_1229,N_27871,N_29359);
nor UO_1230 (O_1230,N_27044,N_29872);
and UO_1231 (O_1231,N_29694,N_28144);
nand UO_1232 (O_1232,N_28089,N_27600);
xor UO_1233 (O_1233,N_27019,N_29355);
xor UO_1234 (O_1234,N_28742,N_28586);
or UO_1235 (O_1235,N_27061,N_29384);
nand UO_1236 (O_1236,N_29801,N_29595);
or UO_1237 (O_1237,N_27325,N_27599);
nand UO_1238 (O_1238,N_27787,N_28010);
or UO_1239 (O_1239,N_29373,N_27144);
nand UO_1240 (O_1240,N_27200,N_28112);
and UO_1241 (O_1241,N_29665,N_27561);
nor UO_1242 (O_1242,N_27991,N_29293);
nand UO_1243 (O_1243,N_29600,N_28510);
or UO_1244 (O_1244,N_27602,N_29214);
nand UO_1245 (O_1245,N_28198,N_29819);
and UO_1246 (O_1246,N_28796,N_29369);
and UO_1247 (O_1247,N_29394,N_28735);
nand UO_1248 (O_1248,N_29651,N_27529);
nand UO_1249 (O_1249,N_27305,N_28076);
xnor UO_1250 (O_1250,N_28751,N_29748);
and UO_1251 (O_1251,N_29714,N_29260);
nand UO_1252 (O_1252,N_28434,N_27349);
or UO_1253 (O_1253,N_29567,N_29024);
xor UO_1254 (O_1254,N_29304,N_29115);
nand UO_1255 (O_1255,N_29166,N_28007);
nand UO_1256 (O_1256,N_29096,N_27713);
xnor UO_1257 (O_1257,N_27541,N_29431);
nand UO_1258 (O_1258,N_29332,N_27709);
xor UO_1259 (O_1259,N_27689,N_28770);
and UO_1260 (O_1260,N_28194,N_28711);
nand UO_1261 (O_1261,N_29379,N_27763);
xnor UO_1262 (O_1262,N_27261,N_29522);
and UO_1263 (O_1263,N_29735,N_28235);
xnor UO_1264 (O_1264,N_27253,N_28767);
nor UO_1265 (O_1265,N_29914,N_27126);
nand UO_1266 (O_1266,N_28528,N_27251);
nor UO_1267 (O_1267,N_28420,N_27733);
nand UO_1268 (O_1268,N_29418,N_29562);
nand UO_1269 (O_1269,N_27028,N_28709);
nor UO_1270 (O_1270,N_28952,N_29586);
and UO_1271 (O_1271,N_29759,N_28097);
and UO_1272 (O_1272,N_28190,N_27847);
nand UO_1273 (O_1273,N_28660,N_29124);
nand UO_1274 (O_1274,N_28736,N_29413);
nor UO_1275 (O_1275,N_28261,N_27540);
nor UO_1276 (O_1276,N_27143,N_27649);
and UO_1277 (O_1277,N_27350,N_28141);
and UO_1278 (O_1278,N_27211,N_27474);
and UO_1279 (O_1279,N_29383,N_27032);
nand UO_1280 (O_1280,N_27481,N_28462);
or UO_1281 (O_1281,N_27499,N_28739);
and UO_1282 (O_1282,N_27115,N_27409);
or UO_1283 (O_1283,N_29781,N_29482);
nand UO_1284 (O_1284,N_29473,N_28049);
or UO_1285 (O_1285,N_28762,N_28149);
xor UO_1286 (O_1286,N_29342,N_27536);
xor UO_1287 (O_1287,N_27149,N_28479);
or UO_1288 (O_1288,N_27375,N_28870);
xnor UO_1289 (O_1289,N_27394,N_27909);
nand UO_1290 (O_1290,N_29387,N_28435);
nand UO_1291 (O_1291,N_29873,N_28727);
nor UO_1292 (O_1292,N_27530,N_29429);
or UO_1293 (O_1293,N_28401,N_28403);
xor UO_1294 (O_1294,N_28157,N_28039);
and UO_1295 (O_1295,N_28673,N_27936);
or UO_1296 (O_1296,N_27467,N_28233);
and UO_1297 (O_1297,N_27630,N_29535);
or UO_1298 (O_1298,N_29426,N_29017);
xor UO_1299 (O_1299,N_27256,N_29465);
or UO_1300 (O_1300,N_29151,N_29437);
nand UO_1301 (O_1301,N_27196,N_27316);
and UO_1302 (O_1302,N_27548,N_27575);
and UO_1303 (O_1303,N_28693,N_29771);
nor UO_1304 (O_1304,N_28780,N_29885);
nor UO_1305 (O_1305,N_27606,N_28485);
nand UO_1306 (O_1306,N_27012,N_28588);
nor UO_1307 (O_1307,N_28712,N_28663);
nand UO_1308 (O_1308,N_29058,N_28241);
xnor UO_1309 (O_1309,N_27020,N_29533);
nor UO_1310 (O_1310,N_28383,N_29305);
nor UO_1311 (O_1311,N_28893,N_28152);
and UO_1312 (O_1312,N_29510,N_29647);
or UO_1313 (O_1313,N_29814,N_29597);
nand UO_1314 (O_1314,N_28226,N_27601);
or UO_1315 (O_1315,N_28064,N_29103);
and UO_1316 (O_1316,N_28651,N_28953);
nand UO_1317 (O_1317,N_27938,N_27056);
nor UO_1318 (O_1318,N_27005,N_27852);
nor UO_1319 (O_1319,N_29184,N_28480);
and UO_1320 (O_1320,N_29154,N_29350);
nand UO_1321 (O_1321,N_28636,N_27199);
nor UO_1322 (O_1322,N_27901,N_27093);
and UO_1323 (O_1323,N_27109,N_27371);
or UO_1324 (O_1324,N_29065,N_27508);
and UO_1325 (O_1325,N_27904,N_27638);
nor UO_1326 (O_1326,N_28449,N_27688);
and UO_1327 (O_1327,N_28165,N_29994);
nor UO_1328 (O_1328,N_29695,N_29760);
or UO_1329 (O_1329,N_27567,N_29941);
nand UO_1330 (O_1330,N_29264,N_28430);
or UO_1331 (O_1331,N_27087,N_29063);
xnor UO_1332 (O_1332,N_27002,N_28524);
xor UO_1333 (O_1333,N_29893,N_27465);
xor UO_1334 (O_1334,N_28497,N_28733);
xnor UO_1335 (O_1335,N_27221,N_27234);
and UO_1336 (O_1336,N_27569,N_29513);
nand UO_1337 (O_1337,N_29345,N_28809);
nor UO_1338 (O_1338,N_28969,N_29370);
nor UO_1339 (O_1339,N_28197,N_27209);
xor UO_1340 (O_1340,N_29825,N_29818);
xor UO_1341 (O_1341,N_27893,N_28183);
nor UO_1342 (O_1342,N_29224,N_27053);
nor UO_1343 (O_1343,N_27237,N_27134);
nor UO_1344 (O_1344,N_27081,N_28730);
or UO_1345 (O_1345,N_29725,N_28312);
or UO_1346 (O_1346,N_28961,N_28371);
xnor UO_1347 (O_1347,N_29803,N_27798);
nand UO_1348 (O_1348,N_28163,N_27067);
nor UO_1349 (O_1349,N_28043,N_27352);
and UO_1350 (O_1350,N_27924,N_27996);
xor UO_1351 (O_1351,N_28635,N_27659);
or UO_1352 (O_1352,N_28933,N_27556);
nor UO_1353 (O_1353,N_29621,N_29505);
and UO_1354 (O_1354,N_27489,N_29126);
nand UO_1355 (O_1355,N_27166,N_27492);
nand UO_1356 (O_1356,N_28363,N_28937);
or UO_1357 (O_1357,N_28826,N_27461);
nand UO_1358 (O_1358,N_27920,N_29815);
and UO_1359 (O_1359,N_28277,N_28318);
nand UO_1360 (O_1360,N_29570,N_27396);
xor UO_1361 (O_1361,N_29285,N_29834);
nor UO_1362 (O_1362,N_29155,N_29375);
or UO_1363 (O_1363,N_28944,N_29773);
nor UO_1364 (O_1364,N_28249,N_29308);
or UO_1365 (O_1365,N_29897,N_27703);
and UO_1366 (O_1366,N_27586,N_27829);
and UO_1367 (O_1367,N_28966,N_28382);
nor UO_1368 (O_1368,N_29036,N_27632);
nor UO_1369 (O_1369,N_28556,N_29743);
xnor UO_1370 (O_1370,N_28763,N_28115);
or UO_1371 (O_1371,N_27574,N_29147);
nor UO_1372 (O_1372,N_28705,N_28410);
and UO_1373 (O_1373,N_27811,N_28683);
nor UO_1374 (O_1374,N_28887,N_29026);
nand UO_1375 (O_1375,N_28187,N_27881);
xor UO_1376 (O_1376,N_28308,N_28650);
and UO_1377 (O_1377,N_28716,N_29618);
nor UO_1378 (O_1378,N_29904,N_29044);
nand UO_1379 (O_1379,N_28110,N_28901);
xnor UO_1380 (O_1380,N_29727,N_27932);
or UO_1381 (O_1381,N_28971,N_29935);
nand UO_1382 (O_1382,N_29441,N_27990);
xor UO_1383 (O_1383,N_27210,N_27383);
nand UO_1384 (O_1384,N_29057,N_28905);
xnor UO_1385 (O_1385,N_29183,N_27027);
or UO_1386 (O_1386,N_29710,N_27819);
nand UO_1387 (O_1387,N_27034,N_28340);
or UO_1388 (O_1388,N_29677,N_27457);
nand UO_1389 (O_1389,N_28116,N_29892);
nand UO_1390 (O_1390,N_29194,N_29257);
nor UO_1391 (O_1391,N_28713,N_28070);
or UO_1392 (O_1392,N_27380,N_29975);
nor UO_1393 (O_1393,N_28096,N_29598);
and UO_1394 (O_1394,N_28810,N_27721);
or UO_1395 (O_1395,N_28515,N_27949);
or UO_1396 (O_1396,N_28481,N_27468);
and UO_1397 (O_1397,N_27857,N_27891);
and UO_1398 (O_1398,N_29900,N_29707);
or UO_1399 (O_1399,N_29854,N_29309);
or UO_1400 (O_1400,N_29034,N_27768);
and UO_1401 (O_1401,N_27879,N_29712);
nor UO_1402 (O_1402,N_29779,N_27459);
or UO_1403 (O_1403,N_27776,N_28790);
and UO_1404 (O_1404,N_29512,N_28994);
or UO_1405 (O_1405,N_29365,N_27315);
nor UO_1406 (O_1406,N_28326,N_29966);
nor UO_1407 (O_1407,N_29196,N_29487);
nand UO_1408 (O_1408,N_29559,N_29947);
xor UO_1409 (O_1409,N_27454,N_28275);
xnor UO_1410 (O_1410,N_29927,N_27266);
nor UO_1411 (O_1411,N_27922,N_29343);
nand UO_1412 (O_1412,N_27364,N_28699);
or UO_1413 (O_1413,N_28425,N_28737);
nand UO_1414 (O_1414,N_28392,N_29075);
xor UO_1415 (O_1415,N_27212,N_27239);
or UO_1416 (O_1416,N_28936,N_28938);
nor UO_1417 (O_1417,N_28455,N_28688);
or UO_1418 (O_1418,N_28444,N_27955);
xor UO_1419 (O_1419,N_29662,N_27531);
and UO_1420 (O_1420,N_28467,N_29730);
nor UO_1421 (O_1421,N_27107,N_29290);
nand UO_1422 (O_1422,N_29744,N_29907);
nand UO_1423 (O_1423,N_28293,N_27362);
and UO_1424 (O_1424,N_28817,N_28924);
or UO_1425 (O_1425,N_29672,N_28877);
and UO_1426 (O_1426,N_27799,N_29245);
nor UO_1427 (O_1427,N_28033,N_28672);
nand UO_1428 (O_1428,N_29696,N_27513);
and UO_1429 (O_1429,N_28267,N_27338);
nand UO_1430 (O_1430,N_27953,N_27385);
and UO_1431 (O_1431,N_27537,N_27511);
nor UO_1432 (O_1432,N_29085,N_28192);
or UO_1433 (O_1433,N_29366,N_28408);
nor UO_1434 (O_1434,N_27075,N_29498);
nand UO_1435 (O_1435,N_28570,N_29040);
or UO_1436 (O_1436,N_29906,N_28882);
nand UO_1437 (O_1437,N_28300,N_29419);
nand UO_1438 (O_1438,N_27151,N_27096);
nor UO_1439 (O_1439,N_27172,N_29053);
nand UO_1440 (O_1440,N_27378,N_28504);
nand UO_1441 (O_1441,N_29128,N_28511);
nor UO_1442 (O_1442,N_29791,N_28829);
nand UO_1443 (O_1443,N_27408,N_29583);
nor UO_1444 (O_1444,N_29389,N_28943);
xor UO_1445 (O_1445,N_29056,N_29093);
nand UO_1446 (O_1446,N_29045,N_27684);
xor UO_1447 (O_1447,N_28466,N_27945);
nand UO_1448 (O_1448,N_27507,N_28993);
or UO_1449 (O_1449,N_27584,N_29972);
xnor UO_1450 (O_1450,N_29889,N_27737);
nand UO_1451 (O_1451,N_27147,N_27797);
xnor UO_1452 (O_1452,N_29659,N_27792);
and UO_1453 (O_1453,N_29099,N_29616);
or UO_1454 (O_1454,N_28464,N_29306);
and UO_1455 (O_1455,N_28062,N_27704);
nor UO_1456 (O_1456,N_29193,N_27416);
nand UO_1457 (O_1457,N_29327,N_28604);
nand UO_1458 (O_1458,N_29980,N_29001);
nand UO_1459 (O_1459,N_29243,N_27735);
xor UO_1460 (O_1460,N_27194,N_27554);
nor UO_1461 (O_1461,N_29684,N_29500);
or UO_1462 (O_1462,N_28600,N_29626);
and UO_1463 (O_1463,N_27386,N_27597);
or UO_1464 (O_1464,N_28682,N_27610);
nand UO_1465 (O_1465,N_27637,N_28044);
or UO_1466 (O_1466,N_27906,N_28012);
or UO_1467 (O_1467,N_29502,N_28385);
nand UO_1468 (O_1468,N_27669,N_28216);
nand UO_1469 (O_1469,N_29592,N_27119);
nor UO_1470 (O_1470,N_29443,N_28398);
nor UO_1471 (O_1471,N_27641,N_29438);
or UO_1472 (O_1472,N_27302,N_27190);
or UO_1473 (O_1473,N_29841,N_29881);
nand UO_1474 (O_1474,N_28507,N_27726);
nand UO_1475 (O_1475,N_28743,N_28626);
nor UO_1476 (O_1476,N_29167,N_29328);
xor UO_1477 (O_1477,N_28337,N_28696);
and UO_1478 (O_1478,N_29638,N_28329);
and UO_1479 (O_1479,N_27921,N_27802);
or UO_1480 (O_1480,N_29209,N_28714);
xnor UO_1481 (O_1481,N_28128,N_29457);
xor UO_1482 (O_1482,N_28803,N_27478);
nor UO_1483 (O_1483,N_29353,N_28268);
nor UO_1484 (O_1484,N_29299,N_29572);
or UO_1485 (O_1485,N_27059,N_28155);
xnor UO_1486 (O_1486,N_27794,N_29558);
nand UO_1487 (O_1487,N_29863,N_27213);
nand UO_1488 (O_1488,N_27856,N_29962);
xnor UO_1489 (O_1489,N_28219,N_29655);
nand UO_1490 (O_1490,N_27913,N_29206);
nand UO_1491 (O_1491,N_29107,N_27907);
nor UO_1492 (O_1492,N_28581,N_27257);
nor UO_1493 (O_1493,N_27273,N_29090);
xnor UO_1494 (O_1494,N_27882,N_28840);
nand UO_1495 (O_1495,N_27354,N_27828);
xnor UO_1496 (O_1496,N_28897,N_29796);
or UO_1497 (O_1497,N_29928,N_27772);
and UO_1498 (O_1498,N_28493,N_28797);
nand UO_1499 (O_1499,N_28053,N_29689);
xor UO_1500 (O_1500,N_27332,N_28765);
and UO_1501 (O_1501,N_28088,N_28293);
xnor UO_1502 (O_1502,N_27127,N_28775);
xnor UO_1503 (O_1503,N_28388,N_29892);
and UO_1504 (O_1504,N_29110,N_28583);
or UO_1505 (O_1505,N_27734,N_28429);
or UO_1506 (O_1506,N_28420,N_28939);
or UO_1507 (O_1507,N_29680,N_28509);
and UO_1508 (O_1508,N_28671,N_28916);
nand UO_1509 (O_1509,N_28945,N_27589);
and UO_1510 (O_1510,N_27242,N_27611);
nor UO_1511 (O_1511,N_29076,N_29561);
or UO_1512 (O_1512,N_29409,N_28688);
nor UO_1513 (O_1513,N_28800,N_27248);
nand UO_1514 (O_1514,N_27093,N_27429);
and UO_1515 (O_1515,N_27244,N_28595);
xnor UO_1516 (O_1516,N_27692,N_29481);
nor UO_1517 (O_1517,N_29199,N_27543);
and UO_1518 (O_1518,N_28181,N_27931);
nand UO_1519 (O_1519,N_27106,N_29657);
or UO_1520 (O_1520,N_29373,N_28338);
nor UO_1521 (O_1521,N_27681,N_27342);
or UO_1522 (O_1522,N_29290,N_29945);
nor UO_1523 (O_1523,N_28065,N_27899);
nand UO_1524 (O_1524,N_27299,N_28907);
nor UO_1525 (O_1525,N_28335,N_29410);
nand UO_1526 (O_1526,N_27103,N_29833);
and UO_1527 (O_1527,N_29794,N_29606);
and UO_1528 (O_1528,N_27163,N_29846);
or UO_1529 (O_1529,N_28304,N_28969);
nand UO_1530 (O_1530,N_28262,N_27036);
or UO_1531 (O_1531,N_27277,N_28325);
or UO_1532 (O_1532,N_29017,N_28726);
xor UO_1533 (O_1533,N_29873,N_28239);
nor UO_1534 (O_1534,N_27019,N_27662);
nand UO_1535 (O_1535,N_29378,N_29333);
and UO_1536 (O_1536,N_27808,N_28475);
and UO_1537 (O_1537,N_27798,N_29575);
nor UO_1538 (O_1538,N_29243,N_27230);
xor UO_1539 (O_1539,N_28435,N_29973);
and UO_1540 (O_1540,N_29691,N_27894);
nand UO_1541 (O_1541,N_28299,N_27799);
nand UO_1542 (O_1542,N_28476,N_29374);
and UO_1543 (O_1543,N_28451,N_28018);
xnor UO_1544 (O_1544,N_28587,N_28273);
nand UO_1545 (O_1545,N_27799,N_27796);
nand UO_1546 (O_1546,N_28680,N_29564);
and UO_1547 (O_1547,N_29363,N_27012);
and UO_1548 (O_1548,N_27079,N_27333);
nor UO_1549 (O_1549,N_27925,N_29678);
or UO_1550 (O_1550,N_28113,N_28905);
or UO_1551 (O_1551,N_28200,N_29167);
and UO_1552 (O_1552,N_29171,N_29643);
or UO_1553 (O_1553,N_28917,N_28393);
nand UO_1554 (O_1554,N_28572,N_29383);
nand UO_1555 (O_1555,N_27981,N_28528);
nor UO_1556 (O_1556,N_27627,N_27007);
and UO_1557 (O_1557,N_29230,N_28231);
nor UO_1558 (O_1558,N_27735,N_28677);
nand UO_1559 (O_1559,N_29172,N_27690);
nand UO_1560 (O_1560,N_29773,N_27191);
nor UO_1561 (O_1561,N_29461,N_28064);
or UO_1562 (O_1562,N_29541,N_28074);
and UO_1563 (O_1563,N_29098,N_28499);
or UO_1564 (O_1564,N_28543,N_28939);
nand UO_1565 (O_1565,N_29197,N_28570);
xor UO_1566 (O_1566,N_27976,N_29501);
nor UO_1567 (O_1567,N_28527,N_29363);
xnor UO_1568 (O_1568,N_27503,N_28187);
nor UO_1569 (O_1569,N_29761,N_27203);
or UO_1570 (O_1570,N_28526,N_29470);
nor UO_1571 (O_1571,N_28662,N_29613);
xor UO_1572 (O_1572,N_29282,N_29044);
xnor UO_1573 (O_1573,N_27321,N_29422);
nand UO_1574 (O_1574,N_28927,N_29239);
nor UO_1575 (O_1575,N_27484,N_29306);
nor UO_1576 (O_1576,N_28657,N_28011);
and UO_1577 (O_1577,N_27703,N_29610);
xor UO_1578 (O_1578,N_27137,N_28554);
xnor UO_1579 (O_1579,N_29955,N_28556);
and UO_1580 (O_1580,N_28986,N_27405);
nand UO_1581 (O_1581,N_28899,N_28093);
nor UO_1582 (O_1582,N_28143,N_28202);
and UO_1583 (O_1583,N_29041,N_28938);
nor UO_1584 (O_1584,N_27026,N_27528);
xor UO_1585 (O_1585,N_27943,N_28735);
or UO_1586 (O_1586,N_27600,N_29183);
xor UO_1587 (O_1587,N_29093,N_28483);
or UO_1588 (O_1588,N_28781,N_28364);
nand UO_1589 (O_1589,N_29398,N_27981);
xor UO_1590 (O_1590,N_29040,N_27589);
nand UO_1591 (O_1591,N_29286,N_28597);
or UO_1592 (O_1592,N_28653,N_29109);
and UO_1593 (O_1593,N_29249,N_29197);
nor UO_1594 (O_1594,N_27167,N_29804);
xor UO_1595 (O_1595,N_27707,N_27052);
nor UO_1596 (O_1596,N_27746,N_28506);
xor UO_1597 (O_1597,N_27959,N_28255);
nor UO_1598 (O_1598,N_28585,N_29311);
xor UO_1599 (O_1599,N_27458,N_29996);
and UO_1600 (O_1600,N_27824,N_28966);
nor UO_1601 (O_1601,N_29626,N_29091);
or UO_1602 (O_1602,N_29711,N_27253);
xor UO_1603 (O_1603,N_27450,N_29410);
or UO_1604 (O_1604,N_29066,N_27707);
nand UO_1605 (O_1605,N_27037,N_27264);
nor UO_1606 (O_1606,N_28271,N_28722);
nor UO_1607 (O_1607,N_27176,N_28168);
or UO_1608 (O_1608,N_29892,N_29760);
nand UO_1609 (O_1609,N_29838,N_28993);
or UO_1610 (O_1610,N_28141,N_29360);
nand UO_1611 (O_1611,N_28261,N_27846);
nand UO_1612 (O_1612,N_27589,N_28144);
and UO_1613 (O_1613,N_29116,N_29823);
or UO_1614 (O_1614,N_28034,N_28283);
xnor UO_1615 (O_1615,N_29225,N_27802);
nand UO_1616 (O_1616,N_29791,N_28210);
nand UO_1617 (O_1617,N_29476,N_29615);
xnor UO_1618 (O_1618,N_29112,N_28802);
or UO_1619 (O_1619,N_27575,N_29386);
nor UO_1620 (O_1620,N_29002,N_27003);
or UO_1621 (O_1621,N_29340,N_29866);
and UO_1622 (O_1622,N_27904,N_29878);
nor UO_1623 (O_1623,N_29291,N_28648);
and UO_1624 (O_1624,N_27746,N_28763);
and UO_1625 (O_1625,N_27420,N_27162);
and UO_1626 (O_1626,N_27501,N_27403);
and UO_1627 (O_1627,N_28153,N_28197);
and UO_1628 (O_1628,N_28602,N_29195);
nor UO_1629 (O_1629,N_27829,N_27622);
nand UO_1630 (O_1630,N_29222,N_27354);
nand UO_1631 (O_1631,N_28243,N_29790);
nand UO_1632 (O_1632,N_29614,N_29441);
and UO_1633 (O_1633,N_27568,N_28233);
and UO_1634 (O_1634,N_27658,N_27864);
or UO_1635 (O_1635,N_29616,N_28770);
or UO_1636 (O_1636,N_27901,N_29127);
nand UO_1637 (O_1637,N_27797,N_27352);
and UO_1638 (O_1638,N_28211,N_27710);
nand UO_1639 (O_1639,N_27727,N_28170);
nor UO_1640 (O_1640,N_28288,N_29556);
or UO_1641 (O_1641,N_28760,N_29159);
and UO_1642 (O_1642,N_29605,N_28833);
and UO_1643 (O_1643,N_29192,N_29460);
and UO_1644 (O_1644,N_27442,N_29817);
and UO_1645 (O_1645,N_29034,N_27196);
xnor UO_1646 (O_1646,N_29490,N_28655);
and UO_1647 (O_1647,N_29152,N_28729);
or UO_1648 (O_1648,N_28006,N_29933);
nand UO_1649 (O_1649,N_27721,N_27884);
nand UO_1650 (O_1650,N_29083,N_27673);
xnor UO_1651 (O_1651,N_27227,N_28470);
nor UO_1652 (O_1652,N_29959,N_29681);
or UO_1653 (O_1653,N_29900,N_28879);
or UO_1654 (O_1654,N_29341,N_29309);
or UO_1655 (O_1655,N_28302,N_27429);
nor UO_1656 (O_1656,N_28810,N_27483);
xnor UO_1657 (O_1657,N_29022,N_27200);
nand UO_1658 (O_1658,N_29159,N_29709);
and UO_1659 (O_1659,N_29858,N_27246);
or UO_1660 (O_1660,N_28464,N_29452);
nand UO_1661 (O_1661,N_27957,N_28303);
nand UO_1662 (O_1662,N_28094,N_28437);
and UO_1663 (O_1663,N_27765,N_27889);
xor UO_1664 (O_1664,N_29311,N_27443);
and UO_1665 (O_1665,N_29708,N_28618);
xor UO_1666 (O_1666,N_28529,N_28496);
nor UO_1667 (O_1667,N_28808,N_28640);
and UO_1668 (O_1668,N_27710,N_27791);
nand UO_1669 (O_1669,N_29210,N_29651);
or UO_1670 (O_1670,N_28066,N_29144);
xor UO_1671 (O_1671,N_29665,N_27013);
xnor UO_1672 (O_1672,N_29914,N_28681);
nand UO_1673 (O_1673,N_27915,N_28375);
and UO_1674 (O_1674,N_29629,N_28572);
and UO_1675 (O_1675,N_28175,N_28437);
nand UO_1676 (O_1676,N_29400,N_28572);
and UO_1677 (O_1677,N_29067,N_28427);
nand UO_1678 (O_1678,N_28639,N_28069);
xor UO_1679 (O_1679,N_29439,N_27492);
xor UO_1680 (O_1680,N_29292,N_28856);
nand UO_1681 (O_1681,N_27128,N_29970);
and UO_1682 (O_1682,N_29625,N_29666);
nand UO_1683 (O_1683,N_29606,N_27719);
xor UO_1684 (O_1684,N_28202,N_29132);
or UO_1685 (O_1685,N_28619,N_29732);
xor UO_1686 (O_1686,N_27778,N_28273);
or UO_1687 (O_1687,N_29755,N_27588);
and UO_1688 (O_1688,N_27297,N_27567);
nand UO_1689 (O_1689,N_28308,N_29136);
nor UO_1690 (O_1690,N_28202,N_28209);
and UO_1691 (O_1691,N_27616,N_27024);
nor UO_1692 (O_1692,N_27188,N_28808);
or UO_1693 (O_1693,N_28141,N_27368);
and UO_1694 (O_1694,N_29557,N_27421);
nand UO_1695 (O_1695,N_29252,N_27731);
and UO_1696 (O_1696,N_27508,N_28902);
and UO_1697 (O_1697,N_29516,N_29935);
nand UO_1698 (O_1698,N_29043,N_29466);
or UO_1699 (O_1699,N_29108,N_29938);
nand UO_1700 (O_1700,N_27387,N_28982);
xor UO_1701 (O_1701,N_28295,N_27894);
xnor UO_1702 (O_1702,N_28021,N_28109);
nand UO_1703 (O_1703,N_28624,N_27167);
or UO_1704 (O_1704,N_28828,N_28417);
nand UO_1705 (O_1705,N_27062,N_29122);
nor UO_1706 (O_1706,N_27813,N_28004);
or UO_1707 (O_1707,N_27539,N_28544);
or UO_1708 (O_1708,N_29591,N_29812);
or UO_1709 (O_1709,N_28557,N_29829);
or UO_1710 (O_1710,N_29018,N_29880);
xnor UO_1711 (O_1711,N_28225,N_27607);
xor UO_1712 (O_1712,N_29517,N_27760);
nor UO_1713 (O_1713,N_27549,N_27330);
xnor UO_1714 (O_1714,N_27823,N_27488);
nor UO_1715 (O_1715,N_28388,N_28681);
xor UO_1716 (O_1716,N_28248,N_29795);
nand UO_1717 (O_1717,N_29970,N_27535);
and UO_1718 (O_1718,N_27857,N_28580);
or UO_1719 (O_1719,N_29790,N_29540);
nand UO_1720 (O_1720,N_28313,N_29486);
xnor UO_1721 (O_1721,N_27937,N_28967);
or UO_1722 (O_1722,N_29312,N_29205);
and UO_1723 (O_1723,N_28719,N_27779);
xnor UO_1724 (O_1724,N_27166,N_28563);
xnor UO_1725 (O_1725,N_29872,N_27193);
or UO_1726 (O_1726,N_27106,N_28636);
nand UO_1727 (O_1727,N_28555,N_27586);
or UO_1728 (O_1728,N_28951,N_29553);
or UO_1729 (O_1729,N_28361,N_29267);
or UO_1730 (O_1730,N_27990,N_27586);
and UO_1731 (O_1731,N_28657,N_29986);
nor UO_1732 (O_1732,N_29085,N_27434);
nand UO_1733 (O_1733,N_28117,N_28343);
nand UO_1734 (O_1734,N_28126,N_28926);
or UO_1735 (O_1735,N_29863,N_29052);
nor UO_1736 (O_1736,N_29506,N_28759);
nand UO_1737 (O_1737,N_28301,N_29943);
xor UO_1738 (O_1738,N_28994,N_29785);
and UO_1739 (O_1739,N_27873,N_29853);
xor UO_1740 (O_1740,N_28592,N_27934);
or UO_1741 (O_1741,N_27141,N_27143);
and UO_1742 (O_1742,N_27768,N_29579);
and UO_1743 (O_1743,N_29935,N_29279);
nor UO_1744 (O_1744,N_29243,N_27842);
nand UO_1745 (O_1745,N_28267,N_28927);
nand UO_1746 (O_1746,N_28410,N_27829);
nor UO_1747 (O_1747,N_29987,N_27917);
nor UO_1748 (O_1748,N_28179,N_28655);
nand UO_1749 (O_1749,N_27794,N_28663);
nand UO_1750 (O_1750,N_29623,N_29855);
xor UO_1751 (O_1751,N_27450,N_29157);
nor UO_1752 (O_1752,N_27865,N_28267);
xor UO_1753 (O_1753,N_27155,N_28705);
nand UO_1754 (O_1754,N_27248,N_27217);
or UO_1755 (O_1755,N_27980,N_27238);
nor UO_1756 (O_1756,N_29921,N_27136);
and UO_1757 (O_1757,N_28843,N_27630);
nand UO_1758 (O_1758,N_28901,N_29145);
nor UO_1759 (O_1759,N_28375,N_28955);
xor UO_1760 (O_1760,N_27039,N_29001);
nand UO_1761 (O_1761,N_29937,N_27986);
or UO_1762 (O_1762,N_27820,N_27315);
and UO_1763 (O_1763,N_28704,N_29623);
and UO_1764 (O_1764,N_29202,N_28310);
and UO_1765 (O_1765,N_28282,N_29757);
nand UO_1766 (O_1766,N_28721,N_27777);
xor UO_1767 (O_1767,N_29969,N_28731);
or UO_1768 (O_1768,N_28899,N_27409);
xor UO_1769 (O_1769,N_27207,N_27184);
xnor UO_1770 (O_1770,N_27208,N_28580);
xor UO_1771 (O_1771,N_29132,N_29660);
nor UO_1772 (O_1772,N_29132,N_29698);
nor UO_1773 (O_1773,N_28027,N_29630);
xnor UO_1774 (O_1774,N_29172,N_27756);
and UO_1775 (O_1775,N_27981,N_28569);
nor UO_1776 (O_1776,N_29112,N_28164);
or UO_1777 (O_1777,N_27191,N_29046);
xor UO_1778 (O_1778,N_28731,N_28497);
nor UO_1779 (O_1779,N_27091,N_29937);
nand UO_1780 (O_1780,N_29814,N_27640);
nand UO_1781 (O_1781,N_29387,N_27607);
nand UO_1782 (O_1782,N_27732,N_27406);
nor UO_1783 (O_1783,N_29505,N_28629);
or UO_1784 (O_1784,N_27979,N_28349);
and UO_1785 (O_1785,N_27873,N_27196);
nand UO_1786 (O_1786,N_29218,N_29060);
xor UO_1787 (O_1787,N_28570,N_27067);
and UO_1788 (O_1788,N_28770,N_28817);
nor UO_1789 (O_1789,N_28986,N_29295);
xnor UO_1790 (O_1790,N_28859,N_27070);
or UO_1791 (O_1791,N_27805,N_29878);
xnor UO_1792 (O_1792,N_28783,N_29039);
and UO_1793 (O_1793,N_28155,N_28141);
and UO_1794 (O_1794,N_27080,N_28029);
or UO_1795 (O_1795,N_28768,N_27783);
nor UO_1796 (O_1796,N_28282,N_29753);
and UO_1797 (O_1797,N_28589,N_29350);
and UO_1798 (O_1798,N_29242,N_27210);
nand UO_1799 (O_1799,N_28461,N_28056);
xnor UO_1800 (O_1800,N_28785,N_27670);
and UO_1801 (O_1801,N_29457,N_27455);
xor UO_1802 (O_1802,N_28951,N_28357);
and UO_1803 (O_1803,N_27601,N_27509);
nor UO_1804 (O_1804,N_27013,N_27560);
nor UO_1805 (O_1805,N_27407,N_28513);
nor UO_1806 (O_1806,N_29640,N_27509);
or UO_1807 (O_1807,N_29904,N_27658);
nor UO_1808 (O_1808,N_28789,N_27968);
or UO_1809 (O_1809,N_29243,N_29835);
and UO_1810 (O_1810,N_29582,N_27561);
or UO_1811 (O_1811,N_29105,N_28440);
nand UO_1812 (O_1812,N_29953,N_27999);
nor UO_1813 (O_1813,N_28735,N_28106);
and UO_1814 (O_1814,N_27812,N_27303);
and UO_1815 (O_1815,N_29058,N_27147);
and UO_1816 (O_1816,N_29981,N_29083);
and UO_1817 (O_1817,N_29289,N_29757);
or UO_1818 (O_1818,N_27275,N_29672);
xnor UO_1819 (O_1819,N_27125,N_28438);
and UO_1820 (O_1820,N_29321,N_29081);
nor UO_1821 (O_1821,N_29526,N_27377);
or UO_1822 (O_1822,N_27251,N_27524);
and UO_1823 (O_1823,N_27133,N_29617);
nand UO_1824 (O_1824,N_28030,N_28659);
nor UO_1825 (O_1825,N_28370,N_28789);
or UO_1826 (O_1826,N_28139,N_27611);
and UO_1827 (O_1827,N_28944,N_28921);
xor UO_1828 (O_1828,N_27263,N_29690);
and UO_1829 (O_1829,N_27304,N_27389);
nand UO_1830 (O_1830,N_27185,N_28156);
nor UO_1831 (O_1831,N_27190,N_28650);
nand UO_1832 (O_1832,N_29171,N_29682);
and UO_1833 (O_1833,N_28807,N_27020);
nor UO_1834 (O_1834,N_27803,N_29487);
nand UO_1835 (O_1835,N_28816,N_29543);
xor UO_1836 (O_1836,N_28167,N_28600);
nor UO_1837 (O_1837,N_29134,N_28725);
and UO_1838 (O_1838,N_28802,N_29035);
nand UO_1839 (O_1839,N_27879,N_27218);
or UO_1840 (O_1840,N_29856,N_29908);
xor UO_1841 (O_1841,N_29749,N_28187);
nor UO_1842 (O_1842,N_27156,N_29528);
nor UO_1843 (O_1843,N_27418,N_29408);
xnor UO_1844 (O_1844,N_28232,N_27878);
nand UO_1845 (O_1845,N_29702,N_28110);
or UO_1846 (O_1846,N_27345,N_28008);
nor UO_1847 (O_1847,N_28028,N_29194);
nor UO_1848 (O_1848,N_27056,N_27947);
or UO_1849 (O_1849,N_28555,N_27611);
and UO_1850 (O_1850,N_29220,N_28734);
and UO_1851 (O_1851,N_29937,N_28093);
or UO_1852 (O_1852,N_28079,N_29208);
nor UO_1853 (O_1853,N_28057,N_28535);
and UO_1854 (O_1854,N_29374,N_28566);
or UO_1855 (O_1855,N_29006,N_28762);
nand UO_1856 (O_1856,N_28047,N_27112);
or UO_1857 (O_1857,N_27256,N_27095);
nand UO_1858 (O_1858,N_29722,N_29634);
nand UO_1859 (O_1859,N_29789,N_27866);
nor UO_1860 (O_1860,N_28416,N_27983);
nand UO_1861 (O_1861,N_28209,N_27377);
xnor UO_1862 (O_1862,N_27999,N_29795);
or UO_1863 (O_1863,N_29006,N_29637);
nand UO_1864 (O_1864,N_27721,N_29757);
or UO_1865 (O_1865,N_29929,N_29413);
or UO_1866 (O_1866,N_28764,N_28565);
xor UO_1867 (O_1867,N_27455,N_28816);
nand UO_1868 (O_1868,N_27383,N_29872);
xor UO_1869 (O_1869,N_27841,N_28687);
and UO_1870 (O_1870,N_29912,N_28615);
and UO_1871 (O_1871,N_29554,N_27694);
nand UO_1872 (O_1872,N_29602,N_27249);
or UO_1873 (O_1873,N_28766,N_29469);
and UO_1874 (O_1874,N_27247,N_27825);
nor UO_1875 (O_1875,N_27876,N_27640);
or UO_1876 (O_1876,N_27487,N_28422);
nand UO_1877 (O_1877,N_27026,N_29981);
or UO_1878 (O_1878,N_29289,N_29991);
and UO_1879 (O_1879,N_28890,N_27415);
xor UO_1880 (O_1880,N_27389,N_29106);
nor UO_1881 (O_1881,N_27815,N_27430);
and UO_1882 (O_1882,N_27135,N_27827);
xnor UO_1883 (O_1883,N_29060,N_28811);
and UO_1884 (O_1884,N_29928,N_29786);
xor UO_1885 (O_1885,N_27122,N_28310);
xor UO_1886 (O_1886,N_29135,N_27048);
nand UO_1887 (O_1887,N_27742,N_28793);
or UO_1888 (O_1888,N_28978,N_28594);
nand UO_1889 (O_1889,N_29279,N_29144);
xor UO_1890 (O_1890,N_29512,N_27009);
xnor UO_1891 (O_1891,N_28342,N_29598);
xor UO_1892 (O_1892,N_28471,N_29950);
xor UO_1893 (O_1893,N_28198,N_29395);
nor UO_1894 (O_1894,N_29209,N_29526);
nand UO_1895 (O_1895,N_27640,N_29619);
xnor UO_1896 (O_1896,N_28184,N_28633);
nand UO_1897 (O_1897,N_27734,N_27057);
nand UO_1898 (O_1898,N_29746,N_28626);
or UO_1899 (O_1899,N_29216,N_27574);
xor UO_1900 (O_1900,N_27779,N_27653);
xnor UO_1901 (O_1901,N_29266,N_29575);
nand UO_1902 (O_1902,N_29401,N_27560);
nor UO_1903 (O_1903,N_28566,N_29092);
nor UO_1904 (O_1904,N_27849,N_27609);
nand UO_1905 (O_1905,N_28529,N_27171);
nand UO_1906 (O_1906,N_27232,N_28634);
or UO_1907 (O_1907,N_29605,N_29074);
and UO_1908 (O_1908,N_28085,N_28531);
nor UO_1909 (O_1909,N_27647,N_28221);
nand UO_1910 (O_1910,N_27282,N_28490);
or UO_1911 (O_1911,N_28428,N_27732);
nor UO_1912 (O_1912,N_29432,N_28986);
xor UO_1913 (O_1913,N_29328,N_27813);
nor UO_1914 (O_1914,N_28421,N_28086);
or UO_1915 (O_1915,N_29636,N_27861);
and UO_1916 (O_1916,N_29288,N_28233);
nor UO_1917 (O_1917,N_27398,N_29718);
xnor UO_1918 (O_1918,N_27141,N_28202);
or UO_1919 (O_1919,N_28734,N_28987);
nand UO_1920 (O_1920,N_28743,N_27176);
and UO_1921 (O_1921,N_28184,N_27615);
nor UO_1922 (O_1922,N_29986,N_27386);
xor UO_1923 (O_1923,N_27690,N_29670);
nor UO_1924 (O_1924,N_27245,N_29925);
or UO_1925 (O_1925,N_28633,N_27938);
or UO_1926 (O_1926,N_28347,N_29400);
nand UO_1927 (O_1927,N_29893,N_27551);
nand UO_1928 (O_1928,N_28905,N_27399);
or UO_1929 (O_1929,N_27148,N_27946);
nor UO_1930 (O_1930,N_27870,N_29310);
nand UO_1931 (O_1931,N_29054,N_29398);
nor UO_1932 (O_1932,N_28750,N_28703);
and UO_1933 (O_1933,N_29181,N_27131);
and UO_1934 (O_1934,N_28526,N_28529);
nand UO_1935 (O_1935,N_29601,N_28243);
and UO_1936 (O_1936,N_29296,N_29038);
xor UO_1937 (O_1937,N_28718,N_29469);
and UO_1938 (O_1938,N_28952,N_29511);
nand UO_1939 (O_1939,N_28755,N_27047);
nor UO_1940 (O_1940,N_29214,N_29080);
nand UO_1941 (O_1941,N_28070,N_29710);
and UO_1942 (O_1942,N_27252,N_28538);
nor UO_1943 (O_1943,N_28058,N_29598);
and UO_1944 (O_1944,N_29665,N_28433);
nor UO_1945 (O_1945,N_29061,N_28684);
xor UO_1946 (O_1946,N_28723,N_29014);
xnor UO_1947 (O_1947,N_28506,N_29968);
nor UO_1948 (O_1948,N_29572,N_27718);
xnor UO_1949 (O_1949,N_28353,N_28888);
or UO_1950 (O_1950,N_29581,N_29777);
nand UO_1951 (O_1951,N_27116,N_29031);
xnor UO_1952 (O_1952,N_28671,N_27628);
and UO_1953 (O_1953,N_29042,N_28640);
nor UO_1954 (O_1954,N_28394,N_27948);
and UO_1955 (O_1955,N_29625,N_27444);
and UO_1956 (O_1956,N_29713,N_28700);
and UO_1957 (O_1957,N_28081,N_29793);
or UO_1958 (O_1958,N_29021,N_28331);
and UO_1959 (O_1959,N_28274,N_28126);
nor UO_1960 (O_1960,N_29359,N_27154);
nor UO_1961 (O_1961,N_27365,N_29332);
and UO_1962 (O_1962,N_29893,N_29825);
and UO_1963 (O_1963,N_27459,N_27449);
and UO_1964 (O_1964,N_27033,N_29563);
or UO_1965 (O_1965,N_28596,N_28743);
xnor UO_1966 (O_1966,N_29215,N_28101);
nor UO_1967 (O_1967,N_29661,N_27666);
nor UO_1968 (O_1968,N_28794,N_29340);
and UO_1969 (O_1969,N_29190,N_28585);
or UO_1970 (O_1970,N_27086,N_27617);
nor UO_1971 (O_1971,N_27605,N_28486);
xnor UO_1972 (O_1972,N_29016,N_29573);
nand UO_1973 (O_1973,N_29338,N_27627);
or UO_1974 (O_1974,N_27554,N_27790);
nand UO_1975 (O_1975,N_28076,N_29340);
nor UO_1976 (O_1976,N_28990,N_29674);
and UO_1977 (O_1977,N_29097,N_27862);
xnor UO_1978 (O_1978,N_28995,N_29669);
and UO_1979 (O_1979,N_27382,N_27205);
and UO_1980 (O_1980,N_27962,N_27354);
or UO_1981 (O_1981,N_27852,N_29675);
or UO_1982 (O_1982,N_29532,N_28643);
and UO_1983 (O_1983,N_29635,N_28575);
nand UO_1984 (O_1984,N_27782,N_28784);
xor UO_1985 (O_1985,N_28656,N_27825);
or UO_1986 (O_1986,N_27445,N_28155);
nor UO_1987 (O_1987,N_27890,N_29180);
nor UO_1988 (O_1988,N_27170,N_29048);
nand UO_1989 (O_1989,N_27251,N_28445);
nand UO_1990 (O_1990,N_27996,N_27063);
xor UO_1991 (O_1991,N_28064,N_29890);
nand UO_1992 (O_1992,N_29489,N_29235);
and UO_1993 (O_1993,N_28621,N_29330);
or UO_1994 (O_1994,N_27691,N_27802);
nand UO_1995 (O_1995,N_27719,N_27003);
nand UO_1996 (O_1996,N_28097,N_28551);
nor UO_1997 (O_1997,N_29844,N_29702);
xor UO_1998 (O_1998,N_27487,N_28027);
nor UO_1999 (O_1999,N_27086,N_28934);
and UO_2000 (O_2000,N_28760,N_27629);
xnor UO_2001 (O_2001,N_28285,N_27511);
xnor UO_2002 (O_2002,N_29480,N_29180);
xnor UO_2003 (O_2003,N_29072,N_29322);
nand UO_2004 (O_2004,N_28696,N_28983);
or UO_2005 (O_2005,N_28603,N_28230);
nand UO_2006 (O_2006,N_27781,N_29407);
and UO_2007 (O_2007,N_27915,N_28350);
or UO_2008 (O_2008,N_28290,N_29400);
or UO_2009 (O_2009,N_28284,N_27878);
nor UO_2010 (O_2010,N_27419,N_27575);
xnor UO_2011 (O_2011,N_28501,N_28185);
or UO_2012 (O_2012,N_29569,N_28306);
or UO_2013 (O_2013,N_28461,N_27032);
nand UO_2014 (O_2014,N_28503,N_28929);
and UO_2015 (O_2015,N_29295,N_29312);
nor UO_2016 (O_2016,N_29371,N_29303);
and UO_2017 (O_2017,N_27383,N_28286);
nand UO_2018 (O_2018,N_28555,N_28966);
nor UO_2019 (O_2019,N_27362,N_27016);
and UO_2020 (O_2020,N_29190,N_28712);
nor UO_2021 (O_2021,N_27766,N_27080);
or UO_2022 (O_2022,N_28181,N_27726);
or UO_2023 (O_2023,N_29486,N_27406);
nor UO_2024 (O_2024,N_29064,N_28106);
and UO_2025 (O_2025,N_28825,N_28385);
and UO_2026 (O_2026,N_27623,N_29365);
nor UO_2027 (O_2027,N_28120,N_29544);
and UO_2028 (O_2028,N_28084,N_28522);
xor UO_2029 (O_2029,N_29535,N_27389);
or UO_2030 (O_2030,N_28630,N_27111);
nor UO_2031 (O_2031,N_27366,N_28253);
or UO_2032 (O_2032,N_29664,N_29265);
nand UO_2033 (O_2033,N_28118,N_28237);
nand UO_2034 (O_2034,N_28935,N_28004);
and UO_2035 (O_2035,N_27277,N_28427);
nand UO_2036 (O_2036,N_28404,N_28911);
or UO_2037 (O_2037,N_27467,N_29318);
or UO_2038 (O_2038,N_27680,N_27294);
and UO_2039 (O_2039,N_27316,N_28161);
nor UO_2040 (O_2040,N_28489,N_28257);
and UO_2041 (O_2041,N_27108,N_27384);
or UO_2042 (O_2042,N_27569,N_28887);
or UO_2043 (O_2043,N_27970,N_28156);
and UO_2044 (O_2044,N_29441,N_27751);
and UO_2045 (O_2045,N_29733,N_29678);
and UO_2046 (O_2046,N_27246,N_27716);
nand UO_2047 (O_2047,N_29629,N_27000);
or UO_2048 (O_2048,N_28536,N_27057);
xnor UO_2049 (O_2049,N_28974,N_27692);
and UO_2050 (O_2050,N_28488,N_27202);
and UO_2051 (O_2051,N_29332,N_27780);
or UO_2052 (O_2052,N_28824,N_28537);
nand UO_2053 (O_2053,N_29634,N_29396);
or UO_2054 (O_2054,N_29449,N_27974);
and UO_2055 (O_2055,N_27286,N_28111);
xor UO_2056 (O_2056,N_29385,N_27327);
and UO_2057 (O_2057,N_29094,N_29346);
nor UO_2058 (O_2058,N_27228,N_27945);
or UO_2059 (O_2059,N_27629,N_27515);
nand UO_2060 (O_2060,N_29352,N_28858);
xnor UO_2061 (O_2061,N_28963,N_27917);
and UO_2062 (O_2062,N_29979,N_29877);
xnor UO_2063 (O_2063,N_27161,N_29695);
and UO_2064 (O_2064,N_27426,N_27787);
nand UO_2065 (O_2065,N_28540,N_28287);
and UO_2066 (O_2066,N_27506,N_28739);
xnor UO_2067 (O_2067,N_28744,N_29477);
and UO_2068 (O_2068,N_29983,N_27513);
nor UO_2069 (O_2069,N_28490,N_28360);
nor UO_2070 (O_2070,N_29135,N_28874);
and UO_2071 (O_2071,N_29781,N_27065);
xnor UO_2072 (O_2072,N_27576,N_28525);
or UO_2073 (O_2073,N_29667,N_27764);
nand UO_2074 (O_2074,N_29712,N_27155);
nor UO_2075 (O_2075,N_29564,N_28749);
xnor UO_2076 (O_2076,N_27175,N_28017);
nor UO_2077 (O_2077,N_29338,N_29373);
or UO_2078 (O_2078,N_29114,N_27685);
or UO_2079 (O_2079,N_28991,N_27646);
or UO_2080 (O_2080,N_29539,N_28997);
or UO_2081 (O_2081,N_28678,N_27750);
and UO_2082 (O_2082,N_28143,N_27718);
nand UO_2083 (O_2083,N_27920,N_28304);
nor UO_2084 (O_2084,N_28073,N_29071);
or UO_2085 (O_2085,N_29500,N_28760);
nand UO_2086 (O_2086,N_27774,N_28520);
xnor UO_2087 (O_2087,N_28266,N_27787);
nand UO_2088 (O_2088,N_28859,N_28985);
and UO_2089 (O_2089,N_29820,N_28960);
nand UO_2090 (O_2090,N_29944,N_29950);
or UO_2091 (O_2091,N_29953,N_28860);
and UO_2092 (O_2092,N_27108,N_28835);
xor UO_2093 (O_2093,N_29979,N_27848);
and UO_2094 (O_2094,N_27938,N_29103);
nand UO_2095 (O_2095,N_28036,N_27409);
and UO_2096 (O_2096,N_28602,N_29413);
nand UO_2097 (O_2097,N_29157,N_28103);
nor UO_2098 (O_2098,N_29181,N_27721);
nor UO_2099 (O_2099,N_29037,N_29141);
nand UO_2100 (O_2100,N_29464,N_29271);
or UO_2101 (O_2101,N_28224,N_27624);
xnor UO_2102 (O_2102,N_28877,N_29216);
nand UO_2103 (O_2103,N_29264,N_27181);
xnor UO_2104 (O_2104,N_27145,N_27826);
nand UO_2105 (O_2105,N_28831,N_28210);
xor UO_2106 (O_2106,N_28991,N_28071);
or UO_2107 (O_2107,N_27856,N_28631);
nor UO_2108 (O_2108,N_28037,N_27846);
or UO_2109 (O_2109,N_27207,N_28124);
xor UO_2110 (O_2110,N_28062,N_27338);
nand UO_2111 (O_2111,N_28911,N_27163);
nor UO_2112 (O_2112,N_27078,N_28421);
and UO_2113 (O_2113,N_27344,N_29360);
or UO_2114 (O_2114,N_28992,N_27427);
xnor UO_2115 (O_2115,N_28826,N_29752);
nand UO_2116 (O_2116,N_28192,N_27658);
or UO_2117 (O_2117,N_27454,N_28008);
nor UO_2118 (O_2118,N_27630,N_27186);
xor UO_2119 (O_2119,N_27507,N_28259);
and UO_2120 (O_2120,N_28275,N_29611);
nand UO_2121 (O_2121,N_27047,N_28285);
and UO_2122 (O_2122,N_27084,N_29898);
nand UO_2123 (O_2123,N_27266,N_29541);
or UO_2124 (O_2124,N_27597,N_27272);
nand UO_2125 (O_2125,N_27157,N_27344);
or UO_2126 (O_2126,N_27312,N_27664);
nand UO_2127 (O_2127,N_27581,N_28922);
xor UO_2128 (O_2128,N_28837,N_28964);
or UO_2129 (O_2129,N_29771,N_27568);
nor UO_2130 (O_2130,N_28632,N_29603);
nand UO_2131 (O_2131,N_28687,N_28293);
or UO_2132 (O_2132,N_29648,N_28884);
nand UO_2133 (O_2133,N_27070,N_27357);
and UO_2134 (O_2134,N_29909,N_29090);
xnor UO_2135 (O_2135,N_29772,N_27855);
and UO_2136 (O_2136,N_29510,N_29578);
or UO_2137 (O_2137,N_29455,N_28034);
and UO_2138 (O_2138,N_29302,N_29143);
nor UO_2139 (O_2139,N_27987,N_28076);
nand UO_2140 (O_2140,N_29451,N_29290);
and UO_2141 (O_2141,N_27213,N_27865);
nand UO_2142 (O_2142,N_29104,N_28135);
nor UO_2143 (O_2143,N_28802,N_27426);
xor UO_2144 (O_2144,N_29467,N_28134);
nor UO_2145 (O_2145,N_28890,N_29798);
and UO_2146 (O_2146,N_28844,N_28469);
xnor UO_2147 (O_2147,N_29314,N_28984);
xor UO_2148 (O_2148,N_27345,N_27872);
nor UO_2149 (O_2149,N_28747,N_29165);
or UO_2150 (O_2150,N_27863,N_28780);
xnor UO_2151 (O_2151,N_27543,N_28279);
and UO_2152 (O_2152,N_29483,N_27728);
nand UO_2153 (O_2153,N_27222,N_27453);
xnor UO_2154 (O_2154,N_28297,N_27365);
nand UO_2155 (O_2155,N_27449,N_28081);
xor UO_2156 (O_2156,N_28908,N_27076);
or UO_2157 (O_2157,N_28142,N_29973);
and UO_2158 (O_2158,N_29843,N_28423);
and UO_2159 (O_2159,N_27730,N_27024);
nand UO_2160 (O_2160,N_29585,N_27497);
xor UO_2161 (O_2161,N_28159,N_28756);
nand UO_2162 (O_2162,N_29566,N_29604);
and UO_2163 (O_2163,N_29751,N_28650);
and UO_2164 (O_2164,N_28078,N_28582);
nand UO_2165 (O_2165,N_27993,N_29799);
xor UO_2166 (O_2166,N_27787,N_27317);
nor UO_2167 (O_2167,N_27189,N_29810);
and UO_2168 (O_2168,N_27258,N_29805);
or UO_2169 (O_2169,N_29646,N_27901);
nor UO_2170 (O_2170,N_28791,N_29050);
and UO_2171 (O_2171,N_27311,N_27285);
nand UO_2172 (O_2172,N_28396,N_27109);
and UO_2173 (O_2173,N_27731,N_28890);
nand UO_2174 (O_2174,N_28223,N_27548);
nor UO_2175 (O_2175,N_28634,N_28115);
nor UO_2176 (O_2176,N_27267,N_28691);
and UO_2177 (O_2177,N_27101,N_29893);
xor UO_2178 (O_2178,N_28062,N_29420);
xnor UO_2179 (O_2179,N_28002,N_29337);
nand UO_2180 (O_2180,N_27912,N_28022);
or UO_2181 (O_2181,N_28603,N_29450);
xor UO_2182 (O_2182,N_29250,N_28502);
xor UO_2183 (O_2183,N_27466,N_27590);
nand UO_2184 (O_2184,N_28532,N_28640);
xor UO_2185 (O_2185,N_28168,N_29237);
and UO_2186 (O_2186,N_28656,N_28512);
and UO_2187 (O_2187,N_28670,N_27231);
nand UO_2188 (O_2188,N_27175,N_29316);
nor UO_2189 (O_2189,N_28534,N_28384);
xor UO_2190 (O_2190,N_27977,N_27465);
and UO_2191 (O_2191,N_29189,N_29718);
nand UO_2192 (O_2192,N_27552,N_28415);
nand UO_2193 (O_2193,N_29234,N_28277);
xnor UO_2194 (O_2194,N_27041,N_27294);
xnor UO_2195 (O_2195,N_29633,N_27934);
xor UO_2196 (O_2196,N_29161,N_29825);
or UO_2197 (O_2197,N_28565,N_29748);
xor UO_2198 (O_2198,N_27032,N_28053);
nor UO_2199 (O_2199,N_27529,N_28534);
and UO_2200 (O_2200,N_29565,N_28104);
xor UO_2201 (O_2201,N_29367,N_29299);
or UO_2202 (O_2202,N_29772,N_28327);
nand UO_2203 (O_2203,N_28981,N_29624);
and UO_2204 (O_2204,N_29989,N_28594);
and UO_2205 (O_2205,N_28447,N_28082);
xor UO_2206 (O_2206,N_27767,N_29104);
and UO_2207 (O_2207,N_27546,N_27568);
and UO_2208 (O_2208,N_28797,N_27756);
or UO_2209 (O_2209,N_27019,N_27782);
xnor UO_2210 (O_2210,N_27142,N_29821);
xnor UO_2211 (O_2211,N_29123,N_28189);
nand UO_2212 (O_2212,N_29139,N_27643);
xor UO_2213 (O_2213,N_29737,N_28785);
or UO_2214 (O_2214,N_27455,N_28243);
nor UO_2215 (O_2215,N_28654,N_27836);
nand UO_2216 (O_2216,N_29563,N_27979);
or UO_2217 (O_2217,N_29987,N_29306);
and UO_2218 (O_2218,N_28235,N_27687);
nor UO_2219 (O_2219,N_27134,N_27347);
and UO_2220 (O_2220,N_28006,N_27176);
and UO_2221 (O_2221,N_28715,N_28669);
nor UO_2222 (O_2222,N_27559,N_27769);
nand UO_2223 (O_2223,N_28056,N_27464);
nand UO_2224 (O_2224,N_27468,N_27447);
or UO_2225 (O_2225,N_29125,N_29402);
xnor UO_2226 (O_2226,N_29123,N_28373);
nand UO_2227 (O_2227,N_29766,N_27660);
or UO_2228 (O_2228,N_28108,N_29506);
nand UO_2229 (O_2229,N_28492,N_27821);
nor UO_2230 (O_2230,N_27052,N_29970);
nand UO_2231 (O_2231,N_27338,N_28489);
nand UO_2232 (O_2232,N_27068,N_27817);
and UO_2233 (O_2233,N_28460,N_28127);
or UO_2234 (O_2234,N_28843,N_29304);
or UO_2235 (O_2235,N_29609,N_27412);
nand UO_2236 (O_2236,N_29520,N_29322);
or UO_2237 (O_2237,N_27525,N_28505);
nand UO_2238 (O_2238,N_27752,N_29873);
nor UO_2239 (O_2239,N_29716,N_29248);
and UO_2240 (O_2240,N_28595,N_29371);
and UO_2241 (O_2241,N_29143,N_29466);
nand UO_2242 (O_2242,N_28696,N_29540);
xor UO_2243 (O_2243,N_28859,N_29873);
nand UO_2244 (O_2244,N_28107,N_28383);
or UO_2245 (O_2245,N_28399,N_29793);
nand UO_2246 (O_2246,N_27715,N_28595);
or UO_2247 (O_2247,N_29160,N_28240);
and UO_2248 (O_2248,N_29488,N_27005);
nand UO_2249 (O_2249,N_29221,N_27036);
nor UO_2250 (O_2250,N_27097,N_27010);
or UO_2251 (O_2251,N_27725,N_27215);
nor UO_2252 (O_2252,N_27086,N_27658);
and UO_2253 (O_2253,N_27795,N_27998);
and UO_2254 (O_2254,N_29127,N_28111);
nand UO_2255 (O_2255,N_29772,N_29060);
nand UO_2256 (O_2256,N_27599,N_29289);
and UO_2257 (O_2257,N_29068,N_29288);
xnor UO_2258 (O_2258,N_29369,N_27567);
or UO_2259 (O_2259,N_27401,N_27561);
xor UO_2260 (O_2260,N_29620,N_28985);
nand UO_2261 (O_2261,N_28552,N_29652);
and UO_2262 (O_2262,N_28206,N_27954);
nor UO_2263 (O_2263,N_29902,N_29693);
and UO_2264 (O_2264,N_28191,N_28333);
nor UO_2265 (O_2265,N_29709,N_28763);
and UO_2266 (O_2266,N_29072,N_28285);
or UO_2267 (O_2267,N_27765,N_27388);
nor UO_2268 (O_2268,N_28584,N_27950);
or UO_2269 (O_2269,N_29841,N_27483);
xnor UO_2270 (O_2270,N_27471,N_28064);
and UO_2271 (O_2271,N_28007,N_27211);
xnor UO_2272 (O_2272,N_29020,N_29144);
nand UO_2273 (O_2273,N_29446,N_27318);
nand UO_2274 (O_2274,N_29077,N_27076);
xnor UO_2275 (O_2275,N_29703,N_29301);
xor UO_2276 (O_2276,N_28477,N_28354);
or UO_2277 (O_2277,N_29482,N_29958);
and UO_2278 (O_2278,N_29870,N_29400);
and UO_2279 (O_2279,N_29516,N_28721);
or UO_2280 (O_2280,N_27879,N_28223);
or UO_2281 (O_2281,N_28033,N_29850);
and UO_2282 (O_2282,N_28359,N_29434);
nor UO_2283 (O_2283,N_28705,N_29280);
xor UO_2284 (O_2284,N_27298,N_28830);
nor UO_2285 (O_2285,N_28285,N_29953);
or UO_2286 (O_2286,N_28732,N_28212);
nor UO_2287 (O_2287,N_29063,N_28753);
nand UO_2288 (O_2288,N_27120,N_29899);
xor UO_2289 (O_2289,N_28290,N_27964);
or UO_2290 (O_2290,N_27036,N_28885);
xor UO_2291 (O_2291,N_29838,N_29506);
nand UO_2292 (O_2292,N_28597,N_28203);
nor UO_2293 (O_2293,N_29275,N_27900);
or UO_2294 (O_2294,N_29871,N_27512);
or UO_2295 (O_2295,N_29175,N_28795);
nand UO_2296 (O_2296,N_29333,N_27327);
and UO_2297 (O_2297,N_29317,N_27244);
or UO_2298 (O_2298,N_28769,N_27281);
and UO_2299 (O_2299,N_27389,N_29737);
nor UO_2300 (O_2300,N_27682,N_27185);
or UO_2301 (O_2301,N_28283,N_27292);
xor UO_2302 (O_2302,N_29713,N_27890);
and UO_2303 (O_2303,N_28164,N_27583);
xor UO_2304 (O_2304,N_28616,N_28859);
and UO_2305 (O_2305,N_28611,N_29872);
xnor UO_2306 (O_2306,N_28058,N_28037);
and UO_2307 (O_2307,N_28340,N_29643);
nor UO_2308 (O_2308,N_27174,N_29232);
nor UO_2309 (O_2309,N_29401,N_28696);
nand UO_2310 (O_2310,N_29357,N_27615);
xnor UO_2311 (O_2311,N_28230,N_28621);
or UO_2312 (O_2312,N_28795,N_27354);
or UO_2313 (O_2313,N_27684,N_28145);
or UO_2314 (O_2314,N_28135,N_29159);
xnor UO_2315 (O_2315,N_28035,N_28391);
or UO_2316 (O_2316,N_29130,N_27288);
nor UO_2317 (O_2317,N_28285,N_29817);
or UO_2318 (O_2318,N_27100,N_28115);
nor UO_2319 (O_2319,N_29997,N_27992);
nand UO_2320 (O_2320,N_27457,N_29389);
nand UO_2321 (O_2321,N_27445,N_27885);
nand UO_2322 (O_2322,N_27969,N_29949);
xnor UO_2323 (O_2323,N_28016,N_28676);
nand UO_2324 (O_2324,N_28923,N_27445);
and UO_2325 (O_2325,N_29179,N_28150);
or UO_2326 (O_2326,N_27087,N_28492);
and UO_2327 (O_2327,N_27347,N_28679);
nand UO_2328 (O_2328,N_29836,N_28854);
and UO_2329 (O_2329,N_28791,N_28069);
nor UO_2330 (O_2330,N_27439,N_27409);
xnor UO_2331 (O_2331,N_27159,N_27833);
nor UO_2332 (O_2332,N_28422,N_29281);
nor UO_2333 (O_2333,N_28777,N_28319);
xnor UO_2334 (O_2334,N_27903,N_29145);
and UO_2335 (O_2335,N_29251,N_29631);
or UO_2336 (O_2336,N_29541,N_28828);
nand UO_2337 (O_2337,N_29901,N_27026);
nor UO_2338 (O_2338,N_27125,N_29243);
nor UO_2339 (O_2339,N_28034,N_29503);
nor UO_2340 (O_2340,N_28601,N_28881);
nor UO_2341 (O_2341,N_29600,N_27313);
xor UO_2342 (O_2342,N_28237,N_28761);
nand UO_2343 (O_2343,N_27321,N_27994);
nor UO_2344 (O_2344,N_28861,N_27275);
nor UO_2345 (O_2345,N_27059,N_28704);
nand UO_2346 (O_2346,N_27118,N_27513);
or UO_2347 (O_2347,N_27448,N_29640);
xor UO_2348 (O_2348,N_29906,N_28154);
nand UO_2349 (O_2349,N_29080,N_27590);
nor UO_2350 (O_2350,N_27099,N_28798);
nor UO_2351 (O_2351,N_27131,N_29318);
or UO_2352 (O_2352,N_29667,N_28265);
and UO_2353 (O_2353,N_29357,N_29676);
xnor UO_2354 (O_2354,N_29150,N_29335);
and UO_2355 (O_2355,N_29529,N_27535);
nor UO_2356 (O_2356,N_29339,N_28088);
and UO_2357 (O_2357,N_29455,N_27281);
nor UO_2358 (O_2358,N_27413,N_29328);
nor UO_2359 (O_2359,N_27463,N_28581);
or UO_2360 (O_2360,N_28764,N_29484);
or UO_2361 (O_2361,N_27391,N_29962);
nor UO_2362 (O_2362,N_27351,N_28316);
or UO_2363 (O_2363,N_29292,N_29732);
nand UO_2364 (O_2364,N_27627,N_29492);
and UO_2365 (O_2365,N_28246,N_28806);
nand UO_2366 (O_2366,N_29144,N_28956);
and UO_2367 (O_2367,N_28369,N_27239);
or UO_2368 (O_2368,N_27578,N_28880);
and UO_2369 (O_2369,N_28769,N_29550);
and UO_2370 (O_2370,N_28642,N_29175);
nand UO_2371 (O_2371,N_28581,N_27983);
or UO_2372 (O_2372,N_27861,N_27960);
xor UO_2373 (O_2373,N_27551,N_28860);
and UO_2374 (O_2374,N_27058,N_27714);
and UO_2375 (O_2375,N_27754,N_28041);
nand UO_2376 (O_2376,N_29509,N_28977);
nor UO_2377 (O_2377,N_27221,N_27323);
nor UO_2378 (O_2378,N_29641,N_28983);
nor UO_2379 (O_2379,N_29553,N_27785);
and UO_2380 (O_2380,N_29385,N_28699);
xor UO_2381 (O_2381,N_28727,N_27303);
and UO_2382 (O_2382,N_29349,N_28464);
xor UO_2383 (O_2383,N_27234,N_28923);
nor UO_2384 (O_2384,N_27283,N_29471);
nor UO_2385 (O_2385,N_28514,N_27711);
and UO_2386 (O_2386,N_28240,N_29635);
or UO_2387 (O_2387,N_29133,N_27000);
nor UO_2388 (O_2388,N_28997,N_27101);
xor UO_2389 (O_2389,N_27107,N_29524);
and UO_2390 (O_2390,N_29722,N_28890);
nand UO_2391 (O_2391,N_27167,N_28224);
nand UO_2392 (O_2392,N_28134,N_28104);
nand UO_2393 (O_2393,N_29031,N_28528);
and UO_2394 (O_2394,N_28622,N_29019);
and UO_2395 (O_2395,N_28559,N_28520);
and UO_2396 (O_2396,N_27222,N_27630);
nor UO_2397 (O_2397,N_29984,N_28147);
nand UO_2398 (O_2398,N_28259,N_27056);
nand UO_2399 (O_2399,N_27248,N_27507);
and UO_2400 (O_2400,N_29664,N_28388);
and UO_2401 (O_2401,N_29185,N_28565);
xor UO_2402 (O_2402,N_28298,N_27235);
nand UO_2403 (O_2403,N_27463,N_27089);
and UO_2404 (O_2404,N_28855,N_27668);
nand UO_2405 (O_2405,N_28383,N_27501);
xor UO_2406 (O_2406,N_29866,N_28739);
nor UO_2407 (O_2407,N_27463,N_29700);
nor UO_2408 (O_2408,N_28994,N_29915);
nor UO_2409 (O_2409,N_28470,N_28747);
and UO_2410 (O_2410,N_29642,N_28923);
and UO_2411 (O_2411,N_29791,N_27092);
xnor UO_2412 (O_2412,N_27895,N_29699);
nor UO_2413 (O_2413,N_29367,N_29052);
and UO_2414 (O_2414,N_28995,N_29506);
nand UO_2415 (O_2415,N_29778,N_28991);
nand UO_2416 (O_2416,N_28833,N_29182);
xor UO_2417 (O_2417,N_28869,N_28753);
and UO_2418 (O_2418,N_27150,N_29187);
nor UO_2419 (O_2419,N_28077,N_29562);
nand UO_2420 (O_2420,N_29683,N_27334);
and UO_2421 (O_2421,N_28993,N_27808);
xnor UO_2422 (O_2422,N_27949,N_27963);
and UO_2423 (O_2423,N_28352,N_29045);
or UO_2424 (O_2424,N_27289,N_29595);
and UO_2425 (O_2425,N_27396,N_28342);
nand UO_2426 (O_2426,N_28563,N_29745);
or UO_2427 (O_2427,N_28734,N_27137);
xnor UO_2428 (O_2428,N_29276,N_27971);
nand UO_2429 (O_2429,N_29769,N_29409);
and UO_2430 (O_2430,N_29792,N_29397);
xnor UO_2431 (O_2431,N_27180,N_28626);
and UO_2432 (O_2432,N_29273,N_27081);
xor UO_2433 (O_2433,N_27652,N_28056);
or UO_2434 (O_2434,N_28287,N_29217);
nand UO_2435 (O_2435,N_29235,N_28981);
and UO_2436 (O_2436,N_29721,N_29563);
or UO_2437 (O_2437,N_28306,N_28366);
xnor UO_2438 (O_2438,N_27057,N_27627);
and UO_2439 (O_2439,N_27512,N_29466);
and UO_2440 (O_2440,N_28184,N_29214);
or UO_2441 (O_2441,N_27534,N_27417);
nand UO_2442 (O_2442,N_28480,N_27296);
nor UO_2443 (O_2443,N_28535,N_29296);
xnor UO_2444 (O_2444,N_29711,N_27020);
xnor UO_2445 (O_2445,N_29128,N_27460);
or UO_2446 (O_2446,N_27815,N_27775);
xor UO_2447 (O_2447,N_28796,N_29641);
and UO_2448 (O_2448,N_28273,N_29464);
xnor UO_2449 (O_2449,N_28147,N_29253);
and UO_2450 (O_2450,N_27423,N_28330);
xor UO_2451 (O_2451,N_27378,N_27219);
or UO_2452 (O_2452,N_28058,N_27508);
nor UO_2453 (O_2453,N_28063,N_27926);
nand UO_2454 (O_2454,N_28710,N_28680);
nand UO_2455 (O_2455,N_27620,N_27787);
or UO_2456 (O_2456,N_29195,N_29424);
nor UO_2457 (O_2457,N_28057,N_27522);
and UO_2458 (O_2458,N_27557,N_27895);
nand UO_2459 (O_2459,N_28835,N_29126);
or UO_2460 (O_2460,N_27118,N_28631);
nor UO_2461 (O_2461,N_27639,N_29459);
nand UO_2462 (O_2462,N_27361,N_29270);
xnor UO_2463 (O_2463,N_29794,N_27470);
and UO_2464 (O_2464,N_28409,N_27940);
or UO_2465 (O_2465,N_29680,N_28401);
nand UO_2466 (O_2466,N_28678,N_27273);
xor UO_2467 (O_2467,N_28774,N_28260);
or UO_2468 (O_2468,N_27376,N_27854);
nor UO_2469 (O_2469,N_29879,N_27966);
xor UO_2470 (O_2470,N_27315,N_29054);
xnor UO_2471 (O_2471,N_27294,N_27874);
xnor UO_2472 (O_2472,N_29509,N_28783);
or UO_2473 (O_2473,N_28384,N_29351);
or UO_2474 (O_2474,N_27148,N_27357);
nor UO_2475 (O_2475,N_28861,N_29186);
nand UO_2476 (O_2476,N_27395,N_27968);
and UO_2477 (O_2477,N_29523,N_28324);
nand UO_2478 (O_2478,N_28960,N_28832);
nand UO_2479 (O_2479,N_28672,N_29700);
nor UO_2480 (O_2480,N_28592,N_27649);
or UO_2481 (O_2481,N_28119,N_27804);
or UO_2482 (O_2482,N_29858,N_29853);
and UO_2483 (O_2483,N_29994,N_28721);
nand UO_2484 (O_2484,N_29911,N_28723);
and UO_2485 (O_2485,N_28158,N_28573);
or UO_2486 (O_2486,N_29294,N_28426);
or UO_2487 (O_2487,N_29061,N_28248);
and UO_2488 (O_2488,N_27425,N_27700);
xor UO_2489 (O_2489,N_27376,N_28314);
xor UO_2490 (O_2490,N_28202,N_29146);
nor UO_2491 (O_2491,N_29542,N_28314);
nand UO_2492 (O_2492,N_28460,N_28619);
and UO_2493 (O_2493,N_29701,N_29521);
and UO_2494 (O_2494,N_29955,N_29450);
or UO_2495 (O_2495,N_29924,N_28468);
nor UO_2496 (O_2496,N_27318,N_28644);
nor UO_2497 (O_2497,N_27672,N_29409);
or UO_2498 (O_2498,N_28289,N_27610);
xnor UO_2499 (O_2499,N_28123,N_29948);
nand UO_2500 (O_2500,N_28723,N_27551);
nand UO_2501 (O_2501,N_28791,N_28337);
or UO_2502 (O_2502,N_29020,N_28645);
nor UO_2503 (O_2503,N_29552,N_28186);
and UO_2504 (O_2504,N_28761,N_27429);
or UO_2505 (O_2505,N_29898,N_27273);
or UO_2506 (O_2506,N_29870,N_28990);
or UO_2507 (O_2507,N_28557,N_29031);
xor UO_2508 (O_2508,N_29293,N_28399);
xor UO_2509 (O_2509,N_27605,N_29200);
nand UO_2510 (O_2510,N_27005,N_28754);
nand UO_2511 (O_2511,N_29045,N_28458);
xor UO_2512 (O_2512,N_29052,N_28767);
nor UO_2513 (O_2513,N_28235,N_27081);
nor UO_2514 (O_2514,N_28655,N_29561);
xor UO_2515 (O_2515,N_29520,N_28261);
and UO_2516 (O_2516,N_29021,N_28373);
xor UO_2517 (O_2517,N_27440,N_29558);
nor UO_2518 (O_2518,N_28094,N_28522);
nor UO_2519 (O_2519,N_28478,N_28586);
and UO_2520 (O_2520,N_27830,N_27302);
xnor UO_2521 (O_2521,N_27265,N_29610);
and UO_2522 (O_2522,N_28201,N_29918);
xor UO_2523 (O_2523,N_29675,N_29760);
and UO_2524 (O_2524,N_28872,N_27028);
and UO_2525 (O_2525,N_28234,N_29768);
nor UO_2526 (O_2526,N_28258,N_27281);
and UO_2527 (O_2527,N_28946,N_27897);
nor UO_2528 (O_2528,N_29537,N_28810);
nor UO_2529 (O_2529,N_27727,N_29094);
nand UO_2530 (O_2530,N_28387,N_29316);
xnor UO_2531 (O_2531,N_27767,N_29939);
or UO_2532 (O_2532,N_28743,N_29429);
and UO_2533 (O_2533,N_27999,N_28003);
nor UO_2534 (O_2534,N_27565,N_27593);
and UO_2535 (O_2535,N_28923,N_27988);
and UO_2536 (O_2536,N_27710,N_29236);
nand UO_2537 (O_2537,N_27402,N_27686);
xnor UO_2538 (O_2538,N_28375,N_29332);
xor UO_2539 (O_2539,N_29256,N_28725);
nor UO_2540 (O_2540,N_28213,N_27738);
and UO_2541 (O_2541,N_28818,N_29963);
xor UO_2542 (O_2542,N_27520,N_28725);
nand UO_2543 (O_2543,N_27465,N_29355);
and UO_2544 (O_2544,N_27349,N_29967);
xor UO_2545 (O_2545,N_28749,N_29994);
xnor UO_2546 (O_2546,N_28632,N_29062);
and UO_2547 (O_2547,N_28909,N_29957);
nand UO_2548 (O_2548,N_27073,N_28504);
nand UO_2549 (O_2549,N_28244,N_28455);
nor UO_2550 (O_2550,N_27643,N_29909);
and UO_2551 (O_2551,N_29504,N_29378);
nand UO_2552 (O_2552,N_28316,N_28074);
xnor UO_2553 (O_2553,N_28236,N_28703);
nor UO_2554 (O_2554,N_28910,N_27695);
or UO_2555 (O_2555,N_29873,N_28448);
xor UO_2556 (O_2556,N_28021,N_29134);
nand UO_2557 (O_2557,N_29836,N_27380);
or UO_2558 (O_2558,N_29597,N_29674);
nor UO_2559 (O_2559,N_27559,N_28200);
nand UO_2560 (O_2560,N_27574,N_28005);
xnor UO_2561 (O_2561,N_28929,N_28788);
xor UO_2562 (O_2562,N_29469,N_29796);
or UO_2563 (O_2563,N_27459,N_28627);
or UO_2564 (O_2564,N_27785,N_27802);
nand UO_2565 (O_2565,N_28867,N_28251);
xnor UO_2566 (O_2566,N_28211,N_29532);
or UO_2567 (O_2567,N_28169,N_27287);
nand UO_2568 (O_2568,N_27093,N_27474);
and UO_2569 (O_2569,N_29742,N_27664);
or UO_2570 (O_2570,N_29260,N_29942);
xor UO_2571 (O_2571,N_29165,N_27488);
or UO_2572 (O_2572,N_29175,N_28283);
or UO_2573 (O_2573,N_29662,N_27504);
nor UO_2574 (O_2574,N_28201,N_27738);
nor UO_2575 (O_2575,N_29792,N_29263);
nand UO_2576 (O_2576,N_29411,N_28363);
or UO_2577 (O_2577,N_28491,N_29753);
nand UO_2578 (O_2578,N_29509,N_29472);
nor UO_2579 (O_2579,N_29192,N_27179);
or UO_2580 (O_2580,N_29313,N_28569);
nor UO_2581 (O_2581,N_27297,N_29379);
or UO_2582 (O_2582,N_27597,N_28047);
xnor UO_2583 (O_2583,N_27872,N_27171);
or UO_2584 (O_2584,N_27191,N_29902);
or UO_2585 (O_2585,N_28358,N_28612);
xor UO_2586 (O_2586,N_28119,N_27820);
or UO_2587 (O_2587,N_29799,N_28577);
and UO_2588 (O_2588,N_27086,N_28804);
and UO_2589 (O_2589,N_27142,N_28609);
xor UO_2590 (O_2590,N_29747,N_27710);
and UO_2591 (O_2591,N_28524,N_28369);
or UO_2592 (O_2592,N_28418,N_29671);
xnor UO_2593 (O_2593,N_29776,N_29277);
and UO_2594 (O_2594,N_29698,N_27318);
and UO_2595 (O_2595,N_27631,N_29459);
or UO_2596 (O_2596,N_27493,N_28759);
xor UO_2597 (O_2597,N_29560,N_28267);
and UO_2598 (O_2598,N_27814,N_27850);
xor UO_2599 (O_2599,N_28582,N_27873);
or UO_2600 (O_2600,N_27045,N_28618);
and UO_2601 (O_2601,N_28163,N_28550);
nand UO_2602 (O_2602,N_29148,N_28613);
and UO_2603 (O_2603,N_29303,N_29358);
nor UO_2604 (O_2604,N_27783,N_27273);
xor UO_2605 (O_2605,N_27945,N_28071);
nor UO_2606 (O_2606,N_29951,N_29754);
nand UO_2607 (O_2607,N_28322,N_27942);
or UO_2608 (O_2608,N_27158,N_28651);
and UO_2609 (O_2609,N_29145,N_27546);
nand UO_2610 (O_2610,N_29724,N_28144);
xor UO_2611 (O_2611,N_29221,N_28806);
xnor UO_2612 (O_2612,N_27460,N_27452);
xor UO_2613 (O_2613,N_27667,N_28616);
nand UO_2614 (O_2614,N_29972,N_27135);
nor UO_2615 (O_2615,N_28451,N_27178);
nand UO_2616 (O_2616,N_28149,N_27574);
and UO_2617 (O_2617,N_29319,N_27899);
xor UO_2618 (O_2618,N_29198,N_28503);
and UO_2619 (O_2619,N_27474,N_28318);
nand UO_2620 (O_2620,N_28821,N_28424);
and UO_2621 (O_2621,N_27221,N_27895);
or UO_2622 (O_2622,N_29193,N_28332);
nand UO_2623 (O_2623,N_29885,N_29108);
nand UO_2624 (O_2624,N_28776,N_27731);
xnor UO_2625 (O_2625,N_28963,N_28214);
and UO_2626 (O_2626,N_28016,N_29184);
or UO_2627 (O_2627,N_27225,N_28930);
nor UO_2628 (O_2628,N_28407,N_28957);
nand UO_2629 (O_2629,N_28703,N_28826);
and UO_2630 (O_2630,N_27570,N_27086);
or UO_2631 (O_2631,N_28307,N_28003);
nand UO_2632 (O_2632,N_28209,N_29710);
and UO_2633 (O_2633,N_29321,N_29019);
or UO_2634 (O_2634,N_28669,N_27628);
nand UO_2635 (O_2635,N_27771,N_29071);
nor UO_2636 (O_2636,N_27620,N_29841);
and UO_2637 (O_2637,N_28347,N_28230);
nor UO_2638 (O_2638,N_29779,N_28759);
and UO_2639 (O_2639,N_28448,N_29991);
and UO_2640 (O_2640,N_29564,N_29375);
xor UO_2641 (O_2641,N_28426,N_27321);
nor UO_2642 (O_2642,N_28579,N_27977);
nor UO_2643 (O_2643,N_27120,N_27670);
xnor UO_2644 (O_2644,N_28369,N_28715);
nor UO_2645 (O_2645,N_28139,N_27064);
or UO_2646 (O_2646,N_27084,N_28372);
nand UO_2647 (O_2647,N_27487,N_29311);
nand UO_2648 (O_2648,N_29449,N_27155);
or UO_2649 (O_2649,N_28610,N_28088);
or UO_2650 (O_2650,N_28895,N_28545);
and UO_2651 (O_2651,N_29632,N_27510);
nand UO_2652 (O_2652,N_27045,N_27813);
nand UO_2653 (O_2653,N_27417,N_27980);
nor UO_2654 (O_2654,N_27065,N_29150);
nor UO_2655 (O_2655,N_27676,N_29193);
nand UO_2656 (O_2656,N_28370,N_27579);
xnor UO_2657 (O_2657,N_28232,N_29584);
or UO_2658 (O_2658,N_29531,N_28329);
and UO_2659 (O_2659,N_29051,N_29477);
and UO_2660 (O_2660,N_27213,N_27894);
nand UO_2661 (O_2661,N_29359,N_29920);
and UO_2662 (O_2662,N_29679,N_29832);
and UO_2663 (O_2663,N_29950,N_29380);
nor UO_2664 (O_2664,N_29893,N_28892);
or UO_2665 (O_2665,N_27865,N_29660);
nand UO_2666 (O_2666,N_28969,N_29307);
xnor UO_2667 (O_2667,N_28467,N_28039);
xnor UO_2668 (O_2668,N_29052,N_29922);
nand UO_2669 (O_2669,N_28169,N_29476);
nand UO_2670 (O_2670,N_29503,N_29277);
xor UO_2671 (O_2671,N_29713,N_29240);
nand UO_2672 (O_2672,N_28065,N_27810);
or UO_2673 (O_2673,N_28033,N_29167);
or UO_2674 (O_2674,N_29912,N_27605);
nand UO_2675 (O_2675,N_27208,N_28094);
nor UO_2676 (O_2676,N_29640,N_28720);
xnor UO_2677 (O_2677,N_28672,N_27994);
nor UO_2678 (O_2678,N_29724,N_28094);
and UO_2679 (O_2679,N_29185,N_27623);
and UO_2680 (O_2680,N_29054,N_28718);
and UO_2681 (O_2681,N_27806,N_29138);
nor UO_2682 (O_2682,N_28803,N_29399);
xor UO_2683 (O_2683,N_28619,N_28988);
nand UO_2684 (O_2684,N_28099,N_29948);
nor UO_2685 (O_2685,N_28046,N_29728);
xor UO_2686 (O_2686,N_29518,N_27251);
xnor UO_2687 (O_2687,N_27996,N_28528);
and UO_2688 (O_2688,N_28183,N_28561);
nand UO_2689 (O_2689,N_27455,N_29810);
xnor UO_2690 (O_2690,N_27367,N_27558);
xnor UO_2691 (O_2691,N_29649,N_27536);
nor UO_2692 (O_2692,N_27982,N_27749);
nor UO_2693 (O_2693,N_28595,N_27643);
and UO_2694 (O_2694,N_28925,N_28952);
nand UO_2695 (O_2695,N_29778,N_28716);
xor UO_2696 (O_2696,N_29836,N_29563);
xor UO_2697 (O_2697,N_27635,N_27162);
nor UO_2698 (O_2698,N_29615,N_27831);
nand UO_2699 (O_2699,N_27459,N_29176);
or UO_2700 (O_2700,N_28672,N_28624);
xor UO_2701 (O_2701,N_29830,N_29618);
xor UO_2702 (O_2702,N_28610,N_27772);
and UO_2703 (O_2703,N_28533,N_27913);
nor UO_2704 (O_2704,N_29310,N_27390);
nor UO_2705 (O_2705,N_28114,N_29627);
xnor UO_2706 (O_2706,N_27761,N_27351);
nand UO_2707 (O_2707,N_27775,N_28036);
or UO_2708 (O_2708,N_27478,N_28721);
nor UO_2709 (O_2709,N_29031,N_29808);
xnor UO_2710 (O_2710,N_27528,N_28791);
and UO_2711 (O_2711,N_29463,N_28250);
or UO_2712 (O_2712,N_29979,N_27526);
xnor UO_2713 (O_2713,N_29180,N_29297);
nand UO_2714 (O_2714,N_28269,N_27082);
nor UO_2715 (O_2715,N_28427,N_27040);
or UO_2716 (O_2716,N_27923,N_29984);
xor UO_2717 (O_2717,N_29569,N_29542);
xor UO_2718 (O_2718,N_29377,N_28538);
xor UO_2719 (O_2719,N_28217,N_27241);
and UO_2720 (O_2720,N_27806,N_27682);
and UO_2721 (O_2721,N_27582,N_28196);
nand UO_2722 (O_2722,N_28450,N_28881);
or UO_2723 (O_2723,N_27353,N_28270);
nand UO_2724 (O_2724,N_27844,N_29764);
nand UO_2725 (O_2725,N_29346,N_29353);
or UO_2726 (O_2726,N_27248,N_29025);
nand UO_2727 (O_2727,N_29910,N_28969);
nor UO_2728 (O_2728,N_28368,N_29434);
or UO_2729 (O_2729,N_29263,N_29402);
nand UO_2730 (O_2730,N_27015,N_28155);
nor UO_2731 (O_2731,N_27550,N_29089);
and UO_2732 (O_2732,N_29769,N_29783);
or UO_2733 (O_2733,N_29296,N_27163);
nor UO_2734 (O_2734,N_29935,N_28681);
xor UO_2735 (O_2735,N_29512,N_27911);
or UO_2736 (O_2736,N_27397,N_27640);
nand UO_2737 (O_2737,N_28889,N_28381);
or UO_2738 (O_2738,N_28964,N_28912);
nor UO_2739 (O_2739,N_28632,N_28093);
nor UO_2740 (O_2740,N_28349,N_28292);
xnor UO_2741 (O_2741,N_27258,N_29100);
nor UO_2742 (O_2742,N_28649,N_28527);
or UO_2743 (O_2743,N_29481,N_27185);
xnor UO_2744 (O_2744,N_28638,N_29166);
xor UO_2745 (O_2745,N_27004,N_28235);
and UO_2746 (O_2746,N_29180,N_28204);
and UO_2747 (O_2747,N_29669,N_29832);
xnor UO_2748 (O_2748,N_28184,N_28564);
nor UO_2749 (O_2749,N_29309,N_29557);
xnor UO_2750 (O_2750,N_29705,N_27065);
xnor UO_2751 (O_2751,N_27805,N_28946);
nand UO_2752 (O_2752,N_28587,N_28767);
and UO_2753 (O_2753,N_29754,N_29737);
nand UO_2754 (O_2754,N_29814,N_27636);
nand UO_2755 (O_2755,N_27545,N_27979);
nand UO_2756 (O_2756,N_28661,N_27900);
nor UO_2757 (O_2757,N_28820,N_28511);
and UO_2758 (O_2758,N_29351,N_29451);
xor UO_2759 (O_2759,N_27815,N_29911);
xnor UO_2760 (O_2760,N_27631,N_29543);
nor UO_2761 (O_2761,N_29752,N_27879);
or UO_2762 (O_2762,N_28953,N_27001);
and UO_2763 (O_2763,N_27674,N_28170);
nand UO_2764 (O_2764,N_29009,N_28356);
nor UO_2765 (O_2765,N_28950,N_28935);
nor UO_2766 (O_2766,N_27171,N_28840);
and UO_2767 (O_2767,N_28916,N_28408);
nand UO_2768 (O_2768,N_29974,N_27599);
nand UO_2769 (O_2769,N_29237,N_27741);
and UO_2770 (O_2770,N_28520,N_27751);
and UO_2771 (O_2771,N_29027,N_29488);
and UO_2772 (O_2772,N_29629,N_29508);
nand UO_2773 (O_2773,N_27596,N_29807);
nor UO_2774 (O_2774,N_28743,N_27891);
or UO_2775 (O_2775,N_27089,N_29312);
xnor UO_2776 (O_2776,N_27210,N_27295);
and UO_2777 (O_2777,N_29791,N_27757);
nor UO_2778 (O_2778,N_29076,N_27305);
nor UO_2779 (O_2779,N_29674,N_29226);
or UO_2780 (O_2780,N_28316,N_27483);
nand UO_2781 (O_2781,N_27295,N_29701);
xnor UO_2782 (O_2782,N_29299,N_28604);
or UO_2783 (O_2783,N_28073,N_27025);
and UO_2784 (O_2784,N_29449,N_27976);
nor UO_2785 (O_2785,N_27526,N_27972);
nor UO_2786 (O_2786,N_27778,N_28663);
xnor UO_2787 (O_2787,N_28052,N_29018);
nand UO_2788 (O_2788,N_27951,N_29230);
nand UO_2789 (O_2789,N_29668,N_28489);
nor UO_2790 (O_2790,N_28519,N_27714);
and UO_2791 (O_2791,N_29560,N_28832);
and UO_2792 (O_2792,N_28234,N_29371);
and UO_2793 (O_2793,N_27883,N_29907);
or UO_2794 (O_2794,N_29599,N_28869);
nand UO_2795 (O_2795,N_27980,N_28695);
nand UO_2796 (O_2796,N_29235,N_27840);
or UO_2797 (O_2797,N_27978,N_27438);
or UO_2798 (O_2798,N_27707,N_29186);
or UO_2799 (O_2799,N_28416,N_28161);
nor UO_2800 (O_2800,N_29836,N_27952);
or UO_2801 (O_2801,N_27838,N_29802);
xor UO_2802 (O_2802,N_28400,N_28081);
nor UO_2803 (O_2803,N_27795,N_29494);
and UO_2804 (O_2804,N_27827,N_28783);
and UO_2805 (O_2805,N_28439,N_28382);
and UO_2806 (O_2806,N_29755,N_29383);
or UO_2807 (O_2807,N_27477,N_29763);
xnor UO_2808 (O_2808,N_28700,N_29264);
xor UO_2809 (O_2809,N_27250,N_27043);
nor UO_2810 (O_2810,N_27338,N_28806);
nand UO_2811 (O_2811,N_28393,N_28776);
xor UO_2812 (O_2812,N_29814,N_29284);
nor UO_2813 (O_2813,N_27602,N_29244);
or UO_2814 (O_2814,N_27944,N_29493);
or UO_2815 (O_2815,N_27166,N_28958);
and UO_2816 (O_2816,N_28864,N_28008);
nand UO_2817 (O_2817,N_28314,N_27955);
nand UO_2818 (O_2818,N_28196,N_29046);
nor UO_2819 (O_2819,N_27033,N_28074);
and UO_2820 (O_2820,N_27276,N_28606);
nor UO_2821 (O_2821,N_28485,N_29316);
and UO_2822 (O_2822,N_29251,N_29904);
nand UO_2823 (O_2823,N_29620,N_29703);
xor UO_2824 (O_2824,N_27157,N_27486);
or UO_2825 (O_2825,N_28344,N_29331);
xor UO_2826 (O_2826,N_29001,N_28169);
nor UO_2827 (O_2827,N_28605,N_27516);
or UO_2828 (O_2828,N_29682,N_29195);
or UO_2829 (O_2829,N_29345,N_29374);
and UO_2830 (O_2830,N_29389,N_29224);
nand UO_2831 (O_2831,N_28538,N_29376);
nand UO_2832 (O_2832,N_28680,N_29559);
xnor UO_2833 (O_2833,N_28876,N_29081);
nor UO_2834 (O_2834,N_27553,N_27293);
nand UO_2835 (O_2835,N_27319,N_29197);
nor UO_2836 (O_2836,N_29236,N_27938);
nor UO_2837 (O_2837,N_29544,N_28053);
and UO_2838 (O_2838,N_28574,N_29136);
and UO_2839 (O_2839,N_28220,N_28887);
xor UO_2840 (O_2840,N_28313,N_28719);
xnor UO_2841 (O_2841,N_27610,N_27242);
or UO_2842 (O_2842,N_27366,N_27125);
nor UO_2843 (O_2843,N_29136,N_28847);
and UO_2844 (O_2844,N_27630,N_27688);
xor UO_2845 (O_2845,N_27619,N_29599);
or UO_2846 (O_2846,N_28903,N_29333);
xnor UO_2847 (O_2847,N_28511,N_27818);
xnor UO_2848 (O_2848,N_27046,N_28934);
nand UO_2849 (O_2849,N_29567,N_28801);
nor UO_2850 (O_2850,N_29603,N_28598);
and UO_2851 (O_2851,N_29282,N_29991);
and UO_2852 (O_2852,N_29710,N_29013);
nand UO_2853 (O_2853,N_28607,N_28230);
nand UO_2854 (O_2854,N_29158,N_28214);
nor UO_2855 (O_2855,N_27369,N_29182);
nor UO_2856 (O_2856,N_28467,N_27112);
xor UO_2857 (O_2857,N_27222,N_28519);
xor UO_2858 (O_2858,N_29330,N_28729);
or UO_2859 (O_2859,N_29599,N_27478);
xor UO_2860 (O_2860,N_27813,N_28639);
or UO_2861 (O_2861,N_27031,N_27947);
and UO_2862 (O_2862,N_27056,N_27304);
nand UO_2863 (O_2863,N_29288,N_29106);
nor UO_2864 (O_2864,N_29365,N_28459);
xnor UO_2865 (O_2865,N_29619,N_28621);
nand UO_2866 (O_2866,N_27797,N_27323);
nand UO_2867 (O_2867,N_28482,N_29879);
and UO_2868 (O_2868,N_27317,N_29113);
or UO_2869 (O_2869,N_28610,N_28762);
xnor UO_2870 (O_2870,N_28879,N_28155);
nor UO_2871 (O_2871,N_27699,N_29275);
and UO_2872 (O_2872,N_28518,N_28151);
nor UO_2873 (O_2873,N_27266,N_29210);
nor UO_2874 (O_2874,N_27325,N_28057);
xnor UO_2875 (O_2875,N_27333,N_29368);
nand UO_2876 (O_2876,N_28182,N_28126);
nor UO_2877 (O_2877,N_28605,N_29584);
and UO_2878 (O_2878,N_27603,N_28897);
or UO_2879 (O_2879,N_29562,N_28676);
or UO_2880 (O_2880,N_29504,N_27616);
nor UO_2881 (O_2881,N_27793,N_29393);
and UO_2882 (O_2882,N_29949,N_29145);
xor UO_2883 (O_2883,N_29645,N_28454);
or UO_2884 (O_2884,N_27007,N_27634);
or UO_2885 (O_2885,N_29027,N_28457);
and UO_2886 (O_2886,N_29054,N_28787);
nor UO_2887 (O_2887,N_27062,N_27652);
nor UO_2888 (O_2888,N_29780,N_27463);
xor UO_2889 (O_2889,N_29075,N_28640);
xor UO_2890 (O_2890,N_27590,N_29563);
or UO_2891 (O_2891,N_28720,N_28501);
nand UO_2892 (O_2892,N_27680,N_28047);
or UO_2893 (O_2893,N_28334,N_28310);
or UO_2894 (O_2894,N_29495,N_28104);
nor UO_2895 (O_2895,N_28124,N_29593);
and UO_2896 (O_2896,N_27070,N_27258);
and UO_2897 (O_2897,N_29783,N_29997);
or UO_2898 (O_2898,N_28939,N_28452);
and UO_2899 (O_2899,N_27914,N_29577);
and UO_2900 (O_2900,N_28041,N_29006);
nor UO_2901 (O_2901,N_27460,N_27793);
and UO_2902 (O_2902,N_27783,N_27706);
nor UO_2903 (O_2903,N_27144,N_27080);
nand UO_2904 (O_2904,N_28628,N_29669);
xor UO_2905 (O_2905,N_29802,N_28698);
xor UO_2906 (O_2906,N_28546,N_29855);
xor UO_2907 (O_2907,N_29239,N_29857);
or UO_2908 (O_2908,N_27978,N_27685);
xnor UO_2909 (O_2909,N_29403,N_28192);
xor UO_2910 (O_2910,N_28543,N_27082);
and UO_2911 (O_2911,N_28841,N_29819);
nor UO_2912 (O_2912,N_27272,N_29155);
or UO_2913 (O_2913,N_28288,N_29112);
nand UO_2914 (O_2914,N_29763,N_28991);
nand UO_2915 (O_2915,N_27991,N_29165);
xor UO_2916 (O_2916,N_29414,N_28578);
nand UO_2917 (O_2917,N_29361,N_28864);
nand UO_2918 (O_2918,N_29567,N_27405);
nand UO_2919 (O_2919,N_27276,N_29630);
nor UO_2920 (O_2920,N_29584,N_27542);
and UO_2921 (O_2921,N_29351,N_28869);
and UO_2922 (O_2922,N_28118,N_27731);
nand UO_2923 (O_2923,N_27922,N_28346);
and UO_2924 (O_2924,N_29515,N_28944);
nand UO_2925 (O_2925,N_28767,N_27090);
nor UO_2926 (O_2926,N_29308,N_28997);
xnor UO_2927 (O_2927,N_27675,N_29945);
and UO_2928 (O_2928,N_29655,N_27444);
xnor UO_2929 (O_2929,N_29565,N_27337);
and UO_2930 (O_2930,N_27385,N_29903);
nand UO_2931 (O_2931,N_27028,N_29178);
nor UO_2932 (O_2932,N_28441,N_28678);
nor UO_2933 (O_2933,N_29984,N_29263);
or UO_2934 (O_2934,N_29100,N_28474);
and UO_2935 (O_2935,N_29745,N_28040);
xnor UO_2936 (O_2936,N_27577,N_27949);
and UO_2937 (O_2937,N_27867,N_29772);
nor UO_2938 (O_2938,N_28659,N_29412);
xor UO_2939 (O_2939,N_29553,N_27548);
and UO_2940 (O_2940,N_28441,N_27776);
or UO_2941 (O_2941,N_28552,N_28793);
nand UO_2942 (O_2942,N_28430,N_27007);
xor UO_2943 (O_2943,N_29082,N_28868);
xor UO_2944 (O_2944,N_28139,N_29821);
xnor UO_2945 (O_2945,N_27579,N_29225);
or UO_2946 (O_2946,N_29380,N_28821);
nor UO_2947 (O_2947,N_28589,N_28798);
nor UO_2948 (O_2948,N_27096,N_28716);
or UO_2949 (O_2949,N_29239,N_27148);
nor UO_2950 (O_2950,N_27023,N_29030);
xor UO_2951 (O_2951,N_28520,N_28954);
and UO_2952 (O_2952,N_28914,N_29375);
xor UO_2953 (O_2953,N_27049,N_29340);
nand UO_2954 (O_2954,N_28101,N_28678);
xnor UO_2955 (O_2955,N_28740,N_29791);
nor UO_2956 (O_2956,N_29326,N_29277);
or UO_2957 (O_2957,N_27638,N_29299);
and UO_2958 (O_2958,N_28213,N_28178);
nor UO_2959 (O_2959,N_27948,N_28742);
or UO_2960 (O_2960,N_29862,N_27600);
xnor UO_2961 (O_2961,N_29414,N_29176);
nor UO_2962 (O_2962,N_27495,N_29260);
nor UO_2963 (O_2963,N_28119,N_28220);
xor UO_2964 (O_2964,N_29091,N_27206);
nand UO_2965 (O_2965,N_29057,N_28631);
and UO_2966 (O_2966,N_29165,N_29105);
and UO_2967 (O_2967,N_27725,N_28044);
or UO_2968 (O_2968,N_28833,N_27547);
nor UO_2969 (O_2969,N_29262,N_29434);
nand UO_2970 (O_2970,N_28534,N_27811);
or UO_2971 (O_2971,N_27658,N_29320);
nor UO_2972 (O_2972,N_27210,N_27865);
nand UO_2973 (O_2973,N_29379,N_27396);
xnor UO_2974 (O_2974,N_28326,N_29533);
or UO_2975 (O_2975,N_29533,N_29896);
nand UO_2976 (O_2976,N_27299,N_27110);
nand UO_2977 (O_2977,N_29607,N_29991);
or UO_2978 (O_2978,N_27918,N_28991);
nand UO_2979 (O_2979,N_29585,N_29293);
nand UO_2980 (O_2980,N_28894,N_29999);
and UO_2981 (O_2981,N_29277,N_29721);
or UO_2982 (O_2982,N_27312,N_27211);
nand UO_2983 (O_2983,N_29150,N_27085);
nor UO_2984 (O_2984,N_27415,N_28595);
and UO_2985 (O_2985,N_28167,N_28211);
nor UO_2986 (O_2986,N_27233,N_29926);
or UO_2987 (O_2987,N_27507,N_28597);
or UO_2988 (O_2988,N_29752,N_27062);
or UO_2989 (O_2989,N_27232,N_29585);
and UO_2990 (O_2990,N_29675,N_29191);
or UO_2991 (O_2991,N_28228,N_29604);
xnor UO_2992 (O_2992,N_29471,N_28678);
xnor UO_2993 (O_2993,N_29937,N_29070);
or UO_2994 (O_2994,N_29334,N_27802);
nand UO_2995 (O_2995,N_29636,N_29464);
or UO_2996 (O_2996,N_28578,N_27416);
and UO_2997 (O_2997,N_27786,N_29461);
or UO_2998 (O_2998,N_28283,N_27824);
nor UO_2999 (O_2999,N_29679,N_27050);
and UO_3000 (O_3000,N_27859,N_28510);
nor UO_3001 (O_3001,N_27617,N_29330);
or UO_3002 (O_3002,N_28781,N_29540);
nor UO_3003 (O_3003,N_29357,N_28873);
xnor UO_3004 (O_3004,N_29398,N_28094);
nor UO_3005 (O_3005,N_27160,N_29710);
or UO_3006 (O_3006,N_28749,N_27784);
nand UO_3007 (O_3007,N_28939,N_28983);
xor UO_3008 (O_3008,N_29013,N_29874);
or UO_3009 (O_3009,N_28479,N_29292);
and UO_3010 (O_3010,N_28833,N_29043);
and UO_3011 (O_3011,N_28181,N_28604);
nor UO_3012 (O_3012,N_28665,N_28458);
nand UO_3013 (O_3013,N_29881,N_28182);
nor UO_3014 (O_3014,N_28846,N_29074);
xnor UO_3015 (O_3015,N_28844,N_28518);
and UO_3016 (O_3016,N_29246,N_27675);
nor UO_3017 (O_3017,N_28992,N_29154);
nand UO_3018 (O_3018,N_29625,N_27034);
and UO_3019 (O_3019,N_29399,N_27812);
nor UO_3020 (O_3020,N_29982,N_28477);
nand UO_3021 (O_3021,N_29459,N_27698);
nand UO_3022 (O_3022,N_29189,N_27412);
nor UO_3023 (O_3023,N_28594,N_27792);
nand UO_3024 (O_3024,N_29443,N_28869);
or UO_3025 (O_3025,N_28611,N_27646);
and UO_3026 (O_3026,N_29853,N_28118);
nor UO_3027 (O_3027,N_29043,N_28459);
or UO_3028 (O_3028,N_29960,N_27373);
nand UO_3029 (O_3029,N_29364,N_29385);
xnor UO_3030 (O_3030,N_29475,N_28945);
or UO_3031 (O_3031,N_28897,N_28534);
nor UO_3032 (O_3032,N_27325,N_28626);
or UO_3033 (O_3033,N_29391,N_28746);
nor UO_3034 (O_3034,N_27543,N_29767);
nand UO_3035 (O_3035,N_29401,N_27932);
and UO_3036 (O_3036,N_27177,N_27532);
nor UO_3037 (O_3037,N_28507,N_28026);
and UO_3038 (O_3038,N_28864,N_27579);
nand UO_3039 (O_3039,N_27525,N_29041);
or UO_3040 (O_3040,N_28452,N_28911);
xor UO_3041 (O_3041,N_27413,N_29873);
nor UO_3042 (O_3042,N_29267,N_28603);
and UO_3043 (O_3043,N_29818,N_27188);
nor UO_3044 (O_3044,N_28800,N_28494);
nor UO_3045 (O_3045,N_28699,N_29281);
or UO_3046 (O_3046,N_27683,N_28177);
and UO_3047 (O_3047,N_28355,N_27121);
and UO_3048 (O_3048,N_29177,N_27519);
or UO_3049 (O_3049,N_29707,N_28184);
and UO_3050 (O_3050,N_29429,N_29484);
nand UO_3051 (O_3051,N_29014,N_28024);
nand UO_3052 (O_3052,N_27638,N_29010);
nor UO_3053 (O_3053,N_29148,N_29539);
nor UO_3054 (O_3054,N_29697,N_27719);
nand UO_3055 (O_3055,N_29338,N_28654);
nor UO_3056 (O_3056,N_28927,N_28014);
xor UO_3057 (O_3057,N_27328,N_27763);
nor UO_3058 (O_3058,N_29392,N_28824);
nor UO_3059 (O_3059,N_28356,N_29613);
nor UO_3060 (O_3060,N_29811,N_27791);
nor UO_3061 (O_3061,N_27368,N_29629);
or UO_3062 (O_3062,N_28079,N_28667);
nand UO_3063 (O_3063,N_27386,N_28017);
and UO_3064 (O_3064,N_27456,N_27957);
nor UO_3065 (O_3065,N_27544,N_29107);
and UO_3066 (O_3066,N_27758,N_28033);
nor UO_3067 (O_3067,N_29436,N_28883);
nor UO_3068 (O_3068,N_29936,N_29767);
nor UO_3069 (O_3069,N_28548,N_29103);
and UO_3070 (O_3070,N_27926,N_29795);
nor UO_3071 (O_3071,N_29601,N_27787);
nor UO_3072 (O_3072,N_29407,N_27079);
and UO_3073 (O_3073,N_28246,N_29530);
xor UO_3074 (O_3074,N_29119,N_28118);
nor UO_3075 (O_3075,N_28475,N_29399);
nand UO_3076 (O_3076,N_27231,N_27663);
xor UO_3077 (O_3077,N_27120,N_27469);
nand UO_3078 (O_3078,N_28722,N_27625);
and UO_3079 (O_3079,N_29962,N_28840);
xnor UO_3080 (O_3080,N_28130,N_28098);
xnor UO_3081 (O_3081,N_29597,N_28166);
xnor UO_3082 (O_3082,N_28365,N_28350);
xnor UO_3083 (O_3083,N_29918,N_29696);
and UO_3084 (O_3084,N_27174,N_29277);
xnor UO_3085 (O_3085,N_29339,N_28034);
nor UO_3086 (O_3086,N_27085,N_28228);
nand UO_3087 (O_3087,N_27176,N_27695);
nor UO_3088 (O_3088,N_28154,N_28800);
xor UO_3089 (O_3089,N_27515,N_27232);
or UO_3090 (O_3090,N_29567,N_28425);
xor UO_3091 (O_3091,N_29670,N_29441);
nor UO_3092 (O_3092,N_29334,N_27951);
xor UO_3093 (O_3093,N_27150,N_28144);
nor UO_3094 (O_3094,N_29186,N_28071);
nor UO_3095 (O_3095,N_27524,N_27288);
nand UO_3096 (O_3096,N_27482,N_27203);
and UO_3097 (O_3097,N_28081,N_27229);
and UO_3098 (O_3098,N_27272,N_28021);
nor UO_3099 (O_3099,N_28229,N_28924);
and UO_3100 (O_3100,N_29469,N_28289);
and UO_3101 (O_3101,N_28481,N_28445);
and UO_3102 (O_3102,N_27054,N_29291);
xnor UO_3103 (O_3103,N_29479,N_27189);
nor UO_3104 (O_3104,N_27199,N_27708);
or UO_3105 (O_3105,N_28795,N_28756);
or UO_3106 (O_3106,N_27431,N_29014);
and UO_3107 (O_3107,N_29377,N_28473);
xor UO_3108 (O_3108,N_29832,N_27213);
or UO_3109 (O_3109,N_29038,N_28549);
or UO_3110 (O_3110,N_29331,N_29535);
and UO_3111 (O_3111,N_28192,N_27979);
or UO_3112 (O_3112,N_28416,N_28926);
xnor UO_3113 (O_3113,N_27681,N_27666);
xor UO_3114 (O_3114,N_29936,N_29321);
xor UO_3115 (O_3115,N_29231,N_29138);
nor UO_3116 (O_3116,N_27649,N_27132);
xor UO_3117 (O_3117,N_29607,N_29236);
nor UO_3118 (O_3118,N_27850,N_28929);
nand UO_3119 (O_3119,N_28080,N_29073);
nor UO_3120 (O_3120,N_28308,N_29902);
or UO_3121 (O_3121,N_27519,N_29899);
nor UO_3122 (O_3122,N_29000,N_27811);
nand UO_3123 (O_3123,N_27108,N_29052);
xor UO_3124 (O_3124,N_27133,N_29525);
nand UO_3125 (O_3125,N_27201,N_28922);
and UO_3126 (O_3126,N_28976,N_29384);
and UO_3127 (O_3127,N_29699,N_29729);
nor UO_3128 (O_3128,N_27436,N_29574);
xnor UO_3129 (O_3129,N_29708,N_27715);
nand UO_3130 (O_3130,N_29059,N_28745);
nand UO_3131 (O_3131,N_29553,N_28281);
or UO_3132 (O_3132,N_27086,N_27383);
nor UO_3133 (O_3133,N_27329,N_27984);
xnor UO_3134 (O_3134,N_29578,N_28277);
or UO_3135 (O_3135,N_27904,N_27103);
or UO_3136 (O_3136,N_29938,N_29822);
nor UO_3137 (O_3137,N_27156,N_28301);
or UO_3138 (O_3138,N_27342,N_29247);
xnor UO_3139 (O_3139,N_28137,N_27485);
and UO_3140 (O_3140,N_28154,N_29566);
nand UO_3141 (O_3141,N_29343,N_27990);
and UO_3142 (O_3142,N_28084,N_29203);
nor UO_3143 (O_3143,N_27061,N_27269);
or UO_3144 (O_3144,N_29058,N_27463);
and UO_3145 (O_3145,N_29892,N_27616);
and UO_3146 (O_3146,N_28539,N_27014);
or UO_3147 (O_3147,N_29562,N_29234);
or UO_3148 (O_3148,N_29309,N_28056);
or UO_3149 (O_3149,N_27000,N_29751);
nand UO_3150 (O_3150,N_28913,N_29750);
nand UO_3151 (O_3151,N_28673,N_27122);
xnor UO_3152 (O_3152,N_28270,N_27672);
and UO_3153 (O_3153,N_29574,N_27295);
xnor UO_3154 (O_3154,N_27465,N_29405);
or UO_3155 (O_3155,N_27645,N_28808);
nand UO_3156 (O_3156,N_28604,N_27582);
nor UO_3157 (O_3157,N_29791,N_29650);
or UO_3158 (O_3158,N_27132,N_29528);
and UO_3159 (O_3159,N_28241,N_27229);
nand UO_3160 (O_3160,N_27699,N_27051);
nand UO_3161 (O_3161,N_29301,N_27995);
and UO_3162 (O_3162,N_27143,N_27205);
xnor UO_3163 (O_3163,N_27102,N_28698);
and UO_3164 (O_3164,N_27281,N_29495);
and UO_3165 (O_3165,N_28093,N_29849);
xnor UO_3166 (O_3166,N_28581,N_29997);
or UO_3167 (O_3167,N_28749,N_28190);
and UO_3168 (O_3168,N_28478,N_29035);
nand UO_3169 (O_3169,N_29524,N_29767);
xor UO_3170 (O_3170,N_28466,N_28000);
nand UO_3171 (O_3171,N_27674,N_29955);
xor UO_3172 (O_3172,N_29685,N_27643);
nand UO_3173 (O_3173,N_29808,N_28765);
and UO_3174 (O_3174,N_28165,N_29737);
nand UO_3175 (O_3175,N_27130,N_29260);
and UO_3176 (O_3176,N_28300,N_28012);
nor UO_3177 (O_3177,N_29130,N_27449);
or UO_3178 (O_3178,N_27467,N_27042);
xnor UO_3179 (O_3179,N_27814,N_29789);
xnor UO_3180 (O_3180,N_27427,N_28096);
nand UO_3181 (O_3181,N_27058,N_28565);
nand UO_3182 (O_3182,N_29862,N_28404);
or UO_3183 (O_3183,N_28894,N_28501);
nor UO_3184 (O_3184,N_28441,N_29973);
and UO_3185 (O_3185,N_28882,N_29176);
or UO_3186 (O_3186,N_29053,N_27769);
nand UO_3187 (O_3187,N_27926,N_29196);
nand UO_3188 (O_3188,N_28599,N_29011);
and UO_3189 (O_3189,N_28729,N_29345);
xnor UO_3190 (O_3190,N_28762,N_29658);
xor UO_3191 (O_3191,N_28465,N_28931);
nor UO_3192 (O_3192,N_28707,N_28838);
or UO_3193 (O_3193,N_27801,N_27740);
nand UO_3194 (O_3194,N_27004,N_28061);
nor UO_3195 (O_3195,N_29386,N_29954);
and UO_3196 (O_3196,N_29077,N_28583);
or UO_3197 (O_3197,N_28175,N_27856);
nand UO_3198 (O_3198,N_27480,N_29975);
nand UO_3199 (O_3199,N_27608,N_28774);
or UO_3200 (O_3200,N_29915,N_29499);
or UO_3201 (O_3201,N_27573,N_29508);
nand UO_3202 (O_3202,N_28458,N_27416);
xor UO_3203 (O_3203,N_28104,N_28813);
or UO_3204 (O_3204,N_27135,N_28891);
and UO_3205 (O_3205,N_27566,N_27423);
or UO_3206 (O_3206,N_27487,N_27922);
nor UO_3207 (O_3207,N_27419,N_29458);
or UO_3208 (O_3208,N_27613,N_28380);
or UO_3209 (O_3209,N_29899,N_28460);
nor UO_3210 (O_3210,N_29667,N_29950);
nor UO_3211 (O_3211,N_27628,N_28118);
or UO_3212 (O_3212,N_29107,N_27106);
and UO_3213 (O_3213,N_27082,N_27072);
or UO_3214 (O_3214,N_27154,N_28330);
nor UO_3215 (O_3215,N_28213,N_28169);
xor UO_3216 (O_3216,N_29745,N_29387);
nand UO_3217 (O_3217,N_29715,N_28092);
nor UO_3218 (O_3218,N_28213,N_28838);
and UO_3219 (O_3219,N_29425,N_28720);
and UO_3220 (O_3220,N_27844,N_29122);
and UO_3221 (O_3221,N_29366,N_28577);
nand UO_3222 (O_3222,N_28568,N_29734);
nor UO_3223 (O_3223,N_27242,N_28372);
or UO_3224 (O_3224,N_29328,N_27368);
nand UO_3225 (O_3225,N_29074,N_29584);
nor UO_3226 (O_3226,N_29789,N_29924);
nor UO_3227 (O_3227,N_27123,N_29229);
xor UO_3228 (O_3228,N_28088,N_28494);
nand UO_3229 (O_3229,N_28602,N_27630);
nor UO_3230 (O_3230,N_28803,N_28501);
xor UO_3231 (O_3231,N_29313,N_28963);
and UO_3232 (O_3232,N_28882,N_28323);
or UO_3233 (O_3233,N_27949,N_27622);
and UO_3234 (O_3234,N_29639,N_27527);
nor UO_3235 (O_3235,N_29184,N_28391);
nor UO_3236 (O_3236,N_27863,N_28478);
and UO_3237 (O_3237,N_28602,N_29880);
and UO_3238 (O_3238,N_28616,N_27342);
and UO_3239 (O_3239,N_28192,N_28690);
and UO_3240 (O_3240,N_27404,N_29605);
nand UO_3241 (O_3241,N_29478,N_29076);
nor UO_3242 (O_3242,N_29200,N_28729);
nand UO_3243 (O_3243,N_29759,N_27061);
xor UO_3244 (O_3244,N_29353,N_27333);
nand UO_3245 (O_3245,N_29846,N_29284);
or UO_3246 (O_3246,N_29358,N_28161);
and UO_3247 (O_3247,N_29143,N_29241);
and UO_3248 (O_3248,N_28936,N_28428);
xnor UO_3249 (O_3249,N_29577,N_29818);
nor UO_3250 (O_3250,N_27818,N_27167);
or UO_3251 (O_3251,N_27783,N_29180);
nand UO_3252 (O_3252,N_28753,N_27313);
and UO_3253 (O_3253,N_28304,N_27172);
xnor UO_3254 (O_3254,N_29490,N_27566);
nor UO_3255 (O_3255,N_27849,N_28866);
xnor UO_3256 (O_3256,N_28059,N_28278);
or UO_3257 (O_3257,N_28789,N_27159);
nand UO_3258 (O_3258,N_28779,N_27831);
nor UO_3259 (O_3259,N_27388,N_27712);
or UO_3260 (O_3260,N_28146,N_29012);
or UO_3261 (O_3261,N_28235,N_27910);
or UO_3262 (O_3262,N_27688,N_28432);
and UO_3263 (O_3263,N_28970,N_29419);
nor UO_3264 (O_3264,N_27880,N_28145);
and UO_3265 (O_3265,N_27354,N_29095);
nor UO_3266 (O_3266,N_28244,N_28067);
nand UO_3267 (O_3267,N_27558,N_28921);
or UO_3268 (O_3268,N_29901,N_29006);
nor UO_3269 (O_3269,N_27137,N_28646);
nand UO_3270 (O_3270,N_29198,N_28385);
or UO_3271 (O_3271,N_28524,N_27012);
xor UO_3272 (O_3272,N_28469,N_28238);
and UO_3273 (O_3273,N_29838,N_27344);
nand UO_3274 (O_3274,N_29778,N_27158);
nand UO_3275 (O_3275,N_27342,N_28316);
or UO_3276 (O_3276,N_27757,N_29606);
or UO_3277 (O_3277,N_28604,N_27984);
nand UO_3278 (O_3278,N_27198,N_29434);
and UO_3279 (O_3279,N_28189,N_27821);
xnor UO_3280 (O_3280,N_27696,N_28569);
nor UO_3281 (O_3281,N_28110,N_27982);
and UO_3282 (O_3282,N_28088,N_27143);
nand UO_3283 (O_3283,N_28992,N_27855);
or UO_3284 (O_3284,N_28699,N_28884);
xor UO_3285 (O_3285,N_28260,N_28489);
nand UO_3286 (O_3286,N_28284,N_27843);
nand UO_3287 (O_3287,N_29683,N_27441);
xor UO_3288 (O_3288,N_27060,N_29595);
xnor UO_3289 (O_3289,N_27057,N_28411);
nand UO_3290 (O_3290,N_27345,N_27488);
and UO_3291 (O_3291,N_29463,N_27844);
nor UO_3292 (O_3292,N_29122,N_28051);
or UO_3293 (O_3293,N_28144,N_28336);
and UO_3294 (O_3294,N_27514,N_28011);
and UO_3295 (O_3295,N_27025,N_27139);
xor UO_3296 (O_3296,N_28401,N_28720);
xnor UO_3297 (O_3297,N_28414,N_29500);
nand UO_3298 (O_3298,N_29085,N_28236);
and UO_3299 (O_3299,N_28830,N_27295);
xnor UO_3300 (O_3300,N_27189,N_29901);
or UO_3301 (O_3301,N_27900,N_28702);
nand UO_3302 (O_3302,N_28293,N_29543);
or UO_3303 (O_3303,N_29489,N_29351);
nor UO_3304 (O_3304,N_28152,N_27528);
and UO_3305 (O_3305,N_29482,N_27287);
and UO_3306 (O_3306,N_27255,N_28438);
nor UO_3307 (O_3307,N_28267,N_27275);
and UO_3308 (O_3308,N_29550,N_29735);
or UO_3309 (O_3309,N_29371,N_28183);
nand UO_3310 (O_3310,N_29962,N_29848);
xnor UO_3311 (O_3311,N_27818,N_28503);
nor UO_3312 (O_3312,N_28726,N_28055);
or UO_3313 (O_3313,N_27132,N_27768);
nor UO_3314 (O_3314,N_28802,N_28296);
xor UO_3315 (O_3315,N_29852,N_29604);
and UO_3316 (O_3316,N_28066,N_27752);
nor UO_3317 (O_3317,N_27521,N_27215);
and UO_3318 (O_3318,N_29941,N_27767);
nand UO_3319 (O_3319,N_27599,N_27724);
or UO_3320 (O_3320,N_27222,N_29093);
and UO_3321 (O_3321,N_27899,N_28562);
or UO_3322 (O_3322,N_28936,N_28459);
and UO_3323 (O_3323,N_28920,N_28302);
xnor UO_3324 (O_3324,N_29044,N_29078);
or UO_3325 (O_3325,N_28648,N_29615);
nand UO_3326 (O_3326,N_27638,N_29467);
nor UO_3327 (O_3327,N_28635,N_28583);
nand UO_3328 (O_3328,N_27907,N_27540);
nand UO_3329 (O_3329,N_28573,N_29214);
xor UO_3330 (O_3330,N_28447,N_27311);
nor UO_3331 (O_3331,N_27717,N_27738);
and UO_3332 (O_3332,N_28472,N_29085);
and UO_3333 (O_3333,N_29508,N_29383);
xnor UO_3334 (O_3334,N_28565,N_28955);
or UO_3335 (O_3335,N_29001,N_28980);
nor UO_3336 (O_3336,N_27084,N_27342);
nor UO_3337 (O_3337,N_28814,N_28104);
nand UO_3338 (O_3338,N_29724,N_29805);
xor UO_3339 (O_3339,N_28352,N_29070);
or UO_3340 (O_3340,N_28987,N_28501);
nor UO_3341 (O_3341,N_28192,N_28102);
nand UO_3342 (O_3342,N_29910,N_28182);
or UO_3343 (O_3343,N_29033,N_28469);
nand UO_3344 (O_3344,N_27015,N_28324);
nand UO_3345 (O_3345,N_29459,N_27164);
or UO_3346 (O_3346,N_28741,N_28173);
xor UO_3347 (O_3347,N_28378,N_28949);
and UO_3348 (O_3348,N_28652,N_28779);
nor UO_3349 (O_3349,N_29779,N_27060);
or UO_3350 (O_3350,N_29455,N_29085);
or UO_3351 (O_3351,N_28477,N_27514);
and UO_3352 (O_3352,N_28587,N_28089);
and UO_3353 (O_3353,N_29634,N_29696);
and UO_3354 (O_3354,N_29559,N_28064);
and UO_3355 (O_3355,N_29002,N_29580);
xnor UO_3356 (O_3356,N_29441,N_27085);
nor UO_3357 (O_3357,N_29219,N_29340);
nand UO_3358 (O_3358,N_28623,N_28608);
or UO_3359 (O_3359,N_27748,N_28001);
nor UO_3360 (O_3360,N_29913,N_27721);
nor UO_3361 (O_3361,N_27314,N_27797);
nand UO_3362 (O_3362,N_27917,N_28398);
nand UO_3363 (O_3363,N_29465,N_27275);
and UO_3364 (O_3364,N_27776,N_28032);
xor UO_3365 (O_3365,N_28031,N_29207);
nand UO_3366 (O_3366,N_28373,N_27972);
xor UO_3367 (O_3367,N_27460,N_28093);
nor UO_3368 (O_3368,N_29000,N_27791);
and UO_3369 (O_3369,N_28892,N_27048);
nand UO_3370 (O_3370,N_29440,N_28167);
and UO_3371 (O_3371,N_29869,N_29926);
nor UO_3372 (O_3372,N_29220,N_29184);
and UO_3373 (O_3373,N_27701,N_28538);
and UO_3374 (O_3374,N_29202,N_28999);
nand UO_3375 (O_3375,N_27639,N_29848);
and UO_3376 (O_3376,N_29619,N_27259);
nor UO_3377 (O_3377,N_28466,N_28067);
nor UO_3378 (O_3378,N_27043,N_27485);
nor UO_3379 (O_3379,N_29172,N_28417);
or UO_3380 (O_3380,N_27270,N_27120);
and UO_3381 (O_3381,N_29075,N_29972);
or UO_3382 (O_3382,N_28710,N_28191);
and UO_3383 (O_3383,N_29496,N_28327);
xor UO_3384 (O_3384,N_29509,N_27206);
and UO_3385 (O_3385,N_29040,N_27067);
and UO_3386 (O_3386,N_29022,N_27157);
or UO_3387 (O_3387,N_29792,N_29628);
xnor UO_3388 (O_3388,N_27193,N_29124);
xnor UO_3389 (O_3389,N_27221,N_27965);
and UO_3390 (O_3390,N_28628,N_29104);
nand UO_3391 (O_3391,N_27872,N_29766);
and UO_3392 (O_3392,N_28432,N_28250);
or UO_3393 (O_3393,N_27086,N_28170);
or UO_3394 (O_3394,N_28571,N_27292);
or UO_3395 (O_3395,N_28717,N_28221);
nand UO_3396 (O_3396,N_27049,N_29222);
xor UO_3397 (O_3397,N_28270,N_28884);
and UO_3398 (O_3398,N_27743,N_29847);
xor UO_3399 (O_3399,N_27211,N_29475);
nand UO_3400 (O_3400,N_28128,N_27642);
or UO_3401 (O_3401,N_27839,N_29272);
or UO_3402 (O_3402,N_29798,N_27272);
or UO_3403 (O_3403,N_29194,N_29163);
and UO_3404 (O_3404,N_28599,N_28988);
or UO_3405 (O_3405,N_29588,N_29225);
or UO_3406 (O_3406,N_29361,N_27696);
nand UO_3407 (O_3407,N_27247,N_28115);
nand UO_3408 (O_3408,N_27308,N_29890);
xor UO_3409 (O_3409,N_29424,N_29122);
or UO_3410 (O_3410,N_29481,N_28636);
nor UO_3411 (O_3411,N_28158,N_28623);
xnor UO_3412 (O_3412,N_28569,N_27393);
and UO_3413 (O_3413,N_29672,N_28685);
and UO_3414 (O_3414,N_28270,N_27094);
nand UO_3415 (O_3415,N_27498,N_27063);
xor UO_3416 (O_3416,N_27528,N_27483);
or UO_3417 (O_3417,N_29942,N_27897);
nand UO_3418 (O_3418,N_27548,N_28051);
and UO_3419 (O_3419,N_28901,N_27925);
or UO_3420 (O_3420,N_28685,N_28928);
xor UO_3421 (O_3421,N_27386,N_27523);
or UO_3422 (O_3422,N_28360,N_29200);
and UO_3423 (O_3423,N_28847,N_29829);
nand UO_3424 (O_3424,N_28717,N_28155);
and UO_3425 (O_3425,N_27929,N_27433);
or UO_3426 (O_3426,N_28012,N_28858);
nand UO_3427 (O_3427,N_29384,N_27480);
xor UO_3428 (O_3428,N_28122,N_28522);
or UO_3429 (O_3429,N_28868,N_27317);
nand UO_3430 (O_3430,N_29749,N_28182);
or UO_3431 (O_3431,N_29605,N_29791);
nor UO_3432 (O_3432,N_28883,N_28658);
or UO_3433 (O_3433,N_27575,N_27629);
nand UO_3434 (O_3434,N_29016,N_29879);
xor UO_3435 (O_3435,N_28612,N_28999);
and UO_3436 (O_3436,N_28819,N_28888);
nor UO_3437 (O_3437,N_28581,N_28133);
and UO_3438 (O_3438,N_28830,N_29056);
or UO_3439 (O_3439,N_27712,N_27756);
nor UO_3440 (O_3440,N_29034,N_29952);
xnor UO_3441 (O_3441,N_29186,N_27411);
nand UO_3442 (O_3442,N_29988,N_27876);
xnor UO_3443 (O_3443,N_28059,N_29080);
or UO_3444 (O_3444,N_29920,N_27527);
or UO_3445 (O_3445,N_29503,N_29971);
and UO_3446 (O_3446,N_29771,N_28195);
or UO_3447 (O_3447,N_27978,N_29979);
nand UO_3448 (O_3448,N_27163,N_29068);
nand UO_3449 (O_3449,N_28822,N_28159);
nand UO_3450 (O_3450,N_29625,N_28398);
nand UO_3451 (O_3451,N_27347,N_29502);
or UO_3452 (O_3452,N_27514,N_28144);
nand UO_3453 (O_3453,N_29142,N_29094);
nor UO_3454 (O_3454,N_27179,N_27318);
and UO_3455 (O_3455,N_29373,N_29897);
or UO_3456 (O_3456,N_29751,N_28781);
or UO_3457 (O_3457,N_27501,N_29040);
nand UO_3458 (O_3458,N_29394,N_28709);
nand UO_3459 (O_3459,N_27169,N_29984);
xnor UO_3460 (O_3460,N_27092,N_28677);
xor UO_3461 (O_3461,N_28554,N_28038);
and UO_3462 (O_3462,N_27198,N_29551);
and UO_3463 (O_3463,N_27247,N_29606);
or UO_3464 (O_3464,N_29769,N_29747);
and UO_3465 (O_3465,N_27045,N_28094);
nor UO_3466 (O_3466,N_28393,N_29100);
or UO_3467 (O_3467,N_28266,N_27090);
nor UO_3468 (O_3468,N_29380,N_29236);
and UO_3469 (O_3469,N_27091,N_27411);
and UO_3470 (O_3470,N_29314,N_29949);
or UO_3471 (O_3471,N_28637,N_27195);
or UO_3472 (O_3472,N_28991,N_27413);
or UO_3473 (O_3473,N_29244,N_27057);
nor UO_3474 (O_3474,N_28889,N_29389);
xnor UO_3475 (O_3475,N_27517,N_28429);
nor UO_3476 (O_3476,N_29628,N_28091);
nor UO_3477 (O_3477,N_28173,N_29610);
and UO_3478 (O_3478,N_27472,N_27245);
or UO_3479 (O_3479,N_29845,N_29076);
xor UO_3480 (O_3480,N_27195,N_29900);
nor UO_3481 (O_3481,N_28446,N_28845);
xnor UO_3482 (O_3482,N_29770,N_27073);
nand UO_3483 (O_3483,N_29042,N_27462);
and UO_3484 (O_3484,N_28881,N_27731);
and UO_3485 (O_3485,N_29235,N_28102);
xnor UO_3486 (O_3486,N_27902,N_28656);
xor UO_3487 (O_3487,N_29156,N_29476);
or UO_3488 (O_3488,N_28128,N_28916);
or UO_3489 (O_3489,N_27134,N_29757);
nand UO_3490 (O_3490,N_28235,N_27516);
or UO_3491 (O_3491,N_28975,N_29561);
xnor UO_3492 (O_3492,N_27540,N_29331);
and UO_3493 (O_3493,N_27077,N_28085);
nand UO_3494 (O_3494,N_27082,N_29649);
nor UO_3495 (O_3495,N_27111,N_28929);
nor UO_3496 (O_3496,N_28942,N_27525);
nor UO_3497 (O_3497,N_28480,N_29032);
xnor UO_3498 (O_3498,N_27329,N_28555);
nand UO_3499 (O_3499,N_29423,N_29759);
endmodule