module basic_500_3000_500_4_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_62,In_176);
nand U1 (N_1,In_14,In_377);
nand U2 (N_2,In_87,In_444);
nor U3 (N_3,In_303,In_250);
and U4 (N_4,In_362,In_197);
or U5 (N_5,In_421,In_224);
or U6 (N_6,In_50,In_277);
and U7 (N_7,In_108,In_376);
nand U8 (N_8,In_297,In_321);
or U9 (N_9,In_429,In_257);
and U10 (N_10,In_229,In_54);
nand U11 (N_11,In_179,In_398);
and U12 (N_12,In_139,In_409);
or U13 (N_13,In_221,In_56);
and U14 (N_14,In_353,In_157);
or U15 (N_15,In_281,In_283);
and U16 (N_16,In_324,In_51);
and U17 (N_17,In_130,In_100);
nand U18 (N_18,In_155,In_147);
or U19 (N_19,In_174,In_180);
and U20 (N_20,In_415,In_170);
xor U21 (N_21,In_269,In_165);
and U22 (N_22,In_472,In_134);
and U23 (N_23,In_191,In_378);
and U24 (N_24,In_138,In_320);
or U25 (N_25,In_309,In_55);
nand U26 (N_26,In_400,In_434);
and U27 (N_27,In_498,In_316);
nor U28 (N_28,In_133,In_368);
nand U29 (N_29,In_346,In_188);
nor U30 (N_30,In_22,In_9);
nand U31 (N_31,In_292,In_274);
and U32 (N_32,In_227,In_384);
and U33 (N_33,In_307,In_311);
nor U34 (N_34,In_351,In_245);
nand U35 (N_35,In_296,In_308);
and U36 (N_36,In_273,In_169);
nand U37 (N_37,In_423,In_266);
and U38 (N_38,In_21,In_26);
nand U39 (N_39,In_68,In_18);
nor U40 (N_40,In_150,In_440);
or U41 (N_41,In_488,In_31);
and U42 (N_42,In_225,In_228);
and U43 (N_43,In_360,In_294);
nor U44 (N_44,In_441,In_70);
or U45 (N_45,In_416,In_348);
or U46 (N_46,In_29,In_48);
nand U47 (N_47,In_23,In_182);
nor U48 (N_48,In_153,In_35);
and U49 (N_49,In_120,In_413);
and U50 (N_50,In_260,In_454);
nor U51 (N_51,In_63,In_226);
nor U52 (N_52,In_331,In_350);
nor U53 (N_53,In_287,In_30);
nor U54 (N_54,In_148,In_37);
or U55 (N_55,In_159,In_58);
or U56 (N_56,In_184,In_220);
and U57 (N_57,In_201,In_473);
and U58 (N_58,In_28,In_330);
or U59 (N_59,In_99,In_49);
xor U60 (N_60,In_397,In_447);
or U61 (N_61,In_73,In_91);
nand U62 (N_62,In_151,In_483);
or U63 (N_63,In_407,In_72);
xor U64 (N_64,In_465,In_450);
nand U65 (N_65,In_299,In_43);
nor U66 (N_66,In_301,In_264);
and U67 (N_67,In_75,In_164);
nor U68 (N_68,In_263,In_86);
nand U69 (N_69,In_90,In_34);
nor U70 (N_70,In_237,In_404);
or U71 (N_71,In_219,In_457);
nor U72 (N_72,In_115,In_71);
nor U73 (N_73,In_298,In_305);
nand U74 (N_74,In_253,In_238);
nor U75 (N_75,In_175,In_322);
or U76 (N_76,In_205,In_116);
nand U77 (N_77,In_342,In_374);
or U78 (N_78,In_209,In_215);
and U79 (N_79,In_442,In_189);
and U80 (N_80,In_93,In_13);
nand U81 (N_81,In_146,In_142);
and U82 (N_82,In_480,In_166);
or U83 (N_83,In_218,In_40);
nor U84 (N_84,In_102,In_438);
or U85 (N_85,In_111,In_363);
nand U86 (N_86,In_185,In_117);
nand U87 (N_87,In_388,In_211);
nor U88 (N_88,In_256,In_354);
and U89 (N_89,In_59,In_381);
nand U90 (N_90,In_328,In_453);
or U91 (N_91,In_19,In_163);
nor U92 (N_92,In_485,In_284);
or U93 (N_93,In_94,In_149);
and U94 (N_94,In_39,In_481);
nand U95 (N_95,In_333,In_95);
and U96 (N_96,In_132,In_206);
and U97 (N_97,In_462,In_231);
nor U98 (N_98,In_3,In_367);
or U99 (N_99,In_390,In_449);
xor U100 (N_100,In_372,In_302);
nor U101 (N_101,In_459,In_448);
or U102 (N_102,In_469,In_255);
nand U103 (N_103,In_208,In_207);
nand U104 (N_104,In_103,In_125);
and U105 (N_105,In_67,In_252);
nor U106 (N_106,In_495,In_338);
and U107 (N_107,In_349,In_172);
or U108 (N_108,In_491,In_233);
nor U109 (N_109,In_16,In_141);
nand U110 (N_110,In_66,In_411);
nand U111 (N_111,In_241,In_344);
nor U112 (N_112,In_2,In_386);
or U113 (N_113,In_8,In_382);
nand U114 (N_114,In_352,In_420);
or U115 (N_115,In_275,In_65);
nand U116 (N_116,In_332,In_119);
or U117 (N_117,In_489,In_437);
and U118 (N_118,In_186,In_410);
and U119 (N_119,In_97,In_78);
and U120 (N_120,In_128,In_80);
xor U121 (N_121,In_312,In_187);
or U122 (N_122,In_474,In_270);
or U123 (N_123,In_236,In_74);
nor U124 (N_124,In_127,In_10);
or U125 (N_125,In_109,In_276);
nor U126 (N_126,In_212,In_279);
or U127 (N_127,In_38,In_17);
nand U128 (N_128,In_11,In_494);
or U129 (N_129,In_20,In_261);
or U130 (N_130,In_248,In_383);
nand U131 (N_131,In_81,In_33);
and U132 (N_132,In_268,In_278);
or U133 (N_133,In_265,In_131);
nor U134 (N_134,In_259,In_183);
nand U135 (N_135,In_479,In_177);
or U136 (N_136,In_0,In_5);
or U137 (N_137,In_171,In_242);
nor U138 (N_138,In_484,In_295);
xor U139 (N_139,In_27,In_458);
or U140 (N_140,In_435,In_249);
nand U141 (N_141,In_232,In_345);
nor U142 (N_142,In_101,In_443);
and U143 (N_143,In_402,In_129);
nor U144 (N_144,In_124,In_327);
nor U145 (N_145,In_408,In_64);
nand U146 (N_146,In_347,In_247);
xnor U147 (N_147,In_464,In_106);
or U148 (N_148,In_452,In_79);
nand U149 (N_149,In_135,In_32);
nor U150 (N_150,In_366,In_190);
xnor U151 (N_151,In_57,In_395);
or U152 (N_152,In_375,In_272);
and U153 (N_153,In_379,In_285);
xnor U154 (N_154,In_267,In_325);
and U155 (N_155,In_422,In_282);
nand U156 (N_156,In_244,In_425);
and U157 (N_157,In_76,In_412);
nor U158 (N_158,In_478,In_405);
nor U159 (N_159,In_318,In_69);
nand U160 (N_160,In_200,In_82);
nor U161 (N_161,In_45,In_160);
nor U162 (N_162,In_192,In_85);
or U163 (N_163,In_162,In_329);
nand U164 (N_164,In_7,In_216);
nor U165 (N_165,In_104,In_313);
or U166 (N_166,In_280,In_36);
xor U167 (N_167,In_492,In_203);
and U168 (N_168,In_471,In_314);
or U169 (N_169,In_291,In_426);
and U170 (N_170,In_84,In_136);
or U171 (N_171,In_83,In_122);
nand U172 (N_172,In_306,In_288);
or U173 (N_173,In_53,In_92);
nand U174 (N_174,In_430,In_335);
or U175 (N_175,In_145,In_343);
and U176 (N_176,In_161,In_123);
or U177 (N_177,In_167,In_389);
nor U178 (N_178,In_392,In_373);
or U179 (N_179,In_475,In_364);
nand U180 (N_180,In_468,In_419);
nor U181 (N_181,In_369,In_198);
or U182 (N_182,In_451,In_436);
or U183 (N_183,In_406,In_262);
nand U184 (N_184,In_380,In_358);
nand U185 (N_185,In_467,In_42);
and U186 (N_186,In_476,In_194);
or U187 (N_187,In_359,In_477);
nand U188 (N_188,In_121,In_433);
and U189 (N_189,In_98,In_213);
or U190 (N_190,In_140,In_286);
or U191 (N_191,In_158,In_496);
or U192 (N_192,In_251,In_417);
nand U193 (N_193,In_156,In_424);
or U194 (N_194,In_12,In_137);
or U195 (N_195,In_455,In_47);
nand U196 (N_196,In_334,In_393);
nor U197 (N_197,In_4,In_210);
or U198 (N_198,In_154,In_52);
and U199 (N_199,In_6,In_493);
nor U200 (N_200,In_470,In_399);
or U201 (N_201,In_173,In_144);
or U202 (N_202,In_193,In_431);
nand U203 (N_203,In_25,In_371);
nor U204 (N_204,In_222,In_60);
nor U205 (N_205,In_497,In_460);
nor U206 (N_206,In_96,In_118);
or U207 (N_207,In_317,In_356);
nand U208 (N_208,In_394,In_112);
nand U209 (N_209,In_304,In_290);
or U210 (N_210,In_289,In_355);
and U211 (N_211,In_77,In_365);
and U212 (N_212,In_217,In_254);
or U213 (N_213,In_44,In_199);
and U214 (N_214,In_181,In_387);
xnor U215 (N_215,In_61,In_427);
nand U216 (N_216,In_499,In_46);
nor U217 (N_217,In_143,In_310);
and U218 (N_218,In_361,In_463);
nand U219 (N_219,In_403,In_337);
nor U220 (N_220,In_195,In_456);
or U221 (N_221,In_88,In_258);
nand U222 (N_222,In_239,In_341);
or U223 (N_223,In_243,In_246);
nand U224 (N_224,In_300,In_1);
or U225 (N_225,In_461,In_15);
nor U226 (N_226,In_105,In_336);
nor U227 (N_227,In_357,In_113);
nor U228 (N_228,In_487,In_24);
or U229 (N_229,In_152,In_271);
or U230 (N_230,In_223,In_126);
xor U231 (N_231,In_204,In_214);
nor U232 (N_232,In_89,In_319);
and U233 (N_233,In_41,In_293);
nor U234 (N_234,In_315,In_391);
or U235 (N_235,In_339,In_326);
xor U236 (N_236,In_486,In_178);
nand U237 (N_237,In_428,In_202);
or U238 (N_238,In_230,In_401);
and U239 (N_239,In_323,In_240);
nand U240 (N_240,In_235,In_482);
nor U241 (N_241,In_107,In_466);
xnor U242 (N_242,In_418,In_196);
and U243 (N_243,In_114,In_446);
nand U244 (N_244,In_490,In_432);
or U245 (N_245,In_340,In_439);
nand U246 (N_246,In_370,In_396);
nor U247 (N_247,In_414,In_385);
nor U248 (N_248,In_168,In_445);
nor U249 (N_249,In_110,In_234);
nand U250 (N_250,In_339,In_398);
nor U251 (N_251,In_410,In_31);
nand U252 (N_252,In_494,In_359);
or U253 (N_253,In_227,In_349);
nor U254 (N_254,In_244,In_489);
and U255 (N_255,In_280,In_89);
and U256 (N_256,In_471,In_468);
and U257 (N_257,In_436,In_282);
and U258 (N_258,In_235,In_398);
and U259 (N_259,In_280,In_204);
or U260 (N_260,In_185,In_275);
nand U261 (N_261,In_116,In_208);
and U262 (N_262,In_222,In_449);
or U263 (N_263,In_229,In_379);
nor U264 (N_264,In_276,In_480);
or U265 (N_265,In_496,In_181);
and U266 (N_266,In_484,In_430);
nand U267 (N_267,In_481,In_319);
or U268 (N_268,In_10,In_91);
nand U269 (N_269,In_254,In_39);
and U270 (N_270,In_44,In_495);
nand U271 (N_271,In_194,In_278);
or U272 (N_272,In_86,In_368);
nand U273 (N_273,In_219,In_354);
nor U274 (N_274,In_203,In_386);
and U275 (N_275,In_48,In_302);
or U276 (N_276,In_171,In_315);
xnor U277 (N_277,In_177,In_18);
or U278 (N_278,In_269,In_141);
or U279 (N_279,In_211,In_492);
nand U280 (N_280,In_47,In_402);
or U281 (N_281,In_137,In_2);
nand U282 (N_282,In_142,In_336);
and U283 (N_283,In_271,In_497);
nand U284 (N_284,In_385,In_474);
or U285 (N_285,In_340,In_421);
or U286 (N_286,In_255,In_455);
nand U287 (N_287,In_196,In_393);
or U288 (N_288,In_30,In_487);
or U289 (N_289,In_386,In_213);
nor U290 (N_290,In_306,In_244);
or U291 (N_291,In_326,In_61);
nor U292 (N_292,In_412,In_131);
or U293 (N_293,In_199,In_130);
nand U294 (N_294,In_434,In_153);
or U295 (N_295,In_404,In_81);
or U296 (N_296,In_152,In_369);
or U297 (N_297,In_232,In_373);
or U298 (N_298,In_192,In_152);
or U299 (N_299,In_484,In_237);
or U300 (N_300,In_98,In_281);
and U301 (N_301,In_387,In_327);
and U302 (N_302,In_108,In_315);
nand U303 (N_303,In_323,In_234);
and U304 (N_304,In_292,In_235);
nand U305 (N_305,In_388,In_45);
nor U306 (N_306,In_319,In_308);
xor U307 (N_307,In_16,In_480);
nor U308 (N_308,In_56,In_461);
nand U309 (N_309,In_422,In_218);
nor U310 (N_310,In_295,In_86);
nor U311 (N_311,In_329,In_433);
and U312 (N_312,In_125,In_330);
and U313 (N_313,In_46,In_82);
and U314 (N_314,In_28,In_21);
or U315 (N_315,In_36,In_384);
and U316 (N_316,In_272,In_284);
nor U317 (N_317,In_15,In_196);
nor U318 (N_318,In_359,In_192);
nor U319 (N_319,In_258,In_493);
or U320 (N_320,In_319,In_65);
nand U321 (N_321,In_224,In_296);
xor U322 (N_322,In_180,In_213);
or U323 (N_323,In_109,In_466);
or U324 (N_324,In_348,In_361);
nor U325 (N_325,In_123,In_399);
nor U326 (N_326,In_398,In_323);
nand U327 (N_327,In_37,In_22);
and U328 (N_328,In_298,In_395);
or U329 (N_329,In_400,In_294);
and U330 (N_330,In_93,In_239);
or U331 (N_331,In_495,In_82);
and U332 (N_332,In_189,In_294);
nand U333 (N_333,In_382,In_92);
or U334 (N_334,In_32,In_37);
nand U335 (N_335,In_46,In_491);
nand U336 (N_336,In_11,In_311);
and U337 (N_337,In_250,In_77);
nand U338 (N_338,In_196,In_261);
nand U339 (N_339,In_452,In_427);
and U340 (N_340,In_386,In_251);
or U341 (N_341,In_138,In_182);
or U342 (N_342,In_17,In_134);
nor U343 (N_343,In_247,In_187);
nor U344 (N_344,In_314,In_125);
nand U345 (N_345,In_281,In_171);
nor U346 (N_346,In_357,In_362);
or U347 (N_347,In_286,In_21);
and U348 (N_348,In_499,In_171);
or U349 (N_349,In_479,In_291);
and U350 (N_350,In_348,In_36);
nand U351 (N_351,In_434,In_269);
nor U352 (N_352,In_10,In_95);
nor U353 (N_353,In_96,In_380);
and U354 (N_354,In_187,In_1);
nor U355 (N_355,In_273,In_210);
nor U356 (N_356,In_134,In_110);
nand U357 (N_357,In_229,In_194);
nor U358 (N_358,In_314,In_194);
xnor U359 (N_359,In_164,In_162);
and U360 (N_360,In_415,In_11);
or U361 (N_361,In_444,In_47);
and U362 (N_362,In_26,In_427);
and U363 (N_363,In_167,In_136);
nand U364 (N_364,In_27,In_272);
nand U365 (N_365,In_264,In_253);
and U366 (N_366,In_451,In_37);
or U367 (N_367,In_141,In_238);
or U368 (N_368,In_23,In_120);
nand U369 (N_369,In_200,In_297);
nor U370 (N_370,In_185,In_268);
or U371 (N_371,In_315,In_1);
and U372 (N_372,In_17,In_25);
nor U373 (N_373,In_410,In_331);
and U374 (N_374,In_32,In_150);
and U375 (N_375,In_3,In_163);
or U376 (N_376,In_397,In_257);
nor U377 (N_377,In_35,In_118);
nor U378 (N_378,In_215,In_161);
xor U379 (N_379,In_39,In_152);
nor U380 (N_380,In_390,In_293);
nor U381 (N_381,In_351,In_56);
or U382 (N_382,In_33,In_175);
and U383 (N_383,In_38,In_235);
nor U384 (N_384,In_35,In_91);
nand U385 (N_385,In_249,In_251);
nand U386 (N_386,In_309,In_231);
nand U387 (N_387,In_102,In_288);
and U388 (N_388,In_453,In_423);
nor U389 (N_389,In_383,In_404);
nor U390 (N_390,In_204,In_441);
nor U391 (N_391,In_402,In_92);
nand U392 (N_392,In_112,In_247);
and U393 (N_393,In_273,In_11);
and U394 (N_394,In_61,In_390);
nand U395 (N_395,In_142,In_320);
nand U396 (N_396,In_202,In_149);
and U397 (N_397,In_451,In_364);
and U398 (N_398,In_235,In_228);
and U399 (N_399,In_412,In_492);
nor U400 (N_400,In_122,In_39);
or U401 (N_401,In_255,In_195);
nor U402 (N_402,In_360,In_81);
or U403 (N_403,In_248,In_273);
nand U404 (N_404,In_207,In_31);
nor U405 (N_405,In_239,In_11);
nor U406 (N_406,In_477,In_415);
and U407 (N_407,In_175,In_128);
and U408 (N_408,In_153,In_155);
nand U409 (N_409,In_169,In_333);
nand U410 (N_410,In_281,In_93);
or U411 (N_411,In_302,In_227);
nand U412 (N_412,In_131,In_279);
and U413 (N_413,In_180,In_63);
and U414 (N_414,In_362,In_318);
nand U415 (N_415,In_156,In_375);
and U416 (N_416,In_93,In_377);
or U417 (N_417,In_368,In_194);
nor U418 (N_418,In_202,In_30);
nand U419 (N_419,In_327,In_233);
nand U420 (N_420,In_412,In_453);
nor U421 (N_421,In_321,In_233);
nor U422 (N_422,In_451,In_36);
nand U423 (N_423,In_52,In_305);
or U424 (N_424,In_483,In_442);
xor U425 (N_425,In_56,In_494);
nor U426 (N_426,In_16,In_261);
nand U427 (N_427,In_334,In_379);
or U428 (N_428,In_252,In_379);
nor U429 (N_429,In_403,In_44);
and U430 (N_430,In_174,In_478);
or U431 (N_431,In_263,In_285);
and U432 (N_432,In_250,In_23);
or U433 (N_433,In_315,In_73);
and U434 (N_434,In_244,In_345);
or U435 (N_435,In_272,In_220);
nor U436 (N_436,In_239,In_294);
nand U437 (N_437,In_437,In_52);
nand U438 (N_438,In_325,In_155);
nand U439 (N_439,In_95,In_142);
nor U440 (N_440,In_265,In_185);
or U441 (N_441,In_463,In_27);
and U442 (N_442,In_250,In_307);
or U443 (N_443,In_458,In_151);
or U444 (N_444,In_471,In_444);
or U445 (N_445,In_460,In_340);
or U446 (N_446,In_318,In_46);
and U447 (N_447,In_167,In_158);
nand U448 (N_448,In_489,In_271);
xnor U449 (N_449,In_108,In_112);
nand U450 (N_450,In_206,In_131);
and U451 (N_451,In_286,In_87);
or U452 (N_452,In_185,In_474);
nand U453 (N_453,In_161,In_15);
and U454 (N_454,In_310,In_311);
or U455 (N_455,In_439,In_321);
or U456 (N_456,In_256,In_3);
nor U457 (N_457,In_4,In_362);
nor U458 (N_458,In_79,In_144);
and U459 (N_459,In_3,In_82);
nand U460 (N_460,In_479,In_218);
nand U461 (N_461,In_198,In_440);
and U462 (N_462,In_472,In_310);
and U463 (N_463,In_220,In_82);
nor U464 (N_464,In_49,In_473);
nand U465 (N_465,In_311,In_170);
and U466 (N_466,In_340,In_60);
or U467 (N_467,In_392,In_119);
and U468 (N_468,In_89,In_311);
nand U469 (N_469,In_440,In_387);
nand U470 (N_470,In_80,In_297);
nor U471 (N_471,In_35,In_383);
nor U472 (N_472,In_289,In_228);
and U473 (N_473,In_138,In_384);
nor U474 (N_474,In_144,In_313);
nor U475 (N_475,In_250,In_411);
or U476 (N_476,In_253,In_295);
nand U477 (N_477,In_427,In_228);
and U478 (N_478,In_23,In_147);
and U479 (N_479,In_260,In_11);
or U480 (N_480,In_367,In_127);
xnor U481 (N_481,In_312,In_128);
nor U482 (N_482,In_48,In_318);
and U483 (N_483,In_350,In_357);
or U484 (N_484,In_174,In_272);
nor U485 (N_485,In_299,In_159);
and U486 (N_486,In_345,In_113);
or U487 (N_487,In_36,In_151);
or U488 (N_488,In_11,In_91);
or U489 (N_489,In_267,In_251);
nand U490 (N_490,In_484,In_90);
nor U491 (N_491,In_476,In_98);
and U492 (N_492,In_476,In_334);
and U493 (N_493,In_412,In_253);
and U494 (N_494,In_445,In_236);
and U495 (N_495,In_410,In_459);
and U496 (N_496,In_90,In_23);
and U497 (N_497,In_1,In_179);
nand U498 (N_498,In_376,In_169);
and U499 (N_499,In_218,In_498);
nand U500 (N_500,In_16,In_9);
nor U501 (N_501,In_194,In_157);
nor U502 (N_502,In_257,In_308);
nor U503 (N_503,In_28,In_164);
xnor U504 (N_504,In_123,In_392);
nand U505 (N_505,In_202,In_467);
and U506 (N_506,In_231,In_272);
and U507 (N_507,In_0,In_71);
nor U508 (N_508,In_178,In_24);
nand U509 (N_509,In_445,In_326);
nor U510 (N_510,In_11,In_405);
and U511 (N_511,In_233,In_310);
or U512 (N_512,In_381,In_126);
nand U513 (N_513,In_160,In_7);
nor U514 (N_514,In_201,In_170);
nand U515 (N_515,In_420,In_498);
nor U516 (N_516,In_38,In_435);
and U517 (N_517,In_348,In_476);
nor U518 (N_518,In_146,In_169);
and U519 (N_519,In_361,In_207);
nor U520 (N_520,In_331,In_256);
nand U521 (N_521,In_385,In_448);
or U522 (N_522,In_370,In_478);
nor U523 (N_523,In_475,In_26);
or U524 (N_524,In_215,In_245);
and U525 (N_525,In_71,In_179);
and U526 (N_526,In_134,In_173);
or U527 (N_527,In_68,In_237);
or U528 (N_528,In_169,In_27);
and U529 (N_529,In_441,In_59);
or U530 (N_530,In_396,In_418);
nor U531 (N_531,In_425,In_437);
nand U532 (N_532,In_256,In_148);
xnor U533 (N_533,In_365,In_187);
and U534 (N_534,In_108,In_2);
or U535 (N_535,In_65,In_199);
nor U536 (N_536,In_308,In_265);
nor U537 (N_537,In_70,In_120);
nand U538 (N_538,In_11,In_295);
nor U539 (N_539,In_93,In_86);
and U540 (N_540,In_264,In_383);
nand U541 (N_541,In_180,In_309);
or U542 (N_542,In_64,In_401);
and U543 (N_543,In_491,In_417);
nand U544 (N_544,In_369,In_288);
and U545 (N_545,In_62,In_427);
and U546 (N_546,In_36,In_94);
nor U547 (N_547,In_164,In_123);
and U548 (N_548,In_281,In_267);
nand U549 (N_549,In_437,In_494);
nand U550 (N_550,In_184,In_111);
nor U551 (N_551,In_26,In_3);
nor U552 (N_552,In_442,In_110);
nor U553 (N_553,In_224,In_404);
nor U554 (N_554,In_402,In_154);
nand U555 (N_555,In_348,In_155);
or U556 (N_556,In_441,In_295);
nand U557 (N_557,In_214,In_27);
and U558 (N_558,In_60,In_208);
or U559 (N_559,In_137,In_96);
nand U560 (N_560,In_100,In_344);
nand U561 (N_561,In_487,In_294);
and U562 (N_562,In_485,In_499);
or U563 (N_563,In_343,In_485);
nand U564 (N_564,In_73,In_114);
nor U565 (N_565,In_453,In_28);
and U566 (N_566,In_383,In_12);
or U567 (N_567,In_100,In_404);
nand U568 (N_568,In_287,In_271);
or U569 (N_569,In_199,In_109);
or U570 (N_570,In_355,In_50);
nand U571 (N_571,In_7,In_114);
and U572 (N_572,In_90,In_76);
nor U573 (N_573,In_473,In_461);
nor U574 (N_574,In_221,In_207);
nor U575 (N_575,In_96,In_326);
nor U576 (N_576,In_223,In_135);
and U577 (N_577,In_108,In_11);
and U578 (N_578,In_258,In_496);
and U579 (N_579,In_378,In_69);
nand U580 (N_580,In_184,In_454);
nand U581 (N_581,In_20,In_39);
xnor U582 (N_582,In_368,In_91);
or U583 (N_583,In_347,In_173);
nand U584 (N_584,In_429,In_298);
and U585 (N_585,In_175,In_137);
nor U586 (N_586,In_185,In_231);
and U587 (N_587,In_323,In_374);
nor U588 (N_588,In_367,In_391);
or U589 (N_589,In_188,In_218);
nand U590 (N_590,In_482,In_161);
nor U591 (N_591,In_208,In_226);
nand U592 (N_592,In_390,In_249);
and U593 (N_593,In_19,In_122);
or U594 (N_594,In_341,In_61);
nand U595 (N_595,In_215,In_244);
nor U596 (N_596,In_36,In_225);
nor U597 (N_597,In_158,In_27);
nor U598 (N_598,In_200,In_414);
and U599 (N_599,In_132,In_217);
or U600 (N_600,In_254,In_396);
nand U601 (N_601,In_308,In_1);
and U602 (N_602,In_30,In_369);
and U603 (N_603,In_303,In_106);
and U604 (N_604,In_98,In_48);
nor U605 (N_605,In_255,In_274);
or U606 (N_606,In_440,In_447);
or U607 (N_607,In_66,In_399);
and U608 (N_608,In_175,In_337);
nor U609 (N_609,In_138,In_250);
and U610 (N_610,In_324,In_373);
nand U611 (N_611,In_128,In_22);
and U612 (N_612,In_316,In_409);
or U613 (N_613,In_359,In_393);
and U614 (N_614,In_390,In_9);
nor U615 (N_615,In_224,In_361);
or U616 (N_616,In_321,In_479);
nand U617 (N_617,In_389,In_462);
nor U618 (N_618,In_211,In_48);
and U619 (N_619,In_499,In_140);
nand U620 (N_620,In_482,In_140);
nor U621 (N_621,In_197,In_210);
xor U622 (N_622,In_381,In_430);
xnor U623 (N_623,In_7,In_395);
nor U624 (N_624,In_24,In_279);
or U625 (N_625,In_410,In_425);
nor U626 (N_626,In_272,In_359);
nor U627 (N_627,In_47,In_77);
and U628 (N_628,In_11,In_142);
nand U629 (N_629,In_247,In_351);
nor U630 (N_630,In_311,In_197);
nand U631 (N_631,In_352,In_266);
or U632 (N_632,In_278,In_433);
nand U633 (N_633,In_213,In_361);
and U634 (N_634,In_251,In_424);
nor U635 (N_635,In_406,In_6);
and U636 (N_636,In_147,In_417);
and U637 (N_637,In_468,In_462);
or U638 (N_638,In_4,In_18);
or U639 (N_639,In_212,In_79);
or U640 (N_640,In_104,In_149);
nor U641 (N_641,In_13,In_173);
xor U642 (N_642,In_406,In_195);
nand U643 (N_643,In_303,In_39);
nand U644 (N_644,In_337,In_297);
and U645 (N_645,In_235,In_433);
nor U646 (N_646,In_219,In_241);
nand U647 (N_647,In_495,In_418);
nor U648 (N_648,In_163,In_161);
and U649 (N_649,In_13,In_82);
nor U650 (N_650,In_365,In_417);
or U651 (N_651,In_202,In_266);
and U652 (N_652,In_22,In_420);
nor U653 (N_653,In_312,In_435);
or U654 (N_654,In_280,In_166);
nor U655 (N_655,In_304,In_215);
or U656 (N_656,In_176,In_115);
nand U657 (N_657,In_37,In_389);
nor U658 (N_658,In_332,In_441);
nand U659 (N_659,In_344,In_101);
nand U660 (N_660,In_273,In_388);
and U661 (N_661,In_435,In_261);
nand U662 (N_662,In_279,In_247);
or U663 (N_663,In_110,In_322);
nand U664 (N_664,In_409,In_103);
nand U665 (N_665,In_229,In_170);
and U666 (N_666,In_296,In_291);
nor U667 (N_667,In_243,In_312);
nor U668 (N_668,In_180,In_163);
and U669 (N_669,In_481,In_32);
nor U670 (N_670,In_61,In_200);
nand U671 (N_671,In_477,In_145);
or U672 (N_672,In_31,In_273);
nor U673 (N_673,In_33,In_211);
or U674 (N_674,In_19,In_476);
nand U675 (N_675,In_483,In_255);
or U676 (N_676,In_454,In_421);
or U677 (N_677,In_416,In_288);
and U678 (N_678,In_479,In_207);
and U679 (N_679,In_64,In_118);
nor U680 (N_680,In_329,In_98);
or U681 (N_681,In_154,In_451);
or U682 (N_682,In_117,In_239);
nand U683 (N_683,In_207,In_269);
and U684 (N_684,In_78,In_314);
nor U685 (N_685,In_191,In_13);
nor U686 (N_686,In_136,In_370);
nor U687 (N_687,In_474,In_493);
nor U688 (N_688,In_20,In_398);
and U689 (N_689,In_484,In_76);
nor U690 (N_690,In_401,In_72);
xor U691 (N_691,In_11,In_145);
nand U692 (N_692,In_179,In_57);
nand U693 (N_693,In_219,In_494);
and U694 (N_694,In_96,In_213);
or U695 (N_695,In_372,In_187);
nor U696 (N_696,In_456,In_286);
and U697 (N_697,In_267,In_168);
and U698 (N_698,In_122,In_461);
or U699 (N_699,In_313,In_335);
nor U700 (N_700,In_345,In_320);
xor U701 (N_701,In_466,In_196);
or U702 (N_702,In_262,In_484);
or U703 (N_703,In_405,In_129);
and U704 (N_704,In_143,In_6);
and U705 (N_705,In_245,In_221);
nand U706 (N_706,In_372,In_121);
or U707 (N_707,In_91,In_427);
or U708 (N_708,In_170,In_345);
nand U709 (N_709,In_96,In_475);
nand U710 (N_710,In_354,In_317);
nand U711 (N_711,In_293,In_299);
and U712 (N_712,In_417,In_479);
and U713 (N_713,In_59,In_6);
or U714 (N_714,In_242,In_183);
nand U715 (N_715,In_57,In_50);
or U716 (N_716,In_157,In_423);
nand U717 (N_717,In_12,In_145);
nand U718 (N_718,In_290,In_228);
nand U719 (N_719,In_272,In_103);
nand U720 (N_720,In_397,In_23);
xnor U721 (N_721,In_464,In_394);
nand U722 (N_722,In_10,In_241);
nand U723 (N_723,In_69,In_459);
nand U724 (N_724,In_183,In_385);
or U725 (N_725,In_334,In_291);
and U726 (N_726,In_209,In_412);
nand U727 (N_727,In_424,In_74);
xor U728 (N_728,In_371,In_440);
or U729 (N_729,In_238,In_183);
nor U730 (N_730,In_223,In_75);
and U731 (N_731,In_129,In_412);
nand U732 (N_732,In_270,In_313);
nor U733 (N_733,In_452,In_23);
or U734 (N_734,In_21,In_287);
or U735 (N_735,In_188,In_424);
and U736 (N_736,In_277,In_64);
or U737 (N_737,In_486,In_385);
nor U738 (N_738,In_354,In_229);
xnor U739 (N_739,In_91,In_103);
nand U740 (N_740,In_63,In_27);
xor U741 (N_741,In_322,In_308);
xor U742 (N_742,In_40,In_395);
nand U743 (N_743,In_15,In_322);
xor U744 (N_744,In_400,In_163);
and U745 (N_745,In_283,In_462);
nand U746 (N_746,In_73,In_64);
nand U747 (N_747,In_55,In_231);
nand U748 (N_748,In_166,In_342);
xor U749 (N_749,In_44,In_168);
nor U750 (N_750,N_294,N_689);
nand U751 (N_751,N_175,N_212);
or U752 (N_752,N_110,N_446);
or U753 (N_753,N_564,N_639);
or U754 (N_754,N_655,N_599);
nand U755 (N_755,N_40,N_198);
or U756 (N_756,N_681,N_0);
and U757 (N_757,N_183,N_744);
or U758 (N_758,N_426,N_72);
and U759 (N_759,N_47,N_596);
or U760 (N_760,N_109,N_589);
and U761 (N_761,N_113,N_66);
or U762 (N_762,N_399,N_277);
xor U763 (N_763,N_76,N_532);
xnor U764 (N_764,N_20,N_11);
or U765 (N_765,N_30,N_497);
and U766 (N_766,N_629,N_613);
nor U767 (N_767,N_59,N_667);
nand U768 (N_768,N_105,N_290);
xnor U769 (N_769,N_563,N_507);
nand U770 (N_770,N_618,N_420);
nor U771 (N_771,N_631,N_389);
and U772 (N_772,N_99,N_575);
nand U773 (N_773,N_202,N_634);
and U774 (N_774,N_423,N_576);
or U775 (N_775,N_508,N_169);
and U776 (N_776,N_482,N_658);
and U777 (N_777,N_236,N_232);
or U778 (N_778,N_41,N_356);
or U779 (N_779,N_354,N_579);
or U780 (N_780,N_644,N_205);
and U781 (N_781,N_250,N_227);
or U782 (N_782,N_612,N_404);
xnor U783 (N_783,N_249,N_359);
nor U784 (N_784,N_546,N_738);
nor U785 (N_785,N_429,N_97);
nor U786 (N_786,N_502,N_338);
or U787 (N_787,N_664,N_69);
nand U788 (N_788,N_188,N_472);
and U789 (N_789,N_272,N_696);
and U790 (N_790,N_263,N_311);
nand U791 (N_791,N_165,N_710);
nand U792 (N_792,N_746,N_28);
nand U793 (N_793,N_75,N_657);
and U794 (N_794,N_641,N_244);
or U795 (N_795,N_112,N_316);
nand U796 (N_796,N_329,N_485);
nand U797 (N_797,N_96,N_384);
nand U798 (N_798,N_585,N_293);
and U799 (N_799,N_600,N_719);
nor U800 (N_800,N_217,N_163);
and U801 (N_801,N_180,N_314);
nor U802 (N_802,N_360,N_184);
nor U803 (N_803,N_385,N_70);
and U804 (N_804,N_684,N_457);
nor U805 (N_805,N_101,N_155);
and U806 (N_806,N_495,N_405);
and U807 (N_807,N_428,N_427);
nand U808 (N_808,N_568,N_661);
and U809 (N_809,N_173,N_619);
and U810 (N_810,N_201,N_477);
nor U811 (N_811,N_79,N_391);
or U812 (N_812,N_462,N_572);
nand U813 (N_813,N_583,N_119);
or U814 (N_814,N_668,N_145);
or U815 (N_815,N_239,N_717);
nand U816 (N_816,N_117,N_274);
nand U817 (N_817,N_56,N_182);
or U818 (N_818,N_256,N_471);
or U819 (N_819,N_143,N_697);
nor U820 (N_820,N_551,N_255);
and U821 (N_821,N_87,N_594);
and U822 (N_822,N_16,N_95);
or U823 (N_823,N_614,N_549);
and U824 (N_824,N_642,N_582);
nor U825 (N_825,N_167,N_622);
and U826 (N_826,N_50,N_677);
nor U827 (N_827,N_139,N_142);
nand U828 (N_828,N_665,N_616);
xnor U829 (N_829,N_211,N_694);
and U830 (N_830,N_104,N_181);
or U831 (N_831,N_645,N_62);
nor U832 (N_832,N_547,N_518);
or U833 (N_833,N_149,N_176);
nor U834 (N_834,N_561,N_410);
and U835 (N_835,N_271,N_504);
or U836 (N_836,N_748,N_269);
nor U837 (N_837,N_83,N_732);
nor U838 (N_838,N_168,N_479);
nor U839 (N_839,N_348,N_610);
nand U840 (N_840,N_45,N_193);
or U841 (N_841,N_353,N_402);
nor U842 (N_842,N_400,N_125);
nand U843 (N_843,N_261,N_206);
nor U844 (N_844,N_510,N_492);
and U845 (N_845,N_682,N_591);
and U846 (N_846,N_73,N_268);
and U847 (N_847,N_628,N_693);
nor U848 (N_848,N_301,N_608);
nor U849 (N_849,N_289,N_185);
xnor U850 (N_850,N_345,N_323);
nand U851 (N_851,N_364,N_299);
xnor U852 (N_852,N_150,N_520);
nor U853 (N_853,N_32,N_553);
or U854 (N_854,N_339,N_539);
and U855 (N_855,N_636,N_230);
and U856 (N_856,N_499,N_229);
nand U857 (N_857,N_52,N_25);
and U858 (N_858,N_533,N_154);
or U859 (N_859,N_308,N_147);
nor U860 (N_860,N_355,N_670);
or U861 (N_861,N_573,N_170);
nand U862 (N_862,N_126,N_254);
nor U863 (N_863,N_525,N_687);
nand U864 (N_864,N_567,N_146);
and U865 (N_865,N_44,N_476);
or U866 (N_866,N_68,N_128);
xnor U867 (N_867,N_243,N_82);
nor U868 (N_868,N_611,N_23);
or U869 (N_869,N_577,N_432);
nand U870 (N_870,N_55,N_559);
and U871 (N_871,N_124,N_24);
nand U872 (N_872,N_447,N_469);
nand U873 (N_873,N_723,N_312);
nor U874 (N_874,N_238,N_392);
xor U875 (N_875,N_709,N_140);
and U876 (N_876,N_463,N_262);
nand U877 (N_877,N_298,N_258);
and U878 (N_878,N_593,N_503);
nand U879 (N_879,N_538,N_341);
nor U880 (N_880,N_587,N_395);
nor U881 (N_881,N_380,N_315);
and U882 (N_882,N_61,N_179);
and U883 (N_883,N_550,N_643);
nand U884 (N_884,N_100,N_376);
nand U885 (N_885,N_248,N_332);
nor U886 (N_886,N_386,N_35);
nand U887 (N_887,N_602,N_541);
nand U888 (N_888,N_333,N_187);
and U889 (N_889,N_204,N_557);
or U890 (N_890,N_725,N_586);
nand U891 (N_891,N_7,N_42);
nor U892 (N_892,N_106,N_451);
or U893 (N_893,N_191,N_77);
nor U894 (N_894,N_449,N_407);
nand U895 (N_895,N_555,N_85);
or U896 (N_896,N_578,N_291);
and U897 (N_897,N_418,N_515);
nor U898 (N_898,N_749,N_127);
nor U899 (N_899,N_220,N_287);
and U900 (N_900,N_344,N_63);
nor U901 (N_901,N_422,N_607);
nand U902 (N_902,N_9,N_114);
or U903 (N_903,N_162,N_718);
or U904 (N_904,N_240,N_200);
or U905 (N_905,N_424,N_413);
and U906 (N_906,N_671,N_226);
nor U907 (N_907,N_715,N_235);
and U908 (N_908,N_158,N_213);
nor U909 (N_909,N_86,N_417);
nor U910 (N_910,N_433,N_488);
or U911 (N_911,N_489,N_686);
or U912 (N_912,N_615,N_527);
or U913 (N_913,N_595,N_306);
nand U914 (N_914,N_703,N_493);
and U915 (N_915,N_328,N_394);
and U916 (N_916,N_490,N_219);
xor U917 (N_917,N_14,N_597);
or U918 (N_918,N_735,N_552);
nand U919 (N_919,N_29,N_509);
nand U920 (N_920,N_635,N_465);
nand U921 (N_921,N_390,N_278);
nor U922 (N_922,N_584,N_27);
nor U923 (N_923,N_171,N_396);
and U924 (N_924,N_729,N_441);
nand U925 (N_925,N_15,N_324);
or U926 (N_926,N_340,N_372);
and U927 (N_927,N_604,N_6);
xor U928 (N_928,N_461,N_253);
or U929 (N_929,N_218,N_406);
nor U930 (N_930,N_517,N_39);
nand U931 (N_931,N_172,N_414);
or U932 (N_932,N_233,N_692);
nand U933 (N_933,N_501,N_444);
nor U934 (N_934,N_470,N_475);
nor U935 (N_935,N_588,N_5);
and U936 (N_936,N_702,N_606);
nand U937 (N_937,N_673,N_565);
nor U938 (N_938,N_474,N_581);
or U939 (N_939,N_483,N_459);
or U940 (N_940,N_535,N_357);
nor U941 (N_941,N_649,N_369);
nor U942 (N_942,N_91,N_295);
or U943 (N_943,N_706,N_279);
and U944 (N_944,N_669,N_53);
nor U945 (N_945,N_231,N_448);
nor U946 (N_946,N_603,N_720);
and U947 (N_947,N_519,N_144);
nand U948 (N_948,N_374,N_280);
and U949 (N_949,N_659,N_487);
or U950 (N_950,N_466,N_51);
nand U951 (N_951,N_209,N_307);
nor U952 (N_952,N_199,N_98);
and U953 (N_953,N_352,N_393);
or U954 (N_954,N_660,N_136);
nand U955 (N_955,N_318,N_327);
nand U956 (N_956,N_652,N_152);
nand U957 (N_957,N_81,N_713);
and U958 (N_958,N_733,N_726);
nand U959 (N_959,N_724,N_92);
nand U960 (N_960,N_54,N_438);
and U961 (N_961,N_467,N_458);
nand U962 (N_962,N_260,N_166);
or U963 (N_963,N_131,N_522);
nor U964 (N_964,N_303,N_672);
nor U965 (N_965,N_305,N_727);
nand U966 (N_966,N_722,N_304);
xor U967 (N_967,N_309,N_129);
and U968 (N_968,N_317,N_580);
nand U969 (N_969,N_464,N_242);
and U970 (N_970,N_58,N_22);
nand U971 (N_971,N_270,N_196);
xor U972 (N_972,N_2,N_452);
or U973 (N_973,N_342,N_688);
nand U974 (N_974,N_273,N_496);
nor U975 (N_975,N_554,N_267);
nand U976 (N_976,N_450,N_118);
nand U977 (N_977,N_536,N_358);
or U978 (N_978,N_26,N_285);
xnor U979 (N_979,N_743,N_494);
nand U980 (N_980,N_313,N_67);
xor U981 (N_981,N_337,N_370);
nand U982 (N_982,N_361,N_210);
nand U983 (N_983,N_111,N_102);
nand U984 (N_984,N_19,N_49);
or U985 (N_985,N_71,N_368);
and U986 (N_986,N_617,N_115);
nor U987 (N_987,N_592,N_569);
nor U988 (N_988,N_730,N_88);
and U989 (N_989,N_473,N_728);
or U990 (N_990,N_431,N_133);
and U991 (N_991,N_506,N_43);
and U992 (N_992,N_731,N_282);
nor U993 (N_993,N_663,N_34);
and U994 (N_994,N_701,N_4);
nor U995 (N_995,N_605,N_46);
nand U996 (N_996,N_284,N_297);
nor U997 (N_997,N_257,N_17);
or U998 (N_998,N_484,N_708);
and U999 (N_999,N_122,N_264);
or U1000 (N_1000,N_695,N_443);
and U1001 (N_1001,N_378,N_350);
nand U1002 (N_1002,N_300,N_624);
nor U1003 (N_1003,N_120,N_135);
nor U1004 (N_1004,N_349,N_178);
or U1005 (N_1005,N_387,N_455);
or U1006 (N_1006,N_534,N_37);
and U1007 (N_1007,N_13,N_521);
nor U1008 (N_1008,N_542,N_132);
and U1009 (N_1009,N_678,N_524);
or U1010 (N_1010,N_78,N_656);
or U1011 (N_1011,N_416,N_151);
and U1012 (N_1012,N_365,N_189);
nor U1013 (N_1013,N_377,N_160);
nand U1014 (N_1014,N_601,N_12);
nor U1015 (N_1015,N_434,N_397);
and U1016 (N_1016,N_570,N_409);
nand U1017 (N_1017,N_445,N_228);
nand U1018 (N_1018,N_453,N_505);
and U1019 (N_1019,N_620,N_225);
nor U1020 (N_1020,N_425,N_736);
or U1021 (N_1021,N_468,N_224);
nor U1022 (N_1022,N_107,N_164);
or U1023 (N_1023,N_711,N_740);
and U1024 (N_1024,N_543,N_215);
nand U1025 (N_1025,N_556,N_566);
and U1026 (N_1026,N_21,N_138);
or U1027 (N_1027,N_203,N_675);
nand U1028 (N_1028,N_331,N_362);
and U1029 (N_1029,N_621,N_121);
nor U1030 (N_1030,N_412,N_383);
nor U1031 (N_1031,N_245,N_545);
or U1032 (N_1032,N_638,N_430);
nand U1033 (N_1033,N_346,N_321);
nand U1034 (N_1034,N_653,N_500);
and U1035 (N_1035,N_286,N_623);
or U1036 (N_1036,N_275,N_174);
nand U1037 (N_1037,N_347,N_266);
nand U1038 (N_1038,N_699,N_363);
or U1039 (N_1039,N_491,N_398);
nand U1040 (N_1040,N_421,N_10);
nand U1041 (N_1041,N_530,N_705);
and U1042 (N_1042,N_640,N_646);
or U1043 (N_1043,N_721,N_288);
nor U1044 (N_1044,N_666,N_153);
and U1045 (N_1045,N_246,N_562);
nand U1046 (N_1046,N_241,N_161);
or U1047 (N_1047,N_265,N_90);
or U1048 (N_1048,N_512,N_190);
nand U1049 (N_1049,N_320,N_237);
or U1050 (N_1050,N_247,N_408);
nor U1051 (N_1051,N_498,N_442);
nor U1052 (N_1052,N_343,N_351);
nand U1053 (N_1053,N_630,N_511);
or U1054 (N_1054,N_537,N_33);
nor U1055 (N_1055,N_330,N_123);
nand U1056 (N_1056,N_326,N_379);
or U1057 (N_1057,N_419,N_283);
nand U1058 (N_1058,N_544,N_439);
nand U1059 (N_1059,N_103,N_222);
and U1060 (N_1060,N_401,N_281);
and U1061 (N_1061,N_214,N_516);
nor U1062 (N_1062,N_64,N_674);
nor U1063 (N_1063,N_745,N_177);
and U1064 (N_1064,N_197,N_1);
nand U1065 (N_1065,N_478,N_251);
or U1066 (N_1066,N_741,N_481);
and U1067 (N_1067,N_676,N_65);
nand U1068 (N_1068,N_8,N_156);
or U1069 (N_1069,N_528,N_3);
xor U1070 (N_1070,N_625,N_80);
nand U1071 (N_1071,N_207,N_371);
nand U1072 (N_1072,N_94,N_513);
nand U1073 (N_1073,N_737,N_325);
nor U1074 (N_1074,N_159,N_707);
and U1075 (N_1075,N_529,N_651);
nor U1076 (N_1076,N_310,N_480);
and U1077 (N_1077,N_195,N_208);
and U1078 (N_1078,N_574,N_366);
and U1079 (N_1079,N_367,N_531);
or U1080 (N_1080,N_335,N_319);
nand U1081 (N_1081,N_252,N_192);
and U1082 (N_1082,N_626,N_704);
nor U1083 (N_1083,N_194,N_747);
nor U1084 (N_1084,N_116,N_685);
and U1085 (N_1085,N_683,N_137);
or U1086 (N_1086,N_662,N_93);
or U1087 (N_1087,N_296,N_571);
nor U1088 (N_1088,N_632,N_540);
and U1089 (N_1089,N_221,N_322);
and U1090 (N_1090,N_700,N_31);
or U1091 (N_1091,N_382,N_691);
nand U1092 (N_1092,N_548,N_698);
nor U1093 (N_1093,N_36,N_60);
or U1094 (N_1094,N_388,N_712);
nor U1095 (N_1095,N_57,N_415);
nand U1096 (N_1096,N_523,N_436);
or U1097 (N_1097,N_292,N_437);
and U1098 (N_1098,N_648,N_690);
nand U1099 (N_1099,N_526,N_460);
nor U1100 (N_1100,N_148,N_627);
and U1101 (N_1101,N_411,N_157);
nor U1102 (N_1102,N_259,N_276);
or U1103 (N_1103,N_440,N_650);
nand U1104 (N_1104,N_734,N_48);
or U1105 (N_1105,N_742,N_590);
or U1106 (N_1106,N_647,N_609);
nand U1107 (N_1107,N_435,N_89);
or U1108 (N_1108,N_714,N_234);
or U1109 (N_1109,N_141,N_403);
or U1110 (N_1110,N_514,N_637);
or U1111 (N_1111,N_375,N_336);
nand U1112 (N_1112,N_186,N_454);
or U1113 (N_1113,N_223,N_302);
nor U1114 (N_1114,N_84,N_598);
nor U1115 (N_1115,N_130,N_381);
nand U1116 (N_1116,N_739,N_108);
or U1117 (N_1117,N_560,N_633);
nor U1118 (N_1118,N_134,N_486);
and U1119 (N_1119,N_38,N_216);
and U1120 (N_1120,N_558,N_456);
and U1121 (N_1121,N_18,N_654);
xor U1122 (N_1122,N_334,N_680);
nand U1123 (N_1123,N_716,N_74);
nand U1124 (N_1124,N_373,N_679);
or U1125 (N_1125,N_733,N_3);
nor U1126 (N_1126,N_464,N_289);
nor U1127 (N_1127,N_20,N_171);
nor U1128 (N_1128,N_528,N_333);
nor U1129 (N_1129,N_524,N_579);
and U1130 (N_1130,N_700,N_697);
and U1131 (N_1131,N_366,N_176);
nor U1132 (N_1132,N_516,N_535);
xor U1133 (N_1133,N_706,N_93);
and U1134 (N_1134,N_85,N_291);
nand U1135 (N_1135,N_20,N_507);
and U1136 (N_1136,N_672,N_486);
or U1137 (N_1137,N_683,N_317);
nand U1138 (N_1138,N_137,N_647);
and U1139 (N_1139,N_37,N_589);
nor U1140 (N_1140,N_216,N_656);
nor U1141 (N_1141,N_639,N_213);
and U1142 (N_1142,N_259,N_202);
nor U1143 (N_1143,N_174,N_344);
nand U1144 (N_1144,N_198,N_654);
nand U1145 (N_1145,N_306,N_362);
nor U1146 (N_1146,N_176,N_274);
and U1147 (N_1147,N_139,N_512);
nor U1148 (N_1148,N_339,N_135);
nor U1149 (N_1149,N_166,N_586);
and U1150 (N_1150,N_332,N_612);
nand U1151 (N_1151,N_567,N_315);
and U1152 (N_1152,N_143,N_739);
nor U1153 (N_1153,N_300,N_188);
nor U1154 (N_1154,N_574,N_406);
or U1155 (N_1155,N_23,N_433);
and U1156 (N_1156,N_652,N_97);
or U1157 (N_1157,N_222,N_209);
and U1158 (N_1158,N_386,N_582);
nand U1159 (N_1159,N_206,N_641);
or U1160 (N_1160,N_538,N_64);
or U1161 (N_1161,N_502,N_105);
and U1162 (N_1162,N_696,N_26);
or U1163 (N_1163,N_713,N_258);
and U1164 (N_1164,N_520,N_303);
nand U1165 (N_1165,N_8,N_650);
and U1166 (N_1166,N_320,N_640);
nor U1167 (N_1167,N_638,N_483);
nand U1168 (N_1168,N_366,N_253);
and U1169 (N_1169,N_715,N_188);
and U1170 (N_1170,N_248,N_45);
and U1171 (N_1171,N_167,N_624);
nor U1172 (N_1172,N_664,N_6);
nor U1173 (N_1173,N_609,N_704);
nor U1174 (N_1174,N_56,N_221);
nor U1175 (N_1175,N_628,N_696);
nor U1176 (N_1176,N_435,N_674);
or U1177 (N_1177,N_726,N_580);
or U1178 (N_1178,N_380,N_332);
and U1179 (N_1179,N_370,N_686);
and U1180 (N_1180,N_583,N_344);
nand U1181 (N_1181,N_455,N_183);
or U1182 (N_1182,N_355,N_23);
nand U1183 (N_1183,N_477,N_257);
or U1184 (N_1184,N_188,N_476);
nand U1185 (N_1185,N_411,N_328);
nor U1186 (N_1186,N_243,N_668);
and U1187 (N_1187,N_184,N_450);
or U1188 (N_1188,N_152,N_63);
nor U1189 (N_1189,N_623,N_327);
nand U1190 (N_1190,N_305,N_738);
or U1191 (N_1191,N_644,N_571);
and U1192 (N_1192,N_100,N_685);
nand U1193 (N_1193,N_40,N_27);
or U1194 (N_1194,N_689,N_377);
and U1195 (N_1195,N_101,N_152);
nand U1196 (N_1196,N_110,N_444);
and U1197 (N_1197,N_561,N_141);
or U1198 (N_1198,N_311,N_179);
nor U1199 (N_1199,N_624,N_437);
or U1200 (N_1200,N_491,N_287);
and U1201 (N_1201,N_270,N_174);
nor U1202 (N_1202,N_603,N_161);
or U1203 (N_1203,N_177,N_530);
nand U1204 (N_1204,N_172,N_330);
nor U1205 (N_1205,N_447,N_134);
nand U1206 (N_1206,N_247,N_719);
nand U1207 (N_1207,N_608,N_236);
and U1208 (N_1208,N_315,N_84);
or U1209 (N_1209,N_209,N_637);
and U1210 (N_1210,N_584,N_423);
or U1211 (N_1211,N_384,N_692);
or U1212 (N_1212,N_578,N_302);
and U1213 (N_1213,N_684,N_327);
or U1214 (N_1214,N_439,N_670);
and U1215 (N_1215,N_590,N_736);
nand U1216 (N_1216,N_162,N_97);
and U1217 (N_1217,N_597,N_715);
and U1218 (N_1218,N_252,N_701);
nor U1219 (N_1219,N_638,N_175);
or U1220 (N_1220,N_324,N_353);
or U1221 (N_1221,N_296,N_159);
nand U1222 (N_1222,N_503,N_510);
xnor U1223 (N_1223,N_429,N_514);
nand U1224 (N_1224,N_431,N_58);
nand U1225 (N_1225,N_50,N_552);
or U1226 (N_1226,N_570,N_519);
nand U1227 (N_1227,N_341,N_520);
nor U1228 (N_1228,N_624,N_421);
nand U1229 (N_1229,N_728,N_59);
nor U1230 (N_1230,N_523,N_422);
and U1231 (N_1231,N_689,N_305);
nor U1232 (N_1232,N_191,N_344);
and U1233 (N_1233,N_204,N_163);
nor U1234 (N_1234,N_502,N_506);
nand U1235 (N_1235,N_282,N_601);
nand U1236 (N_1236,N_69,N_49);
nor U1237 (N_1237,N_129,N_7);
nand U1238 (N_1238,N_662,N_661);
nor U1239 (N_1239,N_749,N_94);
or U1240 (N_1240,N_394,N_619);
and U1241 (N_1241,N_47,N_631);
nor U1242 (N_1242,N_2,N_105);
or U1243 (N_1243,N_748,N_469);
and U1244 (N_1244,N_6,N_74);
and U1245 (N_1245,N_320,N_559);
nor U1246 (N_1246,N_591,N_143);
or U1247 (N_1247,N_6,N_703);
nand U1248 (N_1248,N_126,N_679);
or U1249 (N_1249,N_403,N_139);
or U1250 (N_1250,N_227,N_738);
nor U1251 (N_1251,N_39,N_457);
nand U1252 (N_1252,N_143,N_328);
or U1253 (N_1253,N_498,N_673);
nand U1254 (N_1254,N_509,N_103);
xor U1255 (N_1255,N_663,N_458);
and U1256 (N_1256,N_45,N_295);
nand U1257 (N_1257,N_278,N_5);
and U1258 (N_1258,N_179,N_167);
nor U1259 (N_1259,N_474,N_412);
or U1260 (N_1260,N_174,N_186);
nand U1261 (N_1261,N_296,N_676);
or U1262 (N_1262,N_358,N_614);
or U1263 (N_1263,N_630,N_246);
nand U1264 (N_1264,N_601,N_50);
and U1265 (N_1265,N_278,N_415);
or U1266 (N_1266,N_59,N_307);
nor U1267 (N_1267,N_518,N_200);
and U1268 (N_1268,N_523,N_233);
or U1269 (N_1269,N_210,N_686);
or U1270 (N_1270,N_193,N_282);
nand U1271 (N_1271,N_385,N_602);
and U1272 (N_1272,N_401,N_367);
or U1273 (N_1273,N_3,N_313);
nor U1274 (N_1274,N_9,N_518);
nor U1275 (N_1275,N_458,N_189);
nand U1276 (N_1276,N_591,N_492);
nand U1277 (N_1277,N_589,N_420);
nor U1278 (N_1278,N_590,N_161);
or U1279 (N_1279,N_331,N_701);
and U1280 (N_1280,N_27,N_158);
nor U1281 (N_1281,N_701,N_434);
or U1282 (N_1282,N_745,N_396);
nand U1283 (N_1283,N_654,N_57);
and U1284 (N_1284,N_257,N_494);
nand U1285 (N_1285,N_155,N_505);
nor U1286 (N_1286,N_732,N_559);
or U1287 (N_1287,N_12,N_221);
nand U1288 (N_1288,N_654,N_460);
or U1289 (N_1289,N_564,N_350);
nand U1290 (N_1290,N_447,N_35);
and U1291 (N_1291,N_226,N_556);
or U1292 (N_1292,N_582,N_142);
nand U1293 (N_1293,N_57,N_508);
or U1294 (N_1294,N_535,N_657);
nor U1295 (N_1295,N_668,N_335);
nand U1296 (N_1296,N_123,N_510);
or U1297 (N_1297,N_28,N_329);
and U1298 (N_1298,N_306,N_341);
or U1299 (N_1299,N_631,N_711);
nand U1300 (N_1300,N_89,N_303);
nand U1301 (N_1301,N_123,N_72);
and U1302 (N_1302,N_16,N_382);
nand U1303 (N_1303,N_118,N_344);
nand U1304 (N_1304,N_307,N_435);
nand U1305 (N_1305,N_232,N_9);
nand U1306 (N_1306,N_289,N_734);
nand U1307 (N_1307,N_555,N_515);
nand U1308 (N_1308,N_46,N_57);
and U1309 (N_1309,N_240,N_329);
nor U1310 (N_1310,N_156,N_440);
and U1311 (N_1311,N_372,N_126);
nand U1312 (N_1312,N_429,N_240);
or U1313 (N_1313,N_384,N_169);
nand U1314 (N_1314,N_65,N_734);
or U1315 (N_1315,N_51,N_568);
or U1316 (N_1316,N_70,N_131);
nand U1317 (N_1317,N_611,N_305);
or U1318 (N_1318,N_251,N_325);
and U1319 (N_1319,N_540,N_272);
nor U1320 (N_1320,N_474,N_258);
and U1321 (N_1321,N_313,N_564);
nor U1322 (N_1322,N_409,N_457);
or U1323 (N_1323,N_747,N_90);
nor U1324 (N_1324,N_85,N_180);
or U1325 (N_1325,N_190,N_389);
nand U1326 (N_1326,N_259,N_388);
nor U1327 (N_1327,N_262,N_214);
xor U1328 (N_1328,N_159,N_387);
and U1329 (N_1329,N_661,N_304);
and U1330 (N_1330,N_21,N_668);
nor U1331 (N_1331,N_546,N_6);
nor U1332 (N_1332,N_223,N_681);
or U1333 (N_1333,N_559,N_487);
and U1334 (N_1334,N_123,N_594);
nand U1335 (N_1335,N_575,N_600);
nand U1336 (N_1336,N_414,N_386);
or U1337 (N_1337,N_494,N_515);
xnor U1338 (N_1338,N_67,N_351);
and U1339 (N_1339,N_560,N_691);
nand U1340 (N_1340,N_420,N_295);
nand U1341 (N_1341,N_296,N_13);
or U1342 (N_1342,N_69,N_175);
nor U1343 (N_1343,N_151,N_72);
nor U1344 (N_1344,N_4,N_188);
or U1345 (N_1345,N_195,N_703);
nor U1346 (N_1346,N_671,N_175);
nand U1347 (N_1347,N_237,N_332);
and U1348 (N_1348,N_594,N_372);
or U1349 (N_1349,N_19,N_316);
nor U1350 (N_1350,N_347,N_264);
nand U1351 (N_1351,N_293,N_442);
nand U1352 (N_1352,N_455,N_144);
or U1353 (N_1353,N_729,N_532);
nor U1354 (N_1354,N_77,N_299);
nor U1355 (N_1355,N_446,N_227);
or U1356 (N_1356,N_571,N_531);
nand U1357 (N_1357,N_450,N_191);
nand U1358 (N_1358,N_202,N_340);
nand U1359 (N_1359,N_461,N_388);
or U1360 (N_1360,N_351,N_363);
nor U1361 (N_1361,N_536,N_220);
nor U1362 (N_1362,N_97,N_575);
or U1363 (N_1363,N_70,N_499);
nand U1364 (N_1364,N_249,N_417);
or U1365 (N_1365,N_411,N_219);
nand U1366 (N_1366,N_565,N_651);
or U1367 (N_1367,N_482,N_398);
and U1368 (N_1368,N_246,N_97);
nand U1369 (N_1369,N_100,N_227);
and U1370 (N_1370,N_115,N_431);
or U1371 (N_1371,N_56,N_86);
and U1372 (N_1372,N_171,N_177);
xnor U1373 (N_1373,N_591,N_432);
nor U1374 (N_1374,N_175,N_691);
and U1375 (N_1375,N_572,N_83);
nand U1376 (N_1376,N_706,N_528);
or U1377 (N_1377,N_74,N_704);
or U1378 (N_1378,N_579,N_351);
nor U1379 (N_1379,N_569,N_522);
nand U1380 (N_1380,N_641,N_332);
nand U1381 (N_1381,N_403,N_239);
and U1382 (N_1382,N_455,N_551);
nor U1383 (N_1383,N_433,N_154);
nand U1384 (N_1384,N_307,N_102);
and U1385 (N_1385,N_371,N_536);
nand U1386 (N_1386,N_603,N_706);
nand U1387 (N_1387,N_571,N_318);
and U1388 (N_1388,N_446,N_125);
or U1389 (N_1389,N_704,N_11);
or U1390 (N_1390,N_212,N_88);
and U1391 (N_1391,N_296,N_726);
and U1392 (N_1392,N_117,N_639);
nand U1393 (N_1393,N_144,N_469);
nor U1394 (N_1394,N_527,N_97);
nor U1395 (N_1395,N_192,N_671);
and U1396 (N_1396,N_178,N_50);
and U1397 (N_1397,N_468,N_300);
or U1398 (N_1398,N_586,N_53);
and U1399 (N_1399,N_693,N_495);
nor U1400 (N_1400,N_691,N_496);
or U1401 (N_1401,N_1,N_418);
or U1402 (N_1402,N_605,N_405);
or U1403 (N_1403,N_387,N_308);
nand U1404 (N_1404,N_119,N_416);
or U1405 (N_1405,N_15,N_121);
and U1406 (N_1406,N_679,N_152);
nand U1407 (N_1407,N_575,N_0);
nand U1408 (N_1408,N_167,N_57);
nor U1409 (N_1409,N_176,N_345);
and U1410 (N_1410,N_383,N_535);
or U1411 (N_1411,N_737,N_339);
and U1412 (N_1412,N_735,N_452);
and U1413 (N_1413,N_53,N_207);
or U1414 (N_1414,N_302,N_243);
and U1415 (N_1415,N_522,N_401);
nor U1416 (N_1416,N_188,N_735);
or U1417 (N_1417,N_624,N_693);
and U1418 (N_1418,N_458,N_328);
or U1419 (N_1419,N_285,N_424);
nand U1420 (N_1420,N_388,N_287);
nor U1421 (N_1421,N_154,N_451);
or U1422 (N_1422,N_607,N_386);
and U1423 (N_1423,N_594,N_656);
or U1424 (N_1424,N_177,N_618);
or U1425 (N_1425,N_167,N_99);
nand U1426 (N_1426,N_593,N_332);
nand U1427 (N_1427,N_184,N_122);
nor U1428 (N_1428,N_709,N_226);
nand U1429 (N_1429,N_640,N_664);
nand U1430 (N_1430,N_548,N_677);
and U1431 (N_1431,N_491,N_213);
nand U1432 (N_1432,N_310,N_721);
or U1433 (N_1433,N_451,N_134);
and U1434 (N_1434,N_109,N_10);
nand U1435 (N_1435,N_342,N_134);
and U1436 (N_1436,N_190,N_264);
nor U1437 (N_1437,N_209,N_702);
xor U1438 (N_1438,N_696,N_88);
and U1439 (N_1439,N_59,N_567);
nor U1440 (N_1440,N_394,N_239);
or U1441 (N_1441,N_80,N_594);
and U1442 (N_1442,N_686,N_133);
or U1443 (N_1443,N_382,N_411);
or U1444 (N_1444,N_399,N_623);
nor U1445 (N_1445,N_745,N_618);
or U1446 (N_1446,N_220,N_497);
nor U1447 (N_1447,N_191,N_487);
nor U1448 (N_1448,N_6,N_171);
nand U1449 (N_1449,N_709,N_567);
nand U1450 (N_1450,N_566,N_76);
and U1451 (N_1451,N_133,N_9);
nor U1452 (N_1452,N_606,N_676);
nor U1453 (N_1453,N_523,N_216);
nor U1454 (N_1454,N_518,N_651);
nor U1455 (N_1455,N_376,N_685);
and U1456 (N_1456,N_225,N_69);
xor U1457 (N_1457,N_211,N_202);
or U1458 (N_1458,N_590,N_662);
or U1459 (N_1459,N_368,N_557);
nand U1460 (N_1460,N_527,N_466);
or U1461 (N_1461,N_211,N_119);
nand U1462 (N_1462,N_176,N_640);
nor U1463 (N_1463,N_410,N_692);
or U1464 (N_1464,N_1,N_74);
or U1465 (N_1465,N_149,N_200);
nor U1466 (N_1466,N_565,N_258);
and U1467 (N_1467,N_674,N_156);
nand U1468 (N_1468,N_557,N_689);
and U1469 (N_1469,N_390,N_513);
nor U1470 (N_1470,N_483,N_673);
or U1471 (N_1471,N_309,N_218);
nor U1472 (N_1472,N_426,N_156);
nand U1473 (N_1473,N_405,N_100);
nand U1474 (N_1474,N_539,N_620);
and U1475 (N_1475,N_334,N_42);
nand U1476 (N_1476,N_366,N_716);
or U1477 (N_1477,N_619,N_631);
nor U1478 (N_1478,N_475,N_186);
and U1479 (N_1479,N_650,N_552);
nor U1480 (N_1480,N_256,N_646);
or U1481 (N_1481,N_434,N_499);
nor U1482 (N_1482,N_101,N_602);
nor U1483 (N_1483,N_507,N_637);
or U1484 (N_1484,N_614,N_394);
nor U1485 (N_1485,N_205,N_731);
or U1486 (N_1486,N_655,N_22);
nand U1487 (N_1487,N_485,N_389);
nor U1488 (N_1488,N_633,N_378);
and U1489 (N_1489,N_424,N_2);
xnor U1490 (N_1490,N_512,N_324);
and U1491 (N_1491,N_621,N_5);
and U1492 (N_1492,N_294,N_48);
or U1493 (N_1493,N_507,N_639);
nor U1494 (N_1494,N_477,N_616);
nand U1495 (N_1495,N_414,N_710);
nand U1496 (N_1496,N_536,N_719);
nand U1497 (N_1497,N_519,N_328);
xnor U1498 (N_1498,N_747,N_748);
and U1499 (N_1499,N_510,N_57);
nor U1500 (N_1500,N_1497,N_928);
nand U1501 (N_1501,N_1475,N_1440);
nand U1502 (N_1502,N_992,N_844);
and U1503 (N_1503,N_1446,N_944);
nor U1504 (N_1504,N_938,N_1051);
nand U1505 (N_1505,N_761,N_1039);
nor U1506 (N_1506,N_948,N_1277);
or U1507 (N_1507,N_1182,N_1049);
and U1508 (N_1508,N_1250,N_1476);
nand U1509 (N_1509,N_1268,N_1202);
and U1510 (N_1510,N_805,N_766);
or U1511 (N_1511,N_789,N_1405);
nand U1512 (N_1512,N_1077,N_1161);
and U1513 (N_1513,N_1257,N_1142);
or U1514 (N_1514,N_892,N_1328);
nand U1515 (N_1515,N_1085,N_1139);
or U1516 (N_1516,N_901,N_1288);
nand U1517 (N_1517,N_1419,N_776);
and U1518 (N_1518,N_1170,N_1307);
nand U1519 (N_1519,N_1332,N_1088);
nor U1520 (N_1520,N_1386,N_1353);
nor U1521 (N_1521,N_1279,N_950);
nor U1522 (N_1522,N_1069,N_1094);
nor U1523 (N_1523,N_833,N_873);
nor U1524 (N_1524,N_1424,N_1377);
xnor U1525 (N_1525,N_1123,N_1402);
nor U1526 (N_1526,N_1076,N_1231);
and U1527 (N_1527,N_1205,N_785);
nand U1528 (N_1528,N_955,N_999);
or U1529 (N_1529,N_1201,N_1167);
or U1530 (N_1530,N_1103,N_1152);
xor U1531 (N_1531,N_1482,N_1388);
or U1532 (N_1532,N_1035,N_1158);
nand U1533 (N_1533,N_932,N_918);
nand U1534 (N_1534,N_1130,N_1284);
and U1535 (N_1535,N_1271,N_751);
or U1536 (N_1536,N_1050,N_1412);
and U1537 (N_1537,N_1349,N_890);
nand U1538 (N_1538,N_1404,N_1222);
nand U1539 (N_1539,N_1121,N_973);
xor U1540 (N_1540,N_1255,N_1453);
nand U1541 (N_1541,N_1499,N_1055);
nand U1542 (N_1542,N_753,N_1071);
or U1543 (N_1543,N_1031,N_1192);
or U1544 (N_1544,N_1135,N_957);
nor U1545 (N_1545,N_1263,N_989);
nor U1546 (N_1546,N_1022,N_1163);
nor U1547 (N_1547,N_757,N_1393);
and U1548 (N_1548,N_883,N_756);
or U1549 (N_1549,N_1376,N_1193);
and U1550 (N_1550,N_1299,N_1045);
or U1551 (N_1551,N_1373,N_1477);
or U1552 (N_1552,N_1278,N_1370);
nor U1553 (N_1553,N_900,N_1274);
nor U1554 (N_1554,N_1308,N_1146);
nor U1555 (N_1555,N_1294,N_1430);
or U1556 (N_1556,N_1232,N_1074);
nand U1557 (N_1557,N_1443,N_1003);
and U1558 (N_1558,N_956,N_966);
and U1559 (N_1559,N_1415,N_835);
nor U1560 (N_1560,N_1410,N_803);
nor U1561 (N_1561,N_1454,N_1208);
or U1562 (N_1562,N_878,N_947);
and U1563 (N_1563,N_1262,N_1431);
nor U1564 (N_1564,N_1138,N_1089);
or U1565 (N_1565,N_1168,N_851);
nand U1566 (N_1566,N_983,N_786);
nand U1567 (N_1567,N_880,N_1204);
or U1568 (N_1568,N_1224,N_1064);
or U1569 (N_1569,N_1114,N_929);
nand U1570 (N_1570,N_903,N_1185);
nand U1571 (N_1571,N_1378,N_959);
and U1572 (N_1572,N_1381,N_1399);
nand U1573 (N_1573,N_1119,N_1361);
nand U1574 (N_1574,N_1438,N_933);
nand U1575 (N_1575,N_1061,N_1259);
xnor U1576 (N_1576,N_1156,N_1368);
nand U1577 (N_1577,N_1417,N_870);
nand U1578 (N_1578,N_1219,N_1024);
and U1579 (N_1579,N_779,N_1488);
nor U1580 (N_1580,N_1266,N_927);
nor U1581 (N_1581,N_807,N_1129);
nor U1582 (N_1582,N_931,N_781);
xnor U1583 (N_1583,N_1437,N_1322);
and U1584 (N_1584,N_1043,N_1040);
or U1585 (N_1585,N_1102,N_1218);
or U1586 (N_1586,N_1075,N_1009);
nand U1587 (N_1587,N_846,N_1112);
or U1588 (N_1588,N_904,N_1481);
and U1589 (N_1589,N_1101,N_1291);
and U1590 (N_1590,N_836,N_1293);
nand U1591 (N_1591,N_1418,N_1466);
and U1592 (N_1592,N_1242,N_1362);
and U1593 (N_1593,N_839,N_1046);
and U1594 (N_1594,N_1127,N_1044);
nor U1595 (N_1595,N_1159,N_1191);
nor U1596 (N_1596,N_954,N_930);
xnor U1597 (N_1597,N_1389,N_1305);
nor U1598 (N_1598,N_849,N_1382);
and U1599 (N_1599,N_830,N_912);
and U1600 (N_1600,N_1295,N_969);
nand U1601 (N_1601,N_790,N_1214);
and U1602 (N_1602,N_822,N_1058);
nor U1603 (N_1603,N_1057,N_1011);
and U1604 (N_1604,N_818,N_1326);
nor U1605 (N_1605,N_1487,N_1248);
nand U1606 (N_1606,N_1317,N_917);
or U1607 (N_1607,N_824,N_943);
and U1608 (N_1608,N_1027,N_1400);
or U1609 (N_1609,N_1091,N_1392);
nand U1610 (N_1610,N_1070,N_872);
nor U1611 (N_1611,N_763,N_1169);
or U1612 (N_1612,N_1426,N_1314);
nand U1613 (N_1613,N_1273,N_825);
nand U1614 (N_1614,N_971,N_1434);
and U1615 (N_1615,N_1463,N_1079);
and U1616 (N_1616,N_895,N_850);
and U1617 (N_1617,N_774,N_1017);
or U1618 (N_1618,N_1313,N_1408);
xor U1619 (N_1619,N_936,N_1136);
or U1620 (N_1620,N_1092,N_964);
nand U1621 (N_1621,N_1436,N_1491);
or U1622 (N_1622,N_1217,N_1403);
or U1623 (N_1623,N_962,N_1197);
and U1624 (N_1624,N_1207,N_1090);
nor U1625 (N_1625,N_1281,N_772);
nand U1626 (N_1626,N_1028,N_804);
or U1627 (N_1627,N_847,N_908);
or U1628 (N_1628,N_1254,N_1211);
and U1629 (N_1629,N_1025,N_1387);
nor U1630 (N_1630,N_793,N_843);
or U1631 (N_1631,N_1447,N_1184);
nor U1632 (N_1632,N_784,N_1369);
and U1633 (N_1633,N_1264,N_911);
nand U1634 (N_1634,N_902,N_1016);
nand U1635 (N_1635,N_907,N_1265);
nor U1636 (N_1636,N_1323,N_1343);
and U1637 (N_1637,N_1344,N_1287);
and U1638 (N_1638,N_1486,N_991);
nand U1639 (N_1639,N_1355,N_1199);
nand U1640 (N_1640,N_1238,N_1150);
and U1641 (N_1641,N_1056,N_1173);
nor U1642 (N_1642,N_965,N_1132);
nand U1643 (N_1643,N_1124,N_1128);
nand U1644 (N_1644,N_1458,N_1366);
and U1645 (N_1645,N_1104,N_1483);
xnor U1646 (N_1646,N_993,N_970);
or U1647 (N_1647,N_817,N_820);
or U1648 (N_1648,N_1126,N_975);
or U1649 (N_1649,N_1029,N_1423);
or U1650 (N_1650,N_1367,N_1496);
or U1651 (N_1651,N_1428,N_1144);
and U1652 (N_1652,N_1452,N_968);
or U1653 (N_1653,N_1448,N_762);
nand U1654 (N_1654,N_1109,N_1223);
or U1655 (N_1655,N_1117,N_1106);
and U1656 (N_1656,N_1320,N_1449);
nand U1657 (N_1657,N_888,N_875);
nand U1658 (N_1658,N_865,N_1020);
nand U1659 (N_1659,N_1479,N_1236);
or U1660 (N_1660,N_1472,N_859);
nand U1661 (N_1661,N_1286,N_1176);
nand U1662 (N_1662,N_1283,N_986);
nand U1663 (N_1663,N_1422,N_794);
and U1664 (N_1664,N_831,N_1162);
nand U1665 (N_1665,N_1107,N_1394);
and U1666 (N_1666,N_760,N_979);
nor U1667 (N_1667,N_1354,N_1267);
or U1668 (N_1668,N_915,N_1351);
and U1669 (N_1669,N_1416,N_788);
and U1670 (N_1670,N_868,N_1336);
or U1671 (N_1671,N_990,N_1441);
nand U1672 (N_1672,N_1047,N_1060);
nand U1673 (N_1673,N_1258,N_1494);
nand U1674 (N_1674,N_778,N_1067);
or U1675 (N_1675,N_860,N_1334);
nand U1676 (N_1676,N_893,N_886);
or U1677 (N_1677,N_981,N_1245);
nand U1678 (N_1678,N_1084,N_1301);
nor U1679 (N_1679,N_1350,N_1374);
nor U1680 (N_1680,N_1203,N_1183);
nor U1681 (N_1681,N_1165,N_1498);
and U1682 (N_1682,N_1316,N_1237);
nand U1683 (N_1683,N_1233,N_945);
nand U1684 (N_1684,N_940,N_769);
or U1685 (N_1685,N_1311,N_921);
nor U1686 (N_1686,N_1110,N_1469);
nor U1687 (N_1687,N_827,N_1006);
nor U1688 (N_1688,N_812,N_791);
nand U1689 (N_1689,N_1310,N_1425);
nand U1690 (N_1690,N_1053,N_1181);
and U1691 (N_1691,N_909,N_1246);
and U1692 (N_1692,N_1345,N_840);
nand U1693 (N_1693,N_815,N_1172);
and U1694 (N_1694,N_1166,N_754);
nor U1695 (N_1695,N_814,N_1134);
or U1696 (N_1696,N_806,N_1083);
nor U1697 (N_1697,N_829,N_925);
nand U1698 (N_1698,N_808,N_1113);
nor U1699 (N_1699,N_934,N_1296);
nand U1700 (N_1700,N_1190,N_1082);
or U1701 (N_1701,N_998,N_1234);
nand U1702 (N_1702,N_764,N_1474);
and U1703 (N_1703,N_1215,N_1038);
or U1704 (N_1704,N_1356,N_1140);
and U1705 (N_1705,N_1312,N_1391);
or U1706 (N_1706,N_1010,N_1118);
or U1707 (N_1707,N_1461,N_1068);
and U1708 (N_1708,N_1072,N_802);
nand U1709 (N_1709,N_952,N_1309);
nor U1710 (N_1710,N_1227,N_1340);
or U1711 (N_1711,N_798,N_1013);
nor U1712 (N_1712,N_1493,N_1225);
nor U1713 (N_1713,N_1413,N_1145);
nor U1714 (N_1714,N_792,N_1383);
nand U1715 (N_1715,N_980,N_1209);
nor U1716 (N_1716,N_1052,N_1002);
nor U1717 (N_1717,N_1034,N_838);
and U1718 (N_1718,N_987,N_1063);
nand U1719 (N_1719,N_863,N_899);
nor U1720 (N_1720,N_1252,N_988);
and U1721 (N_1721,N_1086,N_1042);
nand U1722 (N_1722,N_996,N_1253);
and U1723 (N_1723,N_1008,N_1155);
nor U1724 (N_1724,N_914,N_963);
and U1725 (N_1725,N_1188,N_920);
nor U1726 (N_1726,N_832,N_1427);
nor U1727 (N_1727,N_967,N_1276);
nor U1728 (N_1728,N_877,N_871);
nor U1729 (N_1729,N_1235,N_978);
or U1730 (N_1730,N_891,N_1137);
nand U1731 (N_1731,N_995,N_1151);
and U1732 (N_1732,N_1303,N_1442);
nand U1733 (N_1733,N_1212,N_1359);
nand U1734 (N_1734,N_1048,N_1380);
or U1735 (N_1735,N_1465,N_1032);
or U1736 (N_1736,N_801,N_1304);
or U1737 (N_1737,N_1014,N_816);
or U1738 (N_1738,N_857,N_1339);
xnor U1739 (N_1739,N_755,N_800);
nor U1740 (N_1740,N_1347,N_1357);
nand U1741 (N_1741,N_910,N_811);
or U1742 (N_1742,N_1318,N_767);
and U1743 (N_1743,N_922,N_1363);
xor U1744 (N_1744,N_1122,N_897);
nor U1745 (N_1745,N_1398,N_1297);
nand U1746 (N_1746,N_787,N_982);
or U1747 (N_1747,N_1490,N_1021);
and U1748 (N_1748,N_1471,N_1189);
or U1749 (N_1749,N_1030,N_1105);
nand U1750 (N_1750,N_1462,N_977);
nor U1751 (N_1751,N_919,N_1330);
nand U1752 (N_1752,N_1226,N_1179);
nor U1753 (N_1753,N_1484,N_759);
nor U1754 (N_1754,N_1379,N_1247);
and U1755 (N_1755,N_1000,N_1187);
or U1756 (N_1756,N_1433,N_1240);
and U1757 (N_1757,N_1275,N_1435);
nor U1758 (N_1758,N_923,N_885);
and U1759 (N_1759,N_841,N_1100);
or U1760 (N_1760,N_1450,N_819);
and U1761 (N_1761,N_854,N_1116);
and U1762 (N_1762,N_768,N_972);
and U1763 (N_1763,N_1375,N_976);
and U1764 (N_1764,N_1012,N_1489);
nor U1765 (N_1765,N_848,N_1459);
nor U1766 (N_1766,N_1302,N_942);
nand U1767 (N_1767,N_1154,N_821);
and U1768 (N_1768,N_770,N_939);
nand U1769 (N_1769,N_974,N_958);
nor U1770 (N_1770,N_1251,N_926);
or U1771 (N_1771,N_1041,N_896);
or U1772 (N_1772,N_935,N_1337);
xor U1773 (N_1773,N_1473,N_1321);
or U1774 (N_1774,N_782,N_1365);
nand U1775 (N_1775,N_997,N_869);
nand U1776 (N_1776,N_765,N_1464);
nor U1777 (N_1777,N_861,N_1243);
or U1778 (N_1778,N_845,N_905);
and U1779 (N_1779,N_1148,N_1411);
or U1780 (N_1780,N_826,N_1023);
and U1781 (N_1781,N_1371,N_1244);
or U1782 (N_1782,N_1470,N_1319);
or U1783 (N_1783,N_960,N_941);
and U1784 (N_1784,N_876,N_913);
or U1785 (N_1785,N_1198,N_1290);
nand U1786 (N_1786,N_949,N_1282);
or U1787 (N_1787,N_1335,N_889);
nand U1788 (N_1788,N_1325,N_1213);
nand U1789 (N_1789,N_1397,N_879);
nor U1790 (N_1790,N_1439,N_1115);
or U1791 (N_1791,N_1015,N_1099);
and U1792 (N_1792,N_813,N_780);
or U1793 (N_1793,N_1171,N_881);
xor U1794 (N_1794,N_1327,N_809);
and U1795 (N_1795,N_862,N_1005);
or U1796 (N_1796,N_1401,N_1338);
or U1797 (N_1797,N_1007,N_1352);
nor U1798 (N_1798,N_866,N_985);
nand U1799 (N_1799,N_834,N_1406);
or U1800 (N_1800,N_1241,N_1414);
nand U1801 (N_1801,N_1059,N_1432);
nand U1802 (N_1802,N_1270,N_1261);
nand U1803 (N_1803,N_1078,N_1065);
nand U1804 (N_1804,N_1456,N_1256);
or U1805 (N_1805,N_1429,N_1306);
or U1806 (N_1806,N_1125,N_858);
or U1807 (N_1807,N_1485,N_1093);
or U1808 (N_1808,N_810,N_1206);
and U1809 (N_1809,N_1131,N_1157);
or U1810 (N_1810,N_823,N_1186);
nor U1811 (N_1811,N_1495,N_1087);
or U1812 (N_1812,N_894,N_1037);
or U1813 (N_1813,N_1097,N_1174);
nor U1814 (N_1814,N_1229,N_1269);
nand U1815 (N_1815,N_758,N_1285);
or U1816 (N_1816,N_1348,N_837);
nor U1817 (N_1817,N_1396,N_1324);
xor U1818 (N_1818,N_882,N_842);
nand U1819 (N_1819,N_898,N_1341);
and U1820 (N_1820,N_1120,N_1360);
nor U1821 (N_1821,N_1164,N_1384);
or U1822 (N_1822,N_1149,N_1298);
or U1823 (N_1823,N_874,N_946);
or U1824 (N_1824,N_1409,N_1289);
nand U1825 (N_1825,N_1451,N_1468);
nor U1826 (N_1826,N_1062,N_906);
nand U1827 (N_1827,N_961,N_750);
nor U1828 (N_1828,N_1445,N_1210);
or U1829 (N_1829,N_1026,N_799);
or U1830 (N_1830,N_853,N_1004);
nor U1831 (N_1831,N_953,N_1280);
and U1832 (N_1832,N_1478,N_994);
or U1833 (N_1833,N_1033,N_1292);
and U1834 (N_1834,N_1141,N_1178);
and U1835 (N_1835,N_1228,N_777);
nor U1836 (N_1836,N_1420,N_1018);
nor U1837 (N_1837,N_1180,N_1364);
nand U1838 (N_1838,N_1230,N_916);
or U1839 (N_1839,N_1331,N_1073);
and U1840 (N_1840,N_1098,N_984);
or U1841 (N_1841,N_1143,N_1390);
xor U1842 (N_1842,N_867,N_1177);
or U1843 (N_1843,N_1385,N_1315);
or U1844 (N_1844,N_1346,N_1444);
and U1845 (N_1845,N_1457,N_1300);
nand U1846 (N_1846,N_1196,N_1455);
nand U1847 (N_1847,N_924,N_1175);
xnor U1848 (N_1848,N_1036,N_1108);
and U1849 (N_1849,N_1421,N_1160);
or U1850 (N_1850,N_1194,N_937);
or U1851 (N_1851,N_1329,N_1019);
xnor U1852 (N_1852,N_1492,N_771);
nand U1853 (N_1853,N_1147,N_1460);
nor U1854 (N_1854,N_775,N_1001);
nor U1855 (N_1855,N_1333,N_1407);
nand U1856 (N_1856,N_1358,N_1195);
and U1857 (N_1857,N_1096,N_855);
nor U1858 (N_1858,N_1342,N_1249);
nand U1859 (N_1859,N_828,N_1395);
or U1860 (N_1860,N_1066,N_852);
and U1861 (N_1861,N_1133,N_796);
and U1862 (N_1862,N_1200,N_1467);
nand U1863 (N_1863,N_864,N_951);
or U1864 (N_1864,N_1095,N_1080);
and U1865 (N_1865,N_884,N_783);
and U1866 (N_1866,N_1220,N_1221);
nor U1867 (N_1867,N_1260,N_856);
nand U1868 (N_1868,N_797,N_1081);
nor U1869 (N_1869,N_795,N_773);
nor U1870 (N_1870,N_887,N_1372);
nand U1871 (N_1871,N_1239,N_752);
and U1872 (N_1872,N_1480,N_1272);
and U1873 (N_1873,N_1153,N_1111);
or U1874 (N_1874,N_1216,N_1054);
and U1875 (N_1875,N_1333,N_1151);
nor U1876 (N_1876,N_1465,N_1304);
nand U1877 (N_1877,N_1143,N_957);
or U1878 (N_1878,N_900,N_949);
and U1879 (N_1879,N_1125,N_1053);
nand U1880 (N_1880,N_984,N_1022);
or U1881 (N_1881,N_1417,N_914);
nand U1882 (N_1882,N_766,N_1373);
nand U1883 (N_1883,N_756,N_1389);
and U1884 (N_1884,N_1058,N_848);
or U1885 (N_1885,N_1469,N_1310);
nand U1886 (N_1886,N_1111,N_1054);
and U1887 (N_1887,N_1438,N_1357);
or U1888 (N_1888,N_972,N_1087);
nand U1889 (N_1889,N_928,N_1499);
nor U1890 (N_1890,N_1438,N_1356);
or U1891 (N_1891,N_1372,N_1394);
and U1892 (N_1892,N_1028,N_809);
nor U1893 (N_1893,N_1316,N_1012);
or U1894 (N_1894,N_916,N_974);
and U1895 (N_1895,N_1266,N_840);
nor U1896 (N_1896,N_1092,N_1468);
or U1897 (N_1897,N_1109,N_1046);
nor U1898 (N_1898,N_1014,N_1444);
and U1899 (N_1899,N_1202,N_1159);
and U1900 (N_1900,N_1144,N_785);
nor U1901 (N_1901,N_1155,N_1481);
and U1902 (N_1902,N_1478,N_1114);
nand U1903 (N_1903,N_939,N_1401);
xnor U1904 (N_1904,N_1024,N_1361);
nand U1905 (N_1905,N_1348,N_1163);
nand U1906 (N_1906,N_859,N_1292);
and U1907 (N_1907,N_1268,N_1196);
nor U1908 (N_1908,N_1472,N_1345);
and U1909 (N_1909,N_1015,N_1165);
nand U1910 (N_1910,N_1298,N_1137);
nand U1911 (N_1911,N_798,N_873);
nor U1912 (N_1912,N_1469,N_932);
nand U1913 (N_1913,N_1092,N_1355);
nand U1914 (N_1914,N_873,N_946);
nor U1915 (N_1915,N_942,N_1321);
and U1916 (N_1916,N_1192,N_1201);
nor U1917 (N_1917,N_1440,N_1386);
and U1918 (N_1918,N_1378,N_905);
or U1919 (N_1919,N_955,N_905);
or U1920 (N_1920,N_1352,N_1436);
nand U1921 (N_1921,N_835,N_1060);
and U1922 (N_1922,N_1178,N_930);
or U1923 (N_1923,N_1204,N_1155);
nor U1924 (N_1924,N_788,N_1213);
nand U1925 (N_1925,N_946,N_1095);
nand U1926 (N_1926,N_1016,N_810);
or U1927 (N_1927,N_1120,N_1416);
and U1928 (N_1928,N_1229,N_873);
nand U1929 (N_1929,N_1444,N_1211);
nor U1930 (N_1930,N_793,N_1060);
nor U1931 (N_1931,N_795,N_1076);
nand U1932 (N_1932,N_1295,N_771);
nor U1933 (N_1933,N_1468,N_1284);
and U1934 (N_1934,N_823,N_1033);
nand U1935 (N_1935,N_1057,N_802);
nor U1936 (N_1936,N_1081,N_930);
and U1937 (N_1937,N_969,N_1378);
nand U1938 (N_1938,N_1287,N_1075);
or U1939 (N_1939,N_986,N_1030);
nor U1940 (N_1940,N_1372,N_934);
nor U1941 (N_1941,N_1305,N_1113);
nor U1942 (N_1942,N_1486,N_1061);
and U1943 (N_1943,N_848,N_1311);
and U1944 (N_1944,N_1318,N_880);
nor U1945 (N_1945,N_896,N_854);
or U1946 (N_1946,N_798,N_1385);
nand U1947 (N_1947,N_951,N_1164);
nand U1948 (N_1948,N_1261,N_1168);
and U1949 (N_1949,N_1028,N_861);
or U1950 (N_1950,N_1040,N_1352);
or U1951 (N_1951,N_1092,N_1157);
and U1952 (N_1952,N_1322,N_929);
nor U1953 (N_1953,N_1407,N_1467);
and U1954 (N_1954,N_979,N_1021);
nor U1955 (N_1955,N_839,N_1358);
nor U1956 (N_1956,N_1425,N_1239);
nand U1957 (N_1957,N_1259,N_995);
or U1958 (N_1958,N_1012,N_1043);
or U1959 (N_1959,N_1355,N_1446);
or U1960 (N_1960,N_1449,N_811);
nor U1961 (N_1961,N_981,N_1418);
nor U1962 (N_1962,N_1355,N_982);
and U1963 (N_1963,N_1139,N_948);
nand U1964 (N_1964,N_1243,N_1282);
or U1965 (N_1965,N_1459,N_1052);
or U1966 (N_1966,N_1162,N_836);
nor U1967 (N_1967,N_1310,N_1389);
xnor U1968 (N_1968,N_1383,N_1060);
nand U1969 (N_1969,N_973,N_1037);
and U1970 (N_1970,N_876,N_1383);
or U1971 (N_1971,N_1184,N_1397);
or U1972 (N_1972,N_898,N_1416);
nor U1973 (N_1973,N_834,N_1373);
nor U1974 (N_1974,N_1142,N_1367);
and U1975 (N_1975,N_757,N_915);
and U1976 (N_1976,N_1434,N_1395);
nor U1977 (N_1977,N_1442,N_1280);
nor U1978 (N_1978,N_933,N_874);
nor U1979 (N_1979,N_1121,N_981);
nand U1980 (N_1980,N_1235,N_1471);
or U1981 (N_1981,N_806,N_1427);
nor U1982 (N_1982,N_1299,N_785);
and U1983 (N_1983,N_1075,N_1480);
and U1984 (N_1984,N_1405,N_859);
nor U1985 (N_1985,N_1116,N_1019);
xor U1986 (N_1986,N_1249,N_1130);
and U1987 (N_1987,N_1344,N_1318);
nand U1988 (N_1988,N_960,N_1385);
and U1989 (N_1989,N_1325,N_929);
and U1990 (N_1990,N_762,N_1406);
and U1991 (N_1991,N_904,N_1449);
and U1992 (N_1992,N_870,N_923);
and U1993 (N_1993,N_1356,N_1302);
nor U1994 (N_1994,N_1081,N_1042);
nand U1995 (N_1995,N_1402,N_1133);
nor U1996 (N_1996,N_816,N_988);
nor U1997 (N_1997,N_862,N_885);
and U1998 (N_1998,N_1375,N_1490);
nor U1999 (N_1999,N_771,N_783);
nand U2000 (N_2000,N_1285,N_822);
nor U2001 (N_2001,N_1075,N_1219);
and U2002 (N_2002,N_1246,N_1339);
nor U2003 (N_2003,N_834,N_1303);
or U2004 (N_2004,N_1142,N_990);
and U2005 (N_2005,N_1352,N_996);
or U2006 (N_2006,N_950,N_861);
nand U2007 (N_2007,N_958,N_988);
nand U2008 (N_2008,N_1372,N_1255);
nor U2009 (N_2009,N_779,N_1351);
or U2010 (N_2010,N_823,N_1107);
nor U2011 (N_2011,N_1431,N_1347);
nor U2012 (N_2012,N_809,N_1431);
xnor U2013 (N_2013,N_821,N_1341);
and U2014 (N_2014,N_1084,N_1012);
nor U2015 (N_2015,N_1327,N_966);
and U2016 (N_2016,N_775,N_1316);
nand U2017 (N_2017,N_1327,N_1125);
nand U2018 (N_2018,N_1017,N_1021);
nand U2019 (N_2019,N_965,N_878);
nor U2020 (N_2020,N_1399,N_1108);
or U2021 (N_2021,N_821,N_1261);
or U2022 (N_2022,N_1259,N_1346);
and U2023 (N_2023,N_1264,N_781);
nand U2024 (N_2024,N_1497,N_1108);
nand U2025 (N_2025,N_1194,N_1299);
nor U2026 (N_2026,N_1138,N_1206);
or U2027 (N_2027,N_1361,N_870);
or U2028 (N_2028,N_1169,N_796);
xor U2029 (N_2029,N_1108,N_1325);
nand U2030 (N_2030,N_1248,N_880);
nand U2031 (N_2031,N_1409,N_1233);
or U2032 (N_2032,N_831,N_1373);
nand U2033 (N_2033,N_817,N_973);
or U2034 (N_2034,N_1027,N_1352);
or U2035 (N_2035,N_1315,N_1310);
and U2036 (N_2036,N_885,N_1470);
nor U2037 (N_2037,N_1014,N_1244);
and U2038 (N_2038,N_769,N_1144);
and U2039 (N_2039,N_922,N_755);
nand U2040 (N_2040,N_1087,N_1461);
or U2041 (N_2041,N_1444,N_1013);
and U2042 (N_2042,N_1409,N_1013);
and U2043 (N_2043,N_847,N_1140);
or U2044 (N_2044,N_1393,N_1354);
xnor U2045 (N_2045,N_1152,N_1170);
or U2046 (N_2046,N_750,N_1429);
nand U2047 (N_2047,N_1207,N_1325);
nor U2048 (N_2048,N_1091,N_1423);
or U2049 (N_2049,N_937,N_810);
nor U2050 (N_2050,N_1193,N_801);
and U2051 (N_2051,N_980,N_821);
and U2052 (N_2052,N_1258,N_1196);
and U2053 (N_2053,N_906,N_1041);
nor U2054 (N_2054,N_788,N_1497);
and U2055 (N_2055,N_884,N_1212);
nand U2056 (N_2056,N_1356,N_770);
nand U2057 (N_2057,N_1301,N_1011);
nor U2058 (N_2058,N_1487,N_819);
nand U2059 (N_2059,N_971,N_1458);
nor U2060 (N_2060,N_1275,N_1074);
nor U2061 (N_2061,N_809,N_1259);
or U2062 (N_2062,N_1294,N_1318);
nand U2063 (N_2063,N_1308,N_931);
and U2064 (N_2064,N_965,N_889);
nand U2065 (N_2065,N_1333,N_1394);
nor U2066 (N_2066,N_1153,N_1000);
nor U2067 (N_2067,N_1445,N_1318);
and U2068 (N_2068,N_1285,N_1301);
or U2069 (N_2069,N_1042,N_1335);
and U2070 (N_2070,N_1155,N_999);
nor U2071 (N_2071,N_1083,N_1466);
nor U2072 (N_2072,N_1148,N_929);
or U2073 (N_2073,N_1341,N_1252);
nor U2074 (N_2074,N_1010,N_917);
nor U2075 (N_2075,N_1024,N_1180);
nand U2076 (N_2076,N_1336,N_1237);
nand U2077 (N_2077,N_759,N_1000);
nor U2078 (N_2078,N_1476,N_1419);
nor U2079 (N_2079,N_1276,N_828);
and U2080 (N_2080,N_1338,N_789);
and U2081 (N_2081,N_1134,N_1185);
and U2082 (N_2082,N_1393,N_988);
and U2083 (N_2083,N_1163,N_1496);
nand U2084 (N_2084,N_947,N_759);
and U2085 (N_2085,N_1481,N_1176);
and U2086 (N_2086,N_1406,N_1215);
nand U2087 (N_2087,N_953,N_1358);
nand U2088 (N_2088,N_1182,N_1113);
nand U2089 (N_2089,N_1391,N_1161);
or U2090 (N_2090,N_1352,N_1270);
and U2091 (N_2091,N_1225,N_1070);
nor U2092 (N_2092,N_1029,N_1231);
nand U2093 (N_2093,N_1372,N_1042);
and U2094 (N_2094,N_1389,N_1450);
nor U2095 (N_2095,N_1273,N_978);
nor U2096 (N_2096,N_879,N_1237);
or U2097 (N_2097,N_957,N_1234);
xnor U2098 (N_2098,N_1253,N_858);
xor U2099 (N_2099,N_1098,N_788);
and U2100 (N_2100,N_995,N_1381);
nor U2101 (N_2101,N_929,N_788);
nor U2102 (N_2102,N_1327,N_752);
and U2103 (N_2103,N_1061,N_1065);
or U2104 (N_2104,N_1265,N_1196);
nand U2105 (N_2105,N_1486,N_864);
nand U2106 (N_2106,N_763,N_1159);
nand U2107 (N_2107,N_1354,N_1062);
nand U2108 (N_2108,N_1382,N_881);
xor U2109 (N_2109,N_1358,N_1257);
and U2110 (N_2110,N_1016,N_876);
or U2111 (N_2111,N_1169,N_1313);
or U2112 (N_2112,N_1285,N_1354);
and U2113 (N_2113,N_1496,N_938);
nor U2114 (N_2114,N_844,N_811);
nor U2115 (N_2115,N_1160,N_1082);
nor U2116 (N_2116,N_1117,N_1046);
and U2117 (N_2117,N_997,N_1478);
and U2118 (N_2118,N_1207,N_1378);
or U2119 (N_2119,N_1110,N_877);
or U2120 (N_2120,N_1388,N_769);
or U2121 (N_2121,N_1497,N_856);
and U2122 (N_2122,N_1473,N_1073);
nor U2123 (N_2123,N_898,N_1043);
and U2124 (N_2124,N_763,N_970);
nor U2125 (N_2125,N_1044,N_839);
or U2126 (N_2126,N_1214,N_1216);
or U2127 (N_2127,N_896,N_764);
and U2128 (N_2128,N_1427,N_908);
nand U2129 (N_2129,N_1202,N_1157);
nor U2130 (N_2130,N_750,N_1213);
nand U2131 (N_2131,N_817,N_940);
nand U2132 (N_2132,N_1417,N_937);
nor U2133 (N_2133,N_1301,N_995);
nor U2134 (N_2134,N_1181,N_1298);
or U2135 (N_2135,N_1159,N_877);
nor U2136 (N_2136,N_794,N_1257);
nor U2137 (N_2137,N_1271,N_1269);
nor U2138 (N_2138,N_966,N_1249);
or U2139 (N_2139,N_1178,N_1408);
and U2140 (N_2140,N_1376,N_868);
or U2141 (N_2141,N_751,N_925);
xnor U2142 (N_2142,N_1154,N_1292);
or U2143 (N_2143,N_899,N_1436);
and U2144 (N_2144,N_917,N_826);
and U2145 (N_2145,N_1459,N_1018);
and U2146 (N_2146,N_1003,N_761);
nor U2147 (N_2147,N_766,N_1006);
nor U2148 (N_2148,N_947,N_1288);
or U2149 (N_2149,N_866,N_1235);
and U2150 (N_2150,N_844,N_925);
and U2151 (N_2151,N_1095,N_1458);
nand U2152 (N_2152,N_1444,N_790);
nand U2153 (N_2153,N_1419,N_1155);
nor U2154 (N_2154,N_1106,N_1399);
nor U2155 (N_2155,N_927,N_1178);
and U2156 (N_2156,N_1493,N_750);
nand U2157 (N_2157,N_903,N_1265);
nor U2158 (N_2158,N_1349,N_1222);
nor U2159 (N_2159,N_1149,N_877);
and U2160 (N_2160,N_1090,N_1079);
nor U2161 (N_2161,N_762,N_916);
nand U2162 (N_2162,N_804,N_792);
or U2163 (N_2163,N_1425,N_1458);
and U2164 (N_2164,N_1496,N_1395);
nand U2165 (N_2165,N_1002,N_1155);
and U2166 (N_2166,N_1107,N_1140);
nand U2167 (N_2167,N_1013,N_823);
and U2168 (N_2168,N_912,N_1292);
xnor U2169 (N_2169,N_1151,N_812);
and U2170 (N_2170,N_1028,N_820);
nor U2171 (N_2171,N_1081,N_1096);
nor U2172 (N_2172,N_974,N_1476);
nor U2173 (N_2173,N_821,N_864);
nand U2174 (N_2174,N_1330,N_881);
and U2175 (N_2175,N_1116,N_926);
nor U2176 (N_2176,N_1329,N_1098);
nor U2177 (N_2177,N_1433,N_1488);
nand U2178 (N_2178,N_970,N_920);
and U2179 (N_2179,N_1412,N_774);
nand U2180 (N_2180,N_1453,N_1317);
and U2181 (N_2181,N_1389,N_1271);
nor U2182 (N_2182,N_1399,N_825);
nand U2183 (N_2183,N_1129,N_1115);
nand U2184 (N_2184,N_1477,N_793);
nand U2185 (N_2185,N_912,N_1037);
nor U2186 (N_2186,N_1380,N_1460);
nor U2187 (N_2187,N_1236,N_997);
nand U2188 (N_2188,N_769,N_1358);
and U2189 (N_2189,N_1351,N_1499);
and U2190 (N_2190,N_1207,N_945);
or U2191 (N_2191,N_1291,N_777);
or U2192 (N_2192,N_1497,N_1168);
nor U2193 (N_2193,N_958,N_795);
nor U2194 (N_2194,N_1151,N_1279);
or U2195 (N_2195,N_865,N_1362);
or U2196 (N_2196,N_1239,N_1224);
and U2197 (N_2197,N_1299,N_1370);
and U2198 (N_2198,N_814,N_853);
nor U2199 (N_2199,N_1012,N_1275);
and U2200 (N_2200,N_1336,N_999);
nand U2201 (N_2201,N_820,N_1261);
nand U2202 (N_2202,N_1415,N_1267);
nor U2203 (N_2203,N_1334,N_1283);
and U2204 (N_2204,N_1011,N_1174);
and U2205 (N_2205,N_985,N_1314);
nand U2206 (N_2206,N_968,N_785);
or U2207 (N_2207,N_1015,N_931);
nor U2208 (N_2208,N_873,N_1208);
or U2209 (N_2209,N_1148,N_754);
or U2210 (N_2210,N_1471,N_870);
and U2211 (N_2211,N_1496,N_1157);
or U2212 (N_2212,N_853,N_1385);
and U2213 (N_2213,N_1087,N_825);
nor U2214 (N_2214,N_750,N_1457);
nand U2215 (N_2215,N_1152,N_1470);
nand U2216 (N_2216,N_903,N_1462);
and U2217 (N_2217,N_1414,N_1210);
nor U2218 (N_2218,N_1012,N_752);
and U2219 (N_2219,N_833,N_1296);
or U2220 (N_2220,N_1162,N_1250);
and U2221 (N_2221,N_1176,N_878);
nand U2222 (N_2222,N_1117,N_1369);
nor U2223 (N_2223,N_767,N_816);
nor U2224 (N_2224,N_1348,N_1171);
and U2225 (N_2225,N_918,N_1338);
and U2226 (N_2226,N_887,N_1244);
and U2227 (N_2227,N_1185,N_1244);
nand U2228 (N_2228,N_1162,N_898);
nand U2229 (N_2229,N_1063,N_969);
nand U2230 (N_2230,N_1065,N_1191);
nand U2231 (N_2231,N_1098,N_1017);
or U2232 (N_2232,N_1277,N_1211);
xor U2233 (N_2233,N_1108,N_908);
nor U2234 (N_2234,N_1458,N_1014);
nor U2235 (N_2235,N_835,N_1057);
nand U2236 (N_2236,N_914,N_1037);
nand U2237 (N_2237,N_1390,N_1031);
xor U2238 (N_2238,N_1301,N_1091);
nand U2239 (N_2239,N_882,N_1294);
nor U2240 (N_2240,N_1490,N_1340);
nand U2241 (N_2241,N_1481,N_812);
and U2242 (N_2242,N_884,N_1451);
nor U2243 (N_2243,N_1002,N_759);
nor U2244 (N_2244,N_1225,N_1446);
nor U2245 (N_2245,N_820,N_818);
nand U2246 (N_2246,N_857,N_1221);
or U2247 (N_2247,N_1160,N_883);
nor U2248 (N_2248,N_1474,N_765);
nand U2249 (N_2249,N_996,N_912);
and U2250 (N_2250,N_1791,N_1796);
nand U2251 (N_2251,N_2102,N_2214);
nand U2252 (N_2252,N_1529,N_1825);
or U2253 (N_2253,N_2031,N_1827);
or U2254 (N_2254,N_2090,N_2139);
nor U2255 (N_2255,N_1870,N_1808);
nor U2256 (N_2256,N_1832,N_2201);
nand U2257 (N_2257,N_1842,N_1591);
nor U2258 (N_2258,N_1699,N_2147);
nor U2259 (N_2259,N_1918,N_2060);
nand U2260 (N_2260,N_1587,N_1558);
and U2261 (N_2261,N_2081,N_2038);
nand U2262 (N_2262,N_1505,N_1652);
or U2263 (N_2263,N_1608,N_1867);
and U2264 (N_2264,N_1947,N_1923);
nand U2265 (N_2265,N_1741,N_1506);
xor U2266 (N_2266,N_1628,N_1564);
and U2267 (N_2267,N_1881,N_1801);
nand U2268 (N_2268,N_1758,N_1714);
and U2269 (N_2269,N_1710,N_1908);
and U2270 (N_2270,N_1611,N_1956);
nor U2271 (N_2271,N_2200,N_2198);
or U2272 (N_2272,N_1760,N_1862);
nand U2273 (N_2273,N_1643,N_2046);
nand U2274 (N_2274,N_2162,N_1544);
or U2275 (N_2275,N_2230,N_1865);
nand U2276 (N_2276,N_2173,N_2225);
nand U2277 (N_2277,N_1996,N_1509);
nor U2278 (N_2278,N_1823,N_1902);
nor U2279 (N_2279,N_1594,N_1663);
or U2280 (N_2280,N_1550,N_2219);
and U2281 (N_2281,N_2166,N_2109);
or U2282 (N_2282,N_1915,N_2030);
and U2283 (N_2283,N_1998,N_2110);
nor U2284 (N_2284,N_2236,N_1559);
nand U2285 (N_2285,N_2206,N_2155);
nor U2286 (N_2286,N_1524,N_2182);
nor U2287 (N_2287,N_1621,N_1937);
and U2288 (N_2288,N_1855,N_2144);
or U2289 (N_2289,N_1579,N_1879);
or U2290 (N_2290,N_2177,N_1637);
and U2291 (N_2291,N_1868,N_2159);
nand U2292 (N_2292,N_2044,N_1949);
nand U2293 (N_2293,N_1669,N_1647);
nand U2294 (N_2294,N_1935,N_1964);
nand U2295 (N_2295,N_2004,N_2088);
xnor U2296 (N_2296,N_1546,N_2013);
or U2297 (N_2297,N_2240,N_1955);
nand U2298 (N_2298,N_2249,N_1970);
nor U2299 (N_2299,N_1822,N_2014);
nor U2300 (N_2300,N_1689,N_1685);
nand U2301 (N_2301,N_1981,N_1790);
nand U2302 (N_2302,N_1815,N_1730);
or U2303 (N_2303,N_1703,N_2202);
nor U2304 (N_2304,N_1723,N_1891);
nand U2305 (N_2305,N_1805,N_1986);
nor U2306 (N_2306,N_1838,N_2151);
nor U2307 (N_2307,N_1695,N_1934);
nor U2308 (N_2308,N_1993,N_1531);
or U2309 (N_2309,N_1917,N_1535);
or U2310 (N_2310,N_1510,N_2078);
and U2311 (N_2311,N_2197,N_2073);
nor U2312 (N_2312,N_2191,N_2181);
nand U2313 (N_2313,N_1518,N_2023);
or U2314 (N_2314,N_2185,N_1834);
nor U2315 (N_2315,N_1526,N_1795);
nor U2316 (N_2316,N_1675,N_1907);
and U2317 (N_2317,N_2196,N_1893);
and U2318 (N_2318,N_2231,N_1702);
nand U2319 (N_2319,N_2194,N_1916);
or U2320 (N_2320,N_2132,N_2195);
or U2321 (N_2321,N_2061,N_2216);
and U2322 (N_2322,N_2053,N_1646);
nand U2323 (N_2323,N_1682,N_1761);
nand U2324 (N_2324,N_1926,N_1817);
nand U2325 (N_2325,N_1521,N_2146);
nand U2326 (N_2326,N_2076,N_2150);
nand U2327 (N_2327,N_1977,N_2167);
or U2328 (N_2328,N_1786,N_1708);
nand U2329 (N_2329,N_1751,N_1597);
nor U2330 (N_2330,N_2229,N_1542);
nand U2331 (N_2331,N_2108,N_1869);
or U2332 (N_2332,N_1753,N_1960);
nand U2333 (N_2333,N_2169,N_2158);
and U2334 (N_2334,N_1569,N_1684);
and U2335 (N_2335,N_1604,N_1939);
xor U2336 (N_2336,N_1640,N_1552);
nand U2337 (N_2337,N_2099,N_1545);
nor U2338 (N_2338,N_2089,N_1771);
and U2339 (N_2339,N_1861,N_1779);
or U2340 (N_2340,N_1933,N_1700);
nand U2341 (N_2341,N_2000,N_1895);
or U2342 (N_2342,N_1788,N_1976);
and U2343 (N_2343,N_1729,N_1785);
nand U2344 (N_2344,N_1595,N_1953);
nand U2345 (N_2345,N_2207,N_2141);
or U2346 (N_2346,N_2170,N_1909);
and U2347 (N_2347,N_1987,N_1848);
or U2348 (N_2348,N_1880,N_1719);
and U2349 (N_2349,N_1561,N_1890);
nand U2350 (N_2350,N_1994,N_2039);
nand U2351 (N_2351,N_1605,N_2119);
nor U2352 (N_2352,N_1711,N_2002);
xor U2353 (N_2353,N_1578,N_1807);
and U2354 (N_2354,N_1734,N_1773);
nand U2355 (N_2355,N_1568,N_2103);
nor U2356 (N_2356,N_1876,N_2192);
nor U2357 (N_2357,N_2082,N_1845);
nor U2358 (N_2358,N_1792,N_1585);
nor U2359 (N_2359,N_1522,N_1501);
nor U2360 (N_2360,N_1726,N_1820);
or U2361 (N_2361,N_2024,N_2100);
or U2362 (N_2362,N_2041,N_1793);
nand U2363 (N_2363,N_2105,N_1812);
and U2364 (N_2364,N_2032,N_1588);
nor U2365 (N_2365,N_1577,N_1886);
and U2366 (N_2366,N_1581,N_1846);
nor U2367 (N_2367,N_1500,N_2232);
and U2368 (N_2368,N_2153,N_1938);
or U2369 (N_2369,N_2154,N_1819);
and U2370 (N_2370,N_1540,N_1613);
xor U2371 (N_2371,N_1560,N_2126);
and U2372 (N_2372,N_1698,N_2140);
and U2373 (N_2373,N_2127,N_1728);
nand U2374 (N_2374,N_2084,N_1744);
or U2375 (N_2375,N_1514,N_1810);
nor U2376 (N_2376,N_2069,N_1966);
and U2377 (N_2377,N_1688,N_1547);
nor U2378 (N_2378,N_1538,N_2019);
nand U2379 (N_2379,N_2057,N_2247);
or U2380 (N_2380,N_2163,N_1936);
nand U2381 (N_2381,N_2208,N_1602);
nand U2382 (N_2382,N_2106,N_1694);
and U2383 (N_2383,N_1511,N_1950);
and U2384 (N_2384,N_1818,N_2122);
nor U2385 (N_2385,N_1911,N_1580);
nor U2386 (N_2386,N_1746,N_2209);
nand U2387 (N_2387,N_1696,N_1942);
and U2388 (N_2388,N_2016,N_1571);
nand U2389 (N_2389,N_1553,N_1725);
or U2390 (N_2390,N_1623,N_2222);
and U2391 (N_2391,N_1800,N_1831);
and U2392 (N_2392,N_1783,N_1701);
nand U2393 (N_2393,N_1985,N_1704);
and U2394 (N_2394,N_1864,N_2168);
nand U2395 (N_2395,N_2009,N_2010);
nor U2396 (N_2396,N_1666,N_2025);
or U2397 (N_2397,N_1739,N_1978);
nand U2398 (N_2398,N_2234,N_2221);
or U2399 (N_2399,N_1707,N_2174);
and U2400 (N_2400,N_1821,N_1836);
nor U2401 (N_2401,N_1533,N_1828);
or U2402 (N_2402,N_1554,N_2121);
nor U2403 (N_2403,N_1863,N_1636);
nand U2404 (N_2404,N_1990,N_2008);
nor U2405 (N_2405,N_2080,N_2114);
nor U2406 (N_2406,N_1593,N_1984);
nand U2407 (N_2407,N_2165,N_2098);
and U2408 (N_2408,N_1764,N_1523);
and U2409 (N_2409,N_1948,N_1624);
or U2410 (N_2410,N_1639,N_2130);
nor U2411 (N_2411,N_1654,N_1665);
nand U2412 (N_2412,N_1603,N_1859);
nor U2413 (N_2413,N_1872,N_1616);
and U2414 (N_2414,N_1995,N_2187);
and U2415 (N_2415,N_1768,N_1503);
nor U2416 (N_2416,N_1919,N_1574);
and U2417 (N_2417,N_2071,N_1648);
nor U2418 (N_2418,N_2183,N_2026);
or U2419 (N_2419,N_1770,N_1692);
and U2420 (N_2420,N_2021,N_1617);
nand U2421 (N_2421,N_1532,N_2138);
or U2422 (N_2422,N_1737,N_1724);
nand U2423 (N_2423,N_2148,N_2145);
nand U2424 (N_2424,N_1676,N_1678);
or U2425 (N_2425,N_1612,N_2193);
and U2426 (N_2426,N_1833,N_1709);
nor U2427 (N_2427,N_1759,N_1874);
nor U2428 (N_2428,N_1716,N_2043);
nor U2429 (N_2429,N_2129,N_1809);
nor U2430 (N_2430,N_1903,N_1989);
nand U2431 (N_2431,N_1799,N_1727);
nand U2432 (N_2432,N_2131,N_2094);
nor U2433 (N_2433,N_1814,N_2245);
or U2434 (N_2434,N_2142,N_2005);
or U2435 (N_2435,N_1745,N_2086);
or U2436 (N_2436,N_2212,N_1610);
nand U2437 (N_2437,N_2111,N_2246);
nor U2438 (N_2438,N_1972,N_1672);
or U2439 (N_2439,N_1609,N_2243);
or U2440 (N_2440,N_2028,N_1677);
nor U2441 (N_2441,N_1813,N_1536);
nor U2442 (N_2442,N_1614,N_2156);
and U2443 (N_2443,N_1826,N_2157);
nor U2444 (N_2444,N_2035,N_2067);
or U2445 (N_2445,N_2233,N_1873);
nor U2446 (N_2446,N_1959,N_2050);
or U2447 (N_2447,N_2059,N_1887);
nor U2448 (N_2448,N_1988,N_1757);
nand U2449 (N_2449,N_1854,N_2178);
or U2450 (N_2450,N_2218,N_1635);
and U2451 (N_2451,N_1971,N_2242);
nor U2452 (N_2452,N_1735,N_1858);
nand U2453 (N_2453,N_1525,N_2015);
nand U2454 (N_2454,N_1674,N_2093);
or U2455 (N_2455,N_1920,N_1633);
and U2456 (N_2456,N_1655,N_2143);
and U2457 (N_2457,N_1866,N_1681);
nand U2458 (N_2458,N_1963,N_1962);
nand U2459 (N_2459,N_1997,N_1983);
nand U2460 (N_2460,N_1774,N_1556);
nor U2461 (N_2461,N_1824,N_1668);
or U2462 (N_2462,N_1572,N_1721);
or U2463 (N_2463,N_2115,N_1787);
nor U2464 (N_2464,N_2034,N_1747);
nor U2465 (N_2465,N_1583,N_1650);
nor U2466 (N_2466,N_1932,N_2190);
or U2467 (N_2467,N_1905,N_1769);
or U2468 (N_2468,N_2065,N_2124);
nor U2469 (N_2469,N_1914,N_1537);
and U2470 (N_2470,N_1811,N_1910);
and U2471 (N_2471,N_1508,N_1642);
or U2472 (N_2472,N_2220,N_1857);
or U2473 (N_2473,N_1901,N_1922);
nor U2474 (N_2474,N_1921,N_1924);
and U2475 (N_2475,N_1931,N_2049);
or U2476 (N_2476,N_2052,N_2164);
nand U2477 (N_2477,N_1627,N_1667);
and U2478 (N_2478,N_2226,N_2027);
and U2479 (N_2479,N_2118,N_2179);
nor U2480 (N_2480,N_2123,N_1517);
nor U2481 (N_2481,N_1980,N_2136);
and U2482 (N_2482,N_1968,N_1849);
nand U2483 (N_2483,N_1664,N_2228);
nor U2484 (N_2484,N_2215,N_1992);
and U2485 (N_2485,N_1954,N_2075);
or U2486 (N_2486,N_1898,N_1686);
and U2487 (N_2487,N_2244,N_1806);
nor U2488 (N_2488,N_2020,N_1816);
nor U2489 (N_2489,N_1530,N_2188);
or U2490 (N_2490,N_2092,N_2006);
nand U2491 (N_2491,N_1892,N_1776);
nand U2492 (N_2492,N_1875,N_1925);
or U2493 (N_2493,N_1748,N_1638);
and U2494 (N_2494,N_1967,N_1781);
nor U2495 (N_2495,N_1754,N_1527);
or U2496 (N_2496,N_2055,N_1952);
nor U2497 (N_2497,N_2113,N_1520);
nand U2498 (N_2498,N_1878,N_1755);
nor U2499 (N_2499,N_2237,N_2133);
nor U2500 (N_2500,N_1629,N_1899);
nor U2501 (N_2501,N_1645,N_1599);
and U2502 (N_2502,N_2029,N_2087);
and U2503 (N_2503,N_1913,N_2213);
or U2504 (N_2504,N_1961,N_1619);
nand U2505 (N_2505,N_1743,N_1767);
or U2506 (N_2506,N_2018,N_2120);
nor U2507 (N_2507,N_1691,N_1718);
nor U2508 (N_2508,N_2223,N_1973);
nor U2509 (N_2509,N_1670,N_2095);
and U2510 (N_2510,N_1607,N_1940);
nor U2511 (N_2511,N_1660,N_1519);
nor U2512 (N_2512,N_1802,N_1551);
or U2513 (N_2513,N_2058,N_1974);
or U2514 (N_2514,N_1896,N_2003);
nand U2515 (N_2515,N_1644,N_2211);
and U2516 (N_2516,N_1622,N_1661);
nor U2517 (N_2517,N_2210,N_1507);
and U2518 (N_2518,N_1717,N_2248);
xnor U2519 (N_2519,N_1888,N_1693);
and U2520 (N_2520,N_1841,N_1840);
nor U2521 (N_2521,N_2037,N_1601);
or U2522 (N_2522,N_1772,N_1766);
nand U2523 (N_2523,N_1549,N_2104);
nand U2524 (N_2524,N_1502,N_2204);
or U2525 (N_2525,N_1732,N_1982);
nand U2526 (N_2526,N_1586,N_1641);
or U2527 (N_2527,N_2135,N_1570);
and U2528 (N_2528,N_1844,N_1765);
or U2529 (N_2529,N_1662,N_2205);
and U2530 (N_2530,N_2064,N_1632);
or U2531 (N_2531,N_1803,N_2045);
and U2532 (N_2532,N_1625,N_1894);
nor U2533 (N_2533,N_1927,N_1900);
and U2534 (N_2534,N_2152,N_2112);
nor U2535 (N_2535,N_1843,N_1671);
nor U2536 (N_2536,N_2042,N_1543);
and U2537 (N_2537,N_1658,N_2125);
or U2538 (N_2538,N_1763,N_2107);
or U2539 (N_2539,N_1850,N_2074);
nor U2540 (N_2540,N_1516,N_1566);
nor U2541 (N_2541,N_1504,N_1548);
nor U2542 (N_2542,N_2116,N_1713);
xnor U2543 (N_2543,N_1837,N_2077);
xnor U2544 (N_2544,N_1991,N_1946);
and U2545 (N_2545,N_2022,N_1777);
nand U2546 (N_2546,N_1945,N_2007);
or U2547 (N_2547,N_1897,N_1690);
and U2548 (N_2548,N_1943,N_1512);
nor U2549 (N_2549,N_1829,N_1756);
nor U2550 (N_2550,N_2171,N_2033);
nor U2551 (N_2551,N_1798,N_1565);
or U2552 (N_2552,N_1882,N_1742);
and U2553 (N_2553,N_2238,N_1851);
nand U2554 (N_2554,N_1789,N_1541);
and U2555 (N_2555,N_1573,N_1653);
nand U2556 (N_2556,N_1738,N_1852);
nor U2557 (N_2557,N_1539,N_1626);
or U2558 (N_2558,N_2036,N_1576);
or U2559 (N_2559,N_1720,N_1778);
nand U2560 (N_2560,N_2160,N_1780);
and U2561 (N_2561,N_1928,N_2068);
nor U2562 (N_2562,N_1596,N_2083);
and U2563 (N_2563,N_1631,N_1649);
or U2564 (N_2564,N_1680,N_1715);
or U2565 (N_2565,N_1775,N_1871);
and U2566 (N_2566,N_2128,N_1797);
or U2567 (N_2567,N_1733,N_1853);
and U2568 (N_2568,N_1679,N_2066);
and U2569 (N_2569,N_1706,N_1889);
nand U2570 (N_2570,N_1630,N_1590);
nor U2571 (N_2571,N_1534,N_1620);
or U2572 (N_2572,N_1752,N_1659);
nand U2573 (N_2573,N_2241,N_1722);
or U2574 (N_2574,N_1750,N_1562);
or U2575 (N_2575,N_2217,N_1589);
nand U2576 (N_2576,N_2097,N_1582);
and U2577 (N_2577,N_1958,N_1969);
and U2578 (N_2578,N_1705,N_1904);
or U2579 (N_2579,N_1618,N_1885);
or U2580 (N_2580,N_2199,N_1782);
nor U2581 (N_2581,N_2149,N_2239);
xor U2582 (N_2582,N_1912,N_2227);
nand U2583 (N_2583,N_1944,N_1557);
xor U2584 (N_2584,N_2224,N_2070);
or U2585 (N_2585,N_1687,N_1883);
nor U2586 (N_2586,N_1951,N_1839);
nand U2587 (N_2587,N_1563,N_2011);
nand U2588 (N_2588,N_1856,N_1592);
and U2589 (N_2589,N_2001,N_2063);
and U2590 (N_2590,N_1762,N_1567);
nor U2591 (N_2591,N_1860,N_1906);
nor U2592 (N_2592,N_1513,N_1683);
nor U2593 (N_2593,N_1575,N_1979);
nand U2594 (N_2594,N_2079,N_1528);
or U2595 (N_2595,N_1930,N_1929);
and U2596 (N_2596,N_2203,N_2048);
nand U2597 (N_2597,N_1999,N_2012);
xnor U2598 (N_2598,N_1615,N_1957);
or U2599 (N_2599,N_1847,N_1749);
or U2600 (N_2600,N_2085,N_2062);
nor U2601 (N_2601,N_1736,N_1656);
or U2602 (N_2602,N_2051,N_1600);
nand U2603 (N_2603,N_1584,N_2072);
nand U2604 (N_2604,N_2056,N_2117);
or U2605 (N_2605,N_2184,N_2101);
nor U2606 (N_2606,N_1740,N_2047);
nor U2607 (N_2607,N_2096,N_1784);
and U2608 (N_2608,N_1598,N_1830);
or U2609 (N_2609,N_1555,N_2189);
and U2610 (N_2610,N_2137,N_2017);
nand U2611 (N_2611,N_1794,N_1697);
or U2612 (N_2612,N_1634,N_1941);
and U2613 (N_2613,N_1975,N_2175);
or U2614 (N_2614,N_1515,N_1712);
nand U2615 (N_2615,N_2054,N_1804);
nand U2616 (N_2616,N_1606,N_2186);
nand U2617 (N_2617,N_1965,N_2134);
or U2618 (N_2618,N_2176,N_2040);
and U2619 (N_2619,N_1884,N_2091);
xnor U2620 (N_2620,N_1657,N_1731);
nor U2621 (N_2621,N_1877,N_2161);
and U2622 (N_2622,N_2235,N_2180);
nand U2623 (N_2623,N_1651,N_1835);
nand U2624 (N_2624,N_2172,N_1673);
nor U2625 (N_2625,N_1732,N_1832);
nand U2626 (N_2626,N_1943,N_1946);
and U2627 (N_2627,N_1780,N_1536);
xnor U2628 (N_2628,N_1935,N_1804);
nor U2629 (N_2629,N_1813,N_2146);
xor U2630 (N_2630,N_1621,N_1570);
nand U2631 (N_2631,N_1847,N_1523);
and U2632 (N_2632,N_1675,N_2030);
nand U2633 (N_2633,N_1725,N_2132);
nand U2634 (N_2634,N_2157,N_1504);
nor U2635 (N_2635,N_2224,N_1827);
and U2636 (N_2636,N_1638,N_1921);
or U2637 (N_2637,N_2043,N_2110);
nor U2638 (N_2638,N_2207,N_2118);
and U2639 (N_2639,N_1978,N_2176);
nand U2640 (N_2640,N_2183,N_2028);
nand U2641 (N_2641,N_2144,N_2140);
or U2642 (N_2642,N_1920,N_1630);
and U2643 (N_2643,N_2014,N_2113);
and U2644 (N_2644,N_1801,N_1650);
xor U2645 (N_2645,N_1764,N_2170);
nor U2646 (N_2646,N_2001,N_1841);
nand U2647 (N_2647,N_2040,N_2123);
nor U2648 (N_2648,N_2110,N_2220);
nor U2649 (N_2649,N_1760,N_2020);
nor U2650 (N_2650,N_1698,N_1611);
and U2651 (N_2651,N_1788,N_1533);
nor U2652 (N_2652,N_1504,N_1560);
and U2653 (N_2653,N_1558,N_1758);
and U2654 (N_2654,N_1584,N_1992);
nor U2655 (N_2655,N_1853,N_1644);
nor U2656 (N_2656,N_1814,N_2116);
or U2657 (N_2657,N_1534,N_1798);
or U2658 (N_2658,N_1769,N_2180);
nand U2659 (N_2659,N_1943,N_1562);
nand U2660 (N_2660,N_1666,N_1564);
nand U2661 (N_2661,N_2098,N_1777);
and U2662 (N_2662,N_1509,N_1546);
or U2663 (N_2663,N_1615,N_1833);
and U2664 (N_2664,N_2014,N_1934);
nor U2665 (N_2665,N_1639,N_1983);
nand U2666 (N_2666,N_1916,N_1566);
and U2667 (N_2667,N_2105,N_1996);
nand U2668 (N_2668,N_1762,N_1845);
or U2669 (N_2669,N_1557,N_2128);
and U2670 (N_2670,N_2038,N_1963);
and U2671 (N_2671,N_1750,N_1626);
nor U2672 (N_2672,N_1846,N_2092);
nor U2673 (N_2673,N_1831,N_1763);
and U2674 (N_2674,N_2101,N_1674);
and U2675 (N_2675,N_2213,N_2140);
and U2676 (N_2676,N_1657,N_2136);
nand U2677 (N_2677,N_1748,N_1842);
nor U2678 (N_2678,N_2214,N_1658);
nand U2679 (N_2679,N_1973,N_2157);
nand U2680 (N_2680,N_1790,N_1858);
or U2681 (N_2681,N_2148,N_1559);
or U2682 (N_2682,N_1787,N_2070);
nand U2683 (N_2683,N_1804,N_1545);
nor U2684 (N_2684,N_1887,N_1961);
xnor U2685 (N_2685,N_2070,N_1586);
or U2686 (N_2686,N_1651,N_1913);
or U2687 (N_2687,N_2198,N_1971);
and U2688 (N_2688,N_1856,N_1681);
and U2689 (N_2689,N_2085,N_2232);
nor U2690 (N_2690,N_1804,N_1762);
and U2691 (N_2691,N_2162,N_2138);
nor U2692 (N_2692,N_1977,N_1759);
or U2693 (N_2693,N_2048,N_2108);
or U2694 (N_2694,N_1650,N_1633);
and U2695 (N_2695,N_1635,N_2036);
nor U2696 (N_2696,N_1638,N_1585);
and U2697 (N_2697,N_1510,N_1945);
nor U2698 (N_2698,N_1795,N_1554);
and U2699 (N_2699,N_1711,N_1956);
and U2700 (N_2700,N_2023,N_2000);
nor U2701 (N_2701,N_2128,N_1832);
nor U2702 (N_2702,N_2238,N_1697);
and U2703 (N_2703,N_2003,N_2166);
xor U2704 (N_2704,N_1638,N_1818);
nand U2705 (N_2705,N_1835,N_2018);
or U2706 (N_2706,N_1683,N_1728);
and U2707 (N_2707,N_1739,N_1648);
nor U2708 (N_2708,N_1653,N_2204);
and U2709 (N_2709,N_1816,N_1763);
and U2710 (N_2710,N_2094,N_1684);
and U2711 (N_2711,N_2134,N_1902);
nor U2712 (N_2712,N_1825,N_2044);
or U2713 (N_2713,N_2035,N_1808);
or U2714 (N_2714,N_1713,N_2199);
or U2715 (N_2715,N_2244,N_1858);
nand U2716 (N_2716,N_2073,N_2003);
nor U2717 (N_2717,N_1813,N_2027);
nor U2718 (N_2718,N_1548,N_1635);
and U2719 (N_2719,N_2051,N_1525);
nor U2720 (N_2720,N_2169,N_1551);
nor U2721 (N_2721,N_1782,N_1548);
nand U2722 (N_2722,N_1521,N_1924);
and U2723 (N_2723,N_2067,N_1881);
or U2724 (N_2724,N_1987,N_1598);
nor U2725 (N_2725,N_1653,N_2049);
or U2726 (N_2726,N_2182,N_1905);
or U2727 (N_2727,N_1772,N_1871);
nor U2728 (N_2728,N_1700,N_2189);
nand U2729 (N_2729,N_2060,N_1830);
or U2730 (N_2730,N_1870,N_2092);
and U2731 (N_2731,N_2104,N_1743);
and U2732 (N_2732,N_2107,N_1822);
or U2733 (N_2733,N_1720,N_1709);
or U2734 (N_2734,N_2144,N_1880);
nand U2735 (N_2735,N_1724,N_1833);
or U2736 (N_2736,N_1955,N_1527);
nor U2737 (N_2737,N_1507,N_1991);
or U2738 (N_2738,N_2074,N_1796);
nand U2739 (N_2739,N_2105,N_1612);
nand U2740 (N_2740,N_1830,N_1589);
and U2741 (N_2741,N_1662,N_2233);
and U2742 (N_2742,N_1800,N_2134);
nand U2743 (N_2743,N_1831,N_1811);
nor U2744 (N_2744,N_1643,N_2204);
or U2745 (N_2745,N_1781,N_1682);
nand U2746 (N_2746,N_1895,N_1995);
nor U2747 (N_2747,N_1574,N_2159);
nor U2748 (N_2748,N_1568,N_2238);
nand U2749 (N_2749,N_1788,N_1632);
nand U2750 (N_2750,N_2149,N_1778);
nor U2751 (N_2751,N_1950,N_2043);
and U2752 (N_2752,N_2155,N_2027);
nand U2753 (N_2753,N_1868,N_1867);
nand U2754 (N_2754,N_1793,N_1552);
or U2755 (N_2755,N_2108,N_2020);
or U2756 (N_2756,N_2199,N_1840);
nand U2757 (N_2757,N_2101,N_1834);
nand U2758 (N_2758,N_2018,N_1819);
and U2759 (N_2759,N_2249,N_1610);
nand U2760 (N_2760,N_1968,N_1733);
nor U2761 (N_2761,N_2238,N_1558);
or U2762 (N_2762,N_1509,N_1853);
nand U2763 (N_2763,N_1610,N_2034);
and U2764 (N_2764,N_1652,N_2225);
or U2765 (N_2765,N_1928,N_1987);
nor U2766 (N_2766,N_2053,N_1622);
or U2767 (N_2767,N_1610,N_2074);
nor U2768 (N_2768,N_1543,N_1697);
and U2769 (N_2769,N_1504,N_1689);
xor U2770 (N_2770,N_2216,N_2148);
and U2771 (N_2771,N_1751,N_1618);
nor U2772 (N_2772,N_1965,N_1812);
and U2773 (N_2773,N_1572,N_2197);
or U2774 (N_2774,N_1612,N_1856);
nor U2775 (N_2775,N_1741,N_1769);
or U2776 (N_2776,N_2024,N_2146);
nor U2777 (N_2777,N_2075,N_2026);
or U2778 (N_2778,N_1740,N_2010);
nor U2779 (N_2779,N_1896,N_2214);
and U2780 (N_2780,N_1718,N_1906);
and U2781 (N_2781,N_2152,N_1983);
or U2782 (N_2782,N_1627,N_1814);
nand U2783 (N_2783,N_1939,N_2083);
nand U2784 (N_2784,N_1795,N_1661);
and U2785 (N_2785,N_1874,N_1671);
and U2786 (N_2786,N_1542,N_1549);
or U2787 (N_2787,N_1703,N_2004);
nand U2788 (N_2788,N_1843,N_2000);
or U2789 (N_2789,N_2134,N_1523);
and U2790 (N_2790,N_2087,N_1676);
nor U2791 (N_2791,N_1583,N_1954);
nor U2792 (N_2792,N_1680,N_1805);
xor U2793 (N_2793,N_2108,N_1793);
or U2794 (N_2794,N_1636,N_1739);
or U2795 (N_2795,N_1839,N_1908);
nor U2796 (N_2796,N_2106,N_1789);
xor U2797 (N_2797,N_1977,N_1524);
nand U2798 (N_2798,N_2135,N_2156);
nand U2799 (N_2799,N_1806,N_2245);
nor U2800 (N_2800,N_1649,N_1699);
nand U2801 (N_2801,N_1830,N_2117);
or U2802 (N_2802,N_1773,N_1889);
nor U2803 (N_2803,N_1699,N_2028);
or U2804 (N_2804,N_1657,N_2217);
nor U2805 (N_2805,N_1719,N_2055);
and U2806 (N_2806,N_1819,N_2163);
or U2807 (N_2807,N_1993,N_1883);
or U2808 (N_2808,N_1979,N_2168);
nand U2809 (N_2809,N_1954,N_1787);
nor U2810 (N_2810,N_2052,N_2248);
and U2811 (N_2811,N_2055,N_1763);
nand U2812 (N_2812,N_2214,N_2156);
nand U2813 (N_2813,N_1867,N_2240);
nor U2814 (N_2814,N_2077,N_2143);
and U2815 (N_2815,N_1513,N_2121);
nor U2816 (N_2816,N_1772,N_2100);
nor U2817 (N_2817,N_1951,N_2146);
nand U2818 (N_2818,N_1587,N_1683);
and U2819 (N_2819,N_2031,N_1927);
or U2820 (N_2820,N_2169,N_1693);
nand U2821 (N_2821,N_2202,N_1973);
or U2822 (N_2822,N_1528,N_1787);
and U2823 (N_2823,N_1911,N_2163);
nor U2824 (N_2824,N_2208,N_1664);
and U2825 (N_2825,N_1627,N_1941);
or U2826 (N_2826,N_1682,N_1729);
nor U2827 (N_2827,N_1804,N_1590);
and U2828 (N_2828,N_1925,N_1549);
nand U2829 (N_2829,N_1799,N_1612);
or U2830 (N_2830,N_2214,N_1558);
nand U2831 (N_2831,N_1557,N_1868);
nor U2832 (N_2832,N_1704,N_1911);
nor U2833 (N_2833,N_1607,N_1724);
nor U2834 (N_2834,N_1940,N_2110);
or U2835 (N_2835,N_1952,N_1872);
and U2836 (N_2836,N_1703,N_2081);
xor U2837 (N_2837,N_1778,N_1681);
nand U2838 (N_2838,N_2000,N_2014);
or U2839 (N_2839,N_1699,N_1877);
nor U2840 (N_2840,N_2041,N_2055);
nor U2841 (N_2841,N_1618,N_1750);
and U2842 (N_2842,N_2134,N_1908);
nor U2843 (N_2843,N_2114,N_2244);
nand U2844 (N_2844,N_2227,N_1602);
and U2845 (N_2845,N_1862,N_1955);
nor U2846 (N_2846,N_1756,N_1512);
nor U2847 (N_2847,N_2180,N_1908);
nand U2848 (N_2848,N_2181,N_1831);
nand U2849 (N_2849,N_1901,N_1701);
or U2850 (N_2850,N_1987,N_2181);
nor U2851 (N_2851,N_1924,N_1801);
or U2852 (N_2852,N_1903,N_1685);
nand U2853 (N_2853,N_1659,N_2145);
or U2854 (N_2854,N_1956,N_1875);
nor U2855 (N_2855,N_1607,N_1912);
nand U2856 (N_2856,N_2119,N_1517);
or U2857 (N_2857,N_2063,N_1736);
or U2858 (N_2858,N_2158,N_1802);
and U2859 (N_2859,N_2140,N_1706);
or U2860 (N_2860,N_1866,N_1881);
nand U2861 (N_2861,N_1706,N_1651);
nand U2862 (N_2862,N_2172,N_1911);
or U2863 (N_2863,N_2056,N_2085);
or U2864 (N_2864,N_1998,N_2121);
or U2865 (N_2865,N_2239,N_2070);
or U2866 (N_2866,N_1728,N_2148);
nand U2867 (N_2867,N_2120,N_2157);
nand U2868 (N_2868,N_2164,N_1512);
and U2869 (N_2869,N_2178,N_1535);
nor U2870 (N_2870,N_2060,N_1685);
and U2871 (N_2871,N_2134,N_2193);
nor U2872 (N_2872,N_1727,N_1718);
nand U2873 (N_2873,N_2067,N_2125);
nand U2874 (N_2874,N_2098,N_1712);
xnor U2875 (N_2875,N_2167,N_2177);
and U2876 (N_2876,N_2016,N_1896);
nand U2877 (N_2877,N_1911,N_1536);
xor U2878 (N_2878,N_1765,N_1884);
and U2879 (N_2879,N_1835,N_1927);
and U2880 (N_2880,N_2127,N_1792);
and U2881 (N_2881,N_1817,N_1863);
or U2882 (N_2882,N_1885,N_2100);
nand U2883 (N_2883,N_2039,N_2007);
nor U2884 (N_2884,N_1638,N_2200);
nor U2885 (N_2885,N_2210,N_1532);
nand U2886 (N_2886,N_2131,N_2063);
and U2887 (N_2887,N_1500,N_2011);
nor U2888 (N_2888,N_1995,N_2089);
nand U2889 (N_2889,N_2040,N_2154);
or U2890 (N_2890,N_1937,N_2242);
or U2891 (N_2891,N_1522,N_2236);
xnor U2892 (N_2892,N_1532,N_2044);
nor U2893 (N_2893,N_1813,N_1968);
and U2894 (N_2894,N_1949,N_1704);
or U2895 (N_2895,N_2059,N_1952);
nand U2896 (N_2896,N_1721,N_1855);
and U2897 (N_2897,N_1593,N_1735);
nand U2898 (N_2898,N_1918,N_2193);
and U2899 (N_2899,N_1648,N_2163);
nand U2900 (N_2900,N_1738,N_1819);
nand U2901 (N_2901,N_2097,N_1563);
nand U2902 (N_2902,N_2071,N_1705);
nand U2903 (N_2903,N_1614,N_1662);
or U2904 (N_2904,N_2078,N_1788);
and U2905 (N_2905,N_1848,N_1647);
nand U2906 (N_2906,N_2228,N_1527);
nor U2907 (N_2907,N_1708,N_1834);
xor U2908 (N_2908,N_1653,N_1751);
nor U2909 (N_2909,N_2023,N_1764);
and U2910 (N_2910,N_2191,N_2198);
nor U2911 (N_2911,N_1557,N_1608);
or U2912 (N_2912,N_1850,N_1674);
nor U2913 (N_2913,N_1950,N_2151);
nand U2914 (N_2914,N_2182,N_1856);
and U2915 (N_2915,N_2039,N_1984);
and U2916 (N_2916,N_2133,N_1653);
nand U2917 (N_2917,N_1782,N_1576);
or U2918 (N_2918,N_1895,N_1666);
or U2919 (N_2919,N_1552,N_1935);
nor U2920 (N_2920,N_1631,N_2014);
and U2921 (N_2921,N_1719,N_2077);
nor U2922 (N_2922,N_2160,N_2227);
nand U2923 (N_2923,N_1776,N_2059);
and U2924 (N_2924,N_1609,N_1547);
or U2925 (N_2925,N_1775,N_1618);
and U2926 (N_2926,N_1883,N_1679);
nor U2927 (N_2927,N_1981,N_1643);
nor U2928 (N_2928,N_2186,N_2236);
nor U2929 (N_2929,N_1806,N_2177);
nand U2930 (N_2930,N_1695,N_1854);
nand U2931 (N_2931,N_2108,N_1716);
nand U2932 (N_2932,N_1928,N_1925);
or U2933 (N_2933,N_2099,N_1977);
or U2934 (N_2934,N_1767,N_1936);
and U2935 (N_2935,N_1544,N_2215);
nand U2936 (N_2936,N_1513,N_1890);
nor U2937 (N_2937,N_1550,N_1976);
nor U2938 (N_2938,N_1910,N_2070);
nor U2939 (N_2939,N_2194,N_2044);
or U2940 (N_2940,N_2221,N_2007);
or U2941 (N_2941,N_2077,N_2004);
nor U2942 (N_2942,N_1631,N_1768);
xor U2943 (N_2943,N_1775,N_1580);
nor U2944 (N_2944,N_1897,N_2166);
or U2945 (N_2945,N_1525,N_2056);
nor U2946 (N_2946,N_1935,N_2184);
nand U2947 (N_2947,N_1526,N_1639);
and U2948 (N_2948,N_1930,N_1683);
nor U2949 (N_2949,N_2209,N_1908);
nand U2950 (N_2950,N_2186,N_2240);
or U2951 (N_2951,N_2120,N_1835);
nand U2952 (N_2952,N_1525,N_2010);
or U2953 (N_2953,N_1531,N_1931);
or U2954 (N_2954,N_1697,N_2031);
nand U2955 (N_2955,N_1520,N_1536);
nand U2956 (N_2956,N_1548,N_1684);
nand U2957 (N_2957,N_2044,N_1709);
and U2958 (N_2958,N_1706,N_2207);
nand U2959 (N_2959,N_2107,N_2005);
nor U2960 (N_2960,N_2002,N_2240);
nor U2961 (N_2961,N_1773,N_2141);
nand U2962 (N_2962,N_1710,N_1876);
nand U2963 (N_2963,N_1981,N_1987);
nor U2964 (N_2964,N_2132,N_1922);
nand U2965 (N_2965,N_1638,N_2085);
nor U2966 (N_2966,N_2003,N_2115);
nand U2967 (N_2967,N_1925,N_1645);
or U2968 (N_2968,N_2042,N_1810);
or U2969 (N_2969,N_1828,N_2085);
and U2970 (N_2970,N_1580,N_2230);
nand U2971 (N_2971,N_1736,N_2238);
xor U2972 (N_2972,N_2029,N_1832);
nand U2973 (N_2973,N_1921,N_1967);
nor U2974 (N_2974,N_1938,N_1910);
nor U2975 (N_2975,N_1925,N_1598);
nor U2976 (N_2976,N_1715,N_1831);
or U2977 (N_2977,N_1584,N_2192);
nand U2978 (N_2978,N_2229,N_1739);
nand U2979 (N_2979,N_1876,N_1853);
or U2980 (N_2980,N_2136,N_1638);
xor U2981 (N_2981,N_2040,N_1808);
or U2982 (N_2982,N_1612,N_2026);
or U2983 (N_2983,N_1586,N_1553);
nand U2984 (N_2984,N_2161,N_2067);
nor U2985 (N_2985,N_1697,N_2114);
nand U2986 (N_2986,N_2193,N_1917);
or U2987 (N_2987,N_2158,N_2246);
nand U2988 (N_2988,N_1726,N_1745);
and U2989 (N_2989,N_2198,N_1726);
nor U2990 (N_2990,N_2056,N_1707);
and U2991 (N_2991,N_1643,N_1710);
nand U2992 (N_2992,N_1971,N_1661);
and U2993 (N_2993,N_1581,N_2103);
nand U2994 (N_2994,N_2150,N_1554);
or U2995 (N_2995,N_2110,N_1728);
and U2996 (N_2996,N_1708,N_2066);
nor U2997 (N_2997,N_1968,N_1981);
nor U2998 (N_2998,N_1778,N_1500);
or U2999 (N_2999,N_1687,N_1562);
or UO_0 (O_0,N_2625,N_2500);
and UO_1 (O_1,N_2819,N_2435);
or UO_2 (O_2,N_2696,N_2554);
nor UO_3 (O_3,N_2714,N_2637);
or UO_4 (O_4,N_2590,N_2845);
nand UO_5 (O_5,N_2348,N_2759);
or UO_6 (O_6,N_2362,N_2779);
nand UO_7 (O_7,N_2560,N_2765);
nor UO_8 (O_8,N_2720,N_2970);
nand UO_9 (O_9,N_2326,N_2942);
nand UO_10 (O_10,N_2367,N_2470);
or UO_11 (O_11,N_2302,N_2515);
nor UO_12 (O_12,N_2643,N_2337);
or UO_13 (O_13,N_2342,N_2947);
and UO_14 (O_14,N_2962,N_2792);
and UO_15 (O_15,N_2494,N_2938);
and UO_16 (O_16,N_2433,N_2727);
nor UO_17 (O_17,N_2722,N_2730);
nor UO_18 (O_18,N_2859,N_2331);
or UO_19 (O_19,N_2529,N_2275);
nor UO_20 (O_20,N_2370,N_2377);
nand UO_21 (O_21,N_2886,N_2707);
and UO_22 (O_22,N_2907,N_2613);
or UO_23 (O_23,N_2684,N_2545);
nor UO_24 (O_24,N_2624,N_2540);
and UO_25 (O_25,N_2508,N_2833);
and UO_26 (O_26,N_2704,N_2873);
nor UO_27 (O_27,N_2524,N_2852);
and UO_28 (O_28,N_2851,N_2703);
and UO_29 (O_29,N_2677,N_2998);
nor UO_30 (O_30,N_2339,N_2283);
or UO_31 (O_31,N_2816,N_2577);
and UO_32 (O_32,N_2518,N_2454);
or UO_33 (O_33,N_2335,N_2534);
nand UO_34 (O_34,N_2569,N_2300);
or UO_35 (O_35,N_2650,N_2341);
and UO_36 (O_36,N_2604,N_2378);
and UO_37 (O_37,N_2738,N_2394);
nor UO_38 (O_38,N_2736,N_2847);
and UO_39 (O_39,N_2700,N_2880);
and UO_40 (O_40,N_2572,N_2951);
or UO_41 (O_41,N_2799,N_2594);
or UO_42 (O_42,N_2523,N_2877);
or UO_43 (O_43,N_2745,N_2869);
or UO_44 (O_44,N_2413,N_2807);
or UO_45 (O_45,N_2981,N_2739);
xnor UO_46 (O_46,N_2679,N_2855);
and UO_47 (O_47,N_2443,N_2620);
nor UO_48 (O_48,N_2895,N_2626);
nor UO_49 (O_49,N_2393,N_2689);
xnor UO_50 (O_50,N_2610,N_2285);
and UO_51 (O_51,N_2512,N_2871);
nand UO_52 (O_52,N_2860,N_2708);
and UO_53 (O_53,N_2408,N_2657);
nand UO_54 (O_54,N_2823,N_2449);
and UO_55 (O_55,N_2716,N_2828);
and UO_56 (O_56,N_2486,N_2314);
and UO_57 (O_57,N_2972,N_2313);
and UO_58 (O_58,N_2264,N_2281);
nor UO_59 (O_59,N_2891,N_2587);
or UO_60 (O_60,N_2591,N_2784);
and UO_61 (O_61,N_2836,N_2967);
nor UO_62 (O_62,N_2830,N_2905);
nand UO_63 (O_63,N_2582,N_2531);
nor UO_64 (O_64,N_2278,N_2556);
and UO_65 (O_65,N_2287,N_2597);
nor UO_66 (O_66,N_2966,N_2850);
or UO_67 (O_67,N_2919,N_2344);
nor UO_68 (O_68,N_2969,N_2363);
or UO_69 (O_69,N_2780,N_2824);
nor UO_70 (O_70,N_2632,N_2786);
nand UO_71 (O_71,N_2724,N_2544);
and UO_72 (O_72,N_2863,N_2405);
nor UO_73 (O_73,N_2701,N_2996);
nand UO_74 (O_74,N_2472,N_2647);
or UO_75 (O_75,N_2420,N_2955);
nor UO_76 (O_76,N_2915,N_2719);
xnor UO_77 (O_77,N_2878,N_2762);
nand UO_78 (O_78,N_2528,N_2537);
nor UO_79 (O_79,N_2984,N_2491);
or UO_80 (O_80,N_2766,N_2920);
and UO_81 (O_81,N_2261,N_2894);
or UO_82 (O_82,N_2801,N_2434);
nor UO_83 (O_83,N_2777,N_2897);
nand UO_84 (O_84,N_2520,N_2543);
nor UO_85 (O_85,N_2617,N_2715);
nand UO_86 (O_86,N_2676,N_2728);
nor UO_87 (O_87,N_2593,N_2634);
nor UO_88 (O_88,N_2994,N_2619);
and UO_89 (O_89,N_2916,N_2585);
and UO_90 (O_90,N_2459,N_2698);
nor UO_91 (O_91,N_2929,N_2387);
and UO_92 (O_92,N_2546,N_2579);
nor UO_93 (O_93,N_2499,N_2890);
nand UO_94 (O_94,N_2723,N_2813);
and UO_95 (O_95,N_2492,N_2566);
nand UO_96 (O_96,N_2254,N_2710);
or UO_97 (O_97,N_2429,N_2950);
and UO_98 (O_98,N_2640,N_2752);
and UO_99 (O_99,N_2446,N_2810);
or UO_100 (O_100,N_2674,N_2849);
and UO_101 (O_101,N_2959,N_2267);
nor UO_102 (O_102,N_2360,N_2699);
and UO_103 (O_103,N_2359,N_2806);
nor UO_104 (O_104,N_2965,N_2361);
nor UO_105 (O_105,N_2770,N_2404);
and UO_106 (O_106,N_2767,N_2258);
nand UO_107 (O_107,N_2925,N_2776);
and UO_108 (O_108,N_2973,N_2385);
nand UO_109 (O_109,N_2686,N_2474);
or UO_110 (O_110,N_2666,N_2868);
nor UO_111 (O_111,N_2255,N_2865);
nor UO_112 (O_112,N_2516,N_2311);
nor UO_113 (O_113,N_2910,N_2272);
or UO_114 (O_114,N_2366,N_2761);
nand UO_115 (O_115,N_2441,N_2580);
nand UO_116 (O_116,N_2256,N_2940);
nor UO_117 (O_117,N_2747,N_2768);
nor UO_118 (O_118,N_2373,N_2602);
nand UO_119 (O_119,N_2867,N_2416);
nand UO_120 (O_120,N_2286,N_2414);
nand UO_121 (O_121,N_2812,N_2542);
or UO_122 (O_122,N_2844,N_2756);
nor UO_123 (O_123,N_2334,N_2609);
nor UO_124 (O_124,N_2665,N_2980);
and UO_125 (O_125,N_2596,N_2928);
nand UO_126 (O_126,N_2675,N_2588);
and UO_127 (O_127,N_2375,N_2987);
nand UO_128 (O_128,N_2706,N_2406);
nand UO_129 (O_129,N_2646,N_2513);
nand UO_130 (O_130,N_2791,N_2451);
and UO_131 (O_131,N_2858,N_2755);
nand UO_132 (O_132,N_2304,N_2336);
nand UO_133 (O_133,N_2380,N_2427);
nand UO_134 (O_134,N_2993,N_2964);
or UO_135 (O_135,N_2971,N_2896);
and UO_136 (O_136,N_2376,N_2496);
and UO_137 (O_137,N_2997,N_2908);
nand UO_138 (O_138,N_2575,N_2732);
nor UO_139 (O_139,N_2837,N_2517);
or UO_140 (O_140,N_2390,N_2631);
nor UO_141 (O_141,N_2913,N_2794);
and UO_142 (O_142,N_2299,N_2789);
nand UO_143 (O_143,N_2857,N_2511);
nor UO_144 (O_144,N_2750,N_2760);
nand UO_145 (O_145,N_2324,N_2932);
and UO_146 (O_146,N_2442,N_2638);
nor UO_147 (O_147,N_2317,N_2651);
and UO_148 (O_148,N_2384,N_2683);
and UO_149 (O_149,N_2567,N_2338);
or UO_150 (O_150,N_2977,N_2532);
and UO_151 (O_151,N_2729,N_2282);
and UO_152 (O_152,N_2957,N_2288);
nand UO_153 (O_153,N_2424,N_2327);
or UO_154 (O_154,N_2692,N_2548);
and UO_155 (O_155,N_2693,N_2653);
and UO_156 (O_156,N_2725,N_2635);
nor UO_157 (O_157,N_2927,N_2737);
xnor UO_158 (O_158,N_2428,N_2788);
and UO_159 (O_159,N_2892,N_2525);
nand UO_160 (O_160,N_2937,N_2388);
or UO_161 (O_161,N_2347,N_2303);
nand UO_162 (O_162,N_2992,N_2346);
and UO_163 (O_163,N_2445,N_2506);
nor UO_164 (O_164,N_2711,N_2948);
nor UO_165 (O_165,N_2986,N_2589);
nand UO_166 (O_166,N_2349,N_2648);
nand UO_167 (O_167,N_2423,N_2764);
or UO_168 (O_168,N_2259,N_2407);
nand UO_169 (O_169,N_2561,N_2954);
and UO_170 (O_170,N_2583,N_2636);
nand UO_171 (O_171,N_2563,N_2906);
or UO_172 (O_172,N_2505,N_2923);
or UO_173 (O_173,N_2843,N_2773);
nand UO_174 (O_174,N_2562,N_2568);
or UO_175 (O_175,N_2968,N_2945);
and UO_176 (O_176,N_2936,N_2804);
nand UO_177 (O_177,N_2697,N_2252);
nor UO_178 (O_178,N_2774,N_2310);
or UO_179 (O_179,N_2931,N_2976);
and UO_180 (O_180,N_2325,N_2982);
nand UO_181 (O_181,N_2271,N_2622);
and UO_182 (O_182,N_2251,N_2817);
nand UO_183 (O_183,N_2269,N_2262);
nor UO_184 (O_184,N_2538,N_2308);
and UO_185 (O_185,N_2495,N_2498);
and UO_186 (O_186,N_2422,N_2615);
or UO_187 (O_187,N_2547,N_2641);
nor UO_188 (O_188,N_2846,N_2616);
nor UO_189 (O_189,N_2787,N_2879);
nor UO_190 (O_190,N_2821,N_2452);
and UO_191 (O_191,N_2527,N_2260);
or UO_192 (O_192,N_2900,N_2401);
nor UO_193 (O_193,N_2289,N_2914);
or UO_194 (O_194,N_2305,N_2944);
or UO_195 (O_195,N_2270,N_2870);
nor UO_196 (O_196,N_2514,N_2803);
or UO_197 (O_197,N_2555,N_2426);
and UO_198 (O_198,N_2979,N_2618);
or UO_199 (O_199,N_2330,N_2295);
and UO_200 (O_200,N_2864,N_2576);
and UO_201 (O_201,N_2985,N_2328);
and UO_202 (O_202,N_2409,N_2660);
or UO_203 (O_203,N_2383,N_2521);
nand UO_204 (O_204,N_2503,N_2595);
or UO_205 (O_205,N_2705,N_2685);
or UO_206 (O_206,N_2309,N_2306);
xnor UO_207 (O_207,N_2988,N_2802);
or UO_208 (O_208,N_2782,N_2758);
or UO_209 (O_209,N_2291,N_2882);
nand UO_210 (O_210,N_2374,N_2565);
or UO_211 (O_211,N_2436,N_2466);
or UO_212 (O_212,N_2899,N_2898);
nor UO_213 (O_213,N_2365,N_2476);
nand UO_214 (O_214,N_2558,N_2600);
nand UO_215 (O_215,N_2983,N_2838);
and UO_216 (O_216,N_2775,N_2811);
nor UO_217 (O_217,N_2364,N_2746);
and UO_218 (O_218,N_2301,N_2468);
nor UO_219 (O_219,N_2717,N_2276);
and UO_220 (O_220,N_2721,N_2343);
nand UO_221 (O_221,N_2652,N_2961);
nor UO_222 (O_222,N_2471,N_2463);
xor UO_223 (O_223,N_2574,N_2273);
nand UO_224 (O_224,N_2956,N_2805);
and UO_225 (O_225,N_2412,N_2415);
or UO_226 (O_226,N_2818,N_2430);
nor UO_227 (O_227,N_2796,N_2584);
nand UO_228 (O_228,N_2354,N_2733);
nand UO_229 (O_229,N_2389,N_2866);
xnor UO_230 (O_230,N_2448,N_2438);
and UO_231 (O_231,N_2655,N_2355);
or UO_232 (O_232,N_2453,N_2933);
nand UO_233 (O_233,N_2290,N_2629);
or UO_234 (O_234,N_2578,N_2663);
or UO_235 (O_235,N_2601,N_2396);
nand UO_236 (O_236,N_2695,N_2501);
and UO_237 (O_237,N_2307,N_2741);
and UO_238 (O_238,N_2450,N_2599);
xnor UO_239 (O_239,N_2744,N_2671);
or UO_240 (O_240,N_2772,N_2482);
nand UO_241 (O_241,N_2379,N_2297);
or UO_242 (O_242,N_2659,N_2753);
nor UO_243 (O_243,N_2667,N_2460);
or UO_244 (O_244,N_2608,N_2368);
and UO_245 (O_245,N_2483,N_2795);
nor UO_246 (O_246,N_2887,N_2934);
or UO_247 (O_247,N_2645,N_2550);
nor UO_248 (O_248,N_2691,N_2861);
and UO_249 (O_249,N_2834,N_2825);
or UO_250 (O_250,N_2464,N_2778);
nand UO_251 (O_251,N_2842,N_2809);
nor UO_252 (O_252,N_2315,N_2400);
nor UO_253 (O_253,N_2694,N_2841);
nand UO_254 (O_254,N_2351,N_2681);
and UO_255 (O_255,N_2318,N_2353);
and UO_256 (O_256,N_2661,N_2358);
or UO_257 (O_257,N_2356,N_2902);
and UO_258 (O_258,N_2623,N_2382);
nor UO_259 (O_259,N_2439,N_2437);
nor UO_260 (O_260,N_2535,N_2519);
or UO_261 (O_261,N_2510,N_2526);
nor UO_262 (O_262,N_2263,N_2690);
or UO_263 (O_263,N_2876,N_2398);
nor UO_264 (O_264,N_2975,N_2848);
nand UO_265 (O_265,N_2649,N_2952);
or UO_266 (O_266,N_2885,N_2279);
nor UO_267 (O_267,N_2904,N_2820);
or UO_268 (O_268,N_2884,N_2668);
or UO_269 (O_269,N_2477,N_2888);
nand UO_270 (O_270,N_2440,N_2627);
nand UO_271 (O_271,N_2481,N_2901);
nand UO_272 (O_272,N_2431,N_2918);
nor UO_273 (O_273,N_2475,N_2991);
or UO_274 (O_274,N_2487,N_2410);
nor UO_275 (O_275,N_2533,N_2284);
nor UO_276 (O_276,N_2670,N_2332);
nand UO_277 (O_277,N_2573,N_2473);
nand UO_278 (O_278,N_2493,N_2781);
nor UO_279 (O_279,N_2911,N_2357);
nor UO_280 (O_280,N_2656,N_2658);
and UO_281 (O_281,N_2909,N_2614);
nor UO_282 (O_282,N_2989,N_2630);
xor UO_283 (O_283,N_2662,N_2903);
or UO_284 (O_284,N_2922,N_2391);
nand UO_285 (O_285,N_2447,N_2953);
and UO_286 (O_286,N_2266,N_2718);
or UO_287 (O_287,N_2571,N_2417);
nor UO_288 (O_288,N_2322,N_2990);
nand UO_289 (O_289,N_2381,N_2941);
or UO_290 (O_290,N_2606,N_2687);
nor UO_291 (O_291,N_2735,N_2827);
nor UO_292 (O_292,N_2541,N_2960);
nand UO_293 (O_293,N_2444,N_2826);
nor UO_294 (O_294,N_2639,N_2536);
and UO_295 (O_295,N_2369,N_2935);
nor UO_296 (O_296,N_2978,N_2734);
nand UO_297 (O_297,N_2280,N_2628);
nand UO_298 (O_298,N_2250,N_2564);
and UO_299 (O_299,N_2642,N_2712);
and UO_300 (O_300,N_2673,N_2748);
or UO_301 (O_301,N_2999,N_2749);
and UO_302 (O_302,N_2316,N_2467);
and UO_303 (O_303,N_2822,N_2598);
or UO_304 (O_304,N_2553,N_2702);
nand UO_305 (O_305,N_2485,N_2644);
and UO_306 (O_306,N_2603,N_2461);
nand UO_307 (O_307,N_2480,N_2455);
or UO_308 (O_308,N_2839,N_2757);
and UO_309 (O_309,N_2893,N_2680);
or UO_310 (O_310,N_2783,N_2484);
nand UO_311 (O_311,N_2862,N_2539);
nor UO_312 (O_312,N_2958,N_2743);
and UO_313 (O_313,N_2771,N_2465);
nand UO_314 (O_314,N_2489,N_2293);
and UO_315 (O_315,N_2831,N_2411);
or UO_316 (O_316,N_2333,N_2298);
or UO_317 (O_317,N_2522,N_2504);
nand UO_318 (O_318,N_2478,N_2418);
and UO_319 (O_319,N_2319,N_2457);
nand UO_320 (O_320,N_2800,N_2456);
and UO_321 (O_321,N_2881,N_2425);
nand UO_322 (O_322,N_2551,N_2296);
or UO_323 (O_323,N_2949,N_2497);
nand UO_324 (O_324,N_2726,N_2432);
nand UO_325 (O_325,N_2458,N_2633);
or UO_326 (O_326,N_2320,N_2312);
and UO_327 (O_327,N_2557,N_2419);
and UO_328 (O_328,N_2479,N_2672);
nor UO_329 (O_329,N_2856,N_2963);
or UO_330 (O_330,N_2930,N_2939);
nor UO_331 (O_331,N_2399,N_2924);
and UO_332 (O_332,N_2403,N_2840);
nand UO_333 (O_333,N_2507,N_2883);
or UO_334 (O_334,N_2277,N_2386);
nand UO_335 (O_335,N_2581,N_2502);
nand UO_336 (O_336,N_2421,N_2654);
nor UO_337 (O_337,N_2592,N_2292);
and UO_338 (O_338,N_2763,N_2607);
and UO_339 (O_339,N_2321,N_2552);
nor UO_340 (O_340,N_2549,N_2664);
or UO_341 (O_341,N_2874,N_2392);
nand UO_342 (O_342,N_2265,N_2912);
or UO_343 (O_343,N_2509,N_2946);
or UO_344 (O_344,N_2559,N_2350);
and UO_345 (O_345,N_2397,N_2889);
nand UO_346 (O_346,N_2570,N_2257);
or UO_347 (O_347,N_2742,N_2740);
nor UO_348 (O_348,N_2943,N_2323);
xnor UO_349 (O_349,N_2329,N_2974);
nand UO_350 (O_350,N_2854,N_2490);
nor UO_351 (O_351,N_2790,N_2921);
and UO_352 (O_352,N_2754,N_2785);
and UO_353 (O_353,N_2808,N_2352);
nor UO_354 (O_354,N_2835,N_2345);
nand UO_355 (O_355,N_2372,N_2274);
nand UO_356 (O_356,N_2530,N_2832);
and UO_357 (O_357,N_2798,N_2253);
nor UO_358 (O_358,N_2829,N_2462);
or UO_359 (O_359,N_2709,N_2469);
or UO_360 (O_360,N_2488,N_2872);
nor UO_361 (O_361,N_2688,N_2917);
or UO_362 (O_362,N_2793,N_2402);
and UO_363 (O_363,N_2875,N_2926);
or UO_364 (O_364,N_2371,N_2713);
nor UO_365 (O_365,N_2612,N_2268);
and UO_366 (O_366,N_2731,N_2678);
nand UO_367 (O_367,N_2815,N_2611);
nand UO_368 (O_368,N_2769,N_2853);
and UO_369 (O_369,N_2605,N_2621);
or UO_370 (O_370,N_2814,N_2340);
and UO_371 (O_371,N_2294,N_2682);
nand UO_372 (O_372,N_2995,N_2586);
nor UO_373 (O_373,N_2751,N_2395);
or UO_374 (O_374,N_2669,N_2797);
and UO_375 (O_375,N_2712,N_2350);
and UO_376 (O_376,N_2520,N_2749);
or UO_377 (O_377,N_2400,N_2858);
nor UO_378 (O_378,N_2349,N_2546);
or UO_379 (O_379,N_2503,N_2354);
nand UO_380 (O_380,N_2593,N_2472);
or UO_381 (O_381,N_2749,N_2801);
nor UO_382 (O_382,N_2394,N_2592);
or UO_383 (O_383,N_2799,N_2275);
nor UO_384 (O_384,N_2838,N_2857);
nand UO_385 (O_385,N_2960,N_2520);
or UO_386 (O_386,N_2613,N_2426);
nand UO_387 (O_387,N_2451,N_2775);
and UO_388 (O_388,N_2482,N_2951);
xor UO_389 (O_389,N_2725,N_2943);
nand UO_390 (O_390,N_2823,N_2657);
xor UO_391 (O_391,N_2353,N_2594);
nor UO_392 (O_392,N_2332,N_2315);
and UO_393 (O_393,N_2901,N_2709);
or UO_394 (O_394,N_2746,N_2855);
and UO_395 (O_395,N_2641,N_2392);
nand UO_396 (O_396,N_2714,N_2846);
or UO_397 (O_397,N_2471,N_2381);
nor UO_398 (O_398,N_2504,N_2988);
and UO_399 (O_399,N_2611,N_2330);
nand UO_400 (O_400,N_2886,N_2906);
xor UO_401 (O_401,N_2867,N_2306);
nand UO_402 (O_402,N_2847,N_2971);
nand UO_403 (O_403,N_2752,N_2698);
and UO_404 (O_404,N_2481,N_2976);
nand UO_405 (O_405,N_2256,N_2912);
and UO_406 (O_406,N_2697,N_2391);
and UO_407 (O_407,N_2345,N_2624);
and UO_408 (O_408,N_2324,N_2504);
and UO_409 (O_409,N_2422,N_2994);
or UO_410 (O_410,N_2677,N_2992);
and UO_411 (O_411,N_2544,N_2513);
nor UO_412 (O_412,N_2918,N_2258);
or UO_413 (O_413,N_2298,N_2309);
nor UO_414 (O_414,N_2749,N_2423);
nand UO_415 (O_415,N_2349,N_2778);
nor UO_416 (O_416,N_2681,N_2885);
nand UO_417 (O_417,N_2952,N_2766);
and UO_418 (O_418,N_2770,N_2651);
xnor UO_419 (O_419,N_2882,N_2470);
nor UO_420 (O_420,N_2544,N_2940);
nor UO_421 (O_421,N_2558,N_2954);
or UO_422 (O_422,N_2317,N_2448);
or UO_423 (O_423,N_2493,N_2696);
nor UO_424 (O_424,N_2559,N_2844);
nand UO_425 (O_425,N_2827,N_2692);
and UO_426 (O_426,N_2459,N_2373);
nor UO_427 (O_427,N_2597,N_2414);
nand UO_428 (O_428,N_2691,N_2411);
or UO_429 (O_429,N_2655,N_2573);
and UO_430 (O_430,N_2314,N_2496);
nor UO_431 (O_431,N_2302,N_2741);
nor UO_432 (O_432,N_2296,N_2559);
and UO_433 (O_433,N_2913,N_2393);
nor UO_434 (O_434,N_2741,N_2591);
or UO_435 (O_435,N_2458,N_2897);
or UO_436 (O_436,N_2586,N_2698);
or UO_437 (O_437,N_2635,N_2366);
xor UO_438 (O_438,N_2647,N_2542);
or UO_439 (O_439,N_2971,N_2620);
nor UO_440 (O_440,N_2348,N_2295);
or UO_441 (O_441,N_2444,N_2888);
or UO_442 (O_442,N_2862,N_2848);
nor UO_443 (O_443,N_2581,N_2823);
nor UO_444 (O_444,N_2318,N_2799);
nor UO_445 (O_445,N_2411,N_2294);
and UO_446 (O_446,N_2888,N_2324);
or UO_447 (O_447,N_2308,N_2781);
and UO_448 (O_448,N_2620,N_2958);
nand UO_449 (O_449,N_2514,N_2904);
or UO_450 (O_450,N_2319,N_2281);
nand UO_451 (O_451,N_2337,N_2663);
and UO_452 (O_452,N_2338,N_2722);
and UO_453 (O_453,N_2454,N_2520);
and UO_454 (O_454,N_2991,N_2861);
and UO_455 (O_455,N_2649,N_2301);
nand UO_456 (O_456,N_2455,N_2704);
or UO_457 (O_457,N_2774,N_2460);
or UO_458 (O_458,N_2922,N_2838);
nand UO_459 (O_459,N_2503,N_2335);
or UO_460 (O_460,N_2812,N_2934);
or UO_461 (O_461,N_2972,N_2849);
nor UO_462 (O_462,N_2797,N_2491);
nand UO_463 (O_463,N_2615,N_2705);
nor UO_464 (O_464,N_2539,N_2913);
or UO_465 (O_465,N_2761,N_2583);
and UO_466 (O_466,N_2476,N_2866);
nand UO_467 (O_467,N_2394,N_2330);
nand UO_468 (O_468,N_2629,N_2395);
nor UO_469 (O_469,N_2733,N_2766);
nor UO_470 (O_470,N_2932,N_2448);
and UO_471 (O_471,N_2701,N_2931);
or UO_472 (O_472,N_2985,N_2558);
nor UO_473 (O_473,N_2418,N_2775);
and UO_474 (O_474,N_2396,N_2810);
nand UO_475 (O_475,N_2920,N_2709);
nand UO_476 (O_476,N_2779,N_2938);
and UO_477 (O_477,N_2440,N_2411);
or UO_478 (O_478,N_2986,N_2989);
or UO_479 (O_479,N_2856,N_2906);
nor UO_480 (O_480,N_2291,N_2284);
and UO_481 (O_481,N_2569,N_2261);
and UO_482 (O_482,N_2685,N_2763);
or UO_483 (O_483,N_2463,N_2430);
nand UO_484 (O_484,N_2684,N_2510);
and UO_485 (O_485,N_2968,N_2495);
or UO_486 (O_486,N_2587,N_2844);
nand UO_487 (O_487,N_2352,N_2376);
nor UO_488 (O_488,N_2470,N_2746);
nor UO_489 (O_489,N_2581,N_2936);
nor UO_490 (O_490,N_2422,N_2840);
nor UO_491 (O_491,N_2461,N_2844);
and UO_492 (O_492,N_2969,N_2542);
and UO_493 (O_493,N_2890,N_2264);
nor UO_494 (O_494,N_2849,N_2353);
nor UO_495 (O_495,N_2689,N_2762);
nand UO_496 (O_496,N_2374,N_2678);
nor UO_497 (O_497,N_2532,N_2384);
or UO_498 (O_498,N_2355,N_2425);
nor UO_499 (O_499,N_2813,N_2332);
endmodule