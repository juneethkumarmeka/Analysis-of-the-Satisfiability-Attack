module basic_500_3000_500_60_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_357,In_277);
xor U1 (N_1,In_473,In_137);
and U2 (N_2,In_248,In_333);
nor U3 (N_3,In_208,In_356);
nor U4 (N_4,In_396,In_86);
nand U5 (N_5,In_401,In_47);
nor U6 (N_6,In_109,In_1);
and U7 (N_7,In_103,In_278);
nor U8 (N_8,In_451,In_328);
xnor U9 (N_9,In_92,In_161);
nor U10 (N_10,In_130,In_66);
nand U11 (N_11,In_339,In_38);
and U12 (N_12,In_432,In_308);
and U13 (N_13,In_496,In_468);
or U14 (N_14,In_337,In_414);
nand U15 (N_15,In_392,In_388);
nand U16 (N_16,In_228,In_409);
nand U17 (N_17,In_209,In_173);
and U18 (N_18,In_402,In_221);
or U19 (N_19,In_163,In_187);
and U20 (N_20,In_484,In_346);
and U21 (N_21,In_394,In_10);
and U22 (N_22,In_383,In_472);
nor U23 (N_23,In_342,In_4);
and U24 (N_24,In_483,In_118);
or U25 (N_25,In_223,In_139);
nand U26 (N_26,In_309,In_15);
and U27 (N_27,In_271,In_207);
nor U28 (N_28,In_138,In_23);
and U29 (N_29,In_379,In_3);
nand U30 (N_30,In_63,In_53);
and U31 (N_31,In_241,In_97);
and U32 (N_32,In_280,In_167);
and U33 (N_33,In_437,In_49);
or U34 (N_34,In_380,In_0);
and U35 (N_35,In_35,In_311);
and U36 (N_36,In_419,In_366);
and U37 (N_37,In_87,In_417);
nand U38 (N_38,In_205,In_332);
or U39 (N_39,In_41,In_36);
or U40 (N_40,In_470,In_194);
nand U41 (N_41,In_67,In_293);
and U42 (N_42,In_330,In_83);
nor U43 (N_43,In_327,In_183);
and U44 (N_44,In_324,In_261);
nor U45 (N_45,In_389,In_154);
or U46 (N_46,In_292,In_58);
and U47 (N_47,In_34,In_108);
xnor U48 (N_48,In_297,In_129);
and U49 (N_49,In_453,In_478);
or U50 (N_50,In_449,In_158);
nor U51 (N_51,In_263,N_38);
and U52 (N_52,In_233,In_412);
and U53 (N_53,In_82,In_40);
and U54 (N_54,In_455,In_436);
nand U55 (N_55,In_192,In_182);
or U56 (N_56,In_131,In_162);
or U57 (N_57,In_125,In_282);
nand U58 (N_58,In_81,N_26);
or U59 (N_59,In_290,N_3);
nand U60 (N_60,In_353,In_11);
and U61 (N_61,In_224,In_143);
xor U62 (N_62,In_377,In_22);
nand U63 (N_63,In_14,In_313);
and U64 (N_64,In_369,In_135);
nor U65 (N_65,In_355,In_464);
nor U66 (N_66,In_198,N_14);
or U67 (N_67,In_336,In_303);
or U68 (N_68,In_407,In_368);
and U69 (N_69,N_47,In_291);
nand U70 (N_70,In_331,In_210);
or U71 (N_71,In_361,In_146);
and U72 (N_72,In_239,In_364);
and U73 (N_73,N_1,In_150);
nand U74 (N_74,In_463,In_50);
and U75 (N_75,In_180,In_480);
nand U76 (N_76,In_301,In_430);
nand U77 (N_77,In_18,In_254);
nand U78 (N_78,N_16,In_111);
nand U79 (N_79,N_9,In_279);
and U80 (N_80,In_306,In_114);
nand U81 (N_81,In_200,In_80);
nor U82 (N_82,In_462,In_101);
or U83 (N_83,In_486,In_123);
or U84 (N_84,N_17,In_73);
xor U85 (N_85,In_127,In_85);
nand U86 (N_86,In_185,In_189);
nand U87 (N_87,In_244,In_262);
nor U88 (N_88,In_230,In_201);
and U89 (N_89,N_15,In_89);
nor U90 (N_90,In_155,In_323);
nor U91 (N_91,In_457,In_299);
or U92 (N_92,N_49,In_28);
and U93 (N_93,In_497,In_385);
or U94 (N_94,In_264,In_350);
or U95 (N_95,In_266,In_376);
and U96 (N_96,In_12,In_344);
or U97 (N_97,In_491,In_64);
nand U98 (N_98,In_382,In_477);
nor U99 (N_99,In_204,In_426);
nor U100 (N_100,In_226,In_159);
nand U101 (N_101,In_215,N_95);
and U102 (N_102,In_151,In_416);
or U103 (N_103,N_60,In_442);
nand U104 (N_104,In_257,In_287);
or U105 (N_105,In_235,N_84);
nor U106 (N_106,In_298,In_249);
or U107 (N_107,In_395,In_8);
or U108 (N_108,In_196,In_359);
nor U109 (N_109,In_141,In_460);
nor U110 (N_110,In_17,In_433);
or U111 (N_111,In_213,In_120);
nand U112 (N_112,N_66,In_142);
and U113 (N_113,N_36,In_343);
nand U114 (N_114,N_12,In_44);
nor U115 (N_115,In_95,In_267);
nand U116 (N_116,In_372,N_99);
nand U117 (N_117,In_397,In_145);
nor U118 (N_118,In_112,In_371);
nand U119 (N_119,In_466,N_78);
or U120 (N_120,In_321,In_218);
or U121 (N_121,In_485,In_126);
or U122 (N_122,In_77,In_160);
or U123 (N_123,N_4,N_87);
nor U124 (N_124,In_175,In_487);
nor U125 (N_125,In_493,N_41);
and U126 (N_126,N_56,In_5);
nor U127 (N_127,In_441,In_393);
nor U128 (N_128,In_481,In_273);
or U129 (N_129,In_166,In_322);
xor U130 (N_130,In_214,In_105);
or U131 (N_131,In_378,In_459);
or U132 (N_132,In_184,In_448);
nand U133 (N_133,In_72,In_59);
nand U134 (N_134,In_71,N_20);
and U135 (N_135,N_30,In_406);
nand U136 (N_136,N_51,N_69);
nand U137 (N_137,In_489,In_365);
and U138 (N_138,In_21,In_272);
or U139 (N_139,N_82,In_57);
and U140 (N_140,N_80,In_216);
xor U141 (N_141,In_467,In_398);
nand U142 (N_142,N_76,In_147);
or U143 (N_143,N_59,In_136);
xor U144 (N_144,N_34,In_69);
or U145 (N_145,N_71,In_269);
nor U146 (N_146,In_119,In_156);
and U147 (N_147,In_75,In_286);
nor U148 (N_148,In_461,In_107);
nand U149 (N_149,In_479,In_242);
and U150 (N_150,In_31,N_42);
nand U151 (N_151,In_65,In_128);
or U152 (N_152,N_115,In_312);
xor U153 (N_153,In_431,In_20);
nor U154 (N_154,In_317,N_117);
nor U155 (N_155,In_164,In_222);
and U156 (N_156,N_127,N_121);
nor U157 (N_157,In_176,In_229);
nor U158 (N_158,In_42,N_50);
xor U159 (N_159,N_136,N_114);
nor U160 (N_160,In_132,N_43);
and U161 (N_161,In_193,In_281);
and U162 (N_162,In_446,In_447);
nand U163 (N_163,In_240,N_29);
nor U164 (N_164,In_498,In_133);
nand U165 (N_165,N_2,In_51);
nor U166 (N_166,In_304,In_96);
xnor U167 (N_167,In_178,N_48);
and U168 (N_168,In_113,N_63);
or U169 (N_169,N_40,N_124);
nor U170 (N_170,In_29,In_423);
or U171 (N_171,In_212,In_275);
nand U172 (N_172,In_314,In_492);
or U173 (N_173,In_458,In_91);
and U174 (N_174,In_48,N_143);
nor U175 (N_175,In_310,In_102);
and U176 (N_176,In_220,N_104);
or U177 (N_177,In_338,N_11);
nand U178 (N_178,In_400,In_362);
nand U179 (N_179,In_68,N_53);
nand U180 (N_180,In_456,N_32);
nand U181 (N_181,In_219,N_141);
or U182 (N_182,N_138,In_227);
or U183 (N_183,In_19,In_370);
nand U184 (N_184,N_133,N_94);
or U185 (N_185,In_335,N_0);
nand U186 (N_186,In_435,N_86);
nand U187 (N_187,In_268,N_135);
nor U188 (N_188,In_347,In_302);
nand U189 (N_189,In_177,In_100);
or U190 (N_190,N_46,In_56);
nand U191 (N_191,In_39,In_148);
nor U192 (N_192,In_285,In_122);
nand U193 (N_193,In_315,N_70);
or U194 (N_194,In_255,In_46);
or U195 (N_195,In_427,In_172);
nand U196 (N_196,In_454,N_79);
nand U197 (N_197,In_84,In_251);
nand U198 (N_198,In_62,N_92);
nor U199 (N_199,In_345,In_384);
nor U200 (N_200,In_258,In_199);
nor U201 (N_201,In_116,In_60);
and U202 (N_202,In_300,In_289);
or U203 (N_203,In_231,N_64);
and U204 (N_204,In_413,In_482);
and U205 (N_205,In_358,In_94);
and U206 (N_206,In_16,N_6);
and U207 (N_207,N_128,N_179);
or U208 (N_208,N_184,In_334);
nor U209 (N_209,N_146,In_360);
nor U210 (N_210,N_93,In_367);
nor U211 (N_211,N_28,N_85);
nand U212 (N_212,N_123,N_90);
and U213 (N_213,N_52,In_474);
nand U214 (N_214,N_164,N_159);
nor U215 (N_215,In_326,In_43);
or U216 (N_216,N_24,In_2);
nor U217 (N_217,In_283,N_180);
nand U218 (N_218,N_166,N_198);
nor U219 (N_219,In_403,In_452);
nand U220 (N_220,N_174,N_190);
nor U221 (N_221,In_341,In_348);
and U222 (N_222,In_374,In_232);
or U223 (N_223,In_140,In_181);
nor U224 (N_224,In_90,N_96);
nand U225 (N_225,In_197,N_44);
or U226 (N_226,In_475,In_325);
or U227 (N_227,N_165,N_139);
and U228 (N_228,In_405,N_160);
or U229 (N_229,In_363,In_319);
nand U230 (N_230,N_155,N_37);
xor U231 (N_231,In_245,In_354);
xor U232 (N_232,N_107,In_296);
nor U233 (N_233,In_316,In_186);
or U234 (N_234,N_88,In_217);
nor U235 (N_235,N_112,N_142);
or U236 (N_236,In_55,In_418);
and U237 (N_237,N_170,In_259);
nor U238 (N_238,N_97,In_27);
or U239 (N_239,N_118,N_183);
nor U240 (N_240,N_116,N_108);
or U241 (N_241,N_176,In_117);
nand U242 (N_242,In_121,N_18);
xor U243 (N_243,In_76,In_421);
nor U244 (N_244,In_115,N_81);
nand U245 (N_245,In_190,In_33);
nor U246 (N_246,N_109,In_247);
nand U247 (N_247,N_129,In_351);
and U248 (N_248,In_195,In_408);
nand U249 (N_249,In_499,N_103);
nand U250 (N_250,N_236,In_349);
and U251 (N_251,N_163,N_77);
or U252 (N_252,N_45,N_226);
or U253 (N_253,In_434,N_153);
or U254 (N_254,In_93,N_227);
nand U255 (N_255,In_265,In_25);
and U256 (N_256,In_381,N_207);
and U257 (N_257,In_250,In_352);
and U258 (N_258,N_58,In_444);
and U259 (N_259,N_231,N_62);
or U260 (N_260,In_26,In_104);
nand U261 (N_261,N_206,N_235);
or U262 (N_262,N_187,N_229);
nand U263 (N_263,N_185,N_151);
nand U264 (N_264,N_222,N_230);
nand U265 (N_265,N_119,N_172);
or U266 (N_266,In_404,N_175);
nor U267 (N_267,In_243,N_61);
and U268 (N_268,N_186,N_213);
nor U269 (N_269,N_39,In_420);
nand U270 (N_270,In_422,In_6);
nor U271 (N_271,In_74,In_238);
or U272 (N_272,N_238,N_102);
or U273 (N_273,N_137,In_438);
and U274 (N_274,In_234,N_234);
nand U275 (N_275,In_157,N_157);
and U276 (N_276,In_490,N_7);
or U277 (N_277,N_110,N_98);
nand U278 (N_278,N_177,In_424);
or U279 (N_279,In_70,N_246);
nand U280 (N_280,N_31,N_147);
nand U281 (N_281,N_73,N_74);
nor U282 (N_282,In_99,N_245);
or U283 (N_283,N_21,In_152);
and U284 (N_284,N_168,N_232);
nor U285 (N_285,N_65,N_202);
nand U286 (N_286,In_274,N_144);
nor U287 (N_287,In_439,N_192);
nand U288 (N_288,N_239,N_249);
or U289 (N_289,In_110,In_260);
and U290 (N_290,N_134,In_288);
or U291 (N_291,N_220,In_165);
and U292 (N_292,N_126,In_428);
nand U293 (N_293,N_125,In_24);
and U294 (N_294,In_494,N_23);
or U295 (N_295,In_387,N_162);
nor U296 (N_296,N_150,In_54);
nand U297 (N_297,In_153,N_225);
nor U298 (N_298,In_399,N_203);
or U299 (N_299,N_194,N_195);
nor U300 (N_300,N_149,N_278);
nand U301 (N_301,N_256,N_154);
nor U302 (N_302,N_27,N_158);
nand U303 (N_303,N_221,N_264);
and U304 (N_304,N_237,N_75);
and U305 (N_305,In_276,N_72);
and U306 (N_306,In_32,N_274);
xnor U307 (N_307,N_291,N_279);
and U308 (N_308,In_124,N_171);
nor U309 (N_309,In_270,N_210);
nand U310 (N_310,N_156,N_285);
nor U311 (N_311,In_471,N_215);
nor U312 (N_312,In_410,N_233);
and U313 (N_313,In_169,In_225);
nor U314 (N_314,N_167,N_91);
nor U315 (N_315,In_429,N_189);
xnor U316 (N_316,N_259,N_5);
nand U317 (N_317,N_260,In_373);
nor U318 (N_318,N_265,In_295);
nor U319 (N_319,In_37,In_61);
and U320 (N_320,In_106,N_113);
nand U321 (N_321,N_282,In_203);
nor U322 (N_322,In_284,In_390);
or U323 (N_323,In_236,In_329);
or U324 (N_324,In_294,N_223);
and U325 (N_325,In_191,N_57);
or U326 (N_326,In_445,N_55);
or U327 (N_327,In_88,N_100);
nor U328 (N_328,In_211,N_297);
or U329 (N_329,In_174,N_273);
nand U330 (N_330,N_196,N_275);
or U331 (N_331,N_131,N_288);
or U332 (N_332,N_199,In_7);
nand U333 (N_333,In_386,N_205);
or U334 (N_334,N_105,In_476);
and U335 (N_335,N_188,In_488);
nor U336 (N_336,In_78,N_270);
nor U337 (N_337,In_206,N_204);
nand U338 (N_338,N_284,N_271);
nand U339 (N_339,N_268,N_286);
or U340 (N_340,In_495,N_290);
and U341 (N_341,N_280,N_251);
nor U342 (N_342,N_68,N_145);
or U343 (N_343,N_208,In_144);
and U344 (N_344,In_237,N_292);
or U345 (N_345,N_54,N_106);
nand U346 (N_346,In_253,In_134);
xnor U347 (N_347,N_228,N_178);
nand U348 (N_348,In_98,N_182);
nand U349 (N_349,In_391,N_218);
or U350 (N_350,N_314,N_338);
and U351 (N_351,N_120,N_262);
nor U352 (N_352,In_320,N_255);
and U353 (N_353,N_212,N_267);
nand U354 (N_354,N_311,N_348);
nand U355 (N_355,N_122,N_306);
nor U356 (N_356,In_375,N_266);
or U357 (N_357,N_209,In_318);
nand U358 (N_358,N_248,In_425);
or U359 (N_359,N_345,N_253);
and U360 (N_360,N_294,In_443);
and U361 (N_361,In_469,N_303);
nand U362 (N_362,In_252,N_341);
and U363 (N_363,N_272,N_10);
or U364 (N_364,N_241,In_52);
and U365 (N_365,N_325,N_219);
or U366 (N_366,N_258,In_411);
nand U367 (N_367,N_200,N_343);
and U368 (N_368,N_324,N_252);
nand U369 (N_369,N_315,N_216);
nand U370 (N_370,N_250,N_211);
nor U371 (N_371,N_217,N_327);
nand U372 (N_372,N_330,N_313);
nand U373 (N_373,N_140,In_45);
and U374 (N_374,In_171,N_302);
and U375 (N_375,N_269,In_79);
nand U376 (N_376,N_201,N_169);
or U377 (N_377,N_224,N_67);
nor U378 (N_378,N_342,In_168);
nand U379 (N_379,N_254,N_243);
or U380 (N_380,In_13,In_149);
and U381 (N_381,In_465,N_308);
nand U382 (N_382,N_335,In_9);
nor U383 (N_383,N_331,N_333);
and U384 (N_384,N_25,N_35);
nor U385 (N_385,In_202,N_191);
and U386 (N_386,In_307,N_277);
or U387 (N_387,N_310,N_289);
and U388 (N_388,In_179,N_317);
nor U389 (N_389,N_329,N_22);
or U390 (N_390,N_349,N_332);
or U391 (N_391,N_283,N_161);
nand U392 (N_392,N_276,In_256);
or U393 (N_393,In_30,N_300);
and U394 (N_394,N_316,In_246);
nand U395 (N_395,In_440,N_89);
and U396 (N_396,N_320,N_257);
nand U397 (N_397,N_111,N_130);
and U398 (N_398,N_8,N_287);
and U399 (N_399,N_101,In_170);
nor U400 (N_400,N_336,N_399);
nor U401 (N_401,N_344,N_375);
and U402 (N_402,N_304,N_387);
xnor U403 (N_403,N_334,N_193);
or U404 (N_404,N_197,N_378);
and U405 (N_405,N_381,N_366);
or U406 (N_406,N_312,N_328);
nand U407 (N_407,N_152,N_244);
nand U408 (N_408,N_355,N_181);
nor U409 (N_409,N_19,N_353);
and U410 (N_410,N_340,N_379);
nand U411 (N_411,N_13,N_326);
nor U412 (N_412,N_356,N_318);
nor U413 (N_413,N_322,N_392);
xnor U414 (N_414,In_450,N_364);
or U415 (N_415,N_309,N_382);
nand U416 (N_416,N_359,N_307);
or U417 (N_417,N_367,N_296);
and U418 (N_418,N_373,N_240);
nand U419 (N_419,N_354,N_369);
nor U420 (N_420,In_188,N_33);
and U421 (N_421,N_363,N_261);
nor U422 (N_422,N_281,N_380);
or U423 (N_423,N_383,In_340);
and U424 (N_424,N_148,N_337);
nand U425 (N_425,N_214,N_346);
or U426 (N_426,N_397,N_173);
nand U427 (N_427,N_394,N_391);
nor U428 (N_428,N_352,N_298);
and U429 (N_429,N_351,N_395);
and U430 (N_430,N_374,N_372);
or U431 (N_431,N_339,N_299);
and U432 (N_432,N_386,N_389);
nand U433 (N_433,In_305,N_293);
and U434 (N_434,N_370,N_295);
or U435 (N_435,N_319,N_242);
xor U436 (N_436,N_376,N_377);
nand U437 (N_437,N_323,N_347);
nor U438 (N_438,N_83,N_368);
nand U439 (N_439,N_301,N_350);
and U440 (N_440,N_384,N_263);
and U441 (N_441,N_357,In_415);
and U442 (N_442,N_393,N_390);
and U443 (N_443,N_398,N_385);
nor U444 (N_444,N_365,N_371);
nor U445 (N_445,N_305,N_396);
nand U446 (N_446,N_388,N_321);
nand U447 (N_447,N_360,N_132);
and U448 (N_448,N_358,N_362);
and U449 (N_449,N_247,N_361);
and U450 (N_450,N_435,N_415);
nand U451 (N_451,N_438,N_421);
nor U452 (N_452,N_411,N_431);
or U453 (N_453,N_410,N_442);
and U454 (N_454,N_423,N_443);
and U455 (N_455,N_432,N_422);
and U456 (N_456,N_424,N_412);
or U457 (N_457,N_418,N_408);
nand U458 (N_458,N_449,N_403);
nor U459 (N_459,N_416,N_430);
or U460 (N_460,N_426,N_407);
and U461 (N_461,N_441,N_445);
nor U462 (N_462,N_446,N_440);
and U463 (N_463,N_417,N_402);
nand U464 (N_464,N_448,N_429);
nor U465 (N_465,N_400,N_425);
and U466 (N_466,N_436,N_428);
or U467 (N_467,N_427,N_439);
nand U468 (N_468,N_401,N_419);
or U469 (N_469,N_434,N_444);
and U470 (N_470,N_447,N_409);
or U471 (N_471,N_406,N_413);
and U472 (N_472,N_433,N_437);
or U473 (N_473,N_414,N_405);
nor U474 (N_474,N_404,N_420);
nand U475 (N_475,N_423,N_448);
and U476 (N_476,N_447,N_407);
and U477 (N_477,N_420,N_440);
and U478 (N_478,N_401,N_434);
or U479 (N_479,N_418,N_447);
or U480 (N_480,N_447,N_420);
nand U481 (N_481,N_440,N_427);
and U482 (N_482,N_419,N_443);
and U483 (N_483,N_400,N_441);
nand U484 (N_484,N_418,N_436);
nand U485 (N_485,N_414,N_434);
and U486 (N_486,N_407,N_434);
nand U487 (N_487,N_437,N_424);
nor U488 (N_488,N_428,N_410);
nand U489 (N_489,N_415,N_405);
nor U490 (N_490,N_408,N_430);
nor U491 (N_491,N_449,N_423);
and U492 (N_492,N_444,N_429);
and U493 (N_493,N_405,N_444);
or U494 (N_494,N_442,N_407);
or U495 (N_495,N_405,N_413);
nand U496 (N_496,N_441,N_446);
and U497 (N_497,N_413,N_407);
or U498 (N_498,N_401,N_406);
xnor U499 (N_499,N_427,N_403);
nand U500 (N_500,N_477,N_474);
and U501 (N_501,N_450,N_494);
nand U502 (N_502,N_485,N_495);
nor U503 (N_503,N_490,N_462);
and U504 (N_504,N_472,N_493);
xor U505 (N_505,N_498,N_497);
nor U506 (N_506,N_481,N_480);
nor U507 (N_507,N_475,N_469);
and U508 (N_508,N_478,N_491);
nand U509 (N_509,N_487,N_457);
nand U510 (N_510,N_451,N_465);
nand U511 (N_511,N_482,N_467);
xor U512 (N_512,N_479,N_459);
nor U513 (N_513,N_483,N_486);
nand U514 (N_514,N_455,N_471);
and U515 (N_515,N_489,N_468);
nand U516 (N_516,N_460,N_466);
and U517 (N_517,N_453,N_454);
nor U518 (N_518,N_456,N_458);
and U519 (N_519,N_484,N_464);
and U520 (N_520,N_461,N_463);
nand U521 (N_521,N_492,N_496);
nor U522 (N_522,N_470,N_476);
nor U523 (N_523,N_452,N_473);
nor U524 (N_524,N_499,N_488);
or U525 (N_525,N_469,N_456);
nand U526 (N_526,N_465,N_487);
nand U527 (N_527,N_485,N_484);
nor U528 (N_528,N_482,N_484);
nand U529 (N_529,N_468,N_459);
nand U530 (N_530,N_468,N_470);
and U531 (N_531,N_479,N_481);
and U532 (N_532,N_499,N_495);
and U533 (N_533,N_491,N_471);
nor U534 (N_534,N_458,N_459);
nand U535 (N_535,N_460,N_458);
or U536 (N_536,N_475,N_453);
nand U537 (N_537,N_466,N_473);
or U538 (N_538,N_492,N_457);
xnor U539 (N_539,N_478,N_460);
and U540 (N_540,N_485,N_463);
nor U541 (N_541,N_489,N_487);
and U542 (N_542,N_469,N_460);
or U543 (N_543,N_482,N_486);
or U544 (N_544,N_466,N_462);
nor U545 (N_545,N_476,N_460);
or U546 (N_546,N_455,N_450);
nand U547 (N_547,N_491,N_457);
nand U548 (N_548,N_465,N_455);
or U549 (N_549,N_495,N_460);
or U550 (N_550,N_543,N_521);
or U551 (N_551,N_528,N_544);
nor U552 (N_552,N_520,N_540);
and U553 (N_553,N_518,N_546);
and U554 (N_554,N_534,N_505);
nor U555 (N_555,N_512,N_530);
xnor U556 (N_556,N_523,N_527);
nand U557 (N_557,N_542,N_535);
or U558 (N_558,N_506,N_513);
and U559 (N_559,N_537,N_525);
and U560 (N_560,N_547,N_504);
nor U561 (N_561,N_502,N_541);
and U562 (N_562,N_545,N_503);
nand U563 (N_563,N_515,N_508);
or U564 (N_564,N_514,N_526);
xor U565 (N_565,N_532,N_536);
nand U566 (N_566,N_517,N_500);
nor U567 (N_567,N_538,N_549);
and U568 (N_568,N_509,N_529);
nor U569 (N_569,N_524,N_501);
or U570 (N_570,N_548,N_510);
nand U571 (N_571,N_539,N_516);
nand U572 (N_572,N_522,N_507);
xnor U573 (N_573,N_533,N_531);
nand U574 (N_574,N_519,N_511);
and U575 (N_575,N_539,N_546);
nor U576 (N_576,N_527,N_546);
nor U577 (N_577,N_544,N_536);
or U578 (N_578,N_501,N_515);
and U579 (N_579,N_522,N_546);
nand U580 (N_580,N_538,N_547);
or U581 (N_581,N_535,N_544);
and U582 (N_582,N_549,N_519);
nor U583 (N_583,N_516,N_549);
nor U584 (N_584,N_521,N_509);
or U585 (N_585,N_548,N_530);
nand U586 (N_586,N_530,N_520);
nand U587 (N_587,N_543,N_527);
and U588 (N_588,N_529,N_508);
nand U589 (N_589,N_510,N_504);
or U590 (N_590,N_533,N_519);
and U591 (N_591,N_503,N_505);
and U592 (N_592,N_531,N_540);
or U593 (N_593,N_529,N_524);
nor U594 (N_594,N_535,N_506);
nor U595 (N_595,N_546,N_534);
and U596 (N_596,N_532,N_534);
and U597 (N_597,N_510,N_520);
or U598 (N_598,N_537,N_536);
and U599 (N_599,N_516,N_524);
nand U600 (N_600,N_552,N_565);
or U601 (N_601,N_596,N_566);
and U602 (N_602,N_568,N_557);
nor U603 (N_603,N_564,N_584);
nand U604 (N_604,N_583,N_585);
or U605 (N_605,N_567,N_577);
nor U606 (N_606,N_588,N_595);
nor U607 (N_607,N_582,N_576);
nand U608 (N_608,N_570,N_581);
nor U609 (N_609,N_573,N_559);
xnor U610 (N_610,N_574,N_589);
nand U611 (N_611,N_590,N_579);
or U612 (N_612,N_578,N_575);
nor U613 (N_613,N_571,N_554);
or U614 (N_614,N_563,N_586);
and U615 (N_615,N_550,N_597);
or U616 (N_616,N_594,N_562);
nor U617 (N_617,N_580,N_556);
xor U618 (N_618,N_555,N_587);
or U619 (N_619,N_593,N_551);
nor U620 (N_620,N_572,N_569);
nor U621 (N_621,N_553,N_599);
nor U622 (N_622,N_592,N_558);
and U623 (N_623,N_598,N_560);
nor U624 (N_624,N_591,N_561);
nand U625 (N_625,N_558,N_578);
nand U626 (N_626,N_597,N_577);
or U627 (N_627,N_558,N_588);
or U628 (N_628,N_582,N_558);
nand U629 (N_629,N_553,N_594);
and U630 (N_630,N_559,N_586);
nand U631 (N_631,N_565,N_553);
nand U632 (N_632,N_587,N_588);
and U633 (N_633,N_577,N_564);
or U634 (N_634,N_575,N_557);
nand U635 (N_635,N_563,N_571);
xor U636 (N_636,N_554,N_559);
nor U637 (N_637,N_565,N_599);
and U638 (N_638,N_594,N_576);
or U639 (N_639,N_581,N_590);
or U640 (N_640,N_562,N_569);
nand U641 (N_641,N_598,N_556);
and U642 (N_642,N_559,N_585);
nand U643 (N_643,N_594,N_567);
nand U644 (N_644,N_555,N_589);
and U645 (N_645,N_576,N_586);
or U646 (N_646,N_557,N_593);
nand U647 (N_647,N_583,N_570);
nor U648 (N_648,N_554,N_597);
nor U649 (N_649,N_563,N_587);
nor U650 (N_650,N_625,N_603);
or U651 (N_651,N_617,N_630);
or U652 (N_652,N_605,N_648);
and U653 (N_653,N_637,N_613);
nor U654 (N_654,N_646,N_620);
and U655 (N_655,N_618,N_608);
nand U656 (N_656,N_643,N_629);
nor U657 (N_657,N_641,N_614);
and U658 (N_658,N_610,N_635);
or U659 (N_659,N_647,N_622);
nand U660 (N_660,N_611,N_640);
or U661 (N_661,N_627,N_604);
or U662 (N_662,N_649,N_631);
or U663 (N_663,N_619,N_639);
or U664 (N_664,N_602,N_638);
nor U665 (N_665,N_621,N_600);
nand U666 (N_666,N_624,N_632);
nor U667 (N_667,N_628,N_623);
nand U668 (N_668,N_615,N_642);
nor U669 (N_669,N_626,N_645);
or U670 (N_670,N_644,N_633);
or U671 (N_671,N_609,N_634);
and U672 (N_672,N_607,N_616);
xor U673 (N_673,N_601,N_636);
nand U674 (N_674,N_606,N_612);
nand U675 (N_675,N_608,N_641);
or U676 (N_676,N_607,N_637);
or U677 (N_677,N_647,N_614);
nor U678 (N_678,N_627,N_645);
nor U679 (N_679,N_609,N_631);
and U680 (N_680,N_616,N_636);
or U681 (N_681,N_645,N_642);
and U682 (N_682,N_610,N_611);
nand U683 (N_683,N_616,N_624);
or U684 (N_684,N_620,N_644);
and U685 (N_685,N_631,N_616);
nor U686 (N_686,N_641,N_647);
and U687 (N_687,N_648,N_633);
and U688 (N_688,N_633,N_618);
or U689 (N_689,N_631,N_640);
xnor U690 (N_690,N_628,N_602);
or U691 (N_691,N_624,N_614);
nand U692 (N_692,N_612,N_631);
nor U693 (N_693,N_638,N_603);
nor U694 (N_694,N_605,N_635);
or U695 (N_695,N_616,N_632);
or U696 (N_696,N_606,N_610);
xor U697 (N_697,N_605,N_617);
and U698 (N_698,N_618,N_630);
nand U699 (N_699,N_604,N_645);
nand U700 (N_700,N_652,N_678);
nand U701 (N_701,N_670,N_681);
or U702 (N_702,N_693,N_655);
nand U703 (N_703,N_675,N_691);
nor U704 (N_704,N_673,N_665);
and U705 (N_705,N_689,N_658);
nand U706 (N_706,N_653,N_669);
nor U707 (N_707,N_654,N_695);
nand U708 (N_708,N_662,N_668);
nor U709 (N_709,N_680,N_686);
nand U710 (N_710,N_674,N_676);
or U711 (N_711,N_672,N_697);
xor U712 (N_712,N_666,N_677);
or U713 (N_713,N_688,N_679);
or U714 (N_714,N_650,N_659);
and U715 (N_715,N_685,N_661);
nand U716 (N_716,N_651,N_667);
or U717 (N_717,N_696,N_663);
and U718 (N_718,N_694,N_682);
nor U719 (N_719,N_684,N_692);
xnor U720 (N_720,N_698,N_671);
and U721 (N_721,N_660,N_657);
nor U722 (N_722,N_656,N_683);
nand U723 (N_723,N_690,N_699);
nor U724 (N_724,N_687,N_664);
or U725 (N_725,N_695,N_679);
nor U726 (N_726,N_681,N_679);
and U727 (N_727,N_699,N_668);
nor U728 (N_728,N_694,N_652);
and U729 (N_729,N_675,N_654);
or U730 (N_730,N_673,N_687);
nand U731 (N_731,N_669,N_683);
nor U732 (N_732,N_664,N_696);
or U733 (N_733,N_691,N_680);
nand U734 (N_734,N_683,N_665);
nor U735 (N_735,N_683,N_676);
nor U736 (N_736,N_690,N_650);
nor U737 (N_737,N_694,N_677);
and U738 (N_738,N_655,N_675);
or U739 (N_739,N_668,N_654);
or U740 (N_740,N_651,N_692);
nor U741 (N_741,N_691,N_659);
or U742 (N_742,N_659,N_672);
or U743 (N_743,N_697,N_685);
and U744 (N_744,N_659,N_668);
or U745 (N_745,N_666,N_687);
or U746 (N_746,N_694,N_672);
or U747 (N_747,N_670,N_680);
and U748 (N_748,N_667,N_665);
or U749 (N_749,N_653,N_667);
nor U750 (N_750,N_726,N_734);
nor U751 (N_751,N_740,N_711);
xnor U752 (N_752,N_716,N_744);
and U753 (N_753,N_707,N_737);
and U754 (N_754,N_742,N_730);
nand U755 (N_755,N_700,N_743);
nor U756 (N_756,N_724,N_747);
nor U757 (N_757,N_725,N_727);
nand U758 (N_758,N_708,N_729);
xnor U759 (N_759,N_749,N_710);
nor U760 (N_760,N_703,N_731);
and U761 (N_761,N_712,N_718);
or U762 (N_762,N_704,N_705);
nor U763 (N_763,N_733,N_701);
xor U764 (N_764,N_738,N_722);
nor U765 (N_765,N_748,N_715);
nor U766 (N_766,N_723,N_736);
and U767 (N_767,N_732,N_735);
nor U768 (N_768,N_717,N_719);
or U769 (N_769,N_746,N_713);
nand U770 (N_770,N_728,N_720);
or U771 (N_771,N_745,N_709);
and U772 (N_772,N_702,N_741);
and U773 (N_773,N_714,N_721);
nor U774 (N_774,N_739,N_706);
and U775 (N_775,N_712,N_709);
or U776 (N_776,N_742,N_748);
and U777 (N_777,N_704,N_742);
nor U778 (N_778,N_711,N_717);
or U779 (N_779,N_708,N_701);
nor U780 (N_780,N_710,N_713);
and U781 (N_781,N_724,N_714);
or U782 (N_782,N_745,N_702);
nand U783 (N_783,N_700,N_701);
or U784 (N_784,N_724,N_728);
or U785 (N_785,N_704,N_712);
or U786 (N_786,N_745,N_716);
nand U787 (N_787,N_725,N_731);
nor U788 (N_788,N_747,N_723);
and U789 (N_789,N_714,N_728);
or U790 (N_790,N_720,N_701);
nor U791 (N_791,N_706,N_745);
nand U792 (N_792,N_721,N_719);
and U793 (N_793,N_741,N_717);
and U794 (N_794,N_731,N_738);
or U795 (N_795,N_746,N_722);
nor U796 (N_796,N_721,N_727);
nor U797 (N_797,N_704,N_717);
nand U798 (N_798,N_709,N_724);
nor U799 (N_799,N_732,N_749);
nand U800 (N_800,N_759,N_788);
nand U801 (N_801,N_780,N_781);
or U802 (N_802,N_776,N_762);
and U803 (N_803,N_798,N_782);
and U804 (N_804,N_757,N_787);
nand U805 (N_805,N_789,N_766);
nor U806 (N_806,N_772,N_791);
nor U807 (N_807,N_769,N_751);
xnor U808 (N_808,N_773,N_768);
or U809 (N_809,N_794,N_771);
and U810 (N_810,N_778,N_783);
or U811 (N_811,N_796,N_799);
and U812 (N_812,N_774,N_767);
nand U813 (N_813,N_764,N_761);
nand U814 (N_814,N_753,N_793);
or U815 (N_815,N_784,N_777);
and U816 (N_816,N_754,N_763);
and U817 (N_817,N_790,N_775);
nand U818 (N_818,N_779,N_765);
nand U819 (N_819,N_760,N_797);
or U820 (N_820,N_770,N_795);
or U821 (N_821,N_750,N_752);
or U822 (N_822,N_792,N_756);
nor U823 (N_823,N_755,N_785);
and U824 (N_824,N_758,N_786);
or U825 (N_825,N_767,N_781);
nand U826 (N_826,N_757,N_762);
nor U827 (N_827,N_790,N_784);
or U828 (N_828,N_763,N_772);
and U829 (N_829,N_796,N_782);
nand U830 (N_830,N_750,N_773);
and U831 (N_831,N_761,N_759);
nand U832 (N_832,N_776,N_790);
nor U833 (N_833,N_785,N_790);
nand U834 (N_834,N_776,N_795);
and U835 (N_835,N_785,N_799);
nor U836 (N_836,N_790,N_767);
or U837 (N_837,N_796,N_772);
and U838 (N_838,N_787,N_781);
or U839 (N_839,N_797,N_783);
and U840 (N_840,N_755,N_779);
or U841 (N_841,N_783,N_775);
or U842 (N_842,N_793,N_750);
and U843 (N_843,N_753,N_765);
xnor U844 (N_844,N_758,N_759);
nor U845 (N_845,N_787,N_752);
nand U846 (N_846,N_757,N_763);
or U847 (N_847,N_754,N_751);
and U848 (N_848,N_793,N_767);
and U849 (N_849,N_795,N_783);
nor U850 (N_850,N_805,N_813);
nor U851 (N_851,N_826,N_824);
and U852 (N_852,N_808,N_831);
nand U853 (N_853,N_817,N_835);
or U854 (N_854,N_818,N_811);
or U855 (N_855,N_841,N_819);
nor U856 (N_856,N_846,N_845);
and U857 (N_857,N_823,N_802);
nor U858 (N_858,N_810,N_840);
nand U859 (N_859,N_833,N_839);
or U860 (N_860,N_803,N_815);
or U861 (N_861,N_847,N_801);
nor U862 (N_862,N_842,N_838);
or U863 (N_863,N_836,N_843);
or U864 (N_864,N_821,N_812);
and U865 (N_865,N_814,N_809);
nor U866 (N_866,N_825,N_827);
nand U867 (N_867,N_834,N_844);
nand U868 (N_868,N_848,N_816);
nor U869 (N_869,N_828,N_807);
nand U870 (N_870,N_820,N_837);
or U871 (N_871,N_804,N_832);
nand U872 (N_872,N_806,N_830);
nor U873 (N_873,N_849,N_822);
nand U874 (N_874,N_800,N_829);
or U875 (N_875,N_819,N_825);
or U876 (N_876,N_804,N_825);
or U877 (N_877,N_823,N_836);
nor U878 (N_878,N_846,N_843);
and U879 (N_879,N_832,N_810);
or U880 (N_880,N_811,N_806);
and U881 (N_881,N_846,N_800);
or U882 (N_882,N_849,N_830);
or U883 (N_883,N_842,N_846);
or U884 (N_884,N_825,N_848);
or U885 (N_885,N_805,N_847);
nand U886 (N_886,N_828,N_839);
and U887 (N_887,N_833,N_834);
and U888 (N_888,N_807,N_823);
and U889 (N_889,N_844,N_827);
or U890 (N_890,N_824,N_829);
and U891 (N_891,N_839,N_802);
nand U892 (N_892,N_844,N_810);
nor U893 (N_893,N_830,N_827);
nand U894 (N_894,N_823,N_839);
nor U895 (N_895,N_802,N_807);
nor U896 (N_896,N_842,N_817);
nand U897 (N_897,N_822,N_833);
or U898 (N_898,N_842,N_840);
or U899 (N_899,N_840,N_811);
or U900 (N_900,N_894,N_883);
nand U901 (N_901,N_869,N_873);
nand U902 (N_902,N_877,N_898);
and U903 (N_903,N_863,N_885);
nand U904 (N_904,N_855,N_889);
and U905 (N_905,N_851,N_882);
nand U906 (N_906,N_868,N_881);
or U907 (N_907,N_893,N_870);
nor U908 (N_908,N_864,N_892);
and U909 (N_909,N_856,N_876);
or U910 (N_910,N_861,N_858);
and U911 (N_911,N_865,N_899);
and U912 (N_912,N_871,N_860);
nor U913 (N_913,N_850,N_862);
and U914 (N_914,N_888,N_886);
or U915 (N_915,N_857,N_875);
nand U916 (N_916,N_853,N_887);
nand U917 (N_917,N_866,N_854);
or U918 (N_918,N_874,N_890);
or U919 (N_919,N_872,N_879);
and U920 (N_920,N_895,N_897);
nor U921 (N_921,N_852,N_884);
nor U922 (N_922,N_880,N_867);
and U923 (N_923,N_878,N_859);
and U924 (N_924,N_896,N_891);
and U925 (N_925,N_886,N_885);
or U926 (N_926,N_854,N_877);
or U927 (N_927,N_858,N_886);
and U928 (N_928,N_877,N_851);
and U929 (N_929,N_852,N_850);
and U930 (N_930,N_888,N_882);
nor U931 (N_931,N_888,N_853);
nor U932 (N_932,N_897,N_859);
nand U933 (N_933,N_897,N_858);
nor U934 (N_934,N_864,N_898);
and U935 (N_935,N_859,N_890);
nand U936 (N_936,N_853,N_886);
or U937 (N_937,N_861,N_872);
nor U938 (N_938,N_892,N_890);
and U939 (N_939,N_875,N_883);
and U940 (N_940,N_860,N_861);
and U941 (N_941,N_866,N_893);
or U942 (N_942,N_868,N_852);
and U943 (N_943,N_869,N_878);
and U944 (N_944,N_858,N_852);
and U945 (N_945,N_885,N_894);
nand U946 (N_946,N_862,N_868);
and U947 (N_947,N_882,N_876);
nand U948 (N_948,N_893,N_861);
or U949 (N_949,N_873,N_854);
or U950 (N_950,N_938,N_949);
nor U951 (N_951,N_905,N_929);
nand U952 (N_952,N_917,N_935);
xnor U953 (N_953,N_916,N_921);
or U954 (N_954,N_927,N_907);
nand U955 (N_955,N_922,N_902);
and U956 (N_956,N_909,N_933);
nand U957 (N_957,N_913,N_906);
nor U958 (N_958,N_945,N_943);
and U959 (N_959,N_940,N_926);
or U960 (N_960,N_920,N_930);
or U961 (N_961,N_942,N_919);
xor U962 (N_962,N_904,N_944);
and U963 (N_963,N_903,N_910);
or U964 (N_964,N_923,N_932);
and U965 (N_965,N_914,N_936);
and U966 (N_966,N_931,N_947);
and U967 (N_967,N_924,N_915);
or U968 (N_968,N_900,N_928);
nor U969 (N_969,N_918,N_901);
nor U970 (N_970,N_934,N_939);
nor U971 (N_971,N_925,N_908);
and U972 (N_972,N_911,N_941);
nor U973 (N_973,N_946,N_948);
or U974 (N_974,N_937,N_912);
and U975 (N_975,N_934,N_917);
nor U976 (N_976,N_948,N_920);
or U977 (N_977,N_907,N_919);
and U978 (N_978,N_921,N_920);
nand U979 (N_979,N_911,N_942);
nor U980 (N_980,N_931,N_908);
nor U981 (N_981,N_940,N_914);
nand U982 (N_982,N_901,N_940);
nor U983 (N_983,N_909,N_912);
nand U984 (N_984,N_923,N_903);
or U985 (N_985,N_925,N_934);
and U986 (N_986,N_941,N_908);
nor U987 (N_987,N_905,N_906);
and U988 (N_988,N_921,N_914);
nor U989 (N_989,N_920,N_918);
and U990 (N_990,N_902,N_935);
or U991 (N_991,N_919,N_947);
or U992 (N_992,N_926,N_948);
nor U993 (N_993,N_915,N_940);
and U994 (N_994,N_931,N_915);
or U995 (N_995,N_925,N_921);
and U996 (N_996,N_930,N_919);
nor U997 (N_997,N_904,N_922);
and U998 (N_998,N_906,N_939);
and U999 (N_999,N_948,N_932);
nor U1000 (N_1000,N_952,N_959);
or U1001 (N_1001,N_982,N_980);
or U1002 (N_1002,N_955,N_966);
nor U1003 (N_1003,N_951,N_994);
nor U1004 (N_1004,N_979,N_989);
nor U1005 (N_1005,N_968,N_976);
and U1006 (N_1006,N_961,N_970);
nor U1007 (N_1007,N_999,N_975);
or U1008 (N_1008,N_995,N_954);
and U1009 (N_1009,N_974,N_988);
and U1010 (N_1010,N_986,N_991);
nand U1011 (N_1011,N_969,N_978);
or U1012 (N_1012,N_985,N_993);
or U1013 (N_1013,N_958,N_987);
or U1014 (N_1014,N_997,N_983);
and U1015 (N_1015,N_964,N_956);
nor U1016 (N_1016,N_998,N_953);
nor U1017 (N_1017,N_963,N_984);
or U1018 (N_1018,N_973,N_972);
nor U1019 (N_1019,N_967,N_990);
or U1020 (N_1020,N_977,N_992);
nand U1021 (N_1021,N_996,N_971);
or U1022 (N_1022,N_962,N_960);
nand U1023 (N_1023,N_965,N_950);
and U1024 (N_1024,N_957,N_981);
nand U1025 (N_1025,N_970,N_966);
nand U1026 (N_1026,N_951,N_963);
nand U1027 (N_1027,N_951,N_991);
or U1028 (N_1028,N_962,N_951);
nor U1029 (N_1029,N_953,N_990);
or U1030 (N_1030,N_962,N_988);
or U1031 (N_1031,N_983,N_993);
nand U1032 (N_1032,N_967,N_994);
and U1033 (N_1033,N_985,N_979);
or U1034 (N_1034,N_961,N_983);
nand U1035 (N_1035,N_971,N_970);
nand U1036 (N_1036,N_956,N_986);
xor U1037 (N_1037,N_970,N_951);
and U1038 (N_1038,N_996,N_982);
nand U1039 (N_1039,N_971,N_957);
nand U1040 (N_1040,N_963,N_996);
and U1041 (N_1041,N_968,N_957);
and U1042 (N_1042,N_982,N_990);
nor U1043 (N_1043,N_995,N_973);
and U1044 (N_1044,N_975,N_991);
and U1045 (N_1045,N_975,N_954);
and U1046 (N_1046,N_972,N_962);
nor U1047 (N_1047,N_959,N_989);
and U1048 (N_1048,N_979,N_983);
or U1049 (N_1049,N_998,N_951);
nor U1050 (N_1050,N_1014,N_1023);
or U1051 (N_1051,N_1018,N_1003);
or U1052 (N_1052,N_1039,N_1015);
nor U1053 (N_1053,N_1016,N_1032);
nand U1054 (N_1054,N_1021,N_1045);
nand U1055 (N_1055,N_1047,N_1026);
nand U1056 (N_1056,N_1017,N_1011);
and U1057 (N_1057,N_1001,N_1013);
nor U1058 (N_1058,N_1035,N_1005);
nor U1059 (N_1059,N_1025,N_1031);
or U1060 (N_1060,N_1041,N_1004);
or U1061 (N_1061,N_1002,N_1007);
nor U1062 (N_1062,N_1006,N_1012);
or U1063 (N_1063,N_1029,N_1019);
or U1064 (N_1064,N_1022,N_1000);
nor U1065 (N_1065,N_1009,N_1049);
xnor U1066 (N_1066,N_1010,N_1027);
or U1067 (N_1067,N_1020,N_1008);
nand U1068 (N_1068,N_1048,N_1038);
nor U1069 (N_1069,N_1046,N_1024);
nand U1070 (N_1070,N_1030,N_1044);
or U1071 (N_1071,N_1033,N_1042);
or U1072 (N_1072,N_1034,N_1037);
nand U1073 (N_1073,N_1036,N_1040);
and U1074 (N_1074,N_1028,N_1043);
or U1075 (N_1075,N_1018,N_1020);
and U1076 (N_1076,N_1006,N_1010);
nor U1077 (N_1077,N_1023,N_1046);
nand U1078 (N_1078,N_1029,N_1043);
or U1079 (N_1079,N_1024,N_1023);
nand U1080 (N_1080,N_1043,N_1018);
or U1081 (N_1081,N_1000,N_1008);
or U1082 (N_1082,N_1021,N_1042);
nand U1083 (N_1083,N_1027,N_1046);
and U1084 (N_1084,N_1037,N_1001);
nand U1085 (N_1085,N_1039,N_1047);
and U1086 (N_1086,N_1024,N_1011);
and U1087 (N_1087,N_1031,N_1006);
or U1088 (N_1088,N_1034,N_1002);
nor U1089 (N_1089,N_1017,N_1025);
nor U1090 (N_1090,N_1000,N_1028);
nor U1091 (N_1091,N_1011,N_1001);
or U1092 (N_1092,N_1039,N_1004);
nor U1093 (N_1093,N_1048,N_1040);
nand U1094 (N_1094,N_1017,N_1000);
or U1095 (N_1095,N_1013,N_1035);
nand U1096 (N_1096,N_1038,N_1011);
xor U1097 (N_1097,N_1006,N_1008);
or U1098 (N_1098,N_1010,N_1022);
and U1099 (N_1099,N_1041,N_1033);
nor U1100 (N_1100,N_1076,N_1066);
nor U1101 (N_1101,N_1078,N_1063);
nand U1102 (N_1102,N_1064,N_1068);
nand U1103 (N_1103,N_1051,N_1094);
and U1104 (N_1104,N_1072,N_1080);
or U1105 (N_1105,N_1081,N_1054);
and U1106 (N_1106,N_1079,N_1062);
nor U1107 (N_1107,N_1086,N_1089);
nor U1108 (N_1108,N_1070,N_1074);
nand U1109 (N_1109,N_1073,N_1067);
and U1110 (N_1110,N_1060,N_1093);
and U1111 (N_1111,N_1095,N_1096);
nor U1112 (N_1112,N_1050,N_1056);
or U1113 (N_1113,N_1052,N_1061);
and U1114 (N_1114,N_1085,N_1059);
and U1115 (N_1115,N_1053,N_1084);
nor U1116 (N_1116,N_1098,N_1092);
nor U1117 (N_1117,N_1069,N_1055);
and U1118 (N_1118,N_1087,N_1057);
nor U1119 (N_1119,N_1071,N_1088);
nand U1120 (N_1120,N_1065,N_1083);
nor U1121 (N_1121,N_1097,N_1099);
nor U1122 (N_1122,N_1075,N_1058);
nor U1123 (N_1123,N_1091,N_1082);
nor U1124 (N_1124,N_1090,N_1077);
and U1125 (N_1125,N_1070,N_1088);
nand U1126 (N_1126,N_1091,N_1057);
and U1127 (N_1127,N_1053,N_1057);
or U1128 (N_1128,N_1067,N_1090);
or U1129 (N_1129,N_1070,N_1085);
nor U1130 (N_1130,N_1086,N_1081);
and U1131 (N_1131,N_1074,N_1054);
or U1132 (N_1132,N_1050,N_1057);
and U1133 (N_1133,N_1080,N_1062);
nor U1134 (N_1134,N_1081,N_1059);
nor U1135 (N_1135,N_1068,N_1074);
nand U1136 (N_1136,N_1060,N_1083);
and U1137 (N_1137,N_1094,N_1072);
nand U1138 (N_1138,N_1097,N_1071);
or U1139 (N_1139,N_1066,N_1094);
nand U1140 (N_1140,N_1095,N_1093);
nand U1141 (N_1141,N_1058,N_1093);
nand U1142 (N_1142,N_1059,N_1073);
xnor U1143 (N_1143,N_1075,N_1073);
nand U1144 (N_1144,N_1067,N_1056);
nand U1145 (N_1145,N_1084,N_1070);
or U1146 (N_1146,N_1081,N_1099);
nand U1147 (N_1147,N_1084,N_1079);
or U1148 (N_1148,N_1071,N_1057);
or U1149 (N_1149,N_1097,N_1095);
nor U1150 (N_1150,N_1120,N_1129);
nand U1151 (N_1151,N_1136,N_1139);
and U1152 (N_1152,N_1135,N_1107);
or U1153 (N_1153,N_1102,N_1126);
nor U1154 (N_1154,N_1116,N_1140);
xnor U1155 (N_1155,N_1124,N_1146);
nor U1156 (N_1156,N_1143,N_1137);
nor U1157 (N_1157,N_1145,N_1108);
or U1158 (N_1158,N_1127,N_1114);
and U1159 (N_1159,N_1117,N_1133);
nand U1160 (N_1160,N_1112,N_1134);
nand U1161 (N_1161,N_1115,N_1128);
nor U1162 (N_1162,N_1119,N_1105);
and U1163 (N_1163,N_1141,N_1149);
xor U1164 (N_1164,N_1147,N_1110);
nor U1165 (N_1165,N_1106,N_1142);
or U1166 (N_1166,N_1103,N_1113);
nor U1167 (N_1167,N_1123,N_1100);
and U1168 (N_1168,N_1109,N_1132);
nand U1169 (N_1169,N_1148,N_1118);
and U1170 (N_1170,N_1121,N_1104);
and U1171 (N_1171,N_1144,N_1131);
or U1172 (N_1172,N_1125,N_1138);
and U1173 (N_1173,N_1122,N_1101);
nor U1174 (N_1174,N_1130,N_1111);
or U1175 (N_1175,N_1103,N_1143);
and U1176 (N_1176,N_1140,N_1117);
and U1177 (N_1177,N_1119,N_1130);
nor U1178 (N_1178,N_1110,N_1107);
and U1179 (N_1179,N_1142,N_1129);
or U1180 (N_1180,N_1119,N_1135);
nand U1181 (N_1181,N_1140,N_1119);
nor U1182 (N_1182,N_1148,N_1107);
nand U1183 (N_1183,N_1107,N_1132);
nor U1184 (N_1184,N_1100,N_1116);
nand U1185 (N_1185,N_1145,N_1148);
or U1186 (N_1186,N_1143,N_1122);
and U1187 (N_1187,N_1115,N_1114);
and U1188 (N_1188,N_1144,N_1123);
nand U1189 (N_1189,N_1111,N_1119);
and U1190 (N_1190,N_1145,N_1140);
and U1191 (N_1191,N_1138,N_1126);
nand U1192 (N_1192,N_1133,N_1118);
nand U1193 (N_1193,N_1148,N_1121);
nor U1194 (N_1194,N_1104,N_1147);
nor U1195 (N_1195,N_1130,N_1137);
nand U1196 (N_1196,N_1119,N_1120);
or U1197 (N_1197,N_1107,N_1121);
nand U1198 (N_1198,N_1149,N_1117);
nor U1199 (N_1199,N_1114,N_1129);
or U1200 (N_1200,N_1156,N_1175);
or U1201 (N_1201,N_1172,N_1177);
and U1202 (N_1202,N_1162,N_1192);
and U1203 (N_1203,N_1181,N_1179);
nor U1204 (N_1204,N_1168,N_1176);
nor U1205 (N_1205,N_1173,N_1197);
nor U1206 (N_1206,N_1193,N_1157);
nor U1207 (N_1207,N_1169,N_1190);
or U1208 (N_1208,N_1170,N_1152);
or U1209 (N_1209,N_1194,N_1182);
and U1210 (N_1210,N_1151,N_1167);
and U1211 (N_1211,N_1186,N_1161);
and U1212 (N_1212,N_1158,N_1153);
nand U1213 (N_1213,N_1163,N_1171);
or U1214 (N_1214,N_1180,N_1166);
nor U1215 (N_1215,N_1189,N_1155);
or U1216 (N_1216,N_1183,N_1178);
nand U1217 (N_1217,N_1187,N_1184);
nor U1218 (N_1218,N_1160,N_1185);
nor U1219 (N_1219,N_1191,N_1165);
or U1220 (N_1220,N_1174,N_1188);
or U1221 (N_1221,N_1159,N_1198);
nor U1222 (N_1222,N_1195,N_1196);
or U1223 (N_1223,N_1150,N_1154);
and U1224 (N_1224,N_1199,N_1164);
and U1225 (N_1225,N_1150,N_1178);
nor U1226 (N_1226,N_1197,N_1193);
and U1227 (N_1227,N_1167,N_1181);
or U1228 (N_1228,N_1166,N_1199);
or U1229 (N_1229,N_1174,N_1180);
or U1230 (N_1230,N_1157,N_1185);
nor U1231 (N_1231,N_1187,N_1182);
nand U1232 (N_1232,N_1184,N_1197);
or U1233 (N_1233,N_1160,N_1163);
nor U1234 (N_1234,N_1174,N_1197);
nor U1235 (N_1235,N_1162,N_1191);
nor U1236 (N_1236,N_1180,N_1172);
nor U1237 (N_1237,N_1152,N_1164);
nor U1238 (N_1238,N_1170,N_1198);
or U1239 (N_1239,N_1196,N_1162);
and U1240 (N_1240,N_1187,N_1161);
nor U1241 (N_1241,N_1182,N_1163);
and U1242 (N_1242,N_1173,N_1166);
nor U1243 (N_1243,N_1151,N_1154);
nor U1244 (N_1244,N_1193,N_1194);
nand U1245 (N_1245,N_1162,N_1185);
nor U1246 (N_1246,N_1165,N_1193);
nor U1247 (N_1247,N_1185,N_1167);
nor U1248 (N_1248,N_1170,N_1196);
nand U1249 (N_1249,N_1163,N_1178);
nor U1250 (N_1250,N_1232,N_1214);
nor U1251 (N_1251,N_1249,N_1220);
and U1252 (N_1252,N_1236,N_1241);
or U1253 (N_1253,N_1217,N_1226);
or U1254 (N_1254,N_1225,N_1234);
xnor U1255 (N_1255,N_1243,N_1208);
nand U1256 (N_1256,N_1201,N_1248);
nand U1257 (N_1257,N_1230,N_1218);
nor U1258 (N_1258,N_1202,N_1209);
nor U1259 (N_1259,N_1216,N_1221);
and U1260 (N_1260,N_1237,N_1205);
nand U1261 (N_1261,N_1204,N_1244);
or U1262 (N_1262,N_1242,N_1246);
nand U1263 (N_1263,N_1233,N_1239);
nor U1264 (N_1264,N_1247,N_1207);
nand U1265 (N_1265,N_1222,N_1228);
nand U1266 (N_1266,N_1240,N_1200);
nand U1267 (N_1267,N_1229,N_1215);
nor U1268 (N_1268,N_1238,N_1206);
and U1269 (N_1269,N_1211,N_1235);
nor U1270 (N_1270,N_1219,N_1203);
and U1271 (N_1271,N_1210,N_1223);
nand U1272 (N_1272,N_1224,N_1231);
or U1273 (N_1273,N_1212,N_1227);
nor U1274 (N_1274,N_1213,N_1245);
nand U1275 (N_1275,N_1202,N_1222);
nand U1276 (N_1276,N_1236,N_1209);
nor U1277 (N_1277,N_1227,N_1209);
nor U1278 (N_1278,N_1241,N_1209);
nand U1279 (N_1279,N_1230,N_1217);
or U1280 (N_1280,N_1232,N_1241);
and U1281 (N_1281,N_1202,N_1233);
and U1282 (N_1282,N_1203,N_1237);
or U1283 (N_1283,N_1245,N_1212);
and U1284 (N_1284,N_1217,N_1228);
nor U1285 (N_1285,N_1204,N_1236);
nand U1286 (N_1286,N_1200,N_1207);
nand U1287 (N_1287,N_1242,N_1235);
nor U1288 (N_1288,N_1226,N_1208);
nor U1289 (N_1289,N_1246,N_1214);
and U1290 (N_1290,N_1249,N_1202);
nand U1291 (N_1291,N_1222,N_1212);
nor U1292 (N_1292,N_1204,N_1215);
nand U1293 (N_1293,N_1225,N_1249);
nand U1294 (N_1294,N_1206,N_1243);
and U1295 (N_1295,N_1225,N_1214);
and U1296 (N_1296,N_1245,N_1241);
nand U1297 (N_1297,N_1240,N_1205);
nand U1298 (N_1298,N_1219,N_1234);
nor U1299 (N_1299,N_1244,N_1245);
nor U1300 (N_1300,N_1284,N_1280);
or U1301 (N_1301,N_1267,N_1255);
nor U1302 (N_1302,N_1291,N_1260);
nor U1303 (N_1303,N_1292,N_1286);
nand U1304 (N_1304,N_1256,N_1254);
and U1305 (N_1305,N_1266,N_1288);
or U1306 (N_1306,N_1290,N_1298);
nor U1307 (N_1307,N_1274,N_1257);
and U1308 (N_1308,N_1297,N_1294);
and U1309 (N_1309,N_1250,N_1278);
nand U1310 (N_1310,N_1275,N_1276);
or U1311 (N_1311,N_1262,N_1296);
and U1312 (N_1312,N_1252,N_1273);
nor U1313 (N_1313,N_1265,N_1271);
or U1314 (N_1314,N_1261,N_1289);
and U1315 (N_1315,N_1287,N_1285);
or U1316 (N_1316,N_1295,N_1293);
nor U1317 (N_1317,N_1269,N_1279);
and U1318 (N_1318,N_1283,N_1270);
or U1319 (N_1319,N_1264,N_1258);
nand U1320 (N_1320,N_1281,N_1259);
nor U1321 (N_1321,N_1277,N_1268);
nand U1322 (N_1322,N_1299,N_1251);
nor U1323 (N_1323,N_1263,N_1282);
and U1324 (N_1324,N_1272,N_1253);
or U1325 (N_1325,N_1294,N_1295);
nor U1326 (N_1326,N_1263,N_1251);
and U1327 (N_1327,N_1287,N_1260);
and U1328 (N_1328,N_1259,N_1286);
nand U1329 (N_1329,N_1299,N_1276);
or U1330 (N_1330,N_1266,N_1267);
nor U1331 (N_1331,N_1286,N_1277);
nor U1332 (N_1332,N_1280,N_1270);
nand U1333 (N_1333,N_1258,N_1267);
nand U1334 (N_1334,N_1281,N_1269);
or U1335 (N_1335,N_1292,N_1285);
nor U1336 (N_1336,N_1265,N_1293);
nor U1337 (N_1337,N_1255,N_1260);
nand U1338 (N_1338,N_1259,N_1270);
nand U1339 (N_1339,N_1278,N_1270);
xor U1340 (N_1340,N_1274,N_1275);
and U1341 (N_1341,N_1279,N_1264);
and U1342 (N_1342,N_1286,N_1271);
and U1343 (N_1343,N_1283,N_1251);
and U1344 (N_1344,N_1284,N_1273);
and U1345 (N_1345,N_1266,N_1285);
nor U1346 (N_1346,N_1259,N_1271);
and U1347 (N_1347,N_1273,N_1293);
or U1348 (N_1348,N_1288,N_1285);
nor U1349 (N_1349,N_1254,N_1261);
or U1350 (N_1350,N_1306,N_1343);
or U1351 (N_1351,N_1320,N_1310);
nor U1352 (N_1352,N_1312,N_1308);
and U1353 (N_1353,N_1327,N_1326);
nor U1354 (N_1354,N_1341,N_1347);
nor U1355 (N_1355,N_1346,N_1304);
nor U1356 (N_1356,N_1335,N_1349);
nand U1357 (N_1357,N_1334,N_1332);
nand U1358 (N_1358,N_1345,N_1333);
and U1359 (N_1359,N_1322,N_1329);
or U1360 (N_1360,N_1314,N_1302);
nand U1361 (N_1361,N_1321,N_1309);
and U1362 (N_1362,N_1315,N_1316);
and U1363 (N_1363,N_1348,N_1313);
nor U1364 (N_1364,N_1301,N_1319);
or U1365 (N_1365,N_1307,N_1339);
nand U1366 (N_1366,N_1323,N_1325);
and U1367 (N_1367,N_1340,N_1328);
and U1368 (N_1368,N_1342,N_1324);
and U1369 (N_1369,N_1311,N_1305);
nor U1370 (N_1370,N_1300,N_1330);
nor U1371 (N_1371,N_1344,N_1318);
and U1372 (N_1372,N_1337,N_1338);
and U1373 (N_1373,N_1303,N_1317);
nor U1374 (N_1374,N_1331,N_1336);
or U1375 (N_1375,N_1327,N_1310);
nor U1376 (N_1376,N_1309,N_1324);
nand U1377 (N_1377,N_1307,N_1328);
or U1378 (N_1378,N_1322,N_1333);
nor U1379 (N_1379,N_1316,N_1318);
nand U1380 (N_1380,N_1315,N_1322);
xnor U1381 (N_1381,N_1330,N_1346);
nand U1382 (N_1382,N_1325,N_1302);
or U1383 (N_1383,N_1334,N_1345);
and U1384 (N_1384,N_1300,N_1307);
and U1385 (N_1385,N_1325,N_1343);
or U1386 (N_1386,N_1312,N_1320);
and U1387 (N_1387,N_1305,N_1348);
nand U1388 (N_1388,N_1319,N_1331);
and U1389 (N_1389,N_1311,N_1338);
and U1390 (N_1390,N_1324,N_1341);
and U1391 (N_1391,N_1303,N_1342);
and U1392 (N_1392,N_1317,N_1343);
and U1393 (N_1393,N_1318,N_1329);
and U1394 (N_1394,N_1314,N_1301);
or U1395 (N_1395,N_1344,N_1307);
nor U1396 (N_1396,N_1346,N_1344);
or U1397 (N_1397,N_1312,N_1316);
and U1398 (N_1398,N_1309,N_1300);
or U1399 (N_1399,N_1311,N_1332);
nor U1400 (N_1400,N_1392,N_1356);
nand U1401 (N_1401,N_1354,N_1367);
and U1402 (N_1402,N_1359,N_1387);
nand U1403 (N_1403,N_1375,N_1370);
and U1404 (N_1404,N_1378,N_1353);
or U1405 (N_1405,N_1357,N_1364);
or U1406 (N_1406,N_1363,N_1377);
and U1407 (N_1407,N_1373,N_1351);
and U1408 (N_1408,N_1372,N_1384);
and U1409 (N_1409,N_1362,N_1360);
and U1410 (N_1410,N_1396,N_1380);
and U1411 (N_1411,N_1352,N_1365);
nand U1412 (N_1412,N_1383,N_1385);
or U1413 (N_1413,N_1394,N_1388);
nand U1414 (N_1414,N_1399,N_1393);
nand U1415 (N_1415,N_1376,N_1369);
nand U1416 (N_1416,N_1386,N_1379);
and U1417 (N_1417,N_1381,N_1368);
nor U1418 (N_1418,N_1398,N_1366);
nand U1419 (N_1419,N_1350,N_1395);
nor U1420 (N_1420,N_1371,N_1389);
and U1421 (N_1421,N_1397,N_1358);
or U1422 (N_1422,N_1390,N_1355);
or U1423 (N_1423,N_1374,N_1361);
or U1424 (N_1424,N_1382,N_1391);
and U1425 (N_1425,N_1395,N_1351);
nor U1426 (N_1426,N_1355,N_1363);
xnor U1427 (N_1427,N_1386,N_1371);
and U1428 (N_1428,N_1389,N_1378);
nor U1429 (N_1429,N_1390,N_1367);
or U1430 (N_1430,N_1361,N_1364);
nand U1431 (N_1431,N_1366,N_1392);
and U1432 (N_1432,N_1354,N_1392);
and U1433 (N_1433,N_1399,N_1394);
nand U1434 (N_1434,N_1391,N_1355);
and U1435 (N_1435,N_1351,N_1360);
xor U1436 (N_1436,N_1385,N_1395);
nor U1437 (N_1437,N_1377,N_1365);
and U1438 (N_1438,N_1372,N_1381);
and U1439 (N_1439,N_1355,N_1362);
nand U1440 (N_1440,N_1393,N_1377);
nand U1441 (N_1441,N_1377,N_1354);
and U1442 (N_1442,N_1382,N_1376);
or U1443 (N_1443,N_1360,N_1380);
and U1444 (N_1444,N_1351,N_1365);
nand U1445 (N_1445,N_1393,N_1359);
or U1446 (N_1446,N_1388,N_1356);
nand U1447 (N_1447,N_1395,N_1363);
nand U1448 (N_1448,N_1398,N_1377);
or U1449 (N_1449,N_1381,N_1376);
nand U1450 (N_1450,N_1432,N_1418);
or U1451 (N_1451,N_1410,N_1440);
and U1452 (N_1452,N_1419,N_1426);
nor U1453 (N_1453,N_1406,N_1436);
or U1454 (N_1454,N_1429,N_1422);
and U1455 (N_1455,N_1431,N_1448);
nor U1456 (N_1456,N_1449,N_1408);
nor U1457 (N_1457,N_1400,N_1407);
or U1458 (N_1458,N_1433,N_1439);
nand U1459 (N_1459,N_1415,N_1430);
or U1460 (N_1460,N_1401,N_1425);
and U1461 (N_1461,N_1434,N_1403);
and U1462 (N_1462,N_1435,N_1446);
nand U1463 (N_1463,N_1414,N_1412);
or U1464 (N_1464,N_1444,N_1438);
and U1465 (N_1465,N_1445,N_1409);
and U1466 (N_1466,N_1413,N_1443);
and U1467 (N_1467,N_1417,N_1404);
or U1468 (N_1468,N_1420,N_1416);
nand U1469 (N_1469,N_1437,N_1424);
and U1470 (N_1470,N_1428,N_1405);
or U1471 (N_1471,N_1421,N_1442);
or U1472 (N_1472,N_1427,N_1423);
nand U1473 (N_1473,N_1411,N_1402);
and U1474 (N_1474,N_1441,N_1447);
or U1475 (N_1475,N_1445,N_1404);
or U1476 (N_1476,N_1405,N_1408);
and U1477 (N_1477,N_1438,N_1417);
or U1478 (N_1478,N_1428,N_1419);
and U1479 (N_1479,N_1421,N_1435);
or U1480 (N_1480,N_1428,N_1414);
nand U1481 (N_1481,N_1413,N_1434);
nand U1482 (N_1482,N_1443,N_1419);
or U1483 (N_1483,N_1431,N_1422);
xnor U1484 (N_1484,N_1410,N_1435);
nor U1485 (N_1485,N_1413,N_1404);
and U1486 (N_1486,N_1404,N_1447);
and U1487 (N_1487,N_1409,N_1447);
nor U1488 (N_1488,N_1431,N_1403);
or U1489 (N_1489,N_1420,N_1436);
xnor U1490 (N_1490,N_1406,N_1402);
and U1491 (N_1491,N_1415,N_1408);
or U1492 (N_1492,N_1426,N_1418);
nand U1493 (N_1493,N_1421,N_1433);
or U1494 (N_1494,N_1403,N_1404);
nor U1495 (N_1495,N_1431,N_1449);
or U1496 (N_1496,N_1423,N_1401);
or U1497 (N_1497,N_1412,N_1434);
or U1498 (N_1498,N_1418,N_1431);
or U1499 (N_1499,N_1442,N_1425);
nand U1500 (N_1500,N_1461,N_1490);
nand U1501 (N_1501,N_1488,N_1483);
nor U1502 (N_1502,N_1498,N_1452);
xor U1503 (N_1503,N_1451,N_1475);
xnor U1504 (N_1504,N_1470,N_1471);
or U1505 (N_1505,N_1469,N_1493);
or U1506 (N_1506,N_1497,N_1485);
or U1507 (N_1507,N_1479,N_1478);
or U1508 (N_1508,N_1458,N_1460);
and U1509 (N_1509,N_1480,N_1468);
nand U1510 (N_1510,N_1477,N_1484);
nor U1511 (N_1511,N_1492,N_1466);
xor U1512 (N_1512,N_1462,N_1472);
nand U1513 (N_1513,N_1474,N_1489);
xor U1514 (N_1514,N_1456,N_1491);
and U1515 (N_1515,N_1496,N_1482);
or U1516 (N_1516,N_1450,N_1473);
or U1517 (N_1517,N_1453,N_1486);
nand U1518 (N_1518,N_1464,N_1465);
nor U1519 (N_1519,N_1459,N_1481);
nor U1520 (N_1520,N_1455,N_1499);
nand U1521 (N_1521,N_1494,N_1467);
nor U1522 (N_1522,N_1457,N_1454);
or U1523 (N_1523,N_1463,N_1487);
or U1524 (N_1524,N_1495,N_1476);
and U1525 (N_1525,N_1456,N_1480);
nor U1526 (N_1526,N_1452,N_1490);
nand U1527 (N_1527,N_1463,N_1452);
or U1528 (N_1528,N_1486,N_1462);
nand U1529 (N_1529,N_1465,N_1457);
and U1530 (N_1530,N_1466,N_1452);
nor U1531 (N_1531,N_1487,N_1486);
nand U1532 (N_1532,N_1488,N_1494);
or U1533 (N_1533,N_1473,N_1474);
nor U1534 (N_1534,N_1459,N_1484);
nor U1535 (N_1535,N_1461,N_1496);
or U1536 (N_1536,N_1492,N_1477);
nand U1537 (N_1537,N_1493,N_1465);
nand U1538 (N_1538,N_1480,N_1454);
and U1539 (N_1539,N_1484,N_1478);
xnor U1540 (N_1540,N_1492,N_1484);
xor U1541 (N_1541,N_1498,N_1458);
nand U1542 (N_1542,N_1476,N_1483);
nand U1543 (N_1543,N_1495,N_1471);
nor U1544 (N_1544,N_1458,N_1474);
and U1545 (N_1545,N_1490,N_1487);
and U1546 (N_1546,N_1483,N_1497);
nand U1547 (N_1547,N_1450,N_1468);
nor U1548 (N_1548,N_1494,N_1477);
or U1549 (N_1549,N_1489,N_1456);
nor U1550 (N_1550,N_1523,N_1527);
and U1551 (N_1551,N_1533,N_1547);
and U1552 (N_1552,N_1512,N_1525);
or U1553 (N_1553,N_1504,N_1517);
and U1554 (N_1554,N_1548,N_1537);
nand U1555 (N_1555,N_1506,N_1549);
nor U1556 (N_1556,N_1515,N_1510);
or U1557 (N_1557,N_1540,N_1521);
and U1558 (N_1558,N_1529,N_1502);
or U1559 (N_1559,N_1543,N_1524);
nor U1560 (N_1560,N_1544,N_1531);
nand U1561 (N_1561,N_1514,N_1503);
or U1562 (N_1562,N_1532,N_1518);
and U1563 (N_1563,N_1542,N_1508);
nor U1564 (N_1564,N_1522,N_1545);
and U1565 (N_1565,N_1526,N_1535);
nand U1566 (N_1566,N_1507,N_1530);
and U1567 (N_1567,N_1509,N_1539);
nor U1568 (N_1568,N_1541,N_1536);
or U1569 (N_1569,N_1546,N_1501);
nor U1570 (N_1570,N_1519,N_1528);
and U1571 (N_1571,N_1513,N_1500);
or U1572 (N_1572,N_1505,N_1534);
nor U1573 (N_1573,N_1538,N_1511);
and U1574 (N_1574,N_1516,N_1520);
and U1575 (N_1575,N_1526,N_1533);
or U1576 (N_1576,N_1510,N_1505);
nand U1577 (N_1577,N_1513,N_1518);
nor U1578 (N_1578,N_1527,N_1542);
nor U1579 (N_1579,N_1533,N_1535);
nor U1580 (N_1580,N_1531,N_1515);
nor U1581 (N_1581,N_1509,N_1505);
or U1582 (N_1582,N_1500,N_1503);
and U1583 (N_1583,N_1514,N_1510);
nor U1584 (N_1584,N_1500,N_1534);
and U1585 (N_1585,N_1524,N_1531);
nor U1586 (N_1586,N_1517,N_1529);
and U1587 (N_1587,N_1508,N_1548);
or U1588 (N_1588,N_1546,N_1535);
nor U1589 (N_1589,N_1543,N_1519);
or U1590 (N_1590,N_1513,N_1530);
nor U1591 (N_1591,N_1520,N_1511);
and U1592 (N_1592,N_1503,N_1509);
nor U1593 (N_1593,N_1510,N_1524);
or U1594 (N_1594,N_1534,N_1516);
nor U1595 (N_1595,N_1542,N_1540);
nor U1596 (N_1596,N_1524,N_1505);
or U1597 (N_1597,N_1534,N_1543);
nand U1598 (N_1598,N_1547,N_1517);
nor U1599 (N_1599,N_1524,N_1528);
or U1600 (N_1600,N_1550,N_1560);
nand U1601 (N_1601,N_1574,N_1595);
or U1602 (N_1602,N_1596,N_1584);
nand U1603 (N_1603,N_1567,N_1580);
nor U1604 (N_1604,N_1587,N_1581);
nor U1605 (N_1605,N_1568,N_1558);
nor U1606 (N_1606,N_1578,N_1570);
nor U1607 (N_1607,N_1591,N_1556);
and U1608 (N_1608,N_1593,N_1564);
and U1609 (N_1609,N_1562,N_1594);
nand U1610 (N_1610,N_1577,N_1590);
or U1611 (N_1611,N_1575,N_1585);
and U1612 (N_1612,N_1557,N_1552);
or U1613 (N_1613,N_1589,N_1583);
or U1614 (N_1614,N_1598,N_1579);
nand U1615 (N_1615,N_1572,N_1592);
nor U1616 (N_1616,N_1599,N_1563);
and U1617 (N_1617,N_1566,N_1597);
or U1618 (N_1618,N_1554,N_1559);
or U1619 (N_1619,N_1571,N_1569);
and U1620 (N_1620,N_1586,N_1565);
nor U1621 (N_1621,N_1551,N_1561);
and U1622 (N_1622,N_1576,N_1588);
and U1623 (N_1623,N_1553,N_1582);
nand U1624 (N_1624,N_1555,N_1573);
nor U1625 (N_1625,N_1598,N_1577);
or U1626 (N_1626,N_1583,N_1571);
and U1627 (N_1627,N_1598,N_1572);
and U1628 (N_1628,N_1555,N_1553);
nand U1629 (N_1629,N_1551,N_1588);
nand U1630 (N_1630,N_1551,N_1575);
nor U1631 (N_1631,N_1586,N_1556);
nor U1632 (N_1632,N_1554,N_1593);
nand U1633 (N_1633,N_1564,N_1594);
and U1634 (N_1634,N_1577,N_1581);
nand U1635 (N_1635,N_1579,N_1564);
nor U1636 (N_1636,N_1596,N_1575);
and U1637 (N_1637,N_1590,N_1586);
or U1638 (N_1638,N_1550,N_1580);
and U1639 (N_1639,N_1558,N_1590);
nor U1640 (N_1640,N_1554,N_1565);
or U1641 (N_1641,N_1590,N_1559);
nor U1642 (N_1642,N_1561,N_1552);
nand U1643 (N_1643,N_1597,N_1556);
nor U1644 (N_1644,N_1567,N_1586);
and U1645 (N_1645,N_1590,N_1572);
nand U1646 (N_1646,N_1555,N_1566);
nand U1647 (N_1647,N_1594,N_1590);
nor U1648 (N_1648,N_1573,N_1583);
nor U1649 (N_1649,N_1571,N_1588);
or U1650 (N_1650,N_1600,N_1628);
nand U1651 (N_1651,N_1640,N_1619);
nand U1652 (N_1652,N_1609,N_1607);
nor U1653 (N_1653,N_1627,N_1623);
nor U1654 (N_1654,N_1624,N_1626);
nor U1655 (N_1655,N_1641,N_1620);
and U1656 (N_1656,N_1639,N_1621);
nand U1657 (N_1657,N_1616,N_1604);
or U1658 (N_1658,N_1631,N_1642);
nand U1659 (N_1659,N_1649,N_1644);
nand U1660 (N_1660,N_1610,N_1615);
and U1661 (N_1661,N_1637,N_1630);
or U1662 (N_1662,N_1635,N_1645);
nor U1663 (N_1663,N_1638,N_1617);
and U1664 (N_1664,N_1629,N_1612);
nand U1665 (N_1665,N_1602,N_1603);
and U1666 (N_1666,N_1622,N_1606);
nand U1667 (N_1667,N_1643,N_1611);
xor U1668 (N_1668,N_1614,N_1618);
nor U1669 (N_1669,N_1647,N_1648);
or U1670 (N_1670,N_1633,N_1601);
and U1671 (N_1671,N_1605,N_1608);
nand U1672 (N_1672,N_1632,N_1634);
nand U1673 (N_1673,N_1625,N_1646);
nor U1674 (N_1674,N_1613,N_1636);
or U1675 (N_1675,N_1635,N_1606);
and U1676 (N_1676,N_1623,N_1613);
and U1677 (N_1677,N_1638,N_1602);
nor U1678 (N_1678,N_1625,N_1627);
or U1679 (N_1679,N_1644,N_1635);
and U1680 (N_1680,N_1600,N_1609);
or U1681 (N_1681,N_1623,N_1600);
nor U1682 (N_1682,N_1613,N_1619);
or U1683 (N_1683,N_1626,N_1603);
nand U1684 (N_1684,N_1615,N_1617);
nor U1685 (N_1685,N_1608,N_1619);
nand U1686 (N_1686,N_1637,N_1624);
and U1687 (N_1687,N_1627,N_1626);
nand U1688 (N_1688,N_1624,N_1629);
xor U1689 (N_1689,N_1643,N_1640);
or U1690 (N_1690,N_1623,N_1630);
nand U1691 (N_1691,N_1649,N_1614);
xnor U1692 (N_1692,N_1619,N_1609);
nand U1693 (N_1693,N_1628,N_1630);
nand U1694 (N_1694,N_1642,N_1608);
and U1695 (N_1695,N_1608,N_1644);
nor U1696 (N_1696,N_1616,N_1645);
or U1697 (N_1697,N_1624,N_1609);
or U1698 (N_1698,N_1608,N_1641);
and U1699 (N_1699,N_1629,N_1636);
and U1700 (N_1700,N_1661,N_1671);
or U1701 (N_1701,N_1675,N_1662);
and U1702 (N_1702,N_1658,N_1655);
nand U1703 (N_1703,N_1670,N_1663);
or U1704 (N_1704,N_1668,N_1698);
nand U1705 (N_1705,N_1657,N_1677);
and U1706 (N_1706,N_1680,N_1660);
nand U1707 (N_1707,N_1652,N_1683);
and U1708 (N_1708,N_1689,N_1696);
nor U1709 (N_1709,N_1673,N_1651);
nor U1710 (N_1710,N_1682,N_1676);
and U1711 (N_1711,N_1697,N_1659);
or U1712 (N_1712,N_1685,N_1665);
nor U1713 (N_1713,N_1667,N_1681);
nor U1714 (N_1714,N_1656,N_1666);
and U1715 (N_1715,N_1695,N_1674);
and U1716 (N_1716,N_1686,N_1669);
or U1717 (N_1717,N_1678,N_1687);
nand U1718 (N_1718,N_1694,N_1699);
and U1719 (N_1719,N_1650,N_1691);
xnor U1720 (N_1720,N_1664,N_1654);
or U1721 (N_1721,N_1690,N_1693);
nor U1722 (N_1722,N_1688,N_1679);
nor U1723 (N_1723,N_1653,N_1684);
nand U1724 (N_1724,N_1672,N_1692);
nand U1725 (N_1725,N_1671,N_1667);
nand U1726 (N_1726,N_1670,N_1675);
nor U1727 (N_1727,N_1671,N_1675);
nor U1728 (N_1728,N_1661,N_1684);
nand U1729 (N_1729,N_1659,N_1664);
nand U1730 (N_1730,N_1699,N_1686);
nand U1731 (N_1731,N_1654,N_1697);
nand U1732 (N_1732,N_1698,N_1681);
nand U1733 (N_1733,N_1681,N_1653);
nand U1734 (N_1734,N_1673,N_1686);
nor U1735 (N_1735,N_1699,N_1655);
and U1736 (N_1736,N_1688,N_1655);
or U1737 (N_1737,N_1699,N_1657);
and U1738 (N_1738,N_1661,N_1662);
or U1739 (N_1739,N_1667,N_1652);
or U1740 (N_1740,N_1670,N_1659);
nor U1741 (N_1741,N_1657,N_1674);
nand U1742 (N_1742,N_1674,N_1682);
and U1743 (N_1743,N_1655,N_1678);
or U1744 (N_1744,N_1692,N_1694);
and U1745 (N_1745,N_1663,N_1687);
or U1746 (N_1746,N_1689,N_1698);
or U1747 (N_1747,N_1683,N_1672);
or U1748 (N_1748,N_1656,N_1682);
or U1749 (N_1749,N_1655,N_1665);
or U1750 (N_1750,N_1743,N_1717);
or U1751 (N_1751,N_1733,N_1732);
and U1752 (N_1752,N_1701,N_1721);
and U1753 (N_1753,N_1720,N_1738);
nand U1754 (N_1754,N_1702,N_1747);
nand U1755 (N_1755,N_1719,N_1705);
and U1756 (N_1756,N_1749,N_1710);
nor U1757 (N_1757,N_1748,N_1740);
nor U1758 (N_1758,N_1742,N_1722);
nand U1759 (N_1759,N_1744,N_1736);
or U1760 (N_1760,N_1727,N_1704);
or U1761 (N_1761,N_1737,N_1706);
nor U1762 (N_1762,N_1703,N_1746);
nor U1763 (N_1763,N_1739,N_1700);
or U1764 (N_1764,N_1713,N_1735);
nor U1765 (N_1765,N_1707,N_1741);
nor U1766 (N_1766,N_1730,N_1726);
xor U1767 (N_1767,N_1728,N_1745);
or U1768 (N_1768,N_1715,N_1712);
and U1769 (N_1769,N_1731,N_1734);
or U1770 (N_1770,N_1709,N_1725);
nor U1771 (N_1771,N_1729,N_1711);
nand U1772 (N_1772,N_1723,N_1718);
and U1773 (N_1773,N_1708,N_1724);
nor U1774 (N_1774,N_1714,N_1716);
nand U1775 (N_1775,N_1716,N_1733);
or U1776 (N_1776,N_1746,N_1724);
nand U1777 (N_1777,N_1714,N_1735);
nor U1778 (N_1778,N_1708,N_1736);
nor U1779 (N_1779,N_1740,N_1710);
or U1780 (N_1780,N_1720,N_1737);
and U1781 (N_1781,N_1733,N_1747);
and U1782 (N_1782,N_1742,N_1747);
or U1783 (N_1783,N_1715,N_1738);
nand U1784 (N_1784,N_1701,N_1749);
and U1785 (N_1785,N_1708,N_1732);
nor U1786 (N_1786,N_1744,N_1700);
or U1787 (N_1787,N_1717,N_1709);
and U1788 (N_1788,N_1723,N_1714);
and U1789 (N_1789,N_1740,N_1700);
and U1790 (N_1790,N_1709,N_1705);
nand U1791 (N_1791,N_1714,N_1736);
nand U1792 (N_1792,N_1719,N_1738);
nand U1793 (N_1793,N_1747,N_1700);
nand U1794 (N_1794,N_1730,N_1739);
nor U1795 (N_1795,N_1717,N_1701);
nand U1796 (N_1796,N_1740,N_1749);
or U1797 (N_1797,N_1710,N_1719);
nor U1798 (N_1798,N_1707,N_1716);
nor U1799 (N_1799,N_1711,N_1737);
or U1800 (N_1800,N_1769,N_1753);
nor U1801 (N_1801,N_1791,N_1768);
nor U1802 (N_1802,N_1797,N_1779);
nor U1803 (N_1803,N_1774,N_1786);
nor U1804 (N_1804,N_1764,N_1799);
nor U1805 (N_1805,N_1763,N_1790);
nor U1806 (N_1806,N_1782,N_1798);
nand U1807 (N_1807,N_1785,N_1757);
and U1808 (N_1808,N_1788,N_1795);
nand U1809 (N_1809,N_1758,N_1752);
and U1810 (N_1810,N_1793,N_1778);
nand U1811 (N_1811,N_1796,N_1775);
nand U1812 (N_1812,N_1783,N_1780);
or U1813 (N_1813,N_1750,N_1760);
and U1814 (N_1814,N_1759,N_1770);
nand U1815 (N_1815,N_1765,N_1756);
nor U1816 (N_1816,N_1771,N_1772);
or U1817 (N_1817,N_1751,N_1792);
and U1818 (N_1818,N_1781,N_1784);
nor U1819 (N_1819,N_1794,N_1762);
nand U1820 (N_1820,N_1776,N_1767);
and U1821 (N_1821,N_1754,N_1761);
nor U1822 (N_1822,N_1766,N_1755);
and U1823 (N_1823,N_1773,N_1787);
nand U1824 (N_1824,N_1777,N_1789);
nand U1825 (N_1825,N_1750,N_1765);
and U1826 (N_1826,N_1788,N_1751);
nand U1827 (N_1827,N_1769,N_1784);
nand U1828 (N_1828,N_1757,N_1797);
or U1829 (N_1829,N_1764,N_1785);
and U1830 (N_1830,N_1772,N_1780);
and U1831 (N_1831,N_1793,N_1782);
nor U1832 (N_1832,N_1750,N_1779);
or U1833 (N_1833,N_1750,N_1764);
nand U1834 (N_1834,N_1754,N_1772);
and U1835 (N_1835,N_1764,N_1753);
or U1836 (N_1836,N_1764,N_1771);
nand U1837 (N_1837,N_1754,N_1789);
xnor U1838 (N_1838,N_1757,N_1752);
nor U1839 (N_1839,N_1774,N_1799);
or U1840 (N_1840,N_1792,N_1784);
or U1841 (N_1841,N_1796,N_1761);
nor U1842 (N_1842,N_1780,N_1757);
nor U1843 (N_1843,N_1790,N_1754);
nand U1844 (N_1844,N_1784,N_1776);
or U1845 (N_1845,N_1764,N_1780);
or U1846 (N_1846,N_1759,N_1776);
nor U1847 (N_1847,N_1784,N_1783);
nand U1848 (N_1848,N_1769,N_1773);
and U1849 (N_1849,N_1787,N_1768);
xnor U1850 (N_1850,N_1845,N_1829);
nor U1851 (N_1851,N_1837,N_1825);
nor U1852 (N_1852,N_1844,N_1842);
and U1853 (N_1853,N_1834,N_1840);
and U1854 (N_1854,N_1841,N_1801);
and U1855 (N_1855,N_1816,N_1846);
and U1856 (N_1856,N_1843,N_1824);
nor U1857 (N_1857,N_1802,N_1813);
and U1858 (N_1858,N_1822,N_1828);
and U1859 (N_1859,N_1817,N_1810);
nand U1860 (N_1860,N_1839,N_1847);
nand U1861 (N_1861,N_1809,N_1804);
nand U1862 (N_1862,N_1823,N_1827);
or U1863 (N_1863,N_1803,N_1849);
nand U1864 (N_1864,N_1800,N_1814);
and U1865 (N_1865,N_1806,N_1820);
nor U1866 (N_1866,N_1819,N_1831);
nor U1867 (N_1867,N_1835,N_1848);
and U1868 (N_1868,N_1833,N_1807);
nor U1869 (N_1869,N_1821,N_1830);
nand U1870 (N_1870,N_1826,N_1805);
xnor U1871 (N_1871,N_1812,N_1836);
or U1872 (N_1872,N_1832,N_1808);
or U1873 (N_1873,N_1818,N_1811);
nor U1874 (N_1874,N_1815,N_1838);
and U1875 (N_1875,N_1816,N_1848);
or U1876 (N_1876,N_1849,N_1835);
and U1877 (N_1877,N_1841,N_1800);
nand U1878 (N_1878,N_1802,N_1841);
or U1879 (N_1879,N_1836,N_1804);
or U1880 (N_1880,N_1846,N_1830);
or U1881 (N_1881,N_1822,N_1817);
or U1882 (N_1882,N_1812,N_1827);
nand U1883 (N_1883,N_1840,N_1807);
nand U1884 (N_1884,N_1800,N_1822);
nor U1885 (N_1885,N_1825,N_1840);
xor U1886 (N_1886,N_1801,N_1815);
and U1887 (N_1887,N_1815,N_1823);
and U1888 (N_1888,N_1815,N_1817);
nand U1889 (N_1889,N_1819,N_1837);
and U1890 (N_1890,N_1809,N_1845);
and U1891 (N_1891,N_1842,N_1825);
and U1892 (N_1892,N_1841,N_1829);
nor U1893 (N_1893,N_1833,N_1810);
nand U1894 (N_1894,N_1810,N_1838);
and U1895 (N_1895,N_1801,N_1844);
nor U1896 (N_1896,N_1818,N_1803);
nor U1897 (N_1897,N_1809,N_1840);
xor U1898 (N_1898,N_1816,N_1808);
nand U1899 (N_1899,N_1837,N_1839);
and U1900 (N_1900,N_1863,N_1861);
nor U1901 (N_1901,N_1864,N_1882);
or U1902 (N_1902,N_1896,N_1873);
or U1903 (N_1903,N_1898,N_1894);
and U1904 (N_1904,N_1859,N_1878);
nor U1905 (N_1905,N_1875,N_1855);
nand U1906 (N_1906,N_1871,N_1850);
or U1907 (N_1907,N_1854,N_1887);
nor U1908 (N_1908,N_1853,N_1862);
xnor U1909 (N_1909,N_1868,N_1869);
or U1910 (N_1910,N_1851,N_1899);
or U1911 (N_1911,N_1893,N_1870);
or U1912 (N_1912,N_1891,N_1865);
or U1913 (N_1913,N_1895,N_1897);
xor U1914 (N_1914,N_1867,N_1872);
or U1915 (N_1915,N_1880,N_1885);
and U1916 (N_1916,N_1877,N_1890);
nor U1917 (N_1917,N_1883,N_1858);
nor U1918 (N_1918,N_1881,N_1889);
and U1919 (N_1919,N_1888,N_1879);
nand U1920 (N_1920,N_1886,N_1856);
nor U1921 (N_1921,N_1857,N_1884);
or U1922 (N_1922,N_1876,N_1852);
or U1923 (N_1923,N_1874,N_1860);
or U1924 (N_1924,N_1892,N_1866);
or U1925 (N_1925,N_1874,N_1858);
or U1926 (N_1926,N_1879,N_1857);
nand U1927 (N_1927,N_1886,N_1888);
or U1928 (N_1928,N_1883,N_1872);
or U1929 (N_1929,N_1892,N_1874);
nor U1930 (N_1930,N_1890,N_1861);
and U1931 (N_1931,N_1882,N_1893);
nand U1932 (N_1932,N_1877,N_1896);
nand U1933 (N_1933,N_1880,N_1854);
and U1934 (N_1934,N_1864,N_1851);
nand U1935 (N_1935,N_1888,N_1868);
nor U1936 (N_1936,N_1890,N_1855);
xnor U1937 (N_1937,N_1866,N_1894);
nand U1938 (N_1938,N_1883,N_1862);
nand U1939 (N_1939,N_1889,N_1861);
nor U1940 (N_1940,N_1862,N_1897);
or U1941 (N_1941,N_1874,N_1857);
and U1942 (N_1942,N_1899,N_1893);
and U1943 (N_1943,N_1851,N_1874);
nand U1944 (N_1944,N_1891,N_1860);
nor U1945 (N_1945,N_1866,N_1860);
or U1946 (N_1946,N_1895,N_1877);
nor U1947 (N_1947,N_1858,N_1894);
or U1948 (N_1948,N_1893,N_1875);
nor U1949 (N_1949,N_1869,N_1893);
nor U1950 (N_1950,N_1912,N_1924);
nor U1951 (N_1951,N_1938,N_1906);
or U1952 (N_1952,N_1926,N_1932);
nand U1953 (N_1953,N_1941,N_1902);
nand U1954 (N_1954,N_1934,N_1905);
nor U1955 (N_1955,N_1916,N_1940);
nand U1956 (N_1956,N_1915,N_1900);
or U1957 (N_1957,N_1946,N_1909);
or U1958 (N_1958,N_1908,N_1942);
nand U1959 (N_1959,N_1913,N_1937);
and U1960 (N_1960,N_1928,N_1910);
nor U1961 (N_1961,N_1933,N_1945);
xor U1962 (N_1962,N_1944,N_1921);
xnor U1963 (N_1963,N_1949,N_1903);
or U1964 (N_1964,N_1901,N_1918);
and U1965 (N_1965,N_1930,N_1929);
and U1966 (N_1966,N_1907,N_1943);
or U1967 (N_1967,N_1923,N_1927);
or U1968 (N_1968,N_1914,N_1936);
and U1969 (N_1969,N_1948,N_1922);
nor U1970 (N_1970,N_1947,N_1920);
nand U1971 (N_1971,N_1939,N_1917);
nor U1972 (N_1972,N_1904,N_1925);
nand U1973 (N_1973,N_1931,N_1935);
nor U1974 (N_1974,N_1919,N_1911);
or U1975 (N_1975,N_1934,N_1917);
nand U1976 (N_1976,N_1935,N_1907);
xor U1977 (N_1977,N_1923,N_1940);
nand U1978 (N_1978,N_1939,N_1942);
nor U1979 (N_1979,N_1902,N_1935);
nor U1980 (N_1980,N_1921,N_1945);
and U1981 (N_1981,N_1937,N_1925);
nor U1982 (N_1982,N_1922,N_1937);
nor U1983 (N_1983,N_1945,N_1917);
and U1984 (N_1984,N_1920,N_1921);
nor U1985 (N_1985,N_1911,N_1945);
nand U1986 (N_1986,N_1931,N_1927);
nor U1987 (N_1987,N_1915,N_1909);
nor U1988 (N_1988,N_1920,N_1909);
or U1989 (N_1989,N_1931,N_1926);
nor U1990 (N_1990,N_1929,N_1910);
and U1991 (N_1991,N_1945,N_1949);
or U1992 (N_1992,N_1937,N_1901);
or U1993 (N_1993,N_1948,N_1927);
nor U1994 (N_1994,N_1922,N_1924);
and U1995 (N_1995,N_1910,N_1940);
and U1996 (N_1996,N_1922,N_1921);
and U1997 (N_1997,N_1930,N_1938);
nand U1998 (N_1998,N_1901,N_1948);
nor U1999 (N_1999,N_1906,N_1948);
or U2000 (N_2000,N_1989,N_1992);
or U2001 (N_2001,N_1973,N_1986);
nand U2002 (N_2002,N_1977,N_1965);
and U2003 (N_2003,N_1963,N_1982);
or U2004 (N_2004,N_1987,N_1985);
nand U2005 (N_2005,N_1954,N_1970);
nand U2006 (N_2006,N_1998,N_1974);
or U2007 (N_2007,N_1993,N_1972);
nor U2008 (N_2008,N_1961,N_1960);
and U2009 (N_2009,N_1999,N_1956);
nor U2010 (N_2010,N_1983,N_1958);
and U2011 (N_2011,N_1951,N_1955);
xor U2012 (N_2012,N_1997,N_1994);
nand U2013 (N_2013,N_1966,N_1981);
nor U2014 (N_2014,N_1953,N_1990);
xor U2015 (N_2015,N_1952,N_1979);
and U2016 (N_2016,N_1976,N_1991);
nor U2017 (N_2017,N_1980,N_1950);
nand U2018 (N_2018,N_1957,N_1995);
nand U2019 (N_2019,N_1959,N_1964);
and U2020 (N_2020,N_1962,N_1971);
xor U2021 (N_2021,N_1984,N_1988);
nand U2022 (N_2022,N_1969,N_1978);
nor U2023 (N_2023,N_1975,N_1968);
and U2024 (N_2024,N_1996,N_1967);
nand U2025 (N_2025,N_1965,N_1989);
nor U2026 (N_2026,N_1988,N_1955);
nand U2027 (N_2027,N_1956,N_1989);
and U2028 (N_2028,N_1967,N_1975);
nand U2029 (N_2029,N_1990,N_1995);
or U2030 (N_2030,N_1953,N_1950);
nor U2031 (N_2031,N_1980,N_1953);
nand U2032 (N_2032,N_1993,N_1955);
xnor U2033 (N_2033,N_1966,N_1956);
or U2034 (N_2034,N_1973,N_1968);
or U2035 (N_2035,N_1983,N_1987);
nor U2036 (N_2036,N_1983,N_1968);
nand U2037 (N_2037,N_1996,N_1976);
or U2038 (N_2038,N_1952,N_1982);
and U2039 (N_2039,N_1997,N_1951);
nor U2040 (N_2040,N_1957,N_1996);
and U2041 (N_2041,N_1956,N_1967);
and U2042 (N_2042,N_1979,N_1965);
nor U2043 (N_2043,N_1971,N_1969);
and U2044 (N_2044,N_1968,N_1955);
and U2045 (N_2045,N_1981,N_1994);
or U2046 (N_2046,N_1984,N_1959);
nor U2047 (N_2047,N_1977,N_1973);
nand U2048 (N_2048,N_1962,N_1956);
and U2049 (N_2049,N_1992,N_1970);
nand U2050 (N_2050,N_2036,N_2042);
nand U2051 (N_2051,N_2046,N_2020);
nand U2052 (N_2052,N_2005,N_2011);
and U2053 (N_2053,N_2031,N_2019);
and U2054 (N_2054,N_2006,N_2022);
nor U2055 (N_2055,N_2025,N_2017);
xnor U2056 (N_2056,N_2015,N_2044);
nor U2057 (N_2057,N_2026,N_2038);
nor U2058 (N_2058,N_2035,N_2039);
nor U2059 (N_2059,N_2023,N_2034);
and U2060 (N_2060,N_2009,N_2004);
nor U2061 (N_2061,N_2002,N_2045);
nor U2062 (N_2062,N_2048,N_2007);
and U2063 (N_2063,N_2008,N_2018);
and U2064 (N_2064,N_2033,N_2021);
or U2065 (N_2065,N_2047,N_2000);
or U2066 (N_2066,N_2027,N_2028);
nand U2067 (N_2067,N_2003,N_2012);
and U2068 (N_2068,N_2001,N_2013);
and U2069 (N_2069,N_2049,N_2041);
or U2070 (N_2070,N_2014,N_2037);
or U2071 (N_2071,N_2040,N_2024);
nor U2072 (N_2072,N_2030,N_2043);
or U2073 (N_2073,N_2016,N_2010);
and U2074 (N_2074,N_2029,N_2032);
or U2075 (N_2075,N_2031,N_2028);
or U2076 (N_2076,N_2020,N_2000);
and U2077 (N_2077,N_2048,N_2014);
nor U2078 (N_2078,N_2023,N_2005);
nand U2079 (N_2079,N_2009,N_2047);
nand U2080 (N_2080,N_2047,N_2024);
nand U2081 (N_2081,N_2027,N_2031);
nand U2082 (N_2082,N_2014,N_2001);
or U2083 (N_2083,N_2041,N_2013);
nand U2084 (N_2084,N_2038,N_2037);
nand U2085 (N_2085,N_2006,N_2023);
or U2086 (N_2086,N_2025,N_2001);
xor U2087 (N_2087,N_2021,N_2013);
nor U2088 (N_2088,N_2023,N_2016);
nand U2089 (N_2089,N_2048,N_2041);
nor U2090 (N_2090,N_2044,N_2032);
nor U2091 (N_2091,N_2043,N_2029);
or U2092 (N_2092,N_2003,N_2008);
xnor U2093 (N_2093,N_2016,N_2012);
and U2094 (N_2094,N_2045,N_2030);
nor U2095 (N_2095,N_2012,N_2001);
and U2096 (N_2096,N_2010,N_2035);
nand U2097 (N_2097,N_2030,N_2008);
nand U2098 (N_2098,N_2018,N_2004);
nand U2099 (N_2099,N_2011,N_2035);
nor U2100 (N_2100,N_2078,N_2080);
or U2101 (N_2101,N_2064,N_2055);
nand U2102 (N_2102,N_2063,N_2085);
or U2103 (N_2103,N_2054,N_2060);
nor U2104 (N_2104,N_2095,N_2090);
or U2105 (N_2105,N_2077,N_2081);
nor U2106 (N_2106,N_2051,N_2086);
or U2107 (N_2107,N_2059,N_2056);
and U2108 (N_2108,N_2097,N_2053);
nor U2109 (N_2109,N_2072,N_2088);
nand U2110 (N_2110,N_2098,N_2062);
nor U2111 (N_2111,N_2052,N_2087);
and U2112 (N_2112,N_2093,N_2057);
and U2113 (N_2113,N_2076,N_2061);
nor U2114 (N_2114,N_2096,N_2094);
nand U2115 (N_2115,N_2074,N_2073);
or U2116 (N_2116,N_2075,N_2091);
xnor U2117 (N_2117,N_2050,N_2092);
nor U2118 (N_2118,N_2082,N_2066);
nor U2119 (N_2119,N_2079,N_2071);
or U2120 (N_2120,N_2099,N_2065);
nand U2121 (N_2121,N_2067,N_2069);
nor U2122 (N_2122,N_2058,N_2070);
and U2123 (N_2123,N_2084,N_2089);
xor U2124 (N_2124,N_2083,N_2068);
nor U2125 (N_2125,N_2096,N_2054);
nand U2126 (N_2126,N_2096,N_2060);
xor U2127 (N_2127,N_2088,N_2071);
nor U2128 (N_2128,N_2078,N_2059);
or U2129 (N_2129,N_2093,N_2052);
nand U2130 (N_2130,N_2095,N_2072);
xor U2131 (N_2131,N_2050,N_2063);
nand U2132 (N_2132,N_2079,N_2092);
and U2133 (N_2133,N_2051,N_2094);
nor U2134 (N_2134,N_2061,N_2070);
nand U2135 (N_2135,N_2064,N_2061);
nor U2136 (N_2136,N_2056,N_2098);
or U2137 (N_2137,N_2086,N_2094);
nand U2138 (N_2138,N_2090,N_2061);
nor U2139 (N_2139,N_2068,N_2063);
nor U2140 (N_2140,N_2092,N_2054);
nand U2141 (N_2141,N_2060,N_2086);
nor U2142 (N_2142,N_2072,N_2084);
nand U2143 (N_2143,N_2092,N_2097);
nand U2144 (N_2144,N_2069,N_2065);
nor U2145 (N_2145,N_2098,N_2050);
and U2146 (N_2146,N_2054,N_2071);
nor U2147 (N_2147,N_2099,N_2053);
or U2148 (N_2148,N_2053,N_2076);
or U2149 (N_2149,N_2069,N_2058);
or U2150 (N_2150,N_2126,N_2147);
nand U2151 (N_2151,N_2104,N_2102);
and U2152 (N_2152,N_2109,N_2105);
nor U2153 (N_2153,N_2138,N_2128);
and U2154 (N_2154,N_2135,N_2120);
nand U2155 (N_2155,N_2121,N_2145);
or U2156 (N_2156,N_2103,N_2111);
or U2157 (N_2157,N_2118,N_2140);
nor U2158 (N_2158,N_2130,N_2134);
and U2159 (N_2159,N_2123,N_2124);
and U2160 (N_2160,N_2141,N_2136);
and U2161 (N_2161,N_2107,N_2131);
nand U2162 (N_2162,N_2149,N_2106);
nor U2163 (N_2163,N_2115,N_2117);
or U2164 (N_2164,N_2122,N_2143);
nor U2165 (N_2165,N_2137,N_2119);
nor U2166 (N_2166,N_2114,N_2116);
nor U2167 (N_2167,N_2146,N_2142);
or U2168 (N_2168,N_2133,N_2108);
nor U2169 (N_2169,N_2132,N_2148);
and U2170 (N_2170,N_2129,N_2125);
nor U2171 (N_2171,N_2112,N_2110);
nand U2172 (N_2172,N_2127,N_2113);
or U2173 (N_2173,N_2100,N_2139);
nor U2174 (N_2174,N_2101,N_2144);
xnor U2175 (N_2175,N_2105,N_2138);
nand U2176 (N_2176,N_2100,N_2112);
and U2177 (N_2177,N_2138,N_2132);
nand U2178 (N_2178,N_2144,N_2131);
nor U2179 (N_2179,N_2105,N_2139);
nand U2180 (N_2180,N_2113,N_2107);
or U2181 (N_2181,N_2141,N_2111);
or U2182 (N_2182,N_2103,N_2131);
and U2183 (N_2183,N_2110,N_2147);
nor U2184 (N_2184,N_2106,N_2138);
nand U2185 (N_2185,N_2135,N_2100);
nand U2186 (N_2186,N_2136,N_2130);
nand U2187 (N_2187,N_2139,N_2148);
nand U2188 (N_2188,N_2142,N_2141);
or U2189 (N_2189,N_2123,N_2101);
nand U2190 (N_2190,N_2122,N_2147);
xor U2191 (N_2191,N_2101,N_2112);
or U2192 (N_2192,N_2142,N_2114);
and U2193 (N_2193,N_2101,N_2105);
nor U2194 (N_2194,N_2108,N_2122);
nand U2195 (N_2195,N_2127,N_2136);
or U2196 (N_2196,N_2110,N_2125);
nor U2197 (N_2197,N_2114,N_2118);
nor U2198 (N_2198,N_2127,N_2138);
xor U2199 (N_2199,N_2143,N_2149);
and U2200 (N_2200,N_2186,N_2194);
or U2201 (N_2201,N_2174,N_2161);
and U2202 (N_2202,N_2196,N_2182);
or U2203 (N_2203,N_2179,N_2162);
and U2204 (N_2204,N_2157,N_2178);
nor U2205 (N_2205,N_2164,N_2180);
nor U2206 (N_2206,N_2156,N_2198);
nor U2207 (N_2207,N_2160,N_2187);
and U2208 (N_2208,N_2155,N_2195);
nor U2209 (N_2209,N_2183,N_2176);
nor U2210 (N_2210,N_2172,N_2177);
or U2211 (N_2211,N_2191,N_2153);
and U2212 (N_2212,N_2152,N_2189);
nand U2213 (N_2213,N_2150,N_2154);
or U2214 (N_2214,N_2158,N_2168);
nand U2215 (N_2215,N_2159,N_2151);
and U2216 (N_2216,N_2185,N_2190);
and U2217 (N_2217,N_2170,N_2188);
and U2218 (N_2218,N_2163,N_2171);
nor U2219 (N_2219,N_2192,N_2165);
nor U2220 (N_2220,N_2197,N_2167);
nand U2221 (N_2221,N_2181,N_2184);
or U2222 (N_2222,N_2173,N_2175);
and U2223 (N_2223,N_2166,N_2169);
nand U2224 (N_2224,N_2193,N_2199);
nand U2225 (N_2225,N_2151,N_2173);
xnor U2226 (N_2226,N_2185,N_2157);
nor U2227 (N_2227,N_2153,N_2193);
and U2228 (N_2228,N_2196,N_2185);
nor U2229 (N_2229,N_2163,N_2153);
and U2230 (N_2230,N_2185,N_2161);
xor U2231 (N_2231,N_2164,N_2188);
nor U2232 (N_2232,N_2168,N_2188);
nor U2233 (N_2233,N_2172,N_2197);
and U2234 (N_2234,N_2191,N_2183);
or U2235 (N_2235,N_2164,N_2171);
nor U2236 (N_2236,N_2192,N_2168);
nor U2237 (N_2237,N_2152,N_2178);
and U2238 (N_2238,N_2179,N_2156);
or U2239 (N_2239,N_2189,N_2185);
or U2240 (N_2240,N_2185,N_2152);
and U2241 (N_2241,N_2168,N_2173);
xor U2242 (N_2242,N_2181,N_2186);
nand U2243 (N_2243,N_2162,N_2165);
and U2244 (N_2244,N_2165,N_2177);
or U2245 (N_2245,N_2155,N_2158);
or U2246 (N_2246,N_2173,N_2169);
xor U2247 (N_2247,N_2150,N_2184);
nand U2248 (N_2248,N_2162,N_2152);
xor U2249 (N_2249,N_2196,N_2151);
nand U2250 (N_2250,N_2201,N_2215);
nand U2251 (N_2251,N_2206,N_2234);
nand U2252 (N_2252,N_2242,N_2247);
nor U2253 (N_2253,N_2200,N_2232);
nor U2254 (N_2254,N_2224,N_2205);
or U2255 (N_2255,N_2202,N_2237);
nor U2256 (N_2256,N_2214,N_2240);
nor U2257 (N_2257,N_2207,N_2244);
and U2258 (N_2258,N_2223,N_2246);
or U2259 (N_2259,N_2212,N_2213);
nand U2260 (N_2260,N_2219,N_2226);
nand U2261 (N_2261,N_2220,N_2233);
nand U2262 (N_2262,N_2231,N_2227);
nor U2263 (N_2263,N_2225,N_2238);
xnor U2264 (N_2264,N_2208,N_2222);
nand U2265 (N_2265,N_2230,N_2203);
nand U2266 (N_2266,N_2239,N_2235);
nand U2267 (N_2267,N_2210,N_2248);
nand U2268 (N_2268,N_2249,N_2209);
or U2269 (N_2269,N_2243,N_2204);
and U2270 (N_2270,N_2217,N_2216);
nor U2271 (N_2271,N_2221,N_2236);
or U2272 (N_2272,N_2211,N_2218);
and U2273 (N_2273,N_2228,N_2245);
and U2274 (N_2274,N_2229,N_2241);
nand U2275 (N_2275,N_2246,N_2234);
nor U2276 (N_2276,N_2244,N_2205);
xor U2277 (N_2277,N_2236,N_2230);
nand U2278 (N_2278,N_2224,N_2223);
nor U2279 (N_2279,N_2215,N_2233);
nand U2280 (N_2280,N_2241,N_2249);
and U2281 (N_2281,N_2243,N_2217);
and U2282 (N_2282,N_2204,N_2249);
and U2283 (N_2283,N_2204,N_2234);
and U2284 (N_2284,N_2212,N_2203);
nand U2285 (N_2285,N_2230,N_2212);
and U2286 (N_2286,N_2207,N_2233);
or U2287 (N_2287,N_2218,N_2207);
nand U2288 (N_2288,N_2245,N_2207);
nor U2289 (N_2289,N_2226,N_2210);
and U2290 (N_2290,N_2232,N_2205);
and U2291 (N_2291,N_2207,N_2232);
or U2292 (N_2292,N_2220,N_2207);
and U2293 (N_2293,N_2236,N_2233);
or U2294 (N_2294,N_2202,N_2243);
nor U2295 (N_2295,N_2214,N_2210);
and U2296 (N_2296,N_2229,N_2214);
and U2297 (N_2297,N_2217,N_2209);
nand U2298 (N_2298,N_2217,N_2233);
nand U2299 (N_2299,N_2201,N_2212);
nor U2300 (N_2300,N_2295,N_2260);
nor U2301 (N_2301,N_2256,N_2280);
and U2302 (N_2302,N_2294,N_2299);
and U2303 (N_2303,N_2264,N_2272);
nand U2304 (N_2304,N_2273,N_2288);
nor U2305 (N_2305,N_2275,N_2287);
nor U2306 (N_2306,N_2252,N_2266);
nand U2307 (N_2307,N_2283,N_2265);
and U2308 (N_2308,N_2292,N_2277);
or U2309 (N_2309,N_2262,N_2291);
nor U2310 (N_2310,N_2268,N_2276);
and U2311 (N_2311,N_2278,N_2296);
nand U2312 (N_2312,N_2251,N_2298);
or U2313 (N_2313,N_2282,N_2258);
nand U2314 (N_2314,N_2270,N_2279);
nor U2315 (N_2315,N_2269,N_2261);
nor U2316 (N_2316,N_2253,N_2271);
nand U2317 (N_2317,N_2250,N_2254);
and U2318 (N_2318,N_2289,N_2255);
nor U2319 (N_2319,N_2274,N_2286);
and U2320 (N_2320,N_2267,N_2257);
and U2321 (N_2321,N_2263,N_2281);
nor U2322 (N_2322,N_2285,N_2293);
nand U2323 (N_2323,N_2284,N_2259);
and U2324 (N_2324,N_2297,N_2290);
or U2325 (N_2325,N_2288,N_2261);
nor U2326 (N_2326,N_2252,N_2287);
or U2327 (N_2327,N_2264,N_2285);
and U2328 (N_2328,N_2280,N_2261);
and U2329 (N_2329,N_2299,N_2289);
and U2330 (N_2330,N_2263,N_2293);
nor U2331 (N_2331,N_2280,N_2250);
and U2332 (N_2332,N_2266,N_2292);
and U2333 (N_2333,N_2271,N_2259);
and U2334 (N_2334,N_2280,N_2255);
nor U2335 (N_2335,N_2277,N_2294);
nand U2336 (N_2336,N_2278,N_2297);
or U2337 (N_2337,N_2287,N_2250);
nand U2338 (N_2338,N_2262,N_2281);
xor U2339 (N_2339,N_2294,N_2265);
xnor U2340 (N_2340,N_2296,N_2255);
nand U2341 (N_2341,N_2286,N_2285);
nor U2342 (N_2342,N_2293,N_2287);
nor U2343 (N_2343,N_2271,N_2285);
nand U2344 (N_2344,N_2272,N_2297);
and U2345 (N_2345,N_2283,N_2282);
nor U2346 (N_2346,N_2275,N_2292);
or U2347 (N_2347,N_2250,N_2262);
xor U2348 (N_2348,N_2277,N_2291);
xor U2349 (N_2349,N_2285,N_2254);
nand U2350 (N_2350,N_2327,N_2341);
and U2351 (N_2351,N_2312,N_2321);
nand U2352 (N_2352,N_2302,N_2310);
nor U2353 (N_2353,N_2317,N_2332);
nor U2354 (N_2354,N_2308,N_2344);
nand U2355 (N_2355,N_2311,N_2339);
or U2356 (N_2356,N_2349,N_2319);
nor U2357 (N_2357,N_2330,N_2328);
nand U2358 (N_2358,N_2343,N_2315);
nor U2359 (N_2359,N_2326,N_2305);
or U2360 (N_2360,N_2329,N_2325);
nor U2361 (N_2361,N_2348,N_2323);
nor U2362 (N_2362,N_2301,N_2304);
xor U2363 (N_2363,N_2318,N_2324);
or U2364 (N_2364,N_2309,N_2303);
nor U2365 (N_2365,N_2338,N_2314);
nand U2366 (N_2366,N_2335,N_2337);
and U2367 (N_2367,N_2331,N_2333);
or U2368 (N_2368,N_2306,N_2342);
or U2369 (N_2369,N_2316,N_2313);
and U2370 (N_2370,N_2300,N_2345);
nand U2371 (N_2371,N_2307,N_2346);
or U2372 (N_2372,N_2340,N_2334);
nor U2373 (N_2373,N_2322,N_2347);
nand U2374 (N_2374,N_2320,N_2336);
or U2375 (N_2375,N_2348,N_2337);
nor U2376 (N_2376,N_2318,N_2349);
and U2377 (N_2377,N_2327,N_2303);
or U2378 (N_2378,N_2320,N_2315);
nand U2379 (N_2379,N_2340,N_2315);
or U2380 (N_2380,N_2317,N_2347);
nor U2381 (N_2381,N_2305,N_2344);
nor U2382 (N_2382,N_2341,N_2339);
nor U2383 (N_2383,N_2336,N_2345);
nand U2384 (N_2384,N_2339,N_2302);
nand U2385 (N_2385,N_2339,N_2323);
and U2386 (N_2386,N_2337,N_2319);
nor U2387 (N_2387,N_2345,N_2342);
nand U2388 (N_2388,N_2312,N_2335);
or U2389 (N_2389,N_2348,N_2339);
and U2390 (N_2390,N_2321,N_2349);
nor U2391 (N_2391,N_2323,N_2349);
nand U2392 (N_2392,N_2319,N_2310);
and U2393 (N_2393,N_2332,N_2335);
and U2394 (N_2394,N_2343,N_2320);
nor U2395 (N_2395,N_2302,N_2327);
or U2396 (N_2396,N_2337,N_2321);
or U2397 (N_2397,N_2308,N_2347);
and U2398 (N_2398,N_2318,N_2312);
nand U2399 (N_2399,N_2306,N_2332);
and U2400 (N_2400,N_2364,N_2383);
or U2401 (N_2401,N_2397,N_2350);
nor U2402 (N_2402,N_2389,N_2353);
or U2403 (N_2403,N_2379,N_2394);
or U2404 (N_2404,N_2360,N_2376);
and U2405 (N_2405,N_2393,N_2373);
nand U2406 (N_2406,N_2384,N_2390);
nand U2407 (N_2407,N_2378,N_2395);
xor U2408 (N_2408,N_2396,N_2359);
and U2409 (N_2409,N_2388,N_2392);
or U2410 (N_2410,N_2377,N_2354);
xnor U2411 (N_2411,N_2351,N_2386);
and U2412 (N_2412,N_2356,N_2367);
or U2413 (N_2413,N_2385,N_2372);
nand U2414 (N_2414,N_2361,N_2366);
and U2415 (N_2415,N_2370,N_2380);
nand U2416 (N_2416,N_2381,N_2398);
or U2417 (N_2417,N_2363,N_2369);
and U2418 (N_2418,N_2355,N_2365);
and U2419 (N_2419,N_2387,N_2368);
nand U2420 (N_2420,N_2374,N_2352);
or U2421 (N_2421,N_2357,N_2375);
nor U2422 (N_2422,N_2362,N_2358);
nand U2423 (N_2423,N_2382,N_2391);
nor U2424 (N_2424,N_2371,N_2399);
nor U2425 (N_2425,N_2389,N_2369);
nand U2426 (N_2426,N_2381,N_2372);
nor U2427 (N_2427,N_2361,N_2383);
nand U2428 (N_2428,N_2365,N_2387);
or U2429 (N_2429,N_2384,N_2364);
or U2430 (N_2430,N_2378,N_2392);
or U2431 (N_2431,N_2380,N_2387);
and U2432 (N_2432,N_2365,N_2368);
nand U2433 (N_2433,N_2357,N_2379);
or U2434 (N_2434,N_2381,N_2390);
nand U2435 (N_2435,N_2375,N_2350);
nor U2436 (N_2436,N_2352,N_2370);
nand U2437 (N_2437,N_2399,N_2352);
or U2438 (N_2438,N_2367,N_2357);
or U2439 (N_2439,N_2370,N_2359);
or U2440 (N_2440,N_2358,N_2350);
and U2441 (N_2441,N_2375,N_2383);
nand U2442 (N_2442,N_2388,N_2355);
nand U2443 (N_2443,N_2397,N_2371);
nor U2444 (N_2444,N_2397,N_2388);
nor U2445 (N_2445,N_2382,N_2378);
nand U2446 (N_2446,N_2391,N_2371);
xnor U2447 (N_2447,N_2388,N_2375);
xnor U2448 (N_2448,N_2373,N_2392);
or U2449 (N_2449,N_2398,N_2376);
nor U2450 (N_2450,N_2434,N_2401);
or U2451 (N_2451,N_2418,N_2437);
or U2452 (N_2452,N_2408,N_2429);
xnor U2453 (N_2453,N_2428,N_2423);
and U2454 (N_2454,N_2447,N_2446);
nor U2455 (N_2455,N_2443,N_2415);
nor U2456 (N_2456,N_2427,N_2426);
nand U2457 (N_2457,N_2440,N_2403);
xnor U2458 (N_2458,N_2406,N_2414);
and U2459 (N_2459,N_2412,N_2449);
xnor U2460 (N_2460,N_2424,N_2444);
or U2461 (N_2461,N_2411,N_2416);
or U2462 (N_2462,N_2400,N_2422);
and U2463 (N_2463,N_2419,N_2439);
or U2464 (N_2464,N_2421,N_2438);
nand U2465 (N_2465,N_2445,N_2448);
or U2466 (N_2466,N_2442,N_2435);
nand U2467 (N_2467,N_2432,N_2409);
nand U2468 (N_2468,N_2417,N_2430);
nand U2469 (N_2469,N_2436,N_2420);
and U2470 (N_2470,N_2441,N_2425);
nand U2471 (N_2471,N_2431,N_2413);
or U2472 (N_2472,N_2407,N_2402);
nor U2473 (N_2473,N_2433,N_2404);
or U2474 (N_2474,N_2405,N_2410);
xor U2475 (N_2475,N_2430,N_2404);
or U2476 (N_2476,N_2417,N_2429);
nor U2477 (N_2477,N_2425,N_2424);
xor U2478 (N_2478,N_2403,N_2444);
xnor U2479 (N_2479,N_2423,N_2424);
nand U2480 (N_2480,N_2410,N_2441);
nand U2481 (N_2481,N_2418,N_2425);
nor U2482 (N_2482,N_2413,N_2414);
or U2483 (N_2483,N_2433,N_2414);
and U2484 (N_2484,N_2445,N_2414);
nand U2485 (N_2485,N_2428,N_2445);
nor U2486 (N_2486,N_2433,N_2436);
nor U2487 (N_2487,N_2421,N_2412);
nand U2488 (N_2488,N_2436,N_2422);
nor U2489 (N_2489,N_2418,N_2412);
nand U2490 (N_2490,N_2407,N_2412);
or U2491 (N_2491,N_2440,N_2405);
nand U2492 (N_2492,N_2440,N_2449);
and U2493 (N_2493,N_2442,N_2420);
nand U2494 (N_2494,N_2402,N_2400);
nor U2495 (N_2495,N_2446,N_2415);
nand U2496 (N_2496,N_2444,N_2410);
or U2497 (N_2497,N_2432,N_2433);
and U2498 (N_2498,N_2421,N_2425);
and U2499 (N_2499,N_2412,N_2431);
nor U2500 (N_2500,N_2486,N_2452);
nand U2501 (N_2501,N_2492,N_2488);
or U2502 (N_2502,N_2474,N_2460);
or U2503 (N_2503,N_2496,N_2463);
or U2504 (N_2504,N_2465,N_2497);
nand U2505 (N_2505,N_2457,N_2483);
and U2506 (N_2506,N_2482,N_2459);
nor U2507 (N_2507,N_2477,N_2491);
nor U2508 (N_2508,N_2470,N_2489);
nand U2509 (N_2509,N_2468,N_2480);
or U2510 (N_2510,N_2494,N_2478);
nor U2511 (N_2511,N_2484,N_2481);
nor U2512 (N_2512,N_2472,N_2462);
nand U2513 (N_2513,N_2466,N_2451);
nand U2514 (N_2514,N_2454,N_2493);
nor U2515 (N_2515,N_2455,N_2450);
and U2516 (N_2516,N_2479,N_2490);
nor U2517 (N_2517,N_2475,N_2473);
nand U2518 (N_2518,N_2461,N_2469);
or U2519 (N_2519,N_2464,N_2467);
nor U2520 (N_2520,N_2471,N_2498);
nor U2521 (N_2521,N_2485,N_2476);
nand U2522 (N_2522,N_2458,N_2453);
nand U2523 (N_2523,N_2499,N_2456);
nor U2524 (N_2524,N_2487,N_2495);
or U2525 (N_2525,N_2463,N_2456);
nand U2526 (N_2526,N_2460,N_2487);
nand U2527 (N_2527,N_2485,N_2454);
or U2528 (N_2528,N_2489,N_2499);
nor U2529 (N_2529,N_2485,N_2455);
nor U2530 (N_2530,N_2481,N_2495);
and U2531 (N_2531,N_2451,N_2474);
nand U2532 (N_2532,N_2481,N_2478);
or U2533 (N_2533,N_2477,N_2496);
and U2534 (N_2534,N_2494,N_2463);
or U2535 (N_2535,N_2470,N_2481);
nor U2536 (N_2536,N_2470,N_2482);
and U2537 (N_2537,N_2466,N_2450);
nor U2538 (N_2538,N_2454,N_2492);
nand U2539 (N_2539,N_2486,N_2461);
and U2540 (N_2540,N_2480,N_2454);
and U2541 (N_2541,N_2451,N_2497);
nor U2542 (N_2542,N_2454,N_2450);
xor U2543 (N_2543,N_2496,N_2466);
nor U2544 (N_2544,N_2492,N_2461);
and U2545 (N_2545,N_2463,N_2477);
and U2546 (N_2546,N_2471,N_2482);
or U2547 (N_2547,N_2487,N_2497);
and U2548 (N_2548,N_2452,N_2478);
nand U2549 (N_2549,N_2464,N_2499);
nor U2550 (N_2550,N_2531,N_2522);
and U2551 (N_2551,N_2528,N_2545);
nor U2552 (N_2552,N_2532,N_2511);
nand U2553 (N_2553,N_2536,N_2529);
nand U2554 (N_2554,N_2510,N_2516);
nand U2555 (N_2555,N_2542,N_2515);
nor U2556 (N_2556,N_2537,N_2533);
or U2557 (N_2557,N_2526,N_2502);
nand U2558 (N_2558,N_2548,N_2527);
and U2559 (N_2559,N_2543,N_2546);
or U2560 (N_2560,N_2539,N_2521);
nand U2561 (N_2561,N_2504,N_2507);
xor U2562 (N_2562,N_2512,N_2509);
nor U2563 (N_2563,N_2530,N_2534);
nor U2564 (N_2564,N_2514,N_2547);
nor U2565 (N_2565,N_2500,N_2513);
nand U2566 (N_2566,N_2505,N_2506);
and U2567 (N_2567,N_2549,N_2523);
nor U2568 (N_2568,N_2520,N_2544);
nand U2569 (N_2569,N_2503,N_2508);
xor U2570 (N_2570,N_2540,N_2525);
and U2571 (N_2571,N_2538,N_2501);
nor U2572 (N_2572,N_2517,N_2519);
and U2573 (N_2573,N_2518,N_2535);
or U2574 (N_2574,N_2541,N_2524);
nand U2575 (N_2575,N_2534,N_2549);
or U2576 (N_2576,N_2503,N_2516);
or U2577 (N_2577,N_2509,N_2501);
or U2578 (N_2578,N_2545,N_2536);
and U2579 (N_2579,N_2534,N_2522);
and U2580 (N_2580,N_2520,N_2545);
nand U2581 (N_2581,N_2523,N_2522);
and U2582 (N_2582,N_2534,N_2512);
nand U2583 (N_2583,N_2522,N_2515);
or U2584 (N_2584,N_2546,N_2500);
or U2585 (N_2585,N_2533,N_2521);
nor U2586 (N_2586,N_2522,N_2524);
nor U2587 (N_2587,N_2526,N_2527);
and U2588 (N_2588,N_2540,N_2538);
nor U2589 (N_2589,N_2517,N_2531);
nand U2590 (N_2590,N_2542,N_2543);
and U2591 (N_2591,N_2517,N_2502);
nand U2592 (N_2592,N_2546,N_2542);
nor U2593 (N_2593,N_2538,N_2528);
and U2594 (N_2594,N_2534,N_2529);
and U2595 (N_2595,N_2501,N_2506);
nand U2596 (N_2596,N_2533,N_2529);
and U2597 (N_2597,N_2517,N_2540);
or U2598 (N_2598,N_2549,N_2528);
nor U2599 (N_2599,N_2511,N_2547);
and U2600 (N_2600,N_2586,N_2598);
and U2601 (N_2601,N_2584,N_2585);
and U2602 (N_2602,N_2588,N_2557);
nand U2603 (N_2603,N_2561,N_2596);
and U2604 (N_2604,N_2594,N_2564);
nor U2605 (N_2605,N_2581,N_2590);
nor U2606 (N_2606,N_2582,N_2566);
nor U2607 (N_2607,N_2579,N_2560);
nor U2608 (N_2608,N_2578,N_2552);
or U2609 (N_2609,N_2575,N_2553);
and U2610 (N_2610,N_2554,N_2593);
nand U2611 (N_2611,N_2563,N_2595);
and U2612 (N_2612,N_2570,N_2550);
and U2613 (N_2613,N_2556,N_2599);
nor U2614 (N_2614,N_2576,N_2577);
and U2615 (N_2615,N_2572,N_2580);
or U2616 (N_2616,N_2587,N_2573);
and U2617 (N_2617,N_2568,N_2589);
nand U2618 (N_2618,N_2551,N_2592);
and U2619 (N_2619,N_2591,N_2559);
and U2620 (N_2620,N_2571,N_2562);
nor U2621 (N_2621,N_2558,N_2555);
or U2622 (N_2622,N_2569,N_2574);
nand U2623 (N_2623,N_2567,N_2565);
and U2624 (N_2624,N_2597,N_2583);
or U2625 (N_2625,N_2577,N_2560);
nand U2626 (N_2626,N_2550,N_2584);
or U2627 (N_2627,N_2561,N_2592);
and U2628 (N_2628,N_2560,N_2592);
or U2629 (N_2629,N_2578,N_2571);
nand U2630 (N_2630,N_2593,N_2553);
and U2631 (N_2631,N_2562,N_2557);
or U2632 (N_2632,N_2588,N_2563);
and U2633 (N_2633,N_2553,N_2594);
nor U2634 (N_2634,N_2593,N_2583);
or U2635 (N_2635,N_2599,N_2594);
or U2636 (N_2636,N_2595,N_2569);
nor U2637 (N_2637,N_2575,N_2567);
and U2638 (N_2638,N_2585,N_2562);
and U2639 (N_2639,N_2576,N_2588);
nor U2640 (N_2640,N_2577,N_2583);
or U2641 (N_2641,N_2560,N_2581);
nor U2642 (N_2642,N_2566,N_2579);
nand U2643 (N_2643,N_2578,N_2585);
nor U2644 (N_2644,N_2584,N_2568);
or U2645 (N_2645,N_2575,N_2584);
and U2646 (N_2646,N_2560,N_2584);
nand U2647 (N_2647,N_2585,N_2560);
nor U2648 (N_2648,N_2552,N_2597);
and U2649 (N_2649,N_2551,N_2589);
and U2650 (N_2650,N_2604,N_2631);
nor U2651 (N_2651,N_2641,N_2600);
nand U2652 (N_2652,N_2610,N_2606);
nor U2653 (N_2653,N_2627,N_2637);
and U2654 (N_2654,N_2623,N_2632);
nor U2655 (N_2655,N_2636,N_2624);
nor U2656 (N_2656,N_2646,N_2620);
nand U2657 (N_2657,N_2614,N_2615);
nand U2658 (N_2658,N_2639,N_2602);
or U2659 (N_2659,N_2625,N_2616);
and U2660 (N_2660,N_2605,N_2611);
nand U2661 (N_2661,N_2633,N_2645);
or U2662 (N_2662,N_2617,N_2612);
or U2663 (N_2663,N_2648,N_2630);
or U2664 (N_2664,N_2619,N_2613);
nor U2665 (N_2665,N_2608,N_2628);
or U2666 (N_2666,N_2647,N_2618);
and U2667 (N_2667,N_2603,N_2621);
or U2668 (N_2668,N_2634,N_2643);
and U2669 (N_2669,N_2622,N_2626);
nor U2670 (N_2670,N_2629,N_2638);
nand U2671 (N_2671,N_2642,N_2640);
nor U2672 (N_2672,N_2607,N_2635);
nor U2673 (N_2673,N_2649,N_2609);
nor U2674 (N_2674,N_2601,N_2644);
nand U2675 (N_2675,N_2617,N_2605);
or U2676 (N_2676,N_2618,N_2609);
and U2677 (N_2677,N_2640,N_2624);
and U2678 (N_2678,N_2642,N_2611);
and U2679 (N_2679,N_2636,N_2629);
or U2680 (N_2680,N_2617,N_2636);
or U2681 (N_2681,N_2616,N_2606);
nand U2682 (N_2682,N_2643,N_2622);
nand U2683 (N_2683,N_2646,N_2645);
nor U2684 (N_2684,N_2631,N_2618);
and U2685 (N_2685,N_2606,N_2635);
or U2686 (N_2686,N_2611,N_2625);
nor U2687 (N_2687,N_2631,N_2646);
and U2688 (N_2688,N_2635,N_2647);
or U2689 (N_2689,N_2630,N_2633);
nor U2690 (N_2690,N_2607,N_2610);
nand U2691 (N_2691,N_2630,N_2608);
or U2692 (N_2692,N_2647,N_2643);
nand U2693 (N_2693,N_2639,N_2644);
nor U2694 (N_2694,N_2603,N_2626);
and U2695 (N_2695,N_2626,N_2637);
nand U2696 (N_2696,N_2638,N_2646);
or U2697 (N_2697,N_2603,N_2633);
nor U2698 (N_2698,N_2602,N_2629);
nand U2699 (N_2699,N_2631,N_2649);
and U2700 (N_2700,N_2672,N_2687);
nor U2701 (N_2701,N_2688,N_2654);
nor U2702 (N_2702,N_2681,N_2669);
and U2703 (N_2703,N_2676,N_2692);
nor U2704 (N_2704,N_2682,N_2683);
and U2705 (N_2705,N_2695,N_2674);
nand U2706 (N_2706,N_2699,N_2698);
nand U2707 (N_2707,N_2696,N_2660);
or U2708 (N_2708,N_2656,N_2667);
nand U2709 (N_2709,N_2684,N_2693);
nand U2710 (N_2710,N_2668,N_2651);
nand U2711 (N_2711,N_2685,N_2678);
or U2712 (N_2712,N_2690,N_2666);
and U2713 (N_2713,N_2680,N_2661);
nand U2714 (N_2714,N_2658,N_2664);
and U2715 (N_2715,N_2673,N_2689);
nor U2716 (N_2716,N_2691,N_2697);
nand U2717 (N_2717,N_2653,N_2665);
and U2718 (N_2718,N_2655,N_2650);
nor U2719 (N_2719,N_2659,N_2686);
nand U2720 (N_2720,N_2670,N_2657);
nor U2721 (N_2721,N_2675,N_2677);
and U2722 (N_2722,N_2671,N_2679);
and U2723 (N_2723,N_2652,N_2662);
nand U2724 (N_2724,N_2694,N_2663);
nor U2725 (N_2725,N_2665,N_2658);
or U2726 (N_2726,N_2694,N_2699);
nand U2727 (N_2727,N_2671,N_2656);
nor U2728 (N_2728,N_2676,N_2686);
and U2729 (N_2729,N_2657,N_2689);
or U2730 (N_2730,N_2671,N_2658);
or U2731 (N_2731,N_2663,N_2665);
or U2732 (N_2732,N_2683,N_2669);
nand U2733 (N_2733,N_2683,N_2691);
and U2734 (N_2734,N_2698,N_2655);
xor U2735 (N_2735,N_2673,N_2658);
nand U2736 (N_2736,N_2676,N_2673);
nand U2737 (N_2737,N_2691,N_2651);
nor U2738 (N_2738,N_2678,N_2668);
and U2739 (N_2739,N_2650,N_2652);
nor U2740 (N_2740,N_2684,N_2655);
and U2741 (N_2741,N_2695,N_2656);
nor U2742 (N_2742,N_2682,N_2652);
nor U2743 (N_2743,N_2692,N_2664);
nor U2744 (N_2744,N_2671,N_2664);
nand U2745 (N_2745,N_2651,N_2652);
and U2746 (N_2746,N_2691,N_2665);
nand U2747 (N_2747,N_2658,N_2668);
and U2748 (N_2748,N_2653,N_2691);
and U2749 (N_2749,N_2655,N_2689);
and U2750 (N_2750,N_2732,N_2729);
nand U2751 (N_2751,N_2727,N_2718);
or U2752 (N_2752,N_2713,N_2741);
and U2753 (N_2753,N_2740,N_2737);
or U2754 (N_2754,N_2747,N_2721);
and U2755 (N_2755,N_2730,N_2700);
or U2756 (N_2756,N_2733,N_2726);
and U2757 (N_2757,N_2739,N_2734);
xor U2758 (N_2758,N_2701,N_2717);
nand U2759 (N_2759,N_2731,N_2748);
nor U2760 (N_2760,N_2706,N_2704);
nand U2761 (N_2761,N_2728,N_2720);
nor U2762 (N_2762,N_2744,N_2735);
nor U2763 (N_2763,N_2714,N_2724);
xnor U2764 (N_2764,N_2710,N_2749);
or U2765 (N_2765,N_2707,N_2736);
nor U2766 (N_2766,N_2711,N_2712);
and U2767 (N_2767,N_2708,N_2746);
nand U2768 (N_2768,N_2705,N_2719);
and U2769 (N_2769,N_2745,N_2743);
nor U2770 (N_2770,N_2722,N_2702);
nand U2771 (N_2771,N_2703,N_2716);
nand U2772 (N_2772,N_2709,N_2738);
nand U2773 (N_2773,N_2723,N_2742);
nand U2774 (N_2774,N_2715,N_2725);
nor U2775 (N_2775,N_2720,N_2732);
and U2776 (N_2776,N_2712,N_2717);
and U2777 (N_2777,N_2714,N_2740);
nor U2778 (N_2778,N_2742,N_2707);
nor U2779 (N_2779,N_2723,N_2747);
and U2780 (N_2780,N_2704,N_2715);
nor U2781 (N_2781,N_2739,N_2725);
nand U2782 (N_2782,N_2717,N_2703);
nor U2783 (N_2783,N_2746,N_2747);
nor U2784 (N_2784,N_2747,N_2702);
or U2785 (N_2785,N_2704,N_2725);
nor U2786 (N_2786,N_2700,N_2743);
or U2787 (N_2787,N_2715,N_2706);
and U2788 (N_2788,N_2707,N_2709);
xnor U2789 (N_2789,N_2730,N_2707);
nor U2790 (N_2790,N_2741,N_2747);
and U2791 (N_2791,N_2720,N_2746);
nor U2792 (N_2792,N_2707,N_2718);
or U2793 (N_2793,N_2700,N_2706);
and U2794 (N_2794,N_2714,N_2720);
and U2795 (N_2795,N_2749,N_2729);
and U2796 (N_2796,N_2721,N_2712);
or U2797 (N_2797,N_2704,N_2714);
nand U2798 (N_2798,N_2732,N_2718);
and U2799 (N_2799,N_2749,N_2705);
nand U2800 (N_2800,N_2795,N_2782);
nor U2801 (N_2801,N_2785,N_2783);
and U2802 (N_2802,N_2786,N_2797);
nand U2803 (N_2803,N_2779,N_2755);
and U2804 (N_2804,N_2753,N_2762);
nor U2805 (N_2805,N_2788,N_2799);
nand U2806 (N_2806,N_2777,N_2759);
and U2807 (N_2807,N_2767,N_2758);
xnor U2808 (N_2808,N_2793,N_2769);
nor U2809 (N_2809,N_2775,N_2760);
nor U2810 (N_2810,N_2781,N_2774);
or U2811 (N_2811,N_2790,N_2752);
nand U2812 (N_2812,N_2770,N_2765);
and U2813 (N_2813,N_2764,N_2784);
nor U2814 (N_2814,N_2768,N_2791);
nand U2815 (N_2815,N_2778,N_2761);
and U2816 (N_2816,N_2766,N_2754);
nor U2817 (N_2817,N_2756,N_2757);
nor U2818 (N_2818,N_2792,N_2794);
and U2819 (N_2819,N_2780,N_2798);
and U2820 (N_2820,N_2789,N_2787);
nand U2821 (N_2821,N_2750,N_2773);
or U2822 (N_2822,N_2776,N_2763);
and U2823 (N_2823,N_2771,N_2772);
and U2824 (N_2824,N_2796,N_2751);
nor U2825 (N_2825,N_2767,N_2757);
or U2826 (N_2826,N_2762,N_2767);
and U2827 (N_2827,N_2762,N_2755);
or U2828 (N_2828,N_2783,N_2782);
nor U2829 (N_2829,N_2782,N_2775);
nor U2830 (N_2830,N_2769,N_2796);
or U2831 (N_2831,N_2765,N_2766);
and U2832 (N_2832,N_2797,N_2754);
nor U2833 (N_2833,N_2787,N_2769);
nand U2834 (N_2834,N_2762,N_2751);
nor U2835 (N_2835,N_2762,N_2781);
or U2836 (N_2836,N_2771,N_2791);
nand U2837 (N_2837,N_2760,N_2750);
or U2838 (N_2838,N_2791,N_2790);
nor U2839 (N_2839,N_2782,N_2750);
or U2840 (N_2840,N_2759,N_2754);
nand U2841 (N_2841,N_2762,N_2796);
nand U2842 (N_2842,N_2767,N_2780);
or U2843 (N_2843,N_2759,N_2763);
or U2844 (N_2844,N_2793,N_2758);
nor U2845 (N_2845,N_2755,N_2787);
or U2846 (N_2846,N_2752,N_2770);
nand U2847 (N_2847,N_2794,N_2785);
nor U2848 (N_2848,N_2759,N_2781);
or U2849 (N_2849,N_2799,N_2760);
or U2850 (N_2850,N_2821,N_2847);
and U2851 (N_2851,N_2806,N_2848);
and U2852 (N_2852,N_2803,N_2811);
nor U2853 (N_2853,N_2830,N_2810);
or U2854 (N_2854,N_2818,N_2817);
xor U2855 (N_2855,N_2802,N_2827);
nor U2856 (N_2856,N_2849,N_2826);
and U2857 (N_2857,N_2814,N_2840);
or U2858 (N_2858,N_2822,N_2812);
or U2859 (N_2859,N_2836,N_2829);
or U2860 (N_2860,N_2844,N_2831);
or U2861 (N_2861,N_2832,N_2808);
or U2862 (N_2862,N_2820,N_2837);
and U2863 (N_2863,N_2839,N_2828);
nor U2864 (N_2864,N_2846,N_2816);
or U2865 (N_2865,N_2833,N_2804);
nand U2866 (N_2866,N_2815,N_2835);
and U2867 (N_2867,N_2813,N_2823);
and U2868 (N_2868,N_2809,N_2825);
nor U2869 (N_2869,N_2841,N_2834);
or U2870 (N_2870,N_2807,N_2838);
or U2871 (N_2871,N_2843,N_2845);
nand U2872 (N_2872,N_2801,N_2800);
nor U2873 (N_2873,N_2824,N_2819);
or U2874 (N_2874,N_2842,N_2805);
nand U2875 (N_2875,N_2811,N_2841);
nor U2876 (N_2876,N_2803,N_2826);
nor U2877 (N_2877,N_2814,N_2813);
and U2878 (N_2878,N_2804,N_2842);
xnor U2879 (N_2879,N_2832,N_2822);
nor U2880 (N_2880,N_2826,N_2844);
nand U2881 (N_2881,N_2845,N_2821);
nor U2882 (N_2882,N_2832,N_2834);
nor U2883 (N_2883,N_2830,N_2818);
nor U2884 (N_2884,N_2838,N_2804);
or U2885 (N_2885,N_2845,N_2836);
and U2886 (N_2886,N_2812,N_2839);
nor U2887 (N_2887,N_2849,N_2831);
nor U2888 (N_2888,N_2830,N_2804);
nand U2889 (N_2889,N_2818,N_2823);
or U2890 (N_2890,N_2826,N_2836);
nand U2891 (N_2891,N_2847,N_2826);
and U2892 (N_2892,N_2824,N_2848);
nor U2893 (N_2893,N_2817,N_2800);
nand U2894 (N_2894,N_2805,N_2822);
or U2895 (N_2895,N_2822,N_2816);
nor U2896 (N_2896,N_2832,N_2824);
or U2897 (N_2897,N_2849,N_2822);
nand U2898 (N_2898,N_2833,N_2845);
and U2899 (N_2899,N_2817,N_2810);
or U2900 (N_2900,N_2855,N_2869);
xnor U2901 (N_2901,N_2878,N_2899);
nor U2902 (N_2902,N_2851,N_2867);
nand U2903 (N_2903,N_2863,N_2872);
and U2904 (N_2904,N_2865,N_2881);
and U2905 (N_2905,N_2860,N_2893);
xor U2906 (N_2906,N_2894,N_2853);
and U2907 (N_2907,N_2866,N_2898);
or U2908 (N_2908,N_2877,N_2891);
nor U2909 (N_2909,N_2879,N_2883);
nor U2910 (N_2910,N_2889,N_2856);
nand U2911 (N_2911,N_2854,N_2885);
or U2912 (N_2912,N_2871,N_2868);
and U2913 (N_2913,N_2873,N_2875);
and U2914 (N_2914,N_2858,N_2895);
and U2915 (N_2915,N_2880,N_2850);
nand U2916 (N_2916,N_2886,N_2874);
or U2917 (N_2917,N_2861,N_2870);
and U2918 (N_2918,N_2864,N_2892);
nand U2919 (N_2919,N_2852,N_2862);
nor U2920 (N_2920,N_2890,N_2882);
nand U2921 (N_2921,N_2876,N_2887);
nand U2922 (N_2922,N_2859,N_2857);
and U2923 (N_2923,N_2888,N_2897);
or U2924 (N_2924,N_2896,N_2884);
nand U2925 (N_2925,N_2880,N_2868);
nor U2926 (N_2926,N_2855,N_2865);
or U2927 (N_2927,N_2890,N_2877);
nor U2928 (N_2928,N_2863,N_2858);
and U2929 (N_2929,N_2869,N_2865);
nor U2930 (N_2930,N_2887,N_2886);
and U2931 (N_2931,N_2877,N_2889);
nor U2932 (N_2932,N_2885,N_2873);
nand U2933 (N_2933,N_2854,N_2882);
or U2934 (N_2934,N_2867,N_2879);
nor U2935 (N_2935,N_2858,N_2872);
nor U2936 (N_2936,N_2870,N_2876);
nor U2937 (N_2937,N_2858,N_2874);
nand U2938 (N_2938,N_2868,N_2881);
nor U2939 (N_2939,N_2875,N_2854);
nor U2940 (N_2940,N_2896,N_2850);
nor U2941 (N_2941,N_2857,N_2871);
and U2942 (N_2942,N_2885,N_2850);
nand U2943 (N_2943,N_2858,N_2884);
or U2944 (N_2944,N_2861,N_2857);
nand U2945 (N_2945,N_2850,N_2899);
nand U2946 (N_2946,N_2866,N_2875);
xor U2947 (N_2947,N_2869,N_2890);
and U2948 (N_2948,N_2855,N_2898);
and U2949 (N_2949,N_2872,N_2897);
and U2950 (N_2950,N_2925,N_2941);
nor U2951 (N_2951,N_2923,N_2937);
or U2952 (N_2952,N_2935,N_2933);
and U2953 (N_2953,N_2944,N_2901);
nor U2954 (N_2954,N_2932,N_2916);
or U2955 (N_2955,N_2942,N_2911);
nor U2956 (N_2956,N_2920,N_2906);
or U2957 (N_2957,N_2907,N_2903);
and U2958 (N_2958,N_2945,N_2943);
nor U2959 (N_2959,N_2915,N_2927);
and U2960 (N_2960,N_2939,N_2917);
nor U2961 (N_2961,N_2931,N_2902);
or U2962 (N_2962,N_2918,N_2949);
or U2963 (N_2963,N_2908,N_2930);
nand U2964 (N_2964,N_2940,N_2905);
nand U2965 (N_2965,N_2904,N_2948);
nand U2966 (N_2966,N_2900,N_2928);
and U2967 (N_2967,N_2946,N_2913);
nand U2968 (N_2968,N_2938,N_2926);
nor U2969 (N_2969,N_2929,N_2934);
nand U2970 (N_2970,N_2936,N_2914);
or U2971 (N_2971,N_2947,N_2909);
and U2972 (N_2972,N_2912,N_2910);
nand U2973 (N_2973,N_2922,N_2924);
and U2974 (N_2974,N_2919,N_2921);
and U2975 (N_2975,N_2902,N_2917);
nand U2976 (N_2976,N_2928,N_2909);
nand U2977 (N_2977,N_2947,N_2949);
xor U2978 (N_2978,N_2915,N_2907);
nand U2979 (N_2979,N_2919,N_2918);
nand U2980 (N_2980,N_2934,N_2913);
or U2981 (N_2981,N_2910,N_2945);
and U2982 (N_2982,N_2939,N_2945);
nand U2983 (N_2983,N_2900,N_2903);
or U2984 (N_2984,N_2902,N_2944);
nand U2985 (N_2985,N_2917,N_2906);
nor U2986 (N_2986,N_2919,N_2947);
nor U2987 (N_2987,N_2923,N_2927);
or U2988 (N_2988,N_2918,N_2910);
and U2989 (N_2989,N_2909,N_2934);
nor U2990 (N_2990,N_2929,N_2919);
or U2991 (N_2991,N_2916,N_2935);
nand U2992 (N_2992,N_2901,N_2949);
or U2993 (N_2993,N_2938,N_2901);
and U2994 (N_2994,N_2923,N_2911);
nor U2995 (N_2995,N_2905,N_2910);
nor U2996 (N_2996,N_2900,N_2933);
or U2997 (N_2997,N_2938,N_2910);
nor U2998 (N_2998,N_2925,N_2906);
xnor U2999 (N_2999,N_2913,N_2900);
nor UO_0 (O_0,N_2960,N_2969);
or UO_1 (O_1,N_2978,N_2957);
nor UO_2 (O_2,N_2973,N_2988);
nand UO_3 (O_3,N_2980,N_2967);
nand UO_4 (O_4,N_2952,N_2962);
and UO_5 (O_5,N_2972,N_2954);
nand UO_6 (O_6,N_2989,N_2991);
nand UO_7 (O_7,N_2994,N_2982);
nand UO_8 (O_8,N_2981,N_2993);
nor UO_9 (O_9,N_2971,N_2995);
and UO_10 (O_10,N_2983,N_2997);
nand UO_11 (O_11,N_2975,N_2966);
nor UO_12 (O_12,N_2964,N_2986);
or UO_13 (O_13,N_2963,N_2979);
and UO_14 (O_14,N_2974,N_2961);
and UO_15 (O_15,N_2955,N_2987);
nand UO_16 (O_16,N_2992,N_2984);
or UO_17 (O_17,N_2976,N_2965);
or UO_18 (O_18,N_2951,N_2998);
and UO_19 (O_19,N_2985,N_2968);
and UO_20 (O_20,N_2959,N_2956);
nand UO_21 (O_21,N_2970,N_2990);
nor UO_22 (O_22,N_2950,N_2958);
nor UO_23 (O_23,N_2996,N_2999);
and UO_24 (O_24,N_2953,N_2977);
nor UO_25 (O_25,N_2954,N_2966);
and UO_26 (O_26,N_2967,N_2951);
or UO_27 (O_27,N_2973,N_2962);
nor UO_28 (O_28,N_2954,N_2967);
nor UO_29 (O_29,N_2962,N_2959);
or UO_30 (O_30,N_2964,N_2988);
or UO_31 (O_31,N_2991,N_2997);
and UO_32 (O_32,N_2955,N_2952);
or UO_33 (O_33,N_2990,N_2992);
nor UO_34 (O_34,N_2982,N_2981);
nor UO_35 (O_35,N_2981,N_2998);
and UO_36 (O_36,N_2983,N_2992);
or UO_37 (O_37,N_2982,N_2966);
or UO_38 (O_38,N_2985,N_2951);
or UO_39 (O_39,N_2962,N_2990);
and UO_40 (O_40,N_2966,N_2978);
and UO_41 (O_41,N_2970,N_2977);
or UO_42 (O_42,N_2976,N_2994);
nor UO_43 (O_43,N_2992,N_2969);
nand UO_44 (O_44,N_2961,N_2962);
and UO_45 (O_45,N_2983,N_2954);
or UO_46 (O_46,N_2956,N_2988);
and UO_47 (O_47,N_2987,N_2989);
nand UO_48 (O_48,N_2978,N_2997);
nand UO_49 (O_49,N_2993,N_2956);
xnor UO_50 (O_50,N_2966,N_2992);
and UO_51 (O_51,N_2952,N_2983);
nor UO_52 (O_52,N_2994,N_2993);
and UO_53 (O_53,N_2959,N_2982);
nor UO_54 (O_54,N_2961,N_2976);
nor UO_55 (O_55,N_2987,N_2972);
xor UO_56 (O_56,N_2976,N_2975);
or UO_57 (O_57,N_2982,N_2985);
nand UO_58 (O_58,N_2988,N_2952);
and UO_59 (O_59,N_2962,N_2972);
and UO_60 (O_60,N_2962,N_2997);
nand UO_61 (O_61,N_2965,N_2991);
nand UO_62 (O_62,N_2996,N_2956);
xnor UO_63 (O_63,N_2990,N_2997);
nor UO_64 (O_64,N_2971,N_2972);
and UO_65 (O_65,N_2953,N_2968);
and UO_66 (O_66,N_2975,N_2974);
nor UO_67 (O_67,N_2999,N_2954);
nor UO_68 (O_68,N_2954,N_2957);
nor UO_69 (O_69,N_2954,N_2993);
and UO_70 (O_70,N_2951,N_2952);
nand UO_71 (O_71,N_2955,N_2995);
nor UO_72 (O_72,N_2976,N_2999);
nor UO_73 (O_73,N_2951,N_2962);
or UO_74 (O_74,N_2976,N_2955);
nor UO_75 (O_75,N_2996,N_2952);
nor UO_76 (O_76,N_2984,N_2977);
or UO_77 (O_77,N_2999,N_2978);
nand UO_78 (O_78,N_2985,N_2961);
nor UO_79 (O_79,N_2999,N_2967);
and UO_80 (O_80,N_2974,N_2997);
nand UO_81 (O_81,N_2951,N_2979);
or UO_82 (O_82,N_2984,N_2999);
and UO_83 (O_83,N_2999,N_2993);
nor UO_84 (O_84,N_2952,N_2990);
or UO_85 (O_85,N_2997,N_2956);
or UO_86 (O_86,N_2951,N_2996);
and UO_87 (O_87,N_2994,N_2990);
nand UO_88 (O_88,N_2978,N_2958);
xnor UO_89 (O_89,N_2981,N_2971);
nand UO_90 (O_90,N_2994,N_2962);
or UO_91 (O_91,N_2989,N_2954);
nand UO_92 (O_92,N_2968,N_2989);
nor UO_93 (O_93,N_2980,N_2989);
nor UO_94 (O_94,N_2982,N_2978);
nand UO_95 (O_95,N_2955,N_2992);
nand UO_96 (O_96,N_2962,N_2966);
and UO_97 (O_97,N_2994,N_2965);
nand UO_98 (O_98,N_2984,N_2972);
xor UO_99 (O_99,N_2958,N_2984);
nor UO_100 (O_100,N_2956,N_2957);
nor UO_101 (O_101,N_2984,N_2982);
and UO_102 (O_102,N_2992,N_2963);
or UO_103 (O_103,N_2976,N_2960);
nor UO_104 (O_104,N_2968,N_2958);
nand UO_105 (O_105,N_2982,N_2988);
and UO_106 (O_106,N_2990,N_2979);
nor UO_107 (O_107,N_2992,N_2958);
and UO_108 (O_108,N_2968,N_2955);
or UO_109 (O_109,N_2989,N_2998);
nor UO_110 (O_110,N_2994,N_2959);
or UO_111 (O_111,N_2993,N_2969);
or UO_112 (O_112,N_2953,N_2984);
nand UO_113 (O_113,N_2956,N_2965);
nand UO_114 (O_114,N_2969,N_2950);
nor UO_115 (O_115,N_2991,N_2959);
or UO_116 (O_116,N_2991,N_2983);
or UO_117 (O_117,N_2972,N_2976);
or UO_118 (O_118,N_2979,N_2995);
nor UO_119 (O_119,N_2955,N_2991);
nor UO_120 (O_120,N_2958,N_2959);
or UO_121 (O_121,N_2984,N_2985);
and UO_122 (O_122,N_2997,N_2952);
nor UO_123 (O_123,N_2963,N_2958);
or UO_124 (O_124,N_2971,N_2951);
nand UO_125 (O_125,N_2962,N_2978);
nand UO_126 (O_126,N_2975,N_2990);
or UO_127 (O_127,N_2978,N_2952);
nand UO_128 (O_128,N_2983,N_2998);
nor UO_129 (O_129,N_2957,N_2959);
and UO_130 (O_130,N_2970,N_2978);
nand UO_131 (O_131,N_2956,N_2958);
xor UO_132 (O_132,N_2980,N_2994);
nor UO_133 (O_133,N_2986,N_2982);
xnor UO_134 (O_134,N_2984,N_2964);
nor UO_135 (O_135,N_2958,N_2979);
or UO_136 (O_136,N_2952,N_2979);
nand UO_137 (O_137,N_2965,N_2987);
and UO_138 (O_138,N_2999,N_2981);
xor UO_139 (O_139,N_2967,N_2957);
and UO_140 (O_140,N_2962,N_2950);
and UO_141 (O_141,N_2957,N_2984);
xor UO_142 (O_142,N_2981,N_2994);
nor UO_143 (O_143,N_2977,N_2967);
and UO_144 (O_144,N_2974,N_2995);
and UO_145 (O_145,N_2968,N_2952);
nand UO_146 (O_146,N_2992,N_2991);
nand UO_147 (O_147,N_2959,N_2955);
or UO_148 (O_148,N_2997,N_2957);
and UO_149 (O_149,N_2956,N_2973);
nand UO_150 (O_150,N_2965,N_2968);
and UO_151 (O_151,N_2976,N_2997);
and UO_152 (O_152,N_2952,N_2991);
nor UO_153 (O_153,N_2956,N_2991);
and UO_154 (O_154,N_2990,N_2976);
nand UO_155 (O_155,N_2971,N_2975);
and UO_156 (O_156,N_2961,N_2999);
and UO_157 (O_157,N_2959,N_2971);
nand UO_158 (O_158,N_2965,N_2977);
and UO_159 (O_159,N_2955,N_2964);
nor UO_160 (O_160,N_2984,N_2996);
and UO_161 (O_161,N_2996,N_2966);
or UO_162 (O_162,N_2981,N_2967);
nor UO_163 (O_163,N_2997,N_2986);
nor UO_164 (O_164,N_2985,N_2963);
and UO_165 (O_165,N_2955,N_2957);
nand UO_166 (O_166,N_2999,N_2992);
and UO_167 (O_167,N_2958,N_2974);
nor UO_168 (O_168,N_2953,N_2972);
nand UO_169 (O_169,N_2969,N_2995);
nor UO_170 (O_170,N_2962,N_2969);
or UO_171 (O_171,N_2989,N_2970);
nor UO_172 (O_172,N_2954,N_2995);
nand UO_173 (O_173,N_2959,N_2988);
nand UO_174 (O_174,N_2997,N_2998);
nor UO_175 (O_175,N_2995,N_2988);
nand UO_176 (O_176,N_2975,N_2984);
and UO_177 (O_177,N_2963,N_2959);
or UO_178 (O_178,N_2991,N_2994);
or UO_179 (O_179,N_2968,N_2975);
or UO_180 (O_180,N_2982,N_2980);
or UO_181 (O_181,N_2995,N_2987);
or UO_182 (O_182,N_2972,N_2978);
or UO_183 (O_183,N_2992,N_2994);
and UO_184 (O_184,N_2955,N_2970);
nor UO_185 (O_185,N_2955,N_2996);
nor UO_186 (O_186,N_2973,N_2967);
or UO_187 (O_187,N_2998,N_2990);
nand UO_188 (O_188,N_2996,N_2965);
nand UO_189 (O_189,N_2996,N_2954);
nor UO_190 (O_190,N_2993,N_2952);
nor UO_191 (O_191,N_2982,N_2970);
xnor UO_192 (O_192,N_2984,N_2974);
nand UO_193 (O_193,N_2958,N_2951);
and UO_194 (O_194,N_2996,N_2991);
or UO_195 (O_195,N_2979,N_2974);
nor UO_196 (O_196,N_2985,N_2976);
nand UO_197 (O_197,N_2996,N_2994);
or UO_198 (O_198,N_2970,N_2975);
nor UO_199 (O_199,N_2952,N_2966);
nand UO_200 (O_200,N_2958,N_2966);
or UO_201 (O_201,N_2986,N_2956);
and UO_202 (O_202,N_2987,N_2986);
nand UO_203 (O_203,N_2989,N_2975);
or UO_204 (O_204,N_2981,N_2966);
nor UO_205 (O_205,N_2977,N_2956);
or UO_206 (O_206,N_2990,N_2981);
and UO_207 (O_207,N_2966,N_2959);
nand UO_208 (O_208,N_2987,N_2996);
nand UO_209 (O_209,N_2971,N_2966);
nand UO_210 (O_210,N_2968,N_2996);
or UO_211 (O_211,N_2951,N_2963);
nor UO_212 (O_212,N_2980,N_2985);
or UO_213 (O_213,N_2988,N_2967);
nand UO_214 (O_214,N_2961,N_2960);
nor UO_215 (O_215,N_2991,N_2963);
nor UO_216 (O_216,N_2993,N_2957);
and UO_217 (O_217,N_2979,N_2981);
nand UO_218 (O_218,N_2991,N_2974);
nor UO_219 (O_219,N_2956,N_2999);
nand UO_220 (O_220,N_2987,N_2984);
or UO_221 (O_221,N_2996,N_2992);
nor UO_222 (O_222,N_2989,N_2996);
or UO_223 (O_223,N_2990,N_2957);
or UO_224 (O_224,N_2967,N_2982);
xnor UO_225 (O_225,N_2960,N_2972);
and UO_226 (O_226,N_2970,N_2968);
xor UO_227 (O_227,N_2968,N_2974);
or UO_228 (O_228,N_2976,N_2970);
or UO_229 (O_229,N_2976,N_2951);
xnor UO_230 (O_230,N_2972,N_2981);
or UO_231 (O_231,N_2984,N_2970);
and UO_232 (O_232,N_2980,N_2990);
nor UO_233 (O_233,N_2983,N_2964);
and UO_234 (O_234,N_2980,N_2956);
nor UO_235 (O_235,N_2977,N_2951);
nand UO_236 (O_236,N_2951,N_2954);
or UO_237 (O_237,N_2978,N_2960);
and UO_238 (O_238,N_2951,N_2981);
or UO_239 (O_239,N_2995,N_2967);
nor UO_240 (O_240,N_2990,N_2996);
and UO_241 (O_241,N_2976,N_2977);
nor UO_242 (O_242,N_2959,N_2997);
or UO_243 (O_243,N_2970,N_2965);
and UO_244 (O_244,N_2973,N_2975);
and UO_245 (O_245,N_2967,N_2961);
and UO_246 (O_246,N_2961,N_2965);
nor UO_247 (O_247,N_2986,N_2978);
or UO_248 (O_248,N_2996,N_2967);
or UO_249 (O_249,N_2973,N_2981);
nor UO_250 (O_250,N_2968,N_2973);
or UO_251 (O_251,N_2976,N_2988);
nand UO_252 (O_252,N_2971,N_2955);
and UO_253 (O_253,N_2993,N_2992);
or UO_254 (O_254,N_2957,N_2986);
nor UO_255 (O_255,N_2969,N_2983);
xor UO_256 (O_256,N_2950,N_2951);
or UO_257 (O_257,N_2977,N_2969);
nor UO_258 (O_258,N_2984,N_2986);
and UO_259 (O_259,N_2955,N_2966);
nand UO_260 (O_260,N_2955,N_2994);
nand UO_261 (O_261,N_2994,N_2961);
nor UO_262 (O_262,N_2966,N_2985);
and UO_263 (O_263,N_2992,N_2972);
nor UO_264 (O_264,N_2980,N_2993);
nand UO_265 (O_265,N_2970,N_2974);
nand UO_266 (O_266,N_2999,N_2986);
nor UO_267 (O_267,N_2981,N_2961);
xor UO_268 (O_268,N_2988,N_2963);
nand UO_269 (O_269,N_2961,N_2982);
nor UO_270 (O_270,N_2987,N_2991);
and UO_271 (O_271,N_2996,N_2963);
and UO_272 (O_272,N_2983,N_2995);
nand UO_273 (O_273,N_2997,N_2971);
xnor UO_274 (O_274,N_2985,N_2997);
nand UO_275 (O_275,N_2956,N_2964);
and UO_276 (O_276,N_2992,N_2975);
nor UO_277 (O_277,N_2967,N_2991);
and UO_278 (O_278,N_2964,N_2999);
xor UO_279 (O_279,N_2953,N_2956);
nor UO_280 (O_280,N_2960,N_2993);
nor UO_281 (O_281,N_2953,N_2980);
and UO_282 (O_282,N_2974,N_2989);
nand UO_283 (O_283,N_2958,N_2986);
and UO_284 (O_284,N_2999,N_2960);
and UO_285 (O_285,N_2993,N_2974);
nor UO_286 (O_286,N_2995,N_2970);
nor UO_287 (O_287,N_2993,N_2968);
nor UO_288 (O_288,N_2979,N_2960);
nor UO_289 (O_289,N_2960,N_2954);
nor UO_290 (O_290,N_2954,N_2970);
or UO_291 (O_291,N_2999,N_2962);
nor UO_292 (O_292,N_2969,N_2974);
and UO_293 (O_293,N_2985,N_2955);
and UO_294 (O_294,N_2962,N_2985);
nor UO_295 (O_295,N_2956,N_2961);
nand UO_296 (O_296,N_2964,N_2995);
or UO_297 (O_297,N_2950,N_2978);
or UO_298 (O_298,N_2982,N_2990);
xor UO_299 (O_299,N_2958,N_2989);
and UO_300 (O_300,N_2955,N_2977);
nand UO_301 (O_301,N_2975,N_2956);
nand UO_302 (O_302,N_2987,N_2960);
nor UO_303 (O_303,N_2987,N_2994);
nor UO_304 (O_304,N_2972,N_2994);
or UO_305 (O_305,N_2955,N_2961);
nand UO_306 (O_306,N_2958,N_2965);
nor UO_307 (O_307,N_2959,N_2951);
or UO_308 (O_308,N_2996,N_2969);
nand UO_309 (O_309,N_2990,N_2956);
or UO_310 (O_310,N_2993,N_2976);
nor UO_311 (O_311,N_2981,N_2978);
and UO_312 (O_312,N_2989,N_2995);
nor UO_313 (O_313,N_2957,N_2979);
nor UO_314 (O_314,N_2999,N_2977);
and UO_315 (O_315,N_2994,N_2974);
or UO_316 (O_316,N_2990,N_2973);
and UO_317 (O_317,N_2963,N_2986);
and UO_318 (O_318,N_2985,N_2954);
nor UO_319 (O_319,N_2977,N_2979);
or UO_320 (O_320,N_2955,N_2975);
or UO_321 (O_321,N_2983,N_2988);
and UO_322 (O_322,N_2968,N_2969);
and UO_323 (O_323,N_2981,N_2974);
and UO_324 (O_324,N_2981,N_2997);
and UO_325 (O_325,N_2992,N_2953);
or UO_326 (O_326,N_2988,N_2984);
and UO_327 (O_327,N_2956,N_2955);
and UO_328 (O_328,N_2995,N_2976);
nor UO_329 (O_329,N_2983,N_2972);
or UO_330 (O_330,N_2967,N_2987);
or UO_331 (O_331,N_2995,N_2999);
nand UO_332 (O_332,N_2965,N_2984);
nand UO_333 (O_333,N_2989,N_2961);
nand UO_334 (O_334,N_2995,N_2962);
or UO_335 (O_335,N_2999,N_2957);
nand UO_336 (O_336,N_2956,N_2978);
and UO_337 (O_337,N_2980,N_2992);
nand UO_338 (O_338,N_2996,N_2980);
or UO_339 (O_339,N_2952,N_2970);
and UO_340 (O_340,N_2984,N_2998);
and UO_341 (O_341,N_2979,N_2968);
and UO_342 (O_342,N_2961,N_2963);
nand UO_343 (O_343,N_2962,N_2964);
or UO_344 (O_344,N_2967,N_2993);
and UO_345 (O_345,N_2996,N_2977);
nand UO_346 (O_346,N_2984,N_2969);
and UO_347 (O_347,N_2973,N_2959);
and UO_348 (O_348,N_2955,N_2988);
and UO_349 (O_349,N_2961,N_2995);
nand UO_350 (O_350,N_2976,N_2950);
or UO_351 (O_351,N_2965,N_2989);
or UO_352 (O_352,N_2993,N_2982);
or UO_353 (O_353,N_2969,N_2957);
nor UO_354 (O_354,N_2985,N_2986);
nor UO_355 (O_355,N_2963,N_2974);
or UO_356 (O_356,N_2951,N_2989);
or UO_357 (O_357,N_2984,N_2981);
nand UO_358 (O_358,N_2983,N_2962);
nand UO_359 (O_359,N_2960,N_2964);
nor UO_360 (O_360,N_2964,N_2972);
and UO_361 (O_361,N_2965,N_2960);
and UO_362 (O_362,N_2975,N_2959);
and UO_363 (O_363,N_2967,N_2958);
and UO_364 (O_364,N_2997,N_2955);
nor UO_365 (O_365,N_2982,N_2950);
or UO_366 (O_366,N_2971,N_2974);
and UO_367 (O_367,N_2999,N_2970);
xnor UO_368 (O_368,N_2998,N_2964);
nor UO_369 (O_369,N_2958,N_2980);
or UO_370 (O_370,N_2958,N_2969);
or UO_371 (O_371,N_2973,N_2995);
nor UO_372 (O_372,N_2980,N_2981);
and UO_373 (O_373,N_2969,N_2997);
nand UO_374 (O_374,N_2963,N_2960);
nand UO_375 (O_375,N_2961,N_2983);
and UO_376 (O_376,N_2973,N_2960);
nand UO_377 (O_377,N_2982,N_2968);
nor UO_378 (O_378,N_2972,N_2993);
nand UO_379 (O_379,N_2966,N_2969);
and UO_380 (O_380,N_2983,N_2958);
nand UO_381 (O_381,N_2971,N_2987);
nor UO_382 (O_382,N_2958,N_2981);
and UO_383 (O_383,N_2950,N_2965);
nand UO_384 (O_384,N_2950,N_2960);
or UO_385 (O_385,N_2952,N_2985);
and UO_386 (O_386,N_2955,N_2978);
or UO_387 (O_387,N_2986,N_2960);
and UO_388 (O_388,N_2985,N_2964);
and UO_389 (O_389,N_2970,N_2957);
nand UO_390 (O_390,N_2973,N_2976);
nand UO_391 (O_391,N_2951,N_2961);
nor UO_392 (O_392,N_2975,N_2972);
and UO_393 (O_393,N_2985,N_2960);
and UO_394 (O_394,N_2999,N_2985);
nand UO_395 (O_395,N_2995,N_2951);
nand UO_396 (O_396,N_2956,N_2963);
nor UO_397 (O_397,N_2993,N_2986);
and UO_398 (O_398,N_2971,N_2986);
nor UO_399 (O_399,N_2988,N_2958);
nor UO_400 (O_400,N_2976,N_2966);
nand UO_401 (O_401,N_2972,N_2965);
nand UO_402 (O_402,N_2969,N_2961);
or UO_403 (O_403,N_2968,N_2954);
and UO_404 (O_404,N_2985,N_2979);
and UO_405 (O_405,N_2986,N_2962);
nor UO_406 (O_406,N_2971,N_2980);
and UO_407 (O_407,N_2971,N_2990);
nand UO_408 (O_408,N_2977,N_2966);
nand UO_409 (O_409,N_2963,N_2980);
nor UO_410 (O_410,N_2977,N_2960);
or UO_411 (O_411,N_2972,N_2982);
and UO_412 (O_412,N_2991,N_2986);
nor UO_413 (O_413,N_2982,N_2989);
nand UO_414 (O_414,N_2992,N_2968);
nor UO_415 (O_415,N_2982,N_2977);
or UO_416 (O_416,N_2966,N_2995);
nor UO_417 (O_417,N_2970,N_2980);
nor UO_418 (O_418,N_2986,N_2976);
nand UO_419 (O_419,N_2989,N_2990);
nand UO_420 (O_420,N_2953,N_2969);
and UO_421 (O_421,N_2960,N_2951);
and UO_422 (O_422,N_2976,N_2974);
and UO_423 (O_423,N_2996,N_2978);
nand UO_424 (O_424,N_2971,N_2994);
or UO_425 (O_425,N_2972,N_2950);
and UO_426 (O_426,N_2967,N_2968);
xor UO_427 (O_427,N_2973,N_2974);
and UO_428 (O_428,N_2980,N_2962);
or UO_429 (O_429,N_2964,N_2963);
and UO_430 (O_430,N_2977,N_2987);
nand UO_431 (O_431,N_2968,N_2961);
or UO_432 (O_432,N_2952,N_2977);
and UO_433 (O_433,N_2963,N_2999);
nor UO_434 (O_434,N_2983,N_2977);
nor UO_435 (O_435,N_2992,N_2961);
and UO_436 (O_436,N_2995,N_2977);
nand UO_437 (O_437,N_2982,N_2962);
and UO_438 (O_438,N_2983,N_2974);
and UO_439 (O_439,N_2983,N_2985);
and UO_440 (O_440,N_2972,N_2967);
or UO_441 (O_441,N_2969,N_2951);
or UO_442 (O_442,N_2973,N_2952);
and UO_443 (O_443,N_2993,N_2991);
nor UO_444 (O_444,N_2991,N_2979);
nand UO_445 (O_445,N_2966,N_2991);
nor UO_446 (O_446,N_2961,N_2977);
nand UO_447 (O_447,N_2986,N_2995);
and UO_448 (O_448,N_2974,N_2966);
or UO_449 (O_449,N_2957,N_2961);
or UO_450 (O_450,N_2954,N_2955);
or UO_451 (O_451,N_2968,N_2984);
xor UO_452 (O_452,N_2954,N_2997);
and UO_453 (O_453,N_2953,N_2981);
and UO_454 (O_454,N_2983,N_2957);
nor UO_455 (O_455,N_2974,N_2965);
nor UO_456 (O_456,N_2953,N_2974);
xnor UO_457 (O_457,N_2965,N_2980);
or UO_458 (O_458,N_2977,N_2968);
nand UO_459 (O_459,N_2952,N_2987);
nand UO_460 (O_460,N_2976,N_2956);
nor UO_461 (O_461,N_2989,N_2964);
or UO_462 (O_462,N_2974,N_2992);
or UO_463 (O_463,N_2957,N_2952);
or UO_464 (O_464,N_2951,N_2970);
nor UO_465 (O_465,N_2960,N_2953);
nand UO_466 (O_466,N_2995,N_2958);
nor UO_467 (O_467,N_2982,N_2973);
xnor UO_468 (O_468,N_2970,N_2994);
and UO_469 (O_469,N_2961,N_2959);
or UO_470 (O_470,N_2970,N_2964);
nor UO_471 (O_471,N_2993,N_2958);
nor UO_472 (O_472,N_2955,N_2983);
and UO_473 (O_473,N_2984,N_2956);
nand UO_474 (O_474,N_2982,N_2997);
or UO_475 (O_475,N_2960,N_2989);
nand UO_476 (O_476,N_2955,N_2981);
or UO_477 (O_477,N_2967,N_2966);
or UO_478 (O_478,N_2995,N_2994);
or UO_479 (O_479,N_2958,N_2961);
nor UO_480 (O_480,N_2963,N_2952);
or UO_481 (O_481,N_2961,N_2964);
or UO_482 (O_482,N_2993,N_2990);
and UO_483 (O_483,N_2977,N_2973);
and UO_484 (O_484,N_2971,N_2968);
and UO_485 (O_485,N_2986,N_2965);
nor UO_486 (O_486,N_2988,N_2968);
and UO_487 (O_487,N_2989,N_2999);
or UO_488 (O_488,N_2980,N_2952);
nand UO_489 (O_489,N_2950,N_2963);
nor UO_490 (O_490,N_2956,N_2954);
nor UO_491 (O_491,N_2973,N_2966);
nor UO_492 (O_492,N_2963,N_2994);
nor UO_493 (O_493,N_2987,N_2983);
nor UO_494 (O_494,N_2993,N_2964);
and UO_495 (O_495,N_2960,N_2982);
nand UO_496 (O_496,N_2953,N_2993);
and UO_497 (O_497,N_2970,N_2992);
nor UO_498 (O_498,N_2954,N_2952);
or UO_499 (O_499,N_2955,N_2973);
endmodule