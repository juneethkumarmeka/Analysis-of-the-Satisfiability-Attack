module basic_500_3000_500_30_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_66,In_98);
and U1 (N_1,In_231,In_91);
and U2 (N_2,In_203,In_334);
or U3 (N_3,In_264,In_35);
and U4 (N_4,In_87,In_377);
or U5 (N_5,In_415,In_317);
nor U6 (N_6,In_351,In_309);
nor U7 (N_7,In_305,In_330);
nand U8 (N_8,In_451,In_173);
and U9 (N_9,In_482,In_474);
nor U10 (N_10,In_47,In_219);
or U11 (N_11,In_23,In_29);
nor U12 (N_12,In_289,In_45);
or U13 (N_13,In_363,In_357);
or U14 (N_14,In_455,In_112);
or U15 (N_15,In_370,In_142);
nor U16 (N_16,In_46,In_213);
nand U17 (N_17,In_135,In_348);
and U18 (N_18,In_266,In_190);
and U19 (N_19,In_11,In_443);
nand U20 (N_20,In_389,In_332);
or U21 (N_21,In_373,In_324);
nand U22 (N_22,In_485,In_284);
and U23 (N_23,In_210,In_466);
nor U24 (N_24,In_43,In_413);
nand U25 (N_25,In_316,In_378);
nand U26 (N_26,In_115,In_322);
nand U27 (N_27,In_258,In_268);
or U28 (N_28,In_444,In_435);
xnor U29 (N_29,In_420,In_459);
or U30 (N_30,In_68,In_167);
nor U31 (N_31,In_414,In_279);
nand U32 (N_32,In_470,In_165);
or U33 (N_33,In_27,In_181);
and U34 (N_34,In_429,In_49);
and U35 (N_35,In_220,In_382);
and U36 (N_36,In_118,In_410);
nand U37 (N_37,In_411,In_297);
or U38 (N_38,In_217,In_247);
or U39 (N_39,In_280,In_250);
nor U40 (N_40,In_221,In_390);
or U41 (N_41,In_214,In_170);
nor U42 (N_42,In_368,In_67);
or U43 (N_43,In_248,In_261);
nand U44 (N_44,In_344,In_263);
and U45 (N_45,In_33,In_211);
xor U46 (N_46,In_469,In_407);
and U47 (N_47,In_44,In_426);
and U48 (N_48,In_7,In_256);
nand U49 (N_49,In_323,In_273);
nand U50 (N_50,In_207,In_109);
nand U51 (N_51,In_371,In_402);
nor U52 (N_52,In_433,In_171);
nor U53 (N_53,In_141,In_69);
xor U54 (N_54,In_304,In_34);
nor U55 (N_55,In_367,In_14);
or U56 (N_56,In_21,In_326);
nor U57 (N_57,In_137,In_178);
nor U58 (N_58,In_312,In_325);
xnor U59 (N_59,In_65,In_70);
nor U60 (N_60,In_86,In_216);
nor U61 (N_61,In_283,In_10);
nor U62 (N_62,In_270,In_352);
or U63 (N_63,In_193,In_106);
nor U64 (N_64,In_229,In_76);
or U65 (N_65,In_19,In_399);
nand U66 (N_66,In_179,In_240);
nor U67 (N_67,In_476,In_154);
and U68 (N_68,In_204,In_296);
nor U69 (N_69,In_6,In_396);
nand U70 (N_70,In_395,In_276);
or U71 (N_71,In_209,In_468);
or U72 (N_72,In_161,In_475);
xor U73 (N_73,In_483,In_77);
xor U74 (N_74,In_122,In_1);
nand U75 (N_75,In_465,In_132);
nor U76 (N_76,In_271,In_457);
or U77 (N_77,In_13,In_479);
or U78 (N_78,In_252,In_232);
and U79 (N_79,In_498,In_9);
nand U80 (N_80,In_195,In_120);
nor U81 (N_81,In_102,In_292);
nand U82 (N_82,In_405,In_439);
and U83 (N_83,In_484,In_196);
or U84 (N_84,In_274,In_15);
nor U85 (N_85,In_158,In_374);
and U86 (N_86,In_424,In_225);
or U87 (N_87,In_155,In_452);
nor U88 (N_88,In_172,In_152);
nand U89 (N_89,In_131,In_301);
and U90 (N_90,In_226,In_176);
nor U91 (N_91,In_62,In_79);
nand U92 (N_92,In_16,In_20);
nor U93 (N_93,In_281,In_93);
and U94 (N_94,In_480,In_150);
and U95 (N_95,In_146,In_100);
and U96 (N_96,In_477,In_318);
nand U97 (N_97,In_40,In_369);
and U98 (N_98,In_148,In_92);
and U99 (N_99,In_354,In_116);
nand U100 (N_100,In_129,In_398);
nand U101 (N_101,In_299,In_117);
nor U102 (N_102,In_61,N_99);
nand U103 (N_103,In_81,In_486);
and U104 (N_104,In_114,In_64);
or U105 (N_105,N_34,In_208);
and U106 (N_106,In_286,N_63);
nand U107 (N_107,In_104,N_47);
and U108 (N_108,In_139,In_495);
or U109 (N_109,In_244,In_138);
nor U110 (N_110,In_337,In_84);
and U111 (N_111,N_71,N_32);
or U112 (N_112,N_74,N_51);
and U113 (N_113,In_417,In_223);
or U114 (N_114,In_153,N_82);
or U115 (N_115,In_39,In_307);
xor U116 (N_116,In_267,In_5);
xor U117 (N_117,In_177,In_353);
nand U118 (N_118,In_463,In_206);
nor U119 (N_119,In_157,In_241);
nand U120 (N_120,In_434,N_59);
or U121 (N_121,N_37,In_242);
nand U122 (N_122,In_438,In_419);
nand U123 (N_123,In_383,In_50);
nor U124 (N_124,In_392,In_262);
or U125 (N_125,In_107,In_360);
nor U126 (N_126,In_364,N_52);
nand U127 (N_127,In_291,In_97);
nand U128 (N_128,In_487,In_386);
or U129 (N_129,In_57,In_53);
or U130 (N_130,In_460,In_347);
or U131 (N_131,N_97,In_278);
nand U132 (N_132,In_362,N_13);
xnor U133 (N_133,In_99,N_17);
nor U134 (N_134,In_28,In_346);
and U135 (N_135,N_73,N_21);
or U136 (N_136,In_388,In_412);
or U137 (N_137,In_227,In_42);
nand U138 (N_138,In_376,In_350);
or U139 (N_139,In_497,N_2);
or U140 (N_140,N_67,In_126);
or U141 (N_141,In_355,In_356);
and U142 (N_142,In_212,In_265);
or U143 (N_143,N_85,N_38);
or U144 (N_144,In_30,In_385);
nor U145 (N_145,In_272,In_82);
or U146 (N_146,In_427,N_43);
nand U147 (N_147,N_69,In_175);
and U148 (N_148,In_418,In_51);
nand U149 (N_149,In_366,In_311);
and U150 (N_150,In_259,In_313);
or U151 (N_151,In_215,In_111);
and U152 (N_152,In_235,N_70);
or U153 (N_153,In_473,N_15);
xor U154 (N_154,In_253,In_197);
or U155 (N_155,In_401,In_8);
and U156 (N_156,In_394,In_295);
and U157 (N_157,In_492,In_298);
and U158 (N_158,In_124,In_192);
nor U159 (N_159,In_308,In_381);
nand U160 (N_160,In_333,N_9);
or U161 (N_161,In_108,In_127);
and U162 (N_162,In_184,In_319);
nor U163 (N_163,N_96,N_24);
nand U164 (N_164,N_88,In_169);
and U165 (N_165,In_400,N_72);
and U166 (N_166,N_20,In_32);
nand U167 (N_167,In_56,N_62);
nor U168 (N_168,In_224,In_85);
xnor U169 (N_169,In_422,In_496);
nor U170 (N_170,In_423,In_233);
or U171 (N_171,In_60,In_293);
xnor U172 (N_172,In_37,In_163);
or U173 (N_173,In_143,N_91);
and U174 (N_174,In_269,In_257);
nand U175 (N_175,N_93,N_1);
nand U176 (N_176,In_290,In_130);
nor U177 (N_177,In_63,In_202);
or U178 (N_178,In_255,In_343);
nor U179 (N_179,In_52,N_12);
or U180 (N_180,In_391,N_18);
nand U181 (N_181,In_275,In_95);
nor U182 (N_182,In_121,In_431);
and U183 (N_183,In_320,In_321);
and U184 (N_184,In_341,N_10);
or U185 (N_185,N_53,In_440);
nand U186 (N_186,N_95,In_189);
xnor U187 (N_187,N_0,In_445);
nand U188 (N_188,In_285,In_478);
or U189 (N_189,N_83,In_187);
or U190 (N_190,In_234,In_499);
nand U191 (N_191,N_50,In_365);
nor U192 (N_192,In_302,In_294);
nand U193 (N_193,In_75,In_342);
nand U194 (N_194,In_41,In_162);
nor U195 (N_195,In_78,In_489);
or U196 (N_196,In_55,In_372);
and U197 (N_197,N_92,N_68);
nor U198 (N_198,In_4,In_110);
xnor U199 (N_199,In_464,N_28);
nor U200 (N_200,N_146,N_76);
and U201 (N_201,N_195,In_0);
and U202 (N_202,N_120,N_172);
or U203 (N_203,In_222,In_74);
nor U204 (N_204,In_287,N_152);
nor U205 (N_205,In_164,N_183);
xor U206 (N_206,In_144,In_125);
or U207 (N_207,N_94,In_243);
and U208 (N_208,In_387,In_185);
nor U209 (N_209,In_186,In_83);
nand U210 (N_210,In_315,In_228);
and U211 (N_211,In_123,N_30);
or U212 (N_212,N_173,In_218);
nor U213 (N_213,N_56,N_23);
and U214 (N_214,N_131,In_174);
nand U215 (N_215,In_329,N_41);
nand U216 (N_216,In_88,In_182);
nand U217 (N_217,N_167,In_277);
nand U218 (N_218,N_163,N_110);
nor U219 (N_219,In_408,N_144);
and U220 (N_220,N_33,N_44);
nand U221 (N_221,N_189,N_116);
nor U222 (N_222,In_448,N_108);
nand U223 (N_223,In_159,N_151);
and U224 (N_224,N_80,In_432);
and U225 (N_225,N_107,N_165);
nand U226 (N_226,N_86,N_123);
or U227 (N_227,In_38,N_182);
nand U228 (N_228,In_200,In_481);
and U229 (N_229,N_136,In_180);
nand U230 (N_230,In_236,In_441);
nand U231 (N_231,In_359,In_406);
nand U232 (N_232,N_87,In_306);
nor U233 (N_233,N_77,N_142);
nand U234 (N_234,In_430,N_161);
and U235 (N_235,N_104,N_16);
xor U236 (N_236,N_48,In_151);
nand U237 (N_237,In_90,N_155);
or U238 (N_238,N_111,In_17);
and U239 (N_239,In_339,N_178);
or U240 (N_240,N_185,N_78);
or U241 (N_241,N_46,N_19);
or U242 (N_242,In_437,In_336);
and U243 (N_243,In_327,N_115);
xor U244 (N_244,In_328,In_128);
and U245 (N_245,In_436,N_42);
and U246 (N_246,In_403,N_197);
nand U247 (N_247,In_314,N_118);
nor U248 (N_248,N_3,N_114);
nand U249 (N_249,N_58,In_201);
nand U250 (N_250,In_105,N_90);
or U251 (N_251,In_101,In_59);
or U252 (N_252,N_61,In_375);
or U253 (N_253,N_7,N_156);
or U254 (N_254,N_170,In_456);
nand U255 (N_255,In_22,N_127);
nand U256 (N_256,In_461,In_198);
nor U257 (N_257,In_73,N_191);
or U258 (N_258,N_198,N_181);
nor U259 (N_259,N_89,In_282);
nand U260 (N_260,In_380,In_239);
or U261 (N_261,N_22,N_65);
nand U262 (N_262,N_64,N_130);
and U263 (N_263,N_100,N_154);
and U264 (N_264,In_404,N_188);
nor U265 (N_265,N_138,In_71);
and U266 (N_266,N_49,In_446);
and U267 (N_267,In_96,In_349);
nor U268 (N_268,N_137,In_249);
nand U269 (N_269,N_157,In_24);
or U270 (N_270,In_421,In_428);
nor U271 (N_271,N_125,In_288);
or U272 (N_272,N_192,N_139);
and U273 (N_273,In_168,N_55);
nand U274 (N_274,In_133,N_177);
xnor U275 (N_275,In_134,N_147);
nor U276 (N_276,In_379,N_169);
nor U277 (N_277,N_14,N_193);
nor U278 (N_278,In_494,N_8);
nand U279 (N_279,N_171,N_140);
or U280 (N_280,N_54,In_25);
xor U281 (N_281,N_84,N_162);
xnor U282 (N_282,In_26,N_57);
and U283 (N_283,In_260,N_113);
or U284 (N_284,In_335,In_194);
or U285 (N_285,In_453,N_60);
nand U286 (N_286,In_493,N_153);
nor U287 (N_287,N_5,N_143);
nand U288 (N_288,N_4,In_245);
nor U289 (N_289,In_166,In_230);
nand U290 (N_290,N_150,N_36);
nor U291 (N_291,In_490,In_36);
nand U292 (N_292,N_174,N_164);
nor U293 (N_293,N_168,N_184);
and U294 (N_294,In_238,N_40);
nand U295 (N_295,In_358,N_119);
or U296 (N_296,N_102,N_148);
or U297 (N_297,N_196,In_488);
nor U298 (N_298,In_191,In_345);
and U299 (N_299,N_186,In_80);
xor U300 (N_300,N_244,N_226);
or U301 (N_301,N_35,In_393);
nor U302 (N_302,N_145,N_248);
and U303 (N_303,In_160,N_285);
xnor U304 (N_304,N_208,N_233);
and U305 (N_305,N_117,In_310);
nand U306 (N_306,N_290,N_219);
nor U307 (N_307,N_201,N_299);
xor U308 (N_308,N_128,N_75);
and U309 (N_309,N_112,N_133);
or U310 (N_310,In_140,N_293);
nor U311 (N_311,N_149,N_272);
nand U312 (N_312,N_220,In_361);
nor U313 (N_313,In_54,N_105);
or U314 (N_314,N_29,In_467);
nand U315 (N_315,N_209,N_200);
nand U316 (N_316,N_218,In_450);
nor U317 (N_317,In_254,N_269);
and U318 (N_318,In_156,In_58);
nand U319 (N_319,In_18,N_203);
and U320 (N_320,N_242,N_206);
and U321 (N_321,N_238,In_416);
nand U322 (N_322,N_241,N_227);
nor U323 (N_323,N_279,In_462);
nor U324 (N_324,N_225,In_205);
or U325 (N_325,N_45,N_205);
nand U326 (N_326,N_287,In_89);
and U327 (N_327,N_132,N_240);
and U328 (N_328,N_252,N_284);
nor U329 (N_329,N_246,N_271);
nand U330 (N_330,N_158,N_66);
xnor U331 (N_331,N_223,N_292);
and U332 (N_332,N_121,N_264);
and U333 (N_333,N_31,In_246);
nand U334 (N_334,N_190,N_25);
nand U335 (N_335,N_176,N_202);
and U336 (N_336,N_211,N_243);
nand U337 (N_337,N_274,N_249);
xnor U338 (N_338,In_454,N_295);
nor U339 (N_339,N_256,In_136);
or U340 (N_340,In_251,In_384);
nor U341 (N_341,N_278,N_26);
and U342 (N_342,In_397,In_113);
or U343 (N_343,N_263,N_199);
or U344 (N_344,N_257,In_471);
nor U345 (N_345,N_124,In_12);
and U346 (N_346,N_239,N_262);
and U347 (N_347,N_291,N_296);
and U348 (N_348,N_251,N_230);
nand U349 (N_349,N_216,N_222);
nand U350 (N_350,N_273,N_210);
xnor U351 (N_351,In_331,N_180);
and U352 (N_352,N_141,N_267);
xnor U353 (N_353,In_300,In_183);
nor U354 (N_354,In_149,N_6);
or U355 (N_355,N_276,N_126);
xnor U356 (N_356,In_31,N_235);
or U357 (N_357,N_101,In_2);
and U358 (N_358,In_237,N_266);
nor U359 (N_359,N_294,In_199);
nor U360 (N_360,N_259,N_207);
or U361 (N_361,N_237,N_250);
or U362 (N_362,N_98,N_159);
and U363 (N_363,In_472,N_129);
and U364 (N_364,N_275,In_188);
nor U365 (N_365,N_103,N_135);
and U366 (N_366,In_442,N_224);
nand U367 (N_367,N_288,N_234);
nand U368 (N_368,N_11,In_409);
nand U369 (N_369,N_265,N_247);
and U370 (N_370,N_260,N_268);
xnor U371 (N_371,N_286,N_213);
xor U372 (N_372,In_103,N_236);
nand U373 (N_373,In_447,N_254);
or U374 (N_374,N_245,N_214);
or U375 (N_375,In_458,N_27);
and U376 (N_376,N_298,N_166);
and U377 (N_377,N_106,N_229);
xor U378 (N_378,N_281,N_122);
or U379 (N_379,N_134,In_3);
nor U380 (N_380,N_280,N_39);
or U381 (N_381,N_179,In_491);
or U382 (N_382,N_232,N_231);
xnor U383 (N_383,N_277,In_338);
and U384 (N_384,N_175,N_255);
and U385 (N_385,N_282,N_187);
and U386 (N_386,In_145,In_94);
and U387 (N_387,N_261,N_217);
and U388 (N_388,In_425,N_221);
and U389 (N_389,In_303,In_48);
and U390 (N_390,N_215,N_81);
and U391 (N_391,N_253,N_160);
and U392 (N_392,In_340,N_212);
xnor U393 (N_393,N_204,N_228);
nand U394 (N_394,In_119,In_147);
or U395 (N_395,N_270,In_72);
or U396 (N_396,N_297,N_283);
or U397 (N_397,N_79,N_194);
or U398 (N_398,N_289,N_109);
and U399 (N_399,N_258,In_449);
or U400 (N_400,N_378,N_316);
nand U401 (N_401,N_357,N_368);
or U402 (N_402,N_315,N_373);
xor U403 (N_403,N_397,N_348);
and U404 (N_404,N_372,N_389);
nand U405 (N_405,N_331,N_353);
nand U406 (N_406,N_355,N_328);
or U407 (N_407,N_323,N_342);
and U408 (N_408,N_314,N_377);
nand U409 (N_409,N_335,N_366);
nand U410 (N_410,N_394,N_392);
nand U411 (N_411,N_300,N_362);
nand U412 (N_412,N_303,N_320);
nand U413 (N_413,N_390,N_336);
nor U414 (N_414,N_395,N_363);
and U415 (N_415,N_358,N_319);
and U416 (N_416,N_325,N_384);
nand U417 (N_417,N_396,N_354);
nor U418 (N_418,N_371,N_385);
nor U419 (N_419,N_334,N_318);
and U420 (N_420,N_326,N_379);
or U421 (N_421,N_332,N_351);
nand U422 (N_422,N_317,N_337);
and U423 (N_423,N_344,N_322);
and U424 (N_424,N_398,N_321);
nand U425 (N_425,N_393,N_347);
or U426 (N_426,N_391,N_307);
xnor U427 (N_427,N_329,N_330);
and U428 (N_428,N_369,N_356);
and U429 (N_429,N_361,N_375);
or U430 (N_430,N_399,N_388);
or U431 (N_431,N_327,N_360);
or U432 (N_432,N_381,N_309);
or U433 (N_433,N_341,N_349);
nor U434 (N_434,N_370,N_346);
nand U435 (N_435,N_308,N_310);
or U436 (N_436,N_306,N_339);
or U437 (N_437,N_350,N_313);
nand U438 (N_438,N_345,N_305);
or U439 (N_439,N_359,N_364);
and U440 (N_440,N_311,N_340);
nor U441 (N_441,N_301,N_324);
and U442 (N_442,N_365,N_374);
or U443 (N_443,N_343,N_383);
nand U444 (N_444,N_338,N_367);
nand U445 (N_445,N_380,N_382);
nor U446 (N_446,N_312,N_304);
nand U447 (N_447,N_386,N_302);
and U448 (N_448,N_352,N_376);
nand U449 (N_449,N_333,N_387);
nor U450 (N_450,N_368,N_352);
nor U451 (N_451,N_364,N_346);
and U452 (N_452,N_359,N_350);
and U453 (N_453,N_325,N_301);
nand U454 (N_454,N_323,N_343);
or U455 (N_455,N_343,N_308);
xor U456 (N_456,N_307,N_397);
and U457 (N_457,N_370,N_313);
nor U458 (N_458,N_390,N_317);
nor U459 (N_459,N_301,N_305);
nand U460 (N_460,N_301,N_399);
nand U461 (N_461,N_350,N_315);
and U462 (N_462,N_361,N_317);
or U463 (N_463,N_317,N_364);
or U464 (N_464,N_369,N_310);
xnor U465 (N_465,N_392,N_358);
and U466 (N_466,N_336,N_333);
nor U467 (N_467,N_341,N_301);
nor U468 (N_468,N_314,N_330);
xnor U469 (N_469,N_351,N_334);
or U470 (N_470,N_336,N_357);
or U471 (N_471,N_346,N_313);
or U472 (N_472,N_340,N_320);
or U473 (N_473,N_314,N_343);
nand U474 (N_474,N_390,N_323);
and U475 (N_475,N_310,N_331);
or U476 (N_476,N_333,N_337);
nor U477 (N_477,N_315,N_303);
or U478 (N_478,N_324,N_396);
nand U479 (N_479,N_321,N_358);
and U480 (N_480,N_352,N_313);
nand U481 (N_481,N_397,N_374);
and U482 (N_482,N_353,N_321);
and U483 (N_483,N_356,N_362);
xnor U484 (N_484,N_383,N_361);
nand U485 (N_485,N_352,N_367);
and U486 (N_486,N_301,N_316);
or U487 (N_487,N_385,N_352);
or U488 (N_488,N_340,N_309);
nand U489 (N_489,N_382,N_365);
nand U490 (N_490,N_368,N_305);
and U491 (N_491,N_389,N_358);
or U492 (N_492,N_302,N_319);
or U493 (N_493,N_393,N_350);
and U494 (N_494,N_358,N_345);
or U495 (N_495,N_374,N_391);
nand U496 (N_496,N_340,N_355);
nand U497 (N_497,N_322,N_327);
nand U498 (N_498,N_376,N_390);
nand U499 (N_499,N_350,N_306);
and U500 (N_500,N_414,N_491);
and U501 (N_501,N_452,N_499);
nand U502 (N_502,N_442,N_494);
or U503 (N_503,N_453,N_446);
nor U504 (N_504,N_487,N_488);
nor U505 (N_505,N_416,N_431);
or U506 (N_506,N_461,N_405);
xnor U507 (N_507,N_425,N_400);
nand U508 (N_508,N_423,N_426);
nand U509 (N_509,N_479,N_404);
or U510 (N_510,N_433,N_458);
and U511 (N_511,N_412,N_489);
and U512 (N_512,N_401,N_480);
and U513 (N_513,N_485,N_474);
nor U514 (N_514,N_432,N_444);
nand U515 (N_515,N_427,N_477);
nor U516 (N_516,N_492,N_424);
xor U517 (N_517,N_435,N_450);
nor U518 (N_518,N_418,N_476);
and U519 (N_519,N_472,N_436);
and U520 (N_520,N_451,N_484);
and U521 (N_521,N_430,N_454);
xor U522 (N_522,N_441,N_403);
xnor U523 (N_523,N_448,N_496);
nand U524 (N_524,N_420,N_408);
or U525 (N_525,N_490,N_498);
or U526 (N_526,N_466,N_459);
nor U527 (N_527,N_402,N_464);
nor U528 (N_528,N_456,N_468);
and U529 (N_529,N_478,N_439);
and U530 (N_530,N_440,N_481);
nand U531 (N_531,N_419,N_473);
xnor U532 (N_532,N_429,N_469);
xor U533 (N_533,N_475,N_471);
and U534 (N_534,N_437,N_443);
nor U535 (N_535,N_438,N_413);
xor U536 (N_536,N_455,N_465);
or U537 (N_537,N_410,N_409);
and U538 (N_538,N_407,N_495);
xor U539 (N_539,N_462,N_449);
or U540 (N_540,N_415,N_457);
nor U541 (N_541,N_470,N_421);
or U542 (N_542,N_460,N_493);
nor U543 (N_543,N_445,N_497);
xor U544 (N_544,N_482,N_422);
nor U545 (N_545,N_447,N_463);
xnor U546 (N_546,N_417,N_428);
and U547 (N_547,N_434,N_483);
xnor U548 (N_548,N_486,N_411);
and U549 (N_549,N_406,N_467);
and U550 (N_550,N_463,N_489);
nand U551 (N_551,N_408,N_405);
or U552 (N_552,N_418,N_469);
nor U553 (N_553,N_481,N_483);
and U554 (N_554,N_497,N_440);
xnor U555 (N_555,N_483,N_445);
nor U556 (N_556,N_425,N_462);
nand U557 (N_557,N_470,N_451);
xnor U558 (N_558,N_440,N_457);
or U559 (N_559,N_489,N_417);
xnor U560 (N_560,N_453,N_431);
nand U561 (N_561,N_461,N_471);
nand U562 (N_562,N_443,N_420);
and U563 (N_563,N_423,N_460);
or U564 (N_564,N_487,N_421);
nand U565 (N_565,N_403,N_490);
nor U566 (N_566,N_469,N_432);
or U567 (N_567,N_482,N_481);
nand U568 (N_568,N_498,N_404);
or U569 (N_569,N_420,N_428);
and U570 (N_570,N_461,N_463);
and U571 (N_571,N_457,N_404);
nor U572 (N_572,N_476,N_498);
and U573 (N_573,N_435,N_484);
or U574 (N_574,N_429,N_459);
xor U575 (N_575,N_487,N_484);
xnor U576 (N_576,N_495,N_485);
and U577 (N_577,N_457,N_430);
xnor U578 (N_578,N_413,N_441);
nor U579 (N_579,N_409,N_433);
nand U580 (N_580,N_456,N_466);
or U581 (N_581,N_487,N_409);
and U582 (N_582,N_482,N_437);
nor U583 (N_583,N_452,N_425);
nor U584 (N_584,N_462,N_488);
or U585 (N_585,N_452,N_434);
nor U586 (N_586,N_428,N_449);
and U587 (N_587,N_444,N_497);
and U588 (N_588,N_415,N_459);
nand U589 (N_589,N_482,N_406);
and U590 (N_590,N_406,N_483);
nor U591 (N_591,N_411,N_449);
nand U592 (N_592,N_472,N_462);
nor U593 (N_593,N_438,N_410);
nor U594 (N_594,N_464,N_450);
or U595 (N_595,N_406,N_457);
nand U596 (N_596,N_403,N_401);
or U597 (N_597,N_404,N_474);
or U598 (N_598,N_414,N_476);
nand U599 (N_599,N_467,N_466);
nand U600 (N_600,N_599,N_529);
nor U601 (N_601,N_512,N_541);
and U602 (N_602,N_576,N_506);
nand U603 (N_603,N_582,N_536);
xnor U604 (N_604,N_550,N_554);
and U605 (N_605,N_508,N_527);
nor U606 (N_606,N_570,N_589);
xor U607 (N_607,N_533,N_588);
nand U608 (N_608,N_517,N_551);
or U609 (N_609,N_538,N_542);
nand U610 (N_610,N_522,N_586);
and U611 (N_611,N_520,N_592);
xnor U612 (N_612,N_540,N_525);
xor U613 (N_613,N_584,N_562);
nand U614 (N_614,N_552,N_503);
nand U615 (N_615,N_545,N_534);
nor U616 (N_616,N_524,N_532);
and U617 (N_617,N_537,N_531);
nand U618 (N_618,N_567,N_514);
nor U619 (N_619,N_528,N_546);
or U620 (N_620,N_574,N_511);
and U621 (N_621,N_593,N_501);
nand U622 (N_622,N_543,N_547);
nor U623 (N_623,N_580,N_504);
and U624 (N_624,N_594,N_523);
and U625 (N_625,N_569,N_558);
nand U626 (N_626,N_565,N_507);
and U627 (N_627,N_509,N_577);
xnor U628 (N_628,N_557,N_505);
nor U629 (N_629,N_559,N_564);
and U630 (N_630,N_515,N_587);
nand U631 (N_631,N_585,N_573);
and U632 (N_632,N_560,N_553);
and U633 (N_633,N_518,N_563);
and U634 (N_634,N_596,N_578);
or U635 (N_635,N_575,N_549);
nand U636 (N_636,N_566,N_571);
or U637 (N_637,N_595,N_544);
nor U638 (N_638,N_572,N_583);
or U639 (N_639,N_535,N_590);
or U640 (N_640,N_526,N_516);
or U641 (N_641,N_568,N_502);
or U642 (N_642,N_521,N_500);
or U643 (N_643,N_539,N_561);
or U644 (N_644,N_513,N_581);
nor U645 (N_645,N_555,N_510);
and U646 (N_646,N_598,N_597);
and U647 (N_647,N_591,N_548);
nand U648 (N_648,N_579,N_519);
xor U649 (N_649,N_556,N_530);
and U650 (N_650,N_561,N_595);
nand U651 (N_651,N_583,N_511);
and U652 (N_652,N_574,N_597);
nor U653 (N_653,N_583,N_551);
or U654 (N_654,N_557,N_546);
nand U655 (N_655,N_544,N_557);
or U656 (N_656,N_577,N_531);
or U657 (N_657,N_512,N_558);
nand U658 (N_658,N_596,N_590);
nor U659 (N_659,N_528,N_515);
and U660 (N_660,N_528,N_552);
and U661 (N_661,N_570,N_549);
or U662 (N_662,N_502,N_508);
and U663 (N_663,N_570,N_511);
and U664 (N_664,N_599,N_584);
nand U665 (N_665,N_572,N_585);
nor U666 (N_666,N_550,N_542);
nand U667 (N_667,N_513,N_524);
or U668 (N_668,N_504,N_523);
nand U669 (N_669,N_513,N_573);
or U670 (N_670,N_578,N_544);
or U671 (N_671,N_558,N_533);
xnor U672 (N_672,N_598,N_536);
and U673 (N_673,N_576,N_584);
nand U674 (N_674,N_585,N_581);
or U675 (N_675,N_507,N_560);
nand U676 (N_676,N_561,N_503);
xor U677 (N_677,N_574,N_509);
or U678 (N_678,N_586,N_504);
or U679 (N_679,N_527,N_589);
and U680 (N_680,N_536,N_554);
and U681 (N_681,N_501,N_597);
nand U682 (N_682,N_520,N_562);
or U683 (N_683,N_520,N_505);
xnor U684 (N_684,N_518,N_581);
nor U685 (N_685,N_577,N_521);
or U686 (N_686,N_522,N_545);
and U687 (N_687,N_530,N_599);
nand U688 (N_688,N_551,N_570);
or U689 (N_689,N_571,N_524);
nand U690 (N_690,N_561,N_547);
or U691 (N_691,N_515,N_589);
and U692 (N_692,N_548,N_593);
and U693 (N_693,N_579,N_597);
and U694 (N_694,N_530,N_550);
nor U695 (N_695,N_531,N_553);
nand U696 (N_696,N_517,N_557);
and U697 (N_697,N_525,N_584);
xor U698 (N_698,N_578,N_511);
and U699 (N_699,N_587,N_594);
nor U700 (N_700,N_613,N_659);
xor U701 (N_701,N_642,N_697);
nor U702 (N_702,N_631,N_672);
nor U703 (N_703,N_682,N_621);
nor U704 (N_704,N_662,N_634);
nand U705 (N_705,N_615,N_666);
or U706 (N_706,N_687,N_626);
nor U707 (N_707,N_646,N_679);
and U708 (N_708,N_683,N_636);
nand U709 (N_709,N_618,N_614);
nand U710 (N_710,N_698,N_675);
nand U711 (N_711,N_653,N_689);
or U712 (N_712,N_640,N_685);
and U713 (N_713,N_654,N_665);
nand U714 (N_714,N_610,N_620);
nand U715 (N_715,N_612,N_644);
nor U716 (N_716,N_651,N_605);
or U717 (N_717,N_600,N_686);
or U718 (N_718,N_652,N_629);
nand U719 (N_719,N_643,N_630);
and U720 (N_720,N_656,N_657);
or U721 (N_721,N_678,N_695);
and U722 (N_722,N_668,N_649);
and U723 (N_723,N_645,N_641);
and U724 (N_724,N_628,N_676);
or U725 (N_725,N_633,N_655);
nor U726 (N_726,N_663,N_609);
nand U727 (N_727,N_699,N_602);
or U728 (N_728,N_660,N_635);
nor U729 (N_729,N_670,N_650);
and U730 (N_730,N_611,N_625);
or U731 (N_731,N_608,N_658);
or U732 (N_732,N_604,N_677);
nand U733 (N_733,N_693,N_601);
or U734 (N_734,N_638,N_661);
or U735 (N_735,N_688,N_624);
and U736 (N_736,N_632,N_684);
nor U737 (N_737,N_606,N_664);
nor U738 (N_738,N_681,N_674);
or U739 (N_739,N_667,N_671);
and U740 (N_740,N_680,N_648);
nor U741 (N_741,N_692,N_622);
and U742 (N_742,N_696,N_607);
nand U743 (N_743,N_647,N_639);
nand U744 (N_744,N_627,N_694);
nor U745 (N_745,N_690,N_603);
nor U746 (N_746,N_616,N_617);
and U747 (N_747,N_669,N_623);
nor U748 (N_748,N_619,N_673);
xnor U749 (N_749,N_637,N_691);
nand U750 (N_750,N_629,N_628);
and U751 (N_751,N_683,N_668);
nand U752 (N_752,N_655,N_690);
nor U753 (N_753,N_625,N_691);
xor U754 (N_754,N_697,N_644);
or U755 (N_755,N_652,N_656);
or U756 (N_756,N_666,N_632);
nand U757 (N_757,N_621,N_679);
nor U758 (N_758,N_691,N_603);
and U759 (N_759,N_609,N_629);
or U760 (N_760,N_639,N_675);
nor U761 (N_761,N_662,N_620);
xnor U762 (N_762,N_637,N_625);
or U763 (N_763,N_648,N_604);
nor U764 (N_764,N_698,N_603);
or U765 (N_765,N_684,N_680);
nor U766 (N_766,N_636,N_689);
and U767 (N_767,N_664,N_601);
and U768 (N_768,N_612,N_610);
and U769 (N_769,N_689,N_664);
or U770 (N_770,N_698,N_627);
or U771 (N_771,N_626,N_696);
xnor U772 (N_772,N_622,N_634);
nor U773 (N_773,N_612,N_624);
nor U774 (N_774,N_645,N_691);
nand U775 (N_775,N_624,N_678);
xor U776 (N_776,N_602,N_631);
or U777 (N_777,N_680,N_695);
and U778 (N_778,N_652,N_603);
nor U779 (N_779,N_657,N_691);
nand U780 (N_780,N_607,N_642);
nand U781 (N_781,N_669,N_683);
nor U782 (N_782,N_692,N_601);
and U783 (N_783,N_600,N_672);
and U784 (N_784,N_676,N_652);
nor U785 (N_785,N_634,N_686);
nand U786 (N_786,N_668,N_689);
nand U787 (N_787,N_691,N_614);
or U788 (N_788,N_652,N_638);
nand U789 (N_789,N_643,N_636);
or U790 (N_790,N_646,N_697);
xnor U791 (N_791,N_614,N_688);
nand U792 (N_792,N_649,N_689);
and U793 (N_793,N_652,N_690);
or U794 (N_794,N_681,N_644);
or U795 (N_795,N_641,N_692);
and U796 (N_796,N_640,N_649);
nand U797 (N_797,N_610,N_664);
nand U798 (N_798,N_665,N_600);
nand U799 (N_799,N_663,N_645);
nor U800 (N_800,N_798,N_736);
or U801 (N_801,N_785,N_759);
xor U802 (N_802,N_766,N_741);
nor U803 (N_803,N_744,N_796);
nand U804 (N_804,N_762,N_795);
and U805 (N_805,N_764,N_777);
xnor U806 (N_806,N_725,N_786);
or U807 (N_807,N_730,N_780);
nand U808 (N_808,N_720,N_756);
or U809 (N_809,N_700,N_753);
and U810 (N_810,N_746,N_738);
or U811 (N_811,N_767,N_757);
xor U812 (N_812,N_717,N_721);
and U813 (N_813,N_747,N_772);
nand U814 (N_814,N_771,N_793);
nor U815 (N_815,N_731,N_770);
or U816 (N_816,N_781,N_728);
and U817 (N_817,N_775,N_713);
and U818 (N_818,N_740,N_705);
nor U819 (N_819,N_787,N_712);
or U820 (N_820,N_763,N_776);
or U821 (N_821,N_751,N_718);
or U822 (N_822,N_714,N_733);
nand U823 (N_823,N_743,N_749);
and U824 (N_824,N_742,N_709);
or U825 (N_825,N_761,N_719);
nand U826 (N_826,N_782,N_748);
nor U827 (N_827,N_703,N_745);
or U828 (N_828,N_735,N_768);
and U829 (N_829,N_789,N_790);
nor U830 (N_830,N_722,N_704);
nor U831 (N_831,N_773,N_797);
and U832 (N_832,N_702,N_729);
or U833 (N_833,N_755,N_774);
and U834 (N_834,N_708,N_732);
and U835 (N_835,N_727,N_724);
and U836 (N_836,N_715,N_750);
nor U837 (N_837,N_706,N_760);
and U838 (N_838,N_778,N_783);
and U839 (N_839,N_726,N_752);
and U840 (N_840,N_737,N_799);
nor U841 (N_841,N_784,N_711);
nor U842 (N_842,N_723,N_769);
xor U843 (N_843,N_788,N_791);
and U844 (N_844,N_754,N_734);
nor U845 (N_845,N_701,N_716);
or U846 (N_846,N_792,N_779);
or U847 (N_847,N_739,N_794);
and U848 (N_848,N_758,N_765);
and U849 (N_849,N_710,N_707);
xor U850 (N_850,N_728,N_751);
and U851 (N_851,N_713,N_739);
or U852 (N_852,N_786,N_799);
or U853 (N_853,N_793,N_749);
nand U854 (N_854,N_769,N_789);
nor U855 (N_855,N_781,N_798);
xnor U856 (N_856,N_790,N_702);
and U857 (N_857,N_752,N_741);
nor U858 (N_858,N_761,N_799);
or U859 (N_859,N_780,N_729);
and U860 (N_860,N_757,N_768);
nand U861 (N_861,N_754,N_776);
or U862 (N_862,N_771,N_743);
and U863 (N_863,N_767,N_766);
nor U864 (N_864,N_756,N_707);
nand U865 (N_865,N_755,N_747);
nand U866 (N_866,N_753,N_799);
nor U867 (N_867,N_720,N_757);
nor U868 (N_868,N_762,N_711);
nand U869 (N_869,N_734,N_704);
and U870 (N_870,N_785,N_789);
and U871 (N_871,N_724,N_721);
and U872 (N_872,N_759,N_712);
or U873 (N_873,N_757,N_791);
nor U874 (N_874,N_761,N_743);
or U875 (N_875,N_752,N_772);
nand U876 (N_876,N_774,N_720);
or U877 (N_877,N_784,N_772);
nor U878 (N_878,N_737,N_768);
and U879 (N_879,N_759,N_772);
nor U880 (N_880,N_741,N_789);
and U881 (N_881,N_703,N_748);
nand U882 (N_882,N_731,N_723);
or U883 (N_883,N_750,N_704);
nand U884 (N_884,N_702,N_737);
or U885 (N_885,N_762,N_742);
nand U886 (N_886,N_747,N_730);
nor U887 (N_887,N_761,N_720);
or U888 (N_888,N_759,N_711);
nor U889 (N_889,N_748,N_770);
or U890 (N_890,N_748,N_717);
and U891 (N_891,N_799,N_764);
or U892 (N_892,N_787,N_753);
nor U893 (N_893,N_761,N_739);
nand U894 (N_894,N_710,N_729);
or U895 (N_895,N_767,N_761);
nor U896 (N_896,N_737,N_731);
nand U897 (N_897,N_703,N_733);
nor U898 (N_898,N_749,N_737);
nand U899 (N_899,N_740,N_791);
or U900 (N_900,N_848,N_842);
or U901 (N_901,N_851,N_865);
nand U902 (N_902,N_819,N_801);
nor U903 (N_903,N_896,N_859);
nor U904 (N_904,N_890,N_856);
and U905 (N_905,N_818,N_826);
nor U906 (N_906,N_878,N_824);
nand U907 (N_907,N_853,N_832);
or U908 (N_908,N_855,N_829);
nand U909 (N_909,N_807,N_893);
nor U910 (N_910,N_870,N_879);
and U911 (N_911,N_882,N_877);
or U912 (N_912,N_831,N_871);
nand U913 (N_913,N_835,N_872);
nor U914 (N_914,N_899,N_845);
xnor U915 (N_915,N_843,N_867);
or U916 (N_916,N_825,N_897);
or U917 (N_917,N_822,N_874);
and U918 (N_918,N_813,N_892);
nand U919 (N_919,N_849,N_861);
and U920 (N_920,N_894,N_886);
or U921 (N_921,N_891,N_802);
nand U922 (N_922,N_800,N_866);
and U923 (N_923,N_852,N_815);
and U924 (N_924,N_895,N_828);
and U925 (N_925,N_805,N_838);
or U926 (N_926,N_884,N_830);
or U927 (N_927,N_810,N_880);
nand U928 (N_928,N_883,N_841);
or U929 (N_929,N_812,N_876);
xnor U930 (N_930,N_834,N_806);
or U931 (N_931,N_857,N_823);
nand U932 (N_932,N_881,N_814);
and U933 (N_933,N_804,N_833);
or U934 (N_934,N_858,N_817);
or U935 (N_935,N_863,N_811);
or U936 (N_936,N_898,N_887);
nand U937 (N_937,N_808,N_844);
or U938 (N_938,N_840,N_827);
nand U939 (N_939,N_869,N_850);
and U940 (N_940,N_875,N_847);
or U941 (N_941,N_854,N_809);
and U942 (N_942,N_846,N_885);
nand U943 (N_943,N_873,N_888);
and U944 (N_944,N_837,N_862);
nand U945 (N_945,N_821,N_839);
nor U946 (N_946,N_889,N_803);
or U947 (N_947,N_816,N_836);
xor U948 (N_948,N_864,N_820);
nand U949 (N_949,N_860,N_868);
nor U950 (N_950,N_888,N_874);
or U951 (N_951,N_899,N_878);
nor U952 (N_952,N_838,N_872);
or U953 (N_953,N_875,N_878);
nor U954 (N_954,N_855,N_857);
and U955 (N_955,N_899,N_818);
or U956 (N_956,N_887,N_881);
xor U957 (N_957,N_826,N_814);
nand U958 (N_958,N_800,N_855);
nand U959 (N_959,N_818,N_858);
and U960 (N_960,N_810,N_820);
nand U961 (N_961,N_879,N_835);
nand U962 (N_962,N_850,N_830);
or U963 (N_963,N_886,N_811);
nor U964 (N_964,N_848,N_879);
or U965 (N_965,N_833,N_875);
nor U966 (N_966,N_893,N_806);
or U967 (N_967,N_822,N_863);
nor U968 (N_968,N_813,N_845);
xnor U969 (N_969,N_800,N_872);
and U970 (N_970,N_805,N_879);
xor U971 (N_971,N_839,N_891);
nand U972 (N_972,N_854,N_865);
nor U973 (N_973,N_840,N_800);
nor U974 (N_974,N_873,N_823);
nor U975 (N_975,N_890,N_810);
or U976 (N_976,N_892,N_805);
xnor U977 (N_977,N_867,N_825);
nor U978 (N_978,N_866,N_869);
nand U979 (N_979,N_853,N_877);
and U980 (N_980,N_814,N_893);
and U981 (N_981,N_815,N_849);
nand U982 (N_982,N_848,N_808);
nor U983 (N_983,N_850,N_870);
nor U984 (N_984,N_837,N_850);
xor U985 (N_985,N_822,N_895);
nand U986 (N_986,N_833,N_816);
nor U987 (N_987,N_806,N_873);
xnor U988 (N_988,N_846,N_840);
and U989 (N_989,N_837,N_830);
or U990 (N_990,N_810,N_896);
and U991 (N_991,N_806,N_867);
and U992 (N_992,N_852,N_803);
or U993 (N_993,N_864,N_811);
or U994 (N_994,N_851,N_874);
nor U995 (N_995,N_807,N_880);
nand U996 (N_996,N_870,N_818);
nor U997 (N_997,N_848,N_837);
and U998 (N_998,N_839,N_813);
nand U999 (N_999,N_834,N_821);
and U1000 (N_1000,N_949,N_958);
nand U1001 (N_1001,N_935,N_918);
or U1002 (N_1002,N_926,N_960);
and U1003 (N_1003,N_910,N_920);
or U1004 (N_1004,N_955,N_996);
or U1005 (N_1005,N_952,N_993);
nor U1006 (N_1006,N_948,N_900);
nand U1007 (N_1007,N_959,N_997);
or U1008 (N_1008,N_947,N_976);
nand U1009 (N_1009,N_939,N_984);
and U1010 (N_1010,N_905,N_930);
nand U1011 (N_1011,N_956,N_967);
nand U1012 (N_1012,N_973,N_912);
nand U1013 (N_1013,N_914,N_940);
xor U1014 (N_1014,N_980,N_901);
and U1015 (N_1015,N_992,N_968);
or U1016 (N_1016,N_927,N_915);
nor U1017 (N_1017,N_921,N_990);
or U1018 (N_1018,N_931,N_975);
nand U1019 (N_1019,N_928,N_964);
xor U1020 (N_1020,N_936,N_953);
nand U1021 (N_1021,N_961,N_986);
xor U1022 (N_1022,N_954,N_978);
nand U1023 (N_1023,N_962,N_944);
nor U1024 (N_1024,N_904,N_902);
or U1025 (N_1025,N_929,N_938);
and U1026 (N_1026,N_969,N_945);
nand U1027 (N_1027,N_977,N_989);
or U1028 (N_1028,N_922,N_923);
or U1029 (N_1029,N_942,N_908);
nor U1030 (N_1030,N_924,N_972);
nor U1031 (N_1031,N_937,N_983);
nor U1032 (N_1032,N_979,N_965);
nand U1033 (N_1033,N_995,N_932);
nand U1034 (N_1034,N_950,N_966);
or U1035 (N_1035,N_916,N_951);
nand U1036 (N_1036,N_919,N_913);
and U1037 (N_1037,N_987,N_946);
xor U1038 (N_1038,N_925,N_971);
nand U1039 (N_1039,N_985,N_907);
or U1040 (N_1040,N_933,N_998);
nor U1041 (N_1041,N_934,N_909);
and U1042 (N_1042,N_906,N_988);
or U1043 (N_1043,N_974,N_943);
nand U1044 (N_1044,N_982,N_999);
and U1045 (N_1045,N_991,N_903);
nor U1046 (N_1046,N_911,N_970);
xnor U1047 (N_1047,N_994,N_941);
nand U1048 (N_1048,N_917,N_981);
nor U1049 (N_1049,N_963,N_957);
or U1050 (N_1050,N_973,N_958);
and U1051 (N_1051,N_979,N_983);
nand U1052 (N_1052,N_988,N_920);
nand U1053 (N_1053,N_900,N_931);
or U1054 (N_1054,N_970,N_951);
or U1055 (N_1055,N_992,N_950);
nor U1056 (N_1056,N_960,N_937);
nand U1057 (N_1057,N_953,N_992);
or U1058 (N_1058,N_982,N_953);
nor U1059 (N_1059,N_944,N_918);
xnor U1060 (N_1060,N_957,N_978);
nand U1061 (N_1061,N_967,N_915);
nand U1062 (N_1062,N_999,N_994);
and U1063 (N_1063,N_917,N_992);
or U1064 (N_1064,N_958,N_994);
nor U1065 (N_1065,N_916,N_997);
or U1066 (N_1066,N_966,N_989);
nand U1067 (N_1067,N_995,N_946);
xnor U1068 (N_1068,N_944,N_942);
nor U1069 (N_1069,N_989,N_988);
or U1070 (N_1070,N_968,N_931);
nor U1071 (N_1071,N_934,N_978);
nand U1072 (N_1072,N_945,N_928);
xnor U1073 (N_1073,N_918,N_967);
nor U1074 (N_1074,N_981,N_973);
and U1075 (N_1075,N_985,N_972);
or U1076 (N_1076,N_916,N_966);
nand U1077 (N_1077,N_924,N_952);
xnor U1078 (N_1078,N_928,N_960);
or U1079 (N_1079,N_935,N_931);
nand U1080 (N_1080,N_978,N_982);
xor U1081 (N_1081,N_949,N_971);
or U1082 (N_1082,N_933,N_922);
or U1083 (N_1083,N_938,N_936);
nor U1084 (N_1084,N_985,N_997);
xor U1085 (N_1085,N_913,N_997);
nand U1086 (N_1086,N_966,N_978);
nor U1087 (N_1087,N_949,N_900);
and U1088 (N_1088,N_953,N_931);
nor U1089 (N_1089,N_902,N_948);
nor U1090 (N_1090,N_973,N_972);
or U1091 (N_1091,N_960,N_955);
nor U1092 (N_1092,N_986,N_971);
nand U1093 (N_1093,N_991,N_921);
xor U1094 (N_1094,N_990,N_935);
or U1095 (N_1095,N_907,N_992);
nor U1096 (N_1096,N_916,N_939);
xnor U1097 (N_1097,N_937,N_902);
or U1098 (N_1098,N_969,N_982);
nand U1099 (N_1099,N_990,N_925);
nand U1100 (N_1100,N_1035,N_1082);
nand U1101 (N_1101,N_1018,N_1086);
or U1102 (N_1102,N_1005,N_1007);
xnor U1103 (N_1103,N_1092,N_1069);
and U1104 (N_1104,N_1078,N_1034);
and U1105 (N_1105,N_1004,N_1029);
or U1106 (N_1106,N_1085,N_1000);
nand U1107 (N_1107,N_1063,N_1015);
nor U1108 (N_1108,N_1033,N_1026);
nor U1109 (N_1109,N_1023,N_1070);
nand U1110 (N_1110,N_1050,N_1001);
or U1111 (N_1111,N_1012,N_1030);
and U1112 (N_1112,N_1073,N_1055);
or U1113 (N_1113,N_1036,N_1087);
or U1114 (N_1114,N_1088,N_1040);
nor U1115 (N_1115,N_1008,N_1095);
xnor U1116 (N_1116,N_1049,N_1083);
or U1117 (N_1117,N_1051,N_1039);
or U1118 (N_1118,N_1080,N_1081);
nand U1119 (N_1119,N_1038,N_1027);
nor U1120 (N_1120,N_1098,N_1075);
xnor U1121 (N_1121,N_1061,N_1071);
or U1122 (N_1122,N_1043,N_1028);
or U1123 (N_1123,N_1062,N_1094);
nand U1124 (N_1124,N_1019,N_1089);
xor U1125 (N_1125,N_1003,N_1017);
or U1126 (N_1126,N_1074,N_1065);
nand U1127 (N_1127,N_1064,N_1099);
and U1128 (N_1128,N_1054,N_1041);
or U1129 (N_1129,N_1068,N_1010);
nand U1130 (N_1130,N_1076,N_1024);
nor U1131 (N_1131,N_1009,N_1058);
and U1132 (N_1132,N_1025,N_1084);
nor U1133 (N_1133,N_1090,N_1013);
and U1134 (N_1134,N_1011,N_1021);
and U1135 (N_1135,N_1002,N_1067);
nand U1136 (N_1136,N_1044,N_1056);
or U1137 (N_1137,N_1006,N_1066);
or U1138 (N_1138,N_1020,N_1047);
and U1139 (N_1139,N_1091,N_1072);
nand U1140 (N_1140,N_1096,N_1052);
xnor U1141 (N_1141,N_1014,N_1048);
nor U1142 (N_1142,N_1077,N_1045);
and U1143 (N_1143,N_1097,N_1032);
nand U1144 (N_1144,N_1060,N_1093);
xor U1145 (N_1145,N_1031,N_1016);
xnor U1146 (N_1146,N_1053,N_1046);
or U1147 (N_1147,N_1037,N_1057);
nand U1148 (N_1148,N_1059,N_1022);
nor U1149 (N_1149,N_1042,N_1079);
and U1150 (N_1150,N_1024,N_1063);
and U1151 (N_1151,N_1048,N_1001);
or U1152 (N_1152,N_1025,N_1074);
nand U1153 (N_1153,N_1042,N_1000);
nand U1154 (N_1154,N_1058,N_1071);
and U1155 (N_1155,N_1001,N_1017);
and U1156 (N_1156,N_1009,N_1069);
and U1157 (N_1157,N_1042,N_1067);
nor U1158 (N_1158,N_1002,N_1061);
xor U1159 (N_1159,N_1045,N_1086);
nand U1160 (N_1160,N_1099,N_1079);
xnor U1161 (N_1161,N_1006,N_1083);
nand U1162 (N_1162,N_1063,N_1023);
nand U1163 (N_1163,N_1053,N_1060);
nor U1164 (N_1164,N_1013,N_1068);
nand U1165 (N_1165,N_1060,N_1085);
nand U1166 (N_1166,N_1056,N_1092);
xor U1167 (N_1167,N_1020,N_1001);
xnor U1168 (N_1168,N_1010,N_1065);
nor U1169 (N_1169,N_1047,N_1042);
nor U1170 (N_1170,N_1062,N_1079);
or U1171 (N_1171,N_1048,N_1053);
or U1172 (N_1172,N_1038,N_1069);
nand U1173 (N_1173,N_1040,N_1003);
and U1174 (N_1174,N_1001,N_1098);
xor U1175 (N_1175,N_1017,N_1063);
nor U1176 (N_1176,N_1019,N_1039);
nand U1177 (N_1177,N_1054,N_1046);
nor U1178 (N_1178,N_1073,N_1039);
nor U1179 (N_1179,N_1063,N_1061);
xor U1180 (N_1180,N_1042,N_1053);
xnor U1181 (N_1181,N_1037,N_1019);
and U1182 (N_1182,N_1094,N_1059);
nor U1183 (N_1183,N_1007,N_1048);
or U1184 (N_1184,N_1082,N_1069);
xor U1185 (N_1185,N_1056,N_1091);
and U1186 (N_1186,N_1015,N_1098);
nor U1187 (N_1187,N_1047,N_1021);
nand U1188 (N_1188,N_1089,N_1016);
xor U1189 (N_1189,N_1092,N_1052);
nand U1190 (N_1190,N_1057,N_1055);
nor U1191 (N_1191,N_1087,N_1062);
and U1192 (N_1192,N_1074,N_1051);
nor U1193 (N_1193,N_1089,N_1009);
and U1194 (N_1194,N_1012,N_1070);
and U1195 (N_1195,N_1097,N_1017);
and U1196 (N_1196,N_1039,N_1016);
or U1197 (N_1197,N_1031,N_1027);
nor U1198 (N_1198,N_1003,N_1026);
or U1199 (N_1199,N_1040,N_1019);
and U1200 (N_1200,N_1128,N_1148);
xor U1201 (N_1201,N_1170,N_1166);
and U1202 (N_1202,N_1136,N_1134);
nor U1203 (N_1203,N_1145,N_1182);
or U1204 (N_1204,N_1159,N_1175);
nor U1205 (N_1205,N_1196,N_1149);
nand U1206 (N_1206,N_1123,N_1115);
nor U1207 (N_1207,N_1171,N_1199);
nand U1208 (N_1208,N_1185,N_1108);
xnor U1209 (N_1209,N_1156,N_1154);
and U1210 (N_1210,N_1152,N_1127);
nor U1211 (N_1211,N_1193,N_1177);
nand U1212 (N_1212,N_1183,N_1186);
nand U1213 (N_1213,N_1144,N_1167);
or U1214 (N_1214,N_1140,N_1151);
and U1215 (N_1215,N_1181,N_1137);
or U1216 (N_1216,N_1133,N_1110);
or U1217 (N_1217,N_1172,N_1132);
nand U1218 (N_1218,N_1142,N_1104);
xnor U1219 (N_1219,N_1195,N_1153);
nor U1220 (N_1220,N_1117,N_1173);
nor U1221 (N_1221,N_1189,N_1118);
and U1222 (N_1222,N_1163,N_1155);
and U1223 (N_1223,N_1114,N_1116);
or U1224 (N_1224,N_1120,N_1161);
nand U1225 (N_1225,N_1109,N_1174);
and U1226 (N_1226,N_1184,N_1150);
xor U1227 (N_1227,N_1157,N_1121);
or U1228 (N_1228,N_1139,N_1122);
or U1229 (N_1229,N_1165,N_1101);
and U1230 (N_1230,N_1158,N_1105);
nor U1231 (N_1231,N_1112,N_1119);
and U1232 (N_1232,N_1138,N_1194);
nor U1233 (N_1233,N_1188,N_1103);
nand U1234 (N_1234,N_1143,N_1198);
and U1235 (N_1235,N_1169,N_1107);
nor U1236 (N_1236,N_1113,N_1100);
or U1237 (N_1237,N_1106,N_1147);
or U1238 (N_1238,N_1111,N_1190);
and U1239 (N_1239,N_1141,N_1197);
and U1240 (N_1240,N_1176,N_1179);
or U1241 (N_1241,N_1178,N_1146);
and U1242 (N_1242,N_1180,N_1191);
nand U1243 (N_1243,N_1162,N_1192);
and U1244 (N_1244,N_1160,N_1164);
or U1245 (N_1245,N_1126,N_1102);
nand U1246 (N_1246,N_1187,N_1125);
and U1247 (N_1247,N_1129,N_1131);
and U1248 (N_1248,N_1130,N_1168);
or U1249 (N_1249,N_1135,N_1124);
or U1250 (N_1250,N_1142,N_1197);
nor U1251 (N_1251,N_1112,N_1133);
xnor U1252 (N_1252,N_1122,N_1178);
or U1253 (N_1253,N_1193,N_1154);
or U1254 (N_1254,N_1176,N_1121);
nor U1255 (N_1255,N_1177,N_1127);
and U1256 (N_1256,N_1148,N_1171);
and U1257 (N_1257,N_1188,N_1139);
or U1258 (N_1258,N_1185,N_1198);
and U1259 (N_1259,N_1115,N_1157);
and U1260 (N_1260,N_1185,N_1142);
and U1261 (N_1261,N_1109,N_1123);
nor U1262 (N_1262,N_1109,N_1119);
nand U1263 (N_1263,N_1181,N_1168);
or U1264 (N_1264,N_1188,N_1149);
and U1265 (N_1265,N_1127,N_1142);
or U1266 (N_1266,N_1105,N_1155);
or U1267 (N_1267,N_1164,N_1151);
and U1268 (N_1268,N_1171,N_1186);
and U1269 (N_1269,N_1124,N_1103);
nand U1270 (N_1270,N_1149,N_1153);
or U1271 (N_1271,N_1164,N_1149);
nor U1272 (N_1272,N_1177,N_1159);
nor U1273 (N_1273,N_1195,N_1121);
or U1274 (N_1274,N_1148,N_1165);
or U1275 (N_1275,N_1108,N_1186);
nor U1276 (N_1276,N_1129,N_1152);
nor U1277 (N_1277,N_1132,N_1195);
or U1278 (N_1278,N_1144,N_1172);
nor U1279 (N_1279,N_1173,N_1147);
or U1280 (N_1280,N_1154,N_1153);
nand U1281 (N_1281,N_1178,N_1126);
nor U1282 (N_1282,N_1185,N_1138);
or U1283 (N_1283,N_1194,N_1139);
nand U1284 (N_1284,N_1140,N_1196);
or U1285 (N_1285,N_1173,N_1118);
xor U1286 (N_1286,N_1115,N_1122);
nand U1287 (N_1287,N_1166,N_1104);
xor U1288 (N_1288,N_1143,N_1118);
or U1289 (N_1289,N_1194,N_1113);
nor U1290 (N_1290,N_1138,N_1144);
xnor U1291 (N_1291,N_1184,N_1137);
nor U1292 (N_1292,N_1195,N_1189);
or U1293 (N_1293,N_1180,N_1177);
nand U1294 (N_1294,N_1168,N_1164);
xor U1295 (N_1295,N_1198,N_1134);
nand U1296 (N_1296,N_1128,N_1160);
and U1297 (N_1297,N_1110,N_1178);
nand U1298 (N_1298,N_1178,N_1131);
or U1299 (N_1299,N_1124,N_1164);
nand U1300 (N_1300,N_1292,N_1265);
nor U1301 (N_1301,N_1279,N_1210);
and U1302 (N_1302,N_1207,N_1239);
nand U1303 (N_1303,N_1209,N_1244);
nand U1304 (N_1304,N_1232,N_1272);
xor U1305 (N_1305,N_1212,N_1243);
nor U1306 (N_1306,N_1205,N_1219);
or U1307 (N_1307,N_1280,N_1294);
xnor U1308 (N_1308,N_1284,N_1221);
or U1309 (N_1309,N_1249,N_1228);
or U1310 (N_1310,N_1267,N_1213);
nor U1311 (N_1311,N_1214,N_1278);
or U1312 (N_1312,N_1261,N_1256);
or U1313 (N_1313,N_1231,N_1283);
or U1314 (N_1314,N_1201,N_1252);
and U1315 (N_1315,N_1296,N_1206);
and U1316 (N_1316,N_1250,N_1290);
nor U1317 (N_1317,N_1247,N_1200);
nor U1318 (N_1318,N_1226,N_1215);
nor U1319 (N_1319,N_1277,N_1258);
nor U1320 (N_1320,N_1276,N_1240);
nor U1321 (N_1321,N_1237,N_1208);
or U1322 (N_1322,N_1230,N_1217);
xnor U1323 (N_1323,N_1235,N_1211);
nor U1324 (N_1324,N_1248,N_1238);
nand U1325 (N_1325,N_1224,N_1297);
nor U1326 (N_1326,N_1263,N_1289);
nor U1327 (N_1327,N_1233,N_1225);
or U1328 (N_1328,N_1274,N_1227);
or U1329 (N_1329,N_1273,N_1220);
and U1330 (N_1330,N_1236,N_1241);
nor U1331 (N_1331,N_1275,N_1253);
nand U1332 (N_1332,N_1281,N_1271);
xor U1333 (N_1333,N_1223,N_1268);
and U1334 (N_1334,N_1222,N_1266);
and U1335 (N_1335,N_1285,N_1255);
nor U1336 (N_1336,N_1287,N_1262);
xor U1337 (N_1337,N_1257,N_1229);
or U1338 (N_1338,N_1282,N_1270);
nor U1339 (N_1339,N_1246,N_1234);
xnor U1340 (N_1340,N_1264,N_1216);
and U1341 (N_1341,N_1295,N_1202);
xnor U1342 (N_1342,N_1204,N_1259);
nand U1343 (N_1343,N_1291,N_1251);
or U1344 (N_1344,N_1218,N_1269);
or U1345 (N_1345,N_1260,N_1293);
or U1346 (N_1346,N_1286,N_1245);
nand U1347 (N_1347,N_1242,N_1203);
and U1348 (N_1348,N_1254,N_1288);
and U1349 (N_1349,N_1299,N_1298);
or U1350 (N_1350,N_1210,N_1241);
xnor U1351 (N_1351,N_1289,N_1202);
or U1352 (N_1352,N_1223,N_1282);
or U1353 (N_1353,N_1204,N_1271);
and U1354 (N_1354,N_1211,N_1225);
nor U1355 (N_1355,N_1266,N_1293);
nand U1356 (N_1356,N_1285,N_1294);
xnor U1357 (N_1357,N_1216,N_1290);
xnor U1358 (N_1358,N_1205,N_1285);
xnor U1359 (N_1359,N_1295,N_1273);
or U1360 (N_1360,N_1237,N_1235);
and U1361 (N_1361,N_1248,N_1244);
and U1362 (N_1362,N_1239,N_1260);
nor U1363 (N_1363,N_1278,N_1202);
nand U1364 (N_1364,N_1240,N_1226);
or U1365 (N_1365,N_1280,N_1214);
nor U1366 (N_1366,N_1210,N_1229);
and U1367 (N_1367,N_1203,N_1254);
nand U1368 (N_1368,N_1209,N_1298);
or U1369 (N_1369,N_1278,N_1201);
or U1370 (N_1370,N_1255,N_1237);
nand U1371 (N_1371,N_1294,N_1293);
and U1372 (N_1372,N_1265,N_1246);
nand U1373 (N_1373,N_1282,N_1207);
nand U1374 (N_1374,N_1286,N_1209);
nand U1375 (N_1375,N_1295,N_1276);
nand U1376 (N_1376,N_1298,N_1293);
nand U1377 (N_1377,N_1266,N_1287);
nor U1378 (N_1378,N_1238,N_1256);
or U1379 (N_1379,N_1298,N_1235);
nor U1380 (N_1380,N_1256,N_1269);
xor U1381 (N_1381,N_1298,N_1233);
and U1382 (N_1382,N_1258,N_1243);
or U1383 (N_1383,N_1272,N_1237);
nor U1384 (N_1384,N_1201,N_1240);
nor U1385 (N_1385,N_1213,N_1271);
nand U1386 (N_1386,N_1299,N_1241);
and U1387 (N_1387,N_1237,N_1271);
nand U1388 (N_1388,N_1276,N_1272);
and U1389 (N_1389,N_1240,N_1278);
xor U1390 (N_1390,N_1291,N_1281);
xor U1391 (N_1391,N_1200,N_1205);
and U1392 (N_1392,N_1226,N_1273);
or U1393 (N_1393,N_1202,N_1239);
and U1394 (N_1394,N_1298,N_1204);
xnor U1395 (N_1395,N_1280,N_1272);
and U1396 (N_1396,N_1295,N_1236);
or U1397 (N_1397,N_1264,N_1204);
or U1398 (N_1398,N_1212,N_1279);
xnor U1399 (N_1399,N_1253,N_1280);
and U1400 (N_1400,N_1388,N_1396);
nand U1401 (N_1401,N_1355,N_1327);
or U1402 (N_1402,N_1307,N_1311);
nor U1403 (N_1403,N_1370,N_1323);
or U1404 (N_1404,N_1309,N_1363);
and U1405 (N_1405,N_1302,N_1395);
or U1406 (N_1406,N_1352,N_1332);
nor U1407 (N_1407,N_1320,N_1331);
nor U1408 (N_1408,N_1358,N_1350);
nand U1409 (N_1409,N_1360,N_1397);
nor U1410 (N_1410,N_1381,N_1379);
nor U1411 (N_1411,N_1326,N_1303);
nand U1412 (N_1412,N_1305,N_1371);
nor U1413 (N_1413,N_1349,N_1362);
and U1414 (N_1414,N_1384,N_1330);
xor U1415 (N_1415,N_1333,N_1301);
nand U1416 (N_1416,N_1375,N_1342);
and U1417 (N_1417,N_1361,N_1329);
xor U1418 (N_1418,N_1316,N_1345);
or U1419 (N_1419,N_1373,N_1359);
nand U1420 (N_1420,N_1341,N_1368);
or U1421 (N_1421,N_1313,N_1365);
nor U1422 (N_1422,N_1377,N_1337);
and U1423 (N_1423,N_1351,N_1385);
nor U1424 (N_1424,N_1389,N_1340);
nor U1425 (N_1425,N_1339,N_1399);
and U1426 (N_1426,N_1354,N_1328);
and U1427 (N_1427,N_1312,N_1335);
nor U1428 (N_1428,N_1336,N_1324);
nand U1429 (N_1429,N_1394,N_1321);
or U1430 (N_1430,N_1383,N_1391);
nor U1431 (N_1431,N_1357,N_1376);
nand U1432 (N_1432,N_1304,N_1382);
nor U1433 (N_1433,N_1334,N_1378);
or U1434 (N_1434,N_1356,N_1364);
nand U1435 (N_1435,N_1317,N_1398);
nor U1436 (N_1436,N_1314,N_1306);
and U1437 (N_1437,N_1322,N_1392);
or U1438 (N_1438,N_1319,N_1386);
nor U1439 (N_1439,N_1338,N_1346);
nor U1440 (N_1440,N_1344,N_1347);
and U1441 (N_1441,N_1369,N_1325);
nor U1442 (N_1442,N_1315,N_1387);
or U1443 (N_1443,N_1366,N_1348);
nor U1444 (N_1444,N_1372,N_1367);
or U1445 (N_1445,N_1374,N_1343);
nor U1446 (N_1446,N_1353,N_1390);
nor U1447 (N_1447,N_1308,N_1393);
or U1448 (N_1448,N_1310,N_1380);
nor U1449 (N_1449,N_1318,N_1300);
nand U1450 (N_1450,N_1392,N_1350);
or U1451 (N_1451,N_1368,N_1311);
nor U1452 (N_1452,N_1338,N_1354);
nor U1453 (N_1453,N_1359,N_1329);
nand U1454 (N_1454,N_1396,N_1369);
or U1455 (N_1455,N_1319,N_1340);
and U1456 (N_1456,N_1356,N_1334);
xnor U1457 (N_1457,N_1359,N_1317);
and U1458 (N_1458,N_1360,N_1303);
xnor U1459 (N_1459,N_1335,N_1300);
and U1460 (N_1460,N_1368,N_1379);
nand U1461 (N_1461,N_1354,N_1358);
nand U1462 (N_1462,N_1305,N_1369);
nor U1463 (N_1463,N_1395,N_1352);
and U1464 (N_1464,N_1372,N_1363);
and U1465 (N_1465,N_1327,N_1330);
and U1466 (N_1466,N_1393,N_1395);
nand U1467 (N_1467,N_1347,N_1370);
nor U1468 (N_1468,N_1323,N_1335);
and U1469 (N_1469,N_1377,N_1346);
nor U1470 (N_1470,N_1354,N_1382);
xor U1471 (N_1471,N_1361,N_1304);
nand U1472 (N_1472,N_1356,N_1339);
nor U1473 (N_1473,N_1399,N_1360);
nor U1474 (N_1474,N_1336,N_1372);
and U1475 (N_1475,N_1324,N_1321);
or U1476 (N_1476,N_1345,N_1320);
and U1477 (N_1477,N_1356,N_1384);
or U1478 (N_1478,N_1385,N_1376);
and U1479 (N_1479,N_1307,N_1343);
nand U1480 (N_1480,N_1372,N_1396);
xor U1481 (N_1481,N_1326,N_1388);
or U1482 (N_1482,N_1345,N_1308);
and U1483 (N_1483,N_1353,N_1340);
and U1484 (N_1484,N_1363,N_1347);
nor U1485 (N_1485,N_1320,N_1313);
nor U1486 (N_1486,N_1334,N_1335);
and U1487 (N_1487,N_1387,N_1328);
nand U1488 (N_1488,N_1368,N_1313);
nor U1489 (N_1489,N_1386,N_1341);
nand U1490 (N_1490,N_1322,N_1337);
and U1491 (N_1491,N_1312,N_1365);
or U1492 (N_1492,N_1315,N_1385);
nand U1493 (N_1493,N_1379,N_1385);
nor U1494 (N_1494,N_1307,N_1359);
nand U1495 (N_1495,N_1394,N_1328);
nand U1496 (N_1496,N_1327,N_1314);
nand U1497 (N_1497,N_1375,N_1336);
or U1498 (N_1498,N_1337,N_1316);
and U1499 (N_1499,N_1380,N_1378);
xor U1500 (N_1500,N_1455,N_1415);
nor U1501 (N_1501,N_1450,N_1418);
nand U1502 (N_1502,N_1437,N_1425);
nand U1503 (N_1503,N_1493,N_1475);
xnor U1504 (N_1504,N_1491,N_1471);
or U1505 (N_1505,N_1454,N_1453);
and U1506 (N_1506,N_1497,N_1487);
nor U1507 (N_1507,N_1441,N_1424);
xnor U1508 (N_1508,N_1495,N_1488);
nand U1509 (N_1509,N_1414,N_1472);
or U1510 (N_1510,N_1486,N_1461);
nor U1511 (N_1511,N_1481,N_1440);
nand U1512 (N_1512,N_1462,N_1449);
nand U1513 (N_1513,N_1484,N_1445);
xor U1514 (N_1514,N_1436,N_1490);
or U1515 (N_1515,N_1443,N_1404);
or U1516 (N_1516,N_1456,N_1410);
nor U1517 (N_1517,N_1435,N_1431);
and U1518 (N_1518,N_1407,N_1460);
or U1519 (N_1519,N_1419,N_1478);
and U1520 (N_1520,N_1458,N_1479);
or U1521 (N_1521,N_1464,N_1423);
nand U1522 (N_1522,N_1499,N_1476);
nand U1523 (N_1523,N_1451,N_1405);
nand U1524 (N_1524,N_1459,N_1469);
xnor U1525 (N_1525,N_1442,N_1447);
and U1526 (N_1526,N_1463,N_1483);
nand U1527 (N_1527,N_1422,N_1411);
or U1528 (N_1528,N_1485,N_1421);
or U1529 (N_1529,N_1473,N_1465);
nand U1530 (N_1530,N_1428,N_1413);
xor U1531 (N_1531,N_1409,N_1444);
nor U1532 (N_1532,N_1408,N_1489);
xnor U1533 (N_1533,N_1429,N_1482);
xor U1534 (N_1534,N_1467,N_1420);
and U1535 (N_1535,N_1496,N_1434);
or U1536 (N_1536,N_1432,N_1498);
nand U1537 (N_1537,N_1401,N_1417);
and U1538 (N_1538,N_1452,N_1448);
xor U1539 (N_1539,N_1430,N_1466);
or U1540 (N_1540,N_1494,N_1400);
or U1541 (N_1541,N_1468,N_1492);
nor U1542 (N_1542,N_1446,N_1439);
nand U1543 (N_1543,N_1412,N_1470);
nor U1544 (N_1544,N_1457,N_1477);
or U1545 (N_1545,N_1438,N_1402);
xnor U1546 (N_1546,N_1403,N_1427);
nand U1547 (N_1547,N_1406,N_1433);
nor U1548 (N_1548,N_1474,N_1480);
nand U1549 (N_1549,N_1416,N_1426);
nor U1550 (N_1550,N_1481,N_1401);
nand U1551 (N_1551,N_1449,N_1436);
nor U1552 (N_1552,N_1469,N_1416);
and U1553 (N_1553,N_1492,N_1488);
or U1554 (N_1554,N_1410,N_1420);
nor U1555 (N_1555,N_1482,N_1434);
and U1556 (N_1556,N_1441,N_1401);
nor U1557 (N_1557,N_1457,N_1497);
and U1558 (N_1558,N_1481,N_1463);
nand U1559 (N_1559,N_1437,N_1414);
and U1560 (N_1560,N_1458,N_1456);
nor U1561 (N_1561,N_1404,N_1407);
nand U1562 (N_1562,N_1497,N_1422);
and U1563 (N_1563,N_1420,N_1418);
xnor U1564 (N_1564,N_1446,N_1437);
xnor U1565 (N_1565,N_1406,N_1455);
or U1566 (N_1566,N_1495,N_1458);
nor U1567 (N_1567,N_1487,N_1410);
nor U1568 (N_1568,N_1424,N_1499);
nor U1569 (N_1569,N_1436,N_1479);
nor U1570 (N_1570,N_1468,N_1499);
and U1571 (N_1571,N_1476,N_1418);
and U1572 (N_1572,N_1453,N_1431);
or U1573 (N_1573,N_1493,N_1402);
nand U1574 (N_1574,N_1474,N_1468);
and U1575 (N_1575,N_1479,N_1462);
and U1576 (N_1576,N_1412,N_1413);
nor U1577 (N_1577,N_1415,N_1492);
nand U1578 (N_1578,N_1422,N_1455);
or U1579 (N_1579,N_1450,N_1470);
nor U1580 (N_1580,N_1450,N_1426);
nand U1581 (N_1581,N_1424,N_1461);
xnor U1582 (N_1582,N_1484,N_1447);
nor U1583 (N_1583,N_1443,N_1475);
nor U1584 (N_1584,N_1486,N_1438);
or U1585 (N_1585,N_1492,N_1495);
nand U1586 (N_1586,N_1450,N_1437);
nor U1587 (N_1587,N_1457,N_1453);
nand U1588 (N_1588,N_1446,N_1412);
or U1589 (N_1589,N_1417,N_1480);
nand U1590 (N_1590,N_1453,N_1444);
xor U1591 (N_1591,N_1448,N_1435);
and U1592 (N_1592,N_1438,N_1485);
and U1593 (N_1593,N_1432,N_1403);
nand U1594 (N_1594,N_1492,N_1424);
xor U1595 (N_1595,N_1484,N_1480);
nand U1596 (N_1596,N_1471,N_1453);
or U1597 (N_1597,N_1407,N_1451);
nor U1598 (N_1598,N_1488,N_1436);
or U1599 (N_1599,N_1449,N_1482);
and U1600 (N_1600,N_1503,N_1570);
or U1601 (N_1601,N_1545,N_1586);
nand U1602 (N_1602,N_1557,N_1564);
nor U1603 (N_1603,N_1520,N_1597);
or U1604 (N_1604,N_1535,N_1534);
or U1605 (N_1605,N_1538,N_1566);
nor U1606 (N_1606,N_1562,N_1536);
nor U1607 (N_1607,N_1507,N_1589);
and U1608 (N_1608,N_1584,N_1568);
or U1609 (N_1609,N_1574,N_1509);
or U1610 (N_1610,N_1581,N_1513);
or U1611 (N_1611,N_1529,N_1593);
nor U1612 (N_1612,N_1516,N_1549);
or U1613 (N_1613,N_1525,N_1523);
and U1614 (N_1614,N_1576,N_1553);
nor U1615 (N_1615,N_1548,N_1533);
and U1616 (N_1616,N_1541,N_1588);
nand U1617 (N_1617,N_1579,N_1591);
or U1618 (N_1618,N_1505,N_1599);
or U1619 (N_1619,N_1572,N_1531);
and U1620 (N_1620,N_1573,N_1590);
or U1621 (N_1621,N_1506,N_1527);
or U1622 (N_1622,N_1511,N_1580);
or U1623 (N_1623,N_1567,N_1571);
and U1624 (N_1624,N_1550,N_1504);
xor U1625 (N_1625,N_1582,N_1546);
and U1626 (N_1626,N_1592,N_1502);
nand U1627 (N_1627,N_1542,N_1585);
nor U1628 (N_1628,N_1555,N_1594);
nand U1629 (N_1629,N_1543,N_1521);
or U1630 (N_1630,N_1598,N_1596);
or U1631 (N_1631,N_1563,N_1522);
nand U1632 (N_1632,N_1551,N_1547);
and U1633 (N_1633,N_1540,N_1569);
nand U1634 (N_1634,N_1518,N_1528);
and U1635 (N_1635,N_1539,N_1530);
nor U1636 (N_1636,N_1565,N_1517);
or U1637 (N_1637,N_1515,N_1554);
nand U1638 (N_1638,N_1577,N_1552);
and U1639 (N_1639,N_1512,N_1508);
nor U1640 (N_1640,N_1561,N_1575);
and U1641 (N_1641,N_1578,N_1501);
xnor U1642 (N_1642,N_1556,N_1524);
and U1643 (N_1643,N_1510,N_1583);
or U1644 (N_1644,N_1514,N_1587);
nand U1645 (N_1645,N_1558,N_1559);
or U1646 (N_1646,N_1544,N_1526);
nor U1647 (N_1647,N_1500,N_1537);
nor U1648 (N_1648,N_1560,N_1519);
and U1649 (N_1649,N_1532,N_1595);
nor U1650 (N_1650,N_1512,N_1524);
and U1651 (N_1651,N_1595,N_1588);
nor U1652 (N_1652,N_1564,N_1560);
and U1653 (N_1653,N_1554,N_1505);
nor U1654 (N_1654,N_1594,N_1537);
and U1655 (N_1655,N_1586,N_1521);
nor U1656 (N_1656,N_1552,N_1530);
xor U1657 (N_1657,N_1587,N_1552);
nor U1658 (N_1658,N_1518,N_1540);
nand U1659 (N_1659,N_1557,N_1535);
nor U1660 (N_1660,N_1587,N_1538);
xnor U1661 (N_1661,N_1543,N_1523);
nand U1662 (N_1662,N_1573,N_1561);
and U1663 (N_1663,N_1574,N_1566);
or U1664 (N_1664,N_1563,N_1511);
nand U1665 (N_1665,N_1518,N_1531);
and U1666 (N_1666,N_1501,N_1556);
and U1667 (N_1667,N_1533,N_1513);
nand U1668 (N_1668,N_1549,N_1557);
nor U1669 (N_1669,N_1508,N_1517);
xnor U1670 (N_1670,N_1543,N_1589);
or U1671 (N_1671,N_1599,N_1509);
nor U1672 (N_1672,N_1598,N_1552);
or U1673 (N_1673,N_1588,N_1519);
nor U1674 (N_1674,N_1500,N_1599);
nand U1675 (N_1675,N_1530,N_1596);
or U1676 (N_1676,N_1596,N_1556);
nor U1677 (N_1677,N_1506,N_1501);
and U1678 (N_1678,N_1543,N_1519);
nor U1679 (N_1679,N_1538,N_1546);
xnor U1680 (N_1680,N_1529,N_1518);
nand U1681 (N_1681,N_1539,N_1557);
or U1682 (N_1682,N_1526,N_1537);
nor U1683 (N_1683,N_1518,N_1564);
or U1684 (N_1684,N_1580,N_1598);
nand U1685 (N_1685,N_1579,N_1543);
and U1686 (N_1686,N_1586,N_1599);
xor U1687 (N_1687,N_1510,N_1528);
or U1688 (N_1688,N_1507,N_1509);
or U1689 (N_1689,N_1519,N_1554);
or U1690 (N_1690,N_1513,N_1524);
nor U1691 (N_1691,N_1587,N_1546);
and U1692 (N_1692,N_1592,N_1575);
nand U1693 (N_1693,N_1565,N_1505);
or U1694 (N_1694,N_1527,N_1532);
nor U1695 (N_1695,N_1539,N_1566);
xor U1696 (N_1696,N_1582,N_1502);
or U1697 (N_1697,N_1509,N_1591);
or U1698 (N_1698,N_1516,N_1578);
or U1699 (N_1699,N_1505,N_1546);
nand U1700 (N_1700,N_1649,N_1656);
nand U1701 (N_1701,N_1606,N_1674);
or U1702 (N_1702,N_1685,N_1634);
and U1703 (N_1703,N_1638,N_1667);
or U1704 (N_1704,N_1688,N_1619);
nand U1705 (N_1705,N_1684,N_1600);
and U1706 (N_1706,N_1615,N_1612);
nor U1707 (N_1707,N_1694,N_1621);
nor U1708 (N_1708,N_1658,N_1641);
nand U1709 (N_1709,N_1624,N_1692);
or U1710 (N_1710,N_1661,N_1601);
nor U1711 (N_1711,N_1611,N_1603);
nor U1712 (N_1712,N_1698,N_1610);
and U1713 (N_1713,N_1676,N_1617);
nor U1714 (N_1714,N_1648,N_1637);
or U1715 (N_1715,N_1664,N_1643);
and U1716 (N_1716,N_1630,N_1635);
or U1717 (N_1717,N_1652,N_1618);
nor U1718 (N_1718,N_1699,N_1680);
nand U1719 (N_1719,N_1631,N_1696);
nand U1720 (N_1720,N_1689,N_1690);
or U1721 (N_1721,N_1679,N_1670);
nand U1722 (N_1722,N_1636,N_1678);
nand U1723 (N_1723,N_1681,N_1697);
or U1724 (N_1724,N_1626,N_1687);
and U1725 (N_1725,N_1608,N_1673);
and U1726 (N_1726,N_1647,N_1614);
or U1727 (N_1727,N_1682,N_1616);
xor U1728 (N_1728,N_1665,N_1642);
nand U1729 (N_1729,N_1640,N_1651);
nor U1730 (N_1730,N_1604,N_1622);
nor U1731 (N_1731,N_1632,N_1693);
nand U1732 (N_1732,N_1650,N_1683);
or U1733 (N_1733,N_1628,N_1659);
nand U1734 (N_1734,N_1629,N_1675);
nand U1735 (N_1735,N_1645,N_1633);
nand U1736 (N_1736,N_1691,N_1686);
nand U1737 (N_1737,N_1657,N_1669);
or U1738 (N_1738,N_1602,N_1695);
xnor U1739 (N_1739,N_1607,N_1671);
nor U1740 (N_1740,N_1668,N_1666);
and U1741 (N_1741,N_1660,N_1644);
nor U1742 (N_1742,N_1672,N_1653);
or U1743 (N_1743,N_1613,N_1620);
nor U1744 (N_1744,N_1654,N_1639);
xnor U1745 (N_1745,N_1625,N_1662);
or U1746 (N_1746,N_1663,N_1655);
and U1747 (N_1747,N_1623,N_1646);
nor U1748 (N_1748,N_1605,N_1627);
or U1749 (N_1749,N_1609,N_1677);
and U1750 (N_1750,N_1660,N_1627);
and U1751 (N_1751,N_1641,N_1677);
or U1752 (N_1752,N_1662,N_1634);
or U1753 (N_1753,N_1608,N_1680);
or U1754 (N_1754,N_1664,N_1686);
nand U1755 (N_1755,N_1628,N_1632);
nand U1756 (N_1756,N_1684,N_1638);
xnor U1757 (N_1757,N_1648,N_1683);
nor U1758 (N_1758,N_1609,N_1675);
and U1759 (N_1759,N_1660,N_1674);
nor U1760 (N_1760,N_1683,N_1670);
nor U1761 (N_1761,N_1648,N_1632);
and U1762 (N_1762,N_1684,N_1660);
and U1763 (N_1763,N_1657,N_1638);
or U1764 (N_1764,N_1639,N_1657);
nor U1765 (N_1765,N_1622,N_1692);
nand U1766 (N_1766,N_1695,N_1673);
nand U1767 (N_1767,N_1629,N_1655);
xor U1768 (N_1768,N_1693,N_1623);
nor U1769 (N_1769,N_1661,N_1638);
xor U1770 (N_1770,N_1614,N_1667);
nand U1771 (N_1771,N_1600,N_1614);
nand U1772 (N_1772,N_1601,N_1691);
nor U1773 (N_1773,N_1648,N_1680);
or U1774 (N_1774,N_1685,N_1658);
nand U1775 (N_1775,N_1611,N_1680);
nor U1776 (N_1776,N_1686,N_1674);
nor U1777 (N_1777,N_1646,N_1688);
nand U1778 (N_1778,N_1612,N_1655);
or U1779 (N_1779,N_1638,N_1616);
and U1780 (N_1780,N_1652,N_1676);
nand U1781 (N_1781,N_1695,N_1668);
or U1782 (N_1782,N_1630,N_1628);
and U1783 (N_1783,N_1677,N_1685);
nand U1784 (N_1784,N_1659,N_1620);
xor U1785 (N_1785,N_1623,N_1627);
nand U1786 (N_1786,N_1607,N_1633);
and U1787 (N_1787,N_1672,N_1693);
and U1788 (N_1788,N_1604,N_1615);
or U1789 (N_1789,N_1637,N_1674);
nand U1790 (N_1790,N_1641,N_1639);
and U1791 (N_1791,N_1653,N_1670);
nor U1792 (N_1792,N_1638,N_1619);
and U1793 (N_1793,N_1626,N_1677);
nand U1794 (N_1794,N_1615,N_1627);
or U1795 (N_1795,N_1626,N_1632);
nor U1796 (N_1796,N_1662,N_1699);
and U1797 (N_1797,N_1642,N_1689);
or U1798 (N_1798,N_1665,N_1612);
or U1799 (N_1799,N_1635,N_1624);
and U1800 (N_1800,N_1762,N_1765);
and U1801 (N_1801,N_1750,N_1714);
nor U1802 (N_1802,N_1798,N_1717);
nor U1803 (N_1803,N_1758,N_1755);
nor U1804 (N_1804,N_1757,N_1715);
xnor U1805 (N_1805,N_1781,N_1733);
xor U1806 (N_1806,N_1799,N_1764);
nand U1807 (N_1807,N_1761,N_1794);
nor U1808 (N_1808,N_1740,N_1713);
or U1809 (N_1809,N_1707,N_1780);
nor U1810 (N_1810,N_1743,N_1720);
nand U1811 (N_1811,N_1752,N_1741);
xor U1812 (N_1812,N_1775,N_1759);
or U1813 (N_1813,N_1760,N_1788);
or U1814 (N_1814,N_1705,N_1744);
nand U1815 (N_1815,N_1732,N_1790);
nor U1816 (N_1816,N_1769,N_1748);
and U1817 (N_1817,N_1751,N_1789);
and U1818 (N_1818,N_1702,N_1722);
nand U1819 (N_1819,N_1754,N_1779);
nand U1820 (N_1820,N_1776,N_1770);
nand U1821 (N_1821,N_1735,N_1791);
nor U1822 (N_1822,N_1729,N_1785);
and U1823 (N_1823,N_1723,N_1756);
and U1824 (N_1824,N_1768,N_1766);
and U1825 (N_1825,N_1795,N_1739);
or U1826 (N_1826,N_1773,N_1709);
or U1827 (N_1827,N_1728,N_1753);
nand U1828 (N_1828,N_1749,N_1793);
nor U1829 (N_1829,N_1786,N_1763);
or U1830 (N_1830,N_1784,N_1736);
and U1831 (N_1831,N_1703,N_1767);
and U1832 (N_1832,N_1742,N_1727);
nor U1833 (N_1833,N_1772,N_1701);
nor U1834 (N_1834,N_1746,N_1700);
nor U1835 (N_1835,N_1721,N_1724);
nand U1836 (N_1836,N_1719,N_1718);
or U1837 (N_1837,N_1783,N_1708);
and U1838 (N_1838,N_1704,N_1730);
or U1839 (N_1839,N_1782,N_1725);
or U1840 (N_1840,N_1747,N_1796);
nor U1841 (N_1841,N_1738,N_1734);
nor U1842 (N_1842,N_1787,N_1792);
xor U1843 (N_1843,N_1774,N_1777);
nor U1844 (N_1844,N_1737,N_1745);
and U1845 (N_1845,N_1778,N_1711);
nor U1846 (N_1846,N_1710,N_1726);
and U1847 (N_1847,N_1731,N_1771);
nand U1848 (N_1848,N_1706,N_1712);
or U1849 (N_1849,N_1797,N_1716);
nor U1850 (N_1850,N_1701,N_1775);
or U1851 (N_1851,N_1742,N_1796);
or U1852 (N_1852,N_1712,N_1716);
xor U1853 (N_1853,N_1727,N_1753);
and U1854 (N_1854,N_1716,N_1715);
nor U1855 (N_1855,N_1723,N_1772);
and U1856 (N_1856,N_1771,N_1758);
nor U1857 (N_1857,N_1706,N_1732);
nor U1858 (N_1858,N_1705,N_1754);
nor U1859 (N_1859,N_1731,N_1752);
nand U1860 (N_1860,N_1798,N_1768);
nand U1861 (N_1861,N_1730,N_1712);
nand U1862 (N_1862,N_1725,N_1798);
nand U1863 (N_1863,N_1714,N_1758);
or U1864 (N_1864,N_1778,N_1753);
and U1865 (N_1865,N_1716,N_1764);
or U1866 (N_1866,N_1703,N_1706);
nand U1867 (N_1867,N_1770,N_1713);
nor U1868 (N_1868,N_1745,N_1750);
nor U1869 (N_1869,N_1737,N_1705);
nand U1870 (N_1870,N_1759,N_1768);
nand U1871 (N_1871,N_1791,N_1710);
and U1872 (N_1872,N_1736,N_1740);
xor U1873 (N_1873,N_1791,N_1778);
nor U1874 (N_1874,N_1772,N_1786);
or U1875 (N_1875,N_1775,N_1794);
nor U1876 (N_1876,N_1737,N_1778);
and U1877 (N_1877,N_1753,N_1777);
nor U1878 (N_1878,N_1772,N_1739);
or U1879 (N_1879,N_1707,N_1700);
nor U1880 (N_1880,N_1734,N_1701);
xnor U1881 (N_1881,N_1796,N_1774);
and U1882 (N_1882,N_1797,N_1778);
or U1883 (N_1883,N_1751,N_1753);
and U1884 (N_1884,N_1723,N_1739);
nor U1885 (N_1885,N_1748,N_1720);
and U1886 (N_1886,N_1752,N_1798);
nand U1887 (N_1887,N_1768,N_1711);
or U1888 (N_1888,N_1768,N_1701);
or U1889 (N_1889,N_1798,N_1747);
and U1890 (N_1890,N_1770,N_1714);
and U1891 (N_1891,N_1712,N_1742);
or U1892 (N_1892,N_1750,N_1788);
or U1893 (N_1893,N_1798,N_1779);
nor U1894 (N_1894,N_1739,N_1778);
and U1895 (N_1895,N_1755,N_1770);
nand U1896 (N_1896,N_1713,N_1760);
nand U1897 (N_1897,N_1711,N_1741);
xnor U1898 (N_1898,N_1720,N_1714);
and U1899 (N_1899,N_1763,N_1779);
nand U1900 (N_1900,N_1865,N_1888);
or U1901 (N_1901,N_1850,N_1818);
nor U1902 (N_1902,N_1824,N_1806);
nand U1903 (N_1903,N_1879,N_1863);
xor U1904 (N_1904,N_1851,N_1802);
nor U1905 (N_1905,N_1871,N_1856);
or U1906 (N_1906,N_1804,N_1892);
nand U1907 (N_1907,N_1861,N_1897);
xor U1908 (N_1908,N_1822,N_1829);
nor U1909 (N_1909,N_1853,N_1884);
or U1910 (N_1910,N_1858,N_1898);
and U1911 (N_1911,N_1868,N_1881);
nor U1912 (N_1912,N_1876,N_1820);
and U1913 (N_1913,N_1873,N_1852);
nor U1914 (N_1914,N_1813,N_1840);
nor U1915 (N_1915,N_1836,N_1859);
nand U1916 (N_1916,N_1827,N_1831);
xor U1917 (N_1917,N_1855,N_1830);
nand U1918 (N_1918,N_1832,N_1842);
and U1919 (N_1919,N_1886,N_1843);
nand U1920 (N_1920,N_1841,N_1833);
and U1921 (N_1921,N_1870,N_1800);
xor U1922 (N_1922,N_1882,N_1810);
nor U1923 (N_1923,N_1834,N_1819);
nand U1924 (N_1924,N_1809,N_1825);
or U1925 (N_1925,N_1883,N_1846);
nor U1926 (N_1926,N_1838,N_1805);
or U1927 (N_1927,N_1869,N_1889);
nor U1928 (N_1928,N_1862,N_1814);
and U1929 (N_1929,N_1821,N_1885);
and U1930 (N_1930,N_1887,N_1812);
or U1931 (N_1931,N_1864,N_1828);
nand U1932 (N_1932,N_1847,N_1866);
nor U1933 (N_1933,N_1803,N_1880);
and U1934 (N_1934,N_1890,N_1893);
nand U1935 (N_1935,N_1857,N_1867);
nor U1936 (N_1936,N_1811,N_1872);
and U1937 (N_1937,N_1895,N_1826);
or U1938 (N_1938,N_1808,N_1815);
xor U1939 (N_1939,N_1875,N_1845);
and U1940 (N_1940,N_1835,N_1894);
xor U1941 (N_1941,N_1848,N_1844);
and U1942 (N_1942,N_1854,N_1816);
xor U1943 (N_1943,N_1801,N_1896);
or U1944 (N_1944,N_1899,N_1878);
xor U1945 (N_1945,N_1849,N_1860);
nand U1946 (N_1946,N_1837,N_1817);
nor U1947 (N_1947,N_1877,N_1839);
and U1948 (N_1948,N_1823,N_1874);
and U1949 (N_1949,N_1807,N_1891);
nand U1950 (N_1950,N_1842,N_1824);
xnor U1951 (N_1951,N_1896,N_1880);
nor U1952 (N_1952,N_1875,N_1872);
xnor U1953 (N_1953,N_1858,N_1856);
xor U1954 (N_1954,N_1858,N_1890);
and U1955 (N_1955,N_1835,N_1813);
or U1956 (N_1956,N_1833,N_1802);
nor U1957 (N_1957,N_1828,N_1846);
or U1958 (N_1958,N_1819,N_1860);
or U1959 (N_1959,N_1865,N_1854);
and U1960 (N_1960,N_1879,N_1827);
nor U1961 (N_1961,N_1861,N_1885);
and U1962 (N_1962,N_1869,N_1810);
nand U1963 (N_1963,N_1880,N_1891);
or U1964 (N_1964,N_1856,N_1828);
and U1965 (N_1965,N_1809,N_1842);
or U1966 (N_1966,N_1898,N_1819);
nand U1967 (N_1967,N_1842,N_1816);
nor U1968 (N_1968,N_1807,N_1869);
and U1969 (N_1969,N_1844,N_1876);
xnor U1970 (N_1970,N_1876,N_1856);
or U1971 (N_1971,N_1819,N_1817);
xor U1972 (N_1972,N_1893,N_1807);
xor U1973 (N_1973,N_1845,N_1894);
and U1974 (N_1974,N_1881,N_1830);
or U1975 (N_1975,N_1898,N_1864);
or U1976 (N_1976,N_1866,N_1800);
and U1977 (N_1977,N_1807,N_1875);
or U1978 (N_1978,N_1880,N_1820);
or U1979 (N_1979,N_1866,N_1842);
nor U1980 (N_1980,N_1868,N_1839);
nor U1981 (N_1981,N_1835,N_1865);
or U1982 (N_1982,N_1848,N_1852);
nand U1983 (N_1983,N_1872,N_1829);
and U1984 (N_1984,N_1894,N_1812);
nor U1985 (N_1985,N_1849,N_1857);
or U1986 (N_1986,N_1878,N_1898);
and U1987 (N_1987,N_1819,N_1844);
nand U1988 (N_1988,N_1897,N_1829);
xnor U1989 (N_1989,N_1833,N_1847);
or U1990 (N_1990,N_1805,N_1871);
or U1991 (N_1991,N_1844,N_1828);
and U1992 (N_1992,N_1874,N_1853);
and U1993 (N_1993,N_1810,N_1881);
nand U1994 (N_1994,N_1843,N_1815);
nor U1995 (N_1995,N_1816,N_1883);
nor U1996 (N_1996,N_1822,N_1884);
nor U1997 (N_1997,N_1899,N_1806);
nor U1998 (N_1998,N_1869,N_1822);
nand U1999 (N_1999,N_1880,N_1823);
or U2000 (N_2000,N_1942,N_1972);
xor U2001 (N_2001,N_1932,N_1907);
nand U2002 (N_2002,N_1984,N_1902);
or U2003 (N_2003,N_1986,N_1938);
or U2004 (N_2004,N_1922,N_1904);
nand U2005 (N_2005,N_1910,N_1936);
nor U2006 (N_2006,N_1912,N_1920);
or U2007 (N_2007,N_1919,N_1924);
xor U2008 (N_2008,N_1948,N_1909);
or U2009 (N_2009,N_1917,N_1958);
nand U2010 (N_2010,N_1905,N_1908);
nand U2011 (N_2011,N_1933,N_1944);
nand U2012 (N_2012,N_1998,N_1930);
nand U2013 (N_2013,N_1900,N_1973);
nand U2014 (N_2014,N_1969,N_1923);
and U2015 (N_2015,N_1914,N_1927);
xnor U2016 (N_2016,N_1962,N_1937);
nor U2017 (N_2017,N_1964,N_1959);
nand U2018 (N_2018,N_1931,N_1989);
nand U2019 (N_2019,N_1952,N_1915);
or U2020 (N_2020,N_1946,N_1916);
nand U2021 (N_2021,N_1929,N_1971);
or U2022 (N_2022,N_1906,N_1928);
or U2023 (N_2023,N_1979,N_1983);
nor U2024 (N_2024,N_1987,N_1911);
or U2025 (N_2025,N_1975,N_1956);
xnor U2026 (N_2026,N_1992,N_1965);
nand U2027 (N_2027,N_1993,N_1966);
and U2028 (N_2028,N_1926,N_1980);
xnor U2029 (N_2029,N_1985,N_1955);
or U2030 (N_2030,N_1947,N_1918);
and U2031 (N_2031,N_1949,N_1963);
or U2032 (N_2032,N_1941,N_1921);
and U2033 (N_2033,N_1968,N_1943);
xor U2034 (N_2034,N_1960,N_1953);
xnor U2035 (N_2035,N_1957,N_1935);
and U2036 (N_2036,N_1995,N_1951);
and U2037 (N_2037,N_1961,N_1997);
nand U2038 (N_2038,N_1994,N_1981);
or U2039 (N_2039,N_1913,N_1925);
nor U2040 (N_2040,N_1996,N_1934);
and U2041 (N_2041,N_1967,N_1901);
and U2042 (N_2042,N_1940,N_1999);
xor U2043 (N_2043,N_1950,N_1978);
nand U2044 (N_2044,N_1988,N_1939);
and U2045 (N_2045,N_1982,N_1976);
nor U2046 (N_2046,N_1970,N_1974);
nor U2047 (N_2047,N_1903,N_1977);
nor U2048 (N_2048,N_1991,N_1990);
nand U2049 (N_2049,N_1945,N_1954);
and U2050 (N_2050,N_1974,N_1962);
and U2051 (N_2051,N_1968,N_1989);
xnor U2052 (N_2052,N_1988,N_1979);
nor U2053 (N_2053,N_1909,N_1959);
and U2054 (N_2054,N_1998,N_1946);
or U2055 (N_2055,N_1901,N_1980);
xnor U2056 (N_2056,N_1940,N_1926);
nor U2057 (N_2057,N_1991,N_1957);
nor U2058 (N_2058,N_1963,N_1966);
nor U2059 (N_2059,N_1936,N_1999);
xnor U2060 (N_2060,N_1968,N_1942);
and U2061 (N_2061,N_1999,N_1961);
nand U2062 (N_2062,N_1917,N_1951);
or U2063 (N_2063,N_1958,N_1944);
xnor U2064 (N_2064,N_1922,N_1966);
nor U2065 (N_2065,N_1944,N_1975);
and U2066 (N_2066,N_1914,N_1969);
or U2067 (N_2067,N_1975,N_1988);
nand U2068 (N_2068,N_1999,N_1979);
or U2069 (N_2069,N_1922,N_1941);
and U2070 (N_2070,N_1988,N_1911);
nand U2071 (N_2071,N_1950,N_1974);
nor U2072 (N_2072,N_1973,N_1964);
nand U2073 (N_2073,N_1926,N_1925);
nor U2074 (N_2074,N_1978,N_1970);
or U2075 (N_2075,N_1974,N_1927);
nor U2076 (N_2076,N_1928,N_1902);
nor U2077 (N_2077,N_1928,N_1957);
nand U2078 (N_2078,N_1994,N_1919);
nand U2079 (N_2079,N_1971,N_1903);
and U2080 (N_2080,N_1950,N_1910);
xnor U2081 (N_2081,N_1938,N_1987);
nor U2082 (N_2082,N_1952,N_1982);
or U2083 (N_2083,N_1922,N_1954);
and U2084 (N_2084,N_1924,N_1940);
nor U2085 (N_2085,N_1937,N_1911);
nand U2086 (N_2086,N_1937,N_1994);
nor U2087 (N_2087,N_1945,N_1938);
nand U2088 (N_2088,N_1920,N_1903);
or U2089 (N_2089,N_1978,N_1908);
or U2090 (N_2090,N_1988,N_1992);
nor U2091 (N_2091,N_1992,N_1974);
nor U2092 (N_2092,N_1920,N_1985);
nand U2093 (N_2093,N_1917,N_1992);
and U2094 (N_2094,N_1995,N_1918);
or U2095 (N_2095,N_1967,N_1947);
nor U2096 (N_2096,N_1932,N_1940);
nand U2097 (N_2097,N_1921,N_1964);
and U2098 (N_2098,N_1927,N_1966);
and U2099 (N_2099,N_1936,N_1946);
nand U2100 (N_2100,N_2073,N_2062);
or U2101 (N_2101,N_2008,N_2046);
nor U2102 (N_2102,N_2039,N_2069);
and U2103 (N_2103,N_2052,N_2037);
or U2104 (N_2104,N_2047,N_2089);
nor U2105 (N_2105,N_2057,N_2099);
nor U2106 (N_2106,N_2002,N_2095);
or U2107 (N_2107,N_2044,N_2049);
or U2108 (N_2108,N_2055,N_2091);
nor U2109 (N_2109,N_2019,N_2000);
and U2110 (N_2110,N_2074,N_2067);
nor U2111 (N_2111,N_2009,N_2090);
and U2112 (N_2112,N_2027,N_2093);
nand U2113 (N_2113,N_2096,N_2082);
xor U2114 (N_2114,N_2080,N_2065);
nand U2115 (N_2115,N_2066,N_2031);
or U2116 (N_2116,N_2071,N_2064);
nor U2117 (N_2117,N_2059,N_2061);
nand U2118 (N_2118,N_2075,N_2078);
nor U2119 (N_2119,N_2048,N_2021);
nand U2120 (N_2120,N_2053,N_2006);
nand U2121 (N_2121,N_2015,N_2020);
or U2122 (N_2122,N_2038,N_2013);
nand U2123 (N_2123,N_2097,N_2070);
and U2124 (N_2124,N_2088,N_2004);
nor U2125 (N_2125,N_2016,N_2017);
or U2126 (N_2126,N_2086,N_2036);
nand U2127 (N_2127,N_2072,N_2042);
and U2128 (N_2128,N_2087,N_2022);
nor U2129 (N_2129,N_2058,N_2068);
and U2130 (N_2130,N_2040,N_2032);
nand U2131 (N_2131,N_2012,N_2034);
or U2132 (N_2132,N_2084,N_2043);
xor U2133 (N_2133,N_2041,N_2001);
xnor U2134 (N_2134,N_2054,N_2007);
nand U2135 (N_2135,N_2083,N_2014);
nand U2136 (N_2136,N_2005,N_2056);
and U2137 (N_2137,N_2085,N_2033);
and U2138 (N_2138,N_2025,N_2045);
or U2139 (N_2139,N_2011,N_2003);
and U2140 (N_2140,N_2092,N_2076);
nor U2141 (N_2141,N_2063,N_2023);
or U2142 (N_2142,N_2030,N_2077);
nand U2143 (N_2143,N_2010,N_2026);
nor U2144 (N_2144,N_2098,N_2060);
or U2145 (N_2145,N_2081,N_2029);
or U2146 (N_2146,N_2024,N_2051);
nor U2147 (N_2147,N_2018,N_2079);
and U2148 (N_2148,N_2094,N_2035);
nand U2149 (N_2149,N_2028,N_2050);
nor U2150 (N_2150,N_2035,N_2068);
xor U2151 (N_2151,N_2079,N_2040);
xor U2152 (N_2152,N_2013,N_2098);
nor U2153 (N_2153,N_2089,N_2013);
nand U2154 (N_2154,N_2018,N_2044);
xnor U2155 (N_2155,N_2093,N_2085);
or U2156 (N_2156,N_2007,N_2056);
nand U2157 (N_2157,N_2051,N_2034);
nor U2158 (N_2158,N_2081,N_2028);
or U2159 (N_2159,N_2018,N_2012);
xor U2160 (N_2160,N_2085,N_2088);
xor U2161 (N_2161,N_2024,N_2003);
nand U2162 (N_2162,N_2011,N_2082);
or U2163 (N_2163,N_2053,N_2003);
nor U2164 (N_2164,N_2025,N_2000);
nand U2165 (N_2165,N_2073,N_2095);
nand U2166 (N_2166,N_2037,N_2072);
and U2167 (N_2167,N_2095,N_2032);
or U2168 (N_2168,N_2064,N_2023);
and U2169 (N_2169,N_2041,N_2084);
nor U2170 (N_2170,N_2081,N_2032);
nor U2171 (N_2171,N_2033,N_2011);
and U2172 (N_2172,N_2089,N_2075);
or U2173 (N_2173,N_2018,N_2066);
or U2174 (N_2174,N_2099,N_2014);
nand U2175 (N_2175,N_2085,N_2065);
nand U2176 (N_2176,N_2021,N_2009);
and U2177 (N_2177,N_2031,N_2059);
or U2178 (N_2178,N_2076,N_2091);
nand U2179 (N_2179,N_2061,N_2024);
nand U2180 (N_2180,N_2034,N_2038);
nand U2181 (N_2181,N_2026,N_2078);
and U2182 (N_2182,N_2084,N_2075);
xor U2183 (N_2183,N_2096,N_2067);
and U2184 (N_2184,N_2059,N_2044);
xnor U2185 (N_2185,N_2032,N_2023);
xnor U2186 (N_2186,N_2029,N_2052);
nor U2187 (N_2187,N_2013,N_2093);
nor U2188 (N_2188,N_2047,N_2053);
and U2189 (N_2189,N_2012,N_2098);
nor U2190 (N_2190,N_2008,N_2043);
and U2191 (N_2191,N_2026,N_2028);
and U2192 (N_2192,N_2021,N_2064);
or U2193 (N_2193,N_2071,N_2048);
and U2194 (N_2194,N_2004,N_2014);
or U2195 (N_2195,N_2013,N_2057);
xor U2196 (N_2196,N_2030,N_2097);
xnor U2197 (N_2197,N_2047,N_2072);
xor U2198 (N_2198,N_2058,N_2009);
or U2199 (N_2199,N_2046,N_2042);
nor U2200 (N_2200,N_2193,N_2194);
nor U2201 (N_2201,N_2184,N_2106);
and U2202 (N_2202,N_2158,N_2108);
nand U2203 (N_2203,N_2111,N_2172);
nand U2204 (N_2204,N_2154,N_2152);
nand U2205 (N_2205,N_2174,N_2143);
or U2206 (N_2206,N_2173,N_2179);
or U2207 (N_2207,N_2163,N_2162);
xnor U2208 (N_2208,N_2114,N_2121);
or U2209 (N_2209,N_2150,N_2166);
and U2210 (N_2210,N_2170,N_2120);
or U2211 (N_2211,N_2115,N_2185);
and U2212 (N_2212,N_2126,N_2125);
and U2213 (N_2213,N_2103,N_2138);
and U2214 (N_2214,N_2146,N_2104);
and U2215 (N_2215,N_2109,N_2100);
nor U2216 (N_2216,N_2130,N_2144);
or U2217 (N_2217,N_2191,N_2178);
or U2218 (N_2218,N_2189,N_2160);
nand U2219 (N_2219,N_2175,N_2105);
xnor U2220 (N_2220,N_2119,N_2140);
or U2221 (N_2221,N_2139,N_2101);
xor U2222 (N_2222,N_2192,N_2127);
nor U2223 (N_2223,N_2122,N_2168);
or U2224 (N_2224,N_2188,N_2153);
nor U2225 (N_2225,N_2181,N_2137);
and U2226 (N_2226,N_2116,N_2129);
nand U2227 (N_2227,N_2112,N_2124);
or U2228 (N_2228,N_2107,N_2157);
and U2229 (N_2229,N_2136,N_2187);
nand U2230 (N_2230,N_2180,N_2145);
or U2231 (N_2231,N_2123,N_2186);
nor U2232 (N_2232,N_2142,N_2155);
or U2233 (N_2233,N_2196,N_2156);
nor U2234 (N_2234,N_2167,N_2133);
or U2235 (N_2235,N_2161,N_2151);
xnor U2236 (N_2236,N_2131,N_2110);
nand U2237 (N_2237,N_2147,N_2190);
nand U2238 (N_2238,N_2159,N_2171);
or U2239 (N_2239,N_2198,N_2132);
and U2240 (N_2240,N_2199,N_2169);
and U2241 (N_2241,N_2118,N_2113);
or U2242 (N_2242,N_2148,N_2197);
nor U2243 (N_2243,N_2183,N_2176);
or U2244 (N_2244,N_2182,N_2165);
nor U2245 (N_2245,N_2149,N_2117);
nor U2246 (N_2246,N_2141,N_2177);
and U2247 (N_2247,N_2135,N_2164);
and U2248 (N_2248,N_2102,N_2195);
nor U2249 (N_2249,N_2134,N_2128);
or U2250 (N_2250,N_2155,N_2171);
or U2251 (N_2251,N_2175,N_2113);
xnor U2252 (N_2252,N_2125,N_2136);
nor U2253 (N_2253,N_2140,N_2149);
xnor U2254 (N_2254,N_2149,N_2199);
and U2255 (N_2255,N_2177,N_2142);
nand U2256 (N_2256,N_2113,N_2103);
and U2257 (N_2257,N_2148,N_2113);
nand U2258 (N_2258,N_2106,N_2103);
or U2259 (N_2259,N_2109,N_2106);
nor U2260 (N_2260,N_2183,N_2192);
or U2261 (N_2261,N_2156,N_2134);
xor U2262 (N_2262,N_2151,N_2169);
and U2263 (N_2263,N_2191,N_2164);
nor U2264 (N_2264,N_2107,N_2187);
nor U2265 (N_2265,N_2123,N_2195);
or U2266 (N_2266,N_2195,N_2167);
or U2267 (N_2267,N_2173,N_2161);
or U2268 (N_2268,N_2100,N_2174);
or U2269 (N_2269,N_2134,N_2108);
and U2270 (N_2270,N_2143,N_2179);
nor U2271 (N_2271,N_2124,N_2123);
nor U2272 (N_2272,N_2116,N_2190);
nor U2273 (N_2273,N_2101,N_2142);
nor U2274 (N_2274,N_2199,N_2115);
nand U2275 (N_2275,N_2148,N_2164);
nor U2276 (N_2276,N_2105,N_2112);
xor U2277 (N_2277,N_2145,N_2120);
nor U2278 (N_2278,N_2142,N_2169);
nand U2279 (N_2279,N_2184,N_2128);
xnor U2280 (N_2280,N_2187,N_2140);
nand U2281 (N_2281,N_2194,N_2187);
nor U2282 (N_2282,N_2138,N_2153);
and U2283 (N_2283,N_2105,N_2190);
nand U2284 (N_2284,N_2167,N_2152);
or U2285 (N_2285,N_2123,N_2185);
or U2286 (N_2286,N_2160,N_2140);
nor U2287 (N_2287,N_2104,N_2170);
or U2288 (N_2288,N_2165,N_2135);
or U2289 (N_2289,N_2164,N_2168);
or U2290 (N_2290,N_2177,N_2163);
nor U2291 (N_2291,N_2135,N_2101);
and U2292 (N_2292,N_2133,N_2173);
nor U2293 (N_2293,N_2191,N_2105);
nor U2294 (N_2294,N_2137,N_2140);
or U2295 (N_2295,N_2179,N_2129);
or U2296 (N_2296,N_2184,N_2141);
nor U2297 (N_2297,N_2106,N_2111);
nand U2298 (N_2298,N_2193,N_2153);
nand U2299 (N_2299,N_2151,N_2123);
nor U2300 (N_2300,N_2230,N_2244);
or U2301 (N_2301,N_2209,N_2256);
or U2302 (N_2302,N_2223,N_2236);
nand U2303 (N_2303,N_2264,N_2247);
or U2304 (N_2304,N_2219,N_2298);
nand U2305 (N_2305,N_2232,N_2281);
nor U2306 (N_2306,N_2273,N_2225);
and U2307 (N_2307,N_2278,N_2201);
and U2308 (N_2308,N_2259,N_2243);
nor U2309 (N_2309,N_2206,N_2249);
nor U2310 (N_2310,N_2242,N_2292);
xor U2311 (N_2311,N_2272,N_2258);
xor U2312 (N_2312,N_2299,N_2283);
nor U2313 (N_2313,N_2288,N_2240);
and U2314 (N_2314,N_2287,N_2245);
and U2315 (N_2315,N_2294,N_2271);
or U2316 (N_2316,N_2216,N_2285);
or U2317 (N_2317,N_2250,N_2238);
xnor U2318 (N_2318,N_2261,N_2290);
and U2319 (N_2319,N_2212,N_2215);
nand U2320 (N_2320,N_2280,N_2296);
and U2321 (N_2321,N_2295,N_2293);
and U2322 (N_2322,N_2253,N_2282);
nand U2323 (N_2323,N_2224,N_2297);
nor U2324 (N_2324,N_2233,N_2289);
or U2325 (N_2325,N_2246,N_2266);
xor U2326 (N_2326,N_2202,N_2228);
nor U2327 (N_2327,N_2252,N_2276);
xor U2328 (N_2328,N_2214,N_2265);
xor U2329 (N_2329,N_2254,N_2204);
or U2330 (N_2330,N_2213,N_2279);
or U2331 (N_2331,N_2262,N_2229);
nor U2332 (N_2332,N_2270,N_2241);
and U2333 (N_2333,N_2222,N_2248);
nor U2334 (N_2334,N_2226,N_2207);
or U2335 (N_2335,N_2274,N_2251);
or U2336 (N_2336,N_2203,N_2235);
and U2337 (N_2337,N_2239,N_2284);
nor U2338 (N_2338,N_2269,N_2231);
nor U2339 (N_2339,N_2257,N_2267);
or U2340 (N_2340,N_2275,N_2255);
and U2341 (N_2341,N_2217,N_2286);
nor U2342 (N_2342,N_2210,N_2263);
nand U2343 (N_2343,N_2221,N_2220);
and U2344 (N_2344,N_2260,N_2205);
and U2345 (N_2345,N_2237,N_2211);
nor U2346 (N_2346,N_2208,N_2200);
or U2347 (N_2347,N_2268,N_2227);
nor U2348 (N_2348,N_2234,N_2218);
nand U2349 (N_2349,N_2291,N_2277);
nand U2350 (N_2350,N_2296,N_2266);
and U2351 (N_2351,N_2289,N_2228);
or U2352 (N_2352,N_2264,N_2234);
or U2353 (N_2353,N_2230,N_2277);
or U2354 (N_2354,N_2276,N_2297);
nand U2355 (N_2355,N_2244,N_2259);
or U2356 (N_2356,N_2231,N_2242);
nand U2357 (N_2357,N_2290,N_2282);
nor U2358 (N_2358,N_2252,N_2217);
nand U2359 (N_2359,N_2216,N_2250);
nand U2360 (N_2360,N_2252,N_2296);
xnor U2361 (N_2361,N_2259,N_2211);
nand U2362 (N_2362,N_2226,N_2252);
and U2363 (N_2363,N_2209,N_2202);
nand U2364 (N_2364,N_2281,N_2276);
or U2365 (N_2365,N_2290,N_2252);
xor U2366 (N_2366,N_2233,N_2235);
nand U2367 (N_2367,N_2233,N_2236);
or U2368 (N_2368,N_2217,N_2237);
or U2369 (N_2369,N_2234,N_2222);
nand U2370 (N_2370,N_2257,N_2296);
nor U2371 (N_2371,N_2295,N_2220);
nand U2372 (N_2372,N_2282,N_2283);
nor U2373 (N_2373,N_2261,N_2286);
or U2374 (N_2374,N_2215,N_2255);
nor U2375 (N_2375,N_2297,N_2254);
or U2376 (N_2376,N_2261,N_2270);
and U2377 (N_2377,N_2295,N_2200);
nor U2378 (N_2378,N_2263,N_2297);
or U2379 (N_2379,N_2258,N_2233);
or U2380 (N_2380,N_2298,N_2225);
and U2381 (N_2381,N_2257,N_2242);
nand U2382 (N_2382,N_2262,N_2281);
xor U2383 (N_2383,N_2262,N_2288);
nand U2384 (N_2384,N_2236,N_2214);
or U2385 (N_2385,N_2203,N_2270);
nor U2386 (N_2386,N_2266,N_2283);
nand U2387 (N_2387,N_2226,N_2213);
nand U2388 (N_2388,N_2235,N_2210);
and U2389 (N_2389,N_2289,N_2287);
nor U2390 (N_2390,N_2232,N_2255);
nor U2391 (N_2391,N_2202,N_2281);
and U2392 (N_2392,N_2256,N_2255);
nor U2393 (N_2393,N_2242,N_2252);
nand U2394 (N_2394,N_2244,N_2277);
nor U2395 (N_2395,N_2220,N_2293);
and U2396 (N_2396,N_2240,N_2241);
and U2397 (N_2397,N_2287,N_2246);
and U2398 (N_2398,N_2290,N_2211);
nor U2399 (N_2399,N_2262,N_2217);
nand U2400 (N_2400,N_2352,N_2387);
nor U2401 (N_2401,N_2366,N_2309);
and U2402 (N_2402,N_2396,N_2315);
or U2403 (N_2403,N_2306,N_2314);
nand U2404 (N_2404,N_2397,N_2305);
and U2405 (N_2405,N_2361,N_2324);
and U2406 (N_2406,N_2390,N_2383);
nor U2407 (N_2407,N_2393,N_2368);
nand U2408 (N_2408,N_2320,N_2399);
nor U2409 (N_2409,N_2349,N_2338);
nor U2410 (N_2410,N_2332,N_2371);
and U2411 (N_2411,N_2374,N_2312);
and U2412 (N_2412,N_2350,N_2311);
or U2413 (N_2413,N_2355,N_2354);
nor U2414 (N_2414,N_2356,N_2313);
nor U2415 (N_2415,N_2362,N_2318);
nand U2416 (N_2416,N_2398,N_2351);
nand U2417 (N_2417,N_2385,N_2307);
nand U2418 (N_2418,N_2347,N_2346);
and U2419 (N_2419,N_2372,N_2379);
nand U2420 (N_2420,N_2384,N_2317);
and U2421 (N_2421,N_2377,N_2360);
xor U2422 (N_2422,N_2334,N_2304);
and U2423 (N_2423,N_2303,N_2331);
nand U2424 (N_2424,N_2326,N_2382);
or U2425 (N_2425,N_2359,N_2302);
or U2426 (N_2426,N_2337,N_2370);
and U2427 (N_2427,N_2380,N_2373);
nand U2428 (N_2428,N_2375,N_2358);
nand U2429 (N_2429,N_2389,N_2357);
and U2430 (N_2430,N_2369,N_2339);
nor U2431 (N_2431,N_2378,N_2322);
nand U2432 (N_2432,N_2364,N_2344);
nor U2433 (N_2433,N_2330,N_2386);
and U2434 (N_2434,N_2340,N_2308);
nor U2435 (N_2435,N_2395,N_2310);
or U2436 (N_2436,N_2321,N_2391);
nor U2437 (N_2437,N_2348,N_2392);
nor U2438 (N_2438,N_2323,N_2353);
xor U2439 (N_2439,N_2333,N_2327);
nand U2440 (N_2440,N_2328,N_2335);
nor U2441 (N_2441,N_2388,N_2329);
nor U2442 (N_2442,N_2319,N_2336);
nor U2443 (N_2443,N_2325,N_2363);
nor U2444 (N_2444,N_2367,N_2376);
nor U2445 (N_2445,N_2301,N_2365);
or U2446 (N_2446,N_2345,N_2341);
and U2447 (N_2447,N_2343,N_2394);
or U2448 (N_2448,N_2300,N_2381);
xnor U2449 (N_2449,N_2316,N_2342);
xnor U2450 (N_2450,N_2306,N_2301);
nor U2451 (N_2451,N_2309,N_2340);
nand U2452 (N_2452,N_2323,N_2330);
nor U2453 (N_2453,N_2393,N_2333);
nand U2454 (N_2454,N_2379,N_2399);
and U2455 (N_2455,N_2312,N_2379);
nand U2456 (N_2456,N_2322,N_2369);
xor U2457 (N_2457,N_2303,N_2347);
nand U2458 (N_2458,N_2348,N_2309);
and U2459 (N_2459,N_2377,N_2367);
nand U2460 (N_2460,N_2360,N_2355);
nor U2461 (N_2461,N_2389,N_2318);
and U2462 (N_2462,N_2359,N_2397);
nor U2463 (N_2463,N_2333,N_2309);
nand U2464 (N_2464,N_2334,N_2361);
nor U2465 (N_2465,N_2341,N_2376);
nand U2466 (N_2466,N_2358,N_2390);
nand U2467 (N_2467,N_2384,N_2340);
and U2468 (N_2468,N_2311,N_2327);
and U2469 (N_2469,N_2311,N_2305);
nor U2470 (N_2470,N_2351,N_2358);
xnor U2471 (N_2471,N_2341,N_2394);
and U2472 (N_2472,N_2373,N_2389);
nand U2473 (N_2473,N_2353,N_2347);
nand U2474 (N_2474,N_2393,N_2318);
xor U2475 (N_2475,N_2396,N_2342);
nand U2476 (N_2476,N_2384,N_2307);
nor U2477 (N_2477,N_2330,N_2381);
nor U2478 (N_2478,N_2312,N_2390);
and U2479 (N_2479,N_2349,N_2371);
nand U2480 (N_2480,N_2387,N_2380);
xor U2481 (N_2481,N_2363,N_2337);
nand U2482 (N_2482,N_2358,N_2364);
and U2483 (N_2483,N_2398,N_2317);
nand U2484 (N_2484,N_2353,N_2309);
xnor U2485 (N_2485,N_2319,N_2304);
nand U2486 (N_2486,N_2379,N_2361);
xor U2487 (N_2487,N_2384,N_2330);
nand U2488 (N_2488,N_2303,N_2319);
and U2489 (N_2489,N_2380,N_2321);
and U2490 (N_2490,N_2311,N_2394);
nor U2491 (N_2491,N_2352,N_2372);
nand U2492 (N_2492,N_2362,N_2363);
nor U2493 (N_2493,N_2342,N_2314);
xnor U2494 (N_2494,N_2303,N_2354);
and U2495 (N_2495,N_2313,N_2378);
and U2496 (N_2496,N_2324,N_2326);
nand U2497 (N_2497,N_2304,N_2363);
or U2498 (N_2498,N_2394,N_2331);
nand U2499 (N_2499,N_2313,N_2379);
nand U2500 (N_2500,N_2411,N_2427);
nor U2501 (N_2501,N_2424,N_2431);
and U2502 (N_2502,N_2449,N_2445);
nand U2503 (N_2503,N_2487,N_2477);
nor U2504 (N_2504,N_2484,N_2482);
nand U2505 (N_2505,N_2402,N_2466);
and U2506 (N_2506,N_2479,N_2414);
and U2507 (N_2507,N_2441,N_2444);
and U2508 (N_2508,N_2459,N_2493);
or U2509 (N_2509,N_2406,N_2475);
nor U2510 (N_2510,N_2460,N_2409);
and U2511 (N_2511,N_2405,N_2408);
xnor U2512 (N_2512,N_2426,N_2446);
nor U2513 (N_2513,N_2461,N_2462);
and U2514 (N_2514,N_2436,N_2448);
nand U2515 (N_2515,N_2472,N_2421);
or U2516 (N_2516,N_2480,N_2483);
nor U2517 (N_2517,N_2418,N_2463);
nand U2518 (N_2518,N_2455,N_2474);
nor U2519 (N_2519,N_2464,N_2439);
and U2520 (N_2520,N_2451,N_2450);
nor U2521 (N_2521,N_2440,N_2425);
nor U2522 (N_2522,N_2437,N_2417);
or U2523 (N_2523,N_2465,N_2495);
and U2524 (N_2524,N_2478,N_2412);
or U2525 (N_2525,N_2447,N_2476);
or U2526 (N_2526,N_2457,N_2467);
xor U2527 (N_2527,N_2497,N_2423);
and U2528 (N_2528,N_2415,N_2410);
and U2529 (N_2529,N_2492,N_2433);
or U2530 (N_2530,N_2420,N_2429);
or U2531 (N_2531,N_2438,N_2407);
or U2532 (N_2532,N_2453,N_2452);
xor U2533 (N_2533,N_2435,N_2471);
nor U2534 (N_2534,N_2454,N_2456);
and U2535 (N_2535,N_2486,N_2413);
nor U2536 (N_2536,N_2485,N_2498);
nor U2537 (N_2537,N_2428,N_2442);
nor U2538 (N_2538,N_2489,N_2434);
or U2539 (N_2539,N_2496,N_2422);
nor U2540 (N_2540,N_2468,N_2488);
and U2541 (N_2541,N_2490,N_2494);
or U2542 (N_2542,N_2416,N_2401);
nand U2543 (N_2543,N_2443,N_2403);
nor U2544 (N_2544,N_2430,N_2481);
or U2545 (N_2545,N_2469,N_2400);
nor U2546 (N_2546,N_2499,N_2458);
or U2547 (N_2547,N_2470,N_2404);
xor U2548 (N_2548,N_2419,N_2491);
nor U2549 (N_2549,N_2432,N_2473);
nor U2550 (N_2550,N_2476,N_2498);
and U2551 (N_2551,N_2471,N_2420);
and U2552 (N_2552,N_2498,N_2481);
nand U2553 (N_2553,N_2431,N_2461);
nor U2554 (N_2554,N_2477,N_2462);
xnor U2555 (N_2555,N_2417,N_2484);
or U2556 (N_2556,N_2406,N_2400);
and U2557 (N_2557,N_2471,N_2411);
or U2558 (N_2558,N_2491,N_2470);
or U2559 (N_2559,N_2449,N_2476);
or U2560 (N_2560,N_2412,N_2436);
nand U2561 (N_2561,N_2473,N_2407);
and U2562 (N_2562,N_2404,N_2448);
nor U2563 (N_2563,N_2474,N_2454);
nor U2564 (N_2564,N_2406,N_2483);
nor U2565 (N_2565,N_2458,N_2481);
nor U2566 (N_2566,N_2458,N_2448);
nand U2567 (N_2567,N_2482,N_2420);
nor U2568 (N_2568,N_2457,N_2414);
and U2569 (N_2569,N_2476,N_2461);
or U2570 (N_2570,N_2413,N_2406);
nor U2571 (N_2571,N_2423,N_2471);
nand U2572 (N_2572,N_2477,N_2408);
nand U2573 (N_2573,N_2434,N_2494);
xnor U2574 (N_2574,N_2468,N_2478);
and U2575 (N_2575,N_2475,N_2427);
nor U2576 (N_2576,N_2475,N_2497);
or U2577 (N_2577,N_2400,N_2412);
nor U2578 (N_2578,N_2416,N_2422);
nor U2579 (N_2579,N_2429,N_2406);
and U2580 (N_2580,N_2495,N_2433);
nor U2581 (N_2581,N_2471,N_2493);
and U2582 (N_2582,N_2461,N_2425);
nor U2583 (N_2583,N_2446,N_2490);
nor U2584 (N_2584,N_2405,N_2473);
nor U2585 (N_2585,N_2448,N_2476);
nor U2586 (N_2586,N_2481,N_2416);
nand U2587 (N_2587,N_2475,N_2428);
nand U2588 (N_2588,N_2411,N_2447);
nor U2589 (N_2589,N_2437,N_2407);
xor U2590 (N_2590,N_2409,N_2402);
nand U2591 (N_2591,N_2494,N_2438);
and U2592 (N_2592,N_2401,N_2438);
or U2593 (N_2593,N_2458,N_2401);
nand U2594 (N_2594,N_2405,N_2429);
and U2595 (N_2595,N_2403,N_2483);
nand U2596 (N_2596,N_2474,N_2486);
nand U2597 (N_2597,N_2463,N_2493);
nand U2598 (N_2598,N_2452,N_2413);
nand U2599 (N_2599,N_2484,N_2403);
or U2600 (N_2600,N_2543,N_2509);
nand U2601 (N_2601,N_2564,N_2549);
and U2602 (N_2602,N_2541,N_2532);
nor U2603 (N_2603,N_2570,N_2517);
or U2604 (N_2604,N_2513,N_2561);
or U2605 (N_2605,N_2544,N_2523);
or U2606 (N_2606,N_2585,N_2508);
nand U2607 (N_2607,N_2507,N_2581);
or U2608 (N_2608,N_2522,N_2547);
or U2609 (N_2609,N_2559,N_2557);
nor U2610 (N_2610,N_2597,N_2575);
or U2611 (N_2611,N_2537,N_2563);
and U2612 (N_2612,N_2589,N_2566);
nor U2613 (N_2613,N_2568,N_2586);
and U2614 (N_2614,N_2594,N_2503);
nand U2615 (N_2615,N_2593,N_2501);
and U2616 (N_2616,N_2584,N_2558);
nand U2617 (N_2617,N_2536,N_2542);
and U2618 (N_2618,N_2520,N_2550);
and U2619 (N_2619,N_2518,N_2562);
and U2620 (N_2620,N_2506,N_2515);
nor U2621 (N_2621,N_2530,N_2592);
nand U2622 (N_2622,N_2526,N_2546);
and U2623 (N_2623,N_2529,N_2553);
and U2624 (N_2624,N_2582,N_2580);
nor U2625 (N_2625,N_2502,N_2527);
xor U2626 (N_2626,N_2505,N_2521);
and U2627 (N_2627,N_2514,N_2510);
xnor U2628 (N_2628,N_2595,N_2555);
xor U2629 (N_2629,N_2578,N_2590);
or U2630 (N_2630,N_2511,N_2519);
nor U2631 (N_2631,N_2504,N_2571);
or U2632 (N_2632,N_2567,N_2533);
nor U2633 (N_2633,N_2596,N_2569);
nand U2634 (N_2634,N_2556,N_2528);
nand U2635 (N_2635,N_2560,N_2539);
and U2636 (N_2636,N_2587,N_2534);
and U2637 (N_2637,N_2525,N_2599);
nand U2638 (N_2638,N_2588,N_2540);
and U2639 (N_2639,N_2573,N_2512);
nand U2640 (N_2640,N_2576,N_2552);
nor U2641 (N_2641,N_2577,N_2598);
or U2642 (N_2642,N_2572,N_2579);
or U2643 (N_2643,N_2535,N_2554);
and U2644 (N_2644,N_2548,N_2538);
xor U2645 (N_2645,N_2583,N_2531);
nor U2646 (N_2646,N_2591,N_2524);
nand U2647 (N_2647,N_2565,N_2545);
nand U2648 (N_2648,N_2516,N_2500);
and U2649 (N_2649,N_2574,N_2551);
nor U2650 (N_2650,N_2599,N_2554);
and U2651 (N_2651,N_2527,N_2587);
xor U2652 (N_2652,N_2504,N_2513);
and U2653 (N_2653,N_2559,N_2525);
nor U2654 (N_2654,N_2524,N_2554);
nor U2655 (N_2655,N_2545,N_2547);
nand U2656 (N_2656,N_2599,N_2560);
or U2657 (N_2657,N_2516,N_2517);
and U2658 (N_2658,N_2567,N_2549);
xnor U2659 (N_2659,N_2558,N_2536);
or U2660 (N_2660,N_2550,N_2573);
and U2661 (N_2661,N_2527,N_2507);
or U2662 (N_2662,N_2554,N_2529);
nand U2663 (N_2663,N_2562,N_2523);
nand U2664 (N_2664,N_2588,N_2536);
or U2665 (N_2665,N_2506,N_2585);
and U2666 (N_2666,N_2597,N_2593);
or U2667 (N_2667,N_2555,N_2538);
nand U2668 (N_2668,N_2538,N_2510);
and U2669 (N_2669,N_2516,N_2539);
nand U2670 (N_2670,N_2547,N_2533);
and U2671 (N_2671,N_2534,N_2545);
and U2672 (N_2672,N_2530,N_2519);
or U2673 (N_2673,N_2592,N_2563);
nand U2674 (N_2674,N_2580,N_2591);
or U2675 (N_2675,N_2569,N_2510);
and U2676 (N_2676,N_2557,N_2585);
or U2677 (N_2677,N_2511,N_2588);
and U2678 (N_2678,N_2596,N_2508);
xor U2679 (N_2679,N_2510,N_2553);
nand U2680 (N_2680,N_2525,N_2537);
or U2681 (N_2681,N_2586,N_2557);
nor U2682 (N_2682,N_2514,N_2590);
and U2683 (N_2683,N_2565,N_2528);
nand U2684 (N_2684,N_2580,N_2547);
nand U2685 (N_2685,N_2580,N_2550);
and U2686 (N_2686,N_2563,N_2530);
nor U2687 (N_2687,N_2535,N_2521);
or U2688 (N_2688,N_2544,N_2533);
xor U2689 (N_2689,N_2538,N_2518);
nor U2690 (N_2690,N_2557,N_2564);
nor U2691 (N_2691,N_2535,N_2576);
and U2692 (N_2692,N_2574,N_2580);
or U2693 (N_2693,N_2578,N_2591);
xnor U2694 (N_2694,N_2532,N_2581);
nand U2695 (N_2695,N_2571,N_2584);
and U2696 (N_2696,N_2566,N_2507);
and U2697 (N_2697,N_2569,N_2520);
nand U2698 (N_2698,N_2577,N_2568);
xor U2699 (N_2699,N_2537,N_2552);
and U2700 (N_2700,N_2603,N_2608);
or U2701 (N_2701,N_2611,N_2653);
or U2702 (N_2702,N_2699,N_2654);
or U2703 (N_2703,N_2680,N_2630);
or U2704 (N_2704,N_2660,N_2614);
or U2705 (N_2705,N_2617,N_2639);
nand U2706 (N_2706,N_2649,N_2656);
nand U2707 (N_2707,N_2663,N_2685);
nor U2708 (N_2708,N_2691,N_2675);
nand U2709 (N_2709,N_2693,N_2665);
nand U2710 (N_2710,N_2686,N_2633);
xnor U2711 (N_2711,N_2625,N_2668);
or U2712 (N_2712,N_2616,N_2601);
and U2713 (N_2713,N_2610,N_2677);
and U2714 (N_2714,N_2689,N_2658);
or U2715 (N_2715,N_2635,N_2607);
nand U2716 (N_2716,N_2673,N_2672);
nor U2717 (N_2717,N_2666,N_2690);
and U2718 (N_2718,N_2688,N_2604);
nand U2719 (N_2719,N_2657,N_2609);
xnor U2720 (N_2720,N_2619,N_2659);
and U2721 (N_2721,N_2618,N_2683);
or U2722 (N_2722,N_2632,N_2652);
nand U2723 (N_2723,N_2645,N_2692);
nand U2724 (N_2724,N_2687,N_2637);
and U2725 (N_2725,N_2651,N_2621);
nand U2726 (N_2726,N_2600,N_2642);
xor U2727 (N_2727,N_2634,N_2602);
and U2728 (N_2728,N_2647,N_2676);
and U2729 (N_2729,N_2682,N_2644);
nand U2730 (N_2730,N_2674,N_2629);
and U2731 (N_2731,N_2641,N_2650);
or U2732 (N_2732,N_2636,N_2643);
nor U2733 (N_2733,N_2667,N_2679);
nand U2734 (N_2734,N_2661,N_2613);
and U2735 (N_2735,N_2624,N_2626);
xor U2736 (N_2736,N_2605,N_2678);
and U2737 (N_2737,N_2646,N_2648);
nand U2738 (N_2738,N_2696,N_2664);
and U2739 (N_2739,N_2615,N_2627);
or U2740 (N_2740,N_2671,N_2620);
nor U2741 (N_2741,N_2681,N_2622);
nor U2742 (N_2742,N_2640,N_2606);
nor U2743 (N_2743,N_2638,N_2612);
xor U2744 (N_2744,N_2695,N_2655);
xnor U2745 (N_2745,N_2662,N_2628);
nand U2746 (N_2746,N_2670,N_2623);
and U2747 (N_2747,N_2631,N_2694);
or U2748 (N_2748,N_2697,N_2669);
nor U2749 (N_2749,N_2698,N_2684);
nor U2750 (N_2750,N_2674,N_2665);
nand U2751 (N_2751,N_2678,N_2667);
nor U2752 (N_2752,N_2606,N_2634);
and U2753 (N_2753,N_2661,N_2624);
and U2754 (N_2754,N_2692,N_2696);
nand U2755 (N_2755,N_2636,N_2664);
nor U2756 (N_2756,N_2611,N_2616);
nand U2757 (N_2757,N_2665,N_2606);
nand U2758 (N_2758,N_2610,N_2607);
or U2759 (N_2759,N_2602,N_2685);
nand U2760 (N_2760,N_2648,N_2602);
and U2761 (N_2761,N_2678,N_2660);
nand U2762 (N_2762,N_2624,N_2637);
and U2763 (N_2763,N_2659,N_2620);
nand U2764 (N_2764,N_2655,N_2638);
xnor U2765 (N_2765,N_2699,N_2630);
and U2766 (N_2766,N_2644,N_2603);
and U2767 (N_2767,N_2667,N_2697);
or U2768 (N_2768,N_2658,N_2630);
nand U2769 (N_2769,N_2603,N_2696);
nor U2770 (N_2770,N_2611,N_2670);
nor U2771 (N_2771,N_2621,N_2658);
xor U2772 (N_2772,N_2606,N_2659);
nor U2773 (N_2773,N_2651,N_2671);
nor U2774 (N_2774,N_2693,N_2646);
nand U2775 (N_2775,N_2614,N_2641);
or U2776 (N_2776,N_2620,N_2627);
and U2777 (N_2777,N_2660,N_2624);
and U2778 (N_2778,N_2662,N_2690);
xor U2779 (N_2779,N_2647,N_2677);
nor U2780 (N_2780,N_2630,N_2666);
and U2781 (N_2781,N_2674,N_2675);
nand U2782 (N_2782,N_2610,N_2686);
nor U2783 (N_2783,N_2625,N_2671);
or U2784 (N_2784,N_2687,N_2678);
xor U2785 (N_2785,N_2683,N_2626);
and U2786 (N_2786,N_2603,N_2688);
and U2787 (N_2787,N_2617,N_2682);
or U2788 (N_2788,N_2635,N_2661);
or U2789 (N_2789,N_2633,N_2673);
nor U2790 (N_2790,N_2659,N_2677);
and U2791 (N_2791,N_2610,N_2646);
nor U2792 (N_2792,N_2622,N_2639);
nor U2793 (N_2793,N_2688,N_2677);
nor U2794 (N_2794,N_2665,N_2692);
nand U2795 (N_2795,N_2626,N_2635);
and U2796 (N_2796,N_2641,N_2680);
or U2797 (N_2797,N_2621,N_2654);
and U2798 (N_2798,N_2601,N_2670);
or U2799 (N_2799,N_2627,N_2689);
or U2800 (N_2800,N_2796,N_2791);
nand U2801 (N_2801,N_2759,N_2782);
nor U2802 (N_2802,N_2764,N_2752);
or U2803 (N_2803,N_2776,N_2712);
or U2804 (N_2804,N_2738,N_2792);
nor U2805 (N_2805,N_2773,N_2727);
nor U2806 (N_2806,N_2733,N_2728);
nand U2807 (N_2807,N_2704,N_2762);
nand U2808 (N_2808,N_2731,N_2797);
nand U2809 (N_2809,N_2793,N_2730);
or U2810 (N_2810,N_2732,N_2789);
or U2811 (N_2811,N_2736,N_2735);
and U2812 (N_2812,N_2780,N_2765);
nand U2813 (N_2813,N_2768,N_2778);
and U2814 (N_2814,N_2723,N_2749);
or U2815 (N_2815,N_2794,N_2705);
or U2816 (N_2816,N_2743,N_2726);
and U2817 (N_2817,N_2758,N_2729);
or U2818 (N_2818,N_2700,N_2717);
nand U2819 (N_2819,N_2706,N_2741);
nand U2820 (N_2820,N_2719,N_2721);
nor U2821 (N_2821,N_2737,N_2787);
nor U2822 (N_2822,N_2784,N_2724);
nor U2823 (N_2823,N_2748,N_2750);
nand U2824 (N_2824,N_2771,N_2769);
or U2825 (N_2825,N_2775,N_2740);
and U2826 (N_2826,N_2798,N_2746);
xnor U2827 (N_2827,N_2744,N_2799);
or U2828 (N_2828,N_2707,N_2763);
nand U2829 (N_2829,N_2720,N_2722);
xor U2830 (N_2830,N_2790,N_2751);
and U2831 (N_2831,N_2783,N_2777);
or U2832 (N_2832,N_2755,N_2788);
and U2833 (N_2833,N_2718,N_2761);
or U2834 (N_2834,N_2715,N_2754);
xnor U2835 (N_2835,N_2753,N_2795);
nor U2836 (N_2836,N_2702,N_2714);
nor U2837 (N_2837,N_2785,N_2711);
nand U2838 (N_2838,N_2766,N_2725);
xnor U2839 (N_2839,N_2716,N_2703);
and U2840 (N_2840,N_2757,N_2760);
or U2841 (N_2841,N_2713,N_2739);
nand U2842 (N_2842,N_2708,N_2734);
or U2843 (N_2843,N_2774,N_2747);
nand U2844 (N_2844,N_2770,N_2709);
nor U2845 (N_2845,N_2772,N_2756);
and U2846 (N_2846,N_2710,N_2779);
xor U2847 (N_2847,N_2745,N_2742);
nor U2848 (N_2848,N_2767,N_2781);
nand U2849 (N_2849,N_2786,N_2701);
nand U2850 (N_2850,N_2742,N_2774);
and U2851 (N_2851,N_2725,N_2746);
and U2852 (N_2852,N_2785,N_2775);
xnor U2853 (N_2853,N_2733,N_2794);
xnor U2854 (N_2854,N_2735,N_2710);
and U2855 (N_2855,N_2742,N_2778);
or U2856 (N_2856,N_2702,N_2733);
or U2857 (N_2857,N_2783,N_2798);
nand U2858 (N_2858,N_2717,N_2787);
nand U2859 (N_2859,N_2793,N_2776);
or U2860 (N_2860,N_2781,N_2796);
nor U2861 (N_2861,N_2760,N_2747);
or U2862 (N_2862,N_2719,N_2747);
xor U2863 (N_2863,N_2789,N_2707);
nor U2864 (N_2864,N_2703,N_2763);
and U2865 (N_2865,N_2775,N_2764);
nor U2866 (N_2866,N_2705,N_2716);
nand U2867 (N_2867,N_2764,N_2750);
nand U2868 (N_2868,N_2795,N_2731);
and U2869 (N_2869,N_2742,N_2708);
or U2870 (N_2870,N_2781,N_2779);
xnor U2871 (N_2871,N_2736,N_2747);
or U2872 (N_2872,N_2772,N_2776);
nor U2873 (N_2873,N_2765,N_2724);
or U2874 (N_2874,N_2709,N_2749);
nand U2875 (N_2875,N_2716,N_2704);
and U2876 (N_2876,N_2723,N_2772);
and U2877 (N_2877,N_2777,N_2704);
or U2878 (N_2878,N_2789,N_2709);
nand U2879 (N_2879,N_2726,N_2704);
or U2880 (N_2880,N_2719,N_2756);
nand U2881 (N_2881,N_2726,N_2701);
or U2882 (N_2882,N_2788,N_2702);
or U2883 (N_2883,N_2710,N_2796);
xor U2884 (N_2884,N_2744,N_2746);
nand U2885 (N_2885,N_2757,N_2797);
or U2886 (N_2886,N_2793,N_2791);
and U2887 (N_2887,N_2740,N_2748);
and U2888 (N_2888,N_2762,N_2755);
and U2889 (N_2889,N_2757,N_2778);
or U2890 (N_2890,N_2778,N_2765);
xnor U2891 (N_2891,N_2792,N_2770);
and U2892 (N_2892,N_2796,N_2738);
and U2893 (N_2893,N_2774,N_2717);
and U2894 (N_2894,N_2787,N_2782);
and U2895 (N_2895,N_2790,N_2781);
nand U2896 (N_2896,N_2790,N_2716);
nand U2897 (N_2897,N_2748,N_2780);
nand U2898 (N_2898,N_2719,N_2735);
nor U2899 (N_2899,N_2707,N_2738);
nor U2900 (N_2900,N_2883,N_2881);
nand U2901 (N_2901,N_2818,N_2819);
nor U2902 (N_2902,N_2805,N_2873);
xor U2903 (N_2903,N_2884,N_2821);
nand U2904 (N_2904,N_2872,N_2886);
or U2905 (N_2905,N_2844,N_2861);
or U2906 (N_2906,N_2870,N_2849);
xor U2907 (N_2907,N_2828,N_2874);
nand U2908 (N_2908,N_2838,N_2864);
nor U2909 (N_2909,N_2803,N_2880);
nand U2910 (N_2910,N_2800,N_2890);
or U2911 (N_2911,N_2846,N_2895);
nor U2912 (N_2912,N_2852,N_2858);
xnor U2913 (N_2913,N_2871,N_2885);
and U2914 (N_2914,N_2859,N_2866);
xnor U2915 (N_2915,N_2837,N_2845);
xnor U2916 (N_2916,N_2835,N_2831);
nand U2917 (N_2917,N_2812,N_2817);
nor U2918 (N_2918,N_2834,N_2876);
or U2919 (N_2919,N_2836,N_2810);
nand U2920 (N_2920,N_2868,N_2877);
nand U2921 (N_2921,N_2894,N_2804);
and U2922 (N_2922,N_2813,N_2891);
and U2923 (N_2923,N_2825,N_2892);
xor U2924 (N_2924,N_2887,N_2879);
and U2925 (N_2925,N_2814,N_2832);
or U2926 (N_2926,N_2878,N_2897);
nand U2927 (N_2927,N_2851,N_2824);
nor U2928 (N_2928,N_2839,N_2860);
and U2929 (N_2929,N_2842,N_2815);
or U2930 (N_2930,N_2869,N_2809);
nor U2931 (N_2931,N_2833,N_2830);
and U2932 (N_2932,N_2857,N_2855);
nand U2933 (N_2933,N_2862,N_2827);
nand U2934 (N_2934,N_2898,N_2811);
and U2935 (N_2935,N_2826,N_2802);
or U2936 (N_2936,N_2840,N_2841);
nand U2937 (N_2937,N_2816,N_2865);
xor U2938 (N_2938,N_2893,N_2806);
nand U2939 (N_2939,N_2854,N_2856);
nand U2940 (N_2940,N_2808,N_2899);
xor U2941 (N_2941,N_2875,N_2843);
nand U2942 (N_2942,N_2807,N_2863);
nand U2943 (N_2943,N_2822,N_2896);
and U2944 (N_2944,N_2829,N_2882);
or U2945 (N_2945,N_2850,N_2801);
and U2946 (N_2946,N_2853,N_2889);
xnor U2947 (N_2947,N_2820,N_2888);
nor U2948 (N_2948,N_2867,N_2847);
or U2949 (N_2949,N_2848,N_2823);
xor U2950 (N_2950,N_2810,N_2808);
nand U2951 (N_2951,N_2825,N_2887);
and U2952 (N_2952,N_2896,N_2836);
nor U2953 (N_2953,N_2849,N_2888);
or U2954 (N_2954,N_2885,N_2899);
or U2955 (N_2955,N_2891,N_2877);
xor U2956 (N_2956,N_2893,N_2844);
xor U2957 (N_2957,N_2896,N_2862);
xnor U2958 (N_2958,N_2823,N_2820);
nor U2959 (N_2959,N_2841,N_2856);
xor U2960 (N_2960,N_2847,N_2881);
and U2961 (N_2961,N_2855,N_2853);
nand U2962 (N_2962,N_2886,N_2830);
nor U2963 (N_2963,N_2824,N_2880);
or U2964 (N_2964,N_2846,N_2825);
and U2965 (N_2965,N_2817,N_2877);
or U2966 (N_2966,N_2828,N_2885);
nor U2967 (N_2967,N_2898,N_2848);
nor U2968 (N_2968,N_2865,N_2817);
and U2969 (N_2969,N_2899,N_2810);
nand U2970 (N_2970,N_2828,N_2871);
nand U2971 (N_2971,N_2874,N_2816);
and U2972 (N_2972,N_2842,N_2841);
nor U2973 (N_2973,N_2821,N_2866);
nor U2974 (N_2974,N_2853,N_2893);
xor U2975 (N_2975,N_2892,N_2808);
and U2976 (N_2976,N_2840,N_2846);
xor U2977 (N_2977,N_2842,N_2851);
xnor U2978 (N_2978,N_2849,N_2832);
nand U2979 (N_2979,N_2809,N_2847);
or U2980 (N_2980,N_2833,N_2876);
or U2981 (N_2981,N_2848,N_2814);
nand U2982 (N_2982,N_2843,N_2840);
and U2983 (N_2983,N_2833,N_2807);
nor U2984 (N_2984,N_2811,N_2813);
nor U2985 (N_2985,N_2885,N_2876);
nor U2986 (N_2986,N_2871,N_2893);
or U2987 (N_2987,N_2882,N_2855);
and U2988 (N_2988,N_2834,N_2883);
nand U2989 (N_2989,N_2899,N_2827);
nand U2990 (N_2990,N_2816,N_2854);
nand U2991 (N_2991,N_2853,N_2898);
nand U2992 (N_2992,N_2827,N_2838);
or U2993 (N_2993,N_2843,N_2825);
nand U2994 (N_2994,N_2823,N_2870);
or U2995 (N_2995,N_2873,N_2890);
xor U2996 (N_2996,N_2876,N_2810);
nor U2997 (N_2997,N_2820,N_2827);
nor U2998 (N_2998,N_2862,N_2832);
nor U2999 (N_2999,N_2808,N_2825);
nor UO_0 (O_0,N_2986,N_2911);
nor UO_1 (O_1,N_2900,N_2958);
xnor UO_2 (O_2,N_2972,N_2977);
nand UO_3 (O_3,N_2935,N_2988);
and UO_4 (O_4,N_2980,N_2982);
xnor UO_5 (O_5,N_2959,N_2952);
nor UO_6 (O_6,N_2918,N_2995);
nand UO_7 (O_7,N_2954,N_2998);
and UO_8 (O_8,N_2910,N_2932);
xnor UO_9 (O_9,N_2909,N_2926);
and UO_10 (O_10,N_2956,N_2921);
nand UO_11 (O_11,N_2936,N_2940);
and UO_12 (O_12,N_2937,N_2924);
or UO_13 (O_13,N_2922,N_2925);
nor UO_14 (O_14,N_2917,N_2965);
or UO_15 (O_15,N_2974,N_2930);
or UO_16 (O_16,N_2951,N_2913);
nor UO_17 (O_17,N_2978,N_2994);
or UO_18 (O_18,N_2915,N_2955);
xnor UO_19 (O_19,N_2989,N_2999);
and UO_20 (O_20,N_2902,N_2961);
nand UO_21 (O_21,N_2945,N_2985);
or UO_22 (O_22,N_2969,N_2981);
or UO_23 (O_23,N_2967,N_2953);
or UO_24 (O_24,N_2905,N_2957);
nand UO_25 (O_25,N_2928,N_2997);
and UO_26 (O_26,N_2923,N_2971);
or UO_27 (O_27,N_2914,N_2903);
nor UO_28 (O_28,N_2919,N_2983);
nor UO_29 (O_29,N_2963,N_2966);
and UO_30 (O_30,N_2973,N_2907);
or UO_31 (O_31,N_2934,N_2976);
or UO_32 (O_32,N_2979,N_2927);
and UO_33 (O_33,N_2947,N_2964);
nand UO_34 (O_34,N_2991,N_2949);
and UO_35 (O_35,N_2996,N_2933);
or UO_36 (O_36,N_2938,N_2992);
nor UO_37 (O_37,N_2943,N_2939);
and UO_38 (O_38,N_2942,N_2904);
nor UO_39 (O_39,N_2950,N_2912);
xnor UO_40 (O_40,N_2929,N_2987);
nor UO_41 (O_41,N_2984,N_2946);
and UO_42 (O_42,N_2906,N_2944);
and UO_43 (O_43,N_2908,N_2941);
and UO_44 (O_44,N_2960,N_2975);
nor UO_45 (O_45,N_2968,N_2948);
or UO_46 (O_46,N_2901,N_2916);
nor UO_47 (O_47,N_2962,N_2990);
nand UO_48 (O_48,N_2920,N_2931);
nor UO_49 (O_49,N_2993,N_2970);
nor UO_50 (O_50,N_2965,N_2900);
nand UO_51 (O_51,N_2929,N_2913);
or UO_52 (O_52,N_2970,N_2939);
nor UO_53 (O_53,N_2964,N_2968);
nand UO_54 (O_54,N_2908,N_2910);
nand UO_55 (O_55,N_2941,N_2998);
nand UO_56 (O_56,N_2924,N_2941);
nand UO_57 (O_57,N_2997,N_2956);
and UO_58 (O_58,N_2950,N_2932);
nor UO_59 (O_59,N_2993,N_2948);
or UO_60 (O_60,N_2960,N_2982);
or UO_61 (O_61,N_2992,N_2964);
nor UO_62 (O_62,N_2949,N_2904);
or UO_63 (O_63,N_2959,N_2906);
nand UO_64 (O_64,N_2957,N_2909);
nor UO_65 (O_65,N_2911,N_2967);
nand UO_66 (O_66,N_2936,N_2950);
xor UO_67 (O_67,N_2989,N_2926);
nand UO_68 (O_68,N_2912,N_2919);
nand UO_69 (O_69,N_2920,N_2911);
nor UO_70 (O_70,N_2991,N_2912);
or UO_71 (O_71,N_2983,N_2959);
nand UO_72 (O_72,N_2932,N_2962);
nor UO_73 (O_73,N_2970,N_2983);
nand UO_74 (O_74,N_2924,N_2956);
nand UO_75 (O_75,N_2911,N_2970);
nor UO_76 (O_76,N_2977,N_2999);
and UO_77 (O_77,N_2904,N_2905);
and UO_78 (O_78,N_2916,N_2967);
nor UO_79 (O_79,N_2937,N_2967);
and UO_80 (O_80,N_2913,N_2957);
nor UO_81 (O_81,N_2977,N_2937);
or UO_82 (O_82,N_2984,N_2927);
nor UO_83 (O_83,N_2925,N_2953);
nor UO_84 (O_84,N_2957,N_2944);
or UO_85 (O_85,N_2916,N_2900);
and UO_86 (O_86,N_2969,N_2973);
and UO_87 (O_87,N_2932,N_2975);
xor UO_88 (O_88,N_2991,N_2948);
xnor UO_89 (O_89,N_2925,N_2971);
nand UO_90 (O_90,N_2904,N_2979);
and UO_91 (O_91,N_2940,N_2992);
and UO_92 (O_92,N_2959,N_2909);
and UO_93 (O_93,N_2947,N_2941);
nor UO_94 (O_94,N_2914,N_2915);
and UO_95 (O_95,N_2921,N_2995);
and UO_96 (O_96,N_2997,N_2989);
nand UO_97 (O_97,N_2934,N_2945);
nor UO_98 (O_98,N_2918,N_2993);
and UO_99 (O_99,N_2989,N_2967);
nand UO_100 (O_100,N_2983,N_2967);
nand UO_101 (O_101,N_2986,N_2995);
xnor UO_102 (O_102,N_2940,N_2915);
xnor UO_103 (O_103,N_2969,N_2915);
and UO_104 (O_104,N_2995,N_2901);
or UO_105 (O_105,N_2976,N_2931);
nor UO_106 (O_106,N_2952,N_2945);
or UO_107 (O_107,N_2967,N_2905);
and UO_108 (O_108,N_2986,N_2924);
nand UO_109 (O_109,N_2925,N_2937);
or UO_110 (O_110,N_2993,N_2994);
nor UO_111 (O_111,N_2960,N_2976);
nand UO_112 (O_112,N_2958,N_2908);
xor UO_113 (O_113,N_2968,N_2931);
or UO_114 (O_114,N_2935,N_2933);
xor UO_115 (O_115,N_2912,N_2924);
nand UO_116 (O_116,N_2903,N_2930);
nor UO_117 (O_117,N_2992,N_2934);
xnor UO_118 (O_118,N_2944,N_2918);
nor UO_119 (O_119,N_2988,N_2998);
nor UO_120 (O_120,N_2928,N_2948);
or UO_121 (O_121,N_2982,N_2903);
or UO_122 (O_122,N_2997,N_2970);
xnor UO_123 (O_123,N_2905,N_2919);
or UO_124 (O_124,N_2917,N_2915);
nor UO_125 (O_125,N_2950,N_2945);
nor UO_126 (O_126,N_2959,N_2915);
nand UO_127 (O_127,N_2936,N_2998);
nor UO_128 (O_128,N_2978,N_2905);
and UO_129 (O_129,N_2977,N_2933);
nand UO_130 (O_130,N_2922,N_2975);
nor UO_131 (O_131,N_2948,N_2910);
or UO_132 (O_132,N_2959,N_2929);
nor UO_133 (O_133,N_2929,N_2980);
nand UO_134 (O_134,N_2963,N_2943);
xnor UO_135 (O_135,N_2978,N_2984);
or UO_136 (O_136,N_2931,N_2921);
nand UO_137 (O_137,N_2927,N_2987);
and UO_138 (O_138,N_2919,N_2962);
and UO_139 (O_139,N_2965,N_2937);
nor UO_140 (O_140,N_2921,N_2936);
or UO_141 (O_141,N_2984,N_2902);
xor UO_142 (O_142,N_2981,N_2900);
nor UO_143 (O_143,N_2937,N_2985);
or UO_144 (O_144,N_2967,N_2919);
xnor UO_145 (O_145,N_2903,N_2977);
nand UO_146 (O_146,N_2930,N_2918);
nor UO_147 (O_147,N_2926,N_2986);
nand UO_148 (O_148,N_2938,N_2950);
nor UO_149 (O_149,N_2922,N_2984);
xnor UO_150 (O_150,N_2941,N_2913);
and UO_151 (O_151,N_2998,N_2917);
nand UO_152 (O_152,N_2908,N_2921);
nand UO_153 (O_153,N_2945,N_2964);
nand UO_154 (O_154,N_2902,N_2978);
nand UO_155 (O_155,N_2967,N_2955);
nand UO_156 (O_156,N_2926,N_2959);
xnor UO_157 (O_157,N_2966,N_2908);
xor UO_158 (O_158,N_2953,N_2960);
nand UO_159 (O_159,N_2994,N_2961);
nand UO_160 (O_160,N_2918,N_2973);
nor UO_161 (O_161,N_2940,N_2957);
nand UO_162 (O_162,N_2922,N_2969);
nor UO_163 (O_163,N_2940,N_2978);
nand UO_164 (O_164,N_2990,N_2933);
and UO_165 (O_165,N_2965,N_2939);
or UO_166 (O_166,N_2917,N_2972);
and UO_167 (O_167,N_2945,N_2970);
or UO_168 (O_168,N_2917,N_2928);
and UO_169 (O_169,N_2929,N_2955);
and UO_170 (O_170,N_2983,N_2963);
and UO_171 (O_171,N_2984,N_2989);
or UO_172 (O_172,N_2914,N_2958);
nand UO_173 (O_173,N_2917,N_2975);
and UO_174 (O_174,N_2962,N_2904);
or UO_175 (O_175,N_2972,N_2966);
nand UO_176 (O_176,N_2952,N_2956);
nand UO_177 (O_177,N_2917,N_2957);
or UO_178 (O_178,N_2969,N_2918);
nor UO_179 (O_179,N_2979,N_2966);
and UO_180 (O_180,N_2972,N_2985);
nand UO_181 (O_181,N_2936,N_2900);
nor UO_182 (O_182,N_2923,N_2981);
or UO_183 (O_183,N_2962,N_2922);
and UO_184 (O_184,N_2993,N_2904);
nand UO_185 (O_185,N_2940,N_2949);
xnor UO_186 (O_186,N_2902,N_2982);
xor UO_187 (O_187,N_2901,N_2917);
and UO_188 (O_188,N_2953,N_2976);
and UO_189 (O_189,N_2936,N_2926);
and UO_190 (O_190,N_2982,N_2923);
nand UO_191 (O_191,N_2999,N_2968);
nor UO_192 (O_192,N_2951,N_2995);
nor UO_193 (O_193,N_2942,N_2966);
nand UO_194 (O_194,N_2978,N_2937);
xor UO_195 (O_195,N_2920,N_2961);
or UO_196 (O_196,N_2992,N_2996);
and UO_197 (O_197,N_2939,N_2953);
nor UO_198 (O_198,N_2941,N_2914);
nand UO_199 (O_199,N_2984,N_2996);
nor UO_200 (O_200,N_2938,N_2975);
nand UO_201 (O_201,N_2971,N_2966);
xnor UO_202 (O_202,N_2950,N_2962);
nor UO_203 (O_203,N_2960,N_2941);
nand UO_204 (O_204,N_2912,N_2967);
or UO_205 (O_205,N_2991,N_2970);
nand UO_206 (O_206,N_2910,N_2909);
and UO_207 (O_207,N_2929,N_2951);
nor UO_208 (O_208,N_2926,N_2923);
or UO_209 (O_209,N_2942,N_2930);
nor UO_210 (O_210,N_2979,N_2956);
nor UO_211 (O_211,N_2982,N_2968);
nor UO_212 (O_212,N_2975,N_2927);
or UO_213 (O_213,N_2911,N_2927);
nor UO_214 (O_214,N_2972,N_2932);
nand UO_215 (O_215,N_2989,N_2930);
nand UO_216 (O_216,N_2926,N_2996);
nand UO_217 (O_217,N_2941,N_2928);
and UO_218 (O_218,N_2937,N_2941);
xor UO_219 (O_219,N_2999,N_2907);
xor UO_220 (O_220,N_2946,N_2905);
xor UO_221 (O_221,N_2906,N_2928);
and UO_222 (O_222,N_2984,N_2993);
nor UO_223 (O_223,N_2920,N_2986);
nand UO_224 (O_224,N_2958,N_2902);
or UO_225 (O_225,N_2923,N_2963);
or UO_226 (O_226,N_2973,N_2953);
nor UO_227 (O_227,N_2968,N_2949);
or UO_228 (O_228,N_2931,N_2955);
nand UO_229 (O_229,N_2970,N_2960);
or UO_230 (O_230,N_2989,N_2912);
nand UO_231 (O_231,N_2921,N_2951);
or UO_232 (O_232,N_2948,N_2916);
nor UO_233 (O_233,N_2912,N_2916);
or UO_234 (O_234,N_2934,N_2925);
nand UO_235 (O_235,N_2971,N_2993);
and UO_236 (O_236,N_2990,N_2939);
nand UO_237 (O_237,N_2969,N_2954);
or UO_238 (O_238,N_2955,N_2968);
nor UO_239 (O_239,N_2937,N_2945);
nand UO_240 (O_240,N_2928,N_2955);
xor UO_241 (O_241,N_2934,N_2974);
or UO_242 (O_242,N_2921,N_2913);
nor UO_243 (O_243,N_2968,N_2915);
or UO_244 (O_244,N_2951,N_2982);
nor UO_245 (O_245,N_2946,N_2919);
xor UO_246 (O_246,N_2908,N_2988);
or UO_247 (O_247,N_2992,N_2906);
or UO_248 (O_248,N_2968,N_2996);
and UO_249 (O_249,N_2937,N_2934);
xnor UO_250 (O_250,N_2989,N_2905);
nor UO_251 (O_251,N_2979,N_2912);
and UO_252 (O_252,N_2933,N_2974);
nor UO_253 (O_253,N_2990,N_2953);
and UO_254 (O_254,N_2974,N_2967);
nor UO_255 (O_255,N_2990,N_2981);
nor UO_256 (O_256,N_2934,N_2953);
nor UO_257 (O_257,N_2987,N_2963);
or UO_258 (O_258,N_2942,N_2955);
nand UO_259 (O_259,N_2996,N_2973);
nor UO_260 (O_260,N_2960,N_2917);
nor UO_261 (O_261,N_2901,N_2905);
nand UO_262 (O_262,N_2999,N_2911);
nand UO_263 (O_263,N_2918,N_2960);
nor UO_264 (O_264,N_2938,N_2918);
nor UO_265 (O_265,N_2940,N_2948);
nor UO_266 (O_266,N_2929,N_2990);
and UO_267 (O_267,N_2968,N_2998);
and UO_268 (O_268,N_2947,N_2933);
and UO_269 (O_269,N_2921,N_2934);
xnor UO_270 (O_270,N_2951,N_2933);
and UO_271 (O_271,N_2938,N_2920);
or UO_272 (O_272,N_2902,N_2981);
nor UO_273 (O_273,N_2982,N_2944);
nand UO_274 (O_274,N_2961,N_2914);
nor UO_275 (O_275,N_2993,N_2975);
or UO_276 (O_276,N_2948,N_2944);
and UO_277 (O_277,N_2955,N_2958);
and UO_278 (O_278,N_2922,N_2916);
nand UO_279 (O_279,N_2999,N_2990);
or UO_280 (O_280,N_2919,N_2934);
or UO_281 (O_281,N_2962,N_2928);
or UO_282 (O_282,N_2917,N_2999);
or UO_283 (O_283,N_2975,N_2976);
nor UO_284 (O_284,N_2962,N_2964);
or UO_285 (O_285,N_2934,N_2955);
xor UO_286 (O_286,N_2921,N_2969);
or UO_287 (O_287,N_2906,N_2932);
and UO_288 (O_288,N_2927,N_2917);
or UO_289 (O_289,N_2969,N_2980);
nor UO_290 (O_290,N_2905,N_2935);
or UO_291 (O_291,N_2925,N_2980);
and UO_292 (O_292,N_2948,N_2921);
or UO_293 (O_293,N_2921,N_2950);
and UO_294 (O_294,N_2929,N_2939);
nand UO_295 (O_295,N_2983,N_2933);
nor UO_296 (O_296,N_2923,N_2932);
nand UO_297 (O_297,N_2926,N_2997);
xnor UO_298 (O_298,N_2961,N_2983);
xor UO_299 (O_299,N_2905,N_2963);
nor UO_300 (O_300,N_2950,N_2978);
or UO_301 (O_301,N_2926,N_2983);
or UO_302 (O_302,N_2982,N_2958);
and UO_303 (O_303,N_2982,N_2916);
and UO_304 (O_304,N_2982,N_2940);
nand UO_305 (O_305,N_2995,N_2981);
or UO_306 (O_306,N_2907,N_2962);
or UO_307 (O_307,N_2984,N_2982);
nand UO_308 (O_308,N_2968,N_2933);
xor UO_309 (O_309,N_2950,N_2928);
nor UO_310 (O_310,N_2946,N_2936);
nor UO_311 (O_311,N_2918,N_2966);
xor UO_312 (O_312,N_2955,N_2990);
nor UO_313 (O_313,N_2900,N_2901);
and UO_314 (O_314,N_2996,N_2952);
nand UO_315 (O_315,N_2936,N_2952);
nor UO_316 (O_316,N_2921,N_2966);
or UO_317 (O_317,N_2914,N_2945);
xnor UO_318 (O_318,N_2935,N_2982);
or UO_319 (O_319,N_2909,N_2981);
nor UO_320 (O_320,N_2999,N_2933);
or UO_321 (O_321,N_2946,N_2951);
or UO_322 (O_322,N_2901,N_2904);
and UO_323 (O_323,N_2918,N_2974);
nor UO_324 (O_324,N_2985,N_2961);
or UO_325 (O_325,N_2922,N_2971);
nand UO_326 (O_326,N_2906,N_2909);
nand UO_327 (O_327,N_2980,N_2947);
and UO_328 (O_328,N_2909,N_2948);
xnor UO_329 (O_329,N_2984,N_2904);
nor UO_330 (O_330,N_2982,N_2985);
nand UO_331 (O_331,N_2963,N_2903);
and UO_332 (O_332,N_2908,N_2976);
nand UO_333 (O_333,N_2941,N_2958);
nor UO_334 (O_334,N_2966,N_2914);
nor UO_335 (O_335,N_2947,N_2940);
or UO_336 (O_336,N_2961,N_2960);
nor UO_337 (O_337,N_2956,N_2948);
and UO_338 (O_338,N_2950,N_2933);
nor UO_339 (O_339,N_2986,N_2981);
nand UO_340 (O_340,N_2925,N_2912);
nor UO_341 (O_341,N_2978,N_2985);
xor UO_342 (O_342,N_2952,N_2938);
nor UO_343 (O_343,N_2994,N_2930);
or UO_344 (O_344,N_2959,N_2954);
or UO_345 (O_345,N_2997,N_2992);
or UO_346 (O_346,N_2938,N_2980);
and UO_347 (O_347,N_2971,N_2956);
or UO_348 (O_348,N_2963,N_2959);
nand UO_349 (O_349,N_2937,N_2950);
or UO_350 (O_350,N_2923,N_2906);
and UO_351 (O_351,N_2941,N_2987);
and UO_352 (O_352,N_2966,N_2992);
nor UO_353 (O_353,N_2921,N_2976);
nand UO_354 (O_354,N_2942,N_2900);
nor UO_355 (O_355,N_2959,N_2989);
and UO_356 (O_356,N_2978,N_2989);
nor UO_357 (O_357,N_2999,N_2919);
nand UO_358 (O_358,N_2990,N_2952);
xor UO_359 (O_359,N_2988,N_2991);
nor UO_360 (O_360,N_2974,N_2955);
nand UO_361 (O_361,N_2997,N_2953);
nor UO_362 (O_362,N_2957,N_2943);
and UO_363 (O_363,N_2933,N_2942);
nor UO_364 (O_364,N_2929,N_2973);
or UO_365 (O_365,N_2996,N_2921);
or UO_366 (O_366,N_2958,N_2945);
and UO_367 (O_367,N_2979,N_2923);
or UO_368 (O_368,N_2905,N_2924);
and UO_369 (O_369,N_2921,N_2907);
or UO_370 (O_370,N_2986,N_2998);
or UO_371 (O_371,N_2967,N_2914);
nor UO_372 (O_372,N_2947,N_2922);
nand UO_373 (O_373,N_2906,N_2968);
nor UO_374 (O_374,N_2968,N_2987);
or UO_375 (O_375,N_2975,N_2950);
and UO_376 (O_376,N_2964,N_2911);
nand UO_377 (O_377,N_2956,N_2913);
nand UO_378 (O_378,N_2940,N_2943);
or UO_379 (O_379,N_2926,N_2975);
nor UO_380 (O_380,N_2900,N_2919);
xnor UO_381 (O_381,N_2928,N_2952);
and UO_382 (O_382,N_2925,N_2902);
or UO_383 (O_383,N_2979,N_2919);
and UO_384 (O_384,N_2972,N_2955);
nand UO_385 (O_385,N_2945,N_2993);
nor UO_386 (O_386,N_2907,N_2910);
and UO_387 (O_387,N_2913,N_2911);
nand UO_388 (O_388,N_2954,N_2990);
nor UO_389 (O_389,N_2938,N_2949);
or UO_390 (O_390,N_2971,N_2973);
and UO_391 (O_391,N_2918,N_2913);
and UO_392 (O_392,N_2953,N_2916);
nor UO_393 (O_393,N_2940,N_2908);
and UO_394 (O_394,N_2900,N_2998);
nand UO_395 (O_395,N_2995,N_2950);
nor UO_396 (O_396,N_2901,N_2941);
or UO_397 (O_397,N_2979,N_2964);
nor UO_398 (O_398,N_2985,N_2970);
or UO_399 (O_399,N_2930,N_2937);
or UO_400 (O_400,N_2956,N_2976);
nand UO_401 (O_401,N_2953,N_2958);
or UO_402 (O_402,N_2990,N_2994);
nor UO_403 (O_403,N_2954,N_2940);
xor UO_404 (O_404,N_2989,N_2940);
xnor UO_405 (O_405,N_2930,N_2922);
nor UO_406 (O_406,N_2940,N_2996);
nand UO_407 (O_407,N_2971,N_2937);
xor UO_408 (O_408,N_2940,N_2905);
and UO_409 (O_409,N_2978,N_2928);
nand UO_410 (O_410,N_2942,N_2998);
and UO_411 (O_411,N_2963,N_2964);
nand UO_412 (O_412,N_2983,N_2981);
nand UO_413 (O_413,N_2984,N_2985);
nand UO_414 (O_414,N_2903,N_2953);
xnor UO_415 (O_415,N_2944,N_2950);
nor UO_416 (O_416,N_2933,N_2970);
and UO_417 (O_417,N_2963,N_2951);
nand UO_418 (O_418,N_2928,N_2945);
nor UO_419 (O_419,N_2948,N_2900);
or UO_420 (O_420,N_2935,N_2913);
nor UO_421 (O_421,N_2973,N_2978);
and UO_422 (O_422,N_2943,N_2971);
or UO_423 (O_423,N_2929,N_2974);
nor UO_424 (O_424,N_2928,N_2907);
or UO_425 (O_425,N_2970,N_2917);
or UO_426 (O_426,N_2986,N_2909);
nand UO_427 (O_427,N_2970,N_2942);
or UO_428 (O_428,N_2928,N_2966);
nor UO_429 (O_429,N_2936,N_2983);
nand UO_430 (O_430,N_2945,N_2915);
xor UO_431 (O_431,N_2996,N_2929);
xnor UO_432 (O_432,N_2906,N_2965);
and UO_433 (O_433,N_2936,N_2945);
nand UO_434 (O_434,N_2932,N_2901);
or UO_435 (O_435,N_2978,N_2921);
or UO_436 (O_436,N_2957,N_2902);
nand UO_437 (O_437,N_2921,N_2970);
or UO_438 (O_438,N_2931,N_2987);
or UO_439 (O_439,N_2943,N_2931);
nand UO_440 (O_440,N_2997,N_2907);
or UO_441 (O_441,N_2994,N_2902);
nand UO_442 (O_442,N_2911,N_2933);
and UO_443 (O_443,N_2961,N_2935);
nand UO_444 (O_444,N_2987,N_2914);
nand UO_445 (O_445,N_2951,N_2981);
nand UO_446 (O_446,N_2929,N_2919);
or UO_447 (O_447,N_2915,N_2965);
or UO_448 (O_448,N_2999,N_2938);
nand UO_449 (O_449,N_2947,N_2956);
and UO_450 (O_450,N_2975,N_2907);
nand UO_451 (O_451,N_2933,N_2925);
and UO_452 (O_452,N_2947,N_2917);
and UO_453 (O_453,N_2933,N_2900);
and UO_454 (O_454,N_2926,N_2999);
nor UO_455 (O_455,N_2934,N_2988);
nand UO_456 (O_456,N_2990,N_2998);
and UO_457 (O_457,N_2995,N_2923);
and UO_458 (O_458,N_2936,N_2972);
and UO_459 (O_459,N_2968,N_2985);
xor UO_460 (O_460,N_2953,N_2902);
or UO_461 (O_461,N_2974,N_2985);
or UO_462 (O_462,N_2982,N_2981);
and UO_463 (O_463,N_2972,N_2942);
and UO_464 (O_464,N_2978,N_2962);
or UO_465 (O_465,N_2953,N_2956);
nand UO_466 (O_466,N_2953,N_2940);
nor UO_467 (O_467,N_2910,N_2971);
and UO_468 (O_468,N_2915,N_2990);
nor UO_469 (O_469,N_2926,N_2916);
nor UO_470 (O_470,N_2973,N_2964);
nand UO_471 (O_471,N_2935,N_2922);
or UO_472 (O_472,N_2969,N_2976);
nand UO_473 (O_473,N_2990,N_2918);
nor UO_474 (O_474,N_2931,N_2935);
and UO_475 (O_475,N_2999,N_2969);
nor UO_476 (O_476,N_2967,N_2982);
xor UO_477 (O_477,N_2933,N_2997);
and UO_478 (O_478,N_2958,N_2993);
nand UO_479 (O_479,N_2975,N_2965);
nor UO_480 (O_480,N_2946,N_2974);
and UO_481 (O_481,N_2986,N_2927);
xor UO_482 (O_482,N_2984,N_2962);
nand UO_483 (O_483,N_2906,N_2952);
nand UO_484 (O_484,N_2914,N_2920);
and UO_485 (O_485,N_2988,N_2913);
and UO_486 (O_486,N_2982,N_2986);
or UO_487 (O_487,N_2958,N_2969);
nor UO_488 (O_488,N_2909,N_2954);
and UO_489 (O_489,N_2925,N_2901);
nor UO_490 (O_490,N_2956,N_2909);
and UO_491 (O_491,N_2969,N_2908);
nand UO_492 (O_492,N_2949,N_2990);
nand UO_493 (O_493,N_2912,N_2954);
nor UO_494 (O_494,N_2926,N_2942);
nand UO_495 (O_495,N_2912,N_2964);
nor UO_496 (O_496,N_2995,N_2987);
and UO_497 (O_497,N_2907,N_2923);
and UO_498 (O_498,N_2904,N_2972);
xor UO_499 (O_499,N_2944,N_2952);
endmodule