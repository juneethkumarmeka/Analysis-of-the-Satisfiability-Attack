module basic_1500_15000_2000_3_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10035,N_10037,N_10038,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10059,N_10060,N_10061,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10083,N_10084,N_10085,N_10086,N_10088,N_10089,N_10090,N_10093,N_10094,N_10095,N_10096,N_10098,N_10099,N_10100,N_10102,N_10103,N_10104,N_10106,N_10107,N_10108,N_10109,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10121,N_10122,N_10123,N_10124,N_10125,N_10128,N_10130,N_10132,N_10133,N_10135,N_10137,N_10138,N_10139,N_10140,N_10142,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10170,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10193,N_10194,N_10196,N_10197,N_10198,N_10200,N_10201,N_10203,N_10204,N_10205,N_10207,N_10208,N_10210,N_10211,N_10212,N_10214,N_10215,N_10216,N_10218,N_10219,N_10221,N_10222,N_10223,N_10225,N_10227,N_10228,N_10229,N_10231,N_10232,N_10233,N_10236,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10249,N_10250,N_10251,N_10252,N_10253,N_10255,N_10256,N_10257,N_10259,N_10260,N_10261,N_10262,N_10264,N_10265,N_10266,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10297,N_10298,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10309,N_10311,N_10312,N_10313,N_10315,N_10317,N_10318,N_10320,N_10321,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10332,N_10333,N_10334,N_10337,N_10339,N_10340,N_10341,N_10345,N_10347,N_10349,N_10351,N_10352,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10361,N_10362,N_10363,N_10365,N_10366,N_10367,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10379,N_10380,N_10382,N_10383,N_10384,N_10386,N_10387,N_10389,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10400,N_10403,N_10404,N_10405,N_10407,N_10409,N_10410,N_10411,N_10412,N_10415,N_10416,N_10418,N_10419,N_10421,N_10422,N_10423,N_10424,N_10428,N_10429,N_10430,N_10432,N_10434,N_10436,N_10437,N_10438,N_10439,N_10442,N_10443,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10453,N_10454,N_10455,N_10456,N_10458,N_10459,N_10460,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10471,N_10473,N_10474,N_10478,N_10479,N_10480,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10539,N_10540,N_10541,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10554,N_10555,N_10556,N_10558,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10595,N_10596,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10616,N_10617,N_10618,N_10619,N_10620,N_10622,N_10623,N_10624,N_10626,N_10627,N_10628,N_10629,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10640,N_10642,N_10644,N_10645,N_10646,N_10647,N_10649,N_10650,N_10651,N_10652,N_10654,N_10656,N_10657,N_10659,N_10660,N_10661,N_10664,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10684,N_10685,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10721,N_10722,N_10723,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10734,N_10735,N_10736,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10754,N_10755,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10795,N_10796,N_10797,N_10799,N_10801,N_10802,N_10803,N_10805,N_10806,N_10807,N_10808,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10872,N_10873,N_10874,N_10876,N_10877,N_10878,N_10880,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10890,N_10891,N_10892,N_10893,N_10895,N_10896,N_10899,N_10900,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10916,N_10917,N_10919,N_10920,N_10921,N_10922,N_10924,N_10925,N_10926,N_10927,N_10928,N_10931,N_10933,N_10937,N_10938,N_10939,N_10941,N_10943,N_10944,N_10945,N_10946,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10964,N_10967,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10977,N_10979,N_10980,N_10981,N_10982,N_10985,N_10986,N_10988,N_10989,N_10990,N_10991,N_10992,N_10994,N_10996,N_10997,N_10999,N_11002,N_11003,N_11005,N_11008,N_11009,N_11010,N_11011,N_11014,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11023,N_11024,N_11026,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11035,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11047,N_11048,N_11049,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11079,N_11081,N_11082,N_11083,N_11084,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11093,N_11094,N_11095,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11119,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11139,N_11140,N_11141,N_11143,N_11145,N_11146,N_11147,N_11149,N_11150,N_11152,N_11153,N_11154,N_11155,N_11157,N_11158,N_11161,N_11162,N_11163,N_11164,N_11165,N_11167,N_11168,N_11169,N_11171,N_11172,N_11173,N_11175,N_11177,N_11178,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11192,N_11193,N_11194,N_11196,N_11197,N_11199,N_11200,N_11202,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11213,N_11214,N_11216,N_11217,N_11218,N_11219,N_11221,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11230,N_11231,N_11232,N_11233,N_11234,N_11236,N_11237,N_11238,N_11239,N_11241,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11252,N_11253,N_11254,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11265,N_11266,N_11268,N_11269,N_11271,N_11272,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11282,N_11283,N_11285,N_11286,N_11287,N_11291,N_11293,N_11294,N_11297,N_11299,N_11300,N_11301,N_11302,N_11303,N_11306,N_11307,N_11308,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11349,N_11350,N_11352,N_11354,N_11355,N_11356,N_11358,N_11359,N_11360,N_11361,N_11362,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11375,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11387,N_11388,N_11390,N_11391,N_11392,N_11394,N_11395,N_11396,N_11397,N_11398,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11410,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11440,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11454,N_11455,N_11456,N_11458,N_11459,N_11460,N_11461,N_11463,N_11464,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11482,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11508,N_11510,N_11511,N_11512,N_11513,N_11514,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11526,N_11528,N_11529,N_11532,N_11533,N_11536,N_11537,N_11538,N_11539,N_11540,N_11542,N_11543,N_11544,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11555,N_11556,N_11558,N_11559,N_11560,N_11561,N_11562,N_11564,N_11565,N_11566,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11579,N_11580,N_11582,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11612,N_11613,N_11614,N_11617,N_11618,N_11619,N_11620,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11629,N_11630,N_11631,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11650,N_11651,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11693,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11717,N_11718,N_11720,N_11721,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11731,N_11732,N_11733,N_11734,N_11735,N_11737,N_11738,N_11739,N_11740,N_11742,N_11744,N_11745,N_11746,N_11747,N_11748,N_11750,N_11752,N_11753,N_11754,N_11755,N_11756,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11773,N_11774,N_11775,N_11776,N_11778,N_11779,N_11780,N_11781,N_11782,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11793,N_11794,N_11795,N_11796,N_11798,N_11799,N_11800,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11814,N_11815,N_11816,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11826,N_11827,N_11828,N_11829,N_11831,N_11832,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11847,N_11848,N_11849,N_11851,N_11852,N_11854,N_11855,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11865,N_11866,N_11867,N_11868,N_11869,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11881,N_11882,N_11883,N_11885,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11897,N_11899,N_11900,N_11901,N_11902,N_11905,N_11906,N_11908,N_11909,N_11910,N_11912,N_11914,N_11915,N_11916,N_11917,N_11918,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11936,N_11937,N_11938,N_11939,N_11940,N_11942,N_11943,N_11944,N_11945,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11955,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11967,N_11968,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11986,N_11988,N_11989,N_11990,N_11991,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12071,N_12072,N_12073,N_12074,N_12075,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12089,N_12090,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12106,N_12107,N_12108,N_12109,N_12112,N_12113,N_12114,N_12117,N_12118,N_12120,N_12121,N_12124,N_12126,N_12128,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12146,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12161,N_12163,N_12165,N_12167,N_12168,N_12169,N_12171,N_12172,N_12175,N_12178,N_12179,N_12181,N_12182,N_12183,N_12184,N_12186,N_12187,N_12189,N_12190,N_12192,N_12194,N_12195,N_12197,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12217,N_12218,N_12219,N_12220,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12241,N_12242,N_12244,N_12246,N_12247,N_12250,N_12252,N_12253,N_12254,N_12255,N_12257,N_12258,N_12261,N_12262,N_12264,N_12265,N_12267,N_12268,N_12269,N_12270,N_12272,N_12273,N_12274,N_12277,N_12278,N_12279,N_12280,N_12281,N_12283,N_12284,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12316,N_12317,N_12318,N_12319,N_12321,N_12322,N_12324,N_12325,N_12326,N_12327,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12353,N_12354,N_12357,N_12358,N_12359,N_12360,N_12362,N_12363,N_12365,N_12366,N_12367,N_12368,N_12369,N_12371,N_12372,N_12373,N_12374,N_12375,N_12377,N_12378,N_12379,N_12381,N_12382,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12391,N_12392,N_12393,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12404,N_12405,N_12409,N_12410,N_12411,N_12412,N_12413,N_12416,N_12418,N_12419,N_12420,N_12421,N_12422,N_12424,N_12426,N_12427,N_12428,N_12430,N_12431,N_12434,N_12436,N_12437,N_12439,N_12440,N_12441,N_12442,N_12444,N_12445,N_12446,N_12448,N_12450,N_12451,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12462,N_12463,N_12465,N_12468,N_12469,N_12470,N_12471,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12501,N_12502,N_12503,N_12504,N_12506,N_12507,N_12508,N_12510,N_12511,N_12512,N_12513,N_12514,N_12516,N_12517,N_12519,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12531,N_12532,N_12533,N_12534,N_12535,N_12538,N_12539,N_12541,N_12542,N_12543,N_12545,N_12546,N_12547,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12564,N_12566,N_12567,N_12568,N_12569,N_12571,N_12572,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12584,N_12585,N_12587,N_12588,N_12589,N_12590,N_12591,N_12593,N_12594,N_12596,N_12597,N_12599,N_12600,N_12602,N_12603,N_12604,N_12605,N_12606,N_12608,N_12609,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12624,N_12626,N_12627,N_12628,N_12629,N_12631,N_12632,N_12633,N_12634,N_12636,N_12638,N_12639,N_12640,N_12641,N_12643,N_12644,N_12645,N_12646,N_12647,N_12649,N_12650,N_12651,N_12653,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12679,N_12680,N_12681,N_12682,N_12685,N_12686,N_12687,N_12689,N_12690,N_12691,N_12692,N_12693,N_12696,N_12697,N_12698,N_12699,N_12701,N_12702,N_12703,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12735,N_12737,N_12738,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12748,N_12750,N_12751,N_12752,N_12753,N_12754,N_12756,N_12757,N_12758,N_12761,N_12764,N_12765,N_12766,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12779,N_12780,N_12781,N_12782,N_12784,N_12786,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12798,N_12800,N_12802,N_12803,N_12804,N_12805,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12826,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12849,N_12850,N_12851,N_12853,N_12854,N_12855,N_12858,N_12859,N_12860,N_12863,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12892,N_12893,N_12894,N_12895,N_12896,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12932,N_12933,N_12934,N_12937,N_12940,N_12941,N_12942,N_12944,N_12945,N_12946,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12981,N_12983,N_12985,N_12986,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13029,N_13030,N_13031,N_13033,N_13034,N_13035,N_13037,N_13038,N_13039,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13059,N_13060,N_13061,N_13062,N_13063,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13088,N_13090,N_13091,N_13093,N_13094,N_13097,N_13098,N_13102,N_13104,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13133,N_13135,N_13136,N_13137,N_13138,N_13140,N_13141,N_13142,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13153,N_13154,N_13156,N_13158,N_13159,N_13160,N_13161,N_13164,N_13165,N_13166,N_13167,N_13169,N_13170,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13198,N_13199,N_13202,N_13203,N_13204,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13213,N_13214,N_13215,N_13216,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13227,N_13228,N_13230,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13243,N_13244,N_13245,N_13246,N_13248,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13260,N_13261,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13279,N_13280,N_13281,N_13282,N_13284,N_13285,N_13286,N_13287,N_13288,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13357,N_13358,N_13359,N_13360,N_13362,N_13363,N_13364,N_13365,N_13366,N_13368,N_13369,N_13372,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13381,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13393,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13404,N_13405,N_13406,N_13407,N_13410,N_13411,N_13412,N_13414,N_13415,N_13416,N_13417,N_13418,N_13420,N_13421,N_13423,N_13424,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13439,N_13441,N_13442,N_13443,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13454,N_13455,N_13456,N_13457,N_13459,N_13460,N_13462,N_13463,N_13464,N_13465,N_13466,N_13468,N_13469,N_13470,N_13471,N_13472,N_13474,N_13475,N_13476,N_13477,N_13478,N_13481,N_13482,N_13485,N_13486,N_13487,N_13488,N_13490,N_13491,N_13492,N_13495,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13525,N_13526,N_13528,N_13529,N_13530,N_13531,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13542,N_13543,N_13544,N_13545,N_13546,N_13548,N_13549,N_13550,N_13551,N_13552,N_13554,N_13556,N_13557,N_13558,N_13559,N_13560,N_13563,N_13564,N_13565,N_13566,N_13567,N_13569,N_13570,N_13571,N_13572,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13584,N_13587,N_13588,N_13589,N_13592,N_13594,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13612,N_13613,N_13614,N_13618,N_13619,N_13620,N_13621,N_13622,N_13624,N_13625,N_13626,N_13627,N_13629,N_13630,N_13632,N_13633,N_13634,N_13636,N_13637,N_13640,N_13641,N_13643,N_13644,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13663,N_13664,N_13665,N_13666,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13687,N_13688,N_13689,N_13690,N_13691,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13707,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13726,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13795,N_13796,N_13797,N_13799,N_13800,N_13801,N_13802,N_13803,N_13805,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13814,N_13815,N_13816,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13837,N_13838,N_13840,N_13841,N_13842,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13857,N_13858,N_13859,N_13861,N_13862,N_13864,N_13865,N_13867,N_13868,N_13869,N_13870,N_13872,N_13873,N_13876,N_13877,N_13878,N_13880,N_13881,N_13883,N_13884,N_13885,N_13886,N_13887,N_13889,N_13890,N_13892,N_13893,N_13894,N_13895,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13925,N_13927,N_13928,N_13930,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13955,N_13956,N_13958,N_13960,N_13961,N_13962,N_13963,N_13965,N_13967,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13999,N_14000,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14009,N_14010,N_14012,N_14014,N_14017,N_14018,N_14019,N_14020,N_14021,N_14023,N_14024,N_14025,N_14026,N_14028,N_14030,N_14031,N_14032,N_14034,N_14035,N_14036,N_14038,N_14039,N_14040,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14068,N_14069,N_14070,N_14071,N_14074,N_14075,N_14076,N_14078,N_14079,N_14080,N_14081,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14094,N_14095,N_14096,N_14097,N_14099,N_14100,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14134,N_14135,N_14136,N_14137,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14148,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14158,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14180,N_14181,N_14183,N_14185,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14204,N_14206,N_14208,N_14210,N_14211,N_14212,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14231,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14248,N_14251,N_14253,N_14254,N_14256,N_14257,N_14258,N_14259,N_14261,N_14262,N_14263,N_14264,N_14265,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14276,N_14277,N_14278,N_14279,N_14281,N_14283,N_14284,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14304,N_14305,N_14307,N_14308,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14321,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14370,N_14372,N_14375,N_14376,N_14378,N_14379,N_14380,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14389,N_14390,N_14392,N_14393,N_14394,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14405,N_14406,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14444,N_14446,N_14448,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14473,N_14474,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14484,N_14485,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14494,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14504,N_14505,N_14508,N_14509,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14524,N_14525,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14537,N_14538,N_14539,N_14540,N_14541,N_14543,N_14544,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14555,N_14556,N_14557,N_14559,N_14560,N_14561,N_14563,N_14564,N_14567,N_14568,N_14569,N_14570,N_14572,N_14573,N_14574,N_14575,N_14576,N_14578,N_14580,N_14582,N_14583,N_14584,N_14586,N_14587,N_14588,N_14589,N_14590,N_14592,N_14593,N_14594,N_14595,N_14597,N_14599,N_14601,N_14602,N_14603,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14614,N_14615,N_14616,N_14618,N_14619,N_14622,N_14623,N_14624,N_14625,N_14626,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14653,N_14654,N_14655,N_14656,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14665,N_14666,N_14667,N_14668,N_14669,N_14671,N_14672,N_14673,N_14674,N_14675,N_14677,N_14678,N_14680,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14696,N_14697,N_14698,N_14700,N_14702,N_14703,N_14704,N_14707,N_14709,N_14710,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14726,N_14727,N_14728,N_14729,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14742,N_14743,N_14746,N_14747,N_14748,N_14749,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14761,N_14762,N_14763,N_14765,N_14766,N_14767,N_14768,N_14770,N_14771,N_14772,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14787,N_14789,N_14790,N_14791,N_14792,N_14793,N_14795,N_14796,N_14797,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14810,N_14812,N_14813,N_14814,N_14816,N_14817,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14842,N_14843,N_14844,N_14846,N_14847,N_14848,N_14849,N_14850,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14873,N_14875,N_14877,N_14878,N_14880,N_14881,N_14883,N_14884,N_14885,N_14887,N_14888,N_14889,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14898,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14911,N_14912,N_14914,N_14915,N_14916,N_14917,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14937,N_14938,N_14939,N_14940,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14949,N_14950,N_14951,N_14953,N_14954,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14973,N_14974,N_14975,N_14977,N_14978,N_14979,N_14981,N_14982,N_14984,N_14985,N_14986,N_14988,N_14989,N_14990,N_14991,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_760,In_1442);
nand U1 (N_1,In_472,In_1000);
and U2 (N_2,In_247,In_58);
nor U3 (N_3,In_1203,In_1039);
nor U4 (N_4,In_517,In_959);
or U5 (N_5,In_821,In_866);
and U6 (N_6,In_295,In_1051);
or U7 (N_7,In_925,In_28);
nor U8 (N_8,In_1372,In_829);
nand U9 (N_9,In_1440,In_50);
xnor U10 (N_10,In_1156,In_623);
and U11 (N_11,In_108,In_805);
or U12 (N_12,In_1232,In_1395);
nor U13 (N_13,In_605,In_778);
nand U14 (N_14,In_158,In_411);
xor U15 (N_15,In_225,In_318);
nor U16 (N_16,In_569,In_1017);
and U17 (N_17,In_556,In_150);
or U18 (N_18,In_455,In_574);
nand U19 (N_19,In_991,In_835);
or U20 (N_20,In_586,In_1170);
nor U21 (N_21,In_642,In_75);
and U22 (N_22,In_1475,In_815);
nand U23 (N_23,In_794,In_292);
nand U24 (N_24,In_427,In_1464);
nand U25 (N_25,In_369,In_1484);
nor U26 (N_26,In_701,In_1313);
nand U27 (N_27,In_1300,In_1323);
xor U28 (N_28,In_1083,In_1116);
nor U29 (N_29,In_1067,In_1383);
and U30 (N_30,In_618,In_1216);
xnor U31 (N_31,In_1454,In_254);
or U32 (N_32,In_1198,In_1251);
or U33 (N_33,In_1254,In_1416);
and U34 (N_34,In_1191,In_421);
nor U35 (N_35,In_1321,In_613);
xor U36 (N_36,In_130,In_33);
or U37 (N_37,In_974,In_219);
or U38 (N_38,In_432,In_806);
and U39 (N_39,In_984,In_234);
and U40 (N_40,In_624,In_1160);
and U41 (N_41,In_46,In_113);
nand U42 (N_42,In_339,In_1371);
nand U43 (N_43,In_387,In_197);
nor U44 (N_44,In_453,In_338);
nand U45 (N_45,In_350,In_533);
nand U46 (N_46,In_347,In_697);
xnor U47 (N_47,In_633,In_561);
xor U48 (N_48,In_983,In_595);
or U49 (N_49,In_737,In_291);
xor U50 (N_50,In_985,In_930);
nor U51 (N_51,In_1212,In_804);
nand U52 (N_52,In_843,In_980);
nand U53 (N_53,In_1339,In_77);
or U54 (N_54,In_1062,In_1226);
nand U55 (N_55,In_988,In_931);
and U56 (N_56,In_851,In_861);
or U57 (N_57,In_1334,In_721);
or U58 (N_58,In_445,In_43);
nand U59 (N_59,In_252,In_598);
nor U60 (N_60,In_854,In_152);
and U61 (N_61,In_61,In_422);
nor U62 (N_62,In_1043,In_630);
nand U63 (N_63,In_887,In_1024);
or U64 (N_64,In_265,In_731);
nor U65 (N_65,In_536,In_606);
nand U66 (N_66,In_943,In_430);
and U67 (N_67,In_520,In_1081);
nand U68 (N_68,In_1135,In_932);
nand U69 (N_69,In_1301,In_629);
nand U70 (N_70,In_1033,In_85);
nor U71 (N_71,In_1046,In_719);
nor U72 (N_72,In_581,In_329);
or U73 (N_73,In_63,In_636);
and U74 (N_74,In_51,In_740);
nor U75 (N_75,In_24,In_681);
nand U76 (N_76,In_138,In_191);
nor U77 (N_77,In_897,In_1209);
or U78 (N_78,In_249,In_590);
or U79 (N_79,In_129,In_69);
or U80 (N_80,In_15,In_1399);
nand U81 (N_81,In_429,In_706);
and U82 (N_82,In_1435,In_353);
or U83 (N_83,In_196,In_567);
and U84 (N_84,In_954,In_522);
or U85 (N_85,In_74,In_1456);
nand U86 (N_86,In_944,In_71);
and U87 (N_87,In_883,In_1140);
nand U88 (N_88,In_888,In_1279);
nor U89 (N_89,In_386,In_157);
nor U90 (N_90,In_830,In_882);
nand U91 (N_91,In_1034,In_1378);
or U92 (N_92,In_463,In_857);
xor U93 (N_93,In_1109,In_92);
nand U94 (N_94,In_653,In_1218);
nor U95 (N_95,In_299,In_34);
nand U96 (N_96,In_1031,In_457);
nand U97 (N_97,In_631,In_1197);
or U98 (N_98,In_608,In_456);
nor U99 (N_99,In_136,In_782);
or U100 (N_100,In_1326,In_987);
nor U101 (N_101,In_20,In_83);
nand U102 (N_102,In_818,In_1483);
nand U103 (N_103,In_976,In_1286);
nor U104 (N_104,In_290,In_497);
and U105 (N_105,In_436,In_668);
nor U106 (N_106,In_165,In_1258);
or U107 (N_107,In_1108,In_967);
nor U108 (N_108,In_226,In_652);
nor U109 (N_109,In_840,In_377);
and U110 (N_110,In_900,In_1177);
and U111 (N_111,In_529,In_648);
or U112 (N_112,In_998,In_142);
xnor U113 (N_113,In_1432,In_1259);
nor U114 (N_114,In_870,In_268);
nand U115 (N_115,In_696,In_279);
nand U116 (N_116,In_612,In_286);
and U117 (N_117,In_560,In_281);
nand U118 (N_118,In_1136,In_1292);
xor U119 (N_119,In_1101,In_1495);
xnor U120 (N_120,In_104,In_1413);
and U121 (N_121,In_963,In_880);
or U122 (N_122,In_1319,In_534);
and U123 (N_123,In_895,In_1009);
or U124 (N_124,In_1458,In_145);
xnor U125 (N_125,In_1362,In_908);
or U126 (N_126,In_1318,In_1419);
or U127 (N_127,In_32,In_975);
nor U128 (N_128,In_190,In_1436);
or U129 (N_129,In_1246,In_773);
nand U130 (N_130,In_233,In_218);
or U131 (N_131,In_575,In_1146);
and U132 (N_132,In_645,In_968);
or U133 (N_133,In_690,In_126);
or U134 (N_134,In_950,In_1010);
or U135 (N_135,In_564,In_181);
or U136 (N_136,In_1430,In_1186);
or U137 (N_137,In_358,In_966);
nor U138 (N_138,In_559,In_1176);
nor U139 (N_139,In_379,In_651);
nor U140 (N_140,In_1348,In_1283);
nand U141 (N_141,In_1032,In_524);
or U142 (N_142,In_334,In_1478);
xor U143 (N_143,In_867,In_693);
or U144 (N_144,In_712,In_727);
nand U145 (N_145,In_797,In_44);
or U146 (N_146,In_312,In_1200);
xor U147 (N_147,In_444,In_756);
nand U148 (N_148,In_206,In_902);
or U149 (N_149,In_788,In_242);
nand U150 (N_150,In_997,In_549);
nand U151 (N_151,In_1063,In_755);
xnor U152 (N_152,In_765,In_1237);
or U153 (N_153,In_604,In_1414);
nand U154 (N_154,In_1201,In_1139);
xor U155 (N_155,In_443,In_1007);
or U156 (N_156,In_1097,In_232);
or U157 (N_157,In_1470,In_1137);
nand U158 (N_158,In_596,In_1477);
and U159 (N_159,In_1482,In_1335);
nor U160 (N_160,In_1157,In_493);
nor U161 (N_161,In_90,In_514);
and U162 (N_162,In_578,In_949);
nor U163 (N_163,In_924,In_376);
nor U164 (N_164,In_1315,In_656);
nor U165 (N_165,In_128,In_1072);
or U166 (N_166,In_1090,In_717);
nand U167 (N_167,In_1208,In_1274);
and U168 (N_168,In_726,In_1498);
and U169 (N_169,In_1102,In_904);
nand U170 (N_170,In_1266,In_327);
nor U171 (N_171,In_490,In_451);
or U172 (N_172,In_1280,In_1131);
xnor U173 (N_173,In_484,In_698);
nand U174 (N_174,In_29,In_619);
and U175 (N_175,In_1056,In_1341);
nor U176 (N_176,In_532,In_381);
or U177 (N_177,In_1049,In_1337);
xor U178 (N_178,In_607,In_1094);
or U179 (N_179,In_1125,In_396);
or U180 (N_180,In_66,In_30);
or U181 (N_181,In_10,In_97);
and U182 (N_182,In_474,In_343);
nor U183 (N_183,In_222,In_1370);
nor U184 (N_184,In_847,In_1330);
nand U185 (N_185,In_1175,In_48);
and U186 (N_186,In_431,In_912);
and U187 (N_187,In_1181,In_235);
or U188 (N_188,In_101,In_1468);
and U189 (N_189,In_1223,In_1026);
or U190 (N_190,In_280,In_1398);
nor U191 (N_191,In_57,In_1328);
or U192 (N_192,In_1401,In_37);
nand U193 (N_193,In_1023,In_768);
nor U194 (N_194,In_600,In_205);
nor U195 (N_195,In_799,In_1016);
and U196 (N_196,In_25,In_770);
or U197 (N_197,In_1141,In_995);
or U198 (N_198,In_12,In_582);
xnor U199 (N_199,In_135,In_735);
or U200 (N_200,In_494,In_237);
xor U201 (N_201,In_552,In_146);
or U202 (N_202,In_40,In_1096);
nand U203 (N_203,In_223,In_510);
or U204 (N_204,In_89,In_1382);
and U205 (N_205,In_841,In_1297);
nand U206 (N_206,In_438,In_972);
nand U207 (N_207,In_872,In_957);
nand U208 (N_208,In_478,In_858);
and U209 (N_209,In_566,In_419);
nor U210 (N_210,In_1014,In_82);
or U211 (N_211,In_184,In_543);
nor U212 (N_212,In_501,In_397);
xor U213 (N_213,In_124,In_580);
nor U214 (N_214,In_1104,In_625);
nor U215 (N_215,In_8,In_163);
and U216 (N_216,In_70,In_793);
nand U217 (N_217,In_786,In_336);
xnor U218 (N_218,In_321,In_337);
or U219 (N_219,In_182,In_1054);
nor U220 (N_220,In_413,In_248);
nand U221 (N_221,In_39,In_241);
or U222 (N_222,In_1368,In_834);
or U223 (N_223,In_1192,In_907);
xnor U224 (N_224,In_647,In_876);
nand U225 (N_225,In_231,In_850);
nand U226 (N_226,In_951,In_294);
or U227 (N_227,In_415,In_258);
nand U228 (N_228,In_674,In_1367);
xnor U229 (N_229,In_1412,In_1271);
or U230 (N_230,In_477,In_649);
nand U231 (N_231,In_531,In_766);
nand U232 (N_232,In_352,In_1444);
nand U233 (N_233,In_355,In_709);
or U234 (N_234,In_481,In_1317);
and U235 (N_235,In_1188,In_156);
or U236 (N_236,In_1243,In_1343);
nor U237 (N_237,In_1075,In_673);
nor U238 (N_238,In_1278,In_84);
or U239 (N_239,In_111,In_1403);
and U240 (N_240,In_707,In_1047);
nand U241 (N_241,In_592,In_1462);
nor U242 (N_242,In_288,In_588);
and U243 (N_243,In_1205,In_1305);
nor U244 (N_244,In_915,In_1437);
nand U245 (N_245,In_434,In_492);
or U246 (N_246,In_365,In_1418);
nor U247 (N_247,In_500,In_399);
nand U248 (N_248,In_1110,In_22);
and U249 (N_249,In_684,In_420);
nand U250 (N_250,In_485,In_662);
nor U251 (N_251,In_1098,In_742);
or U252 (N_252,In_131,In_1302);
nor U253 (N_253,In_122,In_246);
or U254 (N_254,In_824,In_395);
nand U255 (N_255,In_836,In_779);
or U256 (N_256,In_169,In_1037);
or U257 (N_257,In_732,In_934);
or U258 (N_258,In_76,In_59);
nand U259 (N_259,In_371,In_473);
nand U260 (N_260,In_1429,In_792);
nor U261 (N_261,In_1406,In_127);
or U262 (N_262,In_1185,In_744);
and U263 (N_263,In_209,In_425);
or U264 (N_264,In_1095,In_401);
xor U265 (N_265,In_166,In_784);
xor U266 (N_266,In_1423,In_49);
nor U267 (N_267,In_1189,In_1245);
and U268 (N_268,In_1147,In_133);
nor U269 (N_269,In_270,In_1338);
and U270 (N_270,In_1356,In_911);
nor U271 (N_271,In_547,In_894);
and U272 (N_272,In_1142,In_486);
nand U273 (N_273,In_893,In_573);
xor U274 (N_274,In_919,In_518);
nand U275 (N_275,In_297,In_1115);
nor U276 (N_276,In_585,In_1002);
nand U277 (N_277,In_319,In_713);
and U278 (N_278,In_1447,In_1261);
nor U279 (N_279,In_889,In_535);
nand U280 (N_280,In_0,In_1113);
or U281 (N_281,In_1421,In_817);
nor U282 (N_282,In_67,In_1267);
or U283 (N_283,In_1040,In_667);
or U284 (N_284,In_103,In_459);
xor U285 (N_285,In_1127,In_1018);
and U286 (N_286,In_638,In_78);
and U287 (N_287,In_366,In_1207);
nand U288 (N_288,In_1019,In_545);
nor U289 (N_289,In_999,In_316);
and U290 (N_290,In_1249,In_842);
or U291 (N_291,In_407,In_689);
nor U292 (N_292,In_269,In_198);
nand U293 (N_293,In_368,In_610);
or U294 (N_294,In_21,In_1225);
and U295 (N_295,In_512,In_4);
nor U296 (N_296,In_1304,In_476);
nor U297 (N_297,In_16,In_1182);
nor U298 (N_298,In_1151,In_174);
nor U299 (N_299,In_303,In_121);
xor U300 (N_300,In_1045,In_922);
and U301 (N_301,In_1340,In_351);
nand U302 (N_302,In_1027,In_1263);
or U303 (N_303,In_1298,In_828);
nand U304 (N_304,In_583,In_491);
or U305 (N_305,In_240,In_1349);
or U306 (N_306,In_1076,In_1145);
nand U307 (N_307,In_1048,In_349);
nor U308 (N_308,In_496,In_679);
nor U309 (N_309,In_200,In_302);
nand U310 (N_310,In_960,In_1080);
nand U311 (N_311,In_1257,In_1168);
nand U312 (N_312,In_202,In_989);
or U313 (N_313,In_1250,In_1086);
xnor U314 (N_314,In_1346,In_172);
or U315 (N_315,In_1380,In_741);
xor U316 (N_316,In_1481,In_306);
xor U317 (N_317,In_467,In_1171);
xnor U318 (N_318,In_1415,In_1363);
nand U319 (N_319,In_1091,In_137);
xor U320 (N_320,In_26,In_1264);
and U321 (N_321,In_1473,In_1417);
and U322 (N_322,In_1129,In_204);
or U323 (N_323,In_266,In_282);
nand U324 (N_324,In_958,In_255);
or U325 (N_325,In_1265,In_918);
nand U326 (N_326,In_1052,In_859);
nor U327 (N_327,In_1494,In_60);
nor U328 (N_328,In_1480,In_1314);
nor U329 (N_329,In_916,In_753);
or U330 (N_330,In_783,In_827);
or U331 (N_331,In_1235,In_56);
or U332 (N_332,In_364,In_17);
or U333 (N_333,In_1231,In_1431);
nor U334 (N_334,In_1433,In_764);
nor U335 (N_335,In_965,In_1277);
or U336 (N_336,In_1451,In_822);
nand U337 (N_337,In_1117,In_382);
and U338 (N_338,In_1028,In_856);
nor U339 (N_339,In_99,In_826);
nor U340 (N_340,In_941,In_315);
nand U341 (N_341,In_1163,In_81);
and U342 (N_342,In_1365,In_1238);
nand U343 (N_343,In_171,In_663);
or U344 (N_344,In_936,In_217);
nand U345 (N_345,In_809,In_1122);
or U346 (N_346,In_180,In_1021);
or U347 (N_347,In_1093,In_305);
nand U348 (N_348,In_1386,In_1055);
nand U349 (N_349,In_777,In_93);
and U350 (N_350,In_849,In_47);
and U351 (N_351,In_380,In_27);
nand U352 (N_352,In_700,In_539);
and U353 (N_353,In_3,In_449);
nor U354 (N_354,In_1275,In_1183);
or U355 (N_355,In_1438,In_1461);
xor U356 (N_356,In_757,In_109);
nand U357 (N_357,In_1012,In_340);
or U358 (N_358,In_105,In_626);
nor U359 (N_359,In_439,In_385);
and U360 (N_360,In_1119,In_694);
or U361 (N_361,In_711,In_1471);
and U362 (N_362,In_2,In_729);
nand U363 (N_363,In_589,In_257);
nor U364 (N_364,In_813,In_579);
nor U365 (N_365,In_873,In_141);
nand U366 (N_366,In_1424,In_923);
and U367 (N_367,In_1008,In_724);
xnor U368 (N_368,In_164,In_542);
nand U369 (N_369,In_1357,In_746);
or U370 (N_370,In_929,In_1290);
nor U371 (N_371,In_1044,In_1284);
xnor U372 (N_372,In_1221,In_398);
or U373 (N_373,In_676,In_1397);
or U374 (N_374,In_1224,In_1233);
and U375 (N_375,In_1161,In_417);
nand U376 (N_376,In_1366,In_1344);
or U377 (N_377,In_781,In_937);
or U378 (N_378,In_555,In_1342);
or U379 (N_379,In_52,In_751);
nor U380 (N_380,In_1405,In_1358);
nor U381 (N_381,In_328,In_1079);
nor U382 (N_382,In_1352,In_1213);
nand U383 (N_383,In_309,In_1439);
nor U384 (N_384,In_1490,In_886);
nor U385 (N_385,In_503,In_942);
or U386 (N_386,In_468,In_634);
or U387 (N_387,In_1285,In_409);
xnor U388 (N_388,In_1173,In_394);
and U389 (N_389,In_1179,In_747);
nor U390 (N_390,In_920,In_410);
nor U391 (N_391,In_577,In_260);
nor U392 (N_392,In_1402,In_1428);
xor U393 (N_393,In_769,In_762);
xnor U394 (N_394,In_1474,In_947);
nor U395 (N_395,In_207,In_855);
and U396 (N_396,In_229,In_1303);
and U397 (N_397,In_1020,In_214);
nand U398 (N_398,In_986,In_955);
nand U399 (N_399,In_462,In_183);
nand U400 (N_400,In_1120,In_448);
and U401 (N_401,In_819,In_68);
nor U402 (N_402,In_1331,In_812);
xnor U403 (N_403,In_871,In_1369);
nor U404 (N_404,In_896,In_31);
nor U405 (N_405,In_1228,In_437);
nand U406 (N_406,In_53,In_898);
nor U407 (N_407,In_1379,In_1229);
nor U408 (N_408,In_639,In_990);
and U409 (N_409,In_440,In_345);
and U410 (N_410,In_73,In_1479);
xor U411 (N_411,In_1222,In_483);
or U412 (N_412,In_284,In_1427);
nand U413 (N_413,In_1053,In_509);
nand U414 (N_414,In_901,In_977);
or U415 (N_415,In_332,In_405);
xnor U416 (N_416,In_1488,In_823);
nor U417 (N_417,In_868,In_238);
nor U418 (N_418,In_641,In_227);
xor U419 (N_419,In_271,In_452);
and U420 (N_420,In_553,In_685);
or U421 (N_421,In_333,In_1273);
nand U422 (N_422,In_450,In_928);
nor U423 (N_423,In_1006,In_1111);
nor U424 (N_424,In_134,In_1069);
nor U425 (N_425,In_1153,In_1407);
nor U426 (N_426,In_562,In_616);
and U427 (N_427,In_540,In_185);
and U428 (N_428,In_11,In_454);
and U429 (N_429,In_1184,In_374);
nor U430 (N_430,In_1029,In_356);
and U431 (N_431,In_1022,In_620);
nor U432 (N_432,In_621,In_461);
and U433 (N_433,In_891,In_378);
and U434 (N_434,In_362,In_201);
nand U435 (N_435,In_558,In_1219);
xnor U436 (N_436,In_1389,In_576);
xnor U437 (N_437,In_969,In_464);
nand U438 (N_438,In_153,In_1460);
or U439 (N_439,In_1381,In_62);
and U440 (N_440,In_650,In_1144);
nand U441 (N_441,In_523,In_885);
and U442 (N_442,In_658,In_1404);
nor U443 (N_443,In_1089,In_874);
xor U444 (N_444,In_1118,In_210);
nor U445 (N_445,In_1392,In_100);
and U446 (N_446,In_1036,In_475);
and U447 (N_447,In_1242,In_1071);
xnor U448 (N_448,In_852,In_1085);
nor U449 (N_449,In_403,In_1336);
xor U450 (N_450,In_1322,In_1390);
nor U451 (N_451,In_1138,In_1466);
nand U452 (N_452,In_557,In_890);
or U453 (N_453,In_913,In_1434);
nor U454 (N_454,In_1199,In_703);
nor U455 (N_455,In_1172,In_224);
xnor U456 (N_456,In_441,In_208);
or U457 (N_457,In_115,In_314);
nand U458 (N_458,In_176,In_903);
or U459 (N_459,In_466,In_203);
or U460 (N_460,In_1230,In_41);
nor U461 (N_461,In_892,In_1211);
or U462 (N_462,In_110,In_767);
and U463 (N_463,In_276,In_391);
or U464 (N_464,In_373,In_832);
and U465 (N_465,In_1003,In_98);
xnor U466 (N_466,In_118,In_1152);
nor U467 (N_467,In_938,In_878);
nand U468 (N_468,In_683,In_1041);
nand U469 (N_469,In_123,In_802);
and U470 (N_470,In_584,In_418);
nor U471 (N_471,In_1064,In_846);
nand U472 (N_472,In_563,In_1293);
xor U473 (N_473,In_1355,In_298);
and U474 (N_474,In_372,In_1092);
nand U475 (N_475,In_692,In_962);
nand U476 (N_476,In_1360,In_1409);
nand U477 (N_477,In_771,In_899);
nand U478 (N_478,In_139,In_1347);
and U479 (N_479,In_502,In_116);
and U480 (N_480,In_1167,In_213);
or U481 (N_481,In_617,In_1132);
and U482 (N_482,In_1078,In_1493);
or U483 (N_483,In_708,In_678);
nand U484 (N_484,In_776,In_1408);
nand U485 (N_485,In_637,In_1308);
xor U486 (N_486,In_1320,In_1316);
nor U487 (N_487,In_722,In_1445);
and U488 (N_488,In_671,In_733);
or U489 (N_489,In_1099,In_162);
or U490 (N_490,In_245,In_360);
nand U491 (N_491,In_359,In_743);
nor U492 (N_492,In_504,In_1);
nor U493 (N_493,In_482,In_1296);
nor U494 (N_494,In_796,In_370);
nor U495 (N_495,In_1004,In_1262);
and U496 (N_496,In_261,In_469);
nor U497 (N_497,In_287,In_416);
xnor U498 (N_498,In_905,In_323);
or U499 (N_499,In_313,In_833);
nor U500 (N_500,In_807,In_714);
or U501 (N_501,In_554,In_611);
nand U502 (N_502,In_1105,In_1450);
or U503 (N_503,In_1294,In_38);
or U504 (N_504,In_749,In_798);
nor U505 (N_505,In_243,In_1236);
nor U506 (N_506,In_159,In_1165);
and U507 (N_507,In_1272,In_1291);
nor U508 (N_508,In_194,In_670);
nand U509 (N_509,In_250,In_289);
nor U510 (N_510,In_748,In_154);
nor U511 (N_511,In_479,In_718);
and U512 (N_512,In_808,In_1276);
nand U513 (N_513,In_117,In_790);
nor U514 (N_514,In_716,In_839);
and U515 (N_515,In_1459,In_388);
or U516 (N_516,In_1310,In_1353);
nand U517 (N_517,In_54,In_354);
or U518 (N_518,In_1244,In_521);
xor U519 (N_519,In_632,In_1169);
nor U520 (N_520,In_1359,In_811);
nand U521 (N_521,In_1107,In_1457);
or U522 (N_522,In_643,In_1448);
and U523 (N_523,In_7,In_754);
nor U524 (N_524,In_107,In_42);
nand U525 (N_525,In_917,In_6);
nand U526 (N_526,In_657,In_251);
nor U527 (N_527,In_470,In_230);
nand U528 (N_528,In_1001,In_272);
and U529 (N_529,In_244,In_487);
nand U530 (N_530,In_211,In_283);
xnor U531 (N_531,In_1391,In_734);
nand U532 (N_532,In_831,In_665);
nand U533 (N_533,In_838,In_699);
nor U534 (N_534,In_220,In_423);
nand U535 (N_535,In_363,In_277);
and U536 (N_536,In_346,In_406);
and U537 (N_537,In_79,In_591);
nand U538 (N_538,In_148,In_546);
nand U539 (N_539,In_686,In_155);
and U540 (N_540,In_178,In_527);
nor U541 (N_541,In_1364,In_149);
nand U542 (N_542,In_144,In_55);
xnor U543 (N_543,In_357,In_1394);
nand U544 (N_544,In_926,In_1487);
nand U545 (N_545,In_730,In_1453);
or U546 (N_546,In_1149,In_1057);
or U547 (N_547,In_609,In_627);
nor U548 (N_548,In_511,In_400);
nand U549 (N_549,In_1260,In_1065);
and U550 (N_550,In_428,In_173);
xor U551 (N_551,In_970,In_550);
and U552 (N_552,In_1309,In_992);
nand U553 (N_553,In_87,In_331);
and U554 (N_554,In_568,In_1194);
and U555 (N_555,In_262,In_745);
or U556 (N_556,In_1154,In_837);
or U557 (N_557,In_614,In_739);
xor U558 (N_558,In_412,In_1410);
and U559 (N_559,In_644,In_687);
xor U560 (N_560,In_1074,In_215);
or U561 (N_561,In_1214,In_18);
nor U562 (N_562,In_1035,In_188);
nor U563 (N_563,In_635,In_814);
or U564 (N_564,In_446,In_256);
nand U565 (N_565,In_447,In_19);
nor U566 (N_566,In_816,In_1158);
xnor U567 (N_567,In_325,In_572);
nor U568 (N_568,In_1240,In_170);
and U569 (N_569,In_848,In_758);
and U570 (N_570,In_221,In_1193);
and U571 (N_571,In_274,In_1441);
xnor U572 (N_572,In_1476,In_994);
or U573 (N_573,In_505,In_594);
or U574 (N_574,In_981,In_1281);
nor U575 (N_575,In_1011,In_112);
nand U576 (N_576,In_628,In_800);
nand U577 (N_577,In_1106,In_1206);
nand U578 (N_578,In_1042,In_506);
or U579 (N_579,In_1025,In_300);
nor U580 (N_580,In_1133,In_750);
and U581 (N_581,In_1465,In_143);
nand U582 (N_582,In_1121,In_702);
nand U583 (N_583,In_1082,In_106);
nand U584 (N_584,In_978,In_1307);
nand U585 (N_585,In_508,In_179);
nand U586 (N_586,In_1452,In_940);
nand U587 (N_587,In_761,In_935);
nor U588 (N_588,In_677,In_1060);
nand U589 (N_589,In_367,In_519);
or U590 (N_590,In_317,In_1187);
and U591 (N_591,In_1387,In_1166);
or U592 (N_592,In_1449,In_1299);
or U593 (N_593,In_909,In_1345);
nand U594 (N_594,In_538,In_228);
or U595 (N_595,In_216,In_1388);
nand U596 (N_596,In_1396,In_736);
or U597 (N_597,In_664,In_88);
or U598 (N_598,In_530,In_189);
nand U599 (N_599,In_186,In_1377);
xnor U600 (N_600,In_1247,In_565);
and U601 (N_601,In_23,In_675);
and U602 (N_602,In_785,In_335);
nand U603 (N_603,In_1393,In_1164);
nand U604 (N_604,In_324,In_1070);
nand U605 (N_605,In_1124,In_65);
and U606 (N_606,In_393,In_1162);
nand U607 (N_607,In_1496,In_1174);
or U608 (N_608,In_1373,In_1384);
nand U609 (N_609,In_192,In_801);
xnor U610 (N_610,In_1195,In_780);
or U611 (N_611,In_933,In_168);
nand U612 (N_612,In_212,In_1215);
or U613 (N_613,In_1253,In_1333);
and U614 (N_614,In_308,In_516);
or U615 (N_615,In_513,In_1005);
xnor U616 (N_616,In_320,In_599);
and U617 (N_617,In_1491,In_125);
nor U618 (N_618,In_1443,In_971);
or U619 (N_619,In_1059,In_1077);
or U620 (N_620,In_96,In_442);
and U621 (N_621,In_1227,In_140);
nand U622 (N_622,In_1050,In_1426);
nand U623 (N_623,In_160,In_622);
or U624 (N_624,In_330,In_654);
or U625 (N_625,In_853,In_1180);
nor U626 (N_626,In_1354,In_72);
or U627 (N_627,In_402,In_495);
and U628 (N_628,In_646,In_195);
and U629 (N_629,In_389,In_884);
xor U630 (N_630,In_1100,In_259);
and U631 (N_631,In_95,In_946);
or U632 (N_632,In_1361,In_845);
nor U633 (N_633,In_725,In_795);
nor U634 (N_634,In_498,In_14);
and U635 (N_635,In_375,In_927);
nand U636 (N_636,In_541,In_1128);
and U637 (N_637,In_1469,In_914);
or U638 (N_638,In_825,In_973);
nor U639 (N_639,In_993,In_1066);
and U640 (N_640,In_570,In_1351);
or U641 (N_641,In_810,In_384);
nand U642 (N_642,In_392,In_1038);
and U643 (N_643,In_310,In_161);
or U644 (N_644,In_293,In_253);
nand U645 (N_645,In_1375,In_35);
nand U646 (N_646,In_480,In_548);
and U647 (N_647,In_1013,In_763);
and U648 (N_648,In_489,In_1411);
and U649 (N_649,In_264,In_114);
nor U650 (N_650,In_1030,In_921);
and U651 (N_651,In_952,In_1420);
or U652 (N_652,In_939,In_1126);
and U653 (N_653,In_458,In_1282);
and U654 (N_654,In_1234,In_1324);
nor U655 (N_655,In_659,In_275);
nor U656 (N_656,In_1088,In_1485);
nor U657 (N_657,In_906,In_1327);
or U658 (N_658,In_273,In_285);
nor U659 (N_659,In_1486,In_1400);
or U660 (N_660,In_64,In_544);
nor U661 (N_661,In_666,In_865);
nand U662 (N_662,In_1114,In_1087);
nor U663 (N_663,In_304,In_571);
nor U664 (N_664,In_526,In_881);
and U665 (N_665,In_537,In_787);
nand U666 (N_666,In_13,In_1061);
and U667 (N_667,In_1159,In_525);
and U668 (N_668,In_1103,In_1288);
nor U669 (N_669,In_587,In_1143);
or U670 (N_670,In_738,In_1134);
nand U671 (N_671,In_945,In_296);
xor U672 (N_672,In_1190,In_601);
nor U673 (N_673,In_615,In_759);
xnor U674 (N_674,In_704,In_515);
or U675 (N_675,In_5,In_1385);
or U676 (N_676,In_593,In_715);
nand U677 (N_677,In_311,In_1455);
xnor U678 (N_678,In_661,In_961);
nand U679 (N_679,In_597,In_94);
nand U680 (N_680,In_860,In_383);
nand U681 (N_681,In_789,In_102);
or U682 (N_682,In_956,In_361);
or U683 (N_683,In_1422,In_414);
and U684 (N_684,In_1306,In_1015);
nand U685 (N_685,In_348,In_1329);
or U686 (N_686,In_1202,In_1268);
or U687 (N_687,In_803,In_175);
xor U688 (N_688,In_979,In_879);
xor U689 (N_689,In_326,In_1425);
or U690 (N_690,In_948,In_682);
nand U691 (N_691,In_669,In_1463);
and U692 (N_692,In_1217,In_660);
or U693 (N_693,In_263,In_705);
nand U694 (N_694,In_1497,In_528);
nand U695 (N_695,In_710,In_1269);
nand U696 (N_696,In_507,In_1374);
or U697 (N_697,In_408,In_404);
nand U698 (N_698,In_1270,In_278);
nand U699 (N_699,In_424,In_844);
nand U700 (N_700,In_1178,In_1350);
and U701 (N_701,In_720,In_1289);
nor U702 (N_702,In_45,In_1058);
nor U703 (N_703,In_877,In_1467);
nand U704 (N_704,In_1287,In_1256);
and U705 (N_705,In_307,In_488);
nor U706 (N_706,In_964,In_1311);
and U707 (N_707,In_199,In_1155);
and U708 (N_708,In_322,In_728);
nor U709 (N_709,In_864,In_1295);
nand U710 (N_710,In_80,In_723);
and U711 (N_711,In_1376,In_1210);
nor U712 (N_712,In_695,In_875);
xnor U713 (N_713,In_1123,In_426);
and U714 (N_714,In_1492,In_1150);
nor U715 (N_715,In_680,In_551);
nor U716 (N_716,In_1312,In_1255);
nor U717 (N_717,In_774,In_120);
nor U718 (N_718,In_688,In_1084);
or U719 (N_719,In_791,In_655);
nor U720 (N_720,In_342,In_187);
and U721 (N_721,In_151,In_390);
or U722 (N_722,In_36,In_471);
or U723 (N_723,In_775,In_996);
and U724 (N_724,In_344,In_1248);
nor U725 (N_725,In_1499,In_1252);
nor U726 (N_726,In_167,In_236);
and U727 (N_727,In_1073,In_752);
and U728 (N_728,In_820,In_1241);
and U729 (N_729,In_772,In_132);
xor U730 (N_730,In_301,In_603);
nand U731 (N_731,In_499,In_1239);
or U732 (N_732,In_1112,In_1489);
nor U733 (N_733,In_147,In_119);
nor U734 (N_734,In_1332,In_86);
and U735 (N_735,In_1204,In_863);
or U736 (N_736,In_465,In_640);
nand U737 (N_737,In_982,In_869);
nand U738 (N_738,In_602,In_862);
xnor U739 (N_739,In_9,In_460);
nand U740 (N_740,In_177,In_267);
and U741 (N_741,In_91,In_1130);
or U742 (N_742,In_1196,In_1472);
nand U743 (N_743,In_1325,In_672);
or U744 (N_744,In_435,In_341);
or U745 (N_745,In_1068,In_239);
or U746 (N_746,In_193,In_953);
or U747 (N_747,In_1446,In_691);
xor U748 (N_748,In_1148,In_1220);
nor U749 (N_749,In_433,In_910);
or U750 (N_750,In_1412,In_242);
xor U751 (N_751,In_1424,In_80);
nor U752 (N_752,In_1429,In_911);
and U753 (N_753,In_1189,In_465);
nand U754 (N_754,In_1222,In_68);
and U755 (N_755,In_1190,In_1417);
or U756 (N_756,In_48,In_116);
nand U757 (N_757,In_532,In_616);
or U758 (N_758,In_894,In_255);
or U759 (N_759,In_729,In_1071);
xnor U760 (N_760,In_531,In_1290);
and U761 (N_761,In_411,In_574);
nor U762 (N_762,In_1384,In_1231);
and U763 (N_763,In_271,In_1430);
nand U764 (N_764,In_395,In_259);
and U765 (N_765,In_1355,In_766);
and U766 (N_766,In_198,In_1027);
or U767 (N_767,In_235,In_1386);
nor U768 (N_768,In_1300,In_766);
xor U769 (N_769,In_290,In_680);
and U770 (N_770,In_1343,In_239);
xnor U771 (N_771,In_874,In_1100);
nand U772 (N_772,In_1156,In_1397);
nor U773 (N_773,In_1056,In_147);
and U774 (N_774,In_83,In_750);
nand U775 (N_775,In_42,In_599);
xor U776 (N_776,In_610,In_297);
xor U777 (N_777,In_925,In_157);
nor U778 (N_778,In_665,In_600);
nor U779 (N_779,In_1027,In_368);
nor U780 (N_780,In_867,In_1345);
and U781 (N_781,In_800,In_355);
nor U782 (N_782,In_1309,In_700);
or U783 (N_783,In_1444,In_159);
nor U784 (N_784,In_762,In_468);
nor U785 (N_785,In_743,In_517);
or U786 (N_786,In_12,In_38);
nor U787 (N_787,In_1102,In_629);
xnor U788 (N_788,In_1324,In_968);
nor U789 (N_789,In_1313,In_1459);
and U790 (N_790,In_968,In_1397);
nor U791 (N_791,In_567,In_459);
or U792 (N_792,In_388,In_447);
or U793 (N_793,In_940,In_1291);
xnor U794 (N_794,In_266,In_478);
and U795 (N_795,In_154,In_650);
nand U796 (N_796,In_317,In_483);
xor U797 (N_797,In_1490,In_585);
nor U798 (N_798,In_530,In_351);
nand U799 (N_799,In_1241,In_1407);
or U800 (N_800,In_1052,In_1242);
nand U801 (N_801,In_628,In_1041);
nor U802 (N_802,In_86,In_266);
and U803 (N_803,In_606,In_283);
or U804 (N_804,In_491,In_393);
or U805 (N_805,In_649,In_2);
or U806 (N_806,In_64,In_491);
nand U807 (N_807,In_355,In_779);
nand U808 (N_808,In_1324,In_975);
or U809 (N_809,In_1247,In_108);
nand U810 (N_810,In_1341,In_114);
nor U811 (N_811,In_711,In_557);
or U812 (N_812,In_301,In_311);
nor U813 (N_813,In_1390,In_566);
nor U814 (N_814,In_1258,In_1485);
nand U815 (N_815,In_675,In_748);
nor U816 (N_816,In_539,In_918);
xnor U817 (N_817,In_1215,In_1094);
nand U818 (N_818,In_1182,In_153);
and U819 (N_819,In_1255,In_707);
nor U820 (N_820,In_830,In_1024);
nand U821 (N_821,In_876,In_183);
nor U822 (N_822,In_1139,In_263);
and U823 (N_823,In_641,In_1234);
nand U824 (N_824,In_114,In_744);
and U825 (N_825,In_832,In_120);
nand U826 (N_826,In_1495,In_723);
nand U827 (N_827,In_299,In_1395);
or U828 (N_828,In_1237,In_739);
nor U829 (N_829,In_774,In_1147);
or U830 (N_830,In_819,In_1347);
nand U831 (N_831,In_808,In_430);
or U832 (N_832,In_1389,In_264);
or U833 (N_833,In_491,In_1394);
nor U834 (N_834,In_1380,In_733);
nor U835 (N_835,In_713,In_759);
nand U836 (N_836,In_523,In_1334);
nor U837 (N_837,In_553,In_1185);
nand U838 (N_838,In_450,In_1108);
nor U839 (N_839,In_639,In_163);
or U840 (N_840,In_1158,In_1149);
and U841 (N_841,In_1154,In_509);
and U842 (N_842,In_255,In_70);
nand U843 (N_843,In_1362,In_1443);
nand U844 (N_844,In_1037,In_496);
nand U845 (N_845,In_1338,In_154);
nor U846 (N_846,In_1251,In_1148);
and U847 (N_847,In_754,In_1209);
and U848 (N_848,In_442,In_1038);
xor U849 (N_849,In_619,In_1105);
xor U850 (N_850,In_867,In_518);
or U851 (N_851,In_841,In_326);
and U852 (N_852,In_670,In_307);
or U853 (N_853,In_543,In_753);
nor U854 (N_854,In_351,In_547);
nor U855 (N_855,In_839,In_119);
or U856 (N_856,In_46,In_25);
and U857 (N_857,In_365,In_406);
nand U858 (N_858,In_1330,In_817);
nand U859 (N_859,In_779,In_474);
nor U860 (N_860,In_1136,In_688);
nand U861 (N_861,In_1448,In_1065);
xor U862 (N_862,In_588,In_955);
nor U863 (N_863,In_620,In_1331);
and U864 (N_864,In_126,In_918);
nor U865 (N_865,In_558,In_1078);
or U866 (N_866,In_801,In_935);
and U867 (N_867,In_613,In_806);
or U868 (N_868,In_65,In_356);
nand U869 (N_869,In_738,In_1251);
nor U870 (N_870,In_848,In_666);
and U871 (N_871,In_610,In_1041);
xor U872 (N_872,In_1165,In_893);
nor U873 (N_873,In_514,In_1496);
nor U874 (N_874,In_1185,In_509);
or U875 (N_875,In_447,In_85);
nor U876 (N_876,In_112,In_39);
nor U877 (N_877,In_1481,In_950);
nor U878 (N_878,In_109,In_103);
or U879 (N_879,In_4,In_494);
or U880 (N_880,In_300,In_864);
or U881 (N_881,In_647,In_944);
and U882 (N_882,In_881,In_277);
xnor U883 (N_883,In_367,In_1328);
or U884 (N_884,In_601,In_375);
xnor U885 (N_885,In_1284,In_1028);
xor U886 (N_886,In_456,In_1421);
xor U887 (N_887,In_955,In_1000);
nand U888 (N_888,In_205,In_51);
nand U889 (N_889,In_376,In_963);
nand U890 (N_890,In_1297,In_1432);
and U891 (N_891,In_550,In_1263);
and U892 (N_892,In_533,In_374);
or U893 (N_893,In_591,In_279);
and U894 (N_894,In_251,In_23);
nor U895 (N_895,In_826,In_310);
nor U896 (N_896,In_303,In_53);
or U897 (N_897,In_899,In_100);
and U898 (N_898,In_330,In_933);
nor U899 (N_899,In_754,In_210);
nand U900 (N_900,In_930,In_653);
or U901 (N_901,In_448,In_1261);
nor U902 (N_902,In_757,In_865);
nand U903 (N_903,In_308,In_74);
nor U904 (N_904,In_1324,In_191);
nand U905 (N_905,In_128,In_1107);
nand U906 (N_906,In_638,In_685);
and U907 (N_907,In_987,In_1463);
and U908 (N_908,In_405,In_81);
nand U909 (N_909,In_1242,In_806);
nand U910 (N_910,In_947,In_419);
nor U911 (N_911,In_206,In_818);
or U912 (N_912,In_659,In_219);
and U913 (N_913,In_367,In_692);
and U914 (N_914,In_742,In_437);
nand U915 (N_915,In_1259,In_56);
nand U916 (N_916,In_74,In_593);
or U917 (N_917,In_136,In_1027);
or U918 (N_918,In_1348,In_952);
xor U919 (N_919,In_1194,In_1478);
or U920 (N_920,In_356,In_606);
nor U921 (N_921,In_681,In_467);
nand U922 (N_922,In_644,In_819);
or U923 (N_923,In_736,In_68);
and U924 (N_924,In_750,In_522);
nand U925 (N_925,In_142,In_752);
or U926 (N_926,In_1177,In_1383);
xnor U927 (N_927,In_558,In_385);
and U928 (N_928,In_587,In_185);
nor U929 (N_929,In_1190,In_971);
or U930 (N_930,In_1397,In_1430);
or U931 (N_931,In_1171,In_551);
nand U932 (N_932,In_525,In_1360);
nor U933 (N_933,In_865,In_1339);
or U934 (N_934,In_120,In_1069);
nand U935 (N_935,In_1411,In_236);
nand U936 (N_936,In_915,In_391);
or U937 (N_937,In_152,In_1312);
and U938 (N_938,In_240,In_574);
nand U939 (N_939,In_915,In_276);
nor U940 (N_940,In_232,In_870);
nand U941 (N_941,In_135,In_564);
and U942 (N_942,In_1440,In_1398);
nand U943 (N_943,In_853,In_180);
and U944 (N_944,In_281,In_709);
nor U945 (N_945,In_855,In_728);
or U946 (N_946,In_478,In_902);
nor U947 (N_947,In_739,In_766);
and U948 (N_948,In_933,In_1210);
xor U949 (N_949,In_857,In_1147);
nor U950 (N_950,In_825,In_1150);
nand U951 (N_951,In_872,In_1160);
nand U952 (N_952,In_213,In_237);
xnor U953 (N_953,In_1124,In_231);
nor U954 (N_954,In_1165,In_665);
or U955 (N_955,In_363,In_105);
nor U956 (N_956,In_1143,In_952);
and U957 (N_957,In_1332,In_1331);
and U958 (N_958,In_1441,In_1042);
or U959 (N_959,In_300,In_875);
or U960 (N_960,In_318,In_1371);
nand U961 (N_961,In_400,In_369);
nor U962 (N_962,In_757,In_742);
nand U963 (N_963,In_1215,In_965);
or U964 (N_964,In_1177,In_673);
nand U965 (N_965,In_1480,In_1307);
nand U966 (N_966,In_1056,In_433);
nor U967 (N_967,In_510,In_630);
nand U968 (N_968,In_331,In_537);
and U969 (N_969,In_1403,In_239);
and U970 (N_970,In_1059,In_1213);
nand U971 (N_971,In_1400,In_1464);
or U972 (N_972,In_608,In_424);
and U973 (N_973,In_106,In_1098);
nand U974 (N_974,In_101,In_921);
nand U975 (N_975,In_942,In_680);
and U976 (N_976,In_387,In_1497);
or U977 (N_977,In_200,In_332);
xnor U978 (N_978,In_1208,In_409);
nand U979 (N_979,In_571,In_448);
nor U980 (N_980,In_1339,In_876);
nor U981 (N_981,In_61,In_674);
nand U982 (N_982,In_933,In_881);
nand U983 (N_983,In_1120,In_1388);
and U984 (N_984,In_227,In_970);
nand U985 (N_985,In_240,In_40);
or U986 (N_986,In_1412,In_499);
nor U987 (N_987,In_153,In_984);
nand U988 (N_988,In_762,In_646);
nor U989 (N_989,In_1021,In_1371);
nand U990 (N_990,In_457,In_743);
nand U991 (N_991,In_1261,In_300);
and U992 (N_992,In_321,In_188);
and U993 (N_993,In_859,In_862);
or U994 (N_994,In_1306,In_606);
or U995 (N_995,In_1234,In_242);
nor U996 (N_996,In_1219,In_1167);
and U997 (N_997,In_50,In_1110);
nor U998 (N_998,In_1422,In_1433);
nand U999 (N_999,In_799,In_168);
or U1000 (N_1000,In_379,In_442);
nand U1001 (N_1001,In_753,In_166);
or U1002 (N_1002,In_719,In_579);
nor U1003 (N_1003,In_534,In_1330);
xor U1004 (N_1004,In_224,In_1307);
nor U1005 (N_1005,In_1023,In_1247);
nor U1006 (N_1006,In_1182,In_1141);
and U1007 (N_1007,In_17,In_194);
nand U1008 (N_1008,In_953,In_1451);
and U1009 (N_1009,In_354,In_610);
or U1010 (N_1010,In_221,In_1139);
nand U1011 (N_1011,In_1408,In_1291);
and U1012 (N_1012,In_1255,In_58);
nand U1013 (N_1013,In_46,In_1172);
nor U1014 (N_1014,In_449,In_844);
and U1015 (N_1015,In_1233,In_450);
and U1016 (N_1016,In_481,In_837);
or U1017 (N_1017,In_273,In_815);
and U1018 (N_1018,In_736,In_104);
and U1019 (N_1019,In_1192,In_355);
nor U1020 (N_1020,In_91,In_160);
or U1021 (N_1021,In_984,In_675);
nand U1022 (N_1022,In_310,In_323);
nand U1023 (N_1023,In_540,In_1210);
and U1024 (N_1024,In_211,In_409);
nand U1025 (N_1025,In_1227,In_1114);
or U1026 (N_1026,In_419,In_877);
and U1027 (N_1027,In_330,In_1337);
nand U1028 (N_1028,In_1371,In_539);
and U1029 (N_1029,In_467,In_269);
xor U1030 (N_1030,In_1479,In_475);
xnor U1031 (N_1031,In_103,In_130);
nor U1032 (N_1032,In_1151,In_494);
nor U1033 (N_1033,In_1265,In_331);
and U1034 (N_1034,In_409,In_727);
nand U1035 (N_1035,In_1361,In_1280);
nor U1036 (N_1036,In_1032,In_1402);
and U1037 (N_1037,In_871,In_478);
nor U1038 (N_1038,In_1488,In_1016);
nor U1039 (N_1039,In_494,In_646);
nor U1040 (N_1040,In_1118,In_388);
nor U1041 (N_1041,In_308,In_598);
nor U1042 (N_1042,In_1382,In_434);
nor U1043 (N_1043,In_758,In_1374);
nor U1044 (N_1044,In_586,In_684);
or U1045 (N_1045,In_1118,In_780);
xnor U1046 (N_1046,In_1407,In_799);
nand U1047 (N_1047,In_1269,In_1393);
xor U1048 (N_1048,In_509,In_1048);
and U1049 (N_1049,In_1171,In_644);
xor U1050 (N_1050,In_609,In_372);
xnor U1051 (N_1051,In_908,In_450);
nor U1052 (N_1052,In_395,In_1060);
nand U1053 (N_1053,In_640,In_850);
and U1054 (N_1054,In_533,In_736);
nand U1055 (N_1055,In_1215,In_940);
or U1056 (N_1056,In_1228,In_751);
or U1057 (N_1057,In_550,In_1136);
or U1058 (N_1058,In_1306,In_154);
nor U1059 (N_1059,In_875,In_366);
nand U1060 (N_1060,In_908,In_976);
or U1061 (N_1061,In_664,In_40);
nand U1062 (N_1062,In_1267,In_630);
or U1063 (N_1063,In_663,In_946);
or U1064 (N_1064,In_486,In_1343);
nor U1065 (N_1065,In_1345,In_333);
nor U1066 (N_1066,In_569,In_431);
or U1067 (N_1067,In_1277,In_1137);
nor U1068 (N_1068,In_120,In_611);
and U1069 (N_1069,In_526,In_759);
and U1070 (N_1070,In_48,In_602);
nand U1071 (N_1071,In_187,In_524);
and U1072 (N_1072,In_801,In_364);
nor U1073 (N_1073,In_783,In_50);
nand U1074 (N_1074,In_27,In_1296);
nand U1075 (N_1075,In_323,In_152);
nand U1076 (N_1076,In_1356,In_708);
nand U1077 (N_1077,In_35,In_1101);
nand U1078 (N_1078,In_512,In_369);
xor U1079 (N_1079,In_562,In_1254);
and U1080 (N_1080,In_480,In_1334);
and U1081 (N_1081,In_65,In_1409);
xnor U1082 (N_1082,In_787,In_1373);
and U1083 (N_1083,In_810,In_166);
or U1084 (N_1084,In_1106,In_1037);
or U1085 (N_1085,In_43,In_1316);
and U1086 (N_1086,In_176,In_1307);
and U1087 (N_1087,In_593,In_856);
nand U1088 (N_1088,In_443,In_1010);
xor U1089 (N_1089,In_1469,In_1028);
or U1090 (N_1090,In_790,In_32);
or U1091 (N_1091,In_741,In_1476);
nand U1092 (N_1092,In_1104,In_1107);
nor U1093 (N_1093,In_227,In_5);
xor U1094 (N_1094,In_923,In_606);
or U1095 (N_1095,In_1495,In_128);
xor U1096 (N_1096,In_1132,In_313);
or U1097 (N_1097,In_1078,In_1479);
and U1098 (N_1098,In_710,In_1177);
and U1099 (N_1099,In_518,In_569);
nor U1100 (N_1100,In_244,In_303);
nor U1101 (N_1101,In_1470,In_1035);
and U1102 (N_1102,In_1335,In_848);
nand U1103 (N_1103,In_139,In_27);
nor U1104 (N_1104,In_437,In_21);
nor U1105 (N_1105,In_358,In_757);
nor U1106 (N_1106,In_1194,In_1174);
and U1107 (N_1107,In_1210,In_1303);
nand U1108 (N_1108,In_159,In_244);
nand U1109 (N_1109,In_958,In_975);
xnor U1110 (N_1110,In_809,In_1085);
nand U1111 (N_1111,In_135,In_1305);
or U1112 (N_1112,In_1052,In_221);
or U1113 (N_1113,In_831,In_1380);
nor U1114 (N_1114,In_474,In_417);
and U1115 (N_1115,In_1107,In_1216);
nor U1116 (N_1116,In_479,In_704);
or U1117 (N_1117,In_680,In_96);
or U1118 (N_1118,In_24,In_76);
nand U1119 (N_1119,In_312,In_1359);
nor U1120 (N_1120,In_230,In_472);
or U1121 (N_1121,In_1225,In_1114);
nor U1122 (N_1122,In_845,In_508);
and U1123 (N_1123,In_713,In_1241);
xnor U1124 (N_1124,In_805,In_370);
or U1125 (N_1125,In_277,In_547);
or U1126 (N_1126,In_626,In_98);
nand U1127 (N_1127,In_41,In_1287);
nand U1128 (N_1128,In_612,In_978);
or U1129 (N_1129,In_791,In_291);
and U1130 (N_1130,In_132,In_1042);
or U1131 (N_1131,In_170,In_1107);
nand U1132 (N_1132,In_604,In_1120);
or U1133 (N_1133,In_1254,In_503);
nor U1134 (N_1134,In_1299,In_79);
nor U1135 (N_1135,In_1003,In_81);
nor U1136 (N_1136,In_954,In_929);
nand U1137 (N_1137,In_623,In_1095);
or U1138 (N_1138,In_380,In_1337);
nand U1139 (N_1139,In_1029,In_657);
nor U1140 (N_1140,In_624,In_1052);
nor U1141 (N_1141,In_436,In_605);
and U1142 (N_1142,In_884,In_538);
and U1143 (N_1143,In_1426,In_1119);
nand U1144 (N_1144,In_717,In_1323);
and U1145 (N_1145,In_655,In_904);
and U1146 (N_1146,In_553,In_186);
and U1147 (N_1147,In_1,In_553);
and U1148 (N_1148,In_994,In_1356);
or U1149 (N_1149,In_811,In_508);
or U1150 (N_1150,In_225,In_1022);
nand U1151 (N_1151,In_2,In_1397);
xor U1152 (N_1152,In_965,In_487);
xor U1153 (N_1153,In_1429,In_248);
or U1154 (N_1154,In_567,In_144);
nor U1155 (N_1155,In_628,In_1458);
or U1156 (N_1156,In_1301,In_886);
nand U1157 (N_1157,In_42,In_332);
nor U1158 (N_1158,In_1034,In_645);
or U1159 (N_1159,In_31,In_757);
and U1160 (N_1160,In_761,In_882);
or U1161 (N_1161,In_1142,In_1147);
and U1162 (N_1162,In_917,In_705);
or U1163 (N_1163,In_375,In_1086);
or U1164 (N_1164,In_86,In_282);
and U1165 (N_1165,In_1021,In_1440);
or U1166 (N_1166,In_255,In_166);
and U1167 (N_1167,In_1228,In_493);
nor U1168 (N_1168,In_663,In_725);
or U1169 (N_1169,In_543,In_1448);
nor U1170 (N_1170,In_1130,In_1165);
or U1171 (N_1171,In_712,In_350);
xnor U1172 (N_1172,In_1253,In_1126);
nor U1173 (N_1173,In_303,In_750);
nor U1174 (N_1174,In_124,In_1277);
nand U1175 (N_1175,In_28,In_797);
and U1176 (N_1176,In_945,In_1180);
or U1177 (N_1177,In_331,In_553);
or U1178 (N_1178,In_551,In_322);
xnor U1179 (N_1179,In_862,In_1495);
or U1180 (N_1180,In_1129,In_1378);
nor U1181 (N_1181,In_671,In_98);
nor U1182 (N_1182,In_175,In_525);
and U1183 (N_1183,In_938,In_729);
nor U1184 (N_1184,In_1302,In_611);
or U1185 (N_1185,In_752,In_1232);
nand U1186 (N_1186,In_231,In_1109);
or U1187 (N_1187,In_197,In_257);
or U1188 (N_1188,In_1128,In_936);
nand U1189 (N_1189,In_135,In_1033);
or U1190 (N_1190,In_863,In_1487);
or U1191 (N_1191,In_581,In_1105);
nor U1192 (N_1192,In_524,In_1118);
nand U1193 (N_1193,In_779,In_435);
and U1194 (N_1194,In_297,In_1188);
or U1195 (N_1195,In_65,In_1219);
nor U1196 (N_1196,In_375,In_965);
or U1197 (N_1197,In_240,In_844);
and U1198 (N_1198,In_612,In_521);
or U1199 (N_1199,In_1079,In_969);
nor U1200 (N_1200,In_1074,In_1431);
and U1201 (N_1201,In_1394,In_1018);
nand U1202 (N_1202,In_426,In_1066);
and U1203 (N_1203,In_32,In_188);
nor U1204 (N_1204,In_742,In_10);
nor U1205 (N_1205,In_512,In_964);
and U1206 (N_1206,In_403,In_609);
nand U1207 (N_1207,In_1176,In_872);
nand U1208 (N_1208,In_325,In_1340);
nor U1209 (N_1209,In_1238,In_1404);
or U1210 (N_1210,In_884,In_985);
nand U1211 (N_1211,In_1019,In_1280);
nor U1212 (N_1212,In_1367,In_873);
and U1213 (N_1213,In_1018,In_1317);
or U1214 (N_1214,In_776,In_408);
xor U1215 (N_1215,In_763,In_372);
nor U1216 (N_1216,In_1318,In_90);
or U1217 (N_1217,In_784,In_813);
xor U1218 (N_1218,In_1204,In_927);
nand U1219 (N_1219,In_1178,In_141);
nor U1220 (N_1220,In_1463,In_830);
nand U1221 (N_1221,In_474,In_1271);
nand U1222 (N_1222,In_37,In_831);
xor U1223 (N_1223,In_1097,In_1085);
nand U1224 (N_1224,In_730,In_968);
and U1225 (N_1225,In_371,In_678);
or U1226 (N_1226,In_1320,In_521);
and U1227 (N_1227,In_815,In_387);
and U1228 (N_1228,In_500,In_175);
nor U1229 (N_1229,In_380,In_42);
nor U1230 (N_1230,In_564,In_96);
nor U1231 (N_1231,In_1004,In_540);
and U1232 (N_1232,In_1024,In_678);
nand U1233 (N_1233,In_22,In_566);
nand U1234 (N_1234,In_1476,In_79);
and U1235 (N_1235,In_1424,In_1060);
nor U1236 (N_1236,In_1433,In_476);
xor U1237 (N_1237,In_69,In_157);
nand U1238 (N_1238,In_1162,In_1030);
or U1239 (N_1239,In_432,In_1225);
or U1240 (N_1240,In_1471,In_73);
nor U1241 (N_1241,In_1495,In_112);
nor U1242 (N_1242,In_290,In_131);
nor U1243 (N_1243,In_947,In_941);
nor U1244 (N_1244,In_364,In_430);
and U1245 (N_1245,In_1221,In_734);
nor U1246 (N_1246,In_999,In_1246);
and U1247 (N_1247,In_414,In_629);
and U1248 (N_1248,In_1166,In_397);
or U1249 (N_1249,In_930,In_31);
or U1250 (N_1250,In_582,In_32);
and U1251 (N_1251,In_183,In_1244);
nor U1252 (N_1252,In_867,In_412);
or U1253 (N_1253,In_783,In_869);
nand U1254 (N_1254,In_473,In_1002);
or U1255 (N_1255,In_933,In_604);
or U1256 (N_1256,In_841,In_339);
nand U1257 (N_1257,In_0,In_55);
nor U1258 (N_1258,In_1331,In_1189);
and U1259 (N_1259,In_1270,In_1285);
nand U1260 (N_1260,In_1057,In_1274);
and U1261 (N_1261,In_705,In_1335);
nor U1262 (N_1262,In_509,In_1256);
nand U1263 (N_1263,In_1397,In_519);
nor U1264 (N_1264,In_1358,In_676);
nor U1265 (N_1265,In_52,In_1120);
nand U1266 (N_1266,In_79,In_1071);
nor U1267 (N_1267,In_995,In_576);
nor U1268 (N_1268,In_416,In_466);
or U1269 (N_1269,In_1461,In_107);
and U1270 (N_1270,In_105,In_264);
or U1271 (N_1271,In_88,In_1356);
or U1272 (N_1272,In_1471,In_208);
or U1273 (N_1273,In_1098,In_1393);
and U1274 (N_1274,In_770,In_822);
or U1275 (N_1275,In_1117,In_745);
and U1276 (N_1276,In_1261,In_652);
xor U1277 (N_1277,In_1445,In_184);
or U1278 (N_1278,In_11,In_136);
xnor U1279 (N_1279,In_929,In_1351);
and U1280 (N_1280,In_1072,In_87);
xnor U1281 (N_1281,In_1177,In_1490);
nand U1282 (N_1282,In_29,In_277);
nand U1283 (N_1283,In_631,In_472);
or U1284 (N_1284,In_1213,In_79);
xor U1285 (N_1285,In_646,In_72);
xnor U1286 (N_1286,In_93,In_692);
nand U1287 (N_1287,In_1319,In_1123);
nor U1288 (N_1288,In_1368,In_1283);
nor U1289 (N_1289,In_785,In_384);
or U1290 (N_1290,In_772,In_1492);
or U1291 (N_1291,In_550,In_723);
and U1292 (N_1292,In_113,In_1315);
nor U1293 (N_1293,In_464,In_687);
or U1294 (N_1294,In_490,In_641);
xnor U1295 (N_1295,In_132,In_616);
and U1296 (N_1296,In_1250,In_500);
nand U1297 (N_1297,In_489,In_1365);
and U1298 (N_1298,In_105,In_466);
nand U1299 (N_1299,In_315,In_384);
and U1300 (N_1300,In_392,In_215);
nor U1301 (N_1301,In_446,In_241);
and U1302 (N_1302,In_346,In_5);
nand U1303 (N_1303,In_973,In_587);
or U1304 (N_1304,In_1429,In_450);
nand U1305 (N_1305,In_1311,In_741);
or U1306 (N_1306,In_1395,In_43);
or U1307 (N_1307,In_422,In_380);
or U1308 (N_1308,In_80,In_512);
or U1309 (N_1309,In_661,In_1235);
nor U1310 (N_1310,In_728,In_24);
xor U1311 (N_1311,In_1242,In_1365);
nand U1312 (N_1312,In_1049,In_1388);
nor U1313 (N_1313,In_236,In_1441);
and U1314 (N_1314,In_95,In_1176);
or U1315 (N_1315,In_645,In_1294);
or U1316 (N_1316,In_697,In_45);
nand U1317 (N_1317,In_1032,In_255);
nor U1318 (N_1318,In_445,In_1359);
and U1319 (N_1319,In_1331,In_258);
nor U1320 (N_1320,In_836,In_1287);
nand U1321 (N_1321,In_1292,In_1452);
nor U1322 (N_1322,In_313,In_393);
nand U1323 (N_1323,In_180,In_1301);
or U1324 (N_1324,In_196,In_801);
nand U1325 (N_1325,In_1040,In_125);
nand U1326 (N_1326,In_134,In_1313);
or U1327 (N_1327,In_433,In_1085);
nor U1328 (N_1328,In_1081,In_277);
nor U1329 (N_1329,In_1322,In_6);
or U1330 (N_1330,In_655,In_1250);
nand U1331 (N_1331,In_43,In_657);
or U1332 (N_1332,In_41,In_760);
nor U1333 (N_1333,In_778,In_489);
nor U1334 (N_1334,In_1300,In_428);
xnor U1335 (N_1335,In_86,In_586);
or U1336 (N_1336,In_928,In_1170);
and U1337 (N_1337,In_483,In_1323);
nor U1338 (N_1338,In_752,In_1445);
or U1339 (N_1339,In_140,In_878);
and U1340 (N_1340,In_1061,In_114);
and U1341 (N_1341,In_485,In_1021);
xnor U1342 (N_1342,In_891,In_1474);
nand U1343 (N_1343,In_758,In_487);
nand U1344 (N_1344,In_1239,In_638);
nand U1345 (N_1345,In_657,In_428);
nand U1346 (N_1346,In_226,In_619);
nand U1347 (N_1347,In_383,In_302);
or U1348 (N_1348,In_1412,In_255);
nor U1349 (N_1349,In_1286,In_199);
nand U1350 (N_1350,In_458,In_455);
xnor U1351 (N_1351,In_666,In_394);
and U1352 (N_1352,In_358,In_835);
or U1353 (N_1353,In_508,In_661);
nand U1354 (N_1354,In_50,In_884);
nor U1355 (N_1355,In_470,In_1264);
nand U1356 (N_1356,In_546,In_1264);
nand U1357 (N_1357,In_1131,In_248);
and U1358 (N_1358,In_1492,In_693);
nand U1359 (N_1359,In_273,In_1208);
nand U1360 (N_1360,In_289,In_35);
and U1361 (N_1361,In_950,In_642);
or U1362 (N_1362,In_1063,In_92);
nand U1363 (N_1363,In_1181,In_779);
nand U1364 (N_1364,In_1230,In_1365);
nand U1365 (N_1365,In_1385,In_619);
xor U1366 (N_1366,In_351,In_646);
nand U1367 (N_1367,In_633,In_1085);
or U1368 (N_1368,In_204,In_1342);
or U1369 (N_1369,In_202,In_1238);
nor U1370 (N_1370,In_1172,In_639);
or U1371 (N_1371,In_876,In_1388);
nand U1372 (N_1372,In_329,In_92);
nor U1373 (N_1373,In_411,In_1414);
nor U1374 (N_1374,In_252,In_616);
xor U1375 (N_1375,In_621,In_363);
or U1376 (N_1376,In_226,In_729);
and U1377 (N_1377,In_211,In_545);
and U1378 (N_1378,In_44,In_1138);
or U1379 (N_1379,In_672,In_838);
or U1380 (N_1380,In_108,In_1410);
and U1381 (N_1381,In_484,In_1277);
nand U1382 (N_1382,In_494,In_110);
nor U1383 (N_1383,In_520,In_1164);
and U1384 (N_1384,In_1278,In_514);
nor U1385 (N_1385,In_463,In_394);
nand U1386 (N_1386,In_798,In_1068);
and U1387 (N_1387,In_251,In_857);
xor U1388 (N_1388,In_1065,In_1232);
nor U1389 (N_1389,In_1069,In_1409);
nor U1390 (N_1390,In_241,In_974);
or U1391 (N_1391,In_909,In_280);
nor U1392 (N_1392,In_813,In_960);
nand U1393 (N_1393,In_835,In_983);
nand U1394 (N_1394,In_195,In_828);
nand U1395 (N_1395,In_1372,In_1134);
xnor U1396 (N_1396,In_1044,In_458);
or U1397 (N_1397,In_582,In_856);
or U1398 (N_1398,In_1464,In_1133);
nor U1399 (N_1399,In_109,In_652);
or U1400 (N_1400,In_1479,In_41);
and U1401 (N_1401,In_750,In_441);
nor U1402 (N_1402,In_507,In_1355);
and U1403 (N_1403,In_1449,In_649);
or U1404 (N_1404,In_1158,In_1205);
and U1405 (N_1405,In_1293,In_829);
nor U1406 (N_1406,In_567,In_1175);
nor U1407 (N_1407,In_149,In_212);
nor U1408 (N_1408,In_1063,In_458);
xnor U1409 (N_1409,In_150,In_953);
nor U1410 (N_1410,In_1480,In_424);
or U1411 (N_1411,In_909,In_1453);
or U1412 (N_1412,In_1355,In_495);
nor U1413 (N_1413,In_787,In_1077);
xor U1414 (N_1414,In_911,In_1015);
nor U1415 (N_1415,In_1468,In_242);
nor U1416 (N_1416,In_639,In_1328);
nand U1417 (N_1417,In_1180,In_980);
xnor U1418 (N_1418,In_1205,In_774);
and U1419 (N_1419,In_310,In_406);
xnor U1420 (N_1420,In_44,In_219);
and U1421 (N_1421,In_185,In_1345);
nand U1422 (N_1422,In_1009,In_631);
xor U1423 (N_1423,In_1074,In_174);
or U1424 (N_1424,In_1437,In_1);
or U1425 (N_1425,In_678,In_1183);
nand U1426 (N_1426,In_1248,In_1165);
and U1427 (N_1427,In_762,In_669);
nand U1428 (N_1428,In_1405,In_3);
nand U1429 (N_1429,In_684,In_174);
or U1430 (N_1430,In_122,In_1199);
nand U1431 (N_1431,In_83,In_1415);
nand U1432 (N_1432,In_1001,In_77);
and U1433 (N_1433,In_334,In_175);
nand U1434 (N_1434,In_788,In_1445);
and U1435 (N_1435,In_1305,In_167);
or U1436 (N_1436,In_975,In_92);
or U1437 (N_1437,In_1452,In_518);
nand U1438 (N_1438,In_1392,In_1418);
nand U1439 (N_1439,In_660,In_838);
and U1440 (N_1440,In_679,In_810);
and U1441 (N_1441,In_1266,In_552);
and U1442 (N_1442,In_363,In_924);
nor U1443 (N_1443,In_422,In_888);
nor U1444 (N_1444,In_588,In_1300);
nand U1445 (N_1445,In_902,In_746);
xnor U1446 (N_1446,In_501,In_612);
and U1447 (N_1447,In_361,In_16);
xor U1448 (N_1448,In_1064,In_1289);
nor U1449 (N_1449,In_1228,In_1234);
or U1450 (N_1450,In_1351,In_68);
nand U1451 (N_1451,In_480,In_1018);
and U1452 (N_1452,In_1197,In_1450);
or U1453 (N_1453,In_203,In_1477);
nor U1454 (N_1454,In_230,In_1214);
nand U1455 (N_1455,In_433,In_1117);
xnor U1456 (N_1456,In_301,In_315);
xor U1457 (N_1457,In_758,In_418);
nand U1458 (N_1458,In_1472,In_986);
and U1459 (N_1459,In_1370,In_1312);
xor U1460 (N_1460,In_252,In_725);
nor U1461 (N_1461,In_1287,In_1202);
xor U1462 (N_1462,In_525,In_436);
and U1463 (N_1463,In_335,In_384);
nor U1464 (N_1464,In_658,In_999);
xor U1465 (N_1465,In_609,In_1237);
nand U1466 (N_1466,In_1202,In_1227);
xnor U1467 (N_1467,In_1397,In_1433);
nand U1468 (N_1468,In_1421,In_1262);
and U1469 (N_1469,In_23,In_607);
nor U1470 (N_1470,In_1016,In_1293);
nand U1471 (N_1471,In_346,In_242);
xor U1472 (N_1472,In_1443,In_686);
nand U1473 (N_1473,In_863,In_50);
xor U1474 (N_1474,In_1340,In_959);
or U1475 (N_1475,In_161,In_498);
and U1476 (N_1476,In_1404,In_1478);
and U1477 (N_1477,In_1181,In_1266);
nor U1478 (N_1478,In_1171,In_643);
nand U1479 (N_1479,In_424,In_740);
nand U1480 (N_1480,In_82,In_498);
or U1481 (N_1481,In_675,In_605);
nand U1482 (N_1482,In_461,In_129);
nor U1483 (N_1483,In_276,In_699);
nand U1484 (N_1484,In_374,In_212);
and U1485 (N_1485,In_818,In_5);
nor U1486 (N_1486,In_886,In_1349);
or U1487 (N_1487,In_519,In_1216);
or U1488 (N_1488,In_836,In_1476);
nand U1489 (N_1489,In_310,In_989);
nand U1490 (N_1490,In_262,In_1243);
nor U1491 (N_1491,In_590,In_275);
nor U1492 (N_1492,In_87,In_1382);
and U1493 (N_1493,In_1214,In_246);
nor U1494 (N_1494,In_390,In_772);
and U1495 (N_1495,In_324,In_496);
or U1496 (N_1496,In_833,In_951);
nand U1497 (N_1497,In_1063,In_1135);
nor U1498 (N_1498,In_437,In_1333);
nand U1499 (N_1499,In_582,In_903);
nor U1500 (N_1500,In_77,In_48);
and U1501 (N_1501,In_297,In_351);
and U1502 (N_1502,In_1298,In_48);
xor U1503 (N_1503,In_1202,In_1354);
and U1504 (N_1504,In_95,In_638);
and U1505 (N_1505,In_44,In_1021);
and U1506 (N_1506,In_91,In_427);
and U1507 (N_1507,In_646,In_47);
and U1508 (N_1508,In_1039,In_218);
nor U1509 (N_1509,In_101,In_1265);
nor U1510 (N_1510,In_19,In_983);
nor U1511 (N_1511,In_698,In_1294);
and U1512 (N_1512,In_1433,In_1230);
and U1513 (N_1513,In_131,In_454);
nor U1514 (N_1514,In_942,In_1039);
nor U1515 (N_1515,In_61,In_435);
nand U1516 (N_1516,In_553,In_426);
or U1517 (N_1517,In_187,In_1121);
xor U1518 (N_1518,In_20,In_1346);
nand U1519 (N_1519,In_453,In_1452);
and U1520 (N_1520,In_496,In_862);
nand U1521 (N_1521,In_645,In_1415);
nand U1522 (N_1522,In_338,In_798);
or U1523 (N_1523,In_705,In_26);
xor U1524 (N_1524,In_12,In_570);
nand U1525 (N_1525,In_640,In_602);
or U1526 (N_1526,In_1097,In_296);
nand U1527 (N_1527,In_841,In_953);
and U1528 (N_1528,In_872,In_188);
nand U1529 (N_1529,In_861,In_1279);
nand U1530 (N_1530,In_630,In_102);
or U1531 (N_1531,In_1052,In_242);
and U1532 (N_1532,In_190,In_104);
nor U1533 (N_1533,In_1217,In_115);
nor U1534 (N_1534,In_1158,In_1296);
and U1535 (N_1535,In_508,In_649);
and U1536 (N_1536,In_1492,In_155);
and U1537 (N_1537,In_87,In_738);
nand U1538 (N_1538,In_1074,In_382);
nand U1539 (N_1539,In_646,In_1396);
nand U1540 (N_1540,In_959,In_1311);
nor U1541 (N_1541,In_894,In_1193);
or U1542 (N_1542,In_426,In_399);
and U1543 (N_1543,In_1474,In_1315);
and U1544 (N_1544,In_921,In_1416);
or U1545 (N_1545,In_192,In_1111);
or U1546 (N_1546,In_1012,In_355);
nand U1547 (N_1547,In_864,In_267);
or U1548 (N_1548,In_102,In_638);
xor U1549 (N_1549,In_656,In_38);
nand U1550 (N_1550,In_1447,In_1323);
nor U1551 (N_1551,In_1409,In_605);
and U1552 (N_1552,In_281,In_1239);
xor U1553 (N_1553,In_1051,In_518);
or U1554 (N_1554,In_1438,In_681);
nand U1555 (N_1555,In_706,In_445);
and U1556 (N_1556,In_529,In_1052);
nor U1557 (N_1557,In_699,In_712);
or U1558 (N_1558,In_834,In_842);
xnor U1559 (N_1559,In_141,In_653);
nor U1560 (N_1560,In_202,In_617);
and U1561 (N_1561,In_457,In_644);
or U1562 (N_1562,In_19,In_347);
or U1563 (N_1563,In_1355,In_854);
and U1564 (N_1564,In_1195,In_729);
or U1565 (N_1565,In_922,In_90);
or U1566 (N_1566,In_1489,In_1448);
xnor U1567 (N_1567,In_561,In_557);
nor U1568 (N_1568,In_780,In_472);
and U1569 (N_1569,In_1319,In_602);
nor U1570 (N_1570,In_167,In_548);
nand U1571 (N_1571,In_25,In_1290);
or U1572 (N_1572,In_765,In_1208);
and U1573 (N_1573,In_930,In_525);
nand U1574 (N_1574,In_1007,In_1401);
nor U1575 (N_1575,In_1224,In_1232);
nor U1576 (N_1576,In_694,In_230);
nor U1577 (N_1577,In_1349,In_1271);
nor U1578 (N_1578,In_660,In_461);
and U1579 (N_1579,In_399,In_1091);
nor U1580 (N_1580,In_1014,In_903);
nand U1581 (N_1581,In_1215,In_413);
or U1582 (N_1582,In_109,In_972);
nand U1583 (N_1583,In_355,In_1471);
nor U1584 (N_1584,In_1144,In_368);
nand U1585 (N_1585,In_160,In_885);
and U1586 (N_1586,In_843,In_709);
or U1587 (N_1587,In_869,In_1284);
nor U1588 (N_1588,In_207,In_372);
nand U1589 (N_1589,In_40,In_1093);
or U1590 (N_1590,In_588,In_855);
or U1591 (N_1591,In_419,In_995);
and U1592 (N_1592,In_256,In_527);
nand U1593 (N_1593,In_978,In_491);
nor U1594 (N_1594,In_911,In_178);
xnor U1595 (N_1595,In_1401,In_330);
nand U1596 (N_1596,In_1389,In_780);
nor U1597 (N_1597,In_269,In_1009);
and U1598 (N_1598,In_830,In_1360);
or U1599 (N_1599,In_261,In_606);
nand U1600 (N_1600,In_1056,In_1221);
and U1601 (N_1601,In_291,In_478);
nand U1602 (N_1602,In_542,In_1011);
nor U1603 (N_1603,In_1443,In_521);
nand U1604 (N_1604,In_299,In_536);
xor U1605 (N_1605,In_418,In_71);
or U1606 (N_1606,In_1221,In_915);
and U1607 (N_1607,In_935,In_469);
or U1608 (N_1608,In_1044,In_864);
nor U1609 (N_1609,In_1169,In_676);
nand U1610 (N_1610,In_1309,In_1422);
nand U1611 (N_1611,In_945,In_894);
nand U1612 (N_1612,In_533,In_1105);
nand U1613 (N_1613,In_451,In_575);
xor U1614 (N_1614,In_1489,In_879);
and U1615 (N_1615,In_647,In_248);
nand U1616 (N_1616,In_1412,In_1494);
and U1617 (N_1617,In_902,In_56);
nor U1618 (N_1618,In_228,In_39);
and U1619 (N_1619,In_1498,In_731);
xor U1620 (N_1620,In_904,In_697);
nand U1621 (N_1621,In_469,In_720);
and U1622 (N_1622,In_541,In_308);
nor U1623 (N_1623,In_451,In_1153);
nor U1624 (N_1624,In_77,In_1347);
nor U1625 (N_1625,In_865,In_1488);
nor U1626 (N_1626,In_295,In_201);
nand U1627 (N_1627,In_434,In_604);
nand U1628 (N_1628,In_337,In_296);
nand U1629 (N_1629,In_1454,In_240);
nor U1630 (N_1630,In_248,In_40);
or U1631 (N_1631,In_725,In_832);
nor U1632 (N_1632,In_767,In_1080);
nor U1633 (N_1633,In_1369,In_955);
nor U1634 (N_1634,In_41,In_426);
or U1635 (N_1635,In_577,In_1269);
and U1636 (N_1636,In_1235,In_1483);
nor U1637 (N_1637,In_165,In_706);
nand U1638 (N_1638,In_1025,In_614);
or U1639 (N_1639,In_265,In_1210);
and U1640 (N_1640,In_742,In_802);
or U1641 (N_1641,In_1485,In_971);
nor U1642 (N_1642,In_616,In_570);
nor U1643 (N_1643,In_1118,In_642);
nand U1644 (N_1644,In_1210,In_920);
xor U1645 (N_1645,In_728,In_1428);
nor U1646 (N_1646,In_671,In_900);
or U1647 (N_1647,In_531,In_187);
or U1648 (N_1648,In_584,In_789);
nand U1649 (N_1649,In_42,In_687);
nand U1650 (N_1650,In_700,In_1456);
or U1651 (N_1651,In_1443,In_359);
xor U1652 (N_1652,In_969,In_511);
nor U1653 (N_1653,In_569,In_1219);
and U1654 (N_1654,In_992,In_305);
or U1655 (N_1655,In_1015,In_1190);
xor U1656 (N_1656,In_1132,In_1321);
or U1657 (N_1657,In_77,In_972);
and U1658 (N_1658,In_942,In_440);
nand U1659 (N_1659,In_1136,In_872);
nand U1660 (N_1660,In_1261,In_1414);
or U1661 (N_1661,In_1315,In_1485);
and U1662 (N_1662,In_907,In_313);
or U1663 (N_1663,In_100,In_1324);
and U1664 (N_1664,In_1042,In_1067);
or U1665 (N_1665,In_386,In_44);
nor U1666 (N_1666,In_872,In_1199);
or U1667 (N_1667,In_820,In_1237);
or U1668 (N_1668,In_599,In_143);
and U1669 (N_1669,In_1189,In_664);
nand U1670 (N_1670,In_1332,In_72);
nor U1671 (N_1671,In_54,In_855);
and U1672 (N_1672,In_1429,In_153);
or U1673 (N_1673,In_493,In_1380);
nand U1674 (N_1674,In_331,In_377);
nor U1675 (N_1675,In_1027,In_730);
nor U1676 (N_1676,In_1472,In_505);
and U1677 (N_1677,In_3,In_1119);
nor U1678 (N_1678,In_1128,In_143);
and U1679 (N_1679,In_169,In_891);
or U1680 (N_1680,In_1457,In_1460);
nand U1681 (N_1681,In_1174,In_1440);
and U1682 (N_1682,In_957,In_810);
and U1683 (N_1683,In_535,In_67);
nand U1684 (N_1684,In_1101,In_855);
xor U1685 (N_1685,In_1171,In_55);
nor U1686 (N_1686,In_77,In_1100);
and U1687 (N_1687,In_1240,In_415);
nor U1688 (N_1688,In_1157,In_363);
or U1689 (N_1689,In_313,In_1117);
and U1690 (N_1690,In_822,In_848);
and U1691 (N_1691,In_1378,In_1428);
and U1692 (N_1692,In_1450,In_718);
nand U1693 (N_1693,In_1158,In_724);
or U1694 (N_1694,In_150,In_1130);
nor U1695 (N_1695,In_70,In_768);
nand U1696 (N_1696,In_1153,In_856);
and U1697 (N_1697,In_605,In_773);
and U1698 (N_1698,In_402,In_824);
xnor U1699 (N_1699,In_434,In_667);
and U1700 (N_1700,In_584,In_504);
xnor U1701 (N_1701,In_55,In_863);
or U1702 (N_1702,In_942,In_563);
nor U1703 (N_1703,In_391,In_838);
xor U1704 (N_1704,In_839,In_12);
and U1705 (N_1705,In_1450,In_1428);
and U1706 (N_1706,In_1369,In_55);
or U1707 (N_1707,In_822,In_1420);
or U1708 (N_1708,In_1088,In_344);
nand U1709 (N_1709,In_1265,In_1124);
nor U1710 (N_1710,In_765,In_1479);
xor U1711 (N_1711,In_297,In_1275);
and U1712 (N_1712,In_17,In_867);
and U1713 (N_1713,In_1050,In_654);
nor U1714 (N_1714,In_1078,In_738);
nor U1715 (N_1715,In_837,In_966);
or U1716 (N_1716,In_939,In_623);
nand U1717 (N_1717,In_18,In_181);
or U1718 (N_1718,In_777,In_702);
xnor U1719 (N_1719,In_1251,In_819);
and U1720 (N_1720,In_277,In_824);
nor U1721 (N_1721,In_1490,In_147);
nor U1722 (N_1722,In_1038,In_203);
nor U1723 (N_1723,In_1195,In_1136);
nor U1724 (N_1724,In_782,In_1304);
xnor U1725 (N_1725,In_1020,In_1072);
and U1726 (N_1726,In_900,In_850);
xor U1727 (N_1727,In_554,In_1415);
nand U1728 (N_1728,In_792,In_1356);
and U1729 (N_1729,In_1387,In_396);
nor U1730 (N_1730,In_1122,In_339);
or U1731 (N_1731,In_648,In_783);
nor U1732 (N_1732,In_1395,In_1373);
and U1733 (N_1733,In_774,In_100);
nor U1734 (N_1734,In_1375,In_814);
nand U1735 (N_1735,In_1159,In_677);
nand U1736 (N_1736,In_1049,In_1498);
or U1737 (N_1737,In_1259,In_1240);
nor U1738 (N_1738,In_764,In_598);
nor U1739 (N_1739,In_155,In_1476);
nor U1740 (N_1740,In_838,In_802);
or U1741 (N_1741,In_689,In_1160);
nand U1742 (N_1742,In_384,In_558);
and U1743 (N_1743,In_157,In_1406);
nor U1744 (N_1744,In_481,In_1124);
xor U1745 (N_1745,In_651,In_1431);
xnor U1746 (N_1746,In_1215,In_553);
nor U1747 (N_1747,In_1110,In_1115);
or U1748 (N_1748,In_1099,In_127);
nor U1749 (N_1749,In_1343,In_1163);
nand U1750 (N_1750,In_296,In_290);
xor U1751 (N_1751,In_124,In_123);
nor U1752 (N_1752,In_284,In_61);
nor U1753 (N_1753,In_1321,In_1142);
and U1754 (N_1754,In_1138,In_863);
nand U1755 (N_1755,In_282,In_453);
nand U1756 (N_1756,In_607,In_441);
and U1757 (N_1757,In_318,In_1210);
nand U1758 (N_1758,In_1049,In_794);
xor U1759 (N_1759,In_1420,In_1376);
nor U1760 (N_1760,In_810,In_1044);
nor U1761 (N_1761,In_1163,In_1195);
and U1762 (N_1762,In_411,In_1018);
or U1763 (N_1763,In_613,In_1131);
nor U1764 (N_1764,In_487,In_83);
nand U1765 (N_1765,In_643,In_975);
xnor U1766 (N_1766,In_1493,In_1336);
nor U1767 (N_1767,In_1496,In_46);
or U1768 (N_1768,In_1474,In_712);
or U1769 (N_1769,In_921,In_264);
or U1770 (N_1770,In_41,In_1418);
or U1771 (N_1771,In_704,In_766);
nand U1772 (N_1772,In_62,In_66);
nor U1773 (N_1773,In_1423,In_1434);
xor U1774 (N_1774,In_1290,In_914);
and U1775 (N_1775,In_58,In_1425);
nor U1776 (N_1776,In_166,In_50);
or U1777 (N_1777,In_269,In_1090);
nand U1778 (N_1778,In_1400,In_375);
nand U1779 (N_1779,In_703,In_1179);
and U1780 (N_1780,In_1295,In_1410);
and U1781 (N_1781,In_246,In_906);
nor U1782 (N_1782,In_27,In_731);
nor U1783 (N_1783,In_1479,In_1303);
and U1784 (N_1784,In_1431,In_691);
or U1785 (N_1785,In_1309,In_256);
or U1786 (N_1786,In_939,In_483);
nor U1787 (N_1787,In_923,In_367);
nor U1788 (N_1788,In_462,In_1466);
and U1789 (N_1789,In_292,In_925);
and U1790 (N_1790,In_236,In_738);
and U1791 (N_1791,In_928,In_1029);
nor U1792 (N_1792,In_282,In_1342);
nor U1793 (N_1793,In_206,In_1307);
and U1794 (N_1794,In_157,In_1412);
nor U1795 (N_1795,In_1265,In_314);
or U1796 (N_1796,In_600,In_1278);
or U1797 (N_1797,In_1116,In_875);
and U1798 (N_1798,In_96,In_1076);
nor U1799 (N_1799,In_1015,In_350);
nor U1800 (N_1800,In_319,In_631);
nor U1801 (N_1801,In_1298,In_187);
nand U1802 (N_1802,In_855,In_1402);
nor U1803 (N_1803,In_347,In_247);
and U1804 (N_1804,In_1444,In_762);
or U1805 (N_1805,In_229,In_321);
nor U1806 (N_1806,In_628,In_1315);
and U1807 (N_1807,In_395,In_661);
nor U1808 (N_1808,In_1480,In_408);
nor U1809 (N_1809,In_1388,In_1034);
or U1810 (N_1810,In_95,In_672);
or U1811 (N_1811,In_571,In_222);
or U1812 (N_1812,In_34,In_1324);
xnor U1813 (N_1813,In_75,In_997);
and U1814 (N_1814,In_1066,In_402);
or U1815 (N_1815,In_859,In_891);
nand U1816 (N_1816,In_846,In_30);
nand U1817 (N_1817,In_94,In_44);
nor U1818 (N_1818,In_1031,In_990);
and U1819 (N_1819,In_1352,In_1016);
nor U1820 (N_1820,In_201,In_29);
and U1821 (N_1821,In_549,In_435);
or U1822 (N_1822,In_1427,In_829);
nand U1823 (N_1823,In_815,In_1281);
and U1824 (N_1824,In_13,In_1006);
nor U1825 (N_1825,In_528,In_412);
and U1826 (N_1826,In_862,In_456);
and U1827 (N_1827,In_1425,In_68);
nand U1828 (N_1828,In_904,In_155);
xnor U1829 (N_1829,In_697,In_893);
and U1830 (N_1830,In_193,In_1067);
and U1831 (N_1831,In_50,In_554);
nand U1832 (N_1832,In_481,In_100);
nand U1833 (N_1833,In_314,In_1034);
xor U1834 (N_1834,In_1047,In_1450);
nand U1835 (N_1835,In_741,In_952);
and U1836 (N_1836,In_6,In_1381);
nand U1837 (N_1837,In_63,In_436);
nand U1838 (N_1838,In_275,In_259);
nor U1839 (N_1839,In_443,In_93);
nand U1840 (N_1840,In_485,In_17);
nand U1841 (N_1841,In_353,In_554);
nor U1842 (N_1842,In_712,In_171);
or U1843 (N_1843,In_1238,In_538);
nand U1844 (N_1844,In_483,In_508);
xnor U1845 (N_1845,In_697,In_661);
xor U1846 (N_1846,In_1433,In_888);
xnor U1847 (N_1847,In_488,In_570);
nor U1848 (N_1848,In_1428,In_653);
nor U1849 (N_1849,In_1242,In_1126);
nand U1850 (N_1850,In_744,In_1150);
nand U1851 (N_1851,In_959,In_868);
and U1852 (N_1852,In_90,In_857);
or U1853 (N_1853,In_237,In_306);
nand U1854 (N_1854,In_810,In_358);
nor U1855 (N_1855,In_926,In_1342);
nor U1856 (N_1856,In_616,In_952);
xnor U1857 (N_1857,In_593,In_568);
xor U1858 (N_1858,In_140,In_501);
or U1859 (N_1859,In_17,In_1291);
nor U1860 (N_1860,In_162,In_1418);
and U1861 (N_1861,In_46,In_1365);
nor U1862 (N_1862,In_658,In_1283);
or U1863 (N_1863,In_259,In_942);
nand U1864 (N_1864,In_205,In_788);
nor U1865 (N_1865,In_355,In_1028);
or U1866 (N_1866,In_434,In_967);
and U1867 (N_1867,In_799,In_961);
nand U1868 (N_1868,In_167,In_851);
nand U1869 (N_1869,In_995,In_1207);
and U1870 (N_1870,In_879,In_1456);
xnor U1871 (N_1871,In_1065,In_1355);
nor U1872 (N_1872,In_502,In_552);
or U1873 (N_1873,In_39,In_1273);
nand U1874 (N_1874,In_367,In_671);
xor U1875 (N_1875,In_774,In_1315);
nand U1876 (N_1876,In_613,In_387);
or U1877 (N_1877,In_193,In_1438);
nor U1878 (N_1878,In_171,In_77);
and U1879 (N_1879,In_780,In_406);
or U1880 (N_1880,In_574,In_1055);
xnor U1881 (N_1881,In_332,In_723);
nand U1882 (N_1882,In_190,In_1414);
and U1883 (N_1883,In_1160,In_877);
and U1884 (N_1884,In_938,In_486);
and U1885 (N_1885,In_203,In_216);
nand U1886 (N_1886,In_1311,In_1405);
and U1887 (N_1887,In_1162,In_437);
or U1888 (N_1888,In_383,In_1324);
and U1889 (N_1889,In_980,In_1198);
nor U1890 (N_1890,In_1030,In_169);
nor U1891 (N_1891,In_283,In_561);
or U1892 (N_1892,In_287,In_445);
xor U1893 (N_1893,In_796,In_1424);
and U1894 (N_1894,In_925,In_459);
or U1895 (N_1895,In_647,In_1040);
nor U1896 (N_1896,In_909,In_627);
or U1897 (N_1897,In_1496,In_766);
nand U1898 (N_1898,In_64,In_16);
or U1899 (N_1899,In_528,In_1247);
and U1900 (N_1900,In_834,In_343);
nand U1901 (N_1901,In_1002,In_19);
and U1902 (N_1902,In_1227,In_313);
nor U1903 (N_1903,In_133,In_968);
or U1904 (N_1904,In_1044,In_573);
and U1905 (N_1905,In_255,In_817);
nor U1906 (N_1906,In_172,In_1367);
and U1907 (N_1907,In_1164,In_583);
nor U1908 (N_1908,In_1468,In_520);
or U1909 (N_1909,In_1349,In_1361);
and U1910 (N_1910,In_197,In_924);
nand U1911 (N_1911,In_869,In_1220);
nor U1912 (N_1912,In_1061,In_226);
or U1913 (N_1913,In_1212,In_1331);
nor U1914 (N_1914,In_1447,In_538);
or U1915 (N_1915,In_816,In_818);
nor U1916 (N_1916,In_133,In_926);
xor U1917 (N_1917,In_173,In_593);
or U1918 (N_1918,In_957,In_913);
nand U1919 (N_1919,In_1320,In_1129);
nor U1920 (N_1920,In_1256,In_1347);
nand U1921 (N_1921,In_937,In_864);
and U1922 (N_1922,In_669,In_92);
or U1923 (N_1923,In_563,In_511);
or U1924 (N_1924,In_225,In_400);
nor U1925 (N_1925,In_670,In_1399);
nand U1926 (N_1926,In_850,In_27);
xor U1927 (N_1927,In_407,In_980);
and U1928 (N_1928,In_1115,In_259);
and U1929 (N_1929,In_761,In_378);
nor U1930 (N_1930,In_1104,In_159);
or U1931 (N_1931,In_1084,In_803);
and U1932 (N_1932,In_1025,In_114);
or U1933 (N_1933,In_681,In_529);
nand U1934 (N_1934,In_375,In_129);
or U1935 (N_1935,In_1385,In_697);
nor U1936 (N_1936,In_1143,In_929);
or U1937 (N_1937,In_121,In_1324);
xnor U1938 (N_1938,In_658,In_1337);
nand U1939 (N_1939,In_958,In_1412);
or U1940 (N_1940,In_1109,In_619);
nand U1941 (N_1941,In_380,In_413);
or U1942 (N_1942,In_321,In_1454);
or U1943 (N_1943,In_1478,In_992);
or U1944 (N_1944,In_1400,In_1309);
nor U1945 (N_1945,In_980,In_497);
nand U1946 (N_1946,In_1346,In_939);
and U1947 (N_1947,In_1266,In_0);
and U1948 (N_1948,In_835,In_854);
nor U1949 (N_1949,In_340,In_37);
nor U1950 (N_1950,In_150,In_743);
or U1951 (N_1951,In_1328,In_682);
or U1952 (N_1952,In_1408,In_289);
xnor U1953 (N_1953,In_670,In_654);
and U1954 (N_1954,In_317,In_255);
nor U1955 (N_1955,In_198,In_1497);
or U1956 (N_1956,In_635,In_610);
or U1957 (N_1957,In_22,In_292);
or U1958 (N_1958,In_319,In_216);
nor U1959 (N_1959,In_276,In_1361);
or U1960 (N_1960,In_399,In_728);
nor U1961 (N_1961,In_662,In_763);
xnor U1962 (N_1962,In_1064,In_87);
nand U1963 (N_1963,In_476,In_950);
or U1964 (N_1964,In_1136,In_1186);
nor U1965 (N_1965,In_1277,In_935);
nand U1966 (N_1966,In_486,In_1101);
nor U1967 (N_1967,In_324,In_279);
and U1968 (N_1968,In_132,In_453);
or U1969 (N_1969,In_1161,In_1190);
xor U1970 (N_1970,In_1396,In_1194);
or U1971 (N_1971,In_416,In_1490);
nand U1972 (N_1972,In_187,In_916);
and U1973 (N_1973,In_1400,In_1023);
nand U1974 (N_1974,In_955,In_479);
or U1975 (N_1975,In_592,In_93);
and U1976 (N_1976,In_230,In_724);
nor U1977 (N_1977,In_1105,In_970);
nand U1978 (N_1978,In_1052,In_1240);
and U1979 (N_1979,In_1362,In_519);
nor U1980 (N_1980,In_512,In_1090);
nand U1981 (N_1981,In_1425,In_1352);
nor U1982 (N_1982,In_1029,In_158);
or U1983 (N_1983,In_275,In_1021);
nor U1984 (N_1984,In_230,In_1427);
nor U1985 (N_1985,In_1315,In_897);
nor U1986 (N_1986,In_373,In_781);
nand U1987 (N_1987,In_1085,In_728);
nand U1988 (N_1988,In_1107,In_382);
or U1989 (N_1989,In_306,In_1084);
nor U1990 (N_1990,In_1488,In_572);
or U1991 (N_1991,In_446,In_350);
nand U1992 (N_1992,In_146,In_1242);
xor U1993 (N_1993,In_1454,In_1408);
nand U1994 (N_1994,In_49,In_518);
or U1995 (N_1995,In_450,In_1257);
or U1996 (N_1996,In_833,In_191);
or U1997 (N_1997,In_1473,In_635);
nand U1998 (N_1998,In_1107,In_1212);
and U1999 (N_1999,In_934,In_634);
or U2000 (N_2000,In_118,In_728);
and U2001 (N_2001,In_629,In_380);
nor U2002 (N_2002,In_828,In_603);
or U2003 (N_2003,In_695,In_1478);
nor U2004 (N_2004,In_378,In_663);
or U2005 (N_2005,In_1489,In_1485);
nand U2006 (N_2006,In_1044,In_720);
nor U2007 (N_2007,In_956,In_1223);
nand U2008 (N_2008,In_406,In_1230);
xnor U2009 (N_2009,In_499,In_1236);
nor U2010 (N_2010,In_107,In_992);
and U2011 (N_2011,In_1054,In_1181);
or U2012 (N_2012,In_1384,In_282);
and U2013 (N_2013,In_662,In_674);
nand U2014 (N_2014,In_735,In_569);
nor U2015 (N_2015,In_1142,In_152);
nor U2016 (N_2016,In_1305,In_921);
xor U2017 (N_2017,In_976,In_547);
nor U2018 (N_2018,In_6,In_469);
xnor U2019 (N_2019,In_530,In_1299);
nor U2020 (N_2020,In_252,In_1035);
and U2021 (N_2021,In_591,In_1164);
xor U2022 (N_2022,In_195,In_1091);
nor U2023 (N_2023,In_1339,In_884);
or U2024 (N_2024,In_556,In_1389);
or U2025 (N_2025,In_1433,In_538);
and U2026 (N_2026,In_496,In_1376);
nor U2027 (N_2027,In_1470,In_103);
and U2028 (N_2028,In_186,In_304);
and U2029 (N_2029,In_1420,In_1048);
nor U2030 (N_2030,In_445,In_524);
nand U2031 (N_2031,In_1302,In_1064);
nor U2032 (N_2032,In_347,In_1404);
nand U2033 (N_2033,In_281,In_89);
and U2034 (N_2034,In_48,In_90);
or U2035 (N_2035,In_1347,In_1198);
and U2036 (N_2036,In_863,In_1387);
and U2037 (N_2037,In_969,In_2);
and U2038 (N_2038,In_451,In_613);
and U2039 (N_2039,In_284,In_683);
nor U2040 (N_2040,In_1116,In_1067);
nor U2041 (N_2041,In_19,In_1089);
and U2042 (N_2042,In_46,In_796);
nor U2043 (N_2043,In_96,In_725);
and U2044 (N_2044,In_363,In_1237);
nand U2045 (N_2045,In_1096,In_371);
or U2046 (N_2046,In_669,In_1394);
nor U2047 (N_2047,In_874,In_336);
nand U2048 (N_2048,In_266,In_477);
and U2049 (N_2049,In_188,In_573);
nor U2050 (N_2050,In_671,In_926);
or U2051 (N_2051,In_327,In_459);
or U2052 (N_2052,In_744,In_812);
or U2053 (N_2053,In_54,In_387);
or U2054 (N_2054,In_1073,In_271);
or U2055 (N_2055,In_303,In_1133);
xor U2056 (N_2056,In_374,In_1198);
nor U2057 (N_2057,In_1084,In_995);
nor U2058 (N_2058,In_947,In_618);
nor U2059 (N_2059,In_1297,In_660);
and U2060 (N_2060,In_1042,In_535);
nor U2061 (N_2061,In_1155,In_19);
and U2062 (N_2062,In_744,In_1319);
or U2063 (N_2063,In_822,In_178);
and U2064 (N_2064,In_70,In_557);
nand U2065 (N_2065,In_1171,In_1338);
nor U2066 (N_2066,In_636,In_277);
nor U2067 (N_2067,In_961,In_6);
nand U2068 (N_2068,In_910,In_320);
nand U2069 (N_2069,In_1113,In_369);
nor U2070 (N_2070,In_574,In_345);
nor U2071 (N_2071,In_76,In_517);
and U2072 (N_2072,In_573,In_862);
nand U2073 (N_2073,In_730,In_444);
nor U2074 (N_2074,In_776,In_1161);
and U2075 (N_2075,In_1245,In_1411);
nor U2076 (N_2076,In_274,In_463);
and U2077 (N_2077,In_128,In_604);
xnor U2078 (N_2078,In_375,In_584);
nor U2079 (N_2079,In_873,In_139);
and U2080 (N_2080,In_1154,In_4);
nand U2081 (N_2081,In_468,In_1364);
nor U2082 (N_2082,In_590,In_372);
nand U2083 (N_2083,In_53,In_1127);
nand U2084 (N_2084,In_224,In_1012);
or U2085 (N_2085,In_1042,In_709);
nor U2086 (N_2086,In_1398,In_29);
nor U2087 (N_2087,In_187,In_854);
xnor U2088 (N_2088,In_94,In_261);
nor U2089 (N_2089,In_991,In_893);
nand U2090 (N_2090,In_99,In_1449);
and U2091 (N_2091,In_1473,In_1492);
nand U2092 (N_2092,In_92,In_764);
nand U2093 (N_2093,In_333,In_1394);
and U2094 (N_2094,In_952,In_985);
nand U2095 (N_2095,In_73,In_1400);
and U2096 (N_2096,In_473,In_873);
nand U2097 (N_2097,In_372,In_1106);
or U2098 (N_2098,In_9,In_168);
xnor U2099 (N_2099,In_987,In_597);
or U2100 (N_2100,In_692,In_431);
or U2101 (N_2101,In_1196,In_949);
nand U2102 (N_2102,In_541,In_146);
or U2103 (N_2103,In_701,In_69);
xor U2104 (N_2104,In_850,In_1332);
nor U2105 (N_2105,In_565,In_1429);
nor U2106 (N_2106,In_208,In_818);
nor U2107 (N_2107,In_782,In_867);
nor U2108 (N_2108,In_1140,In_685);
and U2109 (N_2109,In_245,In_776);
nor U2110 (N_2110,In_545,In_620);
or U2111 (N_2111,In_323,In_1153);
nor U2112 (N_2112,In_163,In_431);
or U2113 (N_2113,In_3,In_1415);
nand U2114 (N_2114,In_575,In_1437);
and U2115 (N_2115,In_635,In_692);
nand U2116 (N_2116,In_393,In_5);
and U2117 (N_2117,In_856,In_706);
and U2118 (N_2118,In_980,In_1353);
xnor U2119 (N_2119,In_747,In_553);
nand U2120 (N_2120,In_796,In_354);
or U2121 (N_2121,In_526,In_988);
and U2122 (N_2122,In_108,In_571);
or U2123 (N_2123,In_730,In_520);
xor U2124 (N_2124,In_588,In_265);
or U2125 (N_2125,In_998,In_433);
and U2126 (N_2126,In_211,In_1287);
and U2127 (N_2127,In_1025,In_334);
or U2128 (N_2128,In_986,In_368);
nand U2129 (N_2129,In_435,In_1191);
nor U2130 (N_2130,In_1135,In_1327);
nor U2131 (N_2131,In_234,In_669);
nor U2132 (N_2132,In_608,In_1115);
and U2133 (N_2133,In_1215,In_841);
nor U2134 (N_2134,In_757,In_751);
or U2135 (N_2135,In_1171,In_7);
or U2136 (N_2136,In_839,In_1237);
xor U2137 (N_2137,In_1170,In_718);
and U2138 (N_2138,In_1147,In_1145);
nand U2139 (N_2139,In_607,In_322);
and U2140 (N_2140,In_1029,In_1270);
and U2141 (N_2141,In_1203,In_584);
nor U2142 (N_2142,In_1106,In_428);
nand U2143 (N_2143,In_803,In_1338);
or U2144 (N_2144,In_41,In_640);
and U2145 (N_2145,In_1216,In_1464);
nor U2146 (N_2146,In_936,In_870);
nand U2147 (N_2147,In_324,In_1279);
or U2148 (N_2148,In_382,In_950);
or U2149 (N_2149,In_97,In_856);
or U2150 (N_2150,In_666,In_338);
and U2151 (N_2151,In_1478,In_248);
or U2152 (N_2152,In_739,In_571);
nor U2153 (N_2153,In_933,In_952);
or U2154 (N_2154,In_907,In_1207);
nor U2155 (N_2155,In_1083,In_631);
nor U2156 (N_2156,In_869,In_606);
or U2157 (N_2157,In_1490,In_1355);
nand U2158 (N_2158,In_1041,In_1040);
nor U2159 (N_2159,In_700,In_619);
nand U2160 (N_2160,In_1232,In_445);
nand U2161 (N_2161,In_512,In_86);
nand U2162 (N_2162,In_697,In_278);
or U2163 (N_2163,In_207,In_1454);
or U2164 (N_2164,In_755,In_1034);
and U2165 (N_2165,In_192,In_1218);
and U2166 (N_2166,In_540,In_116);
nor U2167 (N_2167,In_161,In_124);
nor U2168 (N_2168,In_314,In_233);
or U2169 (N_2169,In_463,In_662);
or U2170 (N_2170,In_1283,In_502);
and U2171 (N_2171,In_1386,In_920);
nor U2172 (N_2172,In_195,In_1280);
and U2173 (N_2173,In_457,In_966);
or U2174 (N_2174,In_1097,In_1047);
nor U2175 (N_2175,In_330,In_852);
and U2176 (N_2176,In_766,In_24);
or U2177 (N_2177,In_1426,In_309);
or U2178 (N_2178,In_295,In_1048);
or U2179 (N_2179,In_677,In_1223);
nor U2180 (N_2180,In_444,In_1414);
or U2181 (N_2181,In_219,In_747);
and U2182 (N_2182,In_494,In_58);
and U2183 (N_2183,In_933,In_1457);
or U2184 (N_2184,In_1439,In_575);
xnor U2185 (N_2185,In_1050,In_1243);
or U2186 (N_2186,In_1391,In_1332);
nor U2187 (N_2187,In_1171,In_1071);
or U2188 (N_2188,In_431,In_257);
and U2189 (N_2189,In_582,In_241);
or U2190 (N_2190,In_748,In_9);
or U2191 (N_2191,In_231,In_532);
or U2192 (N_2192,In_1490,In_1219);
nor U2193 (N_2193,In_1400,In_139);
nor U2194 (N_2194,In_950,In_1242);
nor U2195 (N_2195,In_569,In_922);
nand U2196 (N_2196,In_1402,In_1239);
xor U2197 (N_2197,In_989,In_394);
nand U2198 (N_2198,In_1407,In_990);
or U2199 (N_2199,In_1087,In_1097);
xnor U2200 (N_2200,In_673,In_607);
nor U2201 (N_2201,In_477,In_846);
nand U2202 (N_2202,In_838,In_1446);
nor U2203 (N_2203,In_820,In_727);
nand U2204 (N_2204,In_648,In_1018);
and U2205 (N_2205,In_637,In_1046);
nand U2206 (N_2206,In_299,In_562);
nand U2207 (N_2207,In_335,In_693);
and U2208 (N_2208,In_465,In_1149);
or U2209 (N_2209,In_1281,In_114);
nor U2210 (N_2210,In_1444,In_1436);
xnor U2211 (N_2211,In_1449,In_161);
or U2212 (N_2212,In_1225,In_547);
nand U2213 (N_2213,In_503,In_281);
nor U2214 (N_2214,In_255,In_1029);
and U2215 (N_2215,In_394,In_707);
or U2216 (N_2216,In_1408,In_1061);
nand U2217 (N_2217,In_943,In_110);
and U2218 (N_2218,In_719,In_794);
nor U2219 (N_2219,In_936,In_1432);
and U2220 (N_2220,In_422,In_53);
and U2221 (N_2221,In_872,In_801);
or U2222 (N_2222,In_1436,In_1439);
nor U2223 (N_2223,In_303,In_620);
nor U2224 (N_2224,In_151,In_422);
xnor U2225 (N_2225,In_663,In_486);
nand U2226 (N_2226,In_1457,In_906);
and U2227 (N_2227,In_852,In_135);
and U2228 (N_2228,In_897,In_1459);
nor U2229 (N_2229,In_1387,In_1284);
and U2230 (N_2230,In_823,In_214);
nor U2231 (N_2231,In_869,In_1231);
or U2232 (N_2232,In_1465,In_996);
or U2233 (N_2233,In_477,In_214);
nand U2234 (N_2234,In_967,In_924);
and U2235 (N_2235,In_825,In_1016);
or U2236 (N_2236,In_1039,In_295);
or U2237 (N_2237,In_872,In_898);
or U2238 (N_2238,In_1225,In_368);
and U2239 (N_2239,In_785,In_1371);
xor U2240 (N_2240,In_241,In_394);
and U2241 (N_2241,In_1394,In_1461);
nand U2242 (N_2242,In_243,In_765);
nand U2243 (N_2243,In_817,In_955);
nand U2244 (N_2244,In_234,In_642);
and U2245 (N_2245,In_85,In_1287);
and U2246 (N_2246,In_842,In_933);
nand U2247 (N_2247,In_687,In_526);
nor U2248 (N_2248,In_1341,In_774);
or U2249 (N_2249,In_1238,In_247);
nand U2250 (N_2250,In_118,In_100);
and U2251 (N_2251,In_153,In_412);
and U2252 (N_2252,In_680,In_282);
and U2253 (N_2253,In_773,In_845);
nor U2254 (N_2254,In_1465,In_144);
nor U2255 (N_2255,In_959,In_725);
or U2256 (N_2256,In_1462,In_388);
nor U2257 (N_2257,In_907,In_904);
nor U2258 (N_2258,In_848,In_1063);
nor U2259 (N_2259,In_534,In_1048);
xor U2260 (N_2260,In_1266,In_1440);
or U2261 (N_2261,In_737,In_1469);
and U2262 (N_2262,In_680,In_1487);
and U2263 (N_2263,In_223,In_1177);
or U2264 (N_2264,In_1177,In_756);
or U2265 (N_2265,In_113,In_87);
nand U2266 (N_2266,In_657,In_1366);
or U2267 (N_2267,In_449,In_779);
or U2268 (N_2268,In_278,In_1016);
nand U2269 (N_2269,In_1143,In_341);
or U2270 (N_2270,In_37,In_1391);
nor U2271 (N_2271,In_582,In_739);
and U2272 (N_2272,In_862,In_699);
nand U2273 (N_2273,In_1087,In_1355);
nand U2274 (N_2274,In_1071,In_598);
xnor U2275 (N_2275,In_103,In_986);
nand U2276 (N_2276,In_61,In_1183);
nor U2277 (N_2277,In_1216,In_529);
or U2278 (N_2278,In_1249,In_814);
nand U2279 (N_2279,In_215,In_1428);
nor U2280 (N_2280,In_450,In_836);
xor U2281 (N_2281,In_405,In_849);
or U2282 (N_2282,In_589,In_1466);
and U2283 (N_2283,In_799,In_1209);
and U2284 (N_2284,In_670,In_1416);
xnor U2285 (N_2285,In_1453,In_212);
and U2286 (N_2286,In_1494,In_644);
nand U2287 (N_2287,In_1104,In_574);
nand U2288 (N_2288,In_1333,In_1430);
and U2289 (N_2289,In_671,In_506);
nor U2290 (N_2290,In_873,In_636);
nor U2291 (N_2291,In_29,In_712);
nor U2292 (N_2292,In_1449,In_1161);
and U2293 (N_2293,In_455,In_666);
nor U2294 (N_2294,In_134,In_694);
and U2295 (N_2295,In_330,In_287);
or U2296 (N_2296,In_279,In_1352);
or U2297 (N_2297,In_131,In_1415);
and U2298 (N_2298,In_1258,In_1022);
or U2299 (N_2299,In_482,In_1371);
and U2300 (N_2300,In_1389,In_810);
nand U2301 (N_2301,In_949,In_818);
or U2302 (N_2302,In_1410,In_821);
or U2303 (N_2303,In_916,In_661);
nand U2304 (N_2304,In_1320,In_1170);
nand U2305 (N_2305,In_1022,In_695);
nor U2306 (N_2306,In_1342,In_831);
and U2307 (N_2307,In_173,In_1491);
nor U2308 (N_2308,In_470,In_81);
nor U2309 (N_2309,In_1109,In_109);
and U2310 (N_2310,In_386,In_1077);
and U2311 (N_2311,In_646,In_1481);
and U2312 (N_2312,In_398,In_553);
and U2313 (N_2313,In_1179,In_28);
nand U2314 (N_2314,In_1075,In_165);
and U2315 (N_2315,In_24,In_444);
xnor U2316 (N_2316,In_193,In_128);
nand U2317 (N_2317,In_1266,In_412);
and U2318 (N_2318,In_561,In_759);
nand U2319 (N_2319,In_241,In_675);
or U2320 (N_2320,In_466,In_808);
and U2321 (N_2321,In_643,In_1034);
and U2322 (N_2322,In_1403,In_664);
xnor U2323 (N_2323,In_746,In_1251);
nand U2324 (N_2324,In_1246,In_1020);
and U2325 (N_2325,In_499,In_1109);
xnor U2326 (N_2326,In_851,In_63);
nand U2327 (N_2327,In_1121,In_283);
or U2328 (N_2328,In_905,In_1043);
or U2329 (N_2329,In_1392,In_91);
xnor U2330 (N_2330,In_932,In_998);
nor U2331 (N_2331,In_1373,In_322);
and U2332 (N_2332,In_1016,In_1354);
and U2333 (N_2333,In_303,In_1168);
or U2334 (N_2334,In_334,In_1287);
or U2335 (N_2335,In_372,In_1294);
nor U2336 (N_2336,In_1326,In_1200);
and U2337 (N_2337,In_1409,In_161);
and U2338 (N_2338,In_414,In_53);
or U2339 (N_2339,In_797,In_924);
and U2340 (N_2340,In_1481,In_673);
nand U2341 (N_2341,In_57,In_498);
nand U2342 (N_2342,In_696,In_781);
nor U2343 (N_2343,In_398,In_778);
nand U2344 (N_2344,In_304,In_863);
or U2345 (N_2345,In_1021,In_1436);
nor U2346 (N_2346,In_515,In_270);
xor U2347 (N_2347,In_475,In_18);
xor U2348 (N_2348,In_534,In_627);
xor U2349 (N_2349,In_651,In_40);
nand U2350 (N_2350,In_617,In_1458);
nand U2351 (N_2351,In_46,In_1247);
or U2352 (N_2352,In_384,In_832);
nand U2353 (N_2353,In_584,In_385);
nor U2354 (N_2354,In_1421,In_1075);
nor U2355 (N_2355,In_1366,In_1368);
or U2356 (N_2356,In_166,In_1053);
xnor U2357 (N_2357,In_769,In_1356);
nor U2358 (N_2358,In_527,In_317);
nor U2359 (N_2359,In_1121,In_1116);
or U2360 (N_2360,In_62,In_1019);
or U2361 (N_2361,In_434,In_1388);
nor U2362 (N_2362,In_1287,In_438);
nand U2363 (N_2363,In_580,In_1274);
nand U2364 (N_2364,In_727,In_752);
nor U2365 (N_2365,In_1324,In_1371);
and U2366 (N_2366,In_1460,In_574);
and U2367 (N_2367,In_654,In_983);
or U2368 (N_2368,In_44,In_1213);
nor U2369 (N_2369,In_821,In_1188);
and U2370 (N_2370,In_1026,In_376);
or U2371 (N_2371,In_722,In_757);
nor U2372 (N_2372,In_345,In_752);
xor U2373 (N_2373,In_1367,In_216);
or U2374 (N_2374,In_301,In_623);
nand U2375 (N_2375,In_702,In_954);
or U2376 (N_2376,In_1318,In_900);
and U2377 (N_2377,In_782,In_1337);
nand U2378 (N_2378,In_122,In_1070);
nor U2379 (N_2379,In_1038,In_861);
nand U2380 (N_2380,In_1285,In_416);
nor U2381 (N_2381,In_12,In_1057);
and U2382 (N_2382,In_1133,In_343);
nor U2383 (N_2383,In_528,In_691);
and U2384 (N_2384,In_1021,In_1246);
nand U2385 (N_2385,In_144,In_26);
and U2386 (N_2386,In_79,In_745);
and U2387 (N_2387,In_532,In_534);
nand U2388 (N_2388,In_1253,In_101);
nand U2389 (N_2389,In_102,In_190);
nand U2390 (N_2390,In_898,In_672);
and U2391 (N_2391,In_346,In_944);
nor U2392 (N_2392,In_645,In_641);
and U2393 (N_2393,In_542,In_30);
xor U2394 (N_2394,In_126,In_570);
or U2395 (N_2395,In_1356,In_1303);
nor U2396 (N_2396,In_1366,In_1428);
and U2397 (N_2397,In_794,In_294);
nand U2398 (N_2398,In_60,In_817);
nor U2399 (N_2399,In_114,In_1030);
and U2400 (N_2400,In_66,In_268);
or U2401 (N_2401,In_521,In_1333);
nand U2402 (N_2402,In_881,In_1069);
nor U2403 (N_2403,In_702,In_1074);
nand U2404 (N_2404,In_653,In_1436);
nand U2405 (N_2405,In_460,In_526);
nor U2406 (N_2406,In_758,In_1297);
and U2407 (N_2407,In_658,In_1321);
xnor U2408 (N_2408,In_1497,In_990);
and U2409 (N_2409,In_180,In_298);
or U2410 (N_2410,In_365,In_839);
and U2411 (N_2411,In_222,In_175);
nor U2412 (N_2412,In_1320,In_603);
nand U2413 (N_2413,In_810,In_1032);
or U2414 (N_2414,In_1038,In_240);
and U2415 (N_2415,In_1137,In_642);
and U2416 (N_2416,In_1490,In_662);
nor U2417 (N_2417,In_1274,In_1060);
and U2418 (N_2418,In_1465,In_168);
and U2419 (N_2419,In_47,In_904);
xor U2420 (N_2420,In_365,In_1164);
nand U2421 (N_2421,In_1471,In_929);
nor U2422 (N_2422,In_705,In_365);
and U2423 (N_2423,In_1352,In_675);
nor U2424 (N_2424,In_1227,In_777);
and U2425 (N_2425,In_1117,In_683);
nand U2426 (N_2426,In_1159,In_923);
and U2427 (N_2427,In_220,In_551);
nor U2428 (N_2428,In_1493,In_1322);
nor U2429 (N_2429,In_659,In_988);
nor U2430 (N_2430,In_230,In_1241);
nor U2431 (N_2431,In_1448,In_684);
and U2432 (N_2432,In_346,In_755);
and U2433 (N_2433,In_1085,In_1165);
nand U2434 (N_2434,In_1146,In_872);
nor U2435 (N_2435,In_198,In_596);
nand U2436 (N_2436,In_28,In_1024);
nor U2437 (N_2437,In_937,In_898);
and U2438 (N_2438,In_774,In_8);
and U2439 (N_2439,In_127,In_155);
nand U2440 (N_2440,In_701,In_711);
nand U2441 (N_2441,In_1229,In_1202);
nand U2442 (N_2442,In_108,In_523);
or U2443 (N_2443,In_995,In_1461);
or U2444 (N_2444,In_188,In_776);
nand U2445 (N_2445,In_840,In_42);
nor U2446 (N_2446,In_115,In_1200);
or U2447 (N_2447,In_808,In_1111);
nor U2448 (N_2448,In_291,In_1076);
and U2449 (N_2449,In_935,In_86);
nor U2450 (N_2450,In_883,In_36);
nand U2451 (N_2451,In_817,In_885);
or U2452 (N_2452,In_780,In_385);
or U2453 (N_2453,In_1132,In_598);
nor U2454 (N_2454,In_630,In_914);
nor U2455 (N_2455,In_1310,In_52);
nand U2456 (N_2456,In_1272,In_777);
or U2457 (N_2457,In_112,In_1309);
nand U2458 (N_2458,In_853,In_247);
or U2459 (N_2459,In_77,In_289);
and U2460 (N_2460,In_78,In_1358);
or U2461 (N_2461,In_1375,In_819);
nor U2462 (N_2462,In_837,In_541);
nand U2463 (N_2463,In_171,In_463);
nand U2464 (N_2464,In_1012,In_80);
xnor U2465 (N_2465,In_261,In_968);
nor U2466 (N_2466,In_1413,In_34);
or U2467 (N_2467,In_611,In_1068);
nor U2468 (N_2468,In_57,In_1257);
nand U2469 (N_2469,In_868,In_1416);
nor U2470 (N_2470,In_566,In_561);
nand U2471 (N_2471,In_164,In_1108);
and U2472 (N_2472,In_1471,In_1261);
or U2473 (N_2473,In_894,In_1032);
or U2474 (N_2474,In_1025,In_860);
xnor U2475 (N_2475,In_1044,In_1441);
nor U2476 (N_2476,In_1246,In_175);
nand U2477 (N_2477,In_1119,In_1303);
or U2478 (N_2478,In_494,In_1454);
nor U2479 (N_2479,In_150,In_223);
nor U2480 (N_2480,In_712,In_1047);
and U2481 (N_2481,In_458,In_859);
or U2482 (N_2482,In_80,In_319);
or U2483 (N_2483,In_498,In_768);
or U2484 (N_2484,In_166,In_703);
and U2485 (N_2485,In_478,In_1118);
or U2486 (N_2486,In_1308,In_1334);
xor U2487 (N_2487,In_873,In_1446);
nor U2488 (N_2488,In_461,In_446);
and U2489 (N_2489,In_1091,In_179);
or U2490 (N_2490,In_354,In_1372);
or U2491 (N_2491,In_1021,In_1423);
nor U2492 (N_2492,In_513,In_775);
nor U2493 (N_2493,In_392,In_869);
and U2494 (N_2494,In_337,In_1291);
nand U2495 (N_2495,In_30,In_931);
or U2496 (N_2496,In_832,In_396);
nor U2497 (N_2497,In_864,In_1476);
nor U2498 (N_2498,In_986,In_446);
nand U2499 (N_2499,In_915,In_1363);
and U2500 (N_2500,In_288,In_1345);
or U2501 (N_2501,In_1396,In_390);
and U2502 (N_2502,In_508,In_322);
nand U2503 (N_2503,In_81,In_986);
xor U2504 (N_2504,In_882,In_792);
and U2505 (N_2505,In_73,In_381);
and U2506 (N_2506,In_578,In_768);
or U2507 (N_2507,In_98,In_1149);
nor U2508 (N_2508,In_646,In_869);
nor U2509 (N_2509,In_1146,In_914);
xnor U2510 (N_2510,In_1382,In_1108);
and U2511 (N_2511,In_525,In_202);
xor U2512 (N_2512,In_1049,In_1173);
nor U2513 (N_2513,In_230,In_208);
xor U2514 (N_2514,In_1467,In_470);
nand U2515 (N_2515,In_264,In_262);
and U2516 (N_2516,In_687,In_1185);
and U2517 (N_2517,In_1094,In_175);
nor U2518 (N_2518,In_1403,In_1080);
and U2519 (N_2519,In_145,In_1234);
and U2520 (N_2520,In_942,In_1362);
or U2521 (N_2521,In_315,In_360);
nand U2522 (N_2522,In_171,In_818);
nand U2523 (N_2523,In_69,In_243);
or U2524 (N_2524,In_761,In_511);
or U2525 (N_2525,In_253,In_441);
and U2526 (N_2526,In_536,In_680);
nor U2527 (N_2527,In_736,In_208);
and U2528 (N_2528,In_102,In_681);
and U2529 (N_2529,In_11,In_756);
and U2530 (N_2530,In_795,In_696);
and U2531 (N_2531,In_1078,In_196);
and U2532 (N_2532,In_1165,In_234);
nand U2533 (N_2533,In_879,In_1197);
xnor U2534 (N_2534,In_1494,In_303);
nand U2535 (N_2535,In_915,In_1076);
nand U2536 (N_2536,In_465,In_323);
or U2537 (N_2537,In_782,In_453);
nand U2538 (N_2538,In_323,In_1479);
or U2539 (N_2539,In_952,In_1191);
nand U2540 (N_2540,In_359,In_625);
or U2541 (N_2541,In_482,In_601);
nor U2542 (N_2542,In_931,In_1091);
nor U2543 (N_2543,In_1436,In_543);
nand U2544 (N_2544,In_765,In_76);
or U2545 (N_2545,In_1326,In_13);
or U2546 (N_2546,In_1053,In_1271);
and U2547 (N_2547,In_341,In_1025);
or U2548 (N_2548,In_915,In_1176);
nand U2549 (N_2549,In_244,In_1048);
and U2550 (N_2550,In_1222,In_510);
nand U2551 (N_2551,In_240,In_20);
and U2552 (N_2552,In_891,In_119);
nand U2553 (N_2553,In_852,In_1388);
nor U2554 (N_2554,In_498,In_1359);
nand U2555 (N_2555,In_166,In_544);
nor U2556 (N_2556,In_390,In_277);
nand U2557 (N_2557,In_1261,In_990);
nor U2558 (N_2558,In_241,In_1163);
nand U2559 (N_2559,In_1002,In_192);
or U2560 (N_2560,In_262,In_806);
nand U2561 (N_2561,In_986,In_1386);
nor U2562 (N_2562,In_1183,In_210);
nor U2563 (N_2563,In_301,In_1262);
and U2564 (N_2564,In_1258,In_942);
nor U2565 (N_2565,In_1249,In_1407);
or U2566 (N_2566,In_1486,In_378);
nand U2567 (N_2567,In_112,In_386);
nand U2568 (N_2568,In_261,In_1248);
or U2569 (N_2569,In_6,In_1464);
nor U2570 (N_2570,In_496,In_636);
nand U2571 (N_2571,In_1285,In_820);
nand U2572 (N_2572,In_550,In_643);
and U2573 (N_2573,In_174,In_336);
and U2574 (N_2574,In_197,In_955);
nand U2575 (N_2575,In_155,In_1203);
nand U2576 (N_2576,In_698,In_646);
or U2577 (N_2577,In_1304,In_776);
nor U2578 (N_2578,In_62,In_658);
nor U2579 (N_2579,In_1065,In_976);
nand U2580 (N_2580,In_172,In_125);
nand U2581 (N_2581,In_645,In_931);
nor U2582 (N_2582,In_1165,In_181);
or U2583 (N_2583,In_1465,In_446);
nor U2584 (N_2584,In_521,In_464);
or U2585 (N_2585,In_313,In_462);
nor U2586 (N_2586,In_798,In_293);
nor U2587 (N_2587,In_445,In_1239);
nand U2588 (N_2588,In_586,In_657);
or U2589 (N_2589,In_1242,In_753);
nor U2590 (N_2590,In_1476,In_1362);
and U2591 (N_2591,In_1146,In_318);
nand U2592 (N_2592,In_234,In_341);
xor U2593 (N_2593,In_566,In_1320);
nor U2594 (N_2594,In_1103,In_1231);
and U2595 (N_2595,In_955,In_271);
or U2596 (N_2596,In_1431,In_1456);
nand U2597 (N_2597,In_1421,In_834);
nand U2598 (N_2598,In_373,In_1449);
and U2599 (N_2599,In_1063,In_674);
or U2600 (N_2600,In_728,In_481);
or U2601 (N_2601,In_446,In_1482);
and U2602 (N_2602,In_190,In_1289);
nor U2603 (N_2603,In_1274,In_281);
or U2604 (N_2604,In_394,In_865);
nor U2605 (N_2605,In_1345,In_428);
xor U2606 (N_2606,In_287,In_415);
nor U2607 (N_2607,In_1365,In_588);
or U2608 (N_2608,In_838,In_51);
nor U2609 (N_2609,In_877,In_1317);
nor U2610 (N_2610,In_1011,In_490);
nor U2611 (N_2611,In_243,In_900);
or U2612 (N_2612,In_310,In_1466);
or U2613 (N_2613,In_10,In_187);
nand U2614 (N_2614,In_1063,In_902);
nor U2615 (N_2615,In_175,In_386);
or U2616 (N_2616,In_123,In_1242);
nand U2617 (N_2617,In_1139,In_1021);
nand U2618 (N_2618,In_517,In_1079);
nor U2619 (N_2619,In_218,In_572);
or U2620 (N_2620,In_609,In_1068);
or U2621 (N_2621,In_1359,In_362);
xor U2622 (N_2622,In_344,In_1425);
nor U2623 (N_2623,In_691,In_1203);
nor U2624 (N_2624,In_961,In_145);
and U2625 (N_2625,In_392,In_629);
nand U2626 (N_2626,In_907,In_1368);
nor U2627 (N_2627,In_406,In_1006);
nand U2628 (N_2628,In_382,In_346);
nor U2629 (N_2629,In_1154,In_1073);
or U2630 (N_2630,In_782,In_1127);
and U2631 (N_2631,In_754,In_1342);
or U2632 (N_2632,In_357,In_905);
or U2633 (N_2633,In_1458,In_1110);
and U2634 (N_2634,In_667,In_800);
and U2635 (N_2635,In_722,In_969);
nand U2636 (N_2636,In_544,In_1323);
xnor U2637 (N_2637,In_501,In_697);
nor U2638 (N_2638,In_225,In_1479);
nor U2639 (N_2639,In_1474,In_156);
nor U2640 (N_2640,In_208,In_48);
or U2641 (N_2641,In_561,In_1069);
and U2642 (N_2642,In_1073,In_629);
or U2643 (N_2643,In_1220,In_606);
nand U2644 (N_2644,In_520,In_73);
and U2645 (N_2645,In_793,In_513);
and U2646 (N_2646,In_798,In_1485);
nor U2647 (N_2647,In_979,In_46);
nand U2648 (N_2648,In_1421,In_636);
or U2649 (N_2649,In_590,In_852);
nor U2650 (N_2650,In_518,In_184);
xor U2651 (N_2651,In_160,In_450);
nand U2652 (N_2652,In_419,In_871);
nor U2653 (N_2653,In_734,In_258);
xnor U2654 (N_2654,In_783,In_1034);
nor U2655 (N_2655,In_417,In_383);
nand U2656 (N_2656,In_998,In_13);
xnor U2657 (N_2657,In_702,In_533);
and U2658 (N_2658,In_380,In_946);
and U2659 (N_2659,In_912,In_657);
or U2660 (N_2660,In_1421,In_1015);
and U2661 (N_2661,In_723,In_357);
or U2662 (N_2662,In_97,In_1092);
nor U2663 (N_2663,In_1255,In_566);
and U2664 (N_2664,In_623,In_398);
or U2665 (N_2665,In_1368,In_198);
nor U2666 (N_2666,In_865,In_822);
nand U2667 (N_2667,In_318,In_213);
nor U2668 (N_2668,In_1118,In_581);
nor U2669 (N_2669,In_1412,In_15);
xor U2670 (N_2670,In_622,In_1037);
nand U2671 (N_2671,In_353,In_1425);
nor U2672 (N_2672,In_239,In_555);
or U2673 (N_2673,In_701,In_770);
xnor U2674 (N_2674,In_1493,In_173);
or U2675 (N_2675,In_374,In_378);
and U2676 (N_2676,In_721,In_1200);
nor U2677 (N_2677,In_1296,In_340);
nor U2678 (N_2678,In_376,In_249);
nand U2679 (N_2679,In_632,In_162);
nand U2680 (N_2680,In_1010,In_869);
or U2681 (N_2681,In_1467,In_586);
or U2682 (N_2682,In_1123,In_846);
nand U2683 (N_2683,In_1048,In_198);
xnor U2684 (N_2684,In_1253,In_1116);
nand U2685 (N_2685,In_1167,In_442);
xor U2686 (N_2686,In_964,In_1319);
or U2687 (N_2687,In_705,In_1003);
or U2688 (N_2688,In_1173,In_1279);
nand U2689 (N_2689,In_425,In_253);
nor U2690 (N_2690,In_599,In_225);
nor U2691 (N_2691,In_1359,In_77);
nor U2692 (N_2692,In_826,In_1190);
nor U2693 (N_2693,In_211,In_1130);
and U2694 (N_2694,In_1016,In_892);
nand U2695 (N_2695,In_1386,In_1367);
nor U2696 (N_2696,In_160,In_168);
or U2697 (N_2697,In_668,In_969);
nor U2698 (N_2698,In_19,In_898);
xor U2699 (N_2699,In_61,In_1140);
nor U2700 (N_2700,In_580,In_54);
nand U2701 (N_2701,In_1255,In_809);
nor U2702 (N_2702,In_587,In_1304);
nor U2703 (N_2703,In_676,In_1053);
nor U2704 (N_2704,In_540,In_817);
nand U2705 (N_2705,In_1278,In_784);
and U2706 (N_2706,In_590,In_1199);
and U2707 (N_2707,In_949,In_621);
or U2708 (N_2708,In_1378,In_878);
and U2709 (N_2709,In_490,In_20);
and U2710 (N_2710,In_277,In_1419);
xnor U2711 (N_2711,In_1240,In_501);
nor U2712 (N_2712,In_1240,In_599);
or U2713 (N_2713,In_1417,In_631);
and U2714 (N_2714,In_263,In_1261);
nor U2715 (N_2715,In_635,In_975);
and U2716 (N_2716,In_1268,In_1206);
nand U2717 (N_2717,In_175,In_564);
and U2718 (N_2718,In_933,In_1331);
or U2719 (N_2719,In_45,In_1042);
nand U2720 (N_2720,In_1117,In_529);
nor U2721 (N_2721,In_979,In_1284);
nor U2722 (N_2722,In_1470,In_617);
nand U2723 (N_2723,In_1301,In_37);
or U2724 (N_2724,In_1023,In_82);
and U2725 (N_2725,In_182,In_1308);
nor U2726 (N_2726,In_781,In_1181);
and U2727 (N_2727,In_178,In_1383);
and U2728 (N_2728,In_1492,In_1021);
xor U2729 (N_2729,In_0,In_868);
nand U2730 (N_2730,In_73,In_28);
nand U2731 (N_2731,In_713,In_645);
xnor U2732 (N_2732,In_700,In_1057);
and U2733 (N_2733,In_206,In_194);
or U2734 (N_2734,In_1082,In_1318);
nand U2735 (N_2735,In_231,In_1454);
or U2736 (N_2736,In_1226,In_635);
nand U2737 (N_2737,In_1184,In_1490);
nor U2738 (N_2738,In_263,In_291);
nand U2739 (N_2739,In_800,In_981);
and U2740 (N_2740,In_1325,In_1421);
and U2741 (N_2741,In_679,In_839);
xor U2742 (N_2742,In_571,In_1283);
nand U2743 (N_2743,In_24,In_906);
and U2744 (N_2744,In_149,In_292);
nor U2745 (N_2745,In_1461,In_1401);
nor U2746 (N_2746,In_242,In_1095);
nand U2747 (N_2747,In_463,In_152);
and U2748 (N_2748,In_653,In_655);
nand U2749 (N_2749,In_646,In_444);
and U2750 (N_2750,In_918,In_230);
or U2751 (N_2751,In_1119,In_1404);
xor U2752 (N_2752,In_1480,In_47);
nor U2753 (N_2753,In_107,In_311);
or U2754 (N_2754,In_319,In_560);
and U2755 (N_2755,In_362,In_428);
and U2756 (N_2756,In_1101,In_599);
or U2757 (N_2757,In_786,In_192);
xor U2758 (N_2758,In_824,In_378);
nand U2759 (N_2759,In_1320,In_1013);
nand U2760 (N_2760,In_419,In_1347);
nor U2761 (N_2761,In_1090,In_1446);
or U2762 (N_2762,In_1288,In_1127);
xnor U2763 (N_2763,In_1343,In_649);
and U2764 (N_2764,In_947,In_1196);
nor U2765 (N_2765,In_964,In_1012);
and U2766 (N_2766,In_687,In_1364);
xor U2767 (N_2767,In_55,In_1377);
nor U2768 (N_2768,In_963,In_1075);
nor U2769 (N_2769,In_173,In_1198);
nand U2770 (N_2770,In_1278,In_332);
xor U2771 (N_2771,In_968,In_370);
and U2772 (N_2772,In_1013,In_641);
or U2773 (N_2773,In_396,In_1427);
nor U2774 (N_2774,In_1021,In_81);
or U2775 (N_2775,In_1137,In_478);
nor U2776 (N_2776,In_1059,In_630);
nand U2777 (N_2777,In_1459,In_1225);
and U2778 (N_2778,In_1080,In_1448);
nor U2779 (N_2779,In_1447,In_242);
and U2780 (N_2780,In_1029,In_1234);
or U2781 (N_2781,In_193,In_1449);
nand U2782 (N_2782,In_1458,In_308);
nor U2783 (N_2783,In_668,In_112);
xnor U2784 (N_2784,In_548,In_1289);
nor U2785 (N_2785,In_246,In_33);
and U2786 (N_2786,In_424,In_751);
or U2787 (N_2787,In_763,In_544);
xor U2788 (N_2788,In_1345,In_956);
and U2789 (N_2789,In_1426,In_400);
nor U2790 (N_2790,In_1407,In_1481);
nand U2791 (N_2791,In_635,In_582);
xor U2792 (N_2792,In_1393,In_790);
nand U2793 (N_2793,In_131,In_1432);
or U2794 (N_2794,In_277,In_420);
nor U2795 (N_2795,In_307,In_1118);
nand U2796 (N_2796,In_1206,In_816);
nand U2797 (N_2797,In_944,In_870);
nand U2798 (N_2798,In_25,In_28);
nand U2799 (N_2799,In_279,In_551);
nor U2800 (N_2800,In_851,In_900);
and U2801 (N_2801,In_679,In_562);
and U2802 (N_2802,In_803,In_1351);
nor U2803 (N_2803,In_650,In_658);
nand U2804 (N_2804,In_1446,In_1015);
and U2805 (N_2805,In_1043,In_1045);
or U2806 (N_2806,In_528,In_300);
and U2807 (N_2807,In_268,In_278);
nor U2808 (N_2808,In_941,In_687);
nor U2809 (N_2809,In_1448,In_1494);
nor U2810 (N_2810,In_517,In_1395);
or U2811 (N_2811,In_321,In_778);
nor U2812 (N_2812,In_413,In_583);
nor U2813 (N_2813,In_408,In_603);
nor U2814 (N_2814,In_761,In_529);
nor U2815 (N_2815,In_380,In_442);
nor U2816 (N_2816,In_548,In_1453);
or U2817 (N_2817,In_1083,In_1385);
nand U2818 (N_2818,In_1093,In_1128);
nor U2819 (N_2819,In_1493,In_688);
and U2820 (N_2820,In_1005,In_316);
nand U2821 (N_2821,In_321,In_1353);
and U2822 (N_2822,In_263,In_681);
and U2823 (N_2823,In_937,In_1208);
or U2824 (N_2824,In_1362,In_798);
nor U2825 (N_2825,In_1391,In_1146);
or U2826 (N_2826,In_1418,In_293);
nor U2827 (N_2827,In_313,In_627);
or U2828 (N_2828,In_193,In_966);
and U2829 (N_2829,In_5,In_118);
and U2830 (N_2830,In_1107,In_660);
nand U2831 (N_2831,In_532,In_804);
xor U2832 (N_2832,In_267,In_451);
or U2833 (N_2833,In_1076,In_821);
and U2834 (N_2834,In_604,In_688);
or U2835 (N_2835,In_1087,In_834);
and U2836 (N_2836,In_182,In_1012);
and U2837 (N_2837,In_355,In_1191);
nor U2838 (N_2838,In_246,In_1059);
xnor U2839 (N_2839,In_921,In_497);
xor U2840 (N_2840,In_781,In_638);
or U2841 (N_2841,In_991,In_1190);
or U2842 (N_2842,In_153,In_533);
xor U2843 (N_2843,In_984,In_272);
nand U2844 (N_2844,In_1039,In_1172);
or U2845 (N_2845,In_1178,In_1382);
nand U2846 (N_2846,In_1495,In_1436);
or U2847 (N_2847,In_163,In_89);
nand U2848 (N_2848,In_1150,In_990);
nand U2849 (N_2849,In_608,In_1311);
nand U2850 (N_2850,In_947,In_333);
nor U2851 (N_2851,In_826,In_1046);
or U2852 (N_2852,In_1230,In_1318);
nand U2853 (N_2853,In_894,In_168);
and U2854 (N_2854,In_987,In_772);
nor U2855 (N_2855,In_1368,In_945);
and U2856 (N_2856,In_304,In_633);
or U2857 (N_2857,In_1285,In_708);
and U2858 (N_2858,In_968,In_1335);
and U2859 (N_2859,In_826,In_7);
xnor U2860 (N_2860,In_1415,In_427);
xnor U2861 (N_2861,In_487,In_1153);
or U2862 (N_2862,In_526,In_42);
or U2863 (N_2863,In_1405,In_1057);
nor U2864 (N_2864,In_545,In_88);
or U2865 (N_2865,In_921,In_841);
nand U2866 (N_2866,In_433,In_1352);
xnor U2867 (N_2867,In_134,In_378);
or U2868 (N_2868,In_66,In_312);
xor U2869 (N_2869,In_97,In_284);
nor U2870 (N_2870,In_409,In_1047);
nand U2871 (N_2871,In_460,In_1177);
nor U2872 (N_2872,In_340,In_601);
xnor U2873 (N_2873,In_11,In_1412);
nor U2874 (N_2874,In_479,In_702);
and U2875 (N_2875,In_971,In_1200);
and U2876 (N_2876,In_409,In_720);
xor U2877 (N_2877,In_589,In_57);
or U2878 (N_2878,In_221,In_1095);
xnor U2879 (N_2879,In_1123,In_430);
or U2880 (N_2880,In_68,In_494);
nand U2881 (N_2881,In_1285,In_1319);
or U2882 (N_2882,In_626,In_1260);
or U2883 (N_2883,In_1479,In_821);
or U2884 (N_2884,In_954,In_521);
and U2885 (N_2885,In_1442,In_1336);
xor U2886 (N_2886,In_1429,In_1367);
and U2887 (N_2887,In_660,In_1084);
or U2888 (N_2888,In_861,In_181);
nor U2889 (N_2889,In_1438,In_597);
and U2890 (N_2890,In_956,In_358);
nand U2891 (N_2891,In_178,In_1195);
and U2892 (N_2892,In_911,In_720);
nand U2893 (N_2893,In_1040,In_614);
nor U2894 (N_2894,In_1409,In_1126);
and U2895 (N_2895,In_612,In_1019);
nor U2896 (N_2896,In_812,In_1007);
and U2897 (N_2897,In_975,In_1250);
and U2898 (N_2898,In_430,In_36);
nand U2899 (N_2899,In_346,In_741);
nand U2900 (N_2900,In_723,In_313);
nand U2901 (N_2901,In_856,In_950);
nand U2902 (N_2902,In_839,In_785);
and U2903 (N_2903,In_1420,In_342);
and U2904 (N_2904,In_1152,In_509);
or U2905 (N_2905,In_1246,In_1222);
nand U2906 (N_2906,In_305,In_502);
nor U2907 (N_2907,In_1140,In_1097);
or U2908 (N_2908,In_573,In_519);
nor U2909 (N_2909,In_367,In_934);
nor U2910 (N_2910,In_1008,In_268);
nor U2911 (N_2911,In_356,In_455);
or U2912 (N_2912,In_1426,In_1391);
nor U2913 (N_2913,In_837,In_466);
nand U2914 (N_2914,In_1278,In_53);
nand U2915 (N_2915,In_723,In_628);
or U2916 (N_2916,In_861,In_990);
nor U2917 (N_2917,In_722,In_1097);
or U2918 (N_2918,In_1488,In_245);
nor U2919 (N_2919,In_212,In_560);
and U2920 (N_2920,In_1071,In_469);
nor U2921 (N_2921,In_40,In_903);
nor U2922 (N_2922,In_183,In_117);
and U2923 (N_2923,In_415,In_800);
or U2924 (N_2924,In_984,In_1284);
or U2925 (N_2925,In_1095,In_354);
nor U2926 (N_2926,In_1180,In_1011);
nand U2927 (N_2927,In_1254,In_1476);
nor U2928 (N_2928,In_1295,In_742);
nand U2929 (N_2929,In_182,In_404);
nand U2930 (N_2930,In_703,In_1296);
and U2931 (N_2931,In_627,In_1163);
nor U2932 (N_2932,In_926,In_224);
and U2933 (N_2933,In_903,In_616);
and U2934 (N_2934,In_685,In_1379);
nand U2935 (N_2935,In_261,In_114);
nand U2936 (N_2936,In_478,In_758);
or U2937 (N_2937,In_484,In_832);
nor U2938 (N_2938,In_1312,In_883);
nor U2939 (N_2939,In_924,In_1105);
nor U2940 (N_2940,In_1018,In_1203);
or U2941 (N_2941,In_1410,In_818);
and U2942 (N_2942,In_1463,In_564);
or U2943 (N_2943,In_528,In_583);
nor U2944 (N_2944,In_448,In_1170);
nand U2945 (N_2945,In_311,In_1376);
and U2946 (N_2946,In_1228,In_882);
or U2947 (N_2947,In_1105,In_42);
nand U2948 (N_2948,In_1237,In_615);
nor U2949 (N_2949,In_768,In_1412);
nand U2950 (N_2950,In_44,In_249);
nor U2951 (N_2951,In_1346,In_648);
nor U2952 (N_2952,In_204,In_1087);
nor U2953 (N_2953,In_1367,In_506);
nor U2954 (N_2954,In_545,In_455);
nand U2955 (N_2955,In_564,In_1368);
or U2956 (N_2956,In_268,In_354);
nor U2957 (N_2957,In_523,In_51);
or U2958 (N_2958,In_277,In_1349);
and U2959 (N_2959,In_805,In_505);
nand U2960 (N_2960,In_116,In_1287);
nor U2961 (N_2961,In_992,In_309);
nand U2962 (N_2962,In_560,In_660);
and U2963 (N_2963,In_249,In_467);
nor U2964 (N_2964,In_78,In_164);
nor U2965 (N_2965,In_677,In_518);
and U2966 (N_2966,In_1179,In_582);
or U2967 (N_2967,In_611,In_647);
nand U2968 (N_2968,In_859,In_1461);
or U2969 (N_2969,In_1189,In_1020);
or U2970 (N_2970,In_565,In_635);
or U2971 (N_2971,In_1430,In_1044);
and U2972 (N_2972,In_673,In_363);
xnor U2973 (N_2973,In_1120,In_943);
and U2974 (N_2974,In_120,In_777);
nor U2975 (N_2975,In_1314,In_972);
nor U2976 (N_2976,In_1247,In_1181);
and U2977 (N_2977,In_984,In_305);
and U2978 (N_2978,In_978,In_1045);
nor U2979 (N_2979,In_1299,In_1170);
nor U2980 (N_2980,In_1102,In_957);
or U2981 (N_2981,In_399,In_338);
nor U2982 (N_2982,In_974,In_1296);
nor U2983 (N_2983,In_846,In_1486);
or U2984 (N_2984,In_603,In_813);
xor U2985 (N_2985,In_831,In_1439);
nand U2986 (N_2986,In_755,In_609);
and U2987 (N_2987,In_81,In_1397);
nand U2988 (N_2988,In_122,In_720);
nand U2989 (N_2989,In_157,In_964);
nor U2990 (N_2990,In_928,In_992);
or U2991 (N_2991,In_99,In_494);
or U2992 (N_2992,In_1040,In_661);
nand U2993 (N_2993,In_352,In_1178);
nand U2994 (N_2994,In_957,In_1360);
or U2995 (N_2995,In_494,In_817);
nor U2996 (N_2996,In_1045,In_1264);
xor U2997 (N_2997,In_672,In_429);
nand U2998 (N_2998,In_893,In_155);
or U2999 (N_2999,In_1027,In_1253);
and U3000 (N_3000,In_1102,In_1497);
or U3001 (N_3001,In_838,In_762);
or U3002 (N_3002,In_60,In_744);
and U3003 (N_3003,In_238,In_1122);
nor U3004 (N_3004,In_293,In_1105);
and U3005 (N_3005,In_1464,In_1284);
or U3006 (N_3006,In_462,In_86);
or U3007 (N_3007,In_80,In_1289);
and U3008 (N_3008,In_757,In_252);
nand U3009 (N_3009,In_1257,In_302);
and U3010 (N_3010,In_664,In_1055);
xor U3011 (N_3011,In_417,In_814);
nand U3012 (N_3012,In_1263,In_655);
and U3013 (N_3013,In_1002,In_1442);
nor U3014 (N_3014,In_447,In_227);
and U3015 (N_3015,In_339,In_1278);
and U3016 (N_3016,In_564,In_237);
and U3017 (N_3017,In_525,In_1418);
or U3018 (N_3018,In_1041,In_962);
nand U3019 (N_3019,In_658,In_1032);
or U3020 (N_3020,In_1262,In_551);
and U3021 (N_3021,In_1367,In_211);
nor U3022 (N_3022,In_1459,In_1120);
and U3023 (N_3023,In_314,In_1424);
or U3024 (N_3024,In_1152,In_783);
nor U3025 (N_3025,In_113,In_1027);
or U3026 (N_3026,In_489,In_594);
nor U3027 (N_3027,In_1462,In_344);
and U3028 (N_3028,In_1381,In_549);
xnor U3029 (N_3029,In_1309,In_818);
and U3030 (N_3030,In_767,In_649);
xnor U3031 (N_3031,In_446,In_311);
nor U3032 (N_3032,In_1009,In_963);
xnor U3033 (N_3033,In_1355,In_506);
and U3034 (N_3034,In_845,In_811);
or U3035 (N_3035,In_406,In_1118);
nor U3036 (N_3036,In_626,In_611);
nand U3037 (N_3037,In_78,In_1183);
and U3038 (N_3038,In_160,In_948);
nor U3039 (N_3039,In_1077,In_394);
nor U3040 (N_3040,In_617,In_975);
xor U3041 (N_3041,In_1155,In_283);
nor U3042 (N_3042,In_270,In_1037);
nand U3043 (N_3043,In_105,In_1311);
or U3044 (N_3044,In_710,In_388);
nand U3045 (N_3045,In_34,In_1025);
nand U3046 (N_3046,In_556,In_62);
nor U3047 (N_3047,In_76,In_530);
nand U3048 (N_3048,In_623,In_1173);
nand U3049 (N_3049,In_462,In_59);
nand U3050 (N_3050,In_1072,In_555);
or U3051 (N_3051,In_1194,In_1392);
nor U3052 (N_3052,In_717,In_1194);
and U3053 (N_3053,In_82,In_975);
or U3054 (N_3054,In_1492,In_656);
and U3055 (N_3055,In_698,In_99);
xor U3056 (N_3056,In_426,In_1362);
nor U3057 (N_3057,In_283,In_435);
nor U3058 (N_3058,In_1464,In_55);
nor U3059 (N_3059,In_1249,In_365);
or U3060 (N_3060,In_952,In_670);
and U3061 (N_3061,In_359,In_907);
or U3062 (N_3062,In_1295,In_221);
nand U3063 (N_3063,In_1475,In_456);
nand U3064 (N_3064,In_1243,In_971);
nor U3065 (N_3065,In_210,In_1071);
xnor U3066 (N_3066,In_630,In_13);
and U3067 (N_3067,In_913,In_1130);
nand U3068 (N_3068,In_1246,In_0);
nor U3069 (N_3069,In_1206,In_598);
nand U3070 (N_3070,In_1281,In_211);
or U3071 (N_3071,In_195,In_835);
or U3072 (N_3072,In_461,In_634);
and U3073 (N_3073,In_1333,In_469);
and U3074 (N_3074,In_1183,In_104);
nand U3075 (N_3075,In_957,In_820);
nand U3076 (N_3076,In_1099,In_409);
and U3077 (N_3077,In_669,In_1003);
or U3078 (N_3078,In_1404,In_319);
nand U3079 (N_3079,In_1448,In_1423);
nand U3080 (N_3080,In_808,In_141);
xnor U3081 (N_3081,In_380,In_310);
nor U3082 (N_3082,In_1038,In_599);
and U3083 (N_3083,In_147,In_1101);
xnor U3084 (N_3084,In_276,In_315);
or U3085 (N_3085,In_1140,In_467);
nand U3086 (N_3086,In_1081,In_298);
or U3087 (N_3087,In_214,In_904);
and U3088 (N_3088,In_224,In_917);
nand U3089 (N_3089,In_891,In_692);
xor U3090 (N_3090,In_699,In_351);
or U3091 (N_3091,In_138,In_28);
or U3092 (N_3092,In_601,In_237);
or U3093 (N_3093,In_57,In_870);
and U3094 (N_3094,In_431,In_12);
xnor U3095 (N_3095,In_1302,In_591);
xnor U3096 (N_3096,In_830,In_201);
nor U3097 (N_3097,In_470,In_771);
nand U3098 (N_3098,In_168,In_211);
and U3099 (N_3099,In_1348,In_1246);
nand U3100 (N_3100,In_391,In_597);
or U3101 (N_3101,In_1307,In_688);
nand U3102 (N_3102,In_252,In_1484);
nand U3103 (N_3103,In_842,In_1355);
and U3104 (N_3104,In_663,In_710);
or U3105 (N_3105,In_222,In_312);
and U3106 (N_3106,In_1199,In_1083);
nor U3107 (N_3107,In_1039,In_973);
xor U3108 (N_3108,In_322,In_211);
nor U3109 (N_3109,In_1418,In_1031);
nand U3110 (N_3110,In_1021,In_631);
and U3111 (N_3111,In_1348,In_1495);
and U3112 (N_3112,In_254,In_294);
nor U3113 (N_3113,In_948,In_81);
or U3114 (N_3114,In_1085,In_287);
nand U3115 (N_3115,In_113,In_36);
nor U3116 (N_3116,In_489,In_516);
nor U3117 (N_3117,In_1091,In_113);
or U3118 (N_3118,In_694,In_526);
and U3119 (N_3119,In_781,In_1183);
or U3120 (N_3120,In_145,In_756);
nor U3121 (N_3121,In_490,In_618);
nor U3122 (N_3122,In_1139,In_833);
nor U3123 (N_3123,In_843,In_427);
nand U3124 (N_3124,In_502,In_351);
and U3125 (N_3125,In_1185,In_1336);
and U3126 (N_3126,In_242,In_1398);
nor U3127 (N_3127,In_421,In_432);
or U3128 (N_3128,In_55,In_253);
nor U3129 (N_3129,In_901,In_373);
xor U3130 (N_3130,In_1177,In_1235);
or U3131 (N_3131,In_423,In_1345);
or U3132 (N_3132,In_617,In_358);
or U3133 (N_3133,In_1171,In_1061);
nor U3134 (N_3134,In_866,In_598);
nor U3135 (N_3135,In_658,In_704);
nor U3136 (N_3136,In_175,In_117);
or U3137 (N_3137,In_1460,In_1318);
nand U3138 (N_3138,In_32,In_831);
xor U3139 (N_3139,In_411,In_1404);
and U3140 (N_3140,In_1044,In_731);
and U3141 (N_3141,In_284,In_574);
nand U3142 (N_3142,In_1088,In_696);
and U3143 (N_3143,In_1439,In_179);
nand U3144 (N_3144,In_993,In_1146);
nand U3145 (N_3145,In_904,In_1169);
nand U3146 (N_3146,In_1481,In_531);
or U3147 (N_3147,In_750,In_1256);
or U3148 (N_3148,In_551,In_66);
xor U3149 (N_3149,In_1350,In_32);
nor U3150 (N_3150,In_1249,In_1006);
nor U3151 (N_3151,In_1176,In_823);
or U3152 (N_3152,In_1416,In_352);
or U3153 (N_3153,In_1148,In_1087);
nand U3154 (N_3154,In_378,In_822);
nand U3155 (N_3155,In_35,In_408);
nor U3156 (N_3156,In_101,In_629);
or U3157 (N_3157,In_285,In_1424);
or U3158 (N_3158,In_1009,In_731);
or U3159 (N_3159,In_1307,In_951);
or U3160 (N_3160,In_429,In_368);
or U3161 (N_3161,In_397,In_797);
nand U3162 (N_3162,In_993,In_530);
and U3163 (N_3163,In_373,In_171);
nor U3164 (N_3164,In_155,In_1143);
xnor U3165 (N_3165,In_326,In_364);
or U3166 (N_3166,In_1444,In_550);
or U3167 (N_3167,In_736,In_116);
nor U3168 (N_3168,In_653,In_228);
or U3169 (N_3169,In_503,In_1320);
nand U3170 (N_3170,In_392,In_1235);
or U3171 (N_3171,In_552,In_1289);
or U3172 (N_3172,In_252,In_1243);
and U3173 (N_3173,In_511,In_15);
nor U3174 (N_3174,In_365,In_228);
and U3175 (N_3175,In_1328,In_1293);
nor U3176 (N_3176,In_946,In_143);
nand U3177 (N_3177,In_616,In_1209);
or U3178 (N_3178,In_1064,In_159);
nand U3179 (N_3179,In_495,In_606);
and U3180 (N_3180,In_735,In_1330);
nand U3181 (N_3181,In_1187,In_1350);
xnor U3182 (N_3182,In_1311,In_1401);
nor U3183 (N_3183,In_32,In_1108);
or U3184 (N_3184,In_487,In_877);
nand U3185 (N_3185,In_1107,In_1073);
and U3186 (N_3186,In_330,In_671);
nor U3187 (N_3187,In_1365,In_856);
nor U3188 (N_3188,In_676,In_219);
nor U3189 (N_3189,In_348,In_77);
xor U3190 (N_3190,In_825,In_221);
or U3191 (N_3191,In_655,In_906);
nand U3192 (N_3192,In_1425,In_267);
nand U3193 (N_3193,In_220,In_433);
nand U3194 (N_3194,In_1322,In_1303);
or U3195 (N_3195,In_1217,In_556);
or U3196 (N_3196,In_698,In_377);
nand U3197 (N_3197,In_1001,In_172);
and U3198 (N_3198,In_862,In_279);
or U3199 (N_3199,In_1230,In_1393);
or U3200 (N_3200,In_1467,In_1189);
nor U3201 (N_3201,In_1051,In_782);
and U3202 (N_3202,In_1481,In_834);
or U3203 (N_3203,In_1067,In_334);
or U3204 (N_3204,In_427,In_1332);
or U3205 (N_3205,In_1407,In_454);
or U3206 (N_3206,In_1101,In_858);
nand U3207 (N_3207,In_1394,In_571);
nand U3208 (N_3208,In_1148,In_1141);
nand U3209 (N_3209,In_437,In_1343);
nand U3210 (N_3210,In_443,In_79);
or U3211 (N_3211,In_36,In_235);
xnor U3212 (N_3212,In_784,In_806);
or U3213 (N_3213,In_467,In_156);
and U3214 (N_3214,In_441,In_1351);
nand U3215 (N_3215,In_405,In_1257);
nand U3216 (N_3216,In_568,In_932);
and U3217 (N_3217,In_1267,In_1221);
and U3218 (N_3218,In_1466,In_1269);
and U3219 (N_3219,In_1433,In_1293);
nand U3220 (N_3220,In_781,In_939);
and U3221 (N_3221,In_277,In_115);
or U3222 (N_3222,In_590,In_1107);
or U3223 (N_3223,In_193,In_1419);
or U3224 (N_3224,In_269,In_768);
xor U3225 (N_3225,In_399,In_1070);
and U3226 (N_3226,In_182,In_977);
nor U3227 (N_3227,In_1054,In_892);
or U3228 (N_3228,In_735,In_791);
and U3229 (N_3229,In_1466,In_136);
and U3230 (N_3230,In_1363,In_1451);
xnor U3231 (N_3231,In_807,In_554);
and U3232 (N_3232,In_9,In_656);
or U3233 (N_3233,In_461,In_313);
or U3234 (N_3234,In_331,In_1264);
nor U3235 (N_3235,In_372,In_838);
and U3236 (N_3236,In_919,In_423);
and U3237 (N_3237,In_804,In_1090);
xor U3238 (N_3238,In_503,In_1366);
nor U3239 (N_3239,In_1479,In_1389);
or U3240 (N_3240,In_759,In_218);
nor U3241 (N_3241,In_919,In_1473);
nand U3242 (N_3242,In_198,In_500);
nor U3243 (N_3243,In_804,In_1178);
and U3244 (N_3244,In_24,In_331);
or U3245 (N_3245,In_990,In_353);
xnor U3246 (N_3246,In_309,In_474);
nand U3247 (N_3247,In_202,In_696);
nand U3248 (N_3248,In_991,In_932);
or U3249 (N_3249,In_190,In_90);
nor U3250 (N_3250,In_1264,In_1231);
nor U3251 (N_3251,In_389,In_273);
nand U3252 (N_3252,In_816,In_1143);
nor U3253 (N_3253,In_397,In_738);
nor U3254 (N_3254,In_609,In_443);
or U3255 (N_3255,In_541,In_772);
nor U3256 (N_3256,In_452,In_734);
nand U3257 (N_3257,In_1189,In_256);
and U3258 (N_3258,In_279,In_735);
nor U3259 (N_3259,In_1044,In_1004);
or U3260 (N_3260,In_513,In_1482);
and U3261 (N_3261,In_14,In_698);
and U3262 (N_3262,In_698,In_576);
nor U3263 (N_3263,In_888,In_304);
nand U3264 (N_3264,In_543,In_23);
nor U3265 (N_3265,In_675,In_1478);
and U3266 (N_3266,In_611,In_374);
and U3267 (N_3267,In_353,In_746);
or U3268 (N_3268,In_1295,In_956);
or U3269 (N_3269,In_125,In_981);
and U3270 (N_3270,In_1004,In_284);
or U3271 (N_3271,In_108,In_1163);
or U3272 (N_3272,In_333,In_1467);
nor U3273 (N_3273,In_1088,In_106);
xor U3274 (N_3274,In_692,In_612);
and U3275 (N_3275,In_571,In_1242);
nand U3276 (N_3276,In_1133,In_642);
xor U3277 (N_3277,In_22,In_619);
or U3278 (N_3278,In_1218,In_344);
xnor U3279 (N_3279,In_223,In_920);
nand U3280 (N_3280,In_620,In_102);
nand U3281 (N_3281,In_1395,In_401);
and U3282 (N_3282,In_1419,In_703);
and U3283 (N_3283,In_183,In_672);
and U3284 (N_3284,In_486,In_1423);
nand U3285 (N_3285,In_134,In_43);
nor U3286 (N_3286,In_1310,In_601);
or U3287 (N_3287,In_514,In_160);
xnor U3288 (N_3288,In_352,In_649);
and U3289 (N_3289,In_1106,In_206);
nand U3290 (N_3290,In_413,In_1011);
nor U3291 (N_3291,In_78,In_1230);
or U3292 (N_3292,In_676,In_166);
and U3293 (N_3293,In_1341,In_251);
and U3294 (N_3294,In_617,In_744);
nor U3295 (N_3295,In_1100,In_87);
and U3296 (N_3296,In_1304,In_430);
and U3297 (N_3297,In_811,In_489);
nand U3298 (N_3298,In_1354,In_1197);
nand U3299 (N_3299,In_697,In_115);
and U3300 (N_3300,In_908,In_1095);
or U3301 (N_3301,In_731,In_792);
and U3302 (N_3302,In_707,In_1481);
nand U3303 (N_3303,In_952,In_293);
or U3304 (N_3304,In_400,In_1305);
and U3305 (N_3305,In_1461,In_1319);
nor U3306 (N_3306,In_56,In_1499);
nand U3307 (N_3307,In_71,In_595);
and U3308 (N_3308,In_911,In_66);
or U3309 (N_3309,In_48,In_216);
or U3310 (N_3310,In_669,In_497);
nor U3311 (N_3311,In_1316,In_613);
or U3312 (N_3312,In_571,In_1472);
or U3313 (N_3313,In_37,In_1008);
nor U3314 (N_3314,In_1058,In_613);
nor U3315 (N_3315,In_1301,In_1396);
xnor U3316 (N_3316,In_383,In_441);
and U3317 (N_3317,In_1320,In_17);
nand U3318 (N_3318,In_911,In_1046);
nand U3319 (N_3319,In_607,In_104);
nor U3320 (N_3320,In_689,In_1099);
nand U3321 (N_3321,In_747,In_1392);
nand U3322 (N_3322,In_1112,In_170);
nor U3323 (N_3323,In_1453,In_638);
and U3324 (N_3324,In_129,In_200);
or U3325 (N_3325,In_1008,In_1360);
nor U3326 (N_3326,In_978,In_629);
nand U3327 (N_3327,In_578,In_652);
nor U3328 (N_3328,In_475,In_1364);
or U3329 (N_3329,In_1278,In_300);
or U3330 (N_3330,In_1025,In_1040);
nor U3331 (N_3331,In_658,In_472);
and U3332 (N_3332,In_1061,In_345);
nand U3333 (N_3333,In_948,In_1258);
xor U3334 (N_3334,In_361,In_1008);
nand U3335 (N_3335,In_1442,In_34);
nor U3336 (N_3336,In_1317,In_530);
nor U3337 (N_3337,In_806,In_1439);
nor U3338 (N_3338,In_1089,In_654);
nand U3339 (N_3339,In_1341,In_378);
and U3340 (N_3340,In_733,In_940);
nor U3341 (N_3341,In_906,In_711);
and U3342 (N_3342,In_774,In_703);
or U3343 (N_3343,In_402,In_1465);
nor U3344 (N_3344,In_1459,In_1);
or U3345 (N_3345,In_1121,In_542);
xnor U3346 (N_3346,In_94,In_1178);
or U3347 (N_3347,In_41,In_1108);
and U3348 (N_3348,In_90,In_441);
nand U3349 (N_3349,In_1111,In_999);
or U3350 (N_3350,In_608,In_920);
xnor U3351 (N_3351,In_1320,In_697);
nand U3352 (N_3352,In_942,In_114);
and U3353 (N_3353,In_1399,In_924);
nor U3354 (N_3354,In_1489,In_339);
nor U3355 (N_3355,In_178,In_1156);
and U3356 (N_3356,In_210,In_422);
or U3357 (N_3357,In_616,In_1437);
or U3358 (N_3358,In_510,In_613);
or U3359 (N_3359,In_63,In_705);
nand U3360 (N_3360,In_1011,In_573);
and U3361 (N_3361,In_339,In_1125);
and U3362 (N_3362,In_321,In_1115);
xor U3363 (N_3363,In_91,In_1208);
and U3364 (N_3364,In_438,In_270);
nand U3365 (N_3365,In_1080,In_549);
nand U3366 (N_3366,In_721,In_867);
or U3367 (N_3367,In_174,In_158);
nand U3368 (N_3368,In_451,In_892);
and U3369 (N_3369,In_226,In_1458);
or U3370 (N_3370,In_1315,In_465);
and U3371 (N_3371,In_99,In_917);
nor U3372 (N_3372,In_163,In_35);
nor U3373 (N_3373,In_673,In_600);
nand U3374 (N_3374,In_23,In_674);
or U3375 (N_3375,In_374,In_1375);
or U3376 (N_3376,In_532,In_721);
or U3377 (N_3377,In_1065,In_1290);
nor U3378 (N_3378,In_1477,In_566);
nand U3379 (N_3379,In_32,In_458);
and U3380 (N_3380,In_363,In_810);
nor U3381 (N_3381,In_964,In_81);
or U3382 (N_3382,In_609,In_549);
or U3383 (N_3383,In_1152,In_1323);
and U3384 (N_3384,In_987,In_159);
and U3385 (N_3385,In_706,In_1060);
nand U3386 (N_3386,In_1158,In_1216);
or U3387 (N_3387,In_479,In_1179);
or U3388 (N_3388,In_984,In_198);
nor U3389 (N_3389,In_1262,In_774);
nand U3390 (N_3390,In_254,In_129);
or U3391 (N_3391,In_1432,In_142);
xnor U3392 (N_3392,In_594,In_422);
xnor U3393 (N_3393,In_766,In_1477);
xnor U3394 (N_3394,In_1062,In_34);
or U3395 (N_3395,In_660,In_705);
nor U3396 (N_3396,In_1075,In_1341);
xnor U3397 (N_3397,In_107,In_472);
or U3398 (N_3398,In_295,In_700);
or U3399 (N_3399,In_1396,In_142);
or U3400 (N_3400,In_149,In_341);
nor U3401 (N_3401,In_447,In_512);
nor U3402 (N_3402,In_937,In_313);
nand U3403 (N_3403,In_1176,In_259);
xnor U3404 (N_3404,In_381,In_1475);
nor U3405 (N_3405,In_1433,In_756);
nand U3406 (N_3406,In_743,In_1029);
nor U3407 (N_3407,In_1291,In_348);
nor U3408 (N_3408,In_117,In_617);
and U3409 (N_3409,In_395,In_1437);
or U3410 (N_3410,In_1332,In_1048);
or U3411 (N_3411,In_376,In_710);
and U3412 (N_3412,In_975,In_1205);
nand U3413 (N_3413,In_949,In_1071);
xor U3414 (N_3414,In_652,In_176);
nor U3415 (N_3415,In_1479,In_1357);
or U3416 (N_3416,In_1184,In_942);
and U3417 (N_3417,In_1357,In_854);
nor U3418 (N_3418,In_1452,In_1044);
xor U3419 (N_3419,In_515,In_1073);
nand U3420 (N_3420,In_289,In_1106);
or U3421 (N_3421,In_651,In_228);
and U3422 (N_3422,In_444,In_1102);
or U3423 (N_3423,In_76,In_369);
nor U3424 (N_3424,In_851,In_383);
and U3425 (N_3425,In_62,In_939);
and U3426 (N_3426,In_1114,In_160);
or U3427 (N_3427,In_1195,In_184);
and U3428 (N_3428,In_416,In_713);
nand U3429 (N_3429,In_986,In_1302);
nand U3430 (N_3430,In_123,In_914);
nand U3431 (N_3431,In_284,In_1433);
nor U3432 (N_3432,In_112,In_293);
and U3433 (N_3433,In_20,In_942);
or U3434 (N_3434,In_1482,In_125);
or U3435 (N_3435,In_575,In_1110);
or U3436 (N_3436,In_834,In_1429);
nor U3437 (N_3437,In_82,In_1021);
nor U3438 (N_3438,In_1416,In_378);
xnor U3439 (N_3439,In_475,In_1151);
xnor U3440 (N_3440,In_1172,In_172);
or U3441 (N_3441,In_821,In_1199);
nor U3442 (N_3442,In_558,In_145);
nor U3443 (N_3443,In_625,In_882);
nand U3444 (N_3444,In_866,In_253);
and U3445 (N_3445,In_127,In_498);
nand U3446 (N_3446,In_562,In_1117);
nand U3447 (N_3447,In_1409,In_194);
nor U3448 (N_3448,In_528,In_114);
xor U3449 (N_3449,In_922,In_287);
and U3450 (N_3450,In_703,In_857);
nor U3451 (N_3451,In_155,In_1196);
nand U3452 (N_3452,In_604,In_769);
or U3453 (N_3453,In_739,In_839);
nor U3454 (N_3454,In_102,In_691);
or U3455 (N_3455,In_368,In_781);
and U3456 (N_3456,In_351,In_396);
and U3457 (N_3457,In_1347,In_900);
and U3458 (N_3458,In_1427,In_1295);
or U3459 (N_3459,In_223,In_699);
or U3460 (N_3460,In_423,In_142);
xor U3461 (N_3461,In_1202,In_807);
nor U3462 (N_3462,In_559,In_236);
and U3463 (N_3463,In_941,In_41);
nand U3464 (N_3464,In_976,In_334);
or U3465 (N_3465,In_573,In_516);
xor U3466 (N_3466,In_1071,In_1099);
and U3467 (N_3467,In_681,In_846);
or U3468 (N_3468,In_395,In_819);
and U3469 (N_3469,In_601,In_8);
xnor U3470 (N_3470,In_540,In_1337);
nand U3471 (N_3471,In_628,In_657);
and U3472 (N_3472,In_356,In_1246);
nand U3473 (N_3473,In_1078,In_525);
nand U3474 (N_3474,In_834,In_450);
nor U3475 (N_3475,In_916,In_714);
and U3476 (N_3476,In_642,In_19);
and U3477 (N_3477,In_931,In_796);
nor U3478 (N_3478,In_77,In_1352);
nor U3479 (N_3479,In_901,In_501);
and U3480 (N_3480,In_44,In_585);
nor U3481 (N_3481,In_1108,In_252);
nand U3482 (N_3482,In_458,In_172);
nand U3483 (N_3483,In_230,In_905);
nor U3484 (N_3484,In_1080,In_256);
or U3485 (N_3485,In_728,In_1404);
nand U3486 (N_3486,In_634,In_844);
and U3487 (N_3487,In_1267,In_976);
and U3488 (N_3488,In_302,In_564);
and U3489 (N_3489,In_347,In_554);
or U3490 (N_3490,In_1447,In_872);
or U3491 (N_3491,In_140,In_897);
or U3492 (N_3492,In_1365,In_1322);
xor U3493 (N_3493,In_543,In_1443);
xnor U3494 (N_3494,In_881,In_843);
or U3495 (N_3495,In_941,In_1364);
nor U3496 (N_3496,In_1007,In_1467);
nand U3497 (N_3497,In_188,In_272);
and U3498 (N_3498,In_675,In_767);
and U3499 (N_3499,In_1357,In_1200);
nor U3500 (N_3500,In_1004,In_1419);
or U3501 (N_3501,In_1292,In_124);
or U3502 (N_3502,In_247,In_570);
and U3503 (N_3503,In_306,In_276);
and U3504 (N_3504,In_100,In_199);
nor U3505 (N_3505,In_1369,In_900);
nand U3506 (N_3506,In_170,In_1458);
or U3507 (N_3507,In_44,In_346);
nand U3508 (N_3508,In_974,In_552);
nand U3509 (N_3509,In_492,In_1477);
nor U3510 (N_3510,In_1116,In_1356);
xor U3511 (N_3511,In_638,In_482);
or U3512 (N_3512,In_456,In_884);
xor U3513 (N_3513,In_1219,In_983);
nor U3514 (N_3514,In_214,In_306);
nor U3515 (N_3515,In_1323,In_1049);
xor U3516 (N_3516,In_990,In_885);
nand U3517 (N_3517,In_509,In_105);
nand U3518 (N_3518,In_454,In_1414);
nand U3519 (N_3519,In_1263,In_170);
or U3520 (N_3520,In_438,In_941);
nor U3521 (N_3521,In_724,In_35);
nand U3522 (N_3522,In_1179,In_256);
or U3523 (N_3523,In_1051,In_315);
or U3524 (N_3524,In_771,In_248);
nand U3525 (N_3525,In_1349,In_820);
nor U3526 (N_3526,In_484,In_8);
nor U3527 (N_3527,In_519,In_1135);
nor U3528 (N_3528,In_55,In_338);
nand U3529 (N_3529,In_1272,In_1200);
and U3530 (N_3530,In_1253,In_562);
or U3531 (N_3531,In_1105,In_392);
or U3532 (N_3532,In_355,In_76);
nand U3533 (N_3533,In_1448,In_1258);
xor U3534 (N_3534,In_758,In_736);
nand U3535 (N_3535,In_604,In_1179);
nand U3536 (N_3536,In_563,In_789);
and U3537 (N_3537,In_255,In_371);
or U3538 (N_3538,In_303,In_796);
and U3539 (N_3539,In_1399,In_1421);
nand U3540 (N_3540,In_394,In_878);
nand U3541 (N_3541,In_867,In_1287);
or U3542 (N_3542,In_260,In_869);
nand U3543 (N_3543,In_969,In_1178);
nand U3544 (N_3544,In_201,In_1325);
nand U3545 (N_3545,In_369,In_102);
nor U3546 (N_3546,In_1046,In_1205);
nand U3547 (N_3547,In_1180,In_586);
nand U3548 (N_3548,In_162,In_1009);
and U3549 (N_3549,In_435,In_1454);
or U3550 (N_3550,In_1258,In_751);
and U3551 (N_3551,In_1307,In_692);
and U3552 (N_3552,In_30,In_1322);
nor U3553 (N_3553,In_1355,In_1000);
nand U3554 (N_3554,In_459,In_486);
or U3555 (N_3555,In_495,In_181);
and U3556 (N_3556,In_523,In_1083);
nor U3557 (N_3557,In_129,In_1044);
or U3558 (N_3558,In_853,In_469);
or U3559 (N_3559,In_687,In_901);
and U3560 (N_3560,In_908,In_941);
nor U3561 (N_3561,In_509,In_1018);
nor U3562 (N_3562,In_78,In_418);
nand U3563 (N_3563,In_1365,In_648);
nand U3564 (N_3564,In_979,In_229);
and U3565 (N_3565,In_112,In_1292);
nand U3566 (N_3566,In_1455,In_1026);
or U3567 (N_3567,In_871,In_143);
or U3568 (N_3568,In_1174,In_1251);
and U3569 (N_3569,In_1414,In_1153);
nand U3570 (N_3570,In_868,In_928);
nor U3571 (N_3571,In_1299,In_1033);
or U3572 (N_3572,In_1312,In_320);
and U3573 (N_3573,In_1461,In_130);
xnor U3574 (N_3574,In_1467,In_916);
nor U3575 (N_3575,In_276,In_692);
nor U3576 (N_3576,In_549,In_479);
nor U3577 (N_3577,In_821,In_333);
or U3578 (N_3578,In_41,In_728);
and U3579 (N_3579,In_198,In_235);
and U3580 (N_3580,In_997,In_688);
and U3581 (N_3581,In_7,In_1365);
nor U3582 (N_3582,In_566,In_846);
nand U3583 (N_3583,In_1020,In_477);
or U3584 (N_3584,In_102,In_694);
xnor U3585 (N_3585,In_401,In_1453);
and U3586 (N_3586,In_992,In_1375);
or U3587 (N_3587,In_273,In_1165);
nor U3588 (N_3588,In_595,In_166);
or U3589 (N_3589,In_413,In_848);
nand U3590 (N_3590,In_653,In_106);
nand U3591 (N_3591,In_1002,In_314);
nand U3592 (N_3592,In_1087,In_390);
or U3593 (N_3593,In_185,In_455);
and U3594 (N_3594,In_1330,In_1199);
nor U3595 (N_3595,In_938,In_1499);
or U3596 (N_3596,In_344,In_387);
nor U3597 (N_3597,In_1322,In_182);
and U3598 (N_3598,In_965,In_111);
nor U3599 (N_3599,In_303,In_1465);
or U3600 (N_3600,In_657,In_111);
and U3601 (N_3601,In_844,In_157);
nor U3602 (N_3602,In_1078,In_342);
or U3603 (N_3603,In_1356,In_1287);
and U3604 (N_3604,In_677,In_648);
or U3605 (N_3605,In_106,In_218);
or U3606 (N_3606,In_882,In_418);
and U3607 (N_3607,In_1281,In_455);
nand U3608 (N_3608,In_97,In_1416);
xnor U3609 (N_3609,In_380,In_427);
nand U3610 (N_3610,In_726,In_850);
and U3611 (N_3611,In_1193,In_730);
nor U3612 (N_3612,In_598,In_1448);
or U3613 (N_3613,In_3,In_728);
and U3614 (N_3614,In_623,In_701);
nor U3615 (N_3615,In_898,In_271);
or U3616 (N_3616,In_796,In_240);
or U3617 (N_3617,In_1264,In_236);
and U3618 (N_3618,In_960,In_764);
and U3619 (N_3619,In_1446,In_1103);
and U3620 (N_3620,In_349,In_705);
or U3621 (N_3621,In_84,In_882);
and U3622 (N_3622,In_790,In_494);
xnor U3623 (N_3623,In_222,In_115);
nor U3624 (N_3624,In_937,In_585);
xor U3625 (N_3625,In_1380,In_1263);
xnor U3626 (N_3626,In_1258,In_771);
nand U3627 (N_3627,In_1426,In_470);
nand U3628 (N_3628,In_393,In_746);
or U3629 (N_3629,In_1106,In_1159);
and U3630 (N_3630,In_375,In_52);
nand U3631 (N_3631,In_985,In_352);
nor U3632 (N_3632,In_350,In_460);
or U3633 (N_3633,In_550,In_118);
or U3634 (N_3634,In_922,In_403);
nor U3635 (N_3635,In_991,In_561);
nand U3636 (N_3636,In_942,In_62);
and U3637 (N_3637,In_656,In_313);
xor U3638 (N_3638,In_13,In_902);
nor U3639 (N_3639,In_727,In_184);
nand U3640 (N_3640,In_392,In_1317);
or U3641 (N_3641,In_276,In_237);
xor U3642 (N_3642,In_1432,In_1117);
or U3643 (N_3643,In_387,In_99);
xnor U3644 (N_3644,In_750,In_253);
or U3645 (N_3645,In_434,In_758);
nand U3646 (N_3646,In_1030,In_769);
nand U3647 (N_3647,In_550,In_159);
nor U3648 (N_3648,In_1452,In_485);
nor U3649 (N_3649,In_1063,In_598);
or U3650 (N_3650,In_1464,In_727);
nor U3651 (N_3651,In_674,In_545);
and U3652 (N_3652,In_845,In_744);
nor U3653 (N_3653,In_550,In_143);
nand U3654 (N_3654,In_516,In_396);
and U3655 (N_3655,In_565,In_89);
nor U3656 (N_3656,In_910,In_794);
and U3657 (N_3657,In_423,In_651);
nor U3658 (N_3658,In_104,In_25);
nand U3659 (N_3659,In_414,In_993);
nor U3660 (N_3660,In_397,In_216);
and U3661 (N_3661,In_672,In_1164);
and U3662 (N_3662,In_810,In_313);
nor U3663 (N_3663,In_489,In_124);
and U3664 (N_3664,In_1477,In_1490);
and U3665 (N_3665,In_1312,In_1316);
nor U3666 (N_3666,In_258,In_1294);
or U3667 (N_3667,In_1450,In_782);
nand U3668 (N_3668,In_866,In_363);
or U3669 (N_3669,In_923,In_1137);
and U3670 (N_3670,In_585,In_889);
nand U3671 (N_3671,In_1277,In_643);
nand U3672 (N_3672,In_915,In_309);
or U3673 (N_3673,In_476,In_157);
nand U3674 (N_3674,In_219,In_35);
and U3675 (N_3675,In_462,In_530);
nor U3676 (N_3676,In_170,In_734);
nor U3677 (N_3677,In_1310,In_1225);
nand U3678 (N_3678,In_1158,In_301);
or U3679 (N_3679,In_934,In_946);
or U3680 (N_3680,In_1336,In_601);
and U3681 (N_3681,In_1291,In_1115);
nor U3682 (N_3682,In_1085,In_642);
and U3683 (N_3683,In_1102,In_406);
or U3684 (N_3684,In_382,In_647);
nand U3685 (N_3685,In_1487,In_44);
nand U3686 (N_3686,In_1077,In_77);
nand U3687 (N_3687,In_869,In_1030);
nand U3688 (N_3688,In_1212,In_1302);
xnor U3689 (N_3689,In_726,In_1223);
and U3690 (N_3690,In_1143,In_1321);
and U3691 (N_3691,In_134,In_555);
nand U3692 (N_3692,In_1448,In_1474);
xor U3693 (N_3693,In_1221,In_940);
and U3694 (N_3694,In_22,In_144);
and U3695 (N_3695,In_300,In_86);
nand U3696 (N_3696,In_692,In_874);
nand U3697 (N_3697,In_246,In_1039);
nor U3698 (N_3698,In_1028,In_78);
and U3699 (N_3699,In_1424,In_1478);
nand U3700 (N_3700,In_572,In_847);
and U3701 (N_3701,In_837,In_1225);
or U3702 (N_3702,In_338,In_1481);
xor U3703 (N_3703,In_1346,In_201);
and U3704 (N_3704,In_984,In_1041);
nand U3705 (N_3705,In_131,In_1268);
nor U3706 (N_3706,In_1050,In_179);
nor U3707 (N_3707,In_917,In_591);
nor U3708 (N_3708,In_450,In_1057);
and U3709 (N_3709,In_1278,In_509);
or U3710 (N_3710,In_562,In_96);
nand U3711 (N_3711,In_209,In_901);
xnor U3712 (N_3712,In_1234,In_1140);
nand U3713 (N_3713,In_436,In_949);
nand U3714 (N_3714,In_994,In_1142);
or U3715 (N_3715,In_926,In_1273);
nand U3716 (N_3716,In_231,In_1035);
nor U3717 (N_3717,In_140,In_741);
or U3718 (N_3718,In_328,In_994);
and U3719 (N_3719,In_1441,In_746);
or U3720 (N_3720,In_626,In_1129);
nor U3721 (N_3721,In_931,In_902);
or U3722 (N_3722,In_1176,In_348);
xor U3723 (N_3723,In_799,In_680);
nor U3724 (N_3724,In_1076,In_338);
and U3725 (N_3725,In_269,In_730);
nor U3726 (N_3726,In_1200,In_1334);
or U3727 (N_3727,In_219,In_1222);
and U3728 (N_3728,In_564,In_379);
nand U3729 (N_3729,In_353,In_760);
nor U3730 (N_3730,In_1025,In_1180);
and U3731 (N_3731,In_375,In_598);
and U3732 (N_3732,In_415,In_908);
nand U3733 (N_3733,In_1272,In_1042);
nor U3734 (N_3734,In_1248,In_1416);
nand U3735 (N_3735,In_768,In_1254);
nand U3736 (N_3736,In_910,In_994);
or U3737 (N_3737,In_1140,In_397);
nor U3738 (N_3738,In_159,In_607);
and U3739 (N_3739,In_556,In_852);
or U3740 (N_3740,In_1226,In_1087);
nand U3741 (N_3741,In_413,In_749);
and U3742 (N_3742,In_1411,In_1406);
nor U3743 (N_3743,In_460,In_621);
xnor U3744 (N_3744,In_643,In_765);
or U3745 (N_3745,In_433,In_48);
nor U3746 (N_3746,In_60,In_402);
nand U3747 (N_3747,In_442,In_434);
nand U3748 (N_3748,In_74,In_48);
or U3749 (N_3749,In_946,In_1295);
or U3750 (N_3750,In_315,In_1010);
nand U3751 (N_3751,In_1085,In_1261);
or U3752 (N_3752,In_1264,In_365);
or U3753 (N_3753,In_579,In_1348);
nand U3754 (N_3754,In_1080,In_596);
or U3755 (N_3755,In_1290,In_898);
nand U3756 (N_3756,In_1446,In_539);
nand U3757 (N_3757,In_648,In_816);
nor U3758 (N_3758,In_127,In_731);
or U3759 (N_3759,In_1049,In_295);
nand U3760 (N_3760,In_1206,In_861);
nand U3761 (N_3761,In_815,In_1392);
xnor U3762 (N_3762,In_470,In_259);
and U3763 (N_3763,In_1207,In_1445);
and U3764 (N_3764,In_1257,In_1039);
or U3765 (N_3765,In_657,In_557);
or U3766 (N_3766,In_1076,In_1157);
nand U3767 (N_3767,In_1107,In_1317);
nand U3768 (N_3768,In_1166,In_957);
and U3769 (N_3769,In_777,In_599);
nor U3770 (N_3770,In_516,In_1270);
or U3771 (N_3771,In_41,In_6);
and U3772 (N_3772,In_64,In_235);
and U3773 (N_3773,In_589,In_491);
nor U3774 (N_3774,In_1461,In_1120);
nor U3775 (N_3775,In_928,In_58);
nor U3776 (N_3776,In_505,In_980);
and U3777 (N_3777,In_126,In_926);
or U3778 (N_3778,In_160,In_309);
and U3779 (N_3779,In_997,In_365);
nand U3780 (N_3780,In_1161,In_1006);
nor U3781 (N_3781,In_673,In_1184);
or U3782 (N_3782,In_1460,In_540);
xor U3783 (N_3783,In_927,In_53);
xnor U3784 (N_3784,In_1198,In_1155);
and U3785 (N_3785,In_710,In_294);
or U3786 (N_3786,In_80,In_995);
xor U3787 (N_3787,In_204,In_1223);
or U3788 (N_3788,In_1119,In_1031);
nand U3789 (N_3789,In_1403,In_647);
or U3790 (N_3790,In_466,In_323);
nand U3791 (N_3791,In_189,In_301);
or U3792 (N_3792,In_402,In_460);
or U3793 (N_3793,In_1029,In_863);
nor U3794 (N_3794,In_681,In_274);
nand U3795 (N_3795,In_227,In_710);
or U3796 (N_3796,In_691,In_1492);
and U3797 (N_3797,In_980,In_325);
or U3798 (N_3798,In_996,In_1065);
nor U3799 (N_3799,In_1219,In_798);
xnor U3800 (N_3800,In_118,In_1189);
and U3801 (N_3801,In_899,In_594);
nand U3802 (N_3802,In_296,In_588);
nor U3803 (N_3803,In_1133,In_1013);
nor U3804 (N_3804,In_463,In_133);
and U3805 (N_3805,In_352,In_1360);
and U3806 (N_3806,In_24,In_419);
and U3807 (N_3807,In_977,In_851);
or U3808 (N_3808,In_398,In_1412);
nand U3809 (N_3809,In_1009,In_1473);
or U3810 (N_3810,In_1247,In_1418);
nand U3811 (N_3811,In_308,In_1389);
nor U3812 (N_3812,In_1448,In_1249);
and U3813 (N_3813,In_459,In_1098);
or U3814 (N_3814,In_753,In_500);
nand U3815 (N_3815,In_1188,In_1114);
nor U3816 (N_3816,In_946,In_1001);
and U3817 (N_3817,In_382,In_464);
nor U3818 (N_3818,In_915,In_658);
or U3819 (N_3819,In_502,In_682);
nand U3820 (N_3820,In_1489,In_627);
or U3821 (N_3821,In_911,In_148);
or U3822 (N_3822,In_797,In_816);
and U3823 (N_3823,In_1035,In_753);
nand U3824 (N_3824,In_1452,In_1162);
or U3825 (N_3825,In_831,In_595);
and U3826 (N_3826,In_963,In_368);
nand U3827 (N_3827,In_343,In_486);
and U3828 (N_3828,In_854,In_702);
and U3829 (N_3829,In_1450,In_1413);
or U3830 (N_3830,In_591,In_810);
xnor U3831 (N_3831,In_34,In_1235);
nand U3832 (N_3832,In_826,In_704);
nand U3833 (N_3833,In_9,In_1307);
and U3834 (N_3834,In_1403,In_121);
and U3835 (N_3835,In_115,In_124);
nor U3836 (N_3836,In_970,In_1336);
or U3837 (N_3837,In_497,In_300);
or U3838 (N_3838,In_912,In_22);
xnor U3839 (N_3839,In_1384,In_64);
and U3840 (N_3840,In_877,In_581);
nor U3841 (N_3841,In_1398,In_357);
or U3842 (N_3842,In_686,In_1187);
nor U3843 (N_3843,In_29,In_1429);
or U3844 (N_3844,In_474,In_284);
nor U3845 (N_3845,In_239,In_687);
nor U3846 (N_3846,In_12,In_1493);
nor U3847 (N_3847,In_4,In_947);
or U3848 (N_3848,In_825,In_1364);
xnor U3849 (N_3849,In_276,In_294);
nand U3850 (N_3850,In_1297,In_1378);
or U3851 (N_3851,In_968,In_761);
nand U3852 (N_3852,In_996,In_873);
or U3853 (N_3853,In_950,In_855);
nor U3854 (N_3854,In_1197,In_1332);
and U3855 (N_3855,In_858,In_1367);
and U3856 (N_3856,In_935,In_1480);
nand U3857 (N_3857,In_253,In_587);
xnor U3858 (N_3858,In_350,In_1162);
nand U3859 (N_3859,In_94,In_1421);
and U3860 (N_3860,In_1202,In_1064);
nor U3861 (N_3861,In_851,In_1447);
xor U3862 (N_3862,In_1163,In_724);
nor U3863 (N_3863,In_803,In_302);
nand U3864 (N_3864,In_1295,In_1243);
or U3865 (N_3865,In_781,In_1137);
nand U3866 (N_3866,In_319,In_712);
and U3867 (N_3867,In_576,In_133);
nor U3868 (N_3868,In_602,In_1216);
nand U3869 (N_3869,In_8,In_1378);
and U3870 (N_3870,In_966,In_979);
and U3871 (N_3871,In_1024,In_23);
nand U3872 (N_3872,In_149,In_757);
and U3873 (N_3873,In_1070,In_1196);
and U3874 (N_3874,In_906,In_608);
and U3875 (N_3875,In_755,In_912);
or U3876 (N_3876,In_1174,In_539);
or U3877 (N_3877,In_754,In_250);
or U3878 (N_3878,In_1176,In_250);
nand U3879 (N_3879,In_350,In_853);
or U3880 (N_3880,In_95,In_125);
and U3881 (N_3881,In_391,In_1230);
nor U3882 (N_3882,In_1340,In_164);
nor U3883 (N_3883,In_615,In_1189);
nand U3884 (N_3884,In_935,In_88);
nor U3885 (N_3885,In_1050,In_418);
or U3886 (N_3886,In_847,In_457);
nand U3887 (N_3887,In_1386,In_1037);
nor U3888 (N_3888,In_1109,In_800);
or U3889 (N_3889,In_698,In_251);
or U3890 (N_3890,In_142,In_18);
or U3891 (N_3891,In_1023,In_73);
xnor U3892 (N_3892,In_511,In_154);
and U3893 (N_3893,In_1025,In_1458);
and U3894 (N_3894,In_431,In_557);
and U3895 (N_3895,In_729,In_676);
or U3896 (N_3896,In_594,In_652);
nor U3897 (N_3897,In_1483,In_1287);
xor U3898 (N_3898,In_707,In_171);
nor U3899 (N_3899,In_523,In_83);
or U3900 (N_3900,In_451,In_362);
or U3901 (N_3901,In_544,In_587);
nand U3902 (N_3902,In_207,In_94);
nand U3903 (N_3903,In_708,In_301);
nor U3904 (N_3904,In_628,In_791);
and U3905 (N_3905,In_234,In_1238);
or U3906 (N_3906,In_287,In_458);
nand U3907 (N_3907,In_997,In_1108);
nand U3908 (N_3908,In_925,In_253);
or U3909 (N_3909,In_718,In_1419);
and U3910 (N_3910,In_1218,In_923);
and U3911 (N_3911,In_91,In_1246);
and U3912 (N_3912,In_483,In_758);
nor U3913 (N_3913,In_831,In_523);
nand U3914 (N_3914,In_1351,In_342);
and U3915 (N_3915,In_197,In_715);
and U3916 (N_3916,In_685,In_257);
nand U3917 (N_3917,In_1266,In_370);
nor U3918 (N_3918,In_1202,In_1494);
and U3919 (N_3919,In_1234,In_1274);
nor U3920 (N_3920,In_904,In_941);
nand U3921 (N_3921,In_1295,In_544);
nor U3922 (N_3922,In_1136,In_1434);
nor U3923 (N_3923,In_2,In_463);
and U3924 (N_3924,In_566,In_353);
xor U3925 (N_3925,In_1184,In_1028);
nand U3926 (N_3926,In_443,In_1028);
nor U3927 (N_3927,In_186,In_666);
nor U3928 (N_3928,In_953,In_629);
xor U3929 (N_3929,In_778,In_905);
nand U3930 (N_3930,In_564,In_1013);
nand U3931 (N_3931,In_573,In_527);
xor U3932 (N_3932,In_1287,In_879);
and U3933 (N_3933,In_311,In_1444);
and U3934 (N_3934,In_148,In_1079);
xnor U3935 (N_3935,In_976,In_1046);
or U3936 (N_3936,In_260,In_772);
nor U3937 (N_3937,In_940,In_558);
or U3938 (N_3938,In_632,In_723);
or U3939 (N_3939,In_1328,In_1205);
nand U3940 (N_3940,In_1185,In_749);
nor U3941 (N_3941,In_1474,In_615);
nand U3942 (N_3942,In_1050,In_72);
nand U3943 (N_3943,In_1311,In_1233);
and U3944 (N_3944,In_177,In_284);
and U3945 (N_3945,In_801,In_1465);
nor U3946 (N_3946,In_1424,In_1002);
xor U3947 (N_3947,In_804,In_1474);
nand U3948 (N_3948,In_1014,In_716);
nor U3949 (N_3949,In_965,In_1423);
nand U3950 (N_3950,In_830,In_790);
nor U3951 (N_3951,In_3,In_1374);
nand U3952 (N_3952,In_443,In_1375);
nor U3953 (N_3953,In_461,In_155);
nand U3954 (N_3954,In_1088,In_760);
or U3955 (N_3955,In_1093,In_618);
nor U3956 (N_3956,In_1331,In_675);
nor U3957 (N_3957,In_1377,In_303);
nor U3958 (N_3958,In_1319,In_910);
and U3959 (N_3959,In_391,In_122);
nor U3960 (N_3960,In_271,In_1468);
or U3961 (N_3961,In_884,In_123);
and U3962 (N_3962,In_318,In_447);
and U3963 (N_3963,In_47,In_1412);
and U3964 (N_3964,In_1024,In_592);
and U3965 (N_3965,In_940,In_1205);
nor U3966 (N_3966,In_9,In_861);
or U3967 (N_3967,In_1120,In_463);
and U3968 (N_3968,In_59,In_4);
nand U3969 (N_3969,In_252,In_1377);
nor U3970 (N_3970,In_771,In_1454);
nor U3971 (N_3971,In_739,In_783);
xor U3972 (N_3972,In_1323,In_298);
nor U3973 (N_3973,In_878,In_858);
and U3974 (N_3974,In_479,In_1127);
and U3975 (N_3975,In_1071,In_501);
nor U3976 (N_3976,In_1418,In_1269);
or U3977 (N_3977,In_98,In_1290);
nor U3978 (N_3978,In_959,In_395);
and U3979 (N_3979,In_765,In_1389);
nand U3980 (N_3980,In_318,In_62);
and U3981 (N_3981,In_779,In_867);
or U3982 (N_3982,In_15,In_1115);
nor U3983 (N_3983,In_1290,In_130);
xor U3984 (N_3984,In_1241,In_320);
and U3985 (N_3985,In_935,In_422);
nor U3986 (N_3986,In_62,In_1373);
or U3987 (N_3987,In_1347,In_348);
and U3988 (N_3988,In_11,In_898);
nand U3989 (N_3989,In_892,In_251);
or U3990 (N_3990,In_132,In_35);
or U3991 (N_3991,In_373,In_1078);
or U3992 (N_3992,In_1169,In_1354);
or U3993 (N_3993,In_1409,In_588);
nor U3994 (N_3994,In_121,In_583);
or U3995 (N_3995,In_22,In_646);
nand U3996 (N_3996,In_992,In_576);
nand U3997 (N_3997,In_1157,In_306);
nor U3998 (N_3998,In_1097,In_810);
and U3999 (N_3999,In_861,In_883);
or U4000 (N_4000,In_1156,In_891);
xnor U4001 (N_4001,In_870,In_317);
nor U4002 (N_4002,In_996,In_855);
nor U4003 (N_4003,In_462,In_880);
nor U4004 (N_4004,In_1449,In_814);
and U4005 (N_4005,In_104,In_908);
nor U4006 (N_4006,In_1427,In_59);
or U4007 (N_4007,In_573,In_213);
and U4008 (N_4008,In_986,In_794);
xor U4009 (N_4009,In_527,In_5);
nand U4010 (N_4010,In_595,In_109);
nor U4011 (N_4011,In_808,In_909);
or U4012 (N_4012,In_1005,In_864);
and U4013 (N_4013,In_148,In_164);
nor U4014 (N_4014,In_785,In_919);
or U4015 (N_4015,In_1351,In_12);
nor U4016 (N_4016,In_1105,In_764);
and U4017 (N_4017,In_1187,In_897);
nor U4018 (N_4018,In_554,In_1460);
or U4019 (N_4019,In_653,In_782);
or U4020 (N_4020,In_1342,In_381);
and U4021 (N_4021,In_21,In_1065);
and U4022 (N_4022,In_256,In_983);
and U4023 (N_4023,In_594,In_1331);
and U4024 (N_4024,In_353,In_174);
or U4025 (N_4025,In_849,In_894);
or U4026 (N_4026,In_1249,In_1070);
nand U4027 (N_4027,In_327,In_1455);
nor U4028 (N_4028,In_1291,In_1129);
nor U4029 (N_4029,In_760,In_59);
nor U4030 (N_4030,In_427,In_940);
and U4031 (N_4031,In_1036,In_1499);
nand U4032 (N_4032,In_288,In_1440);
or U4033 (N_4033,In_1294,In_1);
and U4034 (N_4034,In_1203,In_1208);
nand U4035 (N_4035,In_1048,In_749);
and U4036 (N_4036,In_432,In_1408);
nand U4037 (N_4037,In_247,In_1247);
nand U4038 (N_4038,In_1348,In_1330);
or U4039 (N_4039,In_797,In_606);
nor U4040 (N_4040,In_760,In_414);
nor U4041 (N_4041,In_1130,In_910);
nand U4042 (N_4042,In_832,In_707);
nand U4043 (N_4043,In_896,In_1452);
nand U4044 (N_4044,In_1138,In_1362);
nand U4045 (N_4045,In_246,In_1379);
and U4046 (N_4046,In_377,In_368);
xor U4047 (N_4047,In_740,In_110);
nor U4048 (N_4048,In_403,In_1105);
nor U4049 (N_4049,In_386,In_198);
nor U4050 (N_4050,In_318,In_927);
nand U4051 (N_4051,In_352,In_211);
nor U4052 (N_4052,In_557,In_948);
and U4053 (N_4053,In_1354,In_1048);
or U4054 (N_4054,In_615,In_1070);
and U4055 (N_4055,In_1332,In_971);
nand U4056 (N_4056,In_1341,In_667);
and U4057 (N_4057,In_24,In_210);
nand U4058 (N_4058,In_1443,In_1082);
and U4059 (N_4059,In_854,In_539);
or U4060 (N_4060,In_837,In_1019);
and U4061 (N_4061,In_303,In_1418);
and U4062 (N_4062,In_622,In_487);
nor U4063 (N_4063,In_965,In_12);
xor U4064 (N_4064,In_579,In_270);
xnor U4065 (N_4065,In_1164,In_851);
and U4066 (N_4066,In_1466,In_535);
nand U4067 (N_4067,In_397,In_1161);
xor U4068 (N_4068,In_1318,In_734);
or U4069 (N_4069,In_1464,In_1006);
nand U4070 (N_4070,In_356,In_1118);
nor U4071 (N_4071,In_648,In_1130);
nand U4072 (N_4072,In_1173,In_368);
and U4073 (N_4073,In_1097,In_1009);
nor U4074 (N_4074,In_697,In_620);
nand U4075 (N_4075,In_1399,In_1368);
or U4076 (N_4076,In_1366,In_1249);
or U4077 (N_4077,In_206,In_1497);
xor U4078 (N_4078,In_28,In_1123);
and U4079 (N_4079,In_1277,In_296);
and U4080 (N_4080,In_432,In_966);
or U4081 (N_4081,In_995,In_906);
xor U4082 (N_4082,In_1422,In_469);
xor U4083 (N_4083,In_65,In_624);
nand U4084 (N_4084,In_303,In_161);
or U4085 (N_4085,In_409,In_803);
or U4086 (N_4086,In_877,In_534);
nand U4087 (N_4087,In_357,In_239);
nor U4088 (N_4088,In_1265,In_454);
nand U4089 (N_4089,In_1371,In_427);
and U4090 (N_4090,In_740,In_1472);
nor U4091 (N_4091,In_36,In_1283);
or U4092 (N_4092,In_730,In_1005);
and U4093 (N_4093,In_130,In_524);
and U4094 (N_4094,In_437,In_727);
nand U4095 (N_4095,In_60,In_694);
and U4096 (N_4096,In_790,In_847);
and U4097 (N_4097,In_1038,In_1228);
or U4098 (N_4098,In_1491,In_322);
or U4099 (N_4099,In_1336,In_1265);
or U4100 (N_4100,In_576,In_427);
nor U4101 (N_4101,In_1022,In_973);
nor U4102 (N_4102,In_381,In_508);
and U4103 (N_4103,In_102,In_1206);
xor U4104 (N_4104,In_629,In_541);
or U4105 (N_4105,In_501,In_1390);
or U4106 (N_4106,In_381,In_289);
nand U4107 (N_4107,In_1009,In_1259);
nor U4108 (N_4108,In_1354,In_859);
nor U4109 (N_4109,In_226,In_37);
nor U4110 (N_4110,In_642,In_478);
xnor U4111 (N_4111,In_4,In_215);
xor U4112 (N_4112,In_285,In_342);
xor U4113 (N_4113,In_65,In_95);
and U4114 (N_4114,In_354,In_917);
or U4115 (N_4115,In_403,In_1492);
nand U4116 (N_4116,In_814,In_884);
and U4117 (N_4117,In_254,In_550);
and U4118 (N_4118,In_267,In_853);
or U4119 (N_4119,In_860,In_146);
or U4120 (N_4120,In_744,In_584);
xor U4121 (N_4121,In_1290,In_871);
or U4122 (N_4122,In_1337,In_1380);
or U4123 (N_4123,In_372,In_477);
xnor U4124 (N_4124,In_944,In_588);
and U4125 (N_4125,In_697,In_405);
or U4126 (N_4126,In_583,In_1232);
and U4127 (N_4127,In_792,In_209);
and U4128 (N_4128,In_747,In_170);
nand U4129 (N_4129,In_285,In_564);
nor U4130 (N_4130,In_589,In_237);
nand U4131 (N_4131,In_875,In_813);
xnor U4132 (N_4132,In_720,In_1036);
nor U4133 (N_4133,In_463,In_982);
nand U4134 (N_4134,In_979,In_618);
or U4135 (N_4135,In_1393,In_860);
nand U4136 (N_4136,In_1189,In_1472);
nor U4137 (N_4137,In_1428,In_1181);
nor U4138 (N_4138,In_1229,In_920);
and U4139 (N_4139,In_1453,In_707);
nand U4140 (N_4140,In_583,In_127);
xor U4141 (N_4141,In_798,In_372);
xor U4142 (N_4142,In_92,In_753);
nor U4143 (N_4143,In_48,In_1356);
nor U4144 (N_4144,In_737,In_425);
or U4145 (N_4145,In_342,In_161);
and U4146 (N_4146,In_993,In_66);
nor U4147 (N_4147,In_621,In_1454);
nor U4148 (N_4148,In_382,In_1489);
xnor U4149 (N_4149,In_1437,In_1235);
nor U4150 (N_4150,In_436,In_1151);
nor U4151 (N_4151,In_1155,In_483);
and U4152 (N_4152,In_297,In_511);
nor U4153 (N_4153,In_562,In_1103);
or U4154 (N_4154,In_979,In_865);
nand U4155 (N_4155,In_278,In_498);
and U4156 (N_4156,In_1232,In_1016);
nor U4157 (N_4157,In_12,In_1445);
or U4158 (N_4158,In_1328,In_302);
nand U4159 (N_4159,In_465,In_1179);
nand U4160 (N_4160,In_652,In_733);
xor U4161 (N_4161,In_872,In_1383);
and U4162 (N_4162,In_800,In_701);
nand U4163 (N_4163,In_237,In_1192);
nor U4164 (N_4164,In_1226,In_1365);
or U4165 (N_4165,In_531,In_424);
nor U4166 (N_4166,In_907,In_435);
or U4167 (N_4167,In_332,In_371);
or U4168 (N_4168,In_906,In_468);
nor U4169 (N_4169,In_76,In_62);
nor U4170 (N_4170,In_1121,In_71);
nand U4171 (N_4171,In_183,In_1092);
nand U4172 (N_4172,In_87,In_741);
or U4173 (N_4173,In_1175,In_165);
xor U4174 (N_4174,In_339,In_1029);
and U4175 (N_4175,In_213,In_636);
and U4176 (N_4176,In_673,In_23);
xor U4177 (N_4177,In_991,In_374);
nor U4178 (N_4178,In_944,In_1409);
or U4179 (N_4179,In_1450,In_548);
and U4180 (N_4180,In_447,In_1199);
and U4181 (N_4181,In_755,In_1036);
and U4182 (N_4182,In_1135,In_294);
nor U4183 (N_4183,In_291,In_1268);
nand U4184 (N_4184,In_652,In_1268);
nor U4185 (N_4185,In_691,In_370);
or U4186 (N_4186,In_1092,In_964);
and U4187 (N_4187,In_563,In_1451);
nor U4188 (N_4188,In_867,In_726);
xnor U4189 (N_4189,In_1281,In_909);
or U4190 (N_4190,In_424,In_678);
nand U4191 (N_4191,In_418,In_273);
or U4192 (N_4192,In_188,In_268);
nor U4193 (N_4193,In_921,In_662);
nor U4194 (N_4194,In_531,In_593);
or U4195 (N_4195,In_129,In_1387);
or U4196 (N_4196,In_424,In_526);
nor U4197 (N_4197,In_1331,In_1133);
and U4198 (N_4198,In_1255,In_335);
or U4199 (N_4199,In_1130,In_1313);
and U4200 (N_4200,In_1377,In_68);
nor U4201 (N_4201,In_1349,In_462);
and U4202 (N_4202,In_649,In_1314);
nor U4203 (N_4203,In_1065,In_1380);
and U4204 (N_4204,In_1060,In_39);
and U4205 (N_4205,In_870,In_176);
or U4206 (N_4206,In_617,In_244);
nor U4207 (N_4207,In_1269,In_1077);
nand U4208 (N_4208,In_1394,In_158);
or U4209 (N_4209,In_912,In_572);
nor U4210 (N_4210,In_199,In_1424);
xnor U4211 (N_4211,In_567,In_850);
and U4212 (N_4212,In_3,In_231);
nor U4213 (N_4213,In_1299,In_262);
nand U4214 (N_4214,In_1200,In_1395);
or U4215 (N_4215,In_1217,In_890);
nand U4216 (N_4216,In_1183,In_327);
nand U4217 (N_4217,In_964,In_1366);
and U4218 (N_4218,In_146,In_598);
nor U4219 (N_4219,In_1482,In_1465);
and U4220 (N_4220,In_669,In_447);
nor U4221 (N_4221,In_888,In_771);
and U4222 (N_4222,In_1085,In_1301);
nand U4223 (N_4223,In_1278,In_1019);
or U4224 (N_4224,In_1078,In_969);
and U4225 (N_4225,In_1492,In_69);
nor U4226 (N_4226,In_849,In_734);
xnor U4227 (N_4227,In_1162,In_1070);
xnor U4228 (N_4228,In_1214,In_1302);
nor U4229 (N_4229,In_822,In_1479);
nand U4230 (N_4230,In_803,In_774);
nor U4231 (N_4231,In_1071,In_1349);
and U4232 (N_4232,In_893,In_1017);
nor U4233 (N_4233,In_1416,In_224);
or U4234 (N_4234,In_649,In_69);
nand U4235 (N_4235,In_1302,In_1174);
nor U4236 (N_4236,In_315,In_117);
nand U4237 (N_4237,In_272,In_194);
xnor U4238 (N_4238,In_1245,In_1033);
and U4239 (N_4239,In_139,In_107);
or U4240 (N_4240,In_699,In_1476);
nor U4241 (N_4241,In_1235,In_1039);
nor U4242 (N_4242,In_811,In_163);
nand U4243 (N_4243,In_1447,In_1207);
nor U4244 (N_4244,In_1020,In_589);
and U4245 (N_4245,In_1050,In_1417);
and U4246 (N_4246,In_1338,In_1099);
nand U4247 (N_4247,In_246,In_1434);
nand U4248 (N_4248,In_1444,In_1064);
or U4249 (N_4249,In_176,In_22);
nor U4250 (N_4250,In_370,In_1488);
nand U4251 (N_4251,In_148,In_1359);
or U4252 (N_4252,In_535,In_126);
nand U4253 (N_4253,In_1130,In_200);
nor U4254 (N_4254,In_1302,In_621);
xor U4255 (N_4255,In_1156,In_214);
and U4256 (N_4256,In_947,In_179);
and U4257 (N_4257,In_677,In_405);
xnor U4258 (N_4258,In_110,In_65);
nor U4259 (N_4259,In_767,In_279);
nand U4260 (N_4260,In_817,In_771);
xor U4261 (N_4261,In_770,In_497);
and U4262 (N_4262,In_54,In_825);
and U4263 (N_4263,In_1327,In_1117);
or U4264 (N_4264,In_1015,In_700);
and U4265 (N_4265,In_213,In_1145);
xor U4266 (N_4266,In_236,In_1381);
nand U4267 (N_4267,In_1295,In_1069);
nor U4268 (N_4268,In_676,In_1408);
nor U4269 (N_4269,In_1217,In_173);
or U4270 (N_4270,In_486,In_113);
and U4271 (N_4271,In_321,In_247);
nand U4272 (N_4272,In_1448,In_583);
or U4273 (N_4273,In_767,In_1213);
or U4274 (N_4274,In_241,In_16);
and U4275 (N_4275,In_1088,In_585);
xnor U4276 (N_4276,In_1436,In_1323);
nor U4277 (N_4277,In_988,In_335);
xnor U4278 (N_4278,In_270,In_273);
xnor U4279 (N_4279,In_141,In_1296);
nand U4280 (N_4280,In_582,In_783);
nand U4281 (N_4281,In_1237,In_1098);
nor U4282 (N_4282,In_94,In_74);
nand U4283 (N_4283,In_1284,In_540);
or U4284 (N_4284,In_1432,In_512);
nor U4285 (N_4285,In_891,In_1389);
and U4286 (N_4286,In_1328,In_1112);
nand U4287 (N_4287,In_358,In_625);
or U4288 (N_4288,In_1438,In_1163);
nand U4289 (N_4289,In_1004,In_534);
or U4290 (N_4290,In_1099,In_760);
or U4291 (N_4291,In_216,In_806);
nand U4292 (N_4292,In_1330,In_801);
or U4293 (N_4293,In_518,In_764);
xnor U4294 (N_4294,In_176,In_545);
nor U4295 (N_4295,In_325,In_568);
or U4296 (N_4296,In_185,In_1021);
and U4297 (N_4297,In_104,In_840);
and U4298 (N_4298,In_47,In_1342);
nand U4299 (N_4299,In_878,In_1012);
or U4300 (N_4300,In_279,In_1309);
or U4301 (N_4301,In_229,In_984);
or U4302 (N_4302,In_1409,In_120);
and U4303 (N_4303,In_1310,In_969);
and U4304 (N_4304,In_1208,In_275);
or U4305 (N_4305,In_97,In_790);
nor U4306 (N_4306,In_437,In_504);
nand U4307 (N_4307,In_116,In_1294);
or U4308 (N_4308,In_1224,In_475);
or U4309 (N_4309,In_367,In_624);
or U4310 (N_4310,In_1445,In_663);
and U4311 (N_4311,In_662,In_145);
nand U4312 (N_4312,In_100,In_207);
nor U4313 (N_4313,In_207,In_270);
or U4314 (N_4314,In_966,In_996);
nor U4315 (N_4315,In_820,In_120);
nor U4316 (N_4316,In_1116,In_458);
and U4317 (N_4317,In_1166,In_862);
or U4318 (N_4318,In_404,In_641);
and U4319 (N_4319,In_1274,In_141);
or U4320 (N_4320,In_993,In_343);
and U4321 (N_4321,In_637,In_415);
and U4322 (N_4322,In_972,In_340);
and U4323 (N_4323,In_553,In_543);
nor U4324 (N_4324,In_705,In_976);
xnor U4325 (N_4325,In_278,In_207);
nor U4326 (N_4326,In_1107,In_41);
or U4327 (N_4327,In_316,In_228);
or U4328 (N_4328,In_528,In_186);
nor U4329 (N_4329,In_1154,In_356);
xor U4330 (N_4330,In_1177,In_1317);
or U4331 (N_4331,In_469,In_839);
and U4332 (N_4332,In_803,In_755);
nand U4333 (N_4333,In_791,In_657);
or U4334 (N_4334,In_666,In_445);
nor U4335 (N_4335,In_213,In_590);
nor U4336 (N_4336,In_371,In_309);
xor U4337 (N_4337,In_1459,In_1326);
or U4338 (N_4338,In_74,In_927);
and U4339 (N_4339,In_1048,In_112);
nor U4340 (N_4340,In_1051,In_512);
or U4341 (N_4341,In_977,In_1310);
xnor U4342 (N_4342,In_41,In_1394);
xnor U4343 (N_4343,In_1473,In_628);
or U4344 (N_4344,In_1280,In_329);
and U4345 (N_4345,In_733,In_919);
nand U4346 (N_4346,In_1226,In_698);
or U4347 (N_4347,In_27,In_384);
or U4348 (N_4348,In_350,In_1219);
nor U4349 (N_4349,In_1054,In_685);
nand U4350 (N_4350,In_1299,In_1298);
or U4351 (N_4351,In_158,In_1452);
nand U4352 (N_4352,In_216,In_816);
nand U4353 (N_4353,In_1051,In_31);
and U4354 (N_4354,In_1264,In_578);
and U4355 (N_4355,In_804,In_837);
xnor U4356 (N_4356,In_1019,In_1015);
and U4357 (N_4357,In_166,In_1456);
or U4358 (N_4358,In_984,In_647);
nor U4359 (N_4359,In_504,In_559);
and U4360 (N_4360,In_663,In_621);
or U4361 (N_4361,In_355,In_406);
nor U4362 (N_4362,In_974,In_998);
nor U4363 (N_4363,In_693,In_457);
and U4364 (N_4364,In_307,In_457);
xor U4365 (N_4365,In_884,In_502);
nor U4366 (N_4366,In_15,In_986);
and U4367 (N_4367,In_638,In_536);
nor U4368 (N_4368,In_97,In_921);
nor U4369 (N_4369,In_1306,In_834);
nor U4370 (N_4370,In_1192,In_842);
nor U4371 (N_4371,In_1140,In_1118);
nand U4372 (N_4372,In_1210,In_528);
or U4373 (N_4373,In_35,In_129);
or U4374 (N_4374,In_290,In_1243);
or U4375 (N_4375,In_944,In_458);
or U4376 (N_4376,In_286,In_1191);
nand U4377 (N_4377,In_896,In_872);
or U4378 (N_4378,In_1432,In_378);
nand U4379 (N_4379,In_1482,In_1349);
nor U4380 (N_4380,In_734,In_655);
nor U4381 (N_4381,In_255,In_1236);
nor U4382 (N_4382,In_74,In_782);
and U4383 (N_4383,In_1442,In_757);
nor U4384 (N_4384,In_457,In_562);
nand U4385 (N_4385,In_549,In_112);
nor U4386 (N_4386,In_418,In_1430);
nand U4387 (N_4387,In_252,In_1146);
nand U4388 (N_4388,In_61,In_494);
or U4389 (N_4389,In_845,In_1453);
and U4390 (N_4390,In_1336,In_1248);
nor U4391 (N_4391,In_564,In_740);
or U4392 (N_4392,In_630,In_1396);
nor U4393 (N_4393,In_699,In_687);
nor U4394 (N_4394,In_389,In_1420);
or U4395 (N_4395,In_1366,In_202);
or U4396 (N_4396,In_757,In_1186);
nor U4397 (N_4397,In_333,In_1425);
and U4398 (N_4398,In_427,In_159);
xor U4399 (N_4399,In_1101,In_370);
and U4400 (N_4400,In_986,In_1080);
and U4401 (N_4401,In_1320,In_1181);
or U4402 (N_4402,In_786,In_549);
and U4403 (N_4403,In_1195,In_113);
and U4404 (N_4404,In_598,In_873);
and U4405 (N_4405,In_291,In_1313);
nand U4406 (N_4406,In_966,In_82);
nand U4407 (N_4407,In_1446,In_713);
nor U4408 (N_4408,In_24,In_1333);
nand U4409 (N_4409,In_45,In_1092);
or U4410 (N_4410,In_877,In_389);
xor U4411 (N_4411,In_46,In_750);
and U4412 (N_4412,In_1148,In_1300);
nor U4413 (N_4413,In_952,In_713);
nand U4414 (N_4414,In_1398,In_460);
nor U4415 (N_4415,In_119,In_1408);
and U4416 (N_4416,In_421,In_548);
or U4417 (N_4417,In_91,In_496);
or U4418 (N_4418,In_1449,In_467);
or U4419 (N_4419,In_17,In_705);
and U4420 (N_4420,In_1487,In_250);
nand U4421 (N_4421,In_356,In_937);
and U4422 (N_4422,In_1002,In_859);
or U4423 (N_4423,In_1353,In_723);
nand U4424 (N_4424,In_213,In_1134);
or U4425 (N_4425,In_357,In_470);
and U4426 (N_4426,In_544,In_1047);
and U4427 (N_4427,In_332,In_1054);
nand U4428 (N_4428,In_88,In_1490);
nand U4429 (N_4429,In_1328,In_686);
nor U4430 (N_4430,In_491,In_37);
or U4431 (N_4431,In_791,In_881);
or U4432 (N_4432,In_205,In_861);
and U4433 (N_4433,In_1134,In_1158);
nor U4434 (N_4434,In_353,In_894);
or U4435 (N_4435,In_267,In_270);
nand U4436 (N_4436,In_1341,In_634);
and U4437 (N_4437,In_1147,In_1091);
or U4438 (N_4438,In_688,In_1160);
or U4439 (N_4439,In_1119,In_655);
and U4440 (N_4440,In_229,In_1230);
nor U4441 (N_4441,In_551,In_1313);
and U4442 (N_4442,In_739,In_581);
nand U4443 (N_4443,In_560,In_810);
nor U4444 (N_4444,In_499,In_939);
xnor U4445 (N_4445,In_1239,In_423);
nor U4446 (N_4446,In_257,In_924);
xor U4447 (N_4447,In_1472,In_663);
or U4448 (N_4448,In_1078,In_417);
nor U4449 (N_4449,In_962,In_1383);
and U4450 (N_4450,In_560,In_945);
or U4451 (N_4451,In_862,In_530);
nor U4452 (N_4452,In_501,In_542);
and U4453 (N_4453,In_87,In_161);
xnor U4454 (N_4454,In_680,In_123);
nor U4455 (N_4455,In_1214,In_379);
nor U4456 (N_4456,In_640,In_118);
and U4457 (N_4457,In_872,In_344);
nand U4458 (N_4458,In_350,In_1283);
xor U4459 (N_4459,In_1365,In_386);
xnor U4460 (N_4460,In_1048,In_782);
and U4461 (N_4461,In_334,In_889);
xnor U4462 (N_4462,In_179,In_191);
nor U4463 (N_4463,In_1001,In_403);
nand U4464 (N_4464,In_311,In_1115);
and U4465 (N_4465,In_679,In_9);
and U4466 (N_4466,In_494,In_693);
nor U4467 (N_4467,In_434,In_1447);
nor U4468 (N_4468,In_1422,In_304);
and U4469 (N_4469,In_592,In_477);
xnor U4470 (N_4470,In_333,In_1400);
or U4471 (N_4471,In_1314,In_846);
nand U4472 (N_4472,In_1220,In_657);
nor U4473 (N_4473,In_398,In_662);
nor U4474 (N_4474,In_341,In_1000);
nor U4475 (N_4475,In_1265,In_305);
nor U4476 (N_4476,In_732,In_536);
nand U4477 (N_4477,In_1081,In_960);
nand U4478 (N_4478,In_924,In_606);
and U4479 (N_4479,In_511,In_391);
nor U4480 (N_4480,In_263,In_140);
or U4481 (N_4481,In_1132,In_284);
nor U4482 (N_4482,In_1275,In_345);
nand U4483 (N_4483,In_489,In_355);
and U4484 (N_4484,In_373,In_1414);
nor U4485 (N_4485,In_1299,In_1252);
or U4486 (N_4486,In_1030,In_720);
and U4487 (N_4487,In_1310,In_1447);
xor U4488 (N_4488,In_909,In_1434);
or U4489 (N_4489,In_951,In_587);
nor U4490 (N_4490,In_881,In_80);
or U4491 (N_4491,In_503,In_1236);
and U4492 (N_4492,In_232,In_939);
nor U4493 (N_4493,In_134,In_1396);
or U4494 (N_4494,In_81,In_36);
and U4495 (N_4495,In_826,In_993);
or U4496 (N_4496,In_291,In_1327);
or U4497 (N_4497,In_235,In_538);
or U4498 (N_4498,In_704,In_277);
nand U4499 (N_4499,In_202,In_1378);
or U4500 (N_4500,In_1231,In_848);
xor U4501 (N_4501,In_621,In_359);
and U4502 (N_4502,In_1109,In_756);
nor U4503 (N_4503,In_453,In_167);
nor U4504 (N_4504,In_631,In_1332);
nand U4505 (N_4505,In_56,In_375);
xor U4506 (N_4506,In_80,In_1293);
or U4507 (N_4507,In_803,In_709);
or U4508 (N_4508,In_1193,In_1073);
nor U4509 (N_4509,In_209,In_806);
or U4510 (N_4510,In_969,In_745);
and U4511 (N_4511,In_1420,In_1128);
nand U4512 (N_4512,In_451,In_97);
or U4513 (N_4513,In_636,In_767);
nor U4514 (N_4514,In_903,In_1201);
nor U4515 (N_4515,In_145,In_677);
or U4516 (N_4516,In_881,In_419);
and U4517 (N_4517,In_458,In_366);
nor U4518 (N_4518,In_344,In_20);
nand U4519 (N_4519,In_1292,In_1282);
nand U4520 (N_4520,In_40,In_1233);
or U4521 (N_4521,In_492,In_1169);
nor U4522 (N_4522,In_347,In_1222);
nor U4523 (N_4523,In_192,In_475);
or U4524 (N_4524,In_125,In_1057);
nor U4525 (N_4525,In_588,In_28);
or U4526 (N_4526,In_1185,In_926);
and U4527 (N_4527,In_671,In_603);
and U4528 (N_4528,In_1175,In_1222);
nand U4529 (N_4529,In_511,In_1111);
and U4530 (N_4530,In_1382,In_279);
nor U4531 (N_4531,In_1059,In_1291);
or U4532 (N_4532,In_1257,In_848);
nor U4533 (N_4533,In_451,In_1496);
nor U4534 (N_4534,In_886,In_127);
or U4535 (N_4535,In_451,In_724);
nand U4536 (N_4536,In_1433,In_293);
or U4537 (N_4537,In_1291,In_577);
or U4538 (N_4538,In_1223,In_1475);
nor U4539 (N_4539,In_281,In_382);
or U4540 (N_4540,In_438,In_147);
nand U4541 (N_4541,In_1056,In_762);
or U4542 (N_4542,In_940,In_1473);
or U4543 (N_4543,In_975,In_205);
nor U4544 (N_4544,In_910,In_319);
and U4545 (N_4545,In_873,In_1183);
nor U4546 (N_4546,In_193,In_656);
nand U4547 (N_4547,In_833,In_1453);
nand U4548 (N_4548,In_433,In_190);
nand U4549 (N_4549,In_972,In_250);
nand U4550 (N_4550,In_6,In_596);
or U4551 (N_4551,In_49,In_558);
nand U4552 (N_4552,In_1190,In_1104);
nand U4553 (N_4553,In_1260,In_49);
nor U4554 (N_4554,In_1012,In_726);
and U4555 (N_4555,In_1272,In_298);
nand U4556 (N_4556,In_585,In_805);
xor U4557 (N_4557,In_1264,In_382);
nor U4558 (N_4558,In_179,In_45);
or U4559 (N_4559,In_131,In_514);
nor U4560 (N_4560,In_686,In_135);
and U4561 (N_4561,In_1221,In_1176);
and U4562 (N_4562,In_319,In_1300);
xor U4563 (N_4563,In_710,In_928);
nand U4564 (N_4564,In_1498,In_1010);
nor U4565 (N_4565,In_942,In_556);
nand U4566 (N_4566,In_567,In_815);
or U4567 (N_4567,In_532,In_603);
and U4568 (N_4568,In_788,In_996);
nand U4569 (N_4569,In_53,In_1446);
xor U4570 (N_4570,In_1126,In_59);
and U4571 (N_4571,In_1194,In_467);
nor U4572 (N_4572,In_437,In_368);
nor U4573 (N_4573,In_426,In_737);
nand U4574 (N_4574,In_463,In_1408);
nor U4575 (N_4575,In_957,In_375);
nand U4576 (N_4576,In_1093,In_1187);
and U4577 (N_4577,In_866,In_663);
nand U4578 (N_4578,In_1384,In_180);
or U4579 (N_4579,In_225,In_926);
nand U4580 (N_4580,In_1499,In_710);
or U4581 (N_4581,In_646,In_676);
nor U4582 (N_4582,In_354,In_1478);
xnor U4583 (N_4583,In_1167,In_966);
or U4584 (N_4584,In_328,In_7);
or U4585 (N_4585,In_1165,In_1330);
and U4586 (N_4586,In_734,In_178);
nor U4587 (N_4587,In_1468,In_977);
or U4588 (N_4588,In_991,In_1430);
and U4589 (N_4589,In_673,In_131);
nor U4590 (N_4590,In_785,In_1452);
nor U4591 (N_4591,In_269,In_123);
or U4592 (N_4592,In_1262,In_554);
xnor U4593 (N_4593,In_1442,In_358);
xor U4594 (N_4594,In_1321,In_290);
nor U4595 (N_4595,In_171,In_238);
nand U4596 (N_4596,In_212,In_1305);
nand U4597 (N_4597,In_83,In_1454);
and U4598 (N_4598,In_404,In_714);
xor U4599 (N_4599,In_969,In_779);
or U4600 (N_4600,In_458,In_113);
nor U4601 (N_4601,In_1138,In_688);
and U4602 (N_4602,In_131,In_97);
and U4603 (N_4603,In_1238,In_1166);
or U4604 (N_4604,In_948,In_1235);
and U4605 (N_4605,In_1127,In_1383);
and U4606 (N_4606,In_283,In_461);
or U4607 (N_4607,In_410,In_841);
nand U4608 (N_4608,In_25,In_314);
or U4609 (N_4609,In_655,In_37);
or U4610 (N_4610,In_725,In_422);
or U4611 (N_4611,In_1065,In_406);
nand U4612 (N_4612,In_44,In_643);
xor U4613 (N_4613,In_1421,In_709);
or U4614 (N_4614,In_370,In_570);
nor U4615 (N_4615,In_1306,In_369);
nand U4616 (N_4616,In_529,In_1415);
and U4617 (N_4617,In_1291,In_825);
nor U4618 (N_4618,In_856,In_512);
nand U4619 (N_4619,In_1346,In_1057);
or U4620 (N_4620,In_110,In_940);
or U4621 (N_4621,In_96,In_956);
and U4622 (N_4622,In_1485,In_1206);
and U4623 (N_4623,In_850,In_1041);
nor U4624 (N_4624,In_297,In_484);
nor U4625 (N_4625,In_517,In_906);
or U4626 (N_4626,In_989,In_788);
or U4627 (N_4627,In_893,In_746);
or U4628 (N_4628,In_1274,In_525);
and U4629 (N_4629,In_1196,In_1086);
and U4630 (N_4630,In_1110,In_1229);
nor U4631 (N_4631,In_1253,In_653);
and U4632 (N_4632,In_727,In_164);
nor U4633 (N_4633,In_126,In_1008);
nand U4634 (N_4634,In_660,In_158);
or U4635 (N_4635,In_1254,In_37);
and U4636 (N_4636,In_558,In_746);
or U4637 (N_4637,In_1121,In_858);
nor U4638 (N_4638,In_249,In_1316);
nor U4639 (N_4639,In_989,In_991);
nand U4640 (N_4640,In_764,In_1358);
or U4641 (N_4641,In_1395,In_384);
nand U4642 (N_4642,In_472,In_19);
and U4643 (N_4643,In_516,In_565);
or U4644 (N_4644,In_1192,In_170);
and U4645 (N_4645,In_666,In_373);
and U4646 (N_4646,In_553,In_809);
and U4647 (N_4647,In_1395,In_745);
and U4648 (N_4648,In_1244,In_541);
nor U4649 (N_4649,In_25,In_632);
nor U4650 (N_4650,In_467,In_547);
nor U4651 (N_4651,In_1022,In_23);
nor U4652 (N_4652,In_160,In_978);
xor U4653 (N_4653,In_1104,In_657);
nor U4654 (N_4654,In_28,In_590);
nand U4655 (N_4655,In_115,In_506);
and U4656 (N_4656,In_103,In_1380);
nor U4657 (N_4657,In_736,In_1124);
or U4658 (N_4658,In_1268,In_625);
and U4659 (N_4659,In_592,In_706);
nor U4660 (N_4660,In_1323,In_897);
nand U4661 (N_4661,In_612,In_1235);
and U4662 (N_4662,In_617,In_203);
nor U4663 (N_4663,In_722,In_245);
and U4664 (N_4664,In_280,In_930);
xor U4665 (N_4665,In_1161,In_1128);
and U4666 (N_4666,In_763,In_70);
or U4667 (N_4667,In_1094,In_1147);
or U4668 (N_4668,In_894,In_1018);
nor U4669 (N_4669,In_1022,In_501);
and U4670 (N_4670,In_1438,In_8);
or U4671 (N_4671,In_254,In_1457);
and U4672 (N_4672,In_1124,In_269);
and U4673 (N_4673,In_1180,In_493);
or U4674 (N_4674,In_1267,In_132);
and U4675 (N_4675,In_847,In_1068);
xnor U4676 (N_4676,In_868,In_766);
and U4677 (N_4677,In_496,In_666);
or U4678 (N_4678,In_305,In_892);
nor U4679 (N_4679,In_1463,In_1209);
or U4680 (N_4680,In_444,In_509);
and U4681 (N_4681,In_1328,In_1418);
xnor U4682 (N_4682,In_1373,In_161);
and U4683 (N_4683,In_992,In_373);
nand U4684 (N_4684,In_66,In_25);
or U4685 (N_4685,In_1031,In_1047);
or U4686 (N_4686,In_107,In_38);
nand U4687 (N_4687,In_35,In_91);
nand U4688 (N_4688,In_908,In_58);
and U4689 (N_4689,In_1302,In_1043);
nor U4690 (N_4690,In_1103,In_459);
and U4691 (N_4691,In_1311,In_453);
or U4692 (N_4692,In_544,In_548);
and U4693 (N_4693,In_58,In_1297);
or U4694 (N_4694,In_1291,In_1355);
or U4695 (N_4695,In_978,In_1088);
or U4696 (N_4696,In_403,In_941);
xnor U4697 (N_4697,In_778,In_503);
or U4698 (N_4698,In_481,In_710);
and U4699 (N_4699,In_1236,In_556);
and U4700 (N_4700,In_162,In_68);
and U4701 (N_4701,In_155,In_813);
xnor U4702 (N_4702,In_1073,In_429);
or U4703 (N_4703,In_323,In_213);
nor U4704 (N_4704,In_1303,In_191);
or U4705 (N_4705,In_1364,In_20);
and U4706 (N_4706,In_1195,In_693);
nand U4707 (N_4707,In_32,In_695);
nor U4708 (N_4708,In_992,In_903);
or U4709 (N_4709,In_1230,In_155);
and U4710 (N_4710,In_560,In_1214);
nor U4711 (N_4711,In_499,In_334);
nand U4712 (N_4712,In_121,In_866);
or U4713 (N_4713,In_1034,In_90);
and U4714 (N_4714,In_125,In_1011);
nand U4715 (N_4715,In_71,In_896);
nor U4716 (N_4716,In_785,In_707);
or U4717 (N_4717,In_1341,In_986);
nand U4718 (N_4718,In_1010,In_885);
nand U4719 (N_4719,In_225,In_833);
xnor U4720 (N_4720,In_73,In_1085);
nor U4721 (N_4721,In_689,In_730);
and U4722 (N_4722,In_1115,In_1220);
nand U4723 (N_4723,In_1235,In_36);
nand U4724 (N_4724,In_769,In_1354);
xnor U4725 (N_4725,In_191,In_652);
or U4726 (N_4726,In_1209,In_934);
nand U4727 (N_4727,In_606,In_1425);
and U4728 (N_4728,In_1188,In_1356);
or U4729 (N_4729,In_169,In_928);
nor U4730 (N_4730,In_963,In_163);
nand U4731 (N_4731,In_371,In_545);
nand U4732 (N_4732,In_642,In_1241);
nor U4733 (N_4733,In_1366,In_404);
nand U4734 (N_4734,In_1173,In_487);
and U4735 (N_4735,In_567,In_380);
nand U4736 (N_4736,In_632,In_1206);
nor U4737 (N_4737,In_1285,In_236);
and U4738 (N_4738,In_1356,In_932);
nand U4739 (N_4739,In_176,In_1214);
nand U4740 (N_4740,In_1483,In_919);
nand U4741 (N_4741,In_958,In_765);
nand U4742 (N_4742,In_495,In_1002);
xor U4743 (N_4743,In_157,In_949);
xnor U4744 (N_4744,In_1411,In_799);
nand U4745 (N_4745,In_994,In_402);
nand U4746 (N_4746,In_1350,In_401);
and U4747 (N_4747,In_467,In_1004);
nand U4748 (N_4748,In_166,In_535);
nand U4749 (N_4749,In_987,In_654);
nand U4750 (N_4750,In_89,In_1467);
nand U4751 (N_4751,In_1198,In_355);
xor U4752 (N_4752,In_184,In_364);
nor U4753 (N_4753,In_608,In_509);
or U4754 (N_4754,In_1295,In_886);
xnor U4755 (N_4755,In_397,In_492);
or U4756 (N_4756,In_215,In_229);
or U4757 (N_4757,In_1095,In_1289);
nand U4758 (N_4758,In_1033,In_620);
and U4759 (N_4759,In_386,In_1458);
xnor U4760 (N_4760,In_927,In_548);
or U4761 (N_4761,In_695,In_1304);
and U4762 (N_4762,In_96,In_1332);
xnor U4763 (N_4763,In_330,In_438);
nand U4764 (N_4764,In_803,In_305);
nand U4765 (N_4765,In_266,In_215);
nand U4766 (N_4766,In_1483,In_1221);
and U4767 (N_4767,In_98,In_767);
and U4768 (N_4768,In_1289,In_818);
and U4769 (N_4769,In_1307,In_155);
xor U4770 (N_4770,In_83,In_305);
nor U4771 (N_4771,In_1333,In_1175);
nor U4772 (N_4772,In_1061,In_899);
nand U4773 (N_4773,In_1144,In_1383);
and U4774 (N_4774,In_1482,In_290);
and U4775 (N_4775,In_1385,In_1398);
or U4776 (N_4776,In_896,In_811);
and U4777 (N_4777,In_174,In_325);
and U4778 (N_4778,In_263,In_997);
and U4779 (N_4779,In_1142,In_888);
or U4780 (N_4780,In_293,In_1419);
nor U4781 (N_4781,In_1352,In_747);
xnor U4782 (N_4782,In_412,In_708);
or U4783 (N_4783,In_1456,In_551);
xor U4784 (N_4784,In_268,In_1328);
xor U4785 (N_4785,In_498,In_641);
and U4786 (N_4786,In_1145,In_276);
nand U4787 (N_4787,In_311,In_657);
nand U4788 (N_4788,In_329,In_836);
and U4789 (N_4789,In_882,In_87);
nand U4790 (N_4790,In_1045,In_1144);
nand U4791 (N_4791,In_1441,In_309);
nor U4792 (N_4792,In_161,In_765);
and U4793 (N_4793,In_364,In_689);
nand U4794 (N_4794,In_233,In_1106);
nor U4795 (N_4795,In_1049,In_439);
xnor U4796 (N_4796,In_1250,In_1252);
and U4797 (N_4797,In_792,In_472);
or U4798 (N_4798,In_764,In_1071);
nor U4799 (N_4799,In_367,In_36);
nor U4800 (N_4800,In_875,In_227);
or U4801 (N_4801,In_770,In_1492);
and U4802 (N_4802,In_1316,In_810);
nand U4803 (N_4803,In_571,In_605);
nor U4804 (N_4804,In_117,In_306);
and U4805 (N_4805,In_1294,In_136);
nand U4806 (N_4806,In_649,In_1349);
nand U4807 (N_4807,In_1102,In_135);
nor U4808 (N_4808,In_1065,In_1066);
and U4809 (N_4809,In_473,In_145);
nor U4810 (N_4810,In_153,In_1426);
and U4811 (N_4811,In_185,In_873);
or U4812 (N_4812,In_997,In_112);
or U4813 (N_4813,In_376,In_1074);
nor U4814 (N_4814,In_1279,In_769);
or U4815 (N_4815,In_1108,In_325);
nand U4816 (N_4816,In_674,In_835);
nor U4817 (N_4817,In_733,In_1361);
nand U4818 (N_4818,In_816,In_804);
nand U4819 (N_4819,In_429,In_337);
nand U4820 (N_4820,In_208,In_78);
nand U4821 (N_4821,In_693,In_1218);
and U4822 (N_4822,In_1324,In_389);
and U4823 (N_4823,In_340,In_1002);
xor U4824 (N_4824,In_1263,In_70);
nand U4825 (N_4825,In_1093,In_192);
nand U4826 (N_4826,In_624,In_485);
nand U4827 (N_4827,In_1058,In_382);
and U4828 (N_4828,In_794,In_280);
xnor U4829 (N_4829,In_1009,In_550);
nand U4830 (N_4830,In_199,In_818);
nand U4831 (N_4831,In_768,In_636);
nor U4832 (N_4832,In_1262,In_837);
nor U4833 (N_4833,In_594,In_189);
nor U4834 (N_4834,In_227,In_1176);
nand U4835 (N_4835,In_872,In_27);
nor U4836 (N_4836,In_730,In_62);
nor U4837 (N_4837,In_99,In_901);
nand U4838 (N_4838,In_643,In_372);
or U4839 (N_4839,In_693,In_386);
or U4840 (N_4840,In_20,In_503);
nand U4841 (N_4841,In_763,In_207);
nand U4842 (N_4842,In_254,In_431);
and U4843 (N_4843,In_1238,In_939);
or U4844 (N_4844,In_60,In_831);
nand U4845 (N_4845,In_1079,In_966);
or U4846 (N_4846,In_154,In_624);
and U4847 (N_4847,In_952,In_1395);
and U4848 (N_4848,In_293,In_845);
nand U4849 (N_4849,In_52,In_74);
nand U4850 (N_4850,In_219,In_850);
nor U4851 (N_4851,In_693,In_745);
nor U4852 (N_4852,In_265,In_544);
nor U4853 (N_4853,In_684,In_695);
or U4854 (N_4854,In_231,In_676);
and U4855 (N_4855,In_1214,In_1446);
and U4856 (N_4856,In_436,In_550);
or U4857 (N_4857,In_851,In_352);
or U4858 (N_4858,In_842,In_1297);
nand U4859 (N_4859,In_860,In_457);
nand U4860 (N_4860,In_797,In_601);
or U4861 (N_4861,In_142,In_1211);
or U4862 (N_4862,In_296,In_729);
or U4863 (N_4863,In_592,In_164);
or U4864 (N_4864,In_1091,In_134);
xnor U4865 (N_4865,In_1019,In_1266);
or U4866 (N_4866,In_307,In_1134);
xor U4867 (N_4867,In_1451,In_605);
xnor U4868 (N_4868,In_1390,In_1134);
and U4869 (N_4869,In_498,In_397);
and U4870 (N_4870,In_989,In_321);
nand U4871 (N_4871,In_4,In_777);
nand U4872 (N_4872,In_1316,In_1215);
or U4873 (N_4873,In_1381,In_802);
nor U4874 (N_4874,In_100,In_877);
nor U4875 (N_4875,In_300,In_20);
nand U4876 (N_4876,In_1111,In_1152);
nor U4877 (N_4877,In_149,In_1097);
nor U4878 (N_4878,In_347,In_185);
and U4879 (N_4879,In_87,In_622);
nand U4880 (N_4880,In_174,In_341);
or U4881 (N_4881,In_823,In_544);
nand U4882 (N_4882,In_1136,In_1197);
or U4883 (N_4883,In_1461,In_1181);
xnor U4884 (N_4884,In_1005,In_488);
xor U4885 (N_4885,In_1292,In_1421);
nand U4886 (N_4886,In_476,In_464);
nor U4887 (N_4887,In_415,In_479);
nor U4888 (N_4888,In_346,In_1164);
or U4889 (N_4889,In_1097,In_882);
nand U4890 (N_4890,In_259,In_1178);
nand U4891 (N_4891,In_167,In_1480);
nor U4892 (N_4892,In_1244,In_363);
and U4893 (N_4893,In_102,In_205);
nand U4894 (N_4894,In_223,In_450);
or U4895 (N_4895,In_849,In_1165);
nor U4896 (N_4896,In_1249,In_1255);
or U4897 (N_4897,In_352,In_354);
nor U4898 (N_4898,In_131,In_981);
xor U4899 (N_4899,In_1305,In_489);
or U4900 (N_4900,In_1057,In_1064);
nor U4901 (N_4901,In_319,In_258);
and U4902 (N_4902,In_7,In_1137);
and U4903 (N_4903,In_261,In_1366);
or U4904 (N_4904,In_344,In_865);
or U4905 (N_4905,In_338,In_992);
nand U4906 (N_4906,In_797,In_354);
xor U4907 (N_4907,In_250,In_1234);
and U4908 (N_4908,In_921,In_680);
and U4909 (N_4909,In_50,In_892);
nor U4910 (N_4910,In_635,In_1021);
or U4911 (N_4911,In_513,In_306);
or U4912 (N_4912,In_1244,In_1390);
and U4913 (N_4913,In_636,In_626);
or U4914 (N_4914,In_878,In_1421);
and U4915 (N_4915,In_885,In_1382);
nor U4916 (N_4916,In_858,In_79);
nor U4917 (N_4917,In_262,In_509);
xnor U4918 (N_4918,In_666,In_281);
and U4919 (N_4919,In_1188,In_452);
nor U4920 (N_4920,In_1176,In_656);
or U4921 (N_4921,In_484,In_118);
or U4922 (N_4922,In_1237,In_213);
xor U4923 (N_4923,In_669,In_857);
or U4924 (N_4924,In_1068,In_1380);
and U4925 (N_4925,In_14,In_1450);
nor U4926 (N_4926,In_1333,In_1189);
or U4927 (N_4927,In_1040,In_384);
and U4928 (N_4928,In_891,In_154);
nand U4929 (N_4929,In_1304,In_1341);
nor U4930 (N_4930,In_66,In_630);
nor U4931 (N_4931,In_238,In_284);
nand U4932 (N_4932,In_1459,In_956);
xnor U4933 (N_4933,In_410,In_837);
xor U4934 (N_4934,In_712,In_360);
nand U4935 (N_4935,In_1132,In_1048);
nand U4936 (N_4936,In_367,In_324);
and U4937 (N_4937,In_326,In_888);
and U4938 (N_4938,In_702,In_1392);
nand U4939 (N_4939,In_131,In_857);
nor U4940 (N_4940,In_650,In_1108);
or U4941 (N_4941,In_234,In_778);
and U4942 (N_4942,In_878,In_862);
and U4943 (N_4943,In_951,In_1231);
and U4944 (N_4944,In_957,In_1222);
nor U4945 (N_4945,In_144,In_359);
and U4946 (N_4946,In_1334,In_844);
or U4947 (N_4947,In_74,In_383);
nand U4948 (N_4948,In_93,In_1389);
xor U4949 (N_4949,In_833,In_1290);
nor U4950 (N_4950,In_1471,In_1495);
or U4951 (N_4951,In_467,In_1435);
and U4952 (N_4952,In_763,In_895);
nand U4953 (N_4953,In_1064,In_349);
or U4954 (N_4954,In_1035,In_138);
or U4955 (N_4955,In_1301,In_1469);
and U4956 (N_4956,In_39,In_1198);
and U4957 (N_4957,In_1412,In_479);
nor U4958 (N_4958,In_265,In_221);
nand U4959 (N_4959,In_190,In_1446);
and U4960 (N_4960,In_404,In_1029);
and U4961 (N_4961,In_914,In_96);
nand U4962 (N_4962,In_8,In_1319);
nor U4963 (N_4963,In_409,In_807);
nor U4964 (N_4964,In_924,In_74);
nor U4965 (N_4965,In_351,In_1293);
nor U4966 (N_4966,In_112,In_405);
nor U4967 (N_4967,In_325,In_104);
or U4968 (N_4968,In_900,In_6);
nand U4969 (N_4969,In_1012,In_713);
xor U4970 (N_4970,In_237,In_1096);
xnor U4971 (N_4971,In_1493,In_303);
and U4972 (N_4972,In_163,In_108);
and U4973 (N_4973,In_1020,In_1083);
xnor U4974 (N_4974,In_29,In_1326);
nand U4975 (N_4975,In_625,In_1099);
nand U4976 (N_4976,In_579,In_1490);
and U4977 (N_4977,In_1494,In_1397);
and U4978 (N_4978,In_1211,In_1312);
xor U4979 (N_4979,In_256,In_1448);
and U4980 (N_4980,In_552,In_549);
and U4981 (N_4981,In_439,In_811);
or U4982 (N_4982,In_1095,In_565);
nand U4983 (N_4983,In_737,In_280);
nand U4984 (N_4984,In_977,In_506);
nand U4985 (N_4985,In_283,In_224);
nand U4986 (N_4986,In_188,In_463);
or U4987 (N_4987,In_483,In_1114);
or U4988 (N_4988,In_1316,In_132);
and U4989 (N_4989,In_752,In_48);
and U4990 (N_4990,In_884,In_101);
and U4991 (N_4991,In_484,In_287);
nand U4992 (N_4992,In_1442,In_1320);
or U4993 (N_4993,In_808,In_849);
xnor U4994 (N_4994,In_842,In_637);
and U4995 (N_4995,In_422,In_732);
nand U4996 (N_4996,In_1002,In_697);
and U4997 (N_4997,In_986,In_314);
or U4998 (N_4998,In_933,In_688);
nand U4999 (N_4999,In_405,In_744);
xnor U5000 (N_5000,N_4608,N_773);
and U5001 (N_5001,N_675,N_3715);
and U5002 (N_5002,N_2505,N_802);
or U5003 (N_5003,N_1760,N_2725);
and U5004 (N_5004,N_4155,N_488);
nor U5005 (N_5005,N_3725,N_3542);
nand U5006 (N_5006,N_4435,N_3385);
nand U5007 (N_5007,N_1471,N_181);
or U5008 (N_5008,N_2634,N_1610);
and U5009 (N_5009,N_4105,N_1524);
nor U5010 (N_5010,N_2040,N_2203);
and U5011 (N_5011,N_487,N_954);
nor U5012 (N_5012,N_3994,N_72);
nand U5013 (N_5013,N_8,N_3489);
nor U5014 (N_5014,N_3632,N_3203);
and U5015 (N_5015,N_4755,N_1789);
xor U5016 (N_5016,N_1539,N_99);
nor U5017 (N_5017,N_3887,N_625);
and U5018 (N_5018,N_1284,N_4416);
or U5019 (N_5019,N_3142,N_447);
nand U5020 (N_5020,N_3791,N_4800);
or U5021 (N_5021,N_321,N_4475);
and U5022 (N_5022,N_93,N_3006);
nand U5023 (N_5023,N_3803,N_4510);
or U5024 (N_5024,N_3447,N_4296);
nand U5025 (N_5025,N_1562,N_4756);
or U5026 (N_5026,N_3174,N_424);
or U5027 (N_5027,N_859,N_393);
or U5028 (N_5028,N_804,N_2525);
nand U5029 (N_5029,N_2822,N_2978);
and U5030 (N_5030,N_3526,N_1341);
and U5031 (N_5031,N_1548,N_388);
nor U5032 (N_5032,N_4266,N_2351);
or U5033 (N_5033,N_4165,N_503);
and U5034 (N_5034,N_735,N_3429);
or U5035 (N_5035,N_452,N_4645);
xor U5036 (N_5036,N_4035,N_3047);
and U5037 (N_5037,N_1234,N_1272);
and U5038 (N_5038,N_1154,N_885);
nor U5039 (N_5039,N_4928,N_3735);
nor U5040 (N_5040,N_3235,N_3727);
and U5041 (N_5041,N_3989,N_1590);
and U5042 (N_5042,N_1630,N_1264);
nor U5043 (N_5043,N_754,N_3305);
xnor U5044 (N_5044,N_600,N_3968);
and U5045 (N_5045,N_2674,N_1681);
nor U5046 (N_5046,N_4770,N_2080);
nand U5047 (N_5047,N_3910,N_3594);
nor U5048 (N_5048,N_1959,N_519);
xnor U5049 (N_5049,N_4917,N_1768);
nor U5050 (N_5050,N_534,N_577);
or U5051 (N_5051,N_4114,N_4984);
and U5052 (N_5052,N_4649,N_1000);
nor U5053 (N_5053,N_1930,N_2032);
and U5054 (N_5054,N_893,N_1770);
or U5055 (N_5055,N_3901,N_1748);
or U5056 (N_5056,N_392,N_3882);
and U5057 (N_5057,N_1433,N_972);
and U5058 (N_5058,N_3605,N_3761);
nor U5059 (N_5059,N_3719,N_2999);
nand U5060 (N_5060,N_3547,N_2554);
xnor U5061 (N_5061,N_1546,N_4113);
nor U5062 (N_5062,N_3581,N_4279);
and U5063 (N_5063,N_286,N_975);
and U5064 (N_5064,N_2762,N_2001);
nor U5065 (N_5065,N_379,N_2852);
nand U5066 (N_5066,N_3330,N_2197);
xnor U5067 (N_5067,N_3357,N_4466);
and U5068 (N_5068,N_4977,N_3474);
nand U5069 (N_5069,N_3313,N_1099);
or U5070 (N_5070,N_3461,N_456);
nor U5071 (N_5071,N_3303,N_3877);
nor U5072 (N_5072,N_2140,N_2814);
nor U5073 (N_5073,N_3158,N_3783);
or U5074 (N_5074,N_1378,N_2177);
or U5075 (N_5075,N_563,N_2403);
and U5076 (N_5076,N_1063,N_4905);
nor U5077 (N_5077,N_2485,N_1321);
xnor U5078 (N_5078,N_2785,N_4093);
and U5079 (N_5079,N_3873,N_4090);
xnor U5080 (N_5080,N_3441,N_3199);
nand U5081 (N_5081,N_2755,N_1822);
and U5082 (N_5082,N_4999,N_3128);
or U5083 (N_5083,N_942,N_2482);
or U5084 (N_5084,N_4257,N_1672);
nor U5085 (N_5085,N_1273,N_2564);
and U5086 (N_5086,N_4620,N_1484);
nand U5087 (N_5087,N_3867,N_1201);
or U5088 (N_5088,N_3374,N_1015);
xor U5089 (N_5089,N_1018,N_3112);
or U5090 (N_5090,N_1737,N_2896);
nor U5091 (N_5091,N_4594,N_4931);
and U5092 (N_5092,N_3551,N_2656);
and U5093 (N_5093,N_2431,N_1830);
nand U5094 (N_5094,N_1485,N_4297);
and U5095 (N_5095,N_4727,N_575);
and U5096 (N_5096,N_3221,N_1310);
nor U5097 (N_5097,N_632,N_2663);
or U5098 (N_5098,N_4473,N_1425);
and U5099 (N_5099,N_3220,N_845);
and U5100 (N_5100,N_4916,N_1659);
and U5101 (N_5101,N_1567,N_892);
nand U5102 (N_5102,N_1337,N_1776);
or U5103 (N_5103,N_1502,N_2085);
or U5104 (N_5104,N_3646,N_949);
and U5105 (N_5105,N_3716,N_597);
nand U5106 (N_5106,N_173,N_3861);
and U5107 (N_5107,N_2865,N_2376);
nor U5108 (N_5108,N_4604,N_4553);
and U5109 (N_5109,N_3696,N_3245);
nand U5110 (N_5110,N_4720,N_700);
and U5111 (N_5111,N_444,N_3236);
and U5112 (N_5112,N_143,N_1331);
or U5113 (N_5113,N_3831,N_2353);
nand U5114 (N_5114,N_2838,N_4794);
nor U5115 (N_5115,N_1315,N_3744);
and U5116 (N_5116,N_4426,N_3216);
or U5117 (N_5117,N_1237,N_2344);
or U5118 (N_5118,N_3491,N_2114);
and U5119 (N_5119,N_355,N_2992);
and U5120 (N_5120,N_1363,N_684);
nor U5121 (N_5121,N_2898,N_3975);
or U5122 (N_5122,N_4764,N_1894);
and U5123 (N_5123,N_4228,N_2159);
or U5124 (N_5124,N_4327,N_4745);
nor U5125 (N_5125,N_4712,N_3611);
nand U5126 (N_5126,N_4486,N_3560);
and U5127 (N_5127,N_4600,N_592);
and U5128 (N_5128,N_959,N_713);
nand U5129 (N_5129,N_2602,N_1816);
nand U5130 (N_5130,N_4425,N_1143);
and U5131 (N_5131,N_50,N_41);
nand U5132 (N_5132,N_2325,N_378);
nor U5133 (N_5133,N_2112,N_1751);
and U5134 (N_5134,N_2954,N_1271);
and U5135 (N_5135,N_2231,N_2976);
and U5136 (N_5136,N_1389,N_2117);
nand U5137 (N_5137,N_188,N_3452);
or U5138 (N_5138,N_1710,N_883);
nor U5139 (N_5139,N_854,N_244);
and U5140 (N_5140,N_1611,N_4543);
nor U5141 (N_5141,N_4660,N_2433);
or U5142 (N_5142,N_331,N_4724);
nand U5143 (N_5143,N_258,N_1219);
and U5144 (N_5144,N_1617,N_4175);
nor U5145 (N_5145,N_3019,N_2448);
nor U5146 (N_5146,N_418,N_2584);
xnor U5147 (N_5147,N_1766,N_1179);
nand U5148 (N_5148,N_1207,N_4926);
or U5149 (N_5149,N_733,N_3002);
xor U5150 (N_5150,N_4786,N_4858);
nor U5151 (N_5151,N_4284,N_2609);
and U5152 (N_5152,N_1633,N_665);
and U5153 (N_5153,N_2710,N_1104);
or U5154 (N_5154,N_2746,N_799);
and U5155 (N_5155,N_3038,N_4803);
nor U5156 (N_5156,N_233,N_4455);
and U5157 (N_5157,N_1314,N_898);
nor U5158 (N_5158,N_4017,N_2851);
nor U5159 (N_5159,N_1288,N_4434);
and U5160 (N_5160,N_4170,N_2147);
nor U5161 (N_5161,N_3520,N_2410);
nor U5162 (N_5162,N_2733,N_1454);
xor U5163 (N_5163,N_4064,N_1616);
nor U5164 (N_5164,N_1754,N_4829);
nor U5165 (N_5165,N_4765,N_2761);
or U5166 (N_5166,N_4976,N_3155);
nand U5167 (N_5167,N_1834,N_2469);
nand U5168 (N_5168,N_4784,N_506);
nand U5169 (N_5169,N_2624,N_2039);
nand U5170 (N_5170,N_1896,N_3712);
or U5171 (N_5171,N_137,N_2421);
xor U5172 (N_5172,N_2628,N_2828);
nand U5173 (N_5173,N_3243,N_1380);
and U5174 (N_5174,N_1646,N_4873);
nor U5175 (N_5175,N_576,N_1108);
or U5176 (N_5176,N_3181,N_4186);
or U5177 (N_5177,N_492,N_4715);
and U5178 (N_5178,N_236,N_3396);
nor U5179 (N_5179,N_4520,N_4541);
nor U5180 (N_5180,N_2200,N_1447);
nor U5181 (N_5181,N_4855,N_1809);
and U5182 (N_5182,N_3763,N_3747);
nor U5183 (N_5183,N_1833,N_3410);
or U5184 (N_5184,N_3556,N_3045);
nand U5185 (N_5185,N_1372,N_421);
nand U5186 (N_5186,N_4337,N_4242);
nand U5187 (N_5187,N_1708,N_2515);
or U5188 (N_5188,N_4643,N_1678);
and U5189 (N_5189,N_3869,N_4082);
or U5190 (N_5190,N_2116,N_2827);
nor U5191 (N_5191,N_4598,N_2030);
nor U5192 (N_5192,N_2437,N_3257);
nor U5193 (N_5193,N_3499,N_2586);
nor U5194 (N_5194,N_510,N_692);
nand U5195 (N_5195,N_1903,N_3033);
nand U5196 (N_5196,N_2715,N_3493);
or U5197 (N_5197,N_2960,N_793);
nor U5198 (N_5198,N_3961,N_4156);
nand U5199 (N_5199,N_1139,N_1963);
nor U5200 (N_5200,N_4397,N_4393);
nor U5201 (N_5201,N_4391,N_3063);
nand U5202 (N_5202,N_4406,N_3490);
and U5203 (N_5203,N_2494,N_4025);
nor U5204 (N_5204,N_3825,N_2356);
nand U5205 (N_5205,N_3164,N_406);
or U5206 (N_5206,N_4813,N_3773);
or U5207 (N_5207,N_3371,N_2417);
nor U5208 (N_5208,N_1387,N_1893);
nor U5209 (N_5209,N_2512,N_4325);
and U5210 (N_5210,N_1037,N_3455);
or U5211 (N_5211,N_4112,N_3375);
xnor U5212 (N_5212,N_4775,N_3913);
nand U5213 (N_5213,N_710,N_1119);
or U5214 (N_5214,N_3933,N_3003);
nand U5215 (N_5215,N_2623,N_285);
nor U5216 (N_5216,N_561,N_4448);
nor U5217 (N_5217,N_3270,N_476);
nand U5218 (N_5218,N_1695,N_3917);
nor U5219 (N_5219,N_2178,N_24);
or U5220 (N_5220,N_4417,N_1427);
and U5221 (N_5221,N_1296,N_4878);
nor U5222 (N_5222,N_982,N_382);
nand U5223 (N_5223,N_2266,N_522);
nor U5224 (N_5224,N_3036,N_497);
nand U5225 (N_5225,N_1826,N_4061);
nor U5226 (N_5226,N_4730,N_477);
nand U5227 (N_5227,N_935,N_3579);
nand U5228 (N_5228,N_4676,N_1658);
xor U5229 (N_5229,N_2267,N_2873);
nor U5230 (N_5230,N_1192,N_475);
and U5231 (N_5231,N_2134,N_4521);
xnor U5232 (N_5232,N_2553,N_2858);
nor U5233 (N_5233,N_1973,N_2475);
and U5234 (N_5234,N_4320,N_1624);
nor U5235 (N_5235,N_3545,N_927);
or U5236 (N_5236,N_4394,N_2980);
nor U5237 (N_5237,N_2837,N_2078);
or U5238 (N_5238,N_3731,N_1482);
xnor U5239 (N_5239,N_4946,N_2043);
nor U5240 (N_5240,N_3781,N_1204);
and U5241 (N_5241,N_2079,N_940);
nand U5242 (N_5242,N_888,N_119);
nand U5243 (N_5243,N_2630,N_200);
and U5244 (N_5244,N_4652,N_2704);
and U5245 (N_5245,N_3765,N_224);
nand U5246 (N_5246,N_824,N_964);
xor U5247 (N_5247,N_5,N_2537);
or U5248 (N_5248,N_4276,N_4133);
nand U5249 (N_5249,N_2190,N_3134);
or U5250 (N_5250,N_2240,N_1325);
or U5251 (N_5251,N_2126,N_3925);
and U5252 (N_5252,N_2793,N_3196);
nand U5253 (N_5253,N_1553,N_3476);
and U5254 (N_5254,N_6,N_363);
and U5255 (N_5255,N_4490,N_2074);
nor U5256 (N_5256,N_4529,N_3207);
nand U5257 (N_5257,N_4566,N_144);
nand U5258 (N_5258,N_1141,N_1511);
and U5259 (N_5259,N_3984,N_4560);
and U5260 (N_5260,N_3934,N_1400);
and U5261 (N_5261,N_250,N_66);
nor U5262 (N_5262,N_243,N_2800);
nand U5263 (N_5263,N_2582,N_4011);
xnor U5264 (N_5264,N_4904,N_1551);
nand U5265 (N_5265,N_3008,N_1463);
and U5266 (N_5266,N_1699,N_4030);
nor U5267 (N_5267,N_607,N_4734);
nor U5268 (N_5268,N_825,N_2075);
xnor U5269 (N_5269,N_3088,N_3955);
or U5270 (N_5270,N_3480,N_221);
or U5271 (N_5271,N_2377,N_1755);
nand U5272 (N_5272,N_4287,N_1625);
and U5273 (N_5273,N_715,N_4439);
or U5274 (N_5274,N_4153,N_4449);
and U5275 (N_5275,N_57,N_208);
nand U5276 (N_5276,N_4331,N_4725);
nand U5277 (N_5277,N_4124,N_2971);
nand U5278 (N_5278,N_4507,N_4695);
or U5279 (N_5279,N_2579,N_1374);
or U5280 (N_5280,N_1905,N_4815);
or U5281 (N_5281,N_3487,N_384);
nand U5282 (N_5282,N_3194,N_235);
xor U5283 (N_5283,N_4733,N_1360);
and U5284 (N_5284,N_2633,N_2681);
nor U5285 (N_5285,N_3321,N_4856);
nand U5286 (N_5286,N_3623,N_1275);
nor U5287 (N_5287,N_3211,N_2990);
nor U5288 (N_5288,N_1815,N_1530);
nor U5289 (N_5289,N_2373,N_3456);
nand U5290 (N_5290,N_2522,N_3826);
nor U5291 (N_5291,N_1690,N_2284);
or U5292 (N_5292,N_2622,N_3509);
nor U5293 (N_5293,N_3760,N_2845);
or U5294 (N_5294,N_1129,N_2765);
or U5295 (N_5295,N_3574,N_2527);
or U5296 (N_5296,N_2955,N_2491);
or U5297 (N_5297,N_2010,N_1174);
and U5298 (N_5298,N_4809,N_2929);
or U5299 (N_5299,N_3732,N_1759);
nand U5300 (N_5300,N_498,N_1342);
nand U5301 (N_5301,N_4177,N_2864);
nor U5302 (N_5302,N_2682,N_2272);
nand U5303 (N_5303,N_861,N_718);
or U5304 (N_5304,N_2042,N_4859);
nand U5305 (N_5305,N_4253,N_1767);
nand U5306 (N_5306,N_971,N_1501);
xnor U5307 (N_5307,N_4833,N_4729);
nand U5308 (N_5308,N_2069,N_4920);
or U5309 (N_5309,N_2277,N_1094);
nand U5310 (N_5310,N_4942,N_4357);
and U5311 (N_5311,N_329,N_3100);
or U5312 (N_5312,N_2620,N_3156);
nor U5313 (N_5313,N_390,N_3498);
xnor U5314 (N_5314,N_4514,N_1067);
or U5315 (N_5315,N_2343,N_2476);
nor U5316 (N_5316,N_1598,N_4877);
or U5317 (N_5317,N_3056,N_2558);
or U5318 (N_5318,N_309,N_1749);
nor U5319 (N_5319,N_2490,N_609);
or U5320 (N_5320,N_1704,N_1361);
nor U5321 (N_5321,N_1895,N_2359);
and U5322 (N_5322,N_91,N_2253);
or U5323 (N_5323,N_4158,N_2795);
or U5324 (N_5324,N_1956,N_4995);
and U5325 (N_5325,N_3558,N_4590);
nand U5326 (N_5326,N_1126,N_3578);
nand U5327 (N_5327,N_1522,N_352);
nor U5328 (N_5328,N_1262,N_3276);
and U5329 (N_5329,N_1718,N_3705);
nand U5330 (N_5330,N_4029,N_1902);
nand U5331 (N_5331,N_3432,N_849);
and U5332 (N_5332,N_3025,N_1137);
nand U5333 (N_5333,N_4741,N_1571);
and U5334 (N_5334,N_4005,N_4094);
nand U5335 (N_5335,N_2939,N_4077);
nand U5336 (N_5336,N_3559,N_2540);
and U5337 (N_5337,N_4147,N_2248);
and U5338 (N_5338,N_1191,N_603);
nor U5339 (N_5339,N_517,N_1281);
and U5340 (N_5340,N_4948,N_3580);
nor U5341 (N_5341,N_1245,N_357);
and U5342 (N_5342,N_88,N_4204);
or U5343 (N_5343,N_225,N_1478);
nand U5344 (N_5344,N_986,N_4459);
nand U5345 (N_5345,N_3401,N_2593);
and U5346 (N_5346,N_3959,N_2199);
nor U5347 (N_5347,N_3141,N_58);
or U5348 (N_5348,N_3513,N_267);
or U5349 (N_5349,N_1451,N_1332);
nor U5350 (N_5350,N_4828,N_4339);
nand U5351 (N_5351,N_3752,N_3706);
xor U5352 (N_5352,N_3876,N_2514);
xor U5353 (N_5353,N_1979,N_1928);
and U5354 (N_5354,N_1879,N_164);
or U5355 (N_5355,N_2568,N_1692);
or U5356 (N_5356,N_75,N_714);
or U5357 (N_5357,N_526,N_4618);
and U5358 (N_5358,N_3845,N_2328);
nor U5359 (N_5359,N_2563,N_4631);
nand U5360 (N_5360,N_3315,N_1212);
nor U5361 (N_5361,N_4360,N_1863);
and U5362 (N_5362,N_3960,N_511);
or U5363 (N_5363,N_4198,N_1838);
or U5364 (N_5364,N_3092,N_4167);
or U5365 (N_5365,N_4440,N_4232);
nor U5366 (N_5366,N_3683,N_2647);
nand U5367 (N_5367,N_3777,N_1085);
or U5368 (N_5368,N_4996,N_1596);
xor U5369 (N_5369,N_3746,N_2830);
nor U5370 (N_5370,N_3399,N_1714);
nand U5371 (N_5371,N_2182,N_4401);
or U5372 (N_5372,N_409,N_4713);
and U5373 (N_5373,N_4988,N_1213);
nand U5374 (N_5374,N_3844,N_2057);
nor U5375 (N_5375,N_3163,N_3981);
xor U5376 (N_5376,N_2481,N_3109);
xor U5377 (N_5377,N_699,N_2108);
nor U5378 (N_5378,N_86,N_3484);
nand U5379 (N_5379,N_3880,N_3479);
nand U5380 (N_5380,N_4328,N_559);
or U5381 (N_5381,N_4958,N_2901);
or U5382 (N_5382,N_1805,N_4666);
xor U5383 (N_5383,N_948,N_3011);
nor U5384 (N_5384,N_3742,N_4497);
xnor U5385 (N_5385,N_633,N_4648);
xor U5386 (N_5386,N_3124,N_4016);
and U5387 (N_5387,N_1856,N_3978);
or U5388 (N_5388,N_3846,N_3685);
nand U5389 (N_5389,N_997,N_4240);
nor U5390 (N_5390,N_1392,N_55);
and U5391 (N_5391,N_2161,N_1664);
or U5392 (N_5392,N_2321,N_3552);
nor U5393 (N_5393,N_3793,N_3443);
nand U5394 (N_5394,N_120,N_455);
or U5395 (N_5395,N_4699,N_2594);
nor U5396 (N_5396,N_900,N_115);
nand U5397 (N_5397,N_1461,N_1350);
and U5398 (N_5398,N_690,N_2903);
nand U5399 (N_5399,N_202,N_59);
or U5400 (N_5400,N_568,N_1801);
and U5401 (N_5401,N_186,N_187);
xor U5402 (N_5402,N_4525,N_4019);
nor U5403 (N_5403,N_4033,N_3932);
or U5404 (N_5404,N_3523,N_70);
or U5405 (N_5405,N_438,N_1800);
or U5406 (N_5406,N_2972,N_794);
nor U5407 (N_5407,N_847,N_4465);
or U5408 (N_5408,N_2347,N_622);
or U5409 (N_5409,N_2011,N_259);
and U5410 (N_5410,N_3347,N_2744);
nor U5411 (N_5411,N_4739,N_3749);
nand U5412 (N_5412,N_4189,N_3833);
or U5413 (N_5413,N_4697,N_247);
or U5414 (N_5414,N_1430,N_2191);
and U5415 (N_5415,N_670,N_509);
and U5416 (N_5416,N_2463,N_3757);
xor U5417 (N_5417,N_3799,N_1700);
or U5418 (N_5418,N_1339,N_274);
or U5419 (N_5419,N_3295,N_201);
or U5420 (N_5420,N_229,N_4506);
nand U5421 (N_5421,N_4385,N_4359);
and U5422 (N_5422,N_3254,N_827);
and U5423 (N_5423,N_3483,N_4683);
or U5424 (N_5424,N_4613,N_4122);
nor U5425 (N_5425,N_2691,N_3848);
or U5426 (N_5426,N_106,N_4661);
nand U5427 (N_5427,N_2677,N_4111);
or U5428 (N_5428,N_2775,N_3979);
xor U5429 (N_5429,N_2638,N_4632);
and U5430 (N_5430,N_1517,N_4131);
and U5431 (N_5431,N_105,N_4312);
xnor U5432 (N_5432,N_2459,N_4126);
xor U5433 (N_5433,N_968,N_462);
nand U5434 (N_5434,N_2504,N_4621);
and U5435 (N_5435,N_4736,N_1428);
nor U5436 (N_5436,N_4623,N_3230);
and U5437 (N_5437,N_4032,N_96);
nand U5438 (N_5438,N_4689,N_3703);
nand U5439 (N_5439,N_4362,N_2879);
xnor U5440 (N_5440,N_1136,N_1937);
nand U5441 (N_5441,N_2872,N_2528);
and U5442 (N_5442,N_4628,N_3435);
and U5443 (N_5443,N_461,N_3114);
xnor U5444 (N_5444,N_2922,N_2397);
xnor U5445 (N_5445,N_3338,N_4280);
xor U5446 (N_5446,N_423,N_1588);
or U5447 (N_5447,N_2849,N_2209);
and U5448 (N_5448,N_1398,N_1939);
and U5449 (N_5449,N_704,N_3774);
nor U5450 (N_5450,N_784,N_1601);
or U5451 (N_5451,N_1906,N_1340);
nand U5452 (N_5452,N_3176,N_541);
nor U5453 (N_5453,N_4914,N_2570);
xor U5454 (N_5454,N_1819,N_4587);
xnor U5455 (N_5455,N_812,N_4959);
nor U5456 (N_5456,N_4669,N_1745);
nor U5457 (N_5457,N_3729,N_4052);
or U5458 (N_5458,N_2918,N_1420);
xor U5459 (N_5459,N_3640,N_151);
nand U5460 (N_5460,N_257,N_2044);
or U5461 (N_5461,N_1852,N_640);
nor U5462 (N_5462,N_434,N_2668);
xnor U5463 (N_5463,N_481,N_4943);
or U5464 (N_5464,N_3726,N_1300);
or U5465 (N_5465,N_3197,N_2041);
nand U5466 (N_5466,N_350,N_1044);
and U5467 (N_5467,N_2627,N_4247);
nor U5468 (N_5468,N_3954,N_3373);
nand U5469 (N_5469,N_3332,N_2866);
nand U5470 (N_5470,N_1265,N_2082);
or U5471 (N_5471,N_2649,N_210);
or U5472 (N_5472,N_3815,N_4622);
nor U5473 (N_5473,N_788,N_389);
nor U5474 (N_5474,N_3039,N_45);
xnor U5475 (N_5475,N_2058,N_1694);
and U5476 (N_5476,N_4120,N_1267);
or U5477 (N_5477,N_4640,N_1597);
nor U5478 (N_5478,N_2832,N_1866);
and U5479 (N_5479,N_3187,N_2149);
and U5480 (N_5480,N_4326,N_4180);
nor U5481 (N_5481,N_3204,N_4009);
or U5482 (N_5482,N_4421,N_4504);
and U5483 (N_5483,N_2234,N_341);
xnor U5484 (N_5484,N_3172,N_94);
or U5485 (N_5485,N_146,N_993);
or U5486 (N_5486,N_613,N_1916);
nand U5487 (N_5487,N_3360,N_3297);
nor U5488 (N_5488,N_3586,N_2840);
or U5489 (N_5489,N_4691,N_3170);
and U5490 (N_5490,N_2263,N_1200);
nor U5491 (N_5491,N_1648,N_275);
and U5492 (N_5492,N_3288,N_1656);
nor U5493 (N_5493,N_1933,N_3445);
and U5494 (N_5494,N_2856,N_454);
and U5495 (N_5495,N_4171,N_649);
and U5496 (N_5496,N_589,N_2261);
or U5497 (N_5497,N_203,N_3054);
or U5498 (N_5498,N_2789,N_272);
and U5499 (N_5499,N_2081,N_3496);
or U5500 (N_5500,N_2868,N_3784);
nand U5501 (N_5501,N_4013,N_2306);
or U5502 (N_5502,N_3267,N_1604);
or U5503 (N_5503,N_4684,N_4740);
or U5504 (N_5504,N_2440,N_2786);
nor U5505 (N_5505,N_4291,N_156);
nand U5506 (N_5506,N_2552,N_2699);
and U5507 (N_5507,N_1958,N_4407);
or U5508 (N_5508,N_3255,N_134);
and U5509 (N_5509,N_4785,N_43);
nor U5510 (N_5510,N_270,N_3262);
and U5511 (N_5511,N_2046,N_2472);
and U5512 (N_5512,N_3677,N_3208);
and U5513 (N_5513,N_1479,N_628);
nor U5514 (N_5514,N_2457,N_4103);
nor U5515 (N_5515,N_4701,N_1936);
nor U5516 (N_5516,N_1460,N_1810);
nor U5517 (N_5517,N_855,N_4488);
or U5518 (N_5518,N_2096,N_3530);
or U5519 (N_5519,N_4709,N_4467);
and U5520 (N_5520,N_4834,N_3521);
nor U5521 (N_5521,N_333,N_2608);
xnor U5522 (N_5522,N_49,N_2395);
or U5523 (N_5523,N_97,N_1515);
and U5524 (N_5524,N_1090,N_2648);
and U5525 (N_5525,N_4883,N_399);
nand U5526 (N_5526,N_771,N_2432);
xor U5527 (N_5527,N_2227,N_1638);
or U5528 (N_5528,N_1124,N_1946);
nor U5529 (N_5529,N_1434,N_3709);
or U5530 (N_5530,N_1279,N_3862);
nor U5531 (N_5531,N_4989,N_4963);
or U5532 (N_5532,N_4896,N_1717);
and U5533 (N_5533,N_1188,N_2927);
or U5534 (N_5534,N_4788,N_3012);
or U5535 (N_5535,N_87,N_3906);
nor U5536 (N_5536,N_3193,N_749);
nor U5537 (N_5537,N_2,N_3004);
and U5538 (N_5538,N_1112,N_3666);
nor U5539 (N_5539,N_3974,N_4731);
or U5540 (N_5540,N_1101,N_2251);
nand U5541 (N_5541,N_167,N_4509);
or U5542 (N_5542,N_4929,N_3770);
or U5543 (N_5543,N_3549,N_2580);
or U5544 (N_5544,N_26,N_1399);
or U5545 (N_5545,N_116,N_3736);
or U5546 (N_5546,N_4722,N_1226);
or U5547 (N_5547,N_4748,N_4454);
or U5548 (N_5548,N_4256,N_1045);
and U5549 (N_5549,N_2520,N_3776);
nor U5550 (N_5550,N_1357,N_1961);
nand U5551 (N_5551,N_2895,N_2592);
or U5552 (N_5552,N_2450,N_2008);
and U5553 (N_5553,N_158,N_51);
or U5554 (N_5554,N_4344,N_2414);
xnor U5555 (N_5555,N_1923,N_1208);
or U5556 (N_5556,N_4261,N_2309);
or U5557 (N_5557,N_2973,N_976);
nor U5558 (N_5558,N_2679,N_276);
nor U5559 (N_5559,N_2033,N_245);
nand U5560 (N_5560,N_223,N_17);
xor U5561 (N_5561,N_3294,N_4168);
nor U5562 (N_5562,N_484,N_1224);
nor U5563 (N_5563,N_4519,N_3237);
nand U5564 (N_5564,N_2363,N_3829);
nand U5565 (N_5565,N_3886,N_3676);
xor U5566 (N_5566,N_3247,N_7);
or U5567 (N_5567,N_1729,N_4481);
or U5568 (N_5568,N_2956,N_2911);
nand U5569 (N_5569,N_4332,N_790);
nor U5570 (N_5570,N_2278,N_4721);
nor U5571 (N_5571,N_1318,N_1202);
xor U5572 (N_5572,N_4562,N_3400);
and U5573 (N_5573,N_1086,N_620);
xor U5574 (N_5574,N_4458,N_3641);
or U5575 (N_5575,N_4670,N_4574);
and U5576 (N_5576,N_1238,N_842);
and U5577 (N_5577,N_2498,N_2768);
and U5578 (N_5578,N_1582,N_734);
and U5579 (N_5579,N_2607,N_951);
or U5580 (N_5580,N_2384,N_4269);
and U5581 (N_5581,N_4318,N_4379);
and U5582 (N_5582,N_4614,N_4906);
xor U5583 (N_5583,N_1869,N_47);
and U5584 (N_5584,N_3782,N_868);
and U5585 (N_5585,N_3367,N_4979);
nor U5586 (N_5586,N_3670,N_108);
nor U5587 (N_5587,N_4162,N_536);
xor U5588 (N_5588,N_4872,N_4096);
or U5589 (N_5589,N_197,N_4068);
nor U5590 (N_5590,N_3963,N_548);
or U5591 (N_5591,N_1716,N_3885);
and U5592 (N_5592,N_4665,N_3541);
and U5593 (N_5593,N_3902,N_3076);
xor U5594 (N_5594,N_819,N_2664);
or U5595 (N_5595,N_3116,N_1579);
or U5596 (N_5596,N_214,N_1075);
or U5597 (N_5597,N_2683,N_4299);
nor U5598 (N_5598,N_1335,N_3673);
nand U5599 (N_5599,N_1413,N_4642);
nand U5600 (N_5600,N_2531,N_783);
and U5601 (N_5601,N_4353,N_4463);
and U5602 (N_5602,N_1367,N_1668);
nor U5603 (N_5603,N_1925,N_1583);
nor U5604 (N_5604,N_2402,N_2862);
and U5605 (N_5605,N_1573,N_3015);
xor U5606 (N_5606,N_4802,N_1701);
nand U5607 (N_5607,N_3206,N_727);
and U5608 (N_5608,N_1613,N_3224);
nor U5609 (N_5609,N_1947,N_2415);
xor U5610 (N_5610,N_4049,N_2219);
and U5611 (N_5611,N_877,N_809);
nor U5612 (N_5612,N_3470,N_2936);
or U5613 (N_5613,N_1159,N_397);
nor U5614 (N_5614,N_2312,N_3477);
and U5615 (N_5615,N_1087,N_2500);
nor U5616 (N_5616,N_1941,N_2556);
nor U5617 (N_5617,N_1263,N_312);
nand U5618 (N_5618,N_1125,N_4107);
and U5619 (N_5619,N_4451,N_601);
and U5620 (N_5620,N_1419,N_283);
and U5621 (N_5621,N_178,N_4647);
or U5622 (N_5622,N_2890,N_4692);
nor U5623 (N_5623,N_565,N_2145);
and U5624 (N_5624,N_3821,N_4098);
nor U5625 (N_5625,N_915,N_3406);
nand U5626 (N_5626,N_1406,N_4235);
nor U5627 (N_5627,N_3263,N_1371);
nand U5628 (N_5628,N_891,N_3044);
xor U5629 (N_5629,N_585,N_2239);
nand U5630 (N_5630,N_4363,N_3524);
xor U5631 (N_5631,N_2925,N_2148);
and U5632 (N_5632,N_4213,N_4974);
nor U5633 (N_5633,N_1679,N_2619);
and U5634 (N_5634,N_3766,N_1870);
nor U5635 (N_5635,N_924,N_1697);
nor U5636 (N_5636,N_1199,N_637);
nand U5637 (N_5637,N_2217,N_90);
nand U5638 (N_5638,N_2232,N_1725);
and U5639 (N_5639,N_405,N_1747);
nand U5640 (N_5640,N_2362,N_1404);
nand U5641 (N_5641,N_2717,N_2212);
nor U5642 (N_5642,N_1877,N_3079);
or U5643 (N_5643,N_4573,N_2269);
nor U5644 (N_5644,N_3890,N_366);
or U5645 (N_5645,N_3278,N_3059);
or U5646 (N_5646,N_4210,N_757);
nor U5647 (N_5647,N_4063,N_4476);
nand U5648 (N_5648,N_1943,N_4078);
nand U5649 (N_5649,N_2213,N_2599);
nor U5650 (N_5650,N_2365,N_2151);
nand U5651 (N_5651,N_2270,N_1525);
nand U5652 (N_5652,N_4278,N_2951);
nor U5653 (N_5653,N_1942,N_792);
or U5654 (N_5654,N_2577,N_1009);
or U5655 (N_5655,N_3273,N_231);
xnor U5656 (N_5656,N_0,N_4460);
or U5657 (N_5657,N_3463,N_3497);
or U5658 (N_5658,N_3430,N_2728);
nand U5659 (N_5659,N_4452,N_3383);
nor U5660 (N_5660,N_2738,N_2012);
nor U5661 (N_5661,N_1720,N_3017);
and U5662 (N_5662,N_1807,N_4453);
nor U5663 (N_5663,N_122,N_3972);
nand U5664 (N_5664,N_4551,N_2439);
nand U5665 (N_5665,N_261,N_4196);
nand U5666 (N_5666,N_2771,N_1259);
nand U5667 (N_5667,N_3929,N_2798);
nand U5668 (N_5668,N_2796,N_1121);
xor U5669 (N_5669,N_1523,N_1170);
or U5670 (N_5670,N_4415,N_1401);
nor U5671 (N_5671,N_4742,N_1538);
nand U5672 (N_5672,N_2610,N_4542);
and U5673 (N_5673,N_3123,N_109);
and U5674 (N_5674,N_182,N_2655);
nor U5675 (N_5675,N_570,N_3593);
and U5676 (N_5676,N_3231,N_1868);
and U5677 (N_5677,N_650,N_4058);
and U5678 (N_5678,N_4879,N_540);
or U5679 (N_5679,N_3022,N_4899);
or U5680 (N_5680,N_4629,N_3723);
and U5681 (N_5681,N_386,N_3185);
and U5682 (N_5682,N_3608,N_1676);
and U5683 (N_5683,N_4143,N_4150);
or U5684 (N_5684,N_3748,N_4997);
or U5685 (N_5685,N_654,N_3688);
and U5686 (N_5686,N_4840,N_2385);
or U5687 (N_5687,N_3292,N_2824);
xor U5688 (N_5688,N_2387,N_1786);
or U5689 (N_5689,N_2706,N_4793);
nor U5690 (N_5690,N_3787,N_789);
nor U5691 (N_5691,N_4501,N_4842);
nand U5692 (N_5692,N_631,N_705);
nor U5693 (N_5693,N_1190,N_445);
or U5694 (N_5694,N_3926,N_4268);
nand U5695 (N_5695,N_2867,N_142);
nor U5696 (N_5696,N_2228,N_1294);
and U5697 (N_5697,N_3965,N_3310);
and U5698 (N_5698,N_2535,N_1057);
or U5699 (N_5699,N_2523,N_1195);
nand U5700 (N_5700,N_2238,N_3319);
nor U5701 (N_5701,N_2835,N_3418);
and U5702 (N_5702,N_779,N_1071);
and U5703 (N_5703,N_3398,N_1004);
and U5704 (N_5704,N_425,N_1945);
or U5705 (N_5705,N_4023,N_3834);
or U5706 (N_5706,N_1519,N_4627);
and U5707 (N_5707,N_1149,N_4042);
and U5708 (N_5708,N_365,N_15);
or U5709 (N_5709,N_3626,N_2425);
nor U5710 (N_5710,N_3153,N_4239);
nor U5711 (N_5711,N_2615,N_2210);
and U5712 (N_5712,N_4681,N_374);
or U5713 (N_5713,N_1727,N_1068);
or U5714 (N_5714,N_159,N_1411);
and U5715 (N_5715,N_2984,N_2792);
xor U5716 (N_5716,N_1825,N_685);
and U5717 (N_5717,N_398,N_1858);
and U5718 (N_5718,N_3812,N_4045);
xor U5719 (N_5719,N_190,N_2413);
nand U5720 (N_5720,N_797,N_598);
or U5721 (N_5721,N_2211,N_3555);
nor U5722 (N_5722,N_1527,N_135);
nand U5723 (N_5723,N_3462,N_1019);
xor U5724 (N_5724,N_562,N_969);
nand U5725 (N_5725,N_4932,N_1088);
nor U5726 (N_5726,N_3261,N_2908);
nand U5727 (N_5727,N_2705,N_703);
nor U5728 (N_5728,N_2479,N_4173);
and U5729 (N_5729,N_2135,N_2870);
and U5730 (N_5730,N_4399,N_1257);
and U5731 (N_5731,N_2567,N_803);
xor U5732 (N_5732,N_4060,N_148);
nor U5733 (N_5733,N_4292,N_4938);
or U5734 (N_5734,N_867,N_450);
nor U5735 (N_5735,N_1351,N_2614);
nor U5736 (N_5736,N_4915,N_912);
xor U5737 (N_5737,N_92,N_2468);
or U5738 (N_5738,N_4558,N_3506);
nor U5739 (N_5739,N_3215,N_4936);
or U5740 (N_5740,N_2855,N_2037);
or U5741 (N_5741,N_903,N_1472);
nor U5742 (N_5742,N_3654,N_1054);
xor U5743 (N_5743,N_485,N_2545);
and U5744 (N_5744,N_4199,N_725);
nand U5745 (N_5745,N_1774,N_1347);
nor U5746 (N_5746,N_1880,N_4726);
xor U5747 (N_5747,N_4650,N_2115);
nand U5748 (N_5748,N_2533,N_4298);
or U5749 (N_5749,N_1097,N_4769);
and U5750 (N_5750,N_2281,N_1240);
nor U5751 (N_5751,N_2300,N_3052);
and U5752 (N_5752,N_3997,N_2934);
nand U5753 (N_5753,N_2051,N_639);
nand U5754 (N_5754,N_3837,N_1053);
and U5755 (N_5755,N_1565,N_3678);
nor U5756 (N_5756,N_501,N_1989);
xnor U5757 (N_5757,N_3192,N_3939);
and U5758 (N_5758,N_2977,N_1301);
xnor U5759 (N_5759,N_4808,N_2829);
xor U5760 (N_5760,N_2639,N_1250);
and U5761 (N_5761,N_1160,N_2686);
xor U5762 (N_5762,N_2685,N_2316);
nor U5763 (N_5763,N_3945,N_2547);
nand U5764 (N_5764,N_1277,N_3789);
nand U5765 (N_5765,N_1602,N_4443);
xnor U5766 (N_5766,N_3021,N_3023);
nand U5767 (N_5767,N_2048,N_3550);
nor U5768 (N_5768,N_691,N_1008);
nor U5769 (N_5769,N_1402,N_4152);
and U5770 (N_5770,N_2027,N_1683);
and U5771 (N_5771,N_1514,N_726);
xor U5772 (N_5772,N_1464,N_3284);
or U5773 (N_5773,N_3378,N_3976);
nor U5774 (N_5774,N_407,N_2902);
nand U5775 (N_5775,N_3495,N_2000);
or U5776 (N_5776,N_1002,N_4099);
nand U5777 (N_5777,N_1924,N_2268);
nor U5778 (N_5778,N_14,N_2398);
or U5779 (N_5779,N_396,N_1290);
nor U5780 (N_5780,N_2905,N_1016);
nand U5781 (N_5781,N_342,N_1113);
and U5782 (N_5782,N_3403,N_3743);
or U5783 (N_5783,N_3690,N_738);
nand U5784 (N_5784,N_1832,N_31);
or U5785 (N_5785,N_3662,N_1652);
and U5786 (N_5786,N_3634,N_1667);
nand U5787 (N_5787,N_1168,N_4797);
xor U5788 (N_5788,N_3584,N_944);
and U5789 (N_5789,N_2657,N_655);
nor U5790 (N_5790,N_3684,N_1261);
nor U5791 (N_5791,N_2777,N_2195);
nand U5792 (N_5792,N_4390,N_2406);
nor U5793 (N_5793,N_2337,N_4998);
and U5794 (N_5794,N_590,N_3691);
or U5795 (N_5795,N_1534,N_4034);
nor U5796 (N_5796,N_3086,N_3702);
and U5797 (N_5797,N_4258,N_1440);
and U5798 (N_5798,N_1220,N_515);
nand U5799 (N_5799,N_539,N_3178);
nor U5800 (N_5800,N_3758,N_4322);
nand U5801 (N_5801,N_1081,N_4527);
nand U5802 (N_5802,N_2390,N_3668);
and U5803 (N_5803,N_2601,N_3428);
nand U5804 (N_5804,N_3391,N_3510);
nand U5805 (N_5805,N_4027,N_956);
and U5806 (N_5806,N_1795,N_1949);
or U5807 (N_5807,N_1410,N_4777);
and U5808 (N_5808,N_544,N_864);
or U5809 (N_5809,N_2979,N_1394);
and U5810 (N_5810,N_3689,N_1684);
nor U5811 (N_5811,N_4822,N_1938);
nand U5812 (N_5812,N_4980,N_1010);
and U5813 (N_5813,N_1186,N_2489);
nor U5814 (N_5814,N_3604,N_3714);
nor U5815 (N_5815,N_2184,N_3824);
or U5816 (N_5816,N_1492,N_4306);
nand U5817 (N_5817,N_4365,N_1954);
xor U5818 (N_5818,N_3337,N_3018);
nor U5819 (N_5819,N_3808,N_3048);
and U5820 (N_5820,N_502,N_2816);
and U5821 (N_5821,N_2790,N_104);
and U5822 (N_5822,N_2511,N_4949);
nor U5823 (N_5823,N_1584,N_4738);
xor U5824 (N_5824,N_3259,N_1653);
nand U5825 (N_5825,N_4549,N_1940);
nor U5826 (N_5826,N_3348,N_4384);
and U5827 (N_5827,N_3177,N_2026);
xor U5828 (N_5828,N_2826,N_2581);
and U5829 (N_5829,N_3639,N_4375);
nand U5830 (N_5830,N_2301,N_4609);
or U5831 (N_5831,N_4356,N_3563);
and U5832 (N_5832,N_4702,N_4148);
and U5833 (N_5833,N_1280,N_249);
or U5834 (N_5834,N_961,N_3372);
xnor U5835 (N_5835,N_1105,N_4135);
and U5836 (N_5836,N_1712,N_3996);
nor U5837 (N_5837,N_1845,N_2062);
or U5838 (N_5838,N_2637,N_448);
or U5839 (N_5839,N_1713,N_831);
or U5840 (N_5840,N_4776,N_518);
nand U5841 (N_5841,N_191,N_4595);
and U5842 (N_5842,N_319,N_4456);
and U5843 (N_5843,N_345,N_3472);
xor U5844 (N_5844,N_4092,N_2391);
nor U5845 (N_5845,N_2983,N_1227);
nor U5846 (N_5846,N_2933,N_1436);
nand U5847 (N_5847,N_651,N_3041);
nor U5848 (N_5848,N_213,N_3333);
and U5849 (N_5849,N_550,N_2645);
and U5850 (N_5850,N_3936,N_35);
and U5851 (N_5851,N_346,N_303);
or U5852 (N_5852,N_1252,N_4238);
or U5853 (N_5853,N_4419,N_1823);
nor U5854 (N_5854,N_2783,N_2952);
nor U5855 (N_5855,N_1591,N_4659);
nand U5856 (N_5856,N_2874,N_3166);
or U5857 (N_5857,N_3918,N_1177);
nor U5858 (N_5858,N_4508,N_4411);
and U5859 (N_5859,N_4222,N_4197);
and U5860 (N_5860,N_2597,N_3150);
nor U5861 (N_5861,N_1662,N_2846);
nor U5862 (N_5862,N_2187,N_907);
and U5863 (N_5863,N_2336,N_2260);
nor U5864 (N_5864,N_782,N_1076);
or U5865 (N_5865,N_4927,N_571);
and U5866 (N_5866,N_354,N_2850);
nor U5867 (N_5867,N_3388,N_4433);
or U5868 (N_5868,N_347,N_856);
nor U5869 (N_5869,N_3359,N_2024);
or U5870 (N_5870,N_4940,N_1426);
nand U5871 (N_5871,N_1365,N_2289);
nand U5872 (N_5872,N_2857,N_1654);
and U5873 (N_5873,N_4990,N_4679);
xnor U5874 (N_5874,N_4293,N_1864);
or U5875 (N_5875,N_2764,N_3612);
nand U5876 (N_5876,N_4678,N_3046);
nor U5877 (N_5877,N_1549,N_192);
xnor U5878 (N_5878,N_4625,N_2428);
nor U5879 (N_5879,N_739,N_2743);
or U5880 (N_5880,N_2471,N_439);
or U5881 (N_5881,N_2769,N_44);
nand U5882 (N_5882,N_4245,N_4596);
nand U5883 (N_5883,N_2456,N_911);
nand U5884 (N_5884,N_920,N_740);
or U5885 (N_5885,N_153,N_2823);
nand U5886 (N_5886,N_1878,N_3794);
nor U5887 (N_5887,N_4480,N_538);
xor U5888 (N_5888,N_1803,N_4857);
or U5889 (N_5889,N_2854,N_1132);
nand U5890 (N_5890,N_572,N_1769);
xor U5891 (N_5891,N_1813,N_4038);
and U5892 (N_5892,N_3136,N_4547);
and U5893 (N_5893,N_2881,N_4234);
xnor U5894 (N_5894,N_1070,N_4003);
nor U5895 (N_5895,N_3842,N_2170);
or U5896 (N_5896,N_2164,N_2404);
nand U5897 (N_5897,N_271,N_1914);
xor U5898 (N_5898,N_4798,N_2716);
and U5899 (N_5899,N_3664,N_65);
and U5900 (N_5900,N_2424,N_3896);
and U5901 (N_5901,N_3522,N_1362);
nand U5902 (N_5902,N_573,N_3508);
nor U5903 (N_5903,N_667,N_431);
or U5904 (N_5904,N_2407,N_4164);
nand U5905 (N_5905,N_4311,N_3717);
nor U5906 (N_5906,N_2818,N_4960);
and U5907 (N_5907,N_4816,N_1952);
nand U5908 (N_5908,N_3318,N_3697);
nand U5909 (N_5909,N_2508,N_2179);
and U5910 (N_5910,N_2778,N_126);
or U5911 (N_5911,N_4225,N_305);
nor U5912 (N_5912,N_1354,N_3577);
nand U5913 (N_5913,N_3037,N_3433);
xnor U5914 (N_5914,N_4151,N_4907);
nand U5915 (N_5915,N_4172,N_1953);
nand U5916 (N_5916,N_3067,N_3700);
nor U5917 (N_5917,N_4534,N_1892);
nand U5918 (N_5918,N_114,N_3883);
nand U5919 (N_5919,N_349,N_3481);
xor U5920 (N_5920,N_3157,N_3110);
nand U5921 (N_5921,N_4799,N_661);
nor U5922 (N_5922,N_619,N_4382);
nor U5923 (N_5923,N_3502,N_1503);
nor U5924 (N_5924,N_4651,N_4637);
xnor U5925 (N_5925,N_269,N_3647);
nor U5926 (N_5926,N_2518,N_4193);
nand U5927 (N_5927,N_2688,N_3500);
nand U5928 (N_5928,N_1999,N_1196);
or U5929 (N_5929,N_4716,N_1123);
nand U5930 (N_5930,N_1997,N_2389);
nand U5931 (N_5931,N_3127,N_1844);
xnor U5932 (N_5932,N_1345,N_2392);
and U5933 (N_5933,N_2174,N_4744);
nand U5934 (N_5934,N_2958,N_4062);
and U5935 (N_5935,N_1439,N_3557);
or U5936 (N_5936,N_3051,N_3453);
nand U5937 (N_5937,N_3860,N_3459);
xor U5938 (N_5938,N_1228,N_2076);
or U5939 (N_5939,N_3511,N_4978);
nor U5940 (N_5940,N_2776,N_1206);
or U5941 (N_5941,N_872,N_1639);
nor U5942 (N_5942,N_3980,N_777);
nand U5943 (N_5943,N_843,N_3139);
or U5944 (N_5944,N_2462,N_1052);
or U5945 (N_5945,N_2871,N_2445);
or U5946 (N_5946,N_2780,N_100);
nor U5947 (N_5947,N_4211,N_3633);
or U5948 (N_5948,N_4442,N_4464);
or U5949 (N_5949,N_1405,N_436);
nand U5950 (N_5950,N_3217,N_32);
and U5951 (N_5951,N_1249,N_2988);
and U5952 (N_5952,N_4139,N_688);
nor U5953 (N_5953,N_1802,N_4646);
xnor U5954 (N_5954,N_4498,N_3589);
or U5955 (N_5955,N_1032,N_3384);
or U5956 (N_5956,N_4693,N_1298);
and U5957 (N_5957,N_4396,N_3970);
nand U5958 (N_5958,N_1151,N_368);
xnor U5959 (N_5959,N_813,N_4212);
xor U5960 (N_5960,N_913,N_1929);
nand U5961 (N_5961,N_4605,N_4271);
and U5962 (N_5962,N_4570,N_2241);
or U5963 (N_5963,N_4237,N_4884);
and U5964 (N_5964,N_4846,N_3656);
nand U5965 (N_5965,N_1978,N_3329);
and U5966 (N_5966,N_3334,N_4444);
xnor U5967 (N_5967,N_2750,N_674);
and U5968 (N_5968,N_4157,N_2970);
or U5969 (N_5969,N_4368,N_2529);
nor U5970 (N_5970,N_1840,N_4513);
and U5971 (N_5971,N_3026,N_2711);
xor U5972 (N_5972,N_4766,N_1457);
and U5973 (N_5973,N_3411,N_2559);
and U5974 (N_5974,N_1817,N_2196);
and U5975 (N_5975,N_1594,N_1230);
or U5976 (N_5976,N_962,N_1414);
nor U5977 (N_5977,N_2418,N_4810);
and U5978 (N_5978,N_4581,N_4804);
nor U5979 (N_5979,N_4835,N_3097);
nor U5980 (N_5980,N_2612,N_2163);
or U5981 (N_5981,N_1303,N_687);
nor U5982 (N_5982,N_1812,N_2698);
nand U5983 (N_5983,N_4791,N_335);
xnor U5984 (N_5984,N_930,N_4778);
or U5985 (N_5985,N_3769,N_1475);
and U5986 (N_5986,N_3020,N_1518);
nand U5987 (N_5987,N_2224,N_54);
nor U5988 (N_5988,N_493,N_4674);
and U5989 (N_5989,N_2825,N_4886);
nand U5990 (N_5990,N_527,N_543);
or U5991 (N_5991,N_4961,N_401);
or U5992 (N_5992,N_242,N_4183);
nor U5993 (N_5993,N_2146,N_2673);
nand U5994 (N_5994,N_4364,N_1761);
and U5995 (N_5995,N_785,N_3269);
xor U5996 (N_5996,N_2441,N_4708);
and U5997 (N_5997,N_950,N_2641);
xor U5998 (N_5998,N_2175,N_1470);
nor U5999 (N_5999,N_2578,N_3140);
nand U6000 (N_6000,N_279,N_2436);
nor U6001 (N_6001,N_593,N_132);
and U6002 (N_6002,N_4658,N_2382);
nor U6003 (N_6003,N_4945,N_987);
nor U6004 (N_6004,N_2307,N_3745);
xor U6005 (N_6005,N_3362,N_402);
and U6006 (N_6006,N_123,N_3130);
nand U6007 (N_6007,N_2346,N_3434);
nor U6008 (N_6008,N_512,N_3394);
or U6009 (N_6009,N_4400,N_1642);
and U6010 (N_6010,N_3652,N_1927);
and U6011 (N_6011,N_4414,N_2452);
or U6012 (N_6012,N_2206,N_1236);
nor U6013 (N_6013,N_2364,N_1266);
xnor U6014 (N_6014,N_266,N_2538);
nand U6015 (N_6015,N_1092,N_1175);
and U6016 (N_6016,N_1663,N_1409);
xnor U6017 (N_6017,N_3952,N_1600);
or U6018 (N_6018,N_1278,N_1006);
nor U6019 (N_6019,N_1061,N_414);
nor U6020 (N_6020,N_2014,N_1396);
xnor U6021 (N_6021,N_442,N_3246);
nor U6022 (N_6022,N_4115,N_3304);
nand U6023 (N_6023,N_2330,N_4346);
and U6024 (N_6024,N_765,N_3820);
nor U6025 (N_6025,N_4491,N_1885);
or U6026 (N_6026,N_3653,N_2618);
and U6027 (N_6027,N_67,N_2763);
and U6028 (N_6028,N_2910,N_1605);
nand U6029 (N_6029,N_170,N_1592);
or U6030 (N_6030,N_3089,N_3516);
and U6031 (N_6031,N_2532,N_1012);
or U6032 (N_6032,N_3819,N_496);
nor U6033 (N_6033,N_551,N_2066);
nor U6034 (N_6034,N_1026,N_3382);
and U6035 (N_6035,N_748,N_1631);
nor U6036 (N_6036,N_566,N_4031);
or U6037 (N_6037,N_742,N_4251);
nor U6038 (N_6038,N_1702,N_449);
xor U6039 (N_6039,N_4201,N_3881);
and U6040 (N_6040,N_490,N_2143);
nand U6041 (N_6041,N_4149,N_2687);
nor U6042 (N_6042,N_3043,N_3250);
nand U6043 (N_6043,N_337,N_474);
nor U6044 (N_6044,N_4685,N_839);
nand U6045 (N_6045,N_1158,N_262);
xnor U6046 (N_6046,N_1072,N_3222);
nand U6047 (N_6047,N_1636,N_1289);
nor U6048 (N_6048,N_1797,N_1305);
nor U6049 (N_6049,N_162,N_4134);
xor U6050 (N_6050,N_1983,N_3228);
and U6051 (N_6051,N_1913,N_3621);
and U6052 (N_6052,N_2394,N_3376);
and U6053 (N_6053,N_372,N_427);
nand U6054 (N_6054,N_3665,N_3985);
and U6055 (N_6055,N_2317,N_2138);
nand U6056 (N_6056,N_3607,N_2128);
and U6057 (N_6057,N_881,N_578);
nand U6058 (N_6058,N_311,N_1229);
or U6059 (N_6059,N_594,N_579);
or U6060 (N_6060,N_4012,N_3438);
xor U6061 (N_6061,N_4606,N_2836);
nor U6062 (N_6062,N_3405,N_1917);
nand U6063 (N_6063,N_2834,N_1533);
and U6064 (N_6064,N_574,N_3943);
or U6065 (N_6065,N_4086,N_1771);
and U6066 (N_6066,N_4868,N_663);
and U6067 (N_6067,N_4820,N_4179);
and U6068 (N_6068,N_3628,N_4441);
xnor U6069 (N_6069,N_1171,N_4117);
and U6070 (N_6070,N_4654,N_4746);
nor U6071 (N_6071,N_638,N_817);
nor U6072 (N_6072,N_4102,N_3390);
nor U6073 (N_6073,N_4260,N_2285);
and U6074 (N_6074,N_2654,N_426);
or U6075 (N_6075,N_4889,N_822);
xnor U6076 (N_6076,N_1311,N_4964);
nand U6077 (N_6077,N_3599,N_3407);
nor U6078 (N_6078,N_1295,N_2084);
nand U6079 (N_6079,N_2296,N_2320);
and U6080 (N_6080,N_2941,N_1256);
or U6081 (N_6081,N_469,N_3942);
nand U6082 (N_6082,N_3540,N_2799);
nor U6083 (N_6083,N_293,N_4413);
and U6084 (N_6084,N_174,N_4137);
xor U6085 (N_6085,N_2675,N_4893);
nand U6086 (N_6086,N_3914,N_2357);
and U6087 (N_6087,N_2693,N_4950);
and U6088 (N_6088,N_2183,N_211);
and U6089 (N_6089,N_3395,N_3811);
nor U6090 (N_6090,N_4546,N_1730);
or U6091 (N_6091,N_2756,N_4830);
nand U6092 (N_6092,N_2788,N_1506);
nand U6093 (N_6093,N_3281,N_2701);
nor U6094 (N_6094,N_4826,N_2526);
nand U6095 (N_6095,N_2652,N_2993);
nand U6096 (N_6096,N_1352,N_1306);
nor U6097 (N_6097,N_154,N_4636);
nor U6098 (N_6098,N_3638,N_1299);
nor U6099 (N_6099,N_1276,N_2517);
or U6100 (N_6100,N_552,N_22);
xnor U6101 (N_6101,N_4370,N_2223);
nor U6102 (N_6102,N_3720,N_4100);
or U6103 (N_6103,N_4208,N_3884);
xor U6104 (N_6104,N_1649,N_176);
nand U6105 (N_6105,N_2551,N_2165);
nor U6106 (N_6106,N_27,N_3264);
and U6107 (N_6107,N_4565,N_325);
or U6108 (N_6108,N_1368,N_4008);
and U6109 (N_6109,N_4163,N_2400);
nor U6110 (N_6110,N_662,N_1147);
xnor U6111 (N_6111,N_3669,N_3408);
and U6112 (N_6112,N_4274,N_4610);
nand U6113 (N_6113,N_3252,N_2246);
nand U6114 (N_6114,N_3009,N_4993);
nand U6115 (N_6115,N_746,N_301);
or U6116 (N_6116,N_3841,N_910);
nor U6117 (N_6117,N_508,N_823);
nor U6118 (N_6118,N_3241,N_2208);
or U6119 (N_6119,N_925,N_1540);
nand U6120 (N_6120,N_3167,N_996);
xor U6121 (N_6121,N_1555,N_1839);
and U6122 (N_6122,N_3571,N_4624);
xnor U6123 (N_6123,N_732,N_3924);
and U6124 (N_6124,N_2283,N_2791);
or U6125 (N_6125,N_2863,N_2806);
xor U6126 (N_6126,N_1285,N_1473);
or U6127 (N_6127,N_635,N_1356);
nand U6128 (N_6128,N_2861,N_4267);
nand U6129 (N_6129,N_4004,N_33);
nand U6130 (N_6130,N_1547,N_4526);
nor U6131 (N_6131,N_2144,N_323);
nand U6132 (N_6132,N_848,N_4430);
and U6133 (N_6133,N_1060,N_2640);
nand U6134 (N_6134,N_4410,N_1382);
nor U6135 (N_6135,N_3323,N_2963);
nand U6136 (N_6136,N_3169,N_3444);
nor U6137 (N_6137,N_3866,N_3421);
nor U6138 (N_6138,N_656,N_1574);
xnor U6139 (N_6139,N_3189,N_441);
and U6140 (N_6140,N_3404,N_2600);
or U6141 (N_6141,N_1650,N_241);
nor U6142 (N_6142,N_2591,N_1934);
and U6143 (N_6143,N_2496,N_4355);
and U6144 (N_6144,N_664,N_1330);
nand U6145 (N_6145,N_816,N_3239);
nand U6146 (N_6146,N_2887,N_2740);
nand U6147 (N_6147,N_3785,N_1117);
xor U6148 (N_6148,N_2426,N_1738);
and U6149 (N_6149,N_3904,N_532);
nand U6150 (N_6150,N_3893,N_4262);
and U6151 (N_6151,N_1353,N_1038);
nand U6152 (N_6152,N_4663,N_2495);
and U6153 (N_6153,N_18,N_582);
and U6154 (N_6154,N_2996,N_1804);
nand U6155 (N_6155,N_4662,N_308);
or U6156 (N_6156,N_521,N_4294);
nor U6157 (N_6157,N_3449,N_2408);
and U6158 (N_6158,N_4123,N_4524);
or U6159 (N_6159,N_3988,N_4617);
nor U6160 (N_6160,N_4767,N_4316);
and U6161 (N_6161,N_69,N_2819);
and U6162 (N_6162,N_2016,N_2737);
xor U6163 (N_6163,N_81,N_4055);
nor U6164 (N_6164,N_1762,N_4072);
and U6165 (N_6165,N_3306,N_1442);
or U6166 (N_6166,N_937,N_4471);
nand U6167 (N_6167,N_1900,N_2022);
and U6168 (N_6168,N_970,N_2326);
nand U6169 (N_6169,N_1182,N_2893);
or U6170 (N_6170,N_1634,N_2625);
nor U6171 (N_6171,N_3958,N_1358);
nor U6172 (N_6172,N_417,N_318);
nor U6173 (N_6173,N_3316,N_889);
xor U6174 (N_6174,N_2381,N_2892);
and U6175 (N_6175,N_1719,N_3287);
nor U6176 (N_6176,N_545,N_385);
nor U6177 (N_6177,N_4705,N_1013);
and U6178 (N_6178,N_420,N_234);
nor U6179 (N_6179,N_2904,N_3324);
or U6180 (N_6180,N_4552,N_3226);
nand U6181 (N_6181,N_4376,N_361);
xnor U6182 (N_6182,N_2658,N_404);
and U6183 (N_6183,N_1563,N_878);
nand U6184 (N_6184,N_2287,N_322);
nor U6185 (N_6185,N_3258,N_1787);
or U6186 (N_6186,N_2606,N_2298);
and U6187 (N_6187,N_3016,N_3469);
or U6188 (N_6188,N_3328,N_3900);
nand U6189 (N_6189,N_2275,N_1260);
and U6190 (N_6190,N_3695,N_4848);
xnor U6191 (N_6191,N_4607,N_4423);
and U6192 (N_6192,N_2229,N_138);
and U6193 (N_6193,N_4140,N_4579);
nand U6194 (N_6194,N_853,N_3195);
or U6195 (N_6195,N_2443,N_4047);
nand U6196 (N_6196,N_3402,N_4493);
and U6197 (N_6197,N_4403,N_3132);
nand U6198 (N_6198,N_2805,N_2703);
nor U6199 (N_6199,N_1465,N_1496);
nand U6200 (N_6200,N_306,N_2264);
nor U6201 (N_6201,N_1047,N_985);
or U6202 (N_6202,N_2729,N_2216);
nand U6203 (N_6203,N_3161,N_1391);
nand U6204 (N_6204,N_3417,N_2784);
or U6205 (N_6205,N_3013,N_2957);
nand U6206 (N_6206,N_1853,N_1388);
xor U6207 (N_6207,N_4205,N_767);
and U6208 (N_6208,N_3266,N_4303);
xor U6209 (N_6209,N_194,N_1320);
or U6210 (N_6210,N_4358,N_608);
xor U6211 (N_6211,N_3661,N_3260);
or U6212 (N_6212,N_4792,N_2294);
or U6213 (N_6213,N_2752,N_3738);
xnor U6214 (N_6214,N_3944,N_2519);
or U6215 (N_6215,N_904,N_3921);
and U6216 (N_6216,N_4944,N_1831);
nor U6217 (N_6217,N_338,N_1778);
and U6218 (N_6218,N_1095,N_316);
and U6219 (N_6219,N_3517,N_1193);
nand U6220 (N_6220,N_362,N_344);
xor U6221 (N_6221,N_2617,N_2942);
nand U6222 (N_6222,N_334,N_1329);
nand U6223 (N_6223,N_2097,N_2781);
or U6224 (N_6224,N_3346,N_1686);
or U6225 (N_6225,N_403,N_1477);
nor U6226 (N_6226,N_1881,N_3949);
or U6227 (N_6227,N_820,N_2843);
nand U6228 (N_6228,N_328,N_1286);
nand U6229 (N_6229,N_3567,N_4875);
nand U6230 (N_6230,N_4593,N_815);
and U6231 (N_6231,N_1628,N_2205);
or U6232 (N_6232,N_2189,N_1225);
or U6233 (N_6233,N_616,N_4771);
nand U6234 (N_6234,N_4601,N_3728);
nand U6235 (N_6235,N_400,N_3614);
nor U6236 (N_6236,N_3753,N_2132);
nand U6237 (N_6237,N_204,N_1703);
nor U6238 (N_6238,N_4970,N_3566);
nand U6239 (N_6239,N_753,N_160);
nand U6240 (N_6240,N_4203,N_973);
and U6241 (N_6241,N_4703,N_1669);
nor U6242 (N_6242,N_4075,N_2340);
nand U6243 (N_6243,N_2546,N_3369);
nor U6244 (N_6244,N_1254,N_4301);
nor U6245 (N_6245,N_1051,N_3244);
nand U6246 (N_6246,N_3082,N_1173);
xnor U6247 (N_6247,N_4341,N_2557);
or U6248 (N_6248,N_3905,N_1859);
nor U6249 (N_6249,N_729,N_863);
and U6250 (N_6250,N_587,N_2945);
or U6251 (N_6251,N_1039,N_1734);
nand U6252 (N_6252,N_4101,N_832);
xnor U6253 (N_6253,N_4516,N_4780);
and U6254 (N_6254,N_1883,N_3466);
or U6255 (N_6255,N_2803,N_1972);
or U6256 (N_6256,N_3625,N_2420);
nor U6257 (N_6257,N_1317,N_644);
nor U6258 (N_6258,N_1848,N_4125);
and U6259 (N_6259,N_3381,N_3450);
nand U6260 (N_6260,N_2745,N_4485);
and U6261 (N_6261,N_4634,N_4295);
nand U6262 (N_6262,N_3597,N_516);
or U6263 (N_6263,N_30,N_2989);
and U6264 (N_6264,N_4760,N_2332);
and U6265 (N_6265,N_615,N_1456);
and U6266 (N_6266,N_4885,N_4911);
and U6267 (N_6267,N_2651,N_3283);
xnor U6268 (N_6268,N_3888,N_2707);
or U6269 (N_6269,N_4825,N_3663);
xnor U6270 (N_6270,N_1307,N_1194);
xnor U6271 (N_6271,N_3713,N_80);
xnor U6272 (N_6272,N_774,N_3120);
nand U6273 (N_6273,N_2405,N_636);
nand U6274 (N_6274,N_129,N_2506);
or U6275 (N_6275,N_3061,N_4867);
and U6276 (N_6276,N_172,N_1384);
and U6277 (N_6277,N_3797,N_4026);
nor U6278 (N_6278,N_1854,N_2722);
xnor U6279 (N_6279,N_706,N_4503);
xnor U6280 (N_6280,N_1750,N_1041);
and U6281 (N_6281,N_4592,N_3962);
nand U6282 (N_6282,N_1964,N_1150);
and U6283 (N_6283,N_4321,N_4367);
and U6284 (N_6284,N_595,N_2644);
xor U6285 (N_6285,N_1127,N_4081);
nand U6286 (N_6286,N_282,N_988);
and U6287 (N_6287,N_4361,N_3536);
nand U6288 (N_6288,N_759,N_627);
and U6289 (N_6289,N_2660,N_1135);
and U6290 (N_6290,N_678,N_4428);
or U6291 (N_6291,N_3615,N_4969);
nor U6292 (N_6292,N_36,N_3422);
nor U6293 (N_6293,N_4630,N_185);
or U6294 (N_6294,N_2369,N_1046);
and U6295 (N_6295,N_4807,N_2388);
nand U6296 (N_6296,N_4097,N_890);
xnor U6297 (N_6297,N_34,N_4902);
nor U6298 (N_6298,N_3818,N_2938);
and U6299 (N_6299,N_310,N_3971);
and U6300 (N_6300,N_4020,N_1077);
nor U6301 (N_6301,N_1283,N_2464);
and U6302 (N_6302,N_3118,N_4313);
and U6303 (N_6303,N_3572,N_307);
xnor U6304 (N_6304,N_4221,N_1635);
nand U6305 (N_6305,N_2136,N_4106);
and U6306 (N_6306,N_4432,N_376);
nor U6307 (N_6307,N_3928,N_2708);
nor U6308 (N_6308,N_4119,N_4578);
nor U6309 (N_6309,N_3863,N_1529);
xnor U6310 (N_6310,N_4795,N_2194);
nor U6311 (N_6311,N_829,N_3101);
and U6312 (N_6312,N_1931,N_3298);
and U6313 (N_6313,N_2222,N_1847);
and U6314 (N_6314,N_1984,N_990);
xnor U6315 (N_6315,N_2930,N_3103);
nand U6316 (N_6316,N_2007,N_1495);
nor U6317 (N_6317,N_4852,N_1623);
nor U6318 (N_6318,N_668,N_4854);
xnor U6319 (N_6319,N_3813,N_626);
nand U6320 (N_6320,N_1003,N_1993);
and U6321 (N_6321,N_1675,N_4723);
nand U6322 (N_6322,N_1950,N_4675);
nor U6323 (N_6323,N_3229,N_3336);
nor U6324 (N_6324,N_2735,N_1497);
and U6325 (N_6325,N_2859,N_2730);
nand U6326 (N_6326,N_3802,N_4283);
nor U6327 (N_6327,N_3916,N_775);
nand U6328 (N_6328,N_2249,N_2379);
xnor U6329 (N_6329,N_2157,N_139);
nand U6330 (N_6330,N_2034,N_1798);
or U6331 (N_6331,N_289,N_460);
and U6332 (N_6332,N_3042,N_38);
nand U6333 (N_6333,N_1007,N_4923);
nor U6334 (N_6334,N_2974,N_2595);
nand U6335 (N_6335,N_4717,N_4559);
nand U6336 (N_6336,N_3296,N_3501);
nor U6337 (N_6337,N_3772,N_1359);
nor U6338 (N_6338,N_3957,N_1185);
nand U6339 (N_6339,N_2713,N_2544);
or U6340 (N_6340,N_1671,N_2311);
nand U6341 (N_6341,N_764,N_2411);
or U6342 (N_6342,N_3655,N_3681);
nor U6343 (N_6343,N_77,N_2804);
nand U6344 (N_6344,N_1102,N_2017);
nand U6345 (N_6345,N_4289,N_2571);
or U6346 (N_6346,N_918,N_3057);
or U6347 (N_6347,N_112,N_40);
nor U6348 (N_6348,N_2760,N_2105);
and U6349 (N_6349,N_1696,N_946);
and U6350 (N_6350,N_530,N_1570);
nor U6351 (N_6351,N_2944,N_4351);
and U6352 (N_6352,N_1665,N_4040);
and U6353 (N_6353,N_3966,N_810);
and U6354 (N_6354,N_3674,N_2643);
and U6355 (N_6355,N_4387,N_800);
xor U6356 (N_6356,N_4431,N_458);
nand U6357 (N_6357,N_520,N_430);
and U6358 (N_6358,N_1443,N_1415);
nor U6359 (N_6359,N_1554,N_2186);
nor U6360 (N_6360,N_3377,N_3458);
or U6361 (N_6361,N_3897,N_4420);
nand U6362 (N_6362,N_3576,N_3969);
nand U6363 (N_6363,N_3686,N_641);
and U6364 (N_6364,N_4474,N_3644);
or U6365 (N_6365,N_1258,N_1327);
and U6366 (N_6366,N_4270,N_2484);
xor U6367 (N_6367,N_2661,N_720);
and U6368 (N_6368,N_1167,N_4309);
nand U6369 (N_6369,N_215,N_1615);
nand U6370 (N_6370,N_2573,N_4909);
or U6371 (N_6371,N_4334,N_4555);
and U6372 (N_6372,N_1643,N_2221);
or U6373 (N_6373,N_4888,N_63);
xor U6374 (N_6374,N_408,N_2603);
nor U6375 (N_6375,N_922,N_4599);
nor U6376 (N_6376,N_253,N_4901);
or U6377 (N_6377,N_3291,N_1585);
or U6378 (N_6378,N_4383,N_4215);
xor U6379 (N_6379,N_1920,N_4288);
and U6380 (N_6380,N_4583,N_4922);
or U6381 (N_6381,N_1967,N_4836);
and U6382 (N_6382,N_3467,N_2454);
or U6383 (N_6383,N_4536,N_2543);
nand U6384 (N_6384,N_3838,N_1886);
nor U6385 (N_6385,N_3915,N_1674);
xor U6386 (N_6386,N_4200,N_3370);
nand U6387 (N_6387,N_3087,N_1871);
and U6388 (N_6388,N_2720,N_1369);
or U6389 (N_6389,N_1505,N_2565);
or U6390 (N_6390,N_743,N_1772);
or U6391 (N_6391,N_4817,N_2982);
nand U6392 (N_6392,N_1687,N_1919);
nand U6393 (N_6393,N_4824,N_3274);
or U6394 (N_6394,N_1078,N_2447);
nor U6395 (N_6395,N_955,N_4427);
and U6396 (N_6396,N_3675,N_3448);
nor U6397 (N_6397,N_1062,N_3151);
nor U6398 (N_6398,N_3084,N_2742);
or U6399 (N_6399,N_1253,N_4371);
or U6400 (N_6400,N_1715,N_2254);
nor U6401 (N_6401,N_2091,N_4577);
or U6402 (N_6402,N_1408,N_2453);
or U6403 (N_6403,N_3878,N_1957);
nor U6404 (N_6404,N_4968,N_3138);
or U6405 (N_6405,N_4837,N_1466);
nor U6406 (N_6406,N_4347,N_4342);
xnor U6407 (N_6407,N_4540,N_666);
nor U6408 (N_6408,N_1589,N_1781);
nand U6409 (N_6409,N_2909,N_564);
nand U6410 (N_6410,N_2458,N_2906);
xnor U6411 (N_6411,N_4866,N_2501);
nor U6412 (N_6412,N_4074,N_840);
and U6413 (N_6413,N_3546,N_1909);
nor U6414 (N_6414,N_2541,N_4892);
nor U6415 (N_6415,N_1724,N_769);
nand U6416 (N_6416,N_4024,N_4898);
xnor U6417 (N_6417,N_2355,N_722);
or U6418 (N_6418,N_73,N_1156);
or U6419 (N_6419,N_967,N_4735);
nand U6420 (N_6420,N_4557,N_2994);
or U6421 (N_6421,N_1765,N_1965);
or U6422 (N_6422,N_1165,N_297);
or U6423 (N_6423,N_4220,N_3354);
and U6424 (N_6424,N_410,N_4169);
or U6425 (N_6425,N_1248,N_3268);
nand U6426 (N_6426,N_3537,N_2470);
nor U6427 (N_6427,N_2598,N_2088);
or U6428 (N_6428,N_1908,N_1103);
nor U6429 (N_6429,N_1073,N_1728);
and U6430 (N_6430,N_3331,N_359);
or U6431 (N_6431,N_25,N_152);
and U6432 (N_6432,N_2305,N_168);
nand U6433 (N_6433,N_1120,N_4429);
or U6434 (N_6434,N_453,N_2218);
xor U6435 (N_6435,N_3040,N_4523);
nor U6436 (N_6436,N_1049,N_852);
nor U6437 (N_6437,N_1904,N_373);
and U6438 (N_6438,N_1764,N_4243);
or U6439 (N_6439,N_3920,N_1606);
and U6440 (N_6440,N_3671,N_914);
nor U6441 (N_6441,N_3425,N_4021);
xor U6442 (N_6442,N_1187,N_4528);
and U6443 (N_6443,N_2031,N_4336);
and U6444 (N_6444,N_4874,N_4751);
and U6445 (N_6445,N_3413,N_1383);
or U6446 (N_6446,N_2348,N_3631);
nand U6447 (N_6447,N_4511,N_3030);
xnor U6448 (N_6448,N_1445,N_4986);
xor U6449 (N_6449,N_3133,N_3482);
xnor U6450 (N_6450,N_3154,N_3104);
and U6451 (N_6451,N_3935,N_4252);
and U6452 (N_6452,N_1948,N_3090);
nor U6453 (N_6453,N_1603,N_2324);
nand U6454 (N_6454,N_2288,N_1799);
and U6455 (N_6455,N_624,N_64);
nor U6456 (N_6456,N_2162,N_1918);
nand U6457 (N_6457,N_4782,N_4714);
and U6458 (N_6458,N_836,N_4405);
and U6459 (N_6459,N_124,N_2875);
and U6460 (N_6460,N_217,N_2150);
nand U6461 (N_6461,N_2590,N_3117);
nor U6462 (N_6462,N_4246,N_3234);
nor U6463 (N_6463,N_3938,N_2429);
nand U6464 (N_6464,N_4881,N_2093);
nor U6465 (N_6465,N_2897,N_3198);
nand U6466 (N_6466,N_4089,N_1557);
or U6467 (N_6467,N_299,N_1898);
nand U6468 (N_6468,N_4522,N_4517);
or U6469 (N_6469,N_381,N_905);
nor U6470 (N_6470,N_3355,N_701);
nand U6471 (N_6471,N_3814,N_2168);
xor U6472 (N_6472,N_4512,N_2692);
or U6473 (N_6473,N_3286,N_4550);
nor U6474 (N_6474,N_391,N_4535);
nor U6475 (N_6475,N_2474,N_1421);
and U6476 (N_6476,N_4264,N_435);
and U6477 (N_6477,N_1779,N_4412);
or U6478 (N_6478,N_2367,N_495);
nand U6479 (N_6479,N_1423,N_413);
nor U6480 (N_6480,N_2444,N_140);
and U6481 (N_6481,N_2166,N_1876);
and U6482 (N_6482,N_2891,N_504);
nand U6483 (N_6483,N_2497,N_4992);
or U6484 (N_6484,N_2894,N_60);
nor U6485 (N_6485,N_3739,N_2455);
nand U6486 (N_6486,N_3947,N_1462);
nand U6487 (N_6487,N_4773,N_4975);
nand U6488 (N_6488,N_4844,N_4495);
and U6489 (N_6489,N_3518,N_226);
nor U6490 (N_6490,N_1274,N_4603);
or U6491 (N_6491,N_908,N_1048);
nand U6492 (N_6492,N_2038,N_2036);
nand U6493 (N_6493,N_1491,N_2680);
nor U6494 (N_6494,N_3205,N_4340);
nand U6495 (N_6495,N_581,N_2749);
and U6496 (N_6496,N_586,N_2350);
and U6497 (N_6497,N_4080,N_3999);
and U6498 (N_6498,N_2966,N_4398);
and U6499 (N_6499,N_1743,N_4505);
nand U6500 (N_6500,N_4127,N_3912);
or U6501 (N_6501,N_4118,N_4821);
nor U6502 (N_6502,N_3602,N_1232);
or U6503 (N_6503,N_3214,N_1785);
and U6504 (N_6504,N_1080,N_724);
nor U6505 (N_6505,N_694,N_2880);
xor U6506 (N_6506,N_981,N_3113);
and U6507 (N_6507,N_3780,N_85);
nor U6508 (N_6508,N_979,N_1403);
or U6509 (N_6509,N_1735,N_1205);
nor U6510 (N_6510,N_2576,N_1333);
nor U6511 (N_6511,N_2808,N_2480);
and U6512 (N_6512,N_673,N_3363);
nor U6513 (N_6513,N_3630,N_4006);
and U6514 (N_6514,N_216,N_680);
nor U6515 (N_6515,N_966,N_4644);
xnor U6516 (N_6516,N_1455,N_4538);
and U6517 (N_6517,N_1458,N_2665);
nor U6518 (N_6518,N_4145,N_149);
and U6519 (N_6519,N_1888,N_3248);
nor U6520 (N_6520,N_4823,N_3667);
or U6521 (N_6521,N_1172,N_3457);
nor U6522 (N_6522,N_478,N_2185);
or U6523 (N_6523,N_1397,N_1543);
nor U6524 (N_6524,N_4710,N_702);
or U6525 (N_6525,N_2466,N_1134);
and U6526 (N_6526,N_183,N_2378);
or U6527 (N_6527,N_2323,N_2412);
and U6528 (N_6528,N_1395,N_3361);
nand U6529 (N_6529,N_3446,N_3233);
nor U6530 (N_6530,N_2666,N_4492);
nand U6531 (N_6531,N_351,N_2065);
nor U6532 (N_6532,N_837,N_4185);
or U6533 (N_6533,N_1849,N_2542);
nand U6534 (N_6534,N_750,N_4472);
or U6535 (N_6535,N_3184,N_1998);
and U6536 (N_6536,N_3810,N_1390);
nor U6537 (N_6537,N_2028,N_3365);
xnor U6538 (N_6538,N_558,N_880);
and U6539 (N_6539,N_557,N_3587);
and U6540 (N_6540,N_3754,N_895);
nand U6541 (N_6541,N_2013,N_1166);
xnor U6542 (N_6542,N_1148,N_2888);
or U6543 (N_6543,N_709,N_4991);
or U6544 (N_6544,N_3740,N_1344);
xnor U6545 (N_6545,N_4752,N_1326);
nor U6546 (N_6546,N_3200,N_3998);
nand U6547 (N_6547,N_2734,N_1043);
nand U6548 (N_6548,N_2167,N_1791);
xor U6549 (N_6549,N_2386,N_3349);
or U6550 (N_6550,N_999,N_150);
or U6551 (N_6551,N_2003,N_2054);
xnor U6552 (N_6552,N_4161,N_2279);
and U6553 (N_6553,N_248,N_3982);
xnor U6554 (N_6554,N_4051,N_1644);
or U6555 (N_6555,N_3853,N_2916);
or U6556 (N_6556,N_1349,N_4897);
nand U6557 (N_6557,N_4972,N_2748);
or U6558 (N_6558,N_1235,N_315);
nand U6559 (N_6559,N_3218,N_4349);
and U6560 (N_6560,N_2636,N_763);
nand U6561 (N_6561,N_850,N_2684);
nor U6562 (N_6562,N_676,N_1014);
and U6563 (N_6563,N_1152,N_1545);
or U6564 (N_6564,N_1422,N_3431);
nand U6565 (N_6565,N_2499,N_2310);
or U6566 (N_6566,N_3010,N_830);
nand U6567 (N_6567,N_457,N_1796);
nand U6568 (N_6568,N_3078,N_2844);
nand U6569 (N_6569,N_1512,N_2995);
or U6570 (N_6570,N_121,N_4372);
nand U6571 (N_6571,N_3569,N_3977);
or U6572 (N_6572,N_844,N_3879);
xnor U6573 (N_6573,N_1677,N_1740);
nand U6574 (N_6574,N_4076,N_1241);
or U6575 (N_6575,N_1244,N_901);
nand U6576 (N_6576,N_1028,N_199);
nor U6577 (N_6577,N_3083,N_2869);
and U6578 (N_6578,N_721,N_2923);
and U6579 (N_6579,N_471,N_1446);
nor U6580 (N_6580,N_4757,N_1850);
or U6581 (N_6581,N_1074,N_1178);
nand U6582 (N_6582,N_133,N_2833);
nand U6583 (N_6583,N_2103,N_161);
nand U6584 (N_6584,N_4947,N_3340);
nand U6585 (N_6585,N_2676,N_3000);
nor U6586 (N_6586,N_205,N_4144);
or U6587 (N_6587,N_4677,N_2801);
and U6588 (N_6588,N_1435,N_2662);
nor U6589 (N_6589,N_4908,N_4195);
and U6590 (N_6590,N_288,N_2265);
nand U6591 (N_6591,N_2250,N_3171);
nor U6592 (N_6592,N_1536,N_3074);
or U6593 (N_6593,N_209,N_2361);
nor U6594 (N_6594,N_2130,N_2015);
or U6595 (N_6595,N_340,N_1922);
or U6596 (N_6596,N_884,N_237);
and U6597 (N_6597,N_3035,N_3864);
nand U6598 (N_6598,N_2907,N_2877);
and U6599 (N_6599,N_1130,N_4315);
xnor U6600 (N_6600,N_4912,N_1614);
or U6601 (N_6601,N_78,N_3007);
or U6602 (N_6602,N_3122,N_1222);
or U6603 (N_6603,N_787,N_4956);
or U6604 (N_6604,N_2575,N_4783);
or U6605 (N_6605,N_945,N_3001);
xnor U6606 (N_6606,N_2086,N_4141);
nor U6607 (N_6607,N_2583,N_240);
xor U6608 (N_6608,N_858,N_682);
nand U6609 (N_6609,N_232,N_1660);
nand U6610 (N_6610,N_1788,N_2154);
or U6611 (N_6611,N_3565,N_300);
and U6612 (N_6612,N_4533,N_280);
nand U6613 (N_6613,N_3827,N_500);
nand U6614 (N_6614,N_3795,N_1528);
nor U6615 (N_6615,N_795,N_4576);
nor U6616 (N_6616,N_4424,N_2672);
nor U6617 (N_6617,N_4190,N_228);
or U6618 (N_6618,N_3210,N_879);
nor U6619 (N_6619,N_2370,N_3426);
xnor U6620 (N_6620,N_2502,N_1297);
or U6621 (N_6621,N_974,N_2853);
and U6622 (N_6622,N_1203,N_3075);
nand U6623 (N_6623,N_3275,N_1621);
and U6624 (N_6624,N_4345,N_3645);
and U6625 (N_6625,N_3922,N_1691);
and U6626 (N_6626,N_643,N_1995);
nor U6627 (N_6627,N_3081,N_1969);
and U6628 (N_6628,N_2106,N_2924);
or U6629 (N_6629,N_2258,N_4487);
and U6630 (N_6630,N_4704,N_4787);
xor U6631 (N_6631,N_1424,N_281);
or U6632 (N_6632,N_3603,N_1140);
nand U6633 (N_6633,N_184,N_2089);
nor U6634 (N_6634,N_3771,N_3080);
xor U6635 (N_6635,N_3168,N_2920);
and U6636 (N_6636,N_4227,N_3439);
nor U6637 (N_6637,N_1846,N_4743);
and U6638 (N_6638,N_4381,N_4095);
and U6639 (N_6639,N_2810,N_419);
and U6640 (N_6640,N_2847,N_4502);
nand U6641 (N_6641,N_4392,N_2366);
nor U6642 (N_6642,N_95,N_3387);
nor U6643 (N_6643,N_3828,N_3762);
and U6644 (N_6644,N_2029,N_324);
nor U6645 (N_6645,N_2334,N_693);
nand U6646 (N_6646,N_3442,N_3515);
nor U6647 (N_6647,N_2071,N_992);
nand U6648 (N_6648,N_2521,N_2252);
and U6649 (N_6649,N_4611,N_1828);
nor U6650 (N_6650,N_4987,N_4827);
xnor U6651 (N_6651,N_3937,N_1027);
nand U6652 (N_6652,N_3271,N_2035);
xor U6653 (N_6653,N_4754,N_2396);
nand U6654 (N_6654,N_4711,N_2176);
xor U6655 (N_6655,N_1144,N_1974);
nand U6656 (N_6656,N_2393,N_1951);
or U6657 (N_6657,N_2111,N_4913);
and U6658 (N_6658,N_294,N_332);
nor U6659 (N_6659,N_2291,N_3420);
nor U6660 (N_6660,N_4633,N_20);
and U6661 (N_6661,N_4281,N_1444);
and U6662 (N_6662,N_3868,N_1083);
and U6663 (N_6663,N_4900,N_2021);
nor U6664 (N_6664,N_3094,N_1814);
nor U6665 (N_6665,N_4307,N_2180);
nor U6666 (N_6666,N_433,N_4462);
nand U6667 (N_6667,N_2090,N_4965);
or U6668 (N_6668,N_1857,N_4223);
or U6669 (N_6669,N_4589,N_4255);
or U6670 (N_6670,N_4404,N_3657);
nor U6671 (N_6671,N_3573,N_3525);
and U6672 (N_6672,N_1566,N_4036);
nor U6673 (N_6673,N_1689,N_1050);
xor U6674 (N_6674,N_2926,N_1115);
and U6675 (N_6675,N_2913,N_698);
or U6676 (N_6676,N_1268,N_4154);
nand U6677 (N_6677,N_1637,N_865);
xnor U6678 (N_6678,N_4494,N_1926);
or U6679 (N_6679,N_916,N_4686);
nand U6680 (N_6680,N_79,N_2718);
or U6681 (N_6681,N_929,N_4819);
xnor U6682 (N_6682,N_4602,N_1851);
xor U6683 (N_6683,N_2807,N_39);
and U6684 (N_6684,N_230,N_395);
or U6685 (N_6685,N_2133,N_3609);
nor U6686 (N_6686,N_3344,N_1233);
nand U6687 (N_6687,N_4249,N_3940);
and U6688 (N_6688,N_3070,N_2339);
nor U6689 (N_6689,N_4626,N_3379);
nor U6690 (N_6690,N_3091,N_857);
or U6691 (N_6691,N_118,N_535);
xnor U6692 (N_6692,N_2101,N_3849);
nand U6693 (N_6693,N_2153,N_4564);
nand U6694 (N_6694,N_728,N_1991);
or U6695 (N_6695,N_3598,N_1169);
nor U6696 (N_6696,N_1100,N_3816);
xor U6697 (N_6697,N_3165,N_1736);
or U6698 (N_6698,N_1291,N_2587);
nand U6699 (N_6699,N_3049,N_1246);
nor U6700 (N_6700,N_360,N_1109);
nor U6701 (N_6701,N_2193,N_1155);
nor U6702 (N_6702,N_3473,N_3724);
or U6703 (N_6703,N_2981,N_1873);
nor U6704 (N_6704,N_4805,N_524);
or U6705 (N_6705,N_42,N_2434);
nand U6706 (N_6706,N_3535,N_336);
or U6707 (N_6707,N_801,N_909);
xor U6708 (N_6708,N_3027,N_1561);
nor U6709 (N_6709,N_896,N_2259);
nand U6710 (N_6710,N_4758,N_1309);
nand U6711 (N_6711,N_1011,N_2004);
or U6712 (N_6712,N_4556,N_4088);
nor U6713 (N_6713,N_3987,N_4044);
nor U6714 (N_6714,N_1578,N_4300);
and U6715 (N_6715,N_4181,N_451);
nand U6716 (N_6716,N_3,N_3159);
nand U6717 (N_6717,N_554,N_2860);
and U6718 (N_6718,N_4954,N_1607);
or U6719 (N_6719,N_1055,N_1504);
nor U6720 (N_6720,N_4569,N_4244);
nand U6721 (N_6721,N_3651,N_1393);
and U6722 (N_6722,N_2129,N_860);
or U6723 (N_6723,N_1346,N_3679);
or U6724 (N_6724,N_2341,N_2931);
or U6725 (N_6725,N_717,N_4747);
or U6726 (N_6726,N_13,N_833);
nor U6727 (N_6727,N_3299,N_1731);
nor U6728 (N_6728,N_965,N_4580);
xor U6729 (N_6729,N_287,N_4259);
and U6730 (N_6730,N_1971,N_273);
or U6731 (N_6731,N_2139,N_1453);
nand U6732 (N_6732,N_4635,N_1657);
or U6733 (N_6733,N_2585,N_4388);
and U6734 (N_6734,N_2181,N_3858);
or U6735 (N_6735,N_1680,N_3931);
nand U6736 (N_6736,N_3755,N_1161);
xnor U6737 (N_6737,N_3967,N_3741);
nand U6738 (N_6738,N_3423,N_1721);
or U6739 (N_6739,N_629,N_4571);
nor U6740 (N_6740,N_4680,N_1323);
and U6741 (N_6741,N_2932,N_531);
and U6742 (N_6742,N_4110,N_1992);
and U6743 (N_6743,N_4302,N_4638);
or U6744 (N_6744,N_3135,N_3891);
nand U6745 (N_6745,N_1483,N_1841);
or U6746 (N_6746,N_4091,N_1560);
and U6747 (N_6747,N_2052,N_2262);
and U6748 (N_6748,N_1324,N_2120);
and U6749 (N_6749,N_2731,N_4109);
nand U6750 (N_6750,N_3941,N_3219);
nand U6751 (N_6751,N_2435,N_953);
or U6752 (N_6752,N_2550,N_295);
and U6753 (N_6753,N_3380,N_375);
nand U6754 (N_6754,N_2723,N_645);
nand U6755 (N_6755,N_2449,N_4847);
or U6756 (N_6756,N_3227,N_591);
nor U6757 (N_6757,N_76,N_4254);
and U6758 (N_6758,N_4468,N_2056);
nor U6759 (N_6759,N_2696,N_781);
and U6760 (N_6760,N_466,N_1897);
or U6761 (N_6761,N_928,N_505);
or U6762 (N_6762,N_3308,N_3352);
and U6763 (N_6763,N_3973,N_3528);
nand U6764 (N_6764,N_4981,N_751);
and U6765 (N_6765,N_2566,N_2338);
and U6766 (N_6766,N_3317,N_1733);
nand U6767 (N_6767,N_1377,N_3851);
xor U6768 (N_6768,N_2124,N_1855);
and U6769 (N_6769,N_1189,N_1500);
nand U6770 (N_6770,N_1875,N_529);
nor U6771 (N_6771,N_4001,N_1608);
or U6772 (N_6772,N_2172,N_465);
or U6773 (N_6773,N_1996,N_3983);
and U6774 (N_6774,N_4749,N_2524);
or U6775 (N_6775,N_252,N_1216);
and U6776 (N_6776,N_736,N_480);
or U6777 (N_6777,N_3209,N_3183);
and U6778 (N_6778,N_264,N_2473);
nor U6779 (N_6779,N_2839,N_353);
or U6780 (N_6780,N_4377,N_4018);
or U6781 (N_6781,N_957,N_3871);
and U6782 (N_6782,N_4250,N_320);
nor U6783 (N_6783,N_3415,N_3801);
nor U6784 (N_6784,N_1024,N_1537);
nand U6785 (N_6785,N_4369,N_2985);
or U6786 (N_6786,N_2293,N_2928);
nand U6787 (N_6787,N_4985,N_2020);
or U6788 (N_6788,N_2914,N_4272);
and U6789 (N_6789,N_2368,N_3488);
nand U6790 (N_6790,N_2946,N_4343);
or U6791 (N_6791,N_1468,N_752);
and U6792 (N_6792,N_3708,N_1784);
or U6793 (N_6793,N_4567,N_886);
nor U6794 (N_6794,N_2549,N_745);
xor U6795 (N_6795,N_2220,N_2092);
nand U6796 (N_6796,N_3533,N_3583);
nand U6797 (N_6797,N_2282,N_4841);
or U6798 (N_6798,N_2244,N_3005);
nand U6799 (N_6799,N_696,N_835);
xor U6800 (N_6800,N_1223,N_2409);
nand U6801 (N_6801,N_3855,N_4483);
or U6802 (N_6802,N_2509,N_4781);
or U6803 (N_6803,N_3290,N_2225);
and U6804 (N_6804,N_1912,N_1985);
and U6805 (N_6805,N_1498,N_1510);
or U6806 (N_6806,N_1355,N_932);
or U6807 (N_6807,N_3956,N_1746);
or U6808 (N_6808,N_2122,N_1595);
nand U6809 (N_6809,N_2286,N_3345);
or U6810 (N_6810,N_1775,N_1753);
or U6811 (N_6811,N_4925,N_339);
or U6812 (N_6812,N_1243,N_4041);
or U6813 (N_6813,N_1976,N_2947);
nand U6814 (N_6814,N_4437,N_2303);
nor U6815 (N_6815,N_4241,N_1418);
and U6816 (N_6816,N_4891,N_2536);
xor U6817 (N_6817,N_2118,N_1911);
nor U6818 (N_6818,N_1651,N_1211);
or U6819 (N_6819,N_1820,N_862);
nand U6820 (N_6820,N_298,N_4772);
nor U6821 (N_6821,N_621,N_4762);
or U6822 (N_6822,N_4806,N_2107);
nand U6823 (N_6823,N_1620,N_731);
or U6824 (N_6824,N_4719,N_3098);
and U6825 (N_6825,N_4142,N_994);
or U6826 (N_6826,N_4226,N_4248);
nor U6827 (N_6827,N_4890,N_3850);
nand U6828 (N_6828,N_3606,N_4037);
nand U6829 (N_6829,N_2604,N_1183);
or U6830 (N_6830,N_4085,N_3507);
nor U6831 (N_6831,N_3066,N_4664);
or U6832 (N_6832,N_3847,N_1693);
and U6833 (N_6833,N_4753,N_4532);
or U6834 (N_6834,N_1836,N_4083);
and U6835 (N_6835,N_370,N_3953);
xor U6836 (N_6836,N_304,N_4966);
nor U6837 (N_6837,N_1128,N_758);
nor U6838 (N_6838,N_1867,N_3992);
nor U6839 (N_6839,N_1709,N_467);
xnor U6840 (N_6840,N_68,N_2782);
nor U6841 (N_6841,N_995,N_3682);
nand U6842 (N_6842,N_4539,N_1023);
and U6843 (N_6843,N_3106,N_2794);
and U6844 (N_6844,N_4690,N_1079);
and U6845 (N_6845,N_1242,N_3358);
nand U6846 (N_6846,N_2171,N_2899);
or U6847 (N_6847,N_2401,N_2256);
nand U6848 (N_6848,N_1901,N_2005);
xnor U6849 (N_6849,N_2236,N_4138);
nand U6850 (N_6850,N_1874,N_2811);
or U6851 (N_6851,N_290,N_102);
and U6852 (N_6852,N_3131,N_4317);
and U6853 (N_6853,N_2137,N_1069);
nor U6854 (N_6854,N_3478,N_3660);
nand U6855 (N_6855,N_2709,N_3596);
nor U6856 (N_6856,N_2700,N_1891);
or U6857 (N_6857,N_3072,N_4065);
xnor U6858 (N_6858,N_1029,N_1486);
or U6859 (N_6859,N_4818,N_2754);
nor U6860 (N_6860,N_4275,N_873);
or U6861 (N_6861,N_2747,N_1025);
or U6862 (N_6862,N_3613,N_3068);
xnor U6863 (N_6863,N_3356,N_3804);
or U6864 (N_6864,N_3146,N_4882);
nand U6865 (N_6865,N_2712,N_1907);
and U6866 (N_6866,N_1861,N_2156);
nor U6867 (N_6867,N_2478,N_926);
and U6868 (N_6868,N_3991,N_343);
nand U6869 (N_6869,N_4887,N_3619);
nor U6870 (N_6870,N_2997,N_747);
nor U6871 (N_6871,N_3946,N_2009);
nor U6872 (N_6872,N_302,N_2953);
nor U6873 (N_6873,N_2099,N_547);
and U6874 (N_6874,N_3108,N_2371);
nor U6875 (N_6875,N_2779,N_770);
or U6876 (N_6876,N_1313,N_3986);
xnor U6877 (N_6877,N_3468,N_3730);
nand U6878 (N_6878,N_4668,N_1577);
nor U6879 (N_6879,N_4304,N_3093);
nand U6880 (N_6880,N_741,N_791);
and U6881 (N_6881,N_277,N_1564);
or U6882 (N_6882,N_2018,N_1507);
and U6883 (N_6883,N_3223,N_869);
nand U6884 (N_6884,N_2399,N_1184);
and U6885 (N_6885,N_4108,N_596);
or U6886 (N_6886,N_960,N_3105);
nand U6887 (N_6887,N_364,N_2430);
xor U6888 (N_6888,N_4839,N_2797);
xnor U6889 (N_6889,N_251,N_2739);
xnor U6890 (N_6890,N_4182,N_814);
and U6891 (N_6891,N_443,N_4518);
nor U6892 (N_6892,N_2921,N_4314);
and U6893 (N_6893,N_4672,N_1042);
nand U6894 (N_6894,N_3053,N_2354);
and U6895 (N_6895,N_2019,N_101);
nand U6896 (N_6896,N_3768,N_2064);
nand U6897 (N_6897,N_1915,N_1163);
nand U6898 (N_6898,N_1093,N_3622);
nor U6899 (N_6899,N_4575,N_653);
nor U6900 (N_6900,N_4,N_3282);
and U6901 (N_6901,N_10,N_4585);
xor U6902 (N_6902,N_4071,N_3531);
nand U6903 (N_6903,N_1508,N_2419);
or U6904 (N_6904,N_1739,N_712);
and U6905 (N_6905,N_2726,N_2949);
and U6906 (N_6906,N_3095,N_2245);
and U6907 (N_6907,N_4136,N_486);
or U6908 (N_6908,N_1977,N_4732);
or U6909 (N_6909,N_2900,N_4450);
and U6910 (N_6910,N_207,N_82);
nand U6911 (N_6911,N_3238,N_157);
nand U6912 (N_6912,N_4422,N_533);
or U6913 (N_6913,N_2642,N_546);
and U6914 (N_6914,N_4955,N_507);
xnor U6915 (N_6915,N_556,N_2884);
or U6916 (N_6916,N_3807,N_3643);
nor U6917 (N_6917,N_1217,N_4484);
or U6918 (N_6918,N_2214,N_623);
nor U6919 (N_6919,N_4273,N_560);
and U6920 (N_6920,N_941,N_3503);
xnor U6921 (N_6921,N_1343,N_3240);
nor U6922 (N_6922,N_2492,N_2158);
nor U6923 (N_6923,N_3427,N_313);
nor U6924 (N_6924,N_3570,N_1932);
nor U6925 (N_6925,N_4612,N_1541);
or U6926 (N_6926,N_3058,N_3701);
nand U6927 (N_6927,N_1065,N_2002);
and U6928 (N_6928,N_169,N_4851);
nor U6929 (N_6929,N_2113,N_4224);
and U6930 (N_6930,N_2315,N_3342);
and U6931 (N_6931,N_1794,N_2314);
or U6932 (N_6932,N_1364,N_2423);
or U6933 (N_6933,N_2273,N_2841);
or U6934 (N_6934,N_3368,N_776);
nor U6935 (N_6935,N_1022,N_2569);
and U6936 (N_6936,N_3911,N_3699);
and U6937 (N_6937,N_1417,N_4461);
and U6938 (N_6938,N_2045,N_1827);
nand U6939 (N_6939,N_358,N_866);
and U6940 (N_6940,N_3636,N_4853);
nand U6941 (N_6941,N_772,N_1962);
or U6942 (N_6942,N_660,N_3024);
or U6943 (N_6943,N_2063,N_125);
nor U6944 (N_6944,N_2646,N_1489);
nor U6945 (N_6945,N_4479,N_1618);
and U6946 (N_6946,N_549,N_744);
and U6947 (N_6947,N_1882,N_1114);
or U6948 (N_6948,N_4656,N_429);
and U6949 (N_6949,N_3440,N_2188);
nor U6950 (N_6950,N_3775,N_3102);
xor U6951 (N_6951,N_3121,N_2967);
or U6952 (N_6952,N_1251,N_1308);
nor U6953 (N_6953,N_2073,N_3836);
or U6954 (N_6954,N_1609,N_1499);
and U6955 (N_6955,N_2292,N_1782);
nand U6956 (N_6956,N_1568,N_1968);
and U6957 (N_6957,N_4860,N_761);
nand U6958 (N_6958,N_1255,N_978);
nor U6959 (N_6959,N_943,N_131);
nor U6960 (N_6960,N_3889,N_1304);
and U6961 (N_6961,N_4982,N_327);
or U6962 (N_6962,N_1860,N_4698);
nand U6963 (N_6963,N_2123,N_4218);
nand U6964 (N_6964,N_2689,N_348);
nor U6965 (N_6965,N_672,N_4768);
and U6966 (N_6966,N_1599,N_4470);
or U6967 (N_6967,N_3649,N_958);
nor U6968 (N_6968,N_1066,N_2155);
nor U6969 (N_6969,N_4718,N_4121);
nor U6970 (N_6970,N_3805,N_614);
and U6971 (N_6971,N_494,N_1379);
nor U6972 (N_6972,N_1829,N_1752);
nand U6973 (N_6973,N_919,N_2383);
xor U6974 (N_6974,N_4478,N_2257);
nor U6975 (N_6975,N_1742,N_4967);
nor U6976 (N_6976,N_4233,N_4409);
or U6977 (N_6977,N_2912,N_2943);
xor U6978 (N_6978,N_2487,N_1312);
nor U6979 (N_6979,N_2758,N_1966);
xnor U6980 (N_6980,N_3629,N_2670);
nand U6981 (N_6981,N_2006,N_3505);
nor U6982 (N_6982,N_4952,N_2773);
xnor U6983 (N_6983,N_1494,N_1180);
and U6984 (N_6984,N_3300,N_2659);
or U6985 (N_6985,N_3711,N_1994);
and U6986 (N_6986,N_2695,N_4007);
nor U6987 (N_6987,N_834,N_1033);
nand U6988 (N_6988,N_2049,N_2109);
nor U6989 (N_6989,N_4146,N_4305);
or U6990 (N_6990,N_1572,N_659);
or U6991 (N_6991,N_1629,N_4655);
nor U6992 (N_6992,N_4994,N_3616);
and U6993 (N_6993,N_4079,N_89);
or U6994 (N_6994,N_2589,N_3527);
nor U6995 (N_6995,N_4591,N_3798);
nor U6996 (N_6996,N_3149,N_2736);
or U6997 (N_6997,N_4050,N_2121);
xnor U6998 (N_6998,N_52,N_3704);
nor U6999 (N_6999,N_2809,N_53);
xnor U7000 (N_7000,N_1493,N_1818);
and U7001 (N_7001,N_657,N_1110);
nor U7002 (N_7002,N_2215,N_906);
and U7003 (N_7003,N_1082,N_3144);
nor U7004 (N_7004,N_3125,N_4188);
or U7005 (N_7005,N_4286,N_3451);
and U7006 (N_7006,N_798,N_984);
or U7007 (N_7007,N_3096,N_3364);
or U7008 (N_7008,N_3600,N_3592);
xnor U7009 (N_7009,N_4639,N_1722);
or U7010 (N_7010,N_1157,N_786);
or U7011 (N_7011,N_3788,N_2935);
xor U7012 (N_7012,N_642,N_3964);
nand U7013 (N_7013,N_1164,N_4682);
nor U7014 (N_7014,N_1247,N_952);
or U7015 (N_7015,N_808,N_882);
nor U7016 (N_7016,N_1162,N_2207);
or U7017 (N_7017,N_610,N_989);
nor U7018 (N_7018,N_1412,N_2308);
nand U7019 (N_7019,N_4202,N_618);
nand U7020 (N_7020,N_1375,N_218);
or U7021 (N_7021,N_1666,N_2422);
and U7022 (N_7022,N_2510,N_3107);
and U7023 (N_7023,N_4457,N_1556);
or U7024 (N_7024,N_2965,N_4812);
nand U7025 (N_7025,N_871,N_1763);
and U7026 (N_7026,N_4500,N_3253);
or U7027 (N_7027,N_4373,N_4285);
nor U7028 (N_7028,N_291,N_2083);
nor U7029 (N_7029,N_4059,N_3279);
and U7030 (N_7030,N_4973,N_2072);
nor U7031 (N_7031,N_1448,N_719);
or U7032 (N_7032,N_2141,N_380);
nor U7033 (N_7033,N_1889,N_2280);
nor U7034 (N_7034,N_737,N_1688);
or U7035 (N_7035,N_3923,N_3064);
and U7036 (N_7036,N_647,N_206);
or U7037 (N_7037,N_2352,N_2313);
and U7038 (N_7038,N_4330,N_1792);
xor U7039 (N_7039,N_46,N_1531);
nor U7040 (N_7040,N_3343,N_3289);
nand U7041 (N_7041,N_411,N_599);
and U7042 (N_7042,N_4216,N_3251);
nor U7043 (N_7043,N_4214,N_1020);
or U7044 (N_7044,N_16,N_1376);
nand U7045 (N_7045,N_1001,N_4290);
or U7046 (N_7046,N_1705,N_4880);
and U7047 (N_7047,N_646,N_3680);
and U7048 (N_7048,N_4128,N_1520);
nand U7049 (N_7049,N_3843,N_2467);
and U7050 (N_7050,N_2626,N_4831);
nand U7051 (N_7051,N_2477,N_292);
nor U7052 (N_7052,N_4838,N_580);
nor U7053 (N_7053,N_998,N_2530);
and U7054 (N_7054,N_2342,N_677);
nor U7055 (N_7055,N_4801,N_1521);
and U7056 (N_7056,N_1986,N_4069);
or U7057 (N_7057,N_1777,N_1098);
nand U7058 (N_7058,N_3990,N_3085);
or U7059 (N_7059,N_4057,N_3285);
nor U7060 (N_7060,N_2611,N_4814);
or U7061 (N_7061,N_917,N_723);
or U7062 (N_7062,N_4582,N_4861);
nand U7063 (N_7063,N_2560,N_1732);
nand U7064 (N_7064,N_1005,N_523);
nor U7065 (N_7065,N_947,N_1960);
nand U7066 (N_7066,N_165,N_1575);
nand U7067 (N_7067,N_1837,N_2751);
and U7068 (N_7068,N_605,N_1887);
nand U7069 (N_7069,N_428,N_1282);
nor U7070 (N_7070,N_479,N_2335);
and U7071 (N_7071,N_111,N_1655);
nor U7072 (N_7072,N_4790,N_3687);
xor U7073 (N_7073,N_2297,N_284);
and U7074 (N_7074,N_1744,N_2345);
or U7075 (N_7075,N_3790,N_4469);
and U7076 (N_7076,N_4561,N_2937);
nor U7077 (N_7077,N_2650,N_4438);
nand U7078 (N_7078,N_4544,N_163);
nor U7079 (N_7079,N_422,N_499);
or U7080 (N_7080,N_2100,N_4386);
nand U7081 (N_7081,N_4545,N_1058);
or U7082 (N_7082,N_806,N_3307);
or U7083 (N_7083,N_4352,N_4129);
and U7084 (N_7084,N_1910,N_3071);
and U7085 (N_7085,N_3722,N_2483);
nand U7086 (N_7086,N_136,N_1842);
nand U7087 (N_7087,N_2940,N_3588);
nand U7088 (N_7088,N_4763,N_222);
or U7089 (N_7089,N_103,N_838);
or U7090 (N_7090,N_899,N_2753);
or U7091 (N_7091,N_4673,N_2882);
xor U7092 (N_7092,N_1935,N_2719);
or U7093 (N_7093,N_1899,N_2950);
nand U7094 (N_7094,N_3060,N_4737);
nand U7095 (N_7095,N_4983,N_1835);
and U7096 (N_7096,N_3111,N_2372);
nor U7097 (N_7097,N_1316,N_1975);
nor U7098 (N_7098,N_446,N_2889);
or U7099 (N_7099,N_2322,N_2302);
nand U7100 (N_7100,N_1450,N_4194);
nor U7101 (N_7101,N_933,N_3175);
nand U7102 (N_7102,N_1017,N_3325);
and U7103 (N_7103,N_611,N_887);
nor U7104 (N_7104,N_1490,N_2770);
nand U7105 (N_7105,N_3694,N_62);
and U7106 (N_7106,N_2812,N_874);
nand U7107 (N_7107,N_2493,N_1587);
nor U7108 (N_7108,N_4073,N_171);
and U7109 (N_7109,N_1138,N_2127);
and U7110 (N_7110,N_4335,N_3424);
nand U7111 (N_7111,N_2025,N_3538);
nand U7112 (N_7112,N_648,N_3034);
nor U7113 (N_7113,N_1429,N_3465);
nor U7114 (N_7114,N_1035,N_3366);
and U7115 (N_7115,N_3856,N_3733);
nor U7116 (N_7116,N_4366,N_3182);
nor U7117 (N_7117,N_2774,N_1437);
or U7118 (N_7118,N_2131,N_4408);
or U7119 (N_7119,N_3322,N_4446);
and U7120 (N_7120,N_1432,N_1467);
nand U7121 (N_7121,N_1215,N_588);
or U7122 (N_7122,N_2915,N_2998);
or U7123 (N_7123,N_145,N_84);
and U7124 (N_7124,N_2068,N_2243);
nand U7125 (N_7125,N_1622,N_2787);
and U7126 (N_7126,N_3710,N_602);
xor U7127 (N_7127,N_1476,N_4728);
and U7128 (N_7128,N_3779,N_686);
nand U7129 (N_7129,N_525,N_470);
or U7130 (N_7130,N_2572,N_3486);
or U7131 (N_7131,N_3562,N_4402);
nor U7132 (N_7132,N_1726,N_707);
nand U7133 (N_7133,N_3437,N_1670);
nor U7134 (N_7134,N_3618,N_2667);
or U7135 (N_7135,N_3277,N_3129);
and U7136 (N_7136,N_3796,N_1133);
or U7137 (N_7137,N_716,N_2331);
and U7138 (N_7138,N_991,N_3302);
nand U7139 (N_7139,N_875,N_3637);
nand U7140 (N_7140,N_1970,N_711);
or U7141 (N_7141,N_4876,N_3232);
nand U7142 (N_7142,N_3188,N_1773);
and U7143 (N_7143,N_939,N_472);
nor U7144 (N_7144,N_147,N_2255);
and U7145 (N_7145,N_923,N_3854);
or U7146 (N_7146,N_1153,N_876);
xnor U7147 (N_7147,N_1146,N_227);
and U7148 (N_7148,N_2968,N_3635);
xor U7149 (N_7149,N_4939,N_220);
xnor U7150 (N_7150,N_367,N_3055);
or U7151 (N_7151,N_3014,N_2486);
or U7152 (N_7152,N_1145,N_1593);
or U7153 (N_7153,N_3792,N_3857);
and U7154 (N_7154,N_2724,N_3397);
xor U7155 (N_7155,N_377,N_4971);
or U7156 (N_7156,N_330,N_604);
nor U7157 (N_7157,N_569,N_4174);
or U7158 (N_7158,N_4845,N_4870);
and U7159 (N_7159,N_3750,N_1302);
nand U7160 (N_7160,N_2596,N_4863);
and U7161 (N_7161,N_2047,N_2635);
nand U7162 (N_7162,N_902,N_1487);
nand U7163 (N_7163,N_482,N_3692);
and U7164 (N_7164,N_3865,N_938);
xor U7165 (N_7165,N_3532,N_4010);
or U7166 (N_7166,N_1673,N_762);
nand U7167 (N_7167,N_1707,N_4489);
and U7168 (N_7168,N_1988,N_1385);
nand U7169 (N_7169,N_4277,N_1758);
nor U7170 (N_7170,N_936,N_870);
nor U7171 (N_7171,N_4843,N_3335);
or U7172 (N_7172,N_1270,N_3436);
nor U7173 (N_7173,N_818,N_1661);
xnor U7174 (N_7174,N_4849,N_2375);
xnor U7175 (N_7175,N_1581,N_4217);
and U7176 (N_7176,N_4084,N_1488);
or U7177 (N_7177,N_2539,N_4323);
or U7178 (N_7178,N_766,N_3823);
nor U7179 (N_7179,N_3650,N_3148);
xnor U7180 (N_7180,N_4584,N_383);
or U7181 (N_7181,N_3548,N_3993);
nor U7182 (N_7182,N_28,N_1862);
or U7183 (N_7183,N_3062,N_1698);
or U7184 (N_7184,N_1682,N_4354);
nand U7185 (N_7185,N_74,N_4554);
nand U7186 (N_7186,N_278,N_2053);
nor U7187 (N_7187,N_697,N_4229);
nand U7188 (N_7188,N_3852,N_1711);
nand U7189 (N_7189,N_491,N_1059);
and U7190 (N_7190,N_2697,N_1843);
xor U7191 (N_7191,N_3069,N_9);
xor U7192 (N_7192,N_394,N_3272);
xnor U7193 (N_7193,N_1516,N_4667);
nor U7194 (N_7194,N_2513,N_265);
nor U7195 (N_7195,N_2669,N_1181);
xor U7196 (N_7196,N_1214,N_489);
or U7197 (N_7197,N_514,N_3353);
nand U7198 (N_7198,N_2588,N_2104);
xnor U7199 (N_7199,N_4053,N_1884);
xnor U7200 (N_7200,N_255,N_3894);
or U7201 (N_7201,N_4022,N_617);
nor U7202 (N_7202,N_1513,N_4687);
nand U7203 (N_7203,N_4619,N_219);
nand U7204 (N_7204,N_3839,N_1064);
nor U7205 (N_7205,N_3180,N_4864);
and U7206 (N_7206,N_4338,N_1509);
and U7207 (N_7207,N_3341,N_1328);
and U7208 (N_7208,N_4184,N_983);
or U7209 (N_7209,N_3892,N_4750);
or U7210 (N_7210,N_2727,N_4350);
and U7211 (N_7211,N_768,N_3512);
nor U7212 (N_7212,N_1865,N_1373);
and U7213 (N_7213,N_3767,N_3147);
or U7214 (N_7214,N_1872,N_1197);
and U7215 (N_7215,N_1084,N_4935);
nor U7216 (N_7216,N_780,N_268);
nor U7217 (N_7217,N_3485,N_3872);
nand U7218 (N_7218,N_37,N_1645);
nand U7219 (N_7219,N_2465,N_2671);
nor U7220 (N_7220,N_2329,N_1987);
and U7221 (N_7221,N_2173,N_2653);
nand U7222 (N_7222,N_3464,N_3875);
or U7223 (N_7223,N_2678,N_3874);
or U7224 (N_7224,N_2060,N_1319);
nor U7225 (N_7225,N_4796,N_1040);
nor U7226 (N_7226,N_3610,N_4066);
or U7227 (N_7227,N_2201,N_2230);
and U7228 (N_7228,N_1210,N_1990);
or U7229 (N_7229,N_3475,N_3564);
nand U7230 (N_7230,N_4166,N_1544);
nor U7231 (N_7231,N_2702,N_3840);
nand U7232 (N_7232,N_98,N_416);
nand U7233 (N_7233,N_1441,N_3126);
and U7234 (N_7234,N_2815,N_3073);
and U7235 (N_7235,N_2055,N_3707);
or U7236 (N_7236,N_4696,N_2333);
nand U7237 (N_7237,N_2318,N_4921);
nand U7238 (N_7238,N_2242,N_4436);
and U7239 (N_7239,N_1890,N_1459);
nor U7240 (N_7240,N_2427,N_1824);
nand U7241 (N_7241,N_1640,N_3201);
nor U7242 (N_7242,N_3907,N_2964);
nand U7243 (N_7243,N_1469,N_4046);
nand U7244 (N_7244,N_652,N_2451);
nand U7245 (N_7245,N_1921,N_4572);
nand U7246 (N_7246,N_3554,N_4563);
or U7247 (N_7247,N_246,N_314);
nor U7248 (N_7248,N_3186,N_3903);
nor U7249 (N_7249,N_3595,N_254);
nand U7250 (N_7250,N_1131,N_553);
and U7251 (N_7251,N_3620,N_811);
nand U7252 (N_7252,N_1955,N_113);
nor U7253 (N_7253,N_3543,N_2621);
nor U7254 (N_7254,N_4159,N_671);
nand U7255 (N_7255,N_468,N_2102);
nand U7256 (N_7256,N_1036,N_846);
or U7257 (N_7257,N_369,N_2198);
nand U7258 (N_7258,N_2631,N_464);
nor U7259 (N_7259,N_2629,N_2358);
or U7260 (N_7260,N_3800,N_239);
nand U7261 (N_7261,N_2152,N_3145);
and U7262 (N_7262,N_1106,N_3721);
xor U7263 (N_7263,N_980,N_463);
nor U7264 (N_7264,N_117,N_2061);
and U7265 (N_7265,N_2023,N_2087);
or U7266 (N_7266,N_3339,N_4706);
nand U7267 (N_7267,N_2975,N_4192);
nand U7268 (N_7268,N_2488,N_1386);
and U7269 (N_7269,N_1632,N_2077);
or U7270 (N_7270,N_2516,N_730);
xor U7271 (N_7271,N_4774,N_528);
and U7272 (N_7272,N_2442,N_4850);
nand U7273 (N_7273,N_1641,N_371);
or U7274 (N_7274,N_1580,N_3393);
nand U7275 (N_7275,N_2233,N_2446);
and U7276 (N_7276,N_1334,N_195);
or U7277 (N_7277,N_3504,N_2295);
xor U7278 (N_7278,N_4957,N_3591);
or U7279 (N_7279,N_2160,N_3756);
nand U7280 (N_7280,N_3454,N_4615);
nor U7281 (N_7281,N_681,N_2438);
nand U7282 (N_7282,N_107,N_542);
or U7283 (N_7283,N_238,N_2095);
or U7284 (N_7284,N_260,N_3870);
nor U7285 (N_7285,N_1821,N_2969);
or U7286 (N_7286,N_3786,N_1031);
or U7287 (N_7287,N_1030,N_4869);
or U7288 (N_7288,N_2714,N_4789);
nand U7289 (N_7289,N_110,N_1480);
nor U7290 (N_7290,N_689,N_567);
and U7291 (N_7291,N_2690,N_513);
nand U7292 (N_7292,N_412,N_3658);
or U7293 (N_7293,N_3173,N_326);
nand U7294 (N_7294,N_4002,N_4937);
nor U7295 (N_7295,N_3778,N_3065);
nand U7296 (N_7296,N_1034,N_4933);
and U7297 (N_7297,N_4207,N_4187);
nand U7298 (N_7298,N_2299,N_127);
nand U7299 (N_7299,N_2948,N_4759);
or U7300 (N_7300,N_2327,N_3119);
and U7301 (N_7301,N_1407,N_1438);
xnor U7302 (N_7302,N_4116,N_3419);
nand U7303 (N_7303,N_634,N_2562);
nor U7304 (N_7304,N_3590,N_4761);
and U7305 (N_7305,N_4039,N_1111);
or U7306 (N_7306,N_1056,N_3293);
nor U7307 (N_7307,N_3514,N_2555);
nand U7308 (N_7308,N_1811,N_1706);
xor U7309 (N_7309,N_3152,N_3280);
and U7310 (N_7310,N_11,N_387);
or U7311 (N_7311,N_29,N_2416);
or U7312 (N_7312,N_3162,N_583);
and U7313 (N_7313,N_3568,N_483);
and U7314 (N_7314,N_130,N_3099);
nor U7315 (N_7315,N_1981,N_2534);
and U7316 (N_7316,N_3539,N_177);
and U7317 (N_7317,N_2842,N_679);
nor U7318 (N_7318,N_1806,N_2360);
nand U7319 (N_7319,N_2274,N_4477);
or U7320 (N_7320,N_3899,N_2125);
or U7321 (N_7321,N_1370,N_3659);
and U7322 (N_7322,N_3898,N_1269);
nand U7323 (N_7323,N_3191,N_4374);
nand U7324 (N_7324,N_1685,N_4548);
and U7325 (N_7325,N_2759,N_166);
nand U7326 (N_7326,N_3327,N_537);
xnor U7327 (N_7327,N_3832,N_2204);
nand U7328 (N_7328,N_3242,N_3202);
nand U7329 (N_7329,N_3492,N_3529);
xor U7330 (N_7330,N_4568,N_1449);
or U7331 (N_7331,N_1552,N_2802);
xnor U7332 (N_7332,N_3249,N_175);
nor U7333 (N_7333,N_3386,N_4070);
and U7334 (N_7334,N_3256,N_2202);
nand U7335 (N_7335,N_1793,N_1116);
and U7336 (N_7336,N_4447,N_4191);
or U7337 (N_7337,N_4641,N_3032);
nor U7338 (N_7338,N_56,N_3627);
or U7339 (N_7339,N_1021,N_1239);
or U7340 (N_7340,N_1336,N_851);
nor U7341 (N_7341,N_3859,N_2304);
nor U7342 (N_7342,N_4515,N_3830);
or U7343 (N_7343,N_4811,N_4445);
nor U7344 (N_7344,N_4862,N_2319);
and U7345 (N_7345,N_4048,N_4378);
nand U7346 (N_7346,N_1627,N_3314);
or U7347 (N_7347,N_4707,N_1287);
or U7348 (N_7348,N_1231,N_1550);
and U7349 (N_7349,N_4178,N_1322);
nand U7350 (N_7350,N_4067,N_1790);
or U7351 (N_7351,N_3806,N_4230);
and U7352 (N_7352,N_1542,N_459);
nand U7353 (N_7353,N_1576,N_584);
nor U7354 (N_7354,N_669,N_2721);
nor U7355 (N_7355,N_4653,N_3160);
and U7356 (N_7356,N_1209,N_1);
nor U7357 (N_7357,N_3028,N_1142);
or U7358 (N_7358,N_3822,N_630);
and U7359 (N_7359,N_606,N_4395);
or U7360 (N_7360,N_155,N_3460);
nor U7361 (N_7361,N_83,N_3582);
nand U7362 (N_7362,N_4919,N_48);
nand U7363 (N_7363,N_189,N_440);
and U7364 (N_7364,N_256,N_1091);
or U7365 (N_7365,N_2574,N_4043);
nor U7366 (N_7366,N_2142,N_1741);
nand U7367 (N_7367,N_3648,N_2917);
xnor U7368 (N_7368,N_2848,N_4779);
or U7369 (N_7369,N_2817,N_180);
and U7370 (N_7370,N_3585,N_4930);
nand U7371 (N_7371,N_4482,N_1122);
nor U7372 (N_7372,N_3414,N_3416);
nand U7373 (N_7373,N_2094,N_2886);
and U7374 (N_7374,N_317,N_3409);
and U7375 (N_7375,N_4496,N_4282);
and U7376 (N_7376,N_179,N_2878);
and U7377 (N_7377,N_2632,N_3534);
or U7378 (N_7378,N_4324,N_4688);
nor U7379 (N_7379,N_2961,N_2461);
or U7380 (N_7380,N_3320,N_1558);
nor U7381 (N_7381,N_755,N_805);
nand U7382 (N_7382,N_4206,N_1089);
or U7383 (N_7383,N_3642,N_2962);
or U7384 (N_7384,N_2067,N_3624);
nand U7385 (N_7385,N_1756,N_212);
nand U7386 (N_7386,N_1416,N_3930);
xor U7387 (N_7387,N_3601,N_1619);
or U7388 (N_7388,N_3809,N_4014);
or U7389 (N_7389,N_3950,N_3948);
nor U7390 (N_7390,N_4015,N_841);
nor U7391 (N_7391,N_3311,N_3494);
and U7392 (N_7392,N_2820,N_1481);
nor U7393 (N_7393,N_3751,N_1198);
nor U7394 (N_7394,N_934,N_3225);
xor U7395 (N_7395,N_2741,N_2959);
and U7396 (N_7396,N_19,N_3392);
or U7397 (N_7397,N_1176,N_756);
and U7398 (N_7398,N_2374,N_193);
nand U7399 (N_7399,N_3909,N_1569);
nand U7400 (N_7400,N_4104,N_4176);
nand U7401 (N_7401,N_4941,N_4054);
nor U7402 (N_7402,N_4597,N_2226);
nor U7403 (N_7403,N_3617,N_1348);
nor U7404 (N_7404,N_612,N_4308);
nand U7405 (N_7405,N_931,N_2098);
or U7406 (N_7406,N_1626,N_296);
nor U7407 (N_7407,N_2694,N_2247);
nor U7408 (N_7408,N_1944,N_3698);
xor U7409 (N_7409,N_2616,N_2503);
or U7410 (N_7410,N_12,N_2050);
nor U7411 (N_7411,N_4380,N_1586);
or U7412 (N_7412,N_3471,N_3031);
or U7413 (N_7413,N_4418,N_4588);
nor U7414 (N_7414,N_21,N_796);
xor U7415 (N_7415,N_4871,N_415);
nor U7416 (N_7416,N_1808,N_2548);
xnor U7417 (N_7417,N_1338,N_3312);
or U7418 (N_7418,N_3050,N_3143);
and U7419 (N_7419,N_3561,N_2349);
and U7420 (N_7420,N_828,N_2276);
nand U7421 (N_7421,N_807,N_2813);
nor U7422 (N_7422,N_2110,N_1723);
or U7423 (N_7423,N_2757,N_4132);
nor U7424 (N_7424,N_3693,N_356);
nand U7425 (N_7425,N_3350,N_4616);
or U7426 (N_7426,N_4329,N_3265);
or U7427 (N_7427,N_4219,N_3115);
or U7428 (N_7428,N_4903,N_3734);
nor U7429 (N_7429,N_4962,N_2732);
xnor U7430 (N_7430,N_2460,N_4657);
or U7431 (N_7431,N_2119,N_4160);
nand U7432 (N_7432,N_4865,N_263);
xnor U7433 (N_7433,N_4000,N_3137);
nor U7434 (N_7434,N_3326,N_3179);
nor U7435 (N_7435,N_3077,N_2271);
or U7436 (N_7436,N_3553,N_4530);
and U7437 (N_7437,N_2876,N_4671);
nor U7438 (N_7438,N_1366,N_4265);
or U7439 (N_7439,N_4934,N_1780);
xnor U7440 (N_7440,N_71,N_198);
nor U7441 (N_7441,N_778,N_3817);
or U7442 (N_7442,N_1535,N_4236);
nand U7443 (N_7443,N_4231,N_4537);
or U7444 (N_7444,N_1218,N_4087);
nor U7445 (N_7445,N_3927,N_1647);
and U7446 (N_7446,N_4028,N_3759);
nand U7447 (N_7447,N_141,N_4209);
nand U7448 (N_7448,N_4700,N_4918);
and U7449 (N_7449,N_2991,N_1612);
nand U7450 (N_7450,N_4531,N_963);
nor U7451 (N_7451,N_3389,N_826);
and U7452 (N_7452,N_3919,N_2169);
nor U7453 (N_7453,N_3575,N_196);
nand U7454 (N_7454,N_3412,N_2885);
and U7455 (N_7455,N_3519,N_1292);
nand U7456 (N_7456,N_1118,N_977);
nand U7457 (N_7457,N_4910,N_432);
or U7458 (N_7458,N_695,N_4310);
or U7459 (N_7459,N_3951,N_2507);
or U7460 (N_7460,N_4389,N_2767);
xor U7461 (N_7461,N_2919,N_4953);
nor U7462 (N_7462,N_3737,N_2772);
nand U7463 (N_7463,N_2192,N_2059);
and U7464 (N_7464,N_1982,N_1559);
or U7465 (N_7465,N_4499,N_3309);
nand U7466 (N_7466,N_4130,N_3190);
and U7467 (N_7467,N_3544,N_2380);
or U7468 (N_7468,N_4056,N_683);
nand U7469 (N_7469,N_3995,N_3351);
nand U7470 (N_7470,N_1096,N_4586);
or U7471 (N_7471,N_3029,N_4832);
nor U7472 (N_7472,N_3835,N_473);
xnor U7473 (N_7473,N_3718,N_4333);
and U7474 (N_7474,N_897,N_3213);
and U7475 (N_7475,N_4348,N_1526);
nand U7476 (N_7476,N_4895,N_1757);
xor U7477 (N_7477,N_2986,N_4319);
or U7478 (N_7478,N_3672,N_921);
nand U7479 (N_7479,N_2766,N_2237);
nand U7480 (N_7480,N_1532,N_3908);
xnor U7481 (N_7481,N_1381,N_4694);
and U7482 (N_7482,N_760,N_23);
or U7483 (N_7483,N_2235,N_4924);
and U7484 (N_7484,N_1452,N_2831);
or U7485 (N_7485,N_1221,N_437);
nor U7486 (N_7486,N_708,N_4894);
nor U7487 (N_7487,N_1293,N_2613);
or U7488 (N_7488,N_1980,N_2605);
nor U7489 (N_7489,N_2070,N_2883);
xnor U7490 (N_7490,N_658,N_555);
or U7491 (N_7491,N_2290,N_3301);
or U7492 (N_7492,N_3764,N_1783);
nor U7493 (N_7493,N_894,N_2821);
nand U7494 (N_7494,N_2987,N_3212);
or U7495 (N_7495,N_1474,N_821);
and U7496 (N_7496,N_4951,N_4263);
and U7497 (N_7497,N_3895,N_128);
or U7498 (N_7498,N_1107,N_61);
nand U7499 (N_7499,N_1431,N_2561);
or U7500 (N_7500,N_231,N_4567);
and U7501 (N_7501,N_2726,N_3541);
nand U7502 (N_7502,N_4536,N_1858);
nor U7503 (N_7503,N_208,N_429);
and U7504 (N_7504,N_3916,N_1349);
and U7505 (N_7505,N_4454,N_685);
nor U7506 (N_7506,N_2714,N_362);
nor U7507 (N_7507,N_3365,N_1744);
nand U7508 (N_7508,N_4584,N_2805);
nand U7509 (N_7509,N_3290,N_543);
nor U7510 (N_7510,N_2214,N_2030);
nand U7511 (N_7511,N_1236,N_4541);
and U7512 (N_7512,N_718,N_4617);
or U7513 (N_7513,N_2158,N_1911);
or U7514 (N_7514,N_2145,N_2202);
and U7515 (N_7515,N_3577,N_4890);
nor U7516 (N_7516,N_226,N_4377);
and U7517 (N_7517,N_4145,N_2201);
and U7518 (N_7518,N_988,N_2207);
or U7519 (N_7519,N_4800,N_1954);
nor U7520 (N_7520,N_1463,N_3637);
or U7521 (N_7521,N_354,N_1727);
or U7522 (N_7522,N_3400,N_4729);
nor U7523 (N_7523,N_2708,N_2292);
nand U7524 (N_7524,N_495,N_924);
and U7525 (N_7525,N_1624,N_3894);
nand U7526 (N_7526,N_365,N_4211);
nand U7527 (N_7527,N_3812,N_3777);
nand U7528 (N_7528,N_1446,N_3483);
and U7529 (N_7529,N_3795,N_1449);
nand U7530 (N_7530,N_2338,N_628);
nor U7531 (N_7531,N_4866,N_3823);
nor U7532 (N_7532,N_581,N_2195);
nor U7533 (N_7533,N_2061,N_1234);
and U7534 (N_7534,N_2226,N_404);
nor U7535 (N_7535,N_4728,N_4576);
and U7536 (N_7536,N_3777,N_1937);
and U7537 (N_7537,N_1463,N_4106);
or U7538 (N_7538,N_509,N_4192);
and U7539 (N_7539,N_340,N_738);
or U7540 (N_7540,N_1713,N_329);
nand U7541 (N_7541,N_4484,N_1948);
and U7542 (N_7542,N_3357,N_3986);
or U7543 (N_7543,N_997,N_3131);
xnor U7544 (N_7544,N_1126,N_2657);
or U7545 (N_7545,N_669,N_2219);
nor U7546 (N_7546,N_1001,N_242);
xnor U7547 (N_7547,N_3830,N_2402);
and U7548 (N_7548,N_3283,N_2124);
or U7549 (N_7549,N_2991,N_3596);
nand U7550 (N_7550,N_304,N_4575);
nand U7551 (N_7551,N_74,N_4593);
nor U7552 (N_7552,N_142,N_4316);
nand U7553 (N_7553,N_950,N_4706);
or U7554 (N_7554,N_3705,N_3028);
nand U7555 (N_7555,N_3696,N_4236);
or U7556 (N_7556,N_4753,N_2848);
and U7557 (N_7557,N_2057,N_4922);
nor U7558 (N_7558,N_1034,N_3109);
nor U7559 (N_7559,N_2599,N_4872);
nand U7560 (N_7560,N_3932,N_4135);
and U7561 (N_7561,N_845,N_469);
nand U7562 (N_7562,N_1173,N_1073);
and U7563 (N_7563,N_4034,N_4338);
or U7564 (N_7564,N_497,N_3621);
nor U7565 (N_7565,N_3428,N_2358);
nor U7566 (N_7566,N_4601,N_2451);
nand U7567 (N_7567,N_791,N_4422);
and U7568 (N_7568,N_741,N_439);
nor U7569 (N_7569,N_4200,N_2186);
and U7570 (N_7570,N_2599,N_2466);
or U7571 (N_7571,N_2667,N_2287);
nand U7572 (N_7572,N_158,N_3073);
or U7573 (N_7573,N_19,N_4181);
and U7574 (N_7574,N_321,N_509);
nand U7575 (N_7575,N_3579,N_1554);
and U7576 (N_7576,N_3353,N_375);
and U7577 (N_7577,N_590,N_4805);
nor U7578 (N_7578,N_2925,N_4979);
nor U7579 (N_7579,N_4594,N_204);
nand U7580 (N_7580,N_3652,N_1754);
or U7581 (N_7581,N_3662,N_1982);
or U7582 (N_7582,N_2126,N_2228);
or U7583 (N_7583,N_4273,N_3610);
nand U7584 (N_7584,N_1561,N_2562);
xnor U7585 (N_7585,N_601,N_3582);
xnor U7586 (N_7586,N_3561,N_3389);
nor U7587 (N_7587,N_1323,N_4841);
nand U7588 (N_7588,N_1337,N_973);
nand U7589 (N_7589,N_2585,N_532);
nor U7590 (N_7590,N_4214,N_1872);
nand U7591 (N_7591,N_467,N_682);
nor U7592 (N_7592,N_4171,N_3434);
and U7593 (N_7593,N_739,N_2695);
or U7594 (N_7594,N_594,N_3525);
or U7595 (N_7595,N_3184,N_1090);
nor U7596 (N_7596,N_4058,N_740);
nand U7597 (N_7597,N_2298,N_465);
and U7598 (N_7598,N_827,N_3435);
xor U7599 (N_7599,N_2899,N_3503);
nand U7600 (N_7600,N_2371,N_3904);
or U7601 (N_7601,N_4528,N_3508);
nand U7602 (N_7602,N_471,N_4887);
nand U7603 (N_7603,N_747,N_3948);
nand U7604 (N_7604,N_1093,N_3619);
or U7605 (N_7605,N_3185,N_1425);
nand U7606 (N_7606,N_2457,N_4966);
or U7607 (N_7607,N_187,N_3782);
or U7608 (N_7608,N_724,N_646);
nand U7609 (N_7609,N_4542,N_354);
and U7610 (N_7610,N_977,N_3471);
xnor U7611 (N_7611,N_3938,N_2112);
and U7612 (N_7612,N_2614,N_312);
or U7613 (N_7613,N_3625,N_3930);
or U7614 (N_7614,N_696,N_1344);
xor U7615 (N_7615,N_4022,N_3162);
or U7616 (N_7616,N_112,N_319);
and U7617 (N_7617,N_1392,N_3097);
and U7618 (N_7618,N_2351,N_352);
or U7619 (N_7619,N_1203,N_4907);
or U7620 (N_7620,N_2613,N_2622);
or U7621 (N_7621,N_2343,N_3487);
nand U7622 (N_7622,N_1962,N_2317);
or U7623 (N_7623,N_1096,N_3051);
and U7624 (N_7624,N_51,N_3805);
nor U7625 (N_7625,N_2245,N_496);
nand U7626 (N_7626,N_2048,N_4013);
and U7627 (N_7627,N_74,N_2031);
and U7628 (N_7628,N_1310,N_1602);
or U7629 (N_7629,N_471,N_3747);
nor U7630 (N_7630,N_1862,N_4353);
nand U7631 (N_7631,N_4093,N_2183);
nand U7632 (N_7632,N_2612,N_4747);
or U7633 (N_7633,N_421,N_1554);
and U7634 (N_7634,N_2178,N_3658);
nand U7635 (N_7635,N_1814,N_4147);
and U7636 (N_7636,N_4157,N_2394);
or U7637 (N_7637,N_3399,N_4465);
and U7638 (N_7638,N_4566,N_2486);
nor U7639 (N_7639,N_3207,N_1296);
nor U7640 (N_7640,N_611,N_1333);
xor U7641 (N_7641,N_4464,N_3757);
or U7642 (N_7642,N_4296,N_3779);
or U7643 (N_7643,N_3632,N_2056);
xnor U7644 (N_7644,N_863,N_1789);
and U7645 (N_7645,N_1016,N_109);
nand U7646 (N_7646,N_3261,N_3268);
or U7647 (N_7647,N_1605,N_3345);
or U7648 (N_7648,N_2662,N_3063);
nand U7649 (N_7649,N_4859,N_1627);
nor U7650 (N_7650,N_1659,N_1303);
and U7651 (N_7651,N_4372,N_4085);
and U7652 (N_7652,N_2570,N_4638);
and U7653 (N_7653,N_3980,N_2459);
or U7654 (N_7654,N_2006,N_3828);
nor U7655 (N_7655,N_1246,N_752);
nand U7656 (N_7656,N_4921,N_4568);
nand U7657 (N_7657,N_606,N_3067);
nand U7658 (N_7658,N_3131,N_403);
and U7659 (N_7659,N_2501,N_1996);
nand U7660 (N_7660,N_2372,N_393);
or U7661 (N_7661,N_4393,N_686);
or U7662 (N_7662,N_3657,N_1005);
nand U7663 (N_7663,N_1608,N_2394);
nor U7664 (N_7664,N_1701,N_3421);
nand U7665 (N_7665,N_3978,N_982);
and U7666 (N_7666,N_2872,N_2984);
or U7667 (N_7667,N_4548,N_3342);
xnor U7668 (N_7668,N_2870,N_504);
or U7669 (N_7669,N_1019,N_4763);
and U7670 (N_7670,N_3543,N_4003);
nand U7671 (N_7671,N_3018,N_4634);
nor U7672 (N_7672,N_655,N_101);
or U7673 (N_7673,N_2066,N_580);
or U7674 (N_7674,N_1081,N_76);
nand U7675 (N_7675,N_1162,N_1954);
xor U7676 (N_7676,N_1424,N_1433);
or U7677 (N_7677,N_4698,N_4052);
xor U7678 (N_7678,N_1952,N_4455);
nand U7679 (N_7679,N_609,N_605);
nand U7680 (N_7680,N_4087,N_1053);
and U7681 (N_7681,N_1594,N_1346);
nand U7682 (N_7682,N_3084,N_3706);
nand U7683 (N_7683,N_4952,N_1453);
or U7684 (N_7684,N_45,N_2960);
or U7685 (N_7685,N_3527,N_2421);
or U7686 (N_7686,N_2179,N_4326);
and U7687 (N_7687,N_160,N_3398);
or U7688 (N_7688,N_2982,N_406);
xor U7689 (N_7689,N_4959,N_3035);
xor U7690 (N_7690,N_4874,N_4032);
or U7691 (N_7691,N_3682,N_1697);
and U7692 (N_7692,N_3135,N_2173);
nand U7693 (N_7693,N_4516,N_3141);
nor U7694 (N_7694,N_4666,N_4892);
or U7695 (N_7695,N_3623,N_2327);
and U7696 (N_7696,N_1931,N_1947);
or U7697 (N_7697,N_1490,N_4570);
and U7698 (N_7698,N_4126,N_3625);
and U7699 (N_7699,N_911,N_1905);
nand U7700 (N_7700,N_2336,N_2171);
and U7701 (N_7701,N_3261,N_1821);
or U7702 (N_7702,N_3337,N_4355);
and U7703 (N_7703,N_3224,N_313);
nand U7704 (N_7704,N_3321,N_4090);
or U7705 (N_7705,N_571,N_2823);
or U7706 (N_7706,N_3483,N_1821);
nor U7707 (N_7707,N_2902,N_4183);
nor U7708 (N_7708,N_2380,N_3454);
and U7709 (N_7709,N_3186,N_2353);
or U7710 (N_7710,N_4277,N_2776);
and U7711 (N_7711,N_4384,N_362);
or U7712 (N_7712,N_4838,N_290);
nand U7713 (N_7713,N_3354,N_4394);
nand U7714 (N_7714,N_4826,N_4766);
nand U7715 (N_7715,N_495,N_2921);
and U7716 (N_7716,N_3381,N_2320);
and U7717 (N_7717,N_2609,N_3912);
or U7718 (N_7718,N_3366,N_2941);
or U7719 (N_7719,N_705,N_4949);
xnor U7720 (N_7720,N_2413,N_2812);
xor U7721 (N_7721,N_2069,N_607);
or U7722 (N_7722,N_2082,N_235);
nor U7723 (N_7723,N_4364,N_2694);
nor U7724 (N_7724,N_752,N_2820);
nand U7725 (N_7725,N_2432,N_1638);
nand U7726 (N_7726,N_3084,N_3328);
or U7727 (N_7727,N_2051,N_1285);
and U7728 (N_7728,N_3260,N_3374);
nand U7729 (N_7729,N_4669,N_2882);
or U7730 (N_7730,N_3324,N_1123);
nor U7731 (N_7731,N_903,N_4415);
nand U7732 (N_7732,N_1926,N_3923);
or U7733 (N_7733,N_3091,N_3379);
or U7734 (N_7734,N_105,N_2958);
or U7735 (N_7735,N_2162,N_2071);
nor U7736 (N_7736,N_3000,N_2922);
or U7737 (N_7737,N_2016,N_1526);
nand U7738 (N_7738,N_2030,N_2015);
nand U7739 (N_7739,N_4848,N_4660);
xnor U7740 (N_7740,N_2222,N_1729);
nand U7741 (N_7741,N_2499,N_4053);
and U7742 (N_7742,N_4656,N_1833);
nor U7743 (N_7743,N_1094,N_842);
nand U7744 (N_7744,N_3805,N_388);
nor U7745 (N_7745,N_1404,N_932);
nand U7746 (N_7746,N_2285,N_340);
or U7747 (N_7747,N_1734,N_2373);
nand U7748 (N_7748,N_31,N_343);
and U7749 (N_7749,N_3885,N_3922);
nor U7750 (N_7750,N_2429,N_4641);
or U7751 (N_7751,N_1110,N_3757);
nand U7752 (N_7752,N_4352,N_4181);
nor U7753 (N_7753,N_4261,N_4724);
and U7754 (N_7754,N_2937,N_2842);
nor U7755 (N_7755,N_1586,N_4401);
nand U7756 (N_7756,N_2593,N_4551);
nor U7757 (N_7757,N_3567,N_4444);
or U7758 (N_7758,N_4353,N_2122);
nor U7759 (N_7759,N_2184,N_2386);
or U7760 (N_7760,N_4932,N_2418);
nor U7761 (N_7761,N_983,N_2355);
nand U7762 (N_7762,N_2693,N_1099);
nand U7763 (N_7763,N_538,N_4568);
xnor U7764 (N_7764,N_560,N_3304);
nor U7765 (N_7765,N_2262,N_2597);
and U7766 (N_7766,N_3618,N_3548);
xor U7767 (N_7767,N_1142,N_897);
nand U7768 (N_7768,N_2395,N_1720);
xnor U7769 (N_7769,N_3159,N_4120);
xor U7770 (N_7770,N_2988,N_4007);
nand U7771 (N_7771,N_4989,N_4149);
nand U7772 (N_7772,N_3435,N_4134);
xor U7773 (N_7773,N_3381,N_64);
or U7774 (N_7774,N_3020,N_1259);
or U7775 (N_7775,N_4840,N_2899);
or U7776 (N_7776,N_4510,N_4231);
and U7777 (N_7777,N_1450,N_3334);
and U7778 (N_7778,N_1627,N_4392);
or U7779 (N_7779,N_1844,N_1713);
nor U7780 (N_7780,N_1536,N_4120);
and U7781 (N_7781,N_736,N_4492);
and U7782 (N_7782,N_7,N_2058);
xor U7783 (N_7783,N_2424,N_3214);
nand U7784 (N_7784,N_3698,N_1860);
xor U7785 (N_7785,N_4607,N_1187);
nand U7786 (N_7786,N_482,N_3172);
nand U7787 (N_7787,N_4600,N_3563);
or U7788 (N_7788,N_4061,N_3982);
nand U7789 (N_7789,N_1591,N_48);
or U7790 (N_7790,N_2241,N_904);
or U7791 (N_7791,N_871,N_3391);
or U7792 (N_7792,N_4100,N_2776);
or U7793 (N_7793,N_13,N_3188);
and U7794 (N_7794,N_2366,N_835);
nand U7795 (N_7795,N_810,N_3548);
and U7796 (N_7796,N_4882,N_2327);
and U7797 (N_7797,N_2836,N_2960);
nor U7798 (N_7798,N_3377,N_3128);
xor U7799 (N_7799,N_4155,N_4456);
and U7800 (N_7800,N_3963,N_950);
or U7801 (N_7801,N_2562,N_1048);
or U7802 (N_7802,N_91,N_2229);
nor U7803 (N_7803,N_147,N_3233);
nor U7804 (N_7804,N_4971,N_3286);
or U7805 (N_7805,N_4540,N_3715);
and U7806 (N_7806,N_1869,N_3827);
nor U7807 (N_7807,N_3780,N_3699);
nand U7808 (N_7808,N_594,N_3741);
and U7809 (N_7809,N_4980,N_3121);
and U7810 (N_7810,N_3330,N_3844);
xor U7811 (N_7811,N_297,N_337);
or U7812 (N_7812,N_3959,N_2600);
and U7813 (N_7813,N_2036,N_4123);
xnor U7814 (N_7814,N_3665,N_4465);
nand U7815 (N_7815,N_2455,N_542);
or U7816 (N_7816,N_814,N_4145);
nor U7817 (N_7817,N_3937,N_1765);
nor U7818 (N_7818,N_3942,N_3484);
or U7819 (N_7819,N_4408,N_452);
and U7820 (N_7820,N_1236,N_721);
xor U7821 (N_7821,N_1084,N_249);
or U7822 (N_7822,N_924,N_1581);
nor U7823 (N_7823,N_2934,N_1602);
or U7824 (N_7824,N_2049,N_4021);
or U7825 (N_7825,N_4759,N_3078);
and U7826 (N_7826,N_3852,N_1454);
and U7827 (N_7827,N_905,N_1749);
or U7828 (N_7828,N_3291,N_4126);
and U7829 (N_7829,N_2741,N_4387);
or U7830 (N_7830,N_3202,N_4050);
xnor U7831 (N_7831,N_3497,N_2267);
xnor U7832 (N_7832,N_4628,N_4248);
nor U7833 (N_7833,N_43,N_3712);
nand U7834 (N_7834,N_3153,N_621);
nor U7835 (N_7835,N_1423,N_3537);
nor U7836 (N_7836,N_4888,N_1292);
xnor U7837 (N_7837,N_4412,N_652);
nor U7838 (N_7838,N_1699,N_4456);
or U7839 (N_7839,N_3945,N_2392);
xnor U7840 (N_7840,N_1886,N_3827);
nand U7841 (N_7841,N_1727,N_4465);
or U7842 (N_7842,N_146,N_1731);
or U7843 (N_7843,N_1578,N_1983);
and U7844 (N_7844,N_2777,N_1619);
or U7845 (N_7845,N_2226,N_538);
or U7846 (N_7846,N_4588,N_1975);
xnor U7847 (N_7847,N_2580,N_1124);
nor U7848 (N_7848,N_1609,N_2568);
or U7849 (N_7849,N_2931,N_960);
nor U7850 (N_7850,N_2035,N_3956);
and U7851 (N_7851,N_3523,N_3401);
xnor U7852 (N_7852,N_4565,N_1079);
or U7853 (N_7853,N_358,N_65);
or U7854 (N_7854,N_2708,N_1136);
nor U7855 (N_7855,N_1875,N_718);
and U7856 (N_7856,N_848,N_2939);
nand U7857 (N_7857,N_2101,N_1285);
and U7858 (N_7858,N_2149,N_4945);
or U7859 (N_7859,N_2599,N_4262);
nor U7860 (N_7860,N_631,N_2812);
and U7861 (N_7861,N_2206,N_4437);
and U7862 (N_7862,N_3147,N_2844);
nand U7863 (N_7863,N_4613,N_2865);
nor U7864 (N_7864,N_4726,N_242);
nand U7865 (N_7865,N_119,N_1453);
nor U7866 (N_7866,N_2945,N_1281);
nand U7867 (N_7867,N_4052,N_4622);
or U7868 (N_7868,N_4509,N_1919);
and U7869 (N_7869,N_3395,N_1212);
nor U7870 (N_7870,N_4203,N_4876);
xnor U7871 (N_7871,N_1357,N_515);
or U7872 (N_7872,N_3485,N_4913);
nor U7873 (N_7873,N_2925,N_3779);
xnor U7874 (N_7874,N_852,N_1959);
and U7875 (N_7875,N_617,N_4568);
xor U7876 (N_7876,N_434,N_3419);
or U7877 (N_7877,N_4188,N_4900);
xor U7878 (N_7878,N_4506,N_1345);
or U7879 (N_7879,N_2098,N_4570);
nor U7880 (N_7880,N_1604,N_917);
nand U7881 (N_7881,N_1029,N_840);
and U7882 (N_7882,N_3466,N_252);
nand U7883 (N_7883,N_1019,N_2369);
nor U7884 (N_7884,N_1338,N_3104);
nor U7885 (N_7885,N_739,N_3000);
xnor U7886 (N_7886,N_2222,N_148);
and U7887 (N_7887,N_2681,N_2866);
xor U7888 (N_7888,N_1336,N_1602);
or U7889 (N_7889,N_4276,N_562);
nor U7890 (N_7890,N_2123,N_851);
nand U7891 (N_7891,N_3707,N_1948);
nor U7892 (N_7892,N_1069,N_1387);
xnor U7893 (N_7893,N_446,N_1074);
nand U7894 (N_7894,N_1589,N_4589);
nor U7895 (N_7895,N_1384,N_885);
nand U7896 (N_7896,N_4089,N_185);
nor U7897 (N_7897,N_2630,N_3641);
nand U7898 (N_7898,N_1619,N_2541);
xnor U7899 (N_7899,N_332,N_4046);
nor U7900 (N_7900,N_3873,N_1958);
xor U7901 (N_7901,N_4128,N_1117);
nand U7902 (N_7902,N_2590,N_2438);
nand U7903 (N_7903,N_2674,N_2710);
or U7904 (N_7904,N_3456,N_4215);
xor U7905 (N_7905,N_3610,N_4034);
nor U7906 (N_7906,N_1217,N_2561);
xnor U7907 (N_7907,N_3511,N_3633);
and U7908 (N_7908,N_3319,N_2758);
or U7909 (N_7909,N_4280,N_3388);
and U7910 (N_7910,N_172,N_2661);
or U7911 (N_7911,N_3355,N_1503);
nor U7912 (N_7912,N_4315,N_1859);
and U7913 (N_7913,N_3867,N_1751);
or U7914 (N_7914,N_4740,N_4817);
and U7915 (N_7915,N_135,N_4128);
or U7916 (N_7916,N_4181,N_4120);
or U7917 (N_7917,N_355,N_2430);
nand U7918 (N_7918,N_1411,N_317);
or U7919 (N_7919,N_868,N_1490);
nand U7920 (N_7920,N_3872,N_364);
and U7921 (N_7921,N_2506,N_921);
nor U7922 (N_7922,N_942,N_3395);
and U7923 (N_7923,N_1139,N_3013);
and U7924 (N_7924,N_1334,N_608);
nor U7925 (N_7925,N_4601,N_3547);
nand U7926 (N_7926,N_982,N_4811);
or U7927 (N_7927,N_2847,N_4464);
nor U7928 (N_7928,N_4126,N_4688);
nand U7929 (N_7929,N_2703,N_857);
or U7930 (N_7930,N_2659,N_3251);
and U7931 (N_7931,N_1731,N_1682);
or U7932 (N_7932,N_2457,N_592);
and U7933 (N_7933,N_658,N_1125);
or U7934 (N_7934,N_1221,N_3458);
and U7935 (N_7935,N_966,N_1508);
and U7936 (N_7936,N_2543,N_1794);
nor U7937 (N_7937,N_1517,N_3309);
or U7938 (N_7938,N_4558,N_3543);
and U7939 (N_7939,N_4554,N_2336);
nand U7940 (N_7940,N_3664,N_4266);
nand U7941 (N_7941,N_3126,N_215);
nor U7942 (N_7942,N_851,N_4972);
and U7943 (N_7943,N_442,N_4410);
and U7944 (N_7944,N_375,N_3568);
xor U7945 (N_7945,N_1566,N_4023);
nand U7946 (N_7946,N_3967,N_1078);
or U7947 (N_7947,N_4347,N_4164);
and U7948 (N_7948,N_3108,N_4291);
nand U7949 (N_7949,N_3682,N_3850);
nand U7950 (N_7950,N_4568,N_1701);
or U7951 (N_7951,N_3899,N_4938);
or U7952 (N_7952,N_2533,N_793);
and U7953 (N_7953,N_2827,N_1142);
nand U7954 (N_7954,N_2171,N_4497);
and U7955 (N_7955,N_4442,N_1180);
nand U7956 (N_7956,N_2081,N_381);
nor U7957 (N_7957,N_1769,N_4);
or U7958 (N_7958,N_4081,N_292);
or U7959 (N_7959,N_359,N_4870);
nand U7960 (N_7960,N_4512,N_4430);
and U7961 (N_7961,N_3949,N_4152);
xnor U7962 (N_7962,N_1634,N_4556);
nor U7963 (N_7963,N_4018,N_2482);
nand U7964 (N_7964,N_2614,N_2391);
or U7965 (N_7965,N_4633,N_2308);
and U7966 (N_7966,N_1692,N_3697);
and U7967 (N_7967,N_590,N_3039);
and U7968 (N_7968,N_4697,N_1590);
xnor U7969 (N_7969,N_1880,N_482);
and U7970 (N_7970,N_984,N_3898);
nand U7971 (N_7971,N_3689,N_750);
nor U7972 (N_7972,N_3794,N_2975);
nand U7973 (N_7973,N_3579,N_1789);
nor U7974 (N_7974,N_1082,N_3868);
nand U7975 (N_7975,N_4318,N_317);
and U7976 (N_7976,N_291,N_3760);
and U7977 (N_7977,N_1136,N_4376);
nor U7978 (N_7978,N_3856,N_4519);
nand U7979 (N_7979,N_1023,N_2994);
and U7980 (N_7980,N_2106,N_1010);
nand U7981 (N_7981,N_1995,N_771);
nor U7982 (N_7982,N_1648,N_4791);
nor U7983 (N_7983,N_337,N_1375);
and U7984 (N_7984,N_267,N_1478);
and U7985 (N_7985,N_1718,N_3067);
nand U7986 (N_7986,N_4466,N_943);
nor U7987 (N_7987,N_2100,N_1933);
nor U7988 (N_7988,N_2983,N_3556);
xnor U7989 (N_7989,N_3461,N_2929);
xnor U7990 (N_7990,N_2577,N_607);
or U7991 (N_7991,N_3844,N_4752);
and U7992 (N_7992,N_2080,N_1281);
nor U7993 (N_7993,N_4971,N_981);
nand U7994 (N_7994,N_2254,N_3420);
nor U7995 (N_7995,N_1184,N_3650);
nand U7996 (N_7996,N_1628,N_2347);
nand U7997 (N_7997,N_578,N_166);
nor U7998 (N_7998,N_2017,N_2931);
and U7999 (N_7999,N_4101,N_868);
xor U8000 (N_8000,N_409,N_3469);
and U8001 (N_8001,N_2524,N_4731);
nand U8002 (N_8002,N_3173,N_4818);
and U8003 (N_8003,N_4107,N_1608);
or U8004 (N_8004,N_1834,N_2778);
nor U8005 (N_8005,N_4661,N_3709);
nand U8006 (N_8006,N_2292,N_4844);
nor U8007 (N_8007,N_4457,N_4595);
and U8008 (N_8008,N_2581,N_102);
or U8009 (N_8009,N_527,N_4971);
nand U8010 (N_8010,N_1939,N_4959);
or U8011 (N_8011,N_2928,N_4460);
and U8012 (N_8012,N_4289,N_4019);
nor U8013 (N_8013,N_4010,N_270);
or U8014 (N_8014,N_3739,N_4786);
and U8015 (N_8015,N_4187,N_4094);
and U8016 (N_8016,N_3341,N_1946);
nand U8017 (N_8017,N_3340,N_2212);
and U8018 (N_8018,N_1849,N_555);
and U8019 (N_8019,N_4178,N_4651);
or U8020 (N_8020,N_2810,N_995);
nand U8021 (N_8021,N_1572,N_730);
or U8022 (N_8022,N_3960,N_4376);
nand U8023 (N_8023,N_3718,N_2549);
nand U8024 (N_8024,N_786,N_1388);
nand U8025 (N_8025,N_1768,N_4310);
and U8026 (N_8026,N_1419,N_3100);
or U8027 (N_8027,N_3774,N_364);
nand U8028 (N_8028,N_3113,N_2835);
nand U8029 (N_8029,N_2215,N_4365);
nand U8030 (N_8030,N_4056,N_3944);
nand U8031 (N_8031,N_2451,N_1151);
or U8032 (N_8032,N_4310,N_854);
nand U8033 (N_8033,N_4746,N_2454);
and U8034 (N_8034,N_3359,N_1345);
nand U8035 (N_8035,N_3888,N_399);
and U8036 (N_8036,N_1779,N_1927);
nor U8037 (N_8037,N_4583,N_1482);
xor U8038 (N_8038,N_4209,N_2924);
nand U8039 (N_8039,N_3083,N_4307);
nor U8040 (N_8040,N_2924,N_4605);
nand U8041 (N_8041,N_3228,N_2182);
nand U8042 (N_8042,N_4646,N_3002);
or U8043 (N_8043,N_4049,N_3010);
nor U8044 (N_8044,N_3797,N_1994);
or U8045 (N_8045,N_4513,N_2748);
and U8046 (N_8046,N_1117,N_3492);
nor U8047 (N_8047,N_1598,N_2666);
nor U8048 (N_8048,N_1663,N_470);
nor U8049 (N_8049,N_275,N_1626);
nor U8050 (N_8050,N_1676,N_1844);
nand U8051 (N_8051,N_2165,N_2696);
and U8052 (N_8052,N_287,N_1642);
and U8053 (N_8053,N_2522,N_3890);
and U8054 (N_8054,N_1711,N_3693);
and U8055 (N_8055,N_3687,N_682);
or U8056 (N_8056,N_3634,N_1648);
xnor U8057 (N_8057,N_3066,N_2295);
nand U8058 (N_8058,N_1499,N_1207);
nor U8059 (N_8059,N_2264,N_911);
xor U8060 (N_8060,N_2934,N_1680);
nor U8061 (N_8061,N_3313,N_1352);
nand U8062 (N_8062,N_3909,N_4608);
and U8063 (N_8063,N_644,N_4462);
and U8064 (N_8064,N_1933,N_4049);
nand U8065 (N_8065,N_2011,N_407);
or U8066 (N_8066,N_4733,N_1580);
nor U8067 (N_8067,N_1658,N_4583);
and U8068 (N_8068,N_644,N_3736);
and U8069 (N_8069,N_206,N_2053);
nor U8070 (N_8070,N_2848,N_2965);
nand U8071 (N_8071,N_2244,N_1072);
nor U8072 (N_8072,N_1049,N_2319);
nor U8073 (N_8073,N_644,N_4879);
nand U8074 (N_8074,N_2615,N_793);
xnor U8075 (N_8075,N_3000,N_4433);
nor U8076 (N_8076,N_228,N_4983);
or U8077 (N_8077,N_3516,N_1175);
nor U8078 (N_8078,N_3177,N_1986);
and U8079 (N_8079,N_4761,N_2838);
or U8080 (N_8080,N_265,N_1550);
xnor U8081 (N_8081,N_3230,N_3245);
nor U8082 (N_8082,N_1461,N_3030);
or U8083 (N_8083,N_3353,N_1337);
and U8084 (N_8084,N_2522,N_307);
or U8085 (N_8085,N_1803,N_4953);
and U8086 (N_8086,N_3422,N_4816);
nor U8087 (N_8087,N_3663,N_485);
and U8088 (N_8088,N_4677,N_4138);
or U8089 (N_8089,N_271,N_3207);
or U8090 (N_8090,N_993,N_4084);
and U8091 (N_8091,N_3062,N_2574);
nand U8092 (N_8092,N_2884,N_4361);
nor U8093 (N_8093,N_4107,N_4490);
nor U8094 (N_8094,N_3760,N_1184);
and U8095 (N_8095,N_3048,N_3490);
and U8096 (N_8096,N_1867,N_3013);
or U8097 (N_8097,N_707,N_2644);
or U8098 (N_8098,N_1351,N_4586);
nor U8099 (N_8099,N_4718,N_169);
or U8100 (N_8100,N_2437,N_3251);
and U8101 (N_8101,N_4808,N_2325);
and U8102 (N_8102,N_320,N_3240);
or U8103 (N_8103,N_1645,N_31);
nand U8104 (N_8104,N_1446,N_3107);
nand U8105 (N_8105,N_4096,N_905);
nor U8106 (N_8106,N_262,N_1070);
nor U8107 (N_8107,N_462,N_3702);
or U8108 (N_8108,N_2965,N_16);
or U8109 (N_8109,N_4210,N_120);
nand U8110 (N_8110,N_1099,N_276);
xnor U8111 (N_8111,N_160,N_1636);
xor U8112 (N_8112,N_4887,N_2244);
or U8113 (N_8113,N_4234,N_1664);
nor U8114 (N_8114,N_2128,N_1084);
or U8115 (N_8115,N_4231,N_3892);
nor U8116 (N_8116,N_4960,N_3170);
xor U8117 (N_8117,N_1851,N_4036);
xnor U8118 (N_8118,N_1494,N_3762);
or U8119 (N_8119,N_1139,N_4491);
xnor U8120 (N_8120,N_3298,N_1796);
and U8121 (N_8121,N_2695,N_4403);
or U8122 (N_8122,N_2030,N_4769);
nor U8123 (N_8123,N_1521,N_2097);
nor U8124 (N_8124,N_2333,N_143);
nand U8125 (N_8125,N_4740,N_4821);
and U8126 (N_8126,N_2868,N_3126);
nor U8127 (N_8127,N_4317,N_2547);
and U8128 (N_8128,N_2626,N_1565);
or U8129 (N_8129,N_1193,N_322);
nand U8130 (N_8130,N_1397,N_2670);
xor U8131 (N_8131,N_743,N_3029);
and U8132 (N_8132,N_3149,N_1903);
nor U8133 (N_8133,N_1174,N_423);
nor U8134 (N_8134,N_168,N_3513);
nand U8135 (N_8135,N_1442,N_422);
or U8136 (N_8136,N_616,N_4523);
or U8137 (N_8137,N_3695,N_3308);
nor U8138 (N_8138,N_2648,N_917);
and U8139 (N_8139,N_646,N_4815);
xor U8140 (N_8140,N_4296,N_4709);
or U8141 (N_8141,N_205,N_1943);
nand U8142 (N_8142,N_3467,N_3342);
xor U8143 (N_8143,N_3350,N_4480);
or U8144 (N_8144,N_4126,N_4893);
or U8145 (N_8145,N_3341,N_2170);
and U8146 (N_8146,N_2602,N_4479);
or U8147 (N_8147,N_501,N_1836);
nand U8148 (N_8148,N_744,N_3322);
nor U8149 (N_8149,N_2783,N_2579);
or U8150 (N_8150,N_1291,N_2194);
nand U8151 (N_8151,N_246,N_4389);
nor U8152 (N_8152,N_4851,N_2276);
nand U8153 (N_8153,N_3746,N_1385);
nor U8154 (N_8154,N_389,N_4639);
xor U8155 (N_8155,N_211,N_1293);
and U8156 (N_8156,N_3220,N_1123);
nand U8157 (N_8157,N_1456,N_1857);
and U8158 (N_8158,N_1363,N_1908);
nor U8159 (N_8159,N_2683,N_2087);
xnor U8160 (N_8160,N_393,N_1329);
and U8161 (N_8161,N_1348,N_2517);
and U8162 (N_8162,N_2007,N_2182);
nand U8163 (N_8163,N_2030,N_1003);
or U8164 (N_8164,N_2864,N_536);
nand U8165 (N_8165,N_2510,N_4049);
or U8166 (N_8166,N_3737,N_620);
and U8167 (N_8167,N_4802,N_3139);
or U8168 (N_8168,N_3068,N_663);
or U8169 (N_8169,N_4040,N_2443);
nand U8170 (N_8170,N_3428,N_1878);
nand U8171 (N_8171,N_3336,N_4665);
nor U8172 (N_8172,N_3464,N_1169);
and U8173 (N_8173,N_4831,N_163);
nand U8174 (N_8174,N_1634,N_1411);
nor U8175 (N_8175,N_2554,N_803);
xor U8176 (N_8176,N_2179,N_3991);
nand U8177 (N_8177,N_8,N_1879);
nand U8178 (N_8178,N_1570,N_1551);
nand U8179 (N_8179,N_107,N_2884);
or U8180 (N_8180,N_4425,N_4551);
and U8181 (N_8181,N_1158,N_1230);
nor U8182 (N_8182,N_793,N_457);
xor U8183 (N_8183,N_3597,N_3821);
nand U8184 (N_8184,N_3609,N_1757);
nor U8185 (N_8185,N_1909,N_3356);
nand U8186 (N_8186,N_1919,N_4967);
or U8187 (N_8187,N_4730,N_4731);
nor U8188 (N_8188,N_3911,N_4764);
or U8189 (N_8189,N_4365,N_744);
and U8190 (N_8190,N_2693,N_2016);
nor U8191 (N_8191,N_2936,N_1143);
nor U8192 (N_8192,N_705,N_1889);
nand U8193 (N_8193,N_66,N_202);
nand U8194 (N_8194,N_854,N_2895);
nor U8195 (N_8195,N_2508,N_3717);
nor U8196 (N_8196,N_2459,N_3306);
nand U8197 (N_8197,N_4361,N_3798);
or U8198 (N_8198,N_1737,N_218);
and U8199 (N_8199,N_1067,N_3300);
or U8200 (N_8200,N_128,N_4087);
or U8201 (N_8201,N_1241,N_1287);
or U8202 (N_8202,N_1366,N_3142);
or U8203 (N_8203,N_745,N_4293);
xor U8204 (N_8204,N_3322,N_308);
xor U8205 (N_8205,N_231,N_1544);
or U8206 (N_8206,N_2426,N_1728);
and U8207 (N_8207,N_1801,N_3048);
xor U8208 (N_8208,N_4922,N_2462);
nor U8209 (N_8209,N_2977,N_4625);
nor U8210 (N_8210,N_3470,N_1465);
and U8211 (N_8211,N_2337,N_4743);
nor U8212 (N_8212,N_1044,N_3325);
nand U8213 (N_8213,N_4684,N_2356);
nand U8214 (N_8214,N_3937,N_3342);
nand U8215 (N_8215,N_728,N_693);
xor U8216 (N_8216,N_1894,N_3838);
and U8217 (N_8217,N_1295,N_2938);
xor U8218 (N_8218,N_3645,N_188);
and U8219 (N_8219,N_1618,N_2754);
xor U8220 (N_8220,N_1602,N_4808);
or U8221 (N_8221,N_1678,N_1661);
or U8222 (N_8222,N_50,N_2195);
nand U8223 (N_8223,N_1248,N_3831);
and U8224 (N_8224,N_758,N_1587);
and U8225 (N_8225,N_2125,N_4689);
and U8226 (N_8226,N_4983,N_680);
and U8227 (N_8227,N_576,N_518);
and U8228 (N_8228,N_1885,N_2972);
nor U8229 (N_8229,N_4627,N_499);
and U8230 (N_8230,N_3583,N_3464);
or U8231 (N_8231,N_736,N_2965);
nand U8232 (N_8232,N_3367,N_4446);
or U8233 (N_8233,N_4327,N_4353);
and U8234 (N_8234,N_1223,N_1626);
xnor U8235 (N_8235,N_355,N_2466);
xnor U8236 (N_8236,N_488,N_2871);
nor U8237 (N_8237,N_2793,N_1820);
or U8238 (N_8238,N_4123,N_513);
nand U8239 (N_8239,N_4109,N_2833);
xnor U8240 (N_8240,N_4899,N_1070);
xor U8241 (N_8241,N_1036,N_3113);
nor U8242 (N_8242,N_3677,N_3674);
and U8243 (N_8243,N_3279,N_4652);
nor U8244 (N_8244,N_1696,N_980);
nand U8245 (N_8245,N_622,N_4029);
and U8246 (N_8246,N_400,N_1315);
nand U8247 (N_8247,N_4719,N_1078);
xnor U8248 (N_8248,N_2217,N_4450);
xnor U8249 (N_8249,N_2241,N_4548);
and U8250 (N_8250,N_2275,N_628);
nand U8251 (N_8251,N_3918,N_3117);
nor U8252 (N_8252,N_2424,N_1790);
nor U8253 (N_8253,N_1628,N_3273);
nor U8254 (N_8254,N_509,N_3583);
xor U8255 (N_8255,N_2337,N_1036);
nand U8256 (N_8256,N_216,N_3553);
nand U8257 (N_8257,N_590,N_3932);
and U8258 (N_8258,N_292,N_881);
xnor U8259 (N_8259,N_4609,N_4376);
nor U8260 (N_8260,N_2694,N_482);
and U8261 (N_8261,N_4709,N_2019);
and U8262 (N_8262,N_4994,N_1764);
or U8263 (N_8263,N_1555,N_3152);
and U8264 (N_8264,N_757,N_2911);
nand U8265 (N_8265,N_1347,N_3608);
xnor U8266 (N_8266,N_76,N_4184);
nand U8267 (N_8267,N_2788,N_1397);
and U8268 (N_8268,N_418,N_4311);
nand U8269 (N_8269,N_4401,N_2234);
nand U8270 (N_8270,N_964,N_3069);
nor U8271 (N_8271,N_1099,N_966);
or U8272 (N_8272,N_1762,N_4936);
nor U8273 (N_8273,N_771,N_1876);
nand U8274 (N_8274,N_3016,N_607);
or U8275 (N_8275,N_2773,N_3353);
and U8276 (N_8276,N_583,N_900);
or U8277 (N_8277,N_4511,N_412);
nor U8278 (N_8278,N_4969,N_1367);
and U8279 (N_8279,N_2304,N_2518);
xor U8280 (N_8280,N_2810,N_3613);
or U8281 (N_8281,N_3694,N_4868);
or U8282 (N_8282,N_30,N_3953);
nand U8283 (N_8283,N_1796,N_116);
or U8284 (N_8284,N_3282,N_1433);
nor U8285 (N_8285,N_3036,N_4739);
nand U8286 (N_8286,N_96,N_595);
or U8287 (N_8287,N_4565,N_1220);
or U8288 (N_8288,N_422,N_2586);
nor U8289 (N_8289,N_4346,N_4751);
nand U8290 (N_8290,N_3558,N_2747);
xnor U8291 (N_8291,N_533,N_2223);
or U8292 (N_8292,N_3417,N_3534);
or U8293 (N_8293,N_4174,N_1886);
or U8294 (N_8294,N_827,N_3058);
or U8295 (N_8295,N_3066,N_3599);
or U8296 (N_8296,N_4199,N_467);
nor U8297 (N_8297,N_1781,N_2464);
nor U8298 (N_8298,N_800,N_1019);
or U8299 (N_8299,N_3495,N_1237);
or U8300 (N_8300,N_4685,N_497);
nand U8301 (N_8301,N_723,N_4294);
xor U8302 (N_8302,N_698,N_1339);
nand U8303 (N_8303,N_4569,N_3691);
nor U8304 (N_8304,N_3042,N_3620);
nand U8305 (N_8305,N_241,N_222);
and U8306 (N_8306,N_1712,N_2996);
nor U8307 (N_8307,N_3090,N_2046);
nor U8308 (N_8308,N_344,N_2444);
nand U8309 (N_8309,N_4185,N_4382);
xnor U8310 (N_8310,N_4415,N_4178);
and U8311 (N_8311,N_3804,N_2912);
nand U8312 (N_8312,N_3059,N_3671);
xnor U8313 (N_8313,N_1194,N_1680);
nor U8314 (N_8314,N_4835,N_888);
nor U8315 (N_8315,N_2423,N_214);
and U8316 (N_8316,N_560,N_1915);
and U8317 (N_8317,N_2781,N_4344);
and U8318 (N_8318,N_2937,N_2444);
or U8319 (N_8319,N_3270,N_4660);
and U8320 (N_8320,N_3218,N_1810);
and U8321 (N_8321,N_532,N_309);
nand U8322 (N_8322,N_1487,N_2142);
nor U8323 (N_8323,N_1792,N_4590);
nand U8324 (N_8324,N_2621,N_3156);
and U8325 (N_8325,N_4634,N_900);
or U8326 (N_8326,N_1479,N_1520);
xor U8327 (N_8327,N_156,N_1300);
and U8328 (N_8328,N_4564,N_1295);
nand U8329 (N_8329,N_1688,N_716);
or U8330 (N_8330,N_80,N_3197);
and U8331 (N_8331,N_652,N_1167);
and U8332 (N_8332,N_4434,N_2911);
and U8333 (N_8333,N_3269,N_2713);
nor U8334 (N_8334,N_1609,N_4512);
nand U8335 (N_8335,N_2275,N_435);
and U8336 (N_8336,N_316,N_2129);
or U8337 (N_8337,N_3131,N_608);
and U8338 (N_8338,N_4943,N_1679);
nand U8339 (N_8339,N_2189,N_4886);
nand U8340 (N_8340,N_1928,N_337);
nor U8341 (N_8341,N_87,N_2851);
xor U8342 (N_8342,N_4056,N_4245);
nand U8343 (N_8343,N_4995,N_1004);
nor U8344 (N_8344,N_3858,N_2002);
nor U8345 (N_8345,N_3414,N_3925);
xnor U8346 (N_8346,N_3570,N_2959);
nor U8347 (N_8347,N_2976,N_2883);
nand U8348 (N_8348,N_4079,N_3368);
or U8349 (N_8349,N_554,N_3736);
or U8350 (N_8350,N_2739,N_3709);
and U8351 (N_8351,N_4783,N_2994);
and U8352 (N_8352,N_2576,N_2033);
or U8353 (N_8353,N_2107,N_1431);
or U8354 (N_8354,N_2199,N_437);
and U8355 (N_8355,N_1811,N_3473);
or U8356 (N_8356,N_3112,N_4668);
nand U8357 (N_8357,N_2785,N_1184);
or U8358 (N_8358,N_435,N_1741);
and U8359 (N_8359,N_2789,N_4404);
and U8360 (N_8360,N_986,N_3676);
or U8361 (N_8361,N_782,N_3867);
nor U8362 (N_8362,N_280,N_1525);
xnor U8363 (N_8363,N_891,N_1919);
xnor U8364 (N_8364,N_1465,N_2775);
and U8365 (N_8365,N_2445,N_512);
nand U8366 (N_8366,N_4890,N_2904);
or U8367 (N_8367,N_3350,N_766);
and U8368 (N_8368,N_554,N_1504);
or U8369 (N_8369,N_3718,N_4695);
nor U8370 (N_8370,N_758,N_3332);
or U8371 (N_8371,N_4083,N_2665);
and U8372 (N_8372,N_4093,N_3839);
and U8373 (N_8373,N_2850,N_3878);
xnor U8374 (N_8374,N_3226,N_1803);
nor U8375 (N_8375,N_4031,N_91);
nor U8376 (N_8376,N_567,N_2947);
nor U8377 (N_8377,N_27,N_3586);
and U8378 (N_8378,N_4271,N_479);
and U8379 (N_8379,N_4836,N_481);
nor U8380 (N_8380,N_4281,N_3502);
nor U8381 (N_8381,N_1753,N_2843);
nor U8382 (N_8382,N_1711,N_3826);
nor U8383 (N_8383,N_4544,N_1950);
nand U8384 (N_8384,N_3910,N_3572);
and U8385 (N_8385,N_3262,N_3247);
nand U8386 (N_8386,N_1839,N_3186);
nor U8387 (N_8387,N_4154,N_950);
nor U8388 (N_8388,N_1242,N_2174);
and U8389 (N_8389,N_4323,N_2503);
xnor U8390 (N_8390,N_4784,N_1980);
or U8391 (N_8391,N_3265,N_2578);
and U8392 (N_8392,N_1,N_1622);
or U8393 (N_8393,N_4812,N_385);
and U8394 (N_8394,N_1940,N_4735);
xnor U8395 (N_8395,N_1600,N_2392);
xnor U8396 (N_8396,N_3316,N_3274);
nor U8397 (N_8397,N_2504,N_1163);
nand U8398 (N_8398,N_2169,N_4988);
nand U8399 (N_8399,N_2992,N_4193);
and U8400 (N_8400,N_553,N_457);
nor U8401 (N_8401,N_4953,N_2419);
nor U8402 (N_8402,N_1557,N_298);
and U8403 (N_8403,N_3378,N_3153);
or U8404 (N_8404,N_479,N_2427);
nor U8405 (N_8405,N_201,N_4911);
and U8406 (N_8406,N_994,N_2594);
nand U8407 (N_8407,N_165,N_3016);
nor U8408 (N_8408,N_2369,N_3873);
nand U8409 (N_8409,N_3500,N_369);
nand U8410 (N_8410,N_59,N_1797);
nor U8411 (N_8411,N_537,N_218);
or U8412 (N_8412,N_2303,N_3668);
xor U8413 (N_8413,N_4293,N_3696);
nand U8414 (N_8414,N_1526,N_357);
and U8415 (N_8415,N_2053,N_3000);
and U8416 (N_8416,N_237,N_2120);
nand U8417 (N_8417,N_4743,N_4321);
xnor U8418 (N_8418,N_1421,N_4967);
and U8419 (N_8419,N_3535,N_1006);
or U8420 (N_8420,N_2226,N_408);
and U8421 (N_8421,N_1630,N_1317);
nand U8422 (N_8422,N_1197,N_3582);
and U8423 (N_8423,N_4119,N_286);
and U8424 (N_8424,N_883,N_4364);
nand U8425 (N_8425,N_1793,N_1415);
and U8426 (N_8426,N_4241,N_4963);
or U8427 (N_8427,N_2418,N_3102);
and U8428 (N_8428,N_2274,N_4834);
nor U8429 (N_8429,N_3851,N_3321);
nor U8430 (N_8430,N_4968,N_2692);
and U8431 (N_8431,N_4933,N_4039);
nor U8432 (N_8432,N_4558,N_2688);
nor U8433 (N_8433,N_2810,N_920);
nor U8434 (N_8434,N_4665,N_3616);
xor U8435 (N_8435,N_3239,N_3993);
and U8436 (N_8436,N_1096,N_991);
xor U8437 (N_8437,N_4480,N_4506);
or U8438 (N_8438,N_2373,N_521);
nor U8439 (N_8439,N_2930,N_4783);
or U8440 (N_8440,N_2724,N_3107);
xor U8441 (N_8441,N_4484,N_3533);
or U8442 (N_8442,N_1708,N_3096);
nor U8443 (N_8443,N_3005,N_3541);
nand U8444 (N_8444,N_2721,N_276);
nand U8445 (N_8445,N_3145,N_2370);
nor U8446 (N_8446,N_836,N_4133);
nor U8447 (N_8447,N_4577,N_3274);
nand U8448 (N_8448,N_2762,N_1296);
and U8449 (N_8449,N_3492,N_1045);
and U8450 (N_8450,N_1897,N_481);
nand U8451 (N_8451,N_1297,N_3889);
and U8452 (N_8452,N_3224,N_1344);
nor U8453 (N_8453,N_3449,N_1740);
and U8454 (N_8454,N_3156,N_4921);
xnor U8455 (N_8455,N_1468,N_4489);
nand U8456 (N_8456,N_2344,N_1574);
nand U8457 (N_8457,N_3555,N_3947);
nor U8458 (N_8458,N_229,N_4577);
nor U8459 (N_8459,N_4623,N_1526);
and U8460 (N_8460,N_2224,N_3305);
or U8461 (N_8461,N_4266,N_1909);
nor U8462 (N_8462,N_3188,N_2088);
or U8463 (N_8463,N_2847,N_4653);
nand U8464 (N_8464,N_3211,N_4002);
and U8465 (N_8465,N_3855,N_1580);
and U8466 (N_8466,N_4935,N_1106);
nor U8467 (N_8467,N_971,N_4496);
and U8468 (N_8468,N_1380,N_1719);
nand U8469 (N_8469,N_3423,N_2690);
nor U8470 (N_8470,N_827,N_1255);
nor U8471 (N_8471,N_3395,N_4123);
or U8472 (N_8472,N_4462,N_1867);
nand U8473 (N_8473,N_1474,N_3736);
nor U8474 (N_8474,N_1093,N_3547);
or U8475 (N_8475,N_3697,N_3101);
nor U8476 (N_8476,N_3464,N_3961);
nand U8477 (N_8477,N_4985,N_769);
xor U8478 (N_8478,N_774,N_4571);
nand U8479 (N_8479,N_3701,N_488);
or U8480 (N_8480,N_3156,N_622);
and U8481 (N_8481,N_3080,N_110);
nor U8482 (N_8482,N_4529,N_1481);
nand U8483 (N_8483,N_3716,N_288);
and U8484 (N_8484,N_1898,N_2389);
or U8485 (N_8485,N_327,N_3522);
or U8486 (N_8486,N_1955,N_2816);
nand U8487 (N_8487,N_4505,N_1879);
and U8488 (N_8488,N_2945,N_3060);
and U8489 (N_8489,N_1333,N_4954);
and U8490 (N_8490,N_4214,N_3857);
nand U8491 (N_8491,N_515,N_1280);
or U8492 (N_8492,N_4346,N_2606);
nand U8493 (N_8493,N_3349,N_2545);
nand U8494 (N_8494,N_1143,N_1824);
and U8495 (N_8495,N_772,N_2139);
and U8496 (N_8496,N_4192,N_809);
nor U8497 (N_8497,N_3542,N_70);
or U8498 (N_8498,N_1371,N_3249);
nor U8499 (N_8499,N_1056,N_187);
nor U8500 (N_8500,N_656,N_3163);
and U8501 (N_8501,N_339,N_4317);
nor U8502 (N_8502,N_3628,N_4479);
or U8503 (N_8503,N_294,N_335);
and U8504 (N_8504,N_1041,N_1295);
nand U8505 (N_8505,N_818,N_3406);
and U8506 (N_8506,N_1330,N_2190);
and U8507 (N_8507,N_2312,N_563);
xnor U8508 (N_8508,N_1652,N_3354);
and U8509 (N_8509,N_773,N_4556);
or U8510 (N_8510,N_3710,N_298);
nor U8511 (N_8511,N_760,N_354);
and U8512 (N_8512,N_1806,N_4622);
nand U8513 (N_8513,N_3105,N_921);
xor U8514 (N_8514,N_3947,N_56);
and U8515 (N_8515,N_697,N_2335);
nand U8516 (N_8516,N_577,N_4887);
nand U8517 (N_8517,N_3647,N_2664);
nand U8518 (N_8518,N_3378,N_4887);
or U8519 (N_8519,N_938,N_3062);
nor U8520 (N_8520,N_2064,N_2074);
nand U8521 (N_8521,N_2247,N_3553);
or U8522 (N_8522,N_3414,N_1314);
and U8523 (N_8523,N_680,N_1261);
or U8524 (N_8524,N_851,N_4618);
nand U8525 (N_8525,N_1230,N_1067);
or U8526 (N_8526,N_865,N_3874);
and U8527 (N_8527,N_4067,N_3109);
nand U8528 (N_8528,N_4719,N_2158);
or U8529 (N_8529,N_3970,N_3247);
nor U8530 (N_8530,N_1392,N_1385);
xnor U8531 (N_8531,N_498,N_3672);
and U8532 (N_8532,N_3320,N_1198);
nand U8533 (N_8533,N_2297,N_1576);
and U8534 (N_8534,N_3776,N_2756);
or U8535 (N_8535,N_2607,N_4470);
nor U8536 (N_8536,N_2518,N_3360);
nor U8537 (N_8537,N_3367,N_1235);
nor U8538 (N_8538,N_4130,N_3642);
or U8539 (N_8539,N_3814,N_4675);
nand U8540 (N_8540,N_3819,N_1705);
and U8541 (N_8541,N_1572,N_1902);
and U8542 (N_8542,N_4762,N_342);
or U8543 (N_8543,N_3285,N_4172);
nand U8544 (N_8544,N_3367,N_1956);
nand U8545 (N_8545,N_1959,N_3884);
and U8546 (N_8546,N_3313,N_4935);
xor U8547 (N_8547,N_907,N_4698);
nor U8548 (N_8548,N_2806,N_2990);
or U8549 (N_8549,N_218,N_861);
or U8550 (N_8550,N_1754,N_3576);
nand U8551 (N_8551,N_4990,N_2551);
and U8552 (N_8552,N_4490,N_2526);
nand U8553 (N_8553,N_4955,N_3432);
nand U8554 (N_8554,N_4876,N_4426);
nand U8555 (N_8555,N_4534,N_4484);
and U8556 (N_8556,N_2187,N_3802);
nand U8557 (N_8557,N_3054,N_1673);
and U8558 (N_8558,N_1763,N_2004);
nand U8559 (N_8559,N_3298,N_2648);
nand U8560 (N_8560,N_3529,N_2501);
xor U8561 (N_8561,N_1233,N_4466);
and U8562 (N_8562,N_886,N_2340);
or U8563 (N_8563,N_1047,N_4711);
nor U8564 (N_8564,N_3012,N_1120);
and U8565 (N_8565,N_1096,N_4120);
and U8566 (N_8566,N_4095,N_4701);
nand U8567 (N_8567,N_3645,N_4988);
or U8568 (N_8568,N_4360,N_3943);
and U8569 (N_8569,N_3581,N_3013);
nor U8570 (N_8570,N_441,N_913);
nor U8571 (N_8571,N_3330,N_201);
and U8572 (N_8572,N_2522,N_2011);
and U8573 (N_8573,N_2123,N_2886);
and U8574 (N_8574,N_4518,N_1891);
nor U8575 (N_8575,N_4163,N_4608);
or U8576 (N_8576,N_2948,N_2482);
nand U8577 (N_8577,N_3976,N_4034);
or U8578 (N_8578,N_4358,N_3216);
and U8579 (N_8579,N_4170,N_3378);
or U8580 (N_8580,N_4236,N_114);
or U8581 (N_8581,N_2987,N_1611);
nor U8582 (N_8582,N_518,N_4252);
nand U8583 (N_8583,N_2886,N_3322);
or U8584 (N_8584,N_4115,N_4442);
and U8585 (N_8585,N_3973,N_3931);
or U8586 (N_8586,N_2950,N_4364);
nor U8587 (N_8587,N_88,N_2042);
nand U8588 (N_8588,N_1327,N_4719);
or U8589 (N_8589,N_2232,N_3675);
nor U8590 (N_8590,N_2501,N_4641);
and U8591 (N_8591,N_4884,N_427);
nor U8592 (N_8592,N_682,N_3600);
and U8593 (N_8593,N_132,N_112);
nor U8594 (N_8594,N_2060,N_4809);
xor U8595 (N_8595,N_4220,N_2681);
and U8596 (N_8596,N_1714,N_1368);
or U8597 (N_8597,N_267,N_223);
nand U8598 (N_8598,N_3213,N_2078);
nand U8599 (N_8599,N_386,N_4941);
nor U8600 (N_8600,N_2713,N_2546);
and U8601 (N_8601,N_2873,N_4312);
and U8602 (N_8602,N_4140,N_3279);
or U8603 (N_8603,N_3906,N_4701);
or U8604 (N_8604,N_4193,N_2596);
and U8605 (N_8605,N_1018,N_2220);
nand U8606 (N_8606,N_3140,N_3762);
nor U8607 (N_8607,N_1343,N_382);
xnor U8608 (N_8608,N_1345,N_2397);
and U8609 (N_8609,N_54,N_2349);
or U8610 (N_8610,N_1007,N_1035);
or U8611 (N_8611,N_4707,N_3104);
nand U8612 (N_8612,N_2226,N_3489);
nand U8613 (N_8613,N_3647,N_4449);
and U8614 (N_8614,N_913,N_344);
xor U8615 (N_8615,N_2545,N_3752);
or U8616 (N_8616,N_2091,N_2418);
or U8617 (N_8617,N_4901,N_820);
xnor U8618 (N_8618,N_1580,N_4045);
or U8619 (N_8619,N_2864,N_4882);
or U8620 (N_8620,N_1383,N_3255);
and U8621 (N_8621,N_4326,N_1143);
and U8622 (N_8622,N_1467,N_2063);
or U8623 (N_8623,N_4764,N_2622);
nand U8624 (N_8624,N_917,N_799);
and U8625 (N_8625,N_4857,N_4228);
and U8626 (N_8626,N_4495,N_50);
and U8627 (N_8627,N_1975,N_2801);
or U8628 (N_8628,N_1758,N_1865);
or U8629 (N_8629,N_2054,N_3519);
and U8630 (N_8630,N_4300,N_1604);
or U8631 (N_8631,N_2817,N_861);
nor U8632 (N_8632,N_661,N_4896);
nand U8633 (N_8633,N_1945,N_1702);
or U8634 (N_8634,N_4029,N_4267);
xnor U8635 (N_8635,N_221,N_2999);
or U8636 (N_8636,N_695,N_3499);
nand U8637 (N_8637,N_4753,N_438);
or U8638 (N_8638,N_4434,N_3830);
nor U8639 (N_8639,N_2337,N_4669);
xnor U8640 (N_8640,N_4970,N_2783);
nor U8641 (N_8641,N_2945,N_4690);
and U8642 (N_8642,N_534,N_2682);
nor U8643 (N_8643,N_654,N_673);
and U8644 (N_8644,N_2916,N_2945);
nor U8645 (N_8645,N_4472,N_3012);
or U8646 (N_8646,N_3214,N_4211);
nor U8647 (N_8647,N_3413,N_293);
nor U8648 (N_8648,N_4395,N_3513);
xor U8649 (N_8649,N_4267,N_2700);
and U8650 (N_8650,N_3073,N_3402);
or U8651 (N_8651,N_297,N_1653);
nor U8652 (N_8652,N_2692,N_1680);
or U8653 (N_8653,N_4679,N_1610);
nand U8654 (N_8654,N_3116,N_2397);
xnor U8655 (N_8655,N_865,N_268);
and U8656 (N_8656,N_2584,N_577);
or U8657 (N_8657,N_130,N_2763);
nand U8658 (N_8658,N_3152,N_4290);
or U8659 (N_8659,N_3770,N_4531);
nand U8660 (N_8660,N_3274,N_3525);
or U8661 (N_8661,N_1284,N_2572);
nor U8662 (N_8662,N_834,N_4841);
xor U8663 (N_8663,N_2763,N_929);
nand U8664 (N_8664,N_2218,N_2576);
or U8665 (N_8665,N_4499,N_3185);
nor U8666 (N_8666,N_283,N_895);
nand U8667 (N_8667,N_4597,N_3197);
and U8668 (N_8668,N_581,N_3681);
nor U8669 (N_8669,N_4485,N_1297);
xor U8670 (N_8670,N_1161,N_3881);
and U8671 (N_8671,N_4173,N_3559);
xor U8672 (N_8672,N_1546,N_3106);
nand U8673 (N_8673,N_2323,N_3458);
xor U8674 (N_8674,N_2398,N_916);
or U8675 (N_8675,N_3435,N_305);
xnor U8676 (N_8676,N_407,N_638);
nand U8677 (N_8677,N_4127,N_943);
and U8678 (N_8678,N_1992,N_2738);
nand U8679 (N_8679,N_1735,N_1705);
nor U8680 (N_8680,N_1020,N_2857);
nor U8681 (N_8681,N_4415,N_2537);
nor U8682 (N_8682,N_4116,N_2565);
and U8683 (N_8683,N_424,N_2833);
nand U8684 (N_8684,N_4401,N_3730);
nand U8685 (N_8685,N_1552,N_4471);
and U8686 (N_8686,N_2041,N_1702);
or U8687 (N_8687,N_1397,N_931);
nor U8688 (N_8688,N_3485,N_4906);
and U8689 (N_8689,N_877,N_377);
nand U8690 (N_8690,N_886,N_4858);
and U8691 (N_8691,N_402,N_2991);
xnor U8692 (N_8692,N_591,N_2103);
or U8693 (N_8693,N_1926,N_852);
nor U8694 (N_8694,N_2837,N_935);
nand U8695 (N_8695,N_504,N_491);
and U8696 (N_8696,N_3969,N_2349);
nand U8697 (N_8697,N_4260,N_2838);
and U8698 (N_8698,N_4712,N_1254);
nor U8699 (N_8699,N_1808,N_442);
nand U8700 (N_8700,N_589,N_836);
nand U8701 (N_8701,N_4718,N_267);
nand U8702 (N_8702,N_767,N_1068);
nand U8703 (N_8703,N_1296,N_1489);
nand U8704 (N_8704,N_169,N_4971);
and U8705 (N_8705,N_3314,N_971);
nor U8706 (N_8706,N_1036,N_2499);
nand U8707 (N_8707,N_293,N_2056);
nand U8708 (N_8708,N_3906,N_1728);
or U8709 (N_8709,N_3493,N_2904);
or U8710 (N_8710,N_4065,N_936);
nand U8711 (N_8711,N_4200,N_2462);
nand U8712 (N_8712,N_3145,N_584);
nor U8713 (N_8713,N_1899,N_4691);
nor U8714 (N_8714,N_2874,N_1969);
and U8715 (N_8715,N_386,N_2883);
nor U8716 (N_8716,N_4575,N_2214);
nand U8717 (N_8717,N_2660,N_369);
xor U8718 (N_8718,N_1214,N_2327);
xnor U8719 (N_8719,N_4793,N_4494);
nor U8720 (N_8720,N_1897,N_74);
and U8721 (N_8721,N_2591,N_3908);
or U8722 (N_8722,N_4956,N_238);
nand U8723 (N_8723,N_4749,N_3967);
nand U8724 (N_8724,N_2039,N_3855);
or U8725 (N_8725,N_434,N_1812);
nand U8726 (N_8726,N_3405,N_4887);
and U8727 (N_8727,N_706,N_1073);
and U8728 (N_8728,N_1495,N_3485);
and U8729 (N_8729,N_107,N_299);
and U8730 (N_8730,N_2254,N_1753);
nor U8731 (N_8731,N_4312,N_1203);
and U8732 (N_8732,N_3040,N_507);
and U8733 (N_8733,N_4571,N_146);
nor U8734 (N_8734,N_968,N_1113);
and U8735 (N_8735,N_890,N_3654);
or U8736 (N_8736,N_1588,N_1913);
and U8737 (N_8737,N_2050,N_3564);
and U8738 (N_8738,N_2455,N_1189);
xor U8739 (N_8739,N_957,N_2719);
nand U8740 (N_8740,N_3910,N_1651);
nand U8741 (N_8741,N_2176,N_4035);
and U8742 (N_8742,N_1661,N_1128);
nor U8743 (N_8743,N_4786,N_2891);
and U8744 (N_8744,N_740,N_216);
and U8745 (N_8745,N_4890,N_2242);
nand U8746 (N_8746,N_4633,N_885);
xnor U8747 (N_8747,N_989,N_2735);
nand U8748 (N_8748,N_4161,N_2506);
nand U8749 (N_8749,N_174,N_2743);
nand U8750 (N_8750,N_4062,N_3659);
and U8751 (N_8751,N_1383,N_4499);
or U8752 (N_8752,N_949,N_3020);
nand U8753 (N_8753,N_2538,N_2898);
and U8754 (N_8754,N_1559,N_1986);
nor U8755 (N_8755,N_3704,N_4399);
nor U8756 (N_8756,N_2660,N_3993);
and U8757 (N_8757,N_664,N_3504);
xor U8758 (N_8758,N_4015,N_91);
nor U8759 (N_8759,N_2033,N_3382);
nor U8760 (N_8760,N_786,N_4146);
nor U8761 (N_8761,N_3887,N_1735);
or U8762 (N_8762,N_4708,N_2886);
or U8763 (N_8763,N_2330,N_3434);
or U8764 (N_8764,N_1081,N_4476);
nor U8765 (N_8765,N_4825,N_4238);
nor U8766 (N_8766,N_956,N_4010);
or U8767 (N_8767,N_4065,N_1762);
and U8768 (N_8768,N_2392,N_705);
xnor U8769 (N_8769,N_173,N_675);
or U8770 (N_8770,N_4596,N_124);
nand U8771 (N_8771,N_2689,N_1524);
nor U8772 (N_8772,N_1916,N_2472);
nand U8773 (N_8773,N_3675,N_3817);
and U8774 (N_8774,N_1088,N_109);
and U8775 (N_8775,N_251,N_2953);
or U8776 (N_8776,N_998,N_1095);
or U8777 (N_8777,N_66,N_2701);
and U8778 (N_8778,N_3411,N_1821);
or U8779 (N_8779,N_2249,N_3503);
or U8780 (N_8780,N_3269,N_2449);
and U8781 (N_8781,N_2860,N_2610);
and U8782 (N_8782,N_3583,N_2208);
nand U8783 (N_8783,N_4129,N_2183);
or U8784 (N_8784,N_3399,N_1229);
and U8785 (N_8785,N_436,N_689);
nand U8786 (N_8786,N_2459,N_1658);
and U8787 (N_8787,N_2005,N_4881);
xnor U8788 (N_8788,N_2704,N_2590);
nor U8789 (N_8789,N_3639,N_4593);
xnor U8790 (N_8790,N_3678,N_3331);
nand U8791 (N_8791,N_2096,N_1649);
or U8792 (N_8792,N_1025,N_3019);
or U8793 (N_8793,N_2617,N_4853);
nand U8794 (N_8794,N_2717,N_3758);
and U8795 (N_8795,N_1542,N_3914);
nor U8796 (N_8796,N_3099,N_1184);
nor U8797 (N_8797,N_2319,N_44);
or U8798 (N_8798,N_1719,N_1292);
and U8799 (N_8799,N_1976,N_2156);
xnor U8800 (N_8800,N_90,N_39);
nor U8801 (N_8801,N_2871,N_1583);
nor U8802 (N_8802,N_4193,N_4678);
xor U8803 (N_8803,N_21,N_359);
nand U8804 (N_8804,N_4641,N_3144);
nand U8805 (N_8805,N_183,N_553);
and U8806 (N_8806,N_2507,N_2230);
or U8807 (N_8807,N_2886,N_3300);
nor U8808 (N_8808,N_1584,N_3341);
nand U8809 (N_8809,N_2214,N_2189);
or U8810 (N_8810,N_2855,N_2160);
nor U8811 (N_8811,N_903,N_1552);
or U8812 (N_8812,N_335,N_3976);
nand U8813 (N_8813,N_3698,N_4896);
and U8814 (N_8814,N_3619,N_4271);
and U8815 (N_8815,N_263,N_1744);
nor U8816 (N_8816,N_4390,N_3983);
or U8817 (N_8817,N_1159,N_1943);
nand U8818 (N_8818,N_3014,N_1708);
and U8819 (N_8819,N_516,N_1154);
nor U8820 (N_8820,N_3670,N_2873);
xor U8821 (N_8821,N_4717,N_4397);
nand U8822 (N_8822,N_1961,N_4993);
xnor U8823 (N_8823,N_1576,N_1210);
nor U8824 (N_8824,N_419,N_2084);
nand U8825 (N_8825,N_3253,N_3884);
xor U8826 (N_8826,N_3423,N_2649);
xor U8827 (N_8827,N_1992,N_2922);
nor U8828 (N_8828,N_4761,N_860);
nor U8829 (N_8829,N_4683,N_1774);
nor U8830 (N_8830,N_1714,N_424);
nand U8831 (N_8831,N_3090,N_3886);
or U8832 (N_8832,N_3631,N_227);
nand U8833 (N_8833,N_2598,N_746);
or U8834 (N_8834,N_3754,N_4797);
nor U8835 (N_8835,N_2644,N_2753);
nor U8836 (N_8836,N_4224,N_4640);
and U8837 (N_8837,N_3560,N_3249);
nand U8838 (N_8838,N_4858,N_3464);
or U8839 (N_8839,N_4006,N_1945);
nand U8840 (N_8840,N_2761,N_2605);
xnor U8841 (N_8841,N_2822,N_3723);
or U8842 (N_8842,N_225,N_2306);
and U8843 (N_8843,N_2533,N_4240);
and U8844 (N_8844,N_2702,N_1305);
or U8845 (N_8845,N_111,N_4742);
or U8846 (N_8846,N_2083,N_1900);
xor U8847 (N_8847,N_4156,N_3156);
nand U8848 (N_8848,N_4468,N_1969);
or U8849 (N_8849,N_4833,N_3908);
nand U8850 (N_8850,N_1948,N_456);
nor U8851 (N_8851,N_1044,N_848);
nor U8852 (N_8852,N_3381,N_3402);
nand U8853 (N_8853,N_258,N_1160);
nor U8854 (N_8854,N_1347,N_4699);
nor U8855 (N_8855,N_1978,N_4611);
and U8856 (N_8856,N_4301,N_4449);
and U8857 (N_8857,N_251,N_35);
nor U8858 (N_8858,N_3280,N_4281);
xnor U8859 (N_8859,N_562,N_1332);
nand U8860 (N_8860,N_3818,N_3941);
or U8861 (N_8861,N_1106,N_1481);
nor U8862 (N_8862,N_2225,N_1474);
or U8863 (N_8863,N_1262,N_3834);
xnor U8864 (N_8864,N_4625,N_1053);
nor U8865 (N_8865,N_4290,N_2114);
nand U8866 (N_8866,N_245,N_1904);
nor U8867 (N_8867,N_4238,N_370);
xor U8868 (N_8868,N_2092,N_853);
nand U8869 (N_8869,N_870,N_2766);
and U8870 (N_8870,N_3723,N_2737);
nand U8871 (N_8871,N_3530,N_3827);
or U8872 (N_8872,N_1556,N_2185);
or U8873 (N_8873,N_3575,N_1400);
nand U8874 (N_8874,N_2412,N_3753);
or U8875 (N_8875,N_3047,N_899);
nand U8876 (N_8876,N_1455,N_2152);
or U8877 (N_8877,N_13,N_2675);
xor U8878 (N_8878,N_659,N_3286);
nand U8879 (N_8879,N_573,N_2493);
and U8880 (N_8880,N_3363,N_611);
nor U8881 (N_8881,N_1878,N_2739);
xnor U8882 (N_8882,N_3490,N_3063);
or U8883 (N_8883,N_3926,N_449);
and U8884 (N_8884,N_4446,N_1610);
nor U8885 (N_8885,N_854,N_2798);
and U8886 (N_8886,N_3854,N_1717);
and U8887 (N_8887,N_311,N_4273);
or U8888 (N_8888,N_3489,N_3274);
nand U8889 (N_8889,N_4249,N_3537);
or U8890 (N_8890,N_288,N_3100);
or U8891 (N_8891,N_2301,N_2969);
xnor U8892 (N_8892,N_3731,N_2399);
nor U8893 (N_8893,N_2181,N_558);
nor U8894 (N_8894,N_4573,N_329);
nand U8895 (N_8895,N_3049,N_4050);
nand U8896 (N_8896,N_4834,N_3145);
and U8897 (N_8897,N_126,N_4218);
nand U8898 (N_8898,N_3900,N_2065);
and U8899 (N_8899,N_1291,N_4767);
nor U8900 (N_8900,N_1526,N_790);
nor U8901 (N_8901,N_4536,N_2697);
nor U8902 (N_8902,N_562,N_75);
or U8903 (N_8903,N_4385,N_4848);
nor U8904 (N_8904,N_440,N_4321);
nand U8905 (N_8905,N_4786,N_4946);
nor U8906 (N_8906,N_2417,N_1759);
nand U8907 (N_8907,N_4920,N_3666);
nand U8908 (N_8908,N_3950,N_115);
nand U8909 (N_8909,N_993,N_3568);
nand U8910 (N_8910,N_4056,N_980);
nor U8911 (N_8911,N_2645,N_2888);
nand U8912 (N_8912,N_1963,N_2280);
and U8913 (N_8913,N_3424,N_4017);
and U8914 (N_8914,N_1480,N_3454);
nand U8915 (N_8915,N_2955,N_1082);
nand U8916 (N_8916,N_4783,N_123);
xnor U8917 (N_8917,N_1908,N_1097);
and U8918 (N_8918,N_1601,N_3256);
nor U8919 (N_8919,N_1270,N_3717);
or U8920 (N_8920,N_4080,N_3952);
xor U8921 (N_8921,N_2104,N_2228);
nor U8922 (N_8922,N_1401,N_1395);
nand U8923 (N_8923,N_2341,N_867);
xnor U8924 (N_8924,N_4014,N_1874);
nor U8925 (N_8925,N_1784,N_1637);
or U8926 (N_8926,N_3267,N_535);
nor U8927 (N_8927,N_1978,N_4825);
nand U8928 (N_8928,N_4177,N_3834);
nor U8929 (N_8929,N_3901,N_2134);
nor U8930 (N_8930,N_2704,N_2364);
or U8931 (N_8931,N_2108,N_4778);
nand U8932 (N_8932,N_767,N_4641);
and U8933 (N_8933,N_2920,N_4495);
xor U8934 (N_8934,N_3556,N_1362);
nand U8935 (N_8935,N_342,N_1482);
xor U8936 (N_8936,N_2416,N_1508);
nor U8937 (N_8937,N_952,N_3099);
nand U8938 (N_8938,N_2339,N_3041);
or U8939 (N_8939,N_2657,N_1011);
and U8940 (N_8940,N_2694,N_4428);
xor U8941 (N_8941,N_3754,N_2092);
or U8942 (N_8942,N_2358,N_1423);
nand U8943 (N_8943,N_2008,N_2614);
nor U8944 (N_8944,N_299,N_1015);
xnor U8945 (N_8945,N_4296,N_611);
or U8946 (N_8946,N_3413,N_1365);
and U8947 (N_8947,N_360,N_3378);
and U8948 (N_8948,N_1807,N_913);
nor U8949 (N_8949,N_4918,N_4579);
nand U8950 (N_8950,N_4121,N_2735);
or U8951 (N_8951,N_1939,N_545);
and U8952 (N_8952,N_2868,N_2274);
nor U8953 (N_8953,N_3104,N_2961);
nand U8954 (N_8954,N_4879,N_3129);
nand U8955 (N_8955,N_4075,N_3044);
and U8956 (N_8956,N_141,N_543);
and U8957 (N_8957,N_3283,N_35);
nand U8958 (N_8958,N_1868,N_1117);
nor U8959 (N_8959,N_1375,N_2855);
or U8960 (N_8960,N_2210,N_94);
xnor U8961 (N_8961,N_4632,N_654);
and U8962 (N_8962,N_3775,N_4818);
or U8963 (N_8963,N_3335,N_772);
or U8964 (N_8964,N_425,N_3676);
or U8965 (N_8965,N_4964,N_4484);
or U8966 (N_8966,N_4206,N_1916);
or U8967 (N_8967,N_4993,N_570);
nor U8968 (N_8968,N_2791,N_1534);
nand U8969 (N_8969,N_2421,N_796);
nand U8970 (N_8970,N_3412,N_4963);
xor U8971 (N_8971,N_4700,N_437);
and U8972 (N_8972,N_4314,N_2847);
nand U8973 (N_8973,N_1523,N_892);
and U8974 (N_8974,N_1032,N_4614);
xor U8975 (N_8975,N_4976,N_1649);
xnor U8976 (N_8976,N_2179,N_3091);
nand U8977 (N_8977,N_4436,N_802);
nor U8978 (N_8978,N_237,N_1134);
nor U8979 (N_8979,N_1591,N_73);
or U8980 (N_8980,N_2318,N_2873);
and U8981 (N_8981,N_3251,N_1456);
nand U8982 (N_8982,N_3701,N_570);
or U8983 (N_8983,N_1479,N_237);
or U8984 (N_8984,N_3745,N_1172);
or U8985 (N_8985,N_4666,N_295);
nand U8986 (N_8986,N_4012,N_3443);
nand U8987 (N_8987,N_291,N_4696);
and U8988 (N_8988,N_1720,N_3559);
nand U8989 (N_8989,N_3965,N_1009);
nand U8990 (N_8990,N_1411,N_3438);
xor U8991 (N_8991,N_3659,N_2030);
nand U8992 (N_8992,N_3173,N_143);
nor U8993 (N_8993,N_1731,N_4884);
nand U8994 (N_8994,N_1172,N_1370);
nand U8995 (N_8995,N_2097,N_394);
or U8996 (N_8996,N_515,N_1581);
or U8997 (N_8997,N_4388,N_2725);
nor U8998 (N_8998,N_4388,N_2720);
or U8999 (N_8999,N_3223,N_4921);
nand U9000 (N_9000,N_1918,N_1571);
or U9001 (N_9001,N_3379,N_1221);
nand U9002 (N_9002,N_2676,N_3187);
and U9003 (N_9003,N_3810,N_2533);
nand U9004 (N_9004,N_3546,N_459);
nand U9005 (N_9005,N_1161,N_4316);
xnor U9006 (N_9006,N_4171,N_1130);
nand U9007 (N_9007,N_945,N_2492);
nor U9008 (N_9008,N_1687,N_1169);
and U9009 (N_9009,N_3921,N_4356);
xor U9010 (N_9010,N_4417,N_4858);
nor U9011 (N_9011,N_1780,N_348);
and U9012 (N_9012,N_2214,N_1306);
nand U9013 (N_9013,N_4331,N_4404);
and U9014 (N_9014,N_373,N_1667);
and U9015 (N_9015,N_2253,N_2056);
and U9016 (N_9016,N_3962,N_2693);
and U9017 (N_9017,N_4923,N_4538);
nor U9018 (N_9018,N_23,N_4085);
nand U9019 (N_9019,N_2966,N_2429);
nand U9020 (N_9020,N_645,N_3903);
nand U9021 (N_9021,N_2792,N_695);
nand U9022 (N_9022,N_3425,N_3706);
nor U9023 (N_9023,N_816,N_3625);
nor U9024 (N_9024,N_809,N_1968);
nor U9025 (N_9025,N_1045,N_3875);
nand U9026 (N_9026,N_838,N_1482);
xnor U9027 (N_9027,N_3765,N_3821);
or U9028 (N_9028,N_3654,N_2307);
nor U9029 (N_9029,N_3036,N_594);
or U9030 (N_9030,N_2514,N_4017);
or U9031 (N_9031,N_717,N_1289);
nand U9032 (N_9032,N_51,N_932);
and U9033 (N_9033,N_184,N_1674);
nor U9034 (N_9034,N_3149,N_4977);
nor U9035 (N_9035,N_4255,N_3138);
xnor U9036 (N_9036,N_1107,N_2885);
or U9037 (N_9037,N_3128,N_2950);
or U9038 (N_9038,N_897,N_4455);
nor U9039 (N_9039,N_2236,N_2866);
nand U9040 (N_9040,N_2873,N_2773);
xor U9041 (N_9041,N_2770,N_2323);
and U9042 (N_9042,N_753,N_618);
xnor U9043 (N_9043,N_2290,N_637);
and U9044 (N_9044,N_411,N_3593);
nand U9045 (N_9045,N_4625,N_518);
or U9046 (N_9046,N_323,N_3353);
and U9047 (N_9047,N_2522,N_198);
and U9048 (N_9048,N_4707,N_2650);
and U9049 (N_9049,N_3889,N_3158);
xnor U9050 (N_9050,N_1497,N_559);
xor U9051 (N_9051,N_3514,N_2918);
and U9052 (N_9052,N_846,N_3560);
or U9053 (N_9053,N_4248,N_3130);
xnor U9054 (N_9054,N_2426,N_2510);
or U9055 (N_9055,N_4932,N_2497);
nand U9056 (N_9056,N_736,N_630);
or U9057 (N_9057,N_4725,N_966);
nor U9058 (N_9058,N_1845,N_3091);
nor U9059 (N_9059,N_2304,N_3933);
nor U9060 (N_9060,N_3537,N_4617);
nor U9061 (N_9061,N_4390,N_2803);
nand U9062 (N_9062,N_2743,N_1789);
nor U9063 (N_9063,N_2214,N_1833);
nor U9064 (N_9064,N_3525,N_1836);
nor U9065 (N_9065,N_1268,N_4808);
nand U9066 (N_9066,N_1121,N_3079);
or U9067 (N_9067,N_4331,N_3371);
or U9068 (N_9068,N_787,N_1107);
nor U9069 (N_9069,N_3612,N_2119);
nor U9070 (N_9070,N_4829,N_1170);
nor U9071 (N_9071,N_4458,N_1602);
nor U9072 (N_9072,N_1625,N_1777);
nor U9073 (N_9073,N_3921,N_4394);
nand U9074 (N_9074,N_3714,N_3729);
nand U9075 (N_9075,N_2321,N_4411);
xnor U9076 (N_9076,N_3757,N_152);
nand U9077 (N_9077,N_1074,N_4602);
or U9078 (N_9078,N_2450,N_243);
nand U9079 (N_9079,N_2046,N_3031);
or U9080 (N_9080,N_4877,N_1384);
or U9081 (N_9081,N_4828,N_622);
xnor U9082 (N_9082,N_3370,N_3087);
or U9083 (N_9083,N_3261,N_786);
nor U9084 (N_9084,N_2018,N_4813);
or U9085 (N_9085,N_369,N_4020);
nor U9086 (N_9086,N_2952,N_389);
nand U9087 (N_9087,N_266,N_3085);
nand U9088 (N_9088,N_2167,N_1729);
nand U9089 (N_9089,N_3624,N_341);
or U9090 (N_9090,N_1908,N_3316);
nand U9091 (N_9091,N_4815,N_3419);
nand U9092 (N_9092,N_486,N_1313);
or U9093 (N_9093,N_611,N_4274);
nor U9094 (N_9094,N_608,N_2407);
or U9095 (N_9095,N_164,N_4941);
or U9096 (N_9096,N_579,N_794);
nand U9097 (N_9097,N_2660,N_4146);
nor U9098 (N_9098,N_4774,N_4226);
nand U9099 (N_9099,N_3393,N_1112);
xnor U9100 (N_9100,N_1833,N_3044);
and U9101 (N_9101,N_3904,N_4915);
nand U9102 (N_9102,N_2288,N_12);
or U9103 (N_9103,N_1404,N_3672);
and U9104 (N_9104,N_2237,N_616);
nand U9105 (N_9105,N_2443,N_2270);
nor U9106 (N_9106,N_2056,N_3261);
nor U9107 (N_9107,N_2922,N_206);
nor U9108 (N_9108,N_3017,N_1401);
nor U9109 (N_9109,N_1098,N_1654);
nand U9110 (N_9110,N_970,N_1714);
nor U9111 (N_9111,N_1794,N_2573);
nor U9112 (N_9112,N_1044,N_1645);
xor U9113 (N_9113,N_2893,N_4835);
nand U9114 (N_9114,N_3457,N_574);
nand U9115 (N_9115,N_981,N_154);
xor U9116 (N_9116,N_905,N_1657);
nor U9117 (N_9117,N_644,N_2971);
or U9118 (N_9118,N_2297,N_4992);
nand U9119 (N_9119,N_37,N_1361);
or U9120 (N_9120,N_144,N_2991);
or U9121 (N_9121,N_1850,N_866);
nand U9122 (N_9122,N_2842,N_158);
nand U9123 (N_9123,N_4464,N_4938);
nor U9124 (N_9124,N_2747,N_2304);
nand U9125 (N_9125,N_640,N_4949);
or U9126 (N_9126,N_2867,N_4363);
and U9127 (N_9127,N_1697,N_970);
nand U9128 (N_9128,N_547,N_4289);
and U9129 (N_9129,N_3695,N_378);
nor U9130 (N_9130,N_1022,N_1507);
or U9131 (N_9131,N_894,N_47);
nor U9132 (N_9132,N_2309,N_3837);
nor U9133 (N_9133,N_4411,N_2112);
nor U9134 (N_9134,N_1064,N_240);
or U9135 (N_9135,N_2103,N_1522);
xor U9136 (N_9136,N_1546,N_4740);
nand U9137 (N_9137,N_4346,N_1185);
or U9138 (N_9138,N_4015,N_251);
nor U9139 (N_9139,N_1294,N_3587);
nor U9140 (N_9140,N_1606,N_90);
or U9141 (N_9141,N_2729,N_1085);
and U9142 (N_9142,N_4985,N_2184);
nand U9143 (N_9143,N_3464,N_4487);
nor U9144 (N_9144,N_1932,N_1359);
and U9145 (N_9145,N_4934,N_3970);
nor U9146 (N_9146,N_2650,N_3496);
nor U9147 (N_9147,N_2656,N_3114);
nor U9148 (N_9148,N_1168,N_934);
xor U9149 (N_9149,N_2247,N_1182);
nor U9150 (N_9150,N_2017,N_4742);
and U9151 (N_9151,N_4186,N_2185);
xnor U9152 (N_9152,N_3774,N_3969);
nor U9153 (N_9153,N_2934,N_4590);
nand U9154 (N_9154,N_3010,N_2040);
nand U9155 (N_9155,N_888,N_4868);
or U9156 (N_9156,N_4108,N_3953);
and U9157 (N_9157,N_4321,N_2161);
or U9158 (N_9158,N_836,N_612);
and U9159 (N_9159,N_3807,N_1015);
nand U9160 (N_9160,N_3099,N_4081);
or U9161 (N_9161,N_682,N_651);
or U9162 (N_9162,N_3982,N_493);
and U9163 (N_9163,N_4969,N_2288);
and U9164 (N_9164,N_3617,N_4717);
and U9165 (N_9165,N_2640,N_538);
nor U9166 (N_9166,N_4496,N_2147);
xor U9167 (N_9167,N_2676,N_3186);
nor U9168 (N_9168,N_3839,N_1473);
nand U9169 (N_9169,N_2145,N_2952);
or U9170 (N_9170,N_4982,N_858);
xor U9171 (N_9171,N_1961,N_3850);
nor U9172 (N_9172,N_2909,N_2530);
and U9173 (N_9173,N_903,N_4878);
nor U9174 (N_9174,N_2291,N_617);
and U9175 (N_9175,N_4803,N_402);
nor U9176 (N_9176,N_4147,N_323);
and U9177 (N_9177,N_3741,N_2726);
or U9178 (N_9178,N_3199,N_559);
and U9179 (N_9179,N_1346,N_498);
nand U9180 (N_9180,N_2497,N_2494);
and U9181 (N_9181,N_4101,N_1898);
nor U9182 (N_9182,N_4678,N_2545);
nand U9183 (N_9183,N_391,N_1535);
xnor U9184 (N_9184,N_3339,N_2235);
and U9185 (N_9185,N_216,N_3711);
nor U9186 (N_9186,N_143,N_2858);
xnor U9187 (N_9187,N_1146,N_4813);
nand U9188 (N_9188,N_2821,N_1487);
nor U9189 (N_9189,N_324,N_3780);
xor U9190 (N_9190,N_4554,N_4567);
nand U9191 (N_9191,N_2195,N_4462);
nand U9192 (N_9192,N_3646,N_690);
xor U9193 (N_9193,N_1324,N_820);
and U9194 (N_9194,N_1012,N_2223);
and U9195 (N_9195,N_2089,N_2904);
or U9196 (N_9196,N_962,N_2702);
nand U9197 (N_9197,N_3625,N_3829);
or U9198 (N_9198,N_1797,N_447);
nand U9199 (N_9199,N_2424,N_930);
xor U9200 (N_9200,N_1331,N_4503);
or U9201 (N_9201,N_3369,N_2544);
and U9202 (N_9202,N_4349,N_4882);
or U9203 (N_9203,N_3580,N_3641);
or U9204 (N_9204,N_3770,N_777);
nand U9205 (N_9205,N_3976,N_323);
nor U9206 (N_9206,N_2762,N_4211);
and U9207 (N_9207,N_2982,N_2637);
or U9208 (N_9208,N_2020,N_733);
and U9209 (N_9209,N_1382,N_3494);
nand U9210 (N_9210,N_1351,N_2500);
and U9211 (N_9211,N_2993,N_699);
nand U9212 (N_9212,N_2979,N_2001);
or U9213 (N_9213,N_24,N_1379);
and U9214 (N_9214,N_1194,N_1365);
and U9215 (N_9215,N_3140,N_4942);
nor U9216 (N_9216,N_3770,N_3154);
nor U9217 (N_9217,N_3094,N_2671);
and U9218 (N_9218,N_4383,N_1123);
and U9219 (N_9219,N_3875,N_4743);
nand U9220 (N_9220,N_3630,N_1266);
xor U9221 (N_9221,N_285,N_3111);
and U9222 (N_9222,N_1596,N_2210);
or U9223 (N_9223,N_3776,N_4321);
or U9224 (N_9224,N_3195,N_4495);
and U9225 (N_9225,N_3303,N_1500);
or U9226 (N_9226,N_2119,N_2256);
nand U9227 (N_9227,N_3826,N_2056);
nand U9228 (N_9228,N_314,N_4118);
nor U9229 (N_9229,N_351,N_1609);
nor U9230 (N_9230,N_4333,N_4173);
nor U9231 (N_9231,N_2790,N_4750);
and U9232 (N_9232,N_1739,N_264);
and U9233 (N_9233,N_2637,N_3055);
nand U9234 (N_9234,N_559,N_3493);
xor U9235 (N_9235,N_2851,N_1658);
nand U9236 (N_9236,N_2845,N_2668);
nand U9237 (N_9237,N_960,N_839);
or U9238 (N_9238,N_3744,N_4038);
or U9239 (N_9239,N_958,N_4887);
or U9240 (N_9240,N_1669,N_1394);
nor U9241 (N_9241,N_3054,N_781);
or U9242 (N_9242,N_236,N_3604);
or U9243 (N_9243,N_758,N_3290);
nor U9244 (N_9244,N_2676,N_4531);
or U9245 (N_9245,N_1682,N_1796);
or U9246 (N_9246,N_552,N_640);
or U9247 (N_9247,N_4098,N_4256);
nand U9248 (N_9248,N_4424,N_2678);
nand U9249 (N_9249,N_1558,N_42);
nor U9250 (N_9250,N_1574,N_695);
or U9251 (N_9251,N_3952,N_1919);
and U9252 (N_9252,N_4572,N_3150);
and U9253 (N_9253,N_3465,N_3832);
and U9254 (N_9254,N_3517,N_1310);
nand U9255 (N_9255,N_1305,N_987);
nor U9256 (N_9256,N_4536,N_1353);
or U9257 (N_9257,N_2229,N_2690);
and U9258 (N_9258,N_1988,N_4069);
nand U9259 (N_9259,N_4850,N_4976);
nand U9260 (N_9260,N_1879,N_4097);
and U9261 (N_9261,N_813,N_4880);
or U9262 (N_9262,N_597,N_3565);
nand U9263 (N_9263,N_610,N_3538);
xor U9264 (N_9264,N_2617,N_1613);
and U9265 (N_9265,N_942,N_3431);
nand U9266 (N_9266,N_840,N_1806);
or U9267 (N_9267,N_4151,N_3859);
nand U9268 (N_9268,N_169,N_1033);
and U9269 (N_9269,N_2565,N_2504);
nor U9270 (N_9270,N_3376,N_4004);
xor U9271 (N_9271,N_1221,N_2968);
and U9272 (N_9272,N_2341,N_4959);
and U9273 (N_9273,N_3862,N_1345);
nand U9274 (N_9274,N_1385,N_3484);
and U9275 (N_9275,N_1535,N_598);
and U9276 (N_9276,N_226,N_4108);
nand U9277 (N_9277,N_2326,N_4805);
nor U9278 (N_9278,N_1308,N_3427);
nor U9279 (N_9279,N_883,N_2693);
or U9280 (N_9280,N_666,N_541);
nor U9281 (N_9281,N_2189,N_2423);
and U9282 (N_9282,N_3067,N_775);
and U9283 (N_9283,N_1684,N_15);
or U9284 (N_9284,N_3700,N_4843);
or U9285 (N_9285,N_1214,N_401);
nor U9286 (N_9286,N_746,N_1125);
nand U9287 (N_9287,N_944,N_3759);
nor U9288 (N_9288,N_1027,N_721);
and U9289 (N_9289,N_1197,N_4556);
nand U9290 (N_9290,N_1522,N_1058);
xor U9291 (N_9291,N_4367,N_4510);
or U9292 (N_9292,N_1163,N_2116);
xnor U9293 (N_9293,N_3072,N_3638);
and U9294 (N_9294,N_1387,N_165);
and U9295 (N_9295,N_4494,N_2740);
or U9296 (N_9296,N_3349,N_669);
nand U9297 (N_9297,N_2081,N_769);
and U9298 (N_9298,N_1286,N_3555);
and U9299 (N_9299,N_740,N_1729);
and U9300 (N_9300,N_2768,N_3680);
and U9301 (N_9301,N_2515,N_2287);
or U9302 (N_9302,N_197,N_214);
nand U9303 (N_9303,N_2837,N_728);
and U9304 (N_9304,N_2660,N_1008);
and U9305 (N_9305,N_1222,N_1766);
nand U9306 (N_9306,N_3806,N_3970);
nor U9307 (N_9307,N_224,N_3884);
and U9308 (N_9308,N_1784,N_4260);
and U9309 (N_9309,N_4553,N_2941);
and U9310 (N_9310,N_890,N_3586);
and U9311 (N_9311,N_2331,N_2544);
and U9312 (N_9312,N_1265,N_2528);
nor U9313 (N_9313,N_3363,N_3922);
nor U9314 (N_9314,N_2116,N_676);
and U9315 (N_9315,N_4376,N_312);
nor U9316 (N_9316,N_558,N_666);
and U9317 (N_9317,N_204,N_577);
nor U9318 (N_9318,N_714,N_259);
nor U9319 (N_9319,N_2822,N_1989);
nand U9320 (N_9320,N_729,N_769);
nor U9321 (N_9321,N_4766,N_629);
nand U9322 (N_9322,N_1963,N_1205);
and U9323 (N_9323,N_951,N_4914);
and U9324 (N_9324,N_1864,N_1344);
and U9325 (N_9325,N_907,N_798);
or U9326 (N_9326,N_3781,N_3824);
or U9327 (N_9327,N_4562,N_1066);
xnor U9328 (N_9328,N_2018,N_3864);
and U9329 (N_9329,N_2749,N_2350);
nand U9330 (N_9330,N_2939,N_1990);
nor U9331 (N_9331,N_3462,N_1115);
or U9332 (N_9332,N_4971,N_2864);
or U9333 (N_9333,N_4643,N_4768);
nor U9334 (N_9334,N_3116,N_2344);
nand U9335 (N_9335,N_510,N_1057);
nor U9336 (N_9336,N_2786,N_2699);
xor U9337 (N_9337,N_24,N_632);
or U9338 (N_9338,N_2112,N_4722);
xor U9339 (N_9339,N_2361,N_139);
and U9340 (N_9340,N_4236,N_4427);
and U9341 (N_9341,N_2577,N_1300);
nand U9342 (N_9342,N_4880,N_4520);
nor U9343 (N_9343,N_853,N_1864);
or U9344 (N_9344,N_4128,N_2593);
and U9345 (N_9345,N_578,N_493);
and U9346 (N_9346,N_1570,N_4763);
or U9347 (N_9347,N_1817,N_4982);
nor U9348 (N_9348,N_2849,N_2079);
and U9349 (N_9349,N_1813,N_4706);
or U9350 (N_9350,N_1365,N_2928);
and U9351 (N_9351,N_3269,N_2386);
nor U9352 (N_9352,N_1266,N_3029);
and U9353 (N_9353,N_4173,N_1607);
or U9354 (N_9354,N_1474,N_3742);
or U9355 (N_9355,N_789,N_2509);
and U9356 (N_9356,N_3967,N_1714);
nand U9357 (N_9357,N_1565,N_2308);
nand U9358 (N_9358,N_1282,N_557);
nor U9359 (N_9359,N_1015,N_964);
xnor U9360 (N_9360,N_1260,N_1450);
or U9361 (N_9361,N_1960,N_4448);
nand U9362 (N_9362,N_67,N_1267);
nand U9363 (N_9363,N_1462,N_1747);
or U9364 (N_9364,N_3346,N_2623);
or U9365 (N_9365,N_3949,N_2750);
and U9366 (N_9366,N_4473,N_3477);
and U9367 (N_9367,N_184,N_604);
nor U9368 (N_9368,N_4910,N_1269);
or U9369 (N_9369,N_3922,N_2296);
nor U9370 (N_9370,N_1330,N_873);
nor U9371 (N_9371,N_3741,N_2514);
nand U9372 (N_9372,N_3728,N_4508);
or U9373 (N_9373,N_4984,N_467);
nand U9374 (N_9374,N_1441,N_4550);
or U9375 (N_9375,N_1990,N_4361);
nand U9376 (N_9376,N_1443,N_4885);
nand U9377 (N_9377,N_2378,N_4464);
nand U9378 (N_9378,N_1005,N_2271);
nor U9379 (N_9379,N_4753,N_2059);
and U9380 (N_9380,N_676,N_4284);
or U9381 (N_9381,N_2650,N_2632);
nand U9382 (N_9382,N_438,N_3849);
or U9383 (N_9383,N_763,N_4526);
and U9384 (N_9384,N_2116,N_465);
and U9385 (N_9385,N_3646,N_116);
nor U9386 (N_9386,N_421,N_628);
or U9387 (N_9387,N_689,N_2078);
nor U9388 (N_9388,N_2763,N_4561);
nor U9389 (N_9389,N_2899,N_4027);
nor U9390 (N_9390,N_2615,N_1295);
or U9391 (N_9391,N_2467,N_2756);
nand U9392 (N_9392,N_4826,N_2988);
and U9393 (N_9393,N_3305,N_554);
or U9394 (N_9394,N_2914,N_396);
nand U9395 (N_9395,N_506,N_2391);
nor U9396 (N_9396,N_386,N_4205);
nand U9397 (N_9397,N_373,N_719);
and U9398 (N_9398,N_135,N_1036);
nor U9399 (N_9399,N_4497,N_4199);
nand U9400 (N_9400,N_967,N_2624);
xnor U9401 (N_9401,N_896,N_3425);
nor U9402 (N_9402,N_2313,N_3360);
nor U9403 (N_9403,N_149,N_854);
and U9404 (N_9404,N_3879,N_4981);
nor U9405 (N_9405,N_1342,N_1004);
and U9406 (N_9406,N_2627,N_1498);
and U9407 (N_9407,N_3840,N_218);
nand U9408 (N_9408,N_4827,N_3436);
nand U9409 (N_9409,N_619,N_1388);
nor U9410 (N_9410,N_3335,N_2285);
xor U9411 (N_9411,N_4730,N_819);
or U9412 (N_9412,N_2851,N_2232);
and U9413 (N_9413,N_1862,N_1873);
nor U9414 (N_9414,N_4729,N_19);
nand U9415 (N_9415,N_3429,N_704);
or U9416 (N_9416,N_1526,N_3133);
nor U9417 (N_9417,N_2546,N_294);
and U9418 (N_9418,N_1625,N_4439);
xor U9419 (N_9419,N_2277,N_1911);
nor U9420 (N_9420,N_4469,N_2878);
nor U9421 (N_9421,N_2485,N_4174);
and U9422 (N_9422,N_3975,N_4064);
or U9423 (N_9423,N_3639,N_3274);
nor U9424 (N_9424,N_2974,N_3712);
or U9425 (N_9425,N_3503,N_4321);
nand U9426 (N_9426,N_1120,N_4262);
or U9427 (N_9427,N_906,N_3637);
xnor U9428 (N_9428,N_4370,N_4683);
or U9429 (N_9429,N_4988,N_2005);
nand U9430 (N_9430,N_4360,N_4001);
nor U9431 (N_9431,N_1133,N_2397);
nor U9432 (N_9432,N_3582,N_2833);
and U9433 (N_9433,N_1067,N_4861);
nor U9434 (N_9434,N_3939,N_3254);
nand U9435 (N_9435,N_2112,N_1263);
nor U9436 (N_9436,N_3014,N_3125);
nor U9437 (N_9437,N_397,N_1464);
nand U9438 (N_9438,N_3771,N_143);
nand U9439 (N_9439,N_3524,N_3301);
and U9440 (N_9440,N_2376,N_3469);
or U9441 (N_9441,N_598,N_555);
and U9442 (N_9442,N_4987,N_3712);
xnor U9443 (N_9443,N_2135,N_3549);
and U9444 (N_9444,N_2613,N_2360);
nand U9445 (N_9445,N_4645,N_1760);
nor U9446 (N_9446,N_1719,N_1972);
nand U9447 (N_9447,N_4628,N_1356);
xor U9448 (N_9448,N_4327,N_4655);
and U9449 (N_9449,N_2561,N_4412);
and U9450 (N_9450,N_2025,N_3143);
nor U9451 (N_9451,N_2201,N_35);
and U9452 (N_9452,N_3583,N_2654);
or U9453 (N_9453,N_4585,N_2469);
xor U9454 (N_9454,N_3595,N_766);
xor U9455 (N_9455,N_2672,N_2046);
nor U9456 (N_9456,N_3575,N_3416);
and U9457 (N_9457,N_2236,N_326);
nand U9458 (N_9458,N_4132,N_1228);
or U9459 (N_9459,N_2563,N_1916);
and U9460 (N_9460,N_1042,N_461);
nor U9461 (N_9461,N_324,N_3269);
and U9462 (N_9462,N_2849,N_4095);
nand U9463 (N_9463,N_1506,N_4286);
nor U9464 (N_9464,N_670,N_1248);
xnor U9465 (N_9465,N_353,N_2315);
or U9466 (N_9466,N_1504,N_1535);
or U9467 (N_9467,N_587,N_3290);
or U9468 (N_9468,N_477,N_1027);
nor U9469 (N_9469,N_3567,N_2893);
or U9470 (N_9470,N_3744,N_357);
or U9471 (N_9471,N_537,N_3631);
and U9472 (N_9472,N_3763,N_4434);
xor U9473 (N_9473,N_3898,N_2198);
xnor U9474 (N_9474,N_1707,N_3111);
and U9475 (N_9475,N_1930,N_973);
or U9476 (N_9476,N_3630,N_1273);
or U9477 (N_9477,N_2573,N_221);
and U9478 (N_9478,N_3393,N_4620);
and U9479 (N_9479,N_3366,N_1824);
and U9480 (N_9480,N_3248,N_2522);
xnor U9481 (N_9481,N_344,N_3407);
nand U9482 (N_9482,N_48,N_1390);
nor U9483 (N_9483,N_4413,N_4500);
and U9484 (N_9484,N_1281,N_388);
or U9485 (N_9485,N_1421,N_91);
or U9486 (N_9486,N_3755,N_420);
or U9487 (N_9487,N_1080,N_2446);
xnor U9488 (N_9488,N_4088,N_2349);
nand U9489 (N_9489,N_3914,N_4178);
nor U9490 (N_9490,N_2148,N_1613);
nor U9491 (N_9491,N_1263,N_2313);
or U9492 (N_9492,N_1683,N_1520);
and U9493 (N_9493,N_372,N_3595);
or U9494 (N_9494,N_3304,N_4958);
and U9495 (N_9495,N_191,N_746);
xor U9496 (N_9496,N_1590,N_1677);
or U9497 (N_9497,N_4347,N_3232);
xor U9498 (N_9498,N_3652,N_473);
nand U9499 (N_9499,N_2441,N_1402);
and U9500 (N_9500,N_2067,N_291);
or U9501 (N_9501,N_1156,N_4527);
or U9502 (N_9502,N_4346,N_1515);
nor U9503 (N_9503,N_3873,N_2294);
xnor U9504 (N_9504,N_2069,N_1885);
nor U9505 (N_9505,N_1450,N_3613);
or U9506 (N_9506,N_65,N_1007);
and U9507 (N_9507,N_2165,N_1297);
nand U9508 (N_9508,N_76,N_455);
and U9509 (N_9509,N_4510,N_3885);
nand U9510 (N_9510,N_4085,N_2031);
nor U9511 (N_9511,N_4438,N_920);
and U9512 (N_9512,N_901,N_3495);
nor U9513 (N_9513,N_3005,N_3759);
nand U9514 (N_9514,N_843,N_3237);
nand U9515 (N_9515,N_2283,N_22);
xnor U9516 (N_9516,N_3432,N_2284);
xor U9517 (N_9517,N_1101,N_4372);
xor U9518 (N_9518,N_3332,N_3260);
nor U9519 (N_9519,N_653,N_1906);
or U9520 (N_9520,N_4730,N_1447);
xnor U9521 (N_9521,N_1394,N_3293);
nor U9522 (N_9522,N_2962,N_2530);
nor U9523 (N_9523,N_1973,N_3970);
nor U9524 (N_9524,N_470,N_4285);
nand U9525 (N_9525,N_4947,N_1262);
nor U9526 (N_9526,N_2444,N_3252);
nor U9527 (N_9527,N_4646,N_1073);
nand U9528 (N_9528,N_931,N_4036);
nand U9529 (N_9529,N_533,N_3344);
or U9530 (N_9530,N_4099,N_3129);
nand U9531 (N_9531,N_2745,N_2447);
nor U9532 (N_9532,N_2032,N_2203);
or U9533 (N_9533,N_4865,N_57);
nand U9534 (N_9534,N_1461,N_4438);
and U9535 (N_9535,N_146,N_4963);
and U9536 (N_9536,N_3628,N_1055);
or U9537 (N_9537,N_197,N_2452);
and U9538 (N_9538,N_2909,N_3053);
nor U9539 (N_9539,N_2565,N_2752);
nor U9540 (N_9540,N_3740,N_2574);
or U9541 (N_9541,N_3696,N_1175);
nand U9542 (N_9542,N_400,N_2443);
nand U9543 (N_9543,N_4716,N_340);
or U9544 (N_9544,N_1892,N_541);
and U9545 (N_9545,N_1753,N_3959);
or U9546 (N_9546,N_3684,N_1547);
or U9547 (N_9547,N_2219,N_330);
nand U9548 (N_9548,N_4333,N_2839);
or U9549 (N_9549,N_2284,N_3404);
or U9550 (N_9550,N_937,N_1036);
and U9551 (N_9551,N_0,N_692);
nand U9552 (N_9552,N_2946,N_3312);
and U9553 (N_9553,N_4231,N_202);
nor U9554 (N_9554,N_2994,N_2032);
or U9555 (N_9555,N_1052,N_2524);
or U9556 (N_9556,N_3448,N_2532);
and U9557 (N_9557,N_283,N_3664);
or U9558 (N_9558,N_1603,N_843);
nand U9559 (N_9559,N_890,N_428);
or U9560 (N_9560,N_4056,N_988);
nand U9561 (N_9561,N_1594,N_2469);
nand U9562 (N_9562,N_2914,N_1427);
nor U9563 (N_9563,N_3783,N_4543);
nand U9564 (N_9564,N_2016,N_700);
and U9565 (N_9565,N_2429,N_2494);
and U9566 (N_9566,N_1178,N_3596);
nor U9567 (N_9567,N_3182,N_278);
or U9568 (N_9568,N_220,N_57);
xor U9569 (N_9569,N_1293,N_1071);
nor U9570 (N_9570,N_3694,N_2186);
nor U9571 (N_9571,N_3408,N_3418);
nor U9572 (N_9572,N_1696,N_2308);
or U9573 (N_9573,N_3278,N_4076);
nor U9574 (N_9574,N_3700,N_3282);
and U9575 (N_9575,N_3985,N_4283);
or U9576 (N_9576,N_2441,N_4782);
nand U9577 (N_9577,N_965,N_2078);
nor U9578 (N_9578,N_3052,N_4081);
nor U9579 (N_9579,N_2832,N_734);
nor U9580 (N_9580,N_2274,N_1668);
nand U9581 (N_9581,N_3842,N_2643);
nor U9582 (N_9582,N_3620,N_197);
and U9583 (N_9583,N_4199,N_2919);
xnor U9584 (N_9584,N_1064,N_3914);
nor U9585 (N_9585,N_2454,N_4108);
and U9586 (N_9586,N_2778,N_3124);
and U9587 (N_9587,N_1945,N_818);
xnor U9588 (N_9588,N_3818,N_1981);
or U9589 (N_9589,N_3158,N_235);
nand U9590 (N_9590,N_1598,N_2991);
xnor U9591 (N_9591,N_1130,N_1580);
or U9592 (N_9592,N_4749,N_3256);
nand U9593 (N_9593,N_4893,N_4991);
nand U9594 (N_9594,N_3909,N_3882);
nor U9595 (N_9595,N_732,N_2719);
nor U9596 (N_9596,N_522,N_2273);
nand U9597 (N_9597,N_1480,N_3125);
nor U9598 (N_9598,N_2198,N_1378);
or U9599 (N_9599,N_1348,N_2874);
nor U9600 (N_9600,N_3905,N_715);
and U9601 (N_9601,N_42,N_4148);
nand U9602 (N_9602,N_437,N_1015);
nand U9603 (N_9603,N_3896,N_311);
nand U9604 (N_9604,N_1708,N_715);
or U9605 (N_9605,N_3935,N_3851);
nand U9606 (N_9606,N_329,N_1129);
and U9607 (N_9607,N_1300,N_864);
and U9608 (N_9608,N_217,N_1075);
nand U9609 (N_9609,N_4974,N_544);
nand U9610 (N_9610,N_4688,N_322);
or U9611 (N_9611,N_2432,N_4368);
nand U9612 (N_9612,N_2585,N_151);
and U9613 (N_9613,N_3823,N_1752);
nor U9614 (N_9614,N_1200,N_4843);
nor U9615 (N_9615,N_2561,N_4271);
nand U9616 (N_9616,N_2369,N_1876);
nand U9617 (N_9617,N_3539,N_3151);
and U9618 (N_9618,N_3142,N_4422);
nand U9619 (N_9619,N_4995,N_1269);
nor U9620 (N_9620,N_2065,N_1183);
nand U9621 (N_9621,N_4973,N_3162);
xnor U9622 (N_9622,N_4829,N_1543);
or U9623 (N_9623,N_2514,N_1065);
nand U9624 (N_9624,N_708,N_3771);
and U9625 (N_9625,N_1125,N_1234);
nor U9626 (N_9626,N_4219,N_2734);
or U9627 (N_9627,N_1350,N_2675);
nand U9628 (N_9628,N_623,N_2063);
nor U9629 (N_9629,N_3326,N_577);
or U9630 (N_9630,N_1414,N_4703);
nand U9631 (N_9631,N_4382,N_3669);
or U9632 (N_9632,N_2810,N_3777);
or U9633 (N_9633,N_3489,N_3840);
nand U9634 (N_9634,N_886,N_745);
nand U9635 (N_9635,N_3886,N_3426);
and U9636 (N_9636,N_4360,N_4351);
or U9637 (N_9637,N_483,N_750);
and U9638 (N_9638,N_1627,N_4568);
nand U9639 (N_9639,N_4267,N_163);
xnor U9640 (N_9640,N_775,N_2269);
or U9641 (N_9641,N_3008,N_4929);
xnor U9642 (N_9642,N_649,N_3777);
nand U9643 (N_9643,N_1097,N_785);
nor U9644 (N_9644,N_3225,N_2044);
or U9645 (N_9645,N_520,N_3838);
or U9646 (N_9646,N_3106,N_1578);
and U9647 (N_9647,N_4194,N_3216);
and U9648 (N_9648,N_4835,N_207);
nand U9649 (N_9649,N_2587,N_3250);
nand U9650 (N_9650,N_1344,N_3691);
and U9651 (N_9651,N_4129,N_1699);
nor U9652 (N_9652,N_579,N_58);
xor U9653 (N_9653,N_1067,N_4785);
nand U9654 (N_9654,N_1991,N_897);
or U9655 (N_9655,N_3856,N_4416);
nor U9656 (N_9656,N_785,N_200);
or U9657 (N_9657,N_75,N_3030);
nand U9658 (N_9658,N_4804,N_4309);
and U9659 (N_9659,N_1172,N_84);
nand U9660 (N_9660,N_2335,N_3804);
nor U9661 (N_9661,N_3027,N_1642);
and U9662 (N_9662,N_1894,N_2111);
nor U9663 (N_9663,N_863,N_53);
or U9664 (N_9664,N_2068,N_992);
nand U9665 (N_9665,N_352,N_3204);
and U9666 (N_9666,N_3565,N_2092);
or U9667 (N_9667,N_2920,N_3770);
and U9668 (N_9668,N_4240,N_2706);
nor U9669 (N_9669,N_3254,N_4277);
and U9670 (N_9670,N_2135,N_4670);
nand U9671 (N_9671,N_248,N_1763);
xor U9672 (N_9672,N_4330,N_312);
or U9673 (N_9673,N_1746,N_594);
nand U9674 (N_9674,N_3176,N_4951);
or U9675 (N_9675,N_735,N_1882);
nor U9676 (N_9676,N_3345,N_671);
nand U9677 (N_9677,N_612,N_1267);
nand U9678 (N_9678,N_3919,N_1909);
or U9679 (N_9679,N_2847,N_1327);
and U9680 (N_9680,N_1026,N_167);
and U9681 (N_9681,N_4548,N_4829);
and U9682 (N_9682,N_1794,N_1316);
or U9683 (N_9683,N_767,N_1357);
xnor U9684 (N_9684,N_2462,N_3063);
xnor U9685 (N_9685,N_1826,N_3768);
xor U9686 (N_9686,N_2052,N_2542);
xor U9687 (N_9687,N_1740,N_4870);
nand U9688 (N_9688,N_3704,N_1351);
and U9689 (N_9689,N_3452,N_1609);
and U9690 (N_9690,N_3219,N_1792);
nor U9691 (N_9691,N_1733,N_3612);
nand U9692 (N_9692,N_4430,N_1351);
or U9693 (N_9693,N_2092,N_69);
or U9694 (N_9694,N_2476,N_1023);
nor U9695 (N_9695,N_3482,N_1275);
or U9696 (N_9696,N_3040,N_4986);
xor U9697 (N_9697,N_2598,N_517);
nand U9698 (N_9698,N_1575,N_4140);
xnor U9699 (N_9699,N_2799,N_3454);
xor U9700 (N_9700,N_4326,N_1022);
nand U9701 (N_9701,N_150,N_742);
nor U9702 (N_9702,N_1967,N_4874);
nand U9703 (N_9703,N_3318,N_632);
nand U9704 (N_9704,N_4630,N_1638);
nand U9705 (N_9705,N_237,N_3771);
nor U9706 (N_9706,N_4282,N_1470);
xnor U9707 (N_9707,N_620,N_4608);
nand U9708 (N_9708,N_2497,N_1200);
and U9709 (N_9709,N_1843,N_3159);
and U9710 (N_9710,N_1335,N_4274);
nor U9711 (N_9711,N_2778,N_3537);
nor U9712 (N_9712,N_699,N_1071);
or U9713 (N_9713,N_1467,N_2790);
nand U9714 (N_9714,N_1531,N_1917);
xnor U9715 (N_9715,N_4798,N_1082);
nor U9716 (N_9716,N_3775,N_4261);
and U9717 (N_9717,N_1653,N_730);
nor U9718 (N_9718,N_2152,N_4518);
nor U9719 (N_9719,N_565,N_105);
and U9720 (N_9720,N_4445,N_2921);
nor U9721 (N_9721,N_1683,N_4268);
nor U9722 (N_9722,N_3542,N_4620);
and U9723 (N_9723,N_943,N_1823);
nor U9724 (N_9724,N_4169,N_2939);
xor U9725 (N_9725,N_2119,N_4504);
nand U9726 (N_9726,N_2422,N_120);
and U9727 (N_9727,N_2146,N_4638);
nand U9728 (N_9728,N_3376,N_157);
or U9729 (N_9729,N_3491,N_4660);
nor U9730 (N_9730,N_3189,N_3631);
nand U9731 (N_9731,N_1365,N_4322);
nand U9732 (N_9732,N_2186,N_1936);
nand U9733 (N_9733,N_981,N_2363);
nand U9734 (N_9734,N_2960,N_1171);
or U9735 (N_9735,N_2453,N_2083);
nor U9736 (N_9736,N_2432,N_3561);
nand U9737 (N_9737,N_1643,N_1843);
or U9738 (N_9738,N_817,N_1873);
xor U9739 (N_9739,N_4285,N_1254);
or U9740 (N_9740,N_3387,N_4052);
xnor U9741 (N_9741,N_677,N_1132);
or U9742 (N_9742,N_3168,N_2279);
or U9743 (N_9743,N_3569,N_4368);
and U9744 (N_9744,N_2297,N_3333);
and U9745 (N_9745,N_4930,N_682);
nand U9746 (N_9746,N_1600,N_727);
or U9747 (N_9747,N_3658,N_3115);
nand U9748 (N_9748,N_2147,N_2654);
or U9749 (N_9749,N_361,N_1770);
nand U9750 (N_9750,N_1519,N_1860);
nand U9751 (N_9751,N_3369,N_560);
nor U9752 (N_9752,N_1532,N_504);
nor U9753 (N_9753,N_4234,N_809);
or U9754 (N_9754,N_19,N_277);
nor U9755 (N_9755,N_3507,N_201);
and U9756 (N_9756,N_4648,N_3652);
and U9757 (N_9757,N_1156,N_2704);
nor U9758 (N_9758,N_4766,N_1297);
xnor U9759 (N_9759,N_1371,N_3762);
and U9760 (N_9760,N_349,N_1267);
nor U9761 (N_9761,N_3327,N_4751);
or U9762 (N_9762,N_387,N_1588);
or U9763 (N_9763,N_954,N_4948);
or U9764 (N_9764,N_1320,N_2688);
nor U9765 (N_9765,N_4990,N_2646);
nand U9766 (N_9766,N_2037,N_3294);
nor U9767 (N_9767,N_1762,N_4710);
nand U9768 (N_9768,N_2131,N_4937);
nand U9769 (N_9769,N_151,N_297);
nor U9770 (N_9770,N_153,N_1070);
or U9771 (N_9771,N_4436,N_2136);
and U9772 (N_9772,N_2235,N_4951);
nand U9773 (N_9773,N_2350,N_4979);
and U9774 (N_9774,N_3265,N_4721);
or U9775 (N_9775,N_2709,N_3660);
and U9776 (N_9776,N_3178,N_1801);
nor U9777 (N_9777,N_1284,N_1560);
and U9778 (N_9778,N_1059,N_62);
or U9779 (N_9779,N_554,N_1642);
nor U9780 (N_9780,N_438,N_248);
nand U9781 (N_9781,N_4265,N_2969);
nand U9782 (N_9782,N_2255,N_2353);
nor U9783 (N_9783,N_4931,N_2079);
nand U9784 (N_9784,N_3345,N_1064);
or U9785 (N_9785,N_3999,N_50);
nor U9786 (N_9786,N_3843,N_4501);
nand U9787 (N_9787,N_4191,N_3948);
and U9788 (N_9788,N_1571,N_1012);
or U9789 (N_9789,N_631,N_1510);
and U9790 (N_9790,N_3815,N_3540);
nand U9791 (N_9791,N_3915,N_4247);
xnor U9792 (N_9792,N_3184,N_4119);
and U9793 (N_9793,N_3869,N_3403);
or U9794 (N_9794,N_3049,N_1608);
nor U9795 (N_9795,N_270,N_453);
xnor U9796 (N_9796,N_4450,N_4138);
and U9797 (N_9797,N_1911,N_3154);
or U9798 (N_9798,N_2921,N_1405);
and U9799 (N_9799,N_439,N_3119);
and U9800 (N_9800,N_2373,N_1640);
or U9801 (N_9801,N_516,N_3604);
nor U9802 (N_9802,N_1205,N_2854);
nand U9803 (N_9803,N_4166,N_4173);
nand U9804 (N_9804,N_2661,N_1793);
nor U9805 (N_9805,N_298,N_4203);
and U9806 (N_9806,N_819,N_1286);
and U9807 (N_9807,N_2012,N_557);
or U9808 (N_9808,N_3103,N_2592);
xor U9809 (N_9809,N_3051,N_263);
or U9810 (N_9810,N_4453,N_688);
or U9811 (N_9811,N_1594,N_2370);
nand U9812 (N_9812,N_771,N_4906);
and U9813 (N_9813,N_4016,N_2458);
nor U9814 (N_9814,N_4175,N_175);
nand U9815 (N_9815,N_2262,N_3803);
nand U9816 (N_9816,N_2475,N_279);
nand U9817 (N_9817,N_1961,N_3549);
nor U9818 (N_9818,N_3910,N_1607);
nor U9819 (N_9819,N_3588,N_1017);
xnor U9820 (N_9820,N_4045,N_2412);
xnor U9821 (N_9821,N_2513,N_3506);
xnor U9822 (N_9822,N_4905,N_2015);
xor U9823 (N_9823,N_1160,N_1791);
or U9824 (N_9824,N_4717,N_759);
xor U9825 (N_9825,N_1433,N_2016);
or U9826 (N_9826,N_2081,N_4290);
nand U9827 (N_9827,N_3396,N_3426);
nor U9828 (N_9828,N_2419,N_394);
and U9829 (N_9829,N_4421,N_1191);
and U9830 (N_9830,N_4473,N_3209);
xnor U9831 (N_9831,N_3856,N_3932);
and U9832 (N_9832,N_12,N_1628);
or U9833 (N_9833,N_4648,N_1956);
nand U9834 (N_9834,N_4597,N_3929);
nand U9835 (N_9835,N_4908,N_1622);
nor U9836 (N_9836,N_4579,N_3364);
xor U9837 (N_9837,N_4164,N_4569);
nand U9838 (N_9838,N_2895,N_2176);
nand U9839 (N_9839,N_4372,N_882);
nor U9840 (N_9840,N_729,N_3566);
nor U9841 (N_9841,N_904,N_118);
or U9842 (N_9842,N_864,N_1362);
or U9843 (N_9843,N_2095,N_4365);
nand U9844 (N_9844,N_2125,N_807);
xor U9845 (N_9845,N_1909,N_3888);
and U9846 (N_9846,N_2919,N_1979);
and U9847 (N_9847,N_455,N_3418);
nand U9848 (N_9848,N_2538,N_4643);
nand U9849 (N_9849,N_851,N_4587);
nand U9850 (N_9850,N_4415,N_247);
and U9851 (N_9851,N_4327,N_1396);
or U9852 (N_9852,N_4337,N_3745);
or U9853 (N_9853,N_977,N_3248);
nand U9854 (N_9854,N_2604,N_2121);
and U9855 (N_9855,N_2647,N_4512);
and U9856 (N_9856,N_1900,N_3899);
nand U9857 (N_9857,N_1574,N_4856);
nor U9858 (N_9858,N_1546,N_3283);
nand U9859 (N_9859,N_3859,N_1316);
and U9860 (N_9860,N_4459,N_4344);
nor U9861 (N_9861,N_3816,N_1976);
or U9862 (N_9862,N_3585,N_2837);
or U9863 (N_9863,N_1212,N_4571);
and U9864 (N_9864,N_4685,N_3780);
and U9865 (N_9865,N_3774,N_4203);
nor U9866 (N_9866,N_2320,N_187);
and U9867 (N_9867,N_2399,N_1131);
nor U9868 (N_9868,N_2044,N_3234);
or U9869 (N_9869,N_4264,N_2532);
and U9870 (N_9870,N_2650,N_2382);
nor U9871 (N_9871,N_48,N_3735);
and U9872 (N_9872,N_1207,N_1032);
and U9873 (N_9873,N_1202,N_2984);
and U9874 (N_9874,N_89,N_4528);
nand U9875 (N_9875,N_4331,N_3567);
nor U9876 (N_9876,N_202,N_1709);
or U9877 (N_9877,N_3015,N_3034);
xnor U9878 (N_9878,N_1969,N_1335);
nand U9879 (N_9879,N_4977,N_4732);
or U9880 (N_9880,N_2384,N_1726);
nand U9881 (N_9881,N_3656,N_3266);
nor U9882 (N_9882,N_4835,N_3897);
or U9883 (N_9883,N_4586,N_3018);
and U9884 (N_9884,N_288,N_1748);
xor U9885 (N_9885,N_3445,N_198);
xor U9886 (N_9886,N_2557,N_3815);
and U9887 (N_9887,N_1918,N_609);
nor U9888 (N_9888,N_4153,N_3537);
nand U9889 (N_9889,N_1154,N_2718);
or U9890 (N_9890,N_2274,N_737);
and U9891 (N_9891,N_3402,N_1755);
nor U9892 (N_9892,N_3350,N_3322);
nor U9893 (N_9893,N_3236,N_2490);
xor U9894 (N_9894,N_4493,N_3090);
nand U9895 (N_9895,N_4030,N_1009);
and U9896 (N_9896,N_868,N_3031);
nor U9897 (N_9897,N_2227,N_1722);
and U9898 (N_9898,N_919,N_935);
nor U9899 (N_9899,N_192,N_4110);
or U9900 (N_9900,N_431,N_2415);
nor U9901 (N_9901,N_1524,N_2128);
nand U9902 (N_9902,N_4742,N_1815);
and U9903 (N_9903,N_1181,N_4128);
nor U9904 (N_9904,N_603,N_3361);
nor U9905 (N_9905,N_83,N_2198);
and U9906 (N_9906,N_1157,N_3482);
or U9907 (N_9907,N_754,N_2314);
nor U9908 (N_9908,N_2091,N_1716);
or U9909 (N_9909,N_4958,N_3811);
and U9910 (N_9910,N_2897,N_947);
or U9911 (N_9911,N_363,N_176);
and U9912 (N_9912,N_4014,N_522);
nor U9913 (N_9913,N_4444,N_3871);
nand U9914 (N_9914,N_2347,N_4572);
nor U9915 (N_9915,N_4044,N_27);
or U9916 (N_9916,N_2081,N_3865);
nor U9917 (N_9917,N_2761,N_2212);
nor U9918 (N_9918,N_345,N_2850);
nand U9919 (N_9919,N_745,N_3332);
nor U9920 (N_9920,N_646,N_4646);
nand U9921 (N_9921,N_3621,N_635);
nor U9922 (N_9922,N_2752,N_4483);
nand U9923 (N_9923,N_3398,N_1135);
nor U9924 (N_9924,N_4423,N_4526);
and U9925 (N_9925,N_3636,N_2499);
and U9926 (N_9926,N_3085,N_1604);
nand U9927 (N_9927,N_4431,N_3785);
nor U9928 (N_9928,N_2238,N_1970);
xnor U9929 (N_9929,N_3850,N_925);
nor U9930 (N_9930,N_1317,N_2052);
nand U9931 (N_9931,N_841,N_1996);
and U9932 (N_9932,N_3309,N_3189);
xor U9933 (N_9933,N_2777,N_3122);
nor U9934 (N_9934,N_3771,N_2335);
or U9935 (N_9935,N_2801,N_3846);
nor U9936 (N_9936,N_3066,N_4150);
nand U9937 (N_9937,N_4922,N_2687);
nor U9938 (N_9938,N_3364,N_4685);
and U9939 (N_9939,N_4002,N_3430);
nor U9940 (N_9940,N_1110,N_442);
nor U9941 (N_9941,N_3874,N_4148);
and U9942 (N_9942,N_1912,N_2923);
or U9943 (N_9943,N_2886,N_3481);
or U9944 (N_9944,N_450,N_2054);
and U9945 (N_9945,N_727,N_1276);
or U9946 (N_9946,N_142,N_3988);
or U9947 (N_9947,N_2062,N_4376);
nand U9948 (N_9948,N_35,N_3835);
xor U9949 (N_9949,N_4596,N_396);
or U9950 (N_9950,N_3513,N_644);
and U9951 (N_9951,N_1217,N_445);
and U9952 (N_9952,N_4590,N_1980);
nor U9953 (N_9953,N_194,N_4509);
xnor U9954 (N_9954,N_2175,N_355);
or U9955 (N_9955,N_2232,N_1853);
nand U9956 (N_9956,N_2481,N_4958);
or U9957 (N_9957,N_2291,N_4213);
xnor U9958 (N_9958,N_940,N_1697);
xor U9959 (N_9959,N_2084,N_3755);
and U9960 (N_9960,N_978,N_2358);
or U9961 (N_9961,N_442,N_2296);
and U9962 (N_9962,N_4191,N_2951);
nor U9963 (N_9963,N_1533,N_4191);
nor U9964 (N_9964,N_1218,N_2572);
nand U9965 (N_9965,N_459,N_3524);
nor U9966 (N_9966,N_1778,N_1472);
and U9967 (N_9967,N_3931,N_4936);
nor U9968 (N_9968,N_4561,N_1045);
nor U9969 (N_9969,N_2676,N_2440);
nor U9970 (N_9970,N_3218,N_1953);
and U9971 (N_9971,N_3908,N_981);
or U9972 (N_9972,N_4035,N_1473);
nor U9973 (N_9973,N_359,N_3499);
or U9974 (N_9974,N_1317,N_2498);
or U9975 (N_9975,N_1157,N_3518);
nand U9976 (N_9976,N_1731,N_1694);
nor U9977 (N_9977,N_3002,N_4150);
nand U9978 (N_9978,N_715,N_2178);
nor U9979 (N_9979,N_2444,N_3149);
nand U9980 (N_9980,N_282,N_1551);
nor U9981 (N_9981,N_1670,N_1347);
nor U9982 (N_9982,N_320,N_364);
or U9983 (N_9983,N_3720,N_2060);
nand U9984 (N_9984,N_4519,N_2923);
or U9985 (N_9985,N_3962,N_823);
nand U9986 (N_9986,N_4893,N_862);
nand U9987 (N_9987,N_4048,N_4162);
and U9988 (N_9988,N_1798,N_2158);
nand U9989 (N_9989,N_4286,N_2689);
or U9990 (N_9990,N_2266,N_4199);
nand U9991 (N_9991,N_2083,N_3656);
and U9992 (N_9992,N_4951,N_4890);
and U9993 (N_9993,N_254,N_1129);
nor U9994 (N_9994,N_311,N_1531);
nor U9995 (N_9995,N_1188,N_4708);
or U9996 (N_9996,N_4194,N_1595);
or U9997 (N_9997,N_2110,N_2895);
nor U9998 (N_9998,N_147,N_2496);
or U9999 (N_9999,N_2119,N_1337);
or U10000 (N_10000,N_9682,N_7820);
and U10001 (N_10001,N_6958,N_6001);
and U10002 (N_10002,N_6455,N_8984);
nor U10003 (N_10003,N_6498,N_7116);
nor U10004 (N_10004,N_8280,N_8756);
nor U10005 (N_10005,N_6643,N_7499);
nand U10006 (N_10006,N_5710,N_7785);
nor U10007 (N_10007,N_8772,N_5997);
and U10008 (N_10008,N_8677,N_5291);
nor U10009 (N_10009,N_5620,N_5435);
xor U10010 (N_10010,N_9901,N_8839);
or U10011 (N_10011,N_6217,N_9271);
nand U10012 (N_10012,N_9146,N_6186);
nand U10013 (N_10013,N_8018,N_9610);
xnor U10014 (N_10014,N_5790,N_9140);
nor U10015 (N_10015,N_5563,N_6552);
nor U10016 (N_10016,N_8279,N_8137);
nand U10017 (N_10017,N_6559,N_6508);
nand U10018 (N_10018,N_7057,N_6737);
and U10019 (N_10019,N_5072,N_9126);
nand U10020 (N_10020,N_5244,N_8288);
nor U10021 (N_10021,N_5248,N_8398);
and U10022 (N_10022,N_7452,N_8173);
or U10023 (N_10023,N_6803,N_6931);
nand U10024 (N_10024,N_7309,N_8913);
nand U10025 (N_10025,N_9362,N_6965);
xor U10026 (N_10026,N_8524,N_6959);
nand U10027 (N_10027,N_8066,N_6124);
and U10028 (N_10028,N_8216,N_7350);
or U10029 (N_10029,N_8065,N_5962);
xnor U10030 (N_10030,N_5334,N_6518);
nand U10031 (N_10031,N_8744,N_8833);
xor U10032 (N_10032,N_5888,N_7394);
or U10033 (N_10033,N_6536,N_8121);
nor U10034 (N_10034,N_5611,N_8424);
or U10035 (N_10035,N_5732,N_9612);
nand U10036 (N_10036,N_7544,N_7869);
nor U10037 (N_10037,N_9613,N_6092);
nand U10038 (N_10038,N_7444,N_6037);
or U10039 (N_10039,N_8969,N_7851);
or U10040 (N_10040,N_8761,N_7050);
nand U10041 (N_10041,N_7790,N_7400);
or U10042 (N_10042,N_7634,N_8584);
nor U10043 (N_10043,N_9514,N_9446);
and U10044 (N_10044,N_8778,N_6054);
and U10045 (N_10045,N_9198,N_9205);
or U10046 (N_10046,N_9403,N_9723);
or U10047 (N_10047,N_8974,N_7362);
or U10048 (N_10048,N_7376,N_6221);
nand U10049 (N_10049,N_5613,N_9677);
or U10050 (N_10050,N_9207,N_8990);
and U10051 (N_10051,N_6975,N_8420);
or U10052 (N_10052,N_7220,N_7558);
and U10053 (N_10053,N_6173,N_6806);
or U10054 (N_10054,N_8836,N_7183);
xor U10055 (N_10055,N_7581,N_6757);
nor U10056 (N_10056,N_8393,N_8391);
or U10057 (N_10057,N_8806,N_5541);
and U10058 (N_10058,N_9987,N_6305);
nand U10059 (N_10059,N_5183,N_9460);
nand U10060 (N_10060,N_5296,N_9011);
nor U10061 (N_10061,N_9255,N_6649);
nor U10062 (N_10062,N_5355,N_9998);
xor U10063 (N_10063,N_9374,N_7886);
xnor U10064 (N_10064,N_7887,N_8988);
nand U10065 (N_10065,N_8951,N_8630);
nand U10066 (N_10066,N_6731,N_6886);
nor U10067 (N_10067,N_5109,N_7804);
or U10068 (N_10068,N_9631,N_6500);
and U10069 (N_10069,N_8129,N_7450);
and U10070 (N_10070,N_6497,N_5975);
nand U10071 (N_10071,N_8725,N_8647);
or U10072 (N_10072,N_6279,N_6687);
xor U10073 (N_10073,N_8535,N_8219);
and U10074 (N_10074,N_7111,N_6726);
nor U10075 (N_10075,N_7020,N_6471);
and U10076 (N_10076,N_6817,N_5893);
and U10077 (N_10077,N_9927,N_8710);
nand U10078 (N_10078,N_6101,N_8205);
nor U10079 (N_10079,N_6983,N_6710);
nand U10080 (N_10080,N_9501,N_6699);
nor U10081 (N_10081,N_8010,N_7734);
nand U10082 (N_10082,N_9201,N_7533);
xnor U10083 (N_10083,N_9357,N_7357);
and U10084 (N_10084,N_8114,N_7512);
or U10085 (N_10085,N_6979,N_7794);
nor U10086 (N_10086,N_7210,N_7181);
and U10087 (N_10087,N_8221,N_8662);
and U10088 (N_10088,N_8374,N_8361);
or U10089 (N_10089,N_5836,N_7714);
or U10090 (N_10090,N_9715,N_5476);
nand U10091 (N_10091,N_8252,N_8898);
nand U10092 (N_10092,N_6602,N_6799);
nand U10093 (N_10093,N_8665,N_7761);
and U10094 (N_10094,N_5969,N_7201);
nand U10095 (N_10095,N_7806,N_6556);
or U10096 (N_10096,N_7212,N_7720);
and U10097 (N_10097,N_6769,N_7705);
and U10098 (N_10098,N_8626,N_7534);
or U10099 (N_10099,N_8599,N_8460);
nand U10100 (N_10100,N_7073,N_6107);
and U10101 (N_10101,N_7426,N_8592);
and U10102 (N_10102,N_5167,N_7055);
nor U10103 (N_10103,N_7800,N_6576);
or U10104 (N_10104,N_8384,N_5775);
nand U10105 (N_10105,N_6473,N_5651);
nor U10106 (N_10106,N_9833,N_7489);
nand U10107 (N_10107,N_5579,N_9949);
and U10108 (N_10108,N_8670,N_8959);
nor U10109 (N_10109,N_7672,N_8946);
or U10110 (N_10110,N_5961,N_6600);
or U10111 (N_10111,N_7843,N_6340);
or U10112 (N_10112,N_9928,N_9830);
and U10113 (N_10113,N_7968,N_7241);
nand U10114 (N_10114,N_5370,N_5091);
nor U10115 (N_10115,N_6812,N_6682);
or U10116 (N_10116,N_6314,N_7121);
and U10117 (N_10117,N_5826,N_8566);
and U10118 (N_10118,N_5509,N_9110);
or U10119 (N_10119,N_8038,N_8166);
or U10120 (N_10120,N_5210,N_7580);
nand U10121 (N_10121,N_9442,N_9798);
nand U10122 (N_10122,N_8433,N_6249);
and U10123 (N_10123,N_5442,N_9107);
nand U10124 (N_10124,N_6328,N_5343);
and U10125 (N_10125,N_6333,N_7891);
or U10126 (N_10126,N_5220,N_9111);
and U10127 (N_10127,N_8943,N_9583);
nor U10128 (N_10128,N_8278,N_8754);
and U10129 (N_10129,N_5900,N_9766);
nand U10130 (N_10130,N_8918,N_5913);
and U10131 (N_10131,N_9737,N_5416);
or U10132 (N_10132,N_6964,N_9371);
xnor U10133 (N_10133,N_7985,N_7051);
nor U10134 (N_10134,N_9741,N_5052);
or U10135 (N_10135,N_7262,N_6447);
nand U10136 (N_10136,N_9988,N_9050);
and U10137 (N_10137,N_8523,N_5389);
nand U10138 (N_10138,N_6651,N_6952);
and U10139 (N_10139,N_8203,N_8053);
nor U10140 (N_10140,N_8285,N_6663);
nor U10141 (N_10141,N_7524,N_8704);
nor U10142 (N_10142,N_7448,N_5705);
or U10143 (N_10143,N_8995,N_8124);
or U10144 (N_10144,N_5313,N_6129);
nand U10145 (N_10145,N_8403,N_7488);
nor U10146 (N_10146,N_7956,N_7110);
nor U10147 (N_10147,N_7955,N_8930);
nand U10148 (N_10148,N_6012,N_9762);
nor U10149 (N_10149,N_7633,N_6857);
nor U10150 (N_10150,N_7497,N_8907);
or U10151 (N_10151,N_8183,N_5851);
or U10152 (N_10152,N_8351,N_5184);
nor U10153 (N_10153,N_9237,N_6715);
and U10154 (N_10154,N_9867,N_9210);
nor U10155 (N_10155,N_6316,N_9367);
and U10156 (N_10156,N_6132,N_7716);
nand U10157 (N_10157,N_6199,N_7638);
nor U10158 (N_10158,N_8552,N_6779);
and U10159 (N_10159,N_6689,N_5817);
and U10160 (N_10160,N_6865,N_8953);
or U10161 (N_10161,N_8540,N_9706);
nand U10162 (N_10162,N_5460,N_7003);
and U10163 (N_10163,N_7341,N_5910);
xnor U10164 (N_10164,N_9535,N_5594);
nand U10165 (N_10165,N_9060,N_6111);
nor U10166 (N_10166,N_7102,N_5825);
nor U10167 (N_10167,N_7908,N_6397);
nand U10168 (N_10168,N_7831,N_9168);
nor U10169 (N_10169,N_5265,N_6103);
xnor U10170 (N_10170,N_7276,N_5873);
or U10171 (N_10171,N_7228,N_8174);
nor U10172 (N_10172,N_9980,N_8645);
and U10173 (N_10173,N_7324,N_6187);
and U10174 (N_10174,N_9490,N_7147);
nand U10175 (N_10175,N_9844,N_9123);
and U10176 (N_10176,N_8215,N_5207);
and U10177 (N_10177,N_7996,N_9686);
nand U10178 (N_10178,N_8354,N_6160);
or U10179 (N_10179,N_7875,N_5443);
nand U10180 (N_10180,N_8964,N_7863);
or U10181 (N_10181,N_7514,N_9983);
nand U10182 (N_10182,N_9398,N_7176);
nor U10183 (N_10183,N_6108,N_6493);
or U10184 (N_10184,N_7391,N_7964);
and U10185 (N_10185,N_5070,N_9187);
or U10186 (N_10186,N_9288,N_9618);
nand U10187 (N_10187,N_5506,N_7841);
or U10188 (N_10188,N_6179,N_7648);
or U10189 (N_10189,N_9790,N_8795);
or U10190 (N_10190,N_6872,N_9658);
nor U10191 (N_10191,N_5305,N_5005);
nand U10192 (N_10192,N_8132,N_8171);
nand U10193 (N_10193,N_9996,N_6570);
or U10194 (N_10194,N_8304,N_5168);
or U10195 (N_10195,N_6693,N_9814);
and U10196 (N_10196,N_8887,N_9345);
xor U10197 (N_10197,N_7257,N_7312);
nor U10198 (N_10198,N_8061,N_8711);
nand U10199 (N_10199,N_9315,N_6479);
nand U10200 (N_10200,N_7365,N_9137);
nor U10201 (N_10201,N_8821,N_8227);
nand U10202 (N_10202,N_6357,N_7923);
xor U10203 (N_10203,N_7502,N_7230);
xnor U10204 (N_10204,N_6875,N_9660);
nor U10205 (N_10205,N_9773,N_7373);
and U10206 (N_10206,N_5874,N_6540);
nor U10207 (N_10207,N_8901,N_9426);
nand U10208 (N_10208,N_5129,N_8505);
nand U10209 (N_10209,N_9907,N_8947);
nand U10210 (N_10210,N_6676,N_6572);
nand U10211 (N_10211,N_7811,N_6346);
nand U10212 (N_10212,N_7295,N_9087);
xnor U10213 (N_10213,N_8130,N_8081);
or U10214 (N_10214,N_6580,N_8360);
nor U10215 (N_10215,N_5409,N_7424);
nor U10216 (N_10216,N_6319,N_7197);
nand U10217 (N_10217,N_7000,N_9815);
nand U10218 (N_10218,N_7782,N_6681);
nand U10219 (N_10219,N_6090,N_7553);
nor U10220 (N_10220,N_9871,N_8759);
and U10221 (N_10221,N_6419,N_5427);
nor U10222 (N_10222,N_7208,N_9633);
nand U10223 (N_10223,N_7728,N_7422);
xnor U10224 (N_10224,N_9789,N_5059);
nand U10225 (N_10225,N_7890,N_8924);
or U10226 (N_10226,N_7756,N_6798);
nand U10227 (N_10227,N_7715,N_5062);
nor U10228 (N_10228,N_7285,N_6423);
or U10229 (N_10229,N_6352,N_9223);
nand U10230 (N_10230,N_8100,N_9689);
xnor U10231 (N_10231,N_5281,N_9391);
nand U10232 (N_10232,N_7946,N_8345);
and U10233 (N_10233,N_9749,N_8311);
xor U10234 (N_10234,N_9655,N_6225);
or U10235 (N_10235,N_6792,N_9589);
nand U10236 (N_10236,N_5286,N_6018);
and U10237 (N_10237,N_5469,N_8276);
and U10238 (N_10238,N_5659,N_6030);
and U10239 (N_10239,N_7509,N_5022);
nand U10240 (N_10240,N_5939,N_7069);
nor U10241 (N_10241,N_5478,N_5392);
nand U10242 (N_10242,N_6313,N_5194);
and U10243 (N_10243,N_6810,N_6547);
nor U10244 (N_10244,N_9020,N_8312);
nand U10245 (N_10245,N_8000,N_7308);
xor U10246 (N_10246,N_8620,N_5208);
nor U10247 (N_10247,N_9122,N_5989);
or U10248 (N_10248,N_6863,N_7904);
nand U10249 (N_10249,N_6442,N_6578);
nand U10250 (N_10250,N_5607,N_6456);
nand U10251 (N_10251,N_5235,N_9319);
or U10252 (N_10252,N_8343,N_5852);
nand U10253 (N_10253,N_6521,N_7472);
and U10254 (N_10254,N_6185,N_6711);
nor U10255 (N_10255,N_7433,N_5857);
and U10256 (N_10256,N_8803,N_9886);
nand U10257 (N_10257,N_9429,N_9997);
xor U10258 (N_10258,N_7918,N_7334);
and U10259 (N_10259,N_5742,N_8815);
or U10260 (N_10260,N_6452,N_6192);
nand U10261 (N_10261,N_6200,N_5677);
or U10262 (N_10262,N_7143,N_6283);
and U10263 (N_10263,N_9885,N_7850);
or U10264 (N_10264,N_5876,N_5864);
or U10265 (N_10265,N_5846,N_7937);
and U10266 (N_10266,N_9413,N_6230);
and U10267 (N_10267,N_6685,N_5717);
nor U10268 (N_10268,N_6234,N_6816);
nand U10269 (N_10269,N_9141,N_8199);
or U10270 (N_10270,N_6970,N_7889);
or U10271 (N_10271,N_7703,N_9694);
nand U10272 (N_10272,N_5369,N_9156);
xor U10273 (N_10273,N_7655,N_5716);
nand U10274 (N_10274,N_6315,N_7838);
nor U10275 (N_10275,N_9826,N_6759);
nor U10276 (N_10276,N_5981,N_5588);
and U10277 (N_10277,N_6375,N_5474);
and U10278 (N_10278,N_8147,N_5557);
and U10279 (N_10279,N_5568,N_6180);
nand U10280 (N_10280,N_7588,N_9545);
or U10281 (N_10281,N_7076,N_8963);
and U10282 (N_10282,N_7883,N_7935);
nand U10283 (N_10283,N_9295,N_6936);
nor U10284 (N_10284,N_9400,N_5947);
or U10285 (N_10285,N_5378,N_9214);
nor U10286 (N_10286,N_8870,N_9034);
or U10287 (N_10287,N_6242,N_5995);
and U10288 (N_10288,N_7459,N_9303);
xor U10289 (N_10289,N_6029,N_7454);
and U10290 (N_10290,N_9528,N_5085);
and U10291 (N_10291,N_9144,N_6477);
and U10292 (N_10292,N_6621,N_9019);
nor U10293 (N_10293,N_5123,N_8416);
and U10294 (N_10294,N_9457,N_8299);
nand U10295 (N_10295,N_8232,N_7769);
or U10296 (N_10296,N_7792,N_5880);
nand U10297 (N_10297,N_9129,N_8889);
nor U10298 (N_10298,N_5928,N_5053);
nand U10299 (N_10299,N_6924,N_5759);
nor U10300 (N_10300,N_8683,N_9880);
and U10301 (N_10301,N_8582,N_9347);
or U10302 (N_10302,N_7070,N_6945);
xnor U10303 (N_10303,N_9572,N_9444);
and U10304 (N_10304,N_9729,N_9099);
nand U10305 (N_10305,N_6392,N_9809);
nand U10306 (N_10306,N_7445,N_6465);
and U10307 (N_10307,N_9620,N_6510);
nor U10308 (N_10308,N_7719,N_9623);
and U10309 (N_10309,N_8218,N_9955);
and U10310 (N_10310,N_6083,N_8306);
or U10311 (N_10311,N_6889,N_5735);
nor U10312 (N_10312,N_7387,N_5591);
xnor U10313 (N_10313,N_7346,N_7817);
xor U10314 (N_10314,N_6300,N_7431);
and U10315 (N_10315,N_6318,N_9592);
and U10316 (N_10316,N_8987,N_9910);
xnor U10317 (N_10317,N_6181,N_6366);
xnor U10318 (N_10318,N_5236,N_6987);
or U10319 (N_10319,N_6066,N_8613);
or U10320 (N_10320,N_6396,N_9561);
or U10321 (N_10321,N_9719,N_9093);
xor U10322 (N_10322,N_7893,N_6106);
nand U10323 (N_10323,N_8217,N_9026);
nand U10324 (N_10324,N_8692,N_5252);
and U10325 (N_10325,N_6067,N_8713);
nand U10326 (N_10326,N_6625,N_9654);
nand U10327 (N_10327,N_8243,N_7271);
and U10328 (N_10328,N_7917,N_6172);
nor U10329 (N_10329,N_9119,N_9092);
or U10330 (N_10330,N_5598,N_8511);
or U10331 (N_10331,N_9325,N_6537);
nand U10332 (N_10332,N_6927,N_5672);
nor U10333 (N_10333,N_8423,N_6360);
nor U10334 (N_10334,N_7546,N_9995);
and U10335 (N_10335,N_6027,N_9632);
and U10336 (N_10336,N_8544,N_7818);
nor U10337 (N_10337,N_8534,N_9601);
nand U10338 (N_10338,N_9625,N_7981);
nand U10339 (N_10339,N_5198,N_8895);
or U10340 (N_10340,N_8012,N_7815);
nand U10341 (N_10341,N_9896,N_8547);
nor U10342 (N_10342,N_5934,N_9709);
and U10343 (N_10343,N_5267,N_7897);
or U10344 (N_10344,N_6126,N_8569);
and U10345 (N_10345,N_7282,N_8188);
xnor U10346 (N_10346,N_8631,N_6099);
or U10347 (N_10347,N_6010,N_7407);
and U10348 (N_10348,N_7381,N_5172);
nor U10349 (N_10349,N_5251,N_8496);
and U10350 (N_10350,N_8741,N_9557);
nand U10351 (N_10351,N_7967,N_6058);
or U10352 (N_10352,N_9624,N_5319);
or U10353 (N_10353,N_6407,N_9898);
or U10354 (N_10354,N_8937,N_6361);
and U10355 (N_10355,N_5081,N_7959);
and U10356 (N_10356,N_5794,N_6169);
nor U10357 (N_10357,N_8452,N_5143);
and U10358 (N_10358,N_9285,N_6207);
xnor U10359 (N_10359,N_7449,N_7235);
and U10360 (N_10360,N_5903,N_7601);
nand U10361 (N_10361,N_9616,N_7292);
nand U10362 (N_10362,N_9656,N_5032);
or U10363 (N_10363,N_6436,N_5314);
or U10364 (N_10364,N_5523,N_5942);
and U10365 (N_10365,N_8255,N_7615);
and U10366 (N_10366,N_5350,N_9563);
and U10367 (N_10367,N_6636,N_5652);
xnor U10368 (N_10368,N_6686,N_7636);
and U10369 (N_10369,N_6581,N_7642);
nor U10370 (N_10370,N_6756,N_9619);
nand U10371 (N_10371,N_7567,N_6331);
and U10372 (N_10372,N_7510,N_5170);
and U10373 (N_10373,N_5728,N_7824);
nand U10374 (N_10374,N_7653,N_9862);
or U10375 (N_10375,N_6631,N_6597);
nand U10376 (N_10376,N_9283,N_6563);
nand U10377 (N_10377,N_6868,N_9991);
nand U10378 (N_10378,N_5468,N_7310);
nand U10379 (N_10379,N_8862,N_5375);
nand U10380 (N_10380,N_9127,N_9639);
xor U10381 (N_10381,N_6386,N_5692);
nor U10382 (N_10382,N_9921,N_5706);
and U10383 (N_10383,N_9016,N_5795);
nor U10384 (N_10384,N_5470,N_9363);
nand U10385 (N_10385,N_9978,N_9990);
and U10386 (N_10386,N_8949,N_5429);
and U10387 (N_10387,N_9153,N_8364);
nor U10388 (N_10388,N_8294,N_9351);
nor U10389 (N_10389,N_5572,N_9594);
and U10390 (N_10390,N_5993,N_5016);
nand U10391 (N_10391,N_6146,N_6697);
or U10392 (N_10392,N_7637,N_5655);
nand U10393 (N_10393,N_9189,N_9470);
or U10394 (N_10394,N_6021,N_8347);
nand U10395 (N_10395,N_8138,N_7945);
or U10396 (N_10396,N_5452,N_5423);
and U10397 (N_10397,N_9775,N_9332);
nor U10398 (N_10398,N_8699,N_6734);
nor U10399 (N_10399,N_7977,N_9423);
nand U10400 (N_10400,N_8986,N_6771);
nand U10401 (N_10401,N_7664,N_7019);
xor U10402 (N_10402,N_6212,N_9744);
xnor U10403 (N_10403,N_8356,N_7694);
and U10404 (N_10404,N_9517,N_9106);
nand U10405 (N_10405,N_9160,N_8079);
or U10406 (N_10406,N_5901,N_9902);
xnor U10407 (N_10407,N_5381,N_5240);
and U10408 (N_10408,N_8527,N_8846);
nor U10409 (N_10409,N_9628,N_8708);
or U10410 (N_10410,N_5885,N_8945);
nor U10411 (N_10411,N_9893,N_7864);
nor U10412 (N_10412,N_9309,N_8720);
or U10413 (N_10413,N_8069,N_9232);
and U10414 (N_10414,N_8333,N_9537);
or U10415 (N_10415,N_5786,N_9443);
nor U10416 (N_10416,N_6087,N_6777);
nor U10417 (N_10417,N_8900,N_7816);
nand U10418 (N_10418,N_6155,N_9783);
xnor U10419 (N_10419,N_9086,N_7048);
nand U10420 (N_10420,N_5708,N_6743);
xnor U10421 (N_10421,N_8159,N_6867);
nand U10422 (N_10422,N_8073,N_5639);
nor U10423 (N_10423,N_7539,N_5188);
nand U10424 (N_10424,N_5228,N_8906);
and U10425 (N_10425,N_5077,N_7754);
nor U10426 (N_10426,N_7947,N_6646);
and U10427 (N_10427,N_9191,N_6745);
or U10428 (N_10428,N_5164,N_7594);
and U10429 (N_10429,N_8113,N_6458);
and U10430 (N_10430,N_6229,N_9266);
and U10431 (N_10431,N_9629,N_7040);
and U10432 (N_10432,N_9568,N_6347);
nor U10433 (N_10433,N_9375,N_6809);
nand U10434 (N_10434,N_5593,N_5104);
and U10435 (N_10435,N_6299,N_6684);
and U10436 (N_10436,N_7130,N_9312);
xor U10437 (N_10437,N_6787,N_9870);
and U10438 (N_10438,N_9548,N_8233);
xor U10439 (N_10439,N_7140,N_9681);
or U10440 (N_10440,N_7304,N_5282);
nor U10441 (N_10441,N_6911,N_9876);
or U10442 (N_10442,N_5436,N_7345);
xor U10443 (N_10443,N_8484,N_7011);
nand U10444 (N_10444,N_8742,N_9108);
or U10445 (N_10445,N_6785,N_8490);
and U10446 (N_10446,N_5952,N_6266);
and U10447 (N_10447,N_5567,N_7411);
nand U10448 (N_10448,N_6840,N_9033);
and U10449 (N_10449,N_5219,N_8220);
nand U10450 (N_10450,N_6295,N_5892);
and U10451 (N_10451,N_6635,N_9407);
or U10452 (N_10452,N_6112,N_7700);
nand U10453 (N_10453,N_5936,N_7690);
xnor U10454 (N_10454,N_7015,N_8330);
and U10455 (N_10455,N_8928,N_9738);
and U10456 (N_10456,N_7884,N_9333);
and U10457 (N_10457,N_8024,N_6401);
nor U10458 (N_10458,N_9077,N_7068);
and U10459 (N_10459,N_7265,N_9196);
nor U10460 (N_10460,N_6399,N_5224);
nor U10461 (N_10461,N_8632,N_7298);
nand U10462 (N_10462,N_8181,N_7092);
and U10463 (N_10463,N_9270,N_8673);
and U10464 (N_10464,N_9573,N_5600);
and U10465 (N_10465,N_8378,N_7646);
or U10466 (N_10466,N_8837,N_8973);
or U10467 (N_10467,N_7321,N_8548);
and U10468 (N_10468,N_5003,N_7932);
or U10469 (N_10469,N_5718,N_9455);
nand U10470 (N_10470,N_6391,N_7253);
nand U10471 (N_10471,N_8435,N_7089);
or U10472 (N_10472,N_7957,N_9839);
nand U10473 (N_10473,N_7024,N_6860);
or U10474 (N_10474,N_9912,N_6878);
or U10475 (N_10475,N_5212,N_5619);
nor U10476 (N_10476,N_6919,N_9970);
nor U10477 (N_10477,N_8648,N_9001);
or U10478 (N_10478,N_8515,N_5529);
nand U10479 (N_10479,N_5973,N_7798);
and U10480 (N_10480,N_8428,N_5616);
xor U10481 (N_10481,N_7773,N_5844);
or U10482 (N_10482,N_7106,N_8904);
and U10483 (N_10483,N_5105,N_7369);
and U10484 (N_10484,N_8848,N_5938);
nor U10485 (N_10485,N_6303,N_6906);
nand U10486 (N_10486,N_6138,N_7389);
and U10487 (N_10487,N_9668,N_8606);
and U10488 (N_10488,N_9946,N_6568);
and U10489 (N_10489,N_7991,N_5428);
nor U10490 (N_10490,N_9310,N_7693);
or U10491 (N_10491,N_5080,N_7084);
nand U10492 (N_10492,N_9418,N_7360);
xor U10493 (N_10493,N_8869,N_9697);
and U10494 (N_10494,N_5100,N_5203);
or U10495 (N_10495,N_6893,N_8014);
nand U10496 (N_10496,N_6453,N_8549);
and U10497 (N_10497,N_8856,N_6457);
nor U10498 (N_10498,N_7857,N_5569);
nor U10499 (N_10499,N_5631,N_7914);
xnor U10500 (N_10500,N_8429,N_8163);
and U10501 (N_10501,N_9888,N_6343);
nor U10502 (N_10502,N_5503,N_5534);
nand U10503 (N_10503,N_7666,N_7248);
or U10504 (N_10504,N_6513,N_9989);
and U10505 (N_10505,N_7049,N_5481);
nor U10506 (N_10506,N_7912,N_9804);
or U10507 (N_10507,N_9349,N_9813);
and U10508 (N_10508,N_9414,N_8493);
nand U10509 (N_10509,N_5634,N_5508);
and U10510 (N_10510,N_5397,N_5119);
and U10511 (N_10511,N_9794,N_8057);
nand U10512 (N_10512,N_6877,N_6943);
and U10513 (N_10513,N_9900,N_5618);
nand U10514 (N_10514,N_9641,N_7556);
nand U10515 (N_10515,N_9580,N_6703);
xor U10516 (N_10516,N_6683,N_7576);
or U10517 (N_10517,N_6938,N_5004);
nor U10518 (N_10518,N_6304,N_9268);
xnor U10519 (N_10519,N_9930,N_6105);
nand U10520 (N_10520,N_6899,N_8929);
nand U10521 (N_10521,N_9691,N_6020);
or U10522 (N_10522,N_9436,N_6036);
nor U10523 (N_10523,N_5801,N_8580);
nand U10524 (N_10524,N_7962,N_9750);
nand U10525 (N_10525,N_5411,N_6739);
and U10526 (N_10526,N_7674,N_7085);
nor U10527 (N_10527,N_6741,N_9139);
or U10528 (N_10528,N_6415,N_5527);
or U10529 (N_10529,N_5514,N_6818);
or U10530 (N_10530,N_9031,N_6384);
and U10531 (N_10531,N_8482,N_9558);
nor U10532 (N_10532,N_5537,N_5384);
and U10533 (N_10533,N_7135,N_6292);
or U10534 (N_10534,N_6424,N_6884);
nand U10535 (N_10535,N_6444,N_7986);
nor U10536 (N_10536,N_8197,N_6434);
nor U10537 (N_10537,N_8871,N_9837);
nor U10538 (N_10538,N_8338,N_9835);
nor U10539 (N_10539,N_7168,N_5241);
nand U10540 (N_10540,N_8178,N_9287);
and U10541 (N_10541,N_8878,N_5983);
or U10542 (N_10542,N_9530,N_5408);
or U10543 (N_10543,N_6031,N_5871);
nor U10544 (N_10544,N_7742,N_7237);
nand U10545 (N_10545,N_9832,N_6463);
nor U10546 (N_10546,N_7795,N_8234);
and U10547 (N_10547,N_5636,N_7108);
or U10548 (N_10548,N_9748,N_7347);
or U10549 (N_10549,N_6940,N_8526);
xor U10550 (N_10550,N_6408,N_8175);
or U10551 (N_10551,N_9204,N_6516);
xor U10552 (N_10552,N_9653,N_8115);
and U10553 (N_10553,N_8244,N_8044);
xnor U10554 (N_10554,N_9133,N_7151);
xor U10555 (N_10555,N_6275,N_8764);
nor U10556 (N_10556,N_6280,N_5299);
or U10557 (N_10557,N_7207,N_6015);
or U10558 (N_10558,N_9387,N_8143);
xnor U10559 (N_10559,N_8767,N_9821);
nor U10560 (N_10560,N_7590,N_6113);
and U10561 (N_10561,N_9569,N_8139);
nand U10562 (N_10562,N_6095,N_5830);
and U10563 (N_10563,N_5917,N_6696);
and U10564 (N_10564,N_7949,N_8853);
nor U10565 (N_10565,N_5342,N_8274);
and U10566 (N_10566,N_8284,N_5891);
and U10567 (N_10567,N_5498,N_7934);
nor U10568 (N_10568,N_9416,N_9702);
nand U10569 (N_10569,N_9074,N_8779);
or U10570 (N_10570,N_8576,N_7430);
and U10571 (N_10571,N_8142,N_6653);
or U10572 (N_10572,N_5524,N_9012);
and U10573 (N_10573,N_6749,N_7215);
and U10574 (N_10574,N_9769,N_9431);
nand U10575 (N_10575,N_8322,N_8735);
and U10576 (N_10576,N_9688,N_9136);
nor U10577 (N_10577,N_5657,N_7120);
nor U10578 (N_10578,N_7498,N_7293);
nand U10579 (N_10579,N_6993,N_9959);
xnor U10580 (N_10580,N_8619,N_9952);
nand U10581 (N_10581,N_8168,N_8908);
nor U10582 (N_10582,N_9021,N_5012);
nor U10583 (N_10583,N_6907,N_9932);
or U10584 (N_10584,N_6835,N_8030);
nor U10585 (N_10585,N_6278,N_7606);
and U10586 (N_10586,N_5178,N_6923);
and U10587 (N_10587,N_5605,N_8983);
nand U10588 (N_10588,N_6606,N_9247);
and U10589 (N_10589,N_9745,N_9599);
nor U10590 (N_10590,N_6057,N_6727);
or U10591 (N_10591,N_9307,N_7175);
and U10592 (N_10592,N_5079,N_9342);
and U10593 (N_10593,N_7583,N_7078);
and U10594 (N_10594,N_6820,N_5287);
and U10595 (N_10595,N_8119,N_5603);
and U10596 (N_10596,N_9974,N_5124);
xor U10597 (N_10597,N_6776,N_5863);
or U10598 (N_10598,N_7368,N_9575);
or U10599 (N_10599,N_7617,N_7349);
or U10600 (N_10600,N_6024,N_5204);
and U10601 (N_10601,N_9385,N_9704);
xor U10602 (N_10602,N_7425,N_7086);
and U10603 (N_10603,N_7840,N_9167);
or U10604 (N_10604,N_8865,N_5150);
and U10605 (N_10605,N_7401,N_8885);
nand U10606 (N_10606,N_9317,N_6664);
or U10607 (N_10607,N_9468,N_9726);
or U10608 (N_10608,N_8157,N_8303);
and U10609 (N_10609,N_8679,N_8530);
nand U10610 (N_10610,N_7245,N_8068);
and U10611 (N_10611,N_6495,N_7320);
or U10612 (N_10612,N_9405,N_5261);
and U10613 (N_10613,N_6862,N_9199);
or U10614 (N_10614,N_8007,N_6584);
and U10615 (N_10615,N_8457,N_7418);
nor U10616 (N_10616,N_7683,N_6752);
xor U10617 (N_10617,N_7468,N_7788);
nor U10618 (N_10618,N_5459,N_6289);
nor U10619 (N_10619,N_7406,N_5043);
nor U10620 (N_10620,N_5711,N_5813);
and U10621 (N_10621,N_5784,N_7236);
nor U10622 (N_10622,N_9734,N_7097);
and U10623 (N_10623,N_5930,N_9277);
nor U10624 (N_10624,N_5226,N_8337);
or U10625 (N_10625,N_5859,N_8230);
or U10626 (N_10626,N_7557,N_7187);
nand U10627 (N_10627,N_8798,N_5816);
or U10628 (N_10628,N_8155,N_9985);
nor U10629 (N_10629,N_6822,N_5028);
or U10630 (N_10630,N_7584,N_5294);
nor U10631 (N_10631,N_7198,N_7860);
xor U10632 (N_10632,N_6788,N_9151);
and U10633 (N_10633,N_8664,N_6220);
nor U10634 (N_10634,N_9101,N_9382);
nand U10635 (N_10635,N_6459,N_8118);
or U10636 (N_10636,N_7340,N_5785);
or U10637 (N_10637,N_9499,N_8323);
xor U10638 (N_10638,N_6454,N_9439);
and U10639 (N_10639,N_7910,N_9577);
nand U10640 (N_10640,N_7410,N_8801);
or U10641 (N_10641,N_6512,N_5833);
and U10642 (N_10642,N_6910,N_9354);
nor U10643 (N_10643,N_7593,N_5078);
and U10644 (N_10644,N_9194,N_5345);
or U10645 (N_10645,N_9510,N_6520);
and U10646 (N_10646,N_7592,N_6897);
nor U10647 (N_10647,N_8872,N_7054);
xnor U10648 (N_10648,N_7808,N_9705);
or U10649 (N_10649,N_9611,N_6364);
or U10650 (N_10650,N_7744,N_8023);
or U10651 (N_10651,N_6484,N_8637);
nor U10652 (N_10652,N_9954,N_7982);
or U10653 (N_10653,N_9329,N_9904);
or U10654 (N_10654,N_8093,N_9296);
and U10655 (N_10655,N_9609,N_9840);
nand U10656 (N_10656,N_5589,N_6336);
or U10657 (N_10657,N_9768,N_5766);
and U10658 (N_10658,N_7170,N_6744);
nand U10659 (N_10659,N_9258,N_5387);
nor U10660 (N_10660,N_5205,N_6933);
nand U10661 (N_10661,N_8531,N_9780);
nand U10662 (N_10662,N_7486,N_9918);
or U10663 (N_10663,N_5215,N_8029);
or U10664 (N_10664,N_8196,N_6690);
or U10665 (N_10665,N_5805,N_7481);
nand U10666 (N_10666,N_6335,N_9117);
xor U10667 (N_10667,N_9846,N_8293);
nor U10668 (N_10668,N_9331,N_7273);
or U10669 (N_10669,N_5686,N_9155);
or U10670 (N_10670,N_8458,N_9712);
and U10671 (N_10671,N_5434,N_5780);
nand U10672 (N_10672,N_5074,N_5363);
and U10673 (N_10673,N_9700,N_5367);
and U10674 (N_10674,N_6732,N_9121);
or U10675 (N_10675,N_8561,N_9588);
nor U10676 (N_10676,N_5041,N_5040);
and U10677 (N_10677,N_8120,N_6309);
and U10678 (N_10678,N_5309,N_6383);
nand U10679 (N_10679,N_9593,N_8257);
xnor U10680 (N_10680,N_8717,N_8840);
nor U10681 (N_10681,N_6592,N_7263);
nor U10682 (N_10682,N_7184,N_5504);
nand U10683 (N_10683,N_5615,N_5929);
or U10684 (N_10684,N_6879,N_5406);
and U10685 (N_10685,N_7755,N_6260);
xnor U10686 (N_10686,N_5561,N_8671);
xnor U10687 (N_10687,N_9130,N_9071);
and U10688 (N_10688,N_7064,N_5758);
or U10689 (N_10689,N_5200,N_7699);
or U10690 (N_10690,N_7153,N_9509);
nand U10691 (N_10691,N_7164,N_5665);
nor U10692 (N_10692,N_9699,N_8989);
nor U10693 (N_10693,N_5823,N_6104);
nand U10694 (N_10694,N_5617,N_9939);
nor U10695 (N_10695,N_6740,N_7178);
nand U10696 (N_10696,N_7663,N_6688);
nand U10697 (N_10697,N_7905,N_7735);
nor U10698 (N_10698,N_6332,N_9878);
nand U10699 (N_10699,N_8604,N_7122);
or U10700 (N_10700,N_5576,N_6937);
or U10701 (N_10701,N_9463,N_6846);
and U10702 (N_10702,N_5610,N_7413);
nand U10703 (N_10703,N_8162,N_5133);
xor U10704 (N_10704,N_6842,N_9526);
nor U10705 (N_10705,N_8618,N_6143);
xnor U10706 (N_10706,N_8198,N_5582);
and U10707 (N_10707,N_9038,N_8650);
or U10708 (N_10708,N_9147,N_8944);
nor U10709 (N_10709,N_7014,N_9067);
and U10710 (N_10710,N_5792,N_7338);
or U10711 (N_10711,N_6470,N_6022);
or U10712 (N_10712,N_9056,N_8058);
or U10713 (N_10713,N_6374,N_8745);
nor U10714 (N_10714,N_8783,N_5925);
and U10715 (N_10715,N_5673,N_8088);
nand U10716 (N_10716,N_5723,N_7760);
and U10717 (N_10717,N_9824,N_8408);
or U10718 (N_10718,N_7574,N_7704);
or U10719 (N_10719,N_9947,N_7723);
nand U10720 (N_10720,N_5746,N_9228);
nor U10721 (N_10721,N_6089,N_6953);
or U10722 (N_10722,N_6645,N_9399);
nand U10723 (N_10723,N_6308,N_6141);
nor U10724 (N_10724,N_9890,N_8655);
nor U10725 (N_10725,N_9234,N_7399);
xor U10726 (N_10726,N_5904,N_7112);
and U10727 (N_10727,N_8316,N_7239);
or U10728 (N_10728,N_6834,N_6698);
and U10729 (N_10729,N_7667,N_7246);
nand U10730 (N_10730,N_6789,N_9104);
or U10731 (N_10731,N_9213,N_5014);
and U10732 (N_10732,N_8451,N_6675);
and U10733 (N_10733,N_6094,N_7903);
or U10734 (N_10734,N_8706,N_5051);
nand U10735 (N_10735,N_6069,N_9145);
xor U10736 (N_10736,N_6102,N_9581);
or U10737 (N_10737,N_6515,N_7087);
nand U10738 (N_10738,N_5463,N_5437);
or U10739 (N_10739,N_6211,N_5991);
or U10740 (N_10740,N_8697,N_6793);
xor U10741 (N_10741,N_6499,N_8852);
xnor U10742 (N_10742,N_7862,N_5256);
nand U10743 (N_10743,N_8858,N_6369);
and U10744 (N_10744,N_9235,N_9648);
and U10745 (N_10745,N_7222,N_5703);
xnor U10746 (N_10746,N_9152,N_6116);
or U10747 (N_10747,N_6322,N_6035);
xor U10748 (N_10748,N_6514,N_7036);
and U10749 (N_10749,N_9822,N_8194);
or U10750 (N_10750,N_5181,N_8200);
nand U10751 (N_10751,N_9497,N_6858);
and U10752 (N_10752,N_7819,N_9516);
nand U10753 (N_10753,N_6504,N_5103);
or U10754 (N_10754,N_7163,N_9269);
nand U10755 (N_10755,N_6669,N_5421);
and U10756 (N_10756,N_6760,N_7527);
xor U10757 (N_10757,N_6705,N_6550);
nor U10758 (N_10758,N_6237,N_5838);
nand U10759 (N_10759,N_5066,N_8577);
nor U10760 (N_10760,N_8389,N_5831);
and U10761 (N_10761,N_7585,N_5979);
nand U10762 (N_10762,N_5811,N_5837);
xor U10763 (N_10763,N_6182,N_8594);
and U10764 (N_10764,N_8617,N_9365);
nand U10765 (N_10765,N_7272,N_9934);
nand U10766 (N_10766,N_6722,N_5869);
or U10767 (N_10767,N_6265,N_9097);
or U10768 (N_10768,N_7277,N_5512);
nor U10769 (N_10769,N_9542,N_7119);
or U10770 (N_10770,N_9771,N_9976);
nand U10771 (N_10771,N_9817,N_8317);
or U10772 (N_10772,N_5698,N_9438);
xor U10773 (N_10773,N_6209,N_7420);
and U10774 (N_10774,N_7953,N_8636);
and U10775 (N_10775,N_8541,N_6794);
nor U10776 (N_10776,N_8241,N_5747);
and U10777 (N_10777,N_6579,N_5690);
nand U10778 (N_10778,N_6511,N_9180);
or U10779 (N_10779,N_7781,N_7823);
and U10780 (N_10780,N_5024,N_9380);
or U10781 (N_10781,N_6390,N_9243);
and U10782 (N_10782,N_6824,N_6900);
and U10783 (N_10783,N_9936,N_9554);
and U10784 (N_10784,N_8103,N_6253);
xnor U10785 (N_10785,N_9208,N_5623);
or U10786 (N_10786,N_8593,N_5417);
or U10787 (N_10787,N_7259,N_7825);
xnor U10788 (N_10788,N_6236,N_8629);
nor U10789 (N_10789,N_7473,N_9458);
nor U10790 (N_10790,N_7463,N_6342);
nand U10791 (N_10791,N_8681,N_7372);
or U10792 (N_10792,N_7763,N_6065);
nand U10793 (N_10793,N_7307,N_6575);
nand U10794 (N_10794,N_8897,N_9883);
nor U10795 (N_10795,N_8657,N_7865);
nand U10796 (N_10796,N_8881,N_6348);
and U10797 (N_10797,N_6638,N_8026);
nor U10798 (N_10798,N_9472,N_5848);
or U10799 (N_10799,N_8208,N_8635);
or U10800 (N_10800,N_8250,N_6898);
nand U10801 (N_10801,N_9163,N_8542);
nand U10802 (N_10802,N_9286,N_7202);
or U10803 (N_10803,N_7283,N_7987);
and U10804 (N_10804,N_5960,N_5325);
nor U10805 (N_10805,N_7126,N_6659);
and U10806 (N_10806,N_8994,N_9401);
xor U10807 (N_10807,N_5788,N_6833);
nor U10808 (N_10808,N_7989,N_6255);
nor U10809 (N_10809,N_5592,N_5097);
and U10810 (N_10810,N_7777,N_6539);
nor U10811 (N_10811,N_7204,N_6014);
xor U10812 (N_10812,N_8453,N_5559);
nand U10813 (N_10813,N_6821,N_6282);
or U10814 (N_10814,N_5490,N_9273);
nor U10815 (N_10815,N_9061,N_7861);
nor U10816 (N_10816,N_7005,N_6201);
and U10817 (N_10817,N_7973,N_9854);
nor U10818 (N_10818,N_6660,N_5357);
nor U10819 (N_10819,N_8290,N_5552);
and U10820 (N_10820,N_9328,N_5632);
and U10821 (N_10821,N_7939,N_8329);
nand U10822 (N_10822,N_8884,N_6607);
or U10823 (N_10823,N_7670,N_6624);
or U10824 (N_10824,N_5755,N_8954);
nand U10825 (N_10825,N_8757,N_6738);
or U10826 (N_10826,N_5719,N_6291);
nor U10827 (N_10827,N_5695,N_9017);
and U10828 (N_10828,N_6425,N_6222);
nor U10829 (N_10829,N_6231,N_9874);
and U10830 (N_10830,N_7998,N_8092);
or U10831 (N_10831,N_5879,N_8567);
and U10832 (N_10832,N_9063,N_9456);
nand U10833 (N_10833,N_5418,N_7453);
and U10834 (N_10834,N_6677,N_8686);
nand U10835 (N_10835,N_9353,N_8955);
and U10836 (N_10836,N_8883,N_8459);
nand U10837 (N_10837,N_5754,N_7545);
and U10838 (N_10838,N_5160,N_8830);
or U10839 (N_10839,N_6673,N_6330);
and U10840 (N_10840,N_6373,N_7995);
or U10841 (N_10841,N_9650,N_9747);
xor U10842 (N_10842,N_8842,N_8857);
and U10843 (N_10843,N_8899,N_5399);
nand U10844 (N_10844,N_6487,N_7098);
or U10845 (N_10845,N_9465,N_5380);
nand U10846 (N_10846,N_6864,N_6531);
and U10847 (N_10847,N_6784,N_8522);
or U10848 (N_10848,N_9066,N_9221);
and U10849 (N_10849,N_9662,N_8775);
xor U10850 (N_10850,N_8078,N_9448);
or U10851 (N_10851,N_8888,N_6403);
and U10852 (N_10852,N_8916,N_5311);
and U10853 (N_10853,N_6585,N_6674);
and U10854 (N_10854,N_5733,N_7254);
nor U10855 (N_10855,N_8753,N_8845);
and U10856 (N_10856,N_6202,N_9049);
and U10857 (N_10857,N_5084,N_7948);
and U10858 (N_10858,N_8529,N_6163);
or U10859 (N_10859,N_5453,N_6198);
nor U10860 (N_10860,N_5186,N_8236);
and U10861 (N_10861,N_5201,N_6854);
nor U10862 (N_10862,N_8893,N_9919);
nor U10863 (N_10863,N_7733,N_8270);
or U10864 (N_10864,N_7711,N_8956);
nor U10865 (N_10865,N_9320,N_8480);
nand U10866 (N_10866,N_6387,N_7194);
and U10867 (N_10867,N_9389,N_9197);
or U10868 (N_10868,N_9437,N_9856);
nand U10869 (N_10869,N_6149,N_8379);
and U10870 (N_10870,N_9791,N_5911);
and U10871 (N_10871,N_9657,N_8562);
and U10872 (N_10872,N_8941,N_5142);
nand U10873 (N_10873,N_7739,N_6825);
nor U10874 (N_10874,N_5666,N_7214);
or U10875 (N_10875,N_5640,N_8473);
nand U10876 (N_10876,N_5625,N_5835);
xor U10877 (N_10877,N_8359,N_9183);
nand U10878 (N_10878,N_9703,N_8222);
nor U10879 (N_10879,N_8812,N_9029);
or U10880 (N_10880,N_7680,N_8497);
and U10881 (N_10881,N_9082,N_9215);
xor U10882 (N_10882,N_5931,N_6586);
nand U10883 (N_10883,N_7722,N_6766);
nor U10884 (N_10884,N_7231,N_6704);
nand U10885 (N_10885,N_8736,N_5669);
xor U10886 (N_10886,N_9924,N_8396);
nor U10887 (N_10887,N_7004,N_7892);
and U10888 (N_10888,N_9850,N_6721);
and U10889 (N_10889,N_6250,N_5922);
and U10890 (N_10890,N_6059,N_5887);
nand U10891 (N_10891,N_8765,N_5714);
nor U10892 (N_10892,N_9687,N_9267);
nor U10893 (N_10893,N_6986,N_7461);
or U10894 (N_10894,N_5691,N_9428);
and U10895 (N_10895,N_5297,N_5454);
or U10896 (N_10896,N_9238,N_5285);
nor U10897 (N_10897,N_7921,N_5401);
nand U10898 (N_10898,N_9666,N_8302);
xor U10899 (N_10899,N_5587,N_9579);
or U10900 (N_10900,N_9427,N_5635);
nor U10901 (N_10901,N_6990,N_8319);
xnor U10902 (N_10902,N_8334,N_9627);
nor U10903 (N_10903,N_5413,N_5222);
nor U10904 (N_10904,N_9925,N_7191);
xnor U10905 (N_10905,N_6405,N_6023);
nand U10906 (N_10906,N_5612,N_9292);
nand U10907 (N_10907,N_8324,N_5430);
and U10908 (N_10908,N_6962,N_5199);
nor U10909 (N_10909,N_6998,N_8309);
nand U10910 (N_10910,N_5762,N_6117);
or U10911 (N_10911,N_6524,N_9828);
nand U10912 (N_10912,N_7503,N_5977);
nor U10913 (N_10913,N_5480,N_8090);
nand U10914 (N_10914,N_7589,N_9742);
or U10915 (N_10915,N_7779,N_6672);
or U10916 (N_10916,N_5528,N_7942);
or U10917 (N_10917,N_5393,N_6241);
nor U10918 (N_10918,N_8977,N_8320);
nor U10919 (N_10919,N_5300,N_8975);
or U10920 (N_10920,N_9290,N_7778);
nand U10921 (N_10921,N_5360,N_8358);
nor U10922 (N_10922,N_5112,N_7396);
or U10923 (N_10923,N_9219,N_9339);
nand U10924 (N_10924,N_6232,N_6971);
and U10925 (N_10925,N_7684,N_6978);
nor U10926 (N_10926,N_8056,N_7894);
or U10927 (N_10927,N_7659,N_6901);
nor U10928 (N_10928,N_8439,N_9531);
xnor U10929 (N_10929,N_7644,N_6505);
xnor U10930 (N_10930,N_6995,N_7495);
nand U10931 (N_10931,N_8472,N_7626);
and U10932 (N_10932,N_9085,N_5566);
or U10933 (N_10933,N_6238,N_5477);
nand U10934 (N_10934,N_9432,N_5633);
nor U10935 (N_10935,N_9651,N_7137);
nor U10936 (N_10936,N_9217,N_6358);
or U10937 (N_10937,N_8950,N_7067);
or U10938 (N_10938,N_9721,N_6839);
nor U10939 (N_10939,N_9582,N_7243);
xnor U10940 (N_10940,N_7535,N_5606);
or U10941 (N_10941,N_7922,N_9743);
nand U10942 (N_10942,N_8981,N_5643);
and U10943 (N_10943,N_7171,N_5779);
or U10944 (N_10944,N_6338,N_7434);
nand U10945 (N_10945,N_5025,N_7035);
and U10946 (N_10946,N_6610,N_8532);
nand U10947 (N_10947,N_7543,N_5658);
xnor U10948 (N_10948,N_9000,N_7034);
or U10949 (N_10949,N_6541,N_7552);
nand U10950 (N_10950,N_5191,N_8729);
nor U10951 (N_10951,N_6713,N_6344);
xnor U10952 (N_10952,N_6474,N_6062);
or U10953 (N_10953,N_5959,N_8667);
nand U10954 (N_10954,N_8514,N_5140);
or U10955 (N_10955,N_8313,N_5675);
and U10956 (N_10956,N_5940,N_6605);
nor U10957 (N_10957,N_5055,N_9984);
or U10958 (N_10958,N_9047,N_8520);
or U10959 (N_10959,N_7319,N_6984);
nor U10960 (N_10960,N_5697,N_5180);
or U10961 (N_10961,N_9895,N_9590);
or U10962 (N_10962,N_6353,N_8261);
or U10963 (N_10963,N_8587,N_6702);
nand U10964 (N_10964,N_9473,N_7105);
xor U10965 (N_10965,N_5667,N_7560);
or U10966 (N_10966,N_8585,N_9209);
nor U10967 (N_10967,N_9647,N_9182);
and U10968 (N_10968,N_5302,N_8380);
and U10969 (N_10969,N_6819,N_7037);
or U10970 (N_10970,N_7506,N_6100);
nor U10971 (N_10971,N_5058,N_6003);
xnor U10972 (N_10972,N_6145,N_9502);
and U10973 (N_10973,N_5685,N_9336);
or U10974 (N_10974,N_8911,N_8321);
or U10975 (N_10975,N_8112,N_9801);
nor U10976 (N_10976,N_6418,N_9511);
xor U10977 (N_10977,N_6564,N_8160);
nand U10978 (N_10978,N_7072,N_5185);
and U10979 (N_10979,N_6385,N_9975);
or U10980 (N_10980,N_8595,N_5553);
or U10981 (N_10981,N_7602,N_5162);
nand U10982 (N_10982,N_8926,N_7058);
or U10983 (N_10983,N_6811,N_9797);
or U10984 (N_10984,N_7847,N_6826);
nor U10985 (N_10985,N_5538,N_9043);
or U10986 (N_10986,N_6678,N_5834);
nor U10987 (N_10987,N_5599,N_8774);
and U10988 (N_10988,N_7925,N_9184);
or U10989 (N_10989,N_5777,N_6655);
nor U10990 (N_10990,N_6929,N_8649);
nor U10991 (N_10991,N_7109,N_9906);
and U10992 (N_10992,N_7582,N_9968);
nand U10993 (N_10993,N_7686,N_8751);
and U10994 (N_10994,N_6085,N_6560);
and U10995 (N_10995,N_9479,N_5963);
nand U10996 (N_10996,N_8340,N_6502);
nand U10997 (N_10997,N_7866,N_8447);
and U10998 (N_10998,N_7104,N_9202);
nand U10999 (N_10999,N_7358,N_5361);
nor U11000 (N_11000,N_5584,N_8982);
or U11001 (N_11001,N_5560,N_7500);
nand U11002 (N_11002,N_8247,N_6311);
and U11003 (N_11003,N_6650,N_6701);
nand U11004 (N_11004,N_8478,N_9233);
nand U11005 (N_11005,N_9960,N_6748);
and U11006 (N_11006,N_5254,N_6081);
nor U11007 (N_11007,N_5280,N_6052);
nand U11008 (N_11008,N_8554,N_9305);
or U11009 (N_11009,N_8060,N_8651);
and U11010 (N_11010,N_8962,N_8033);
nand U11011 (N_11011,N_9177,N_7620);
nor U11012 (N_11012,N_6733,N_6074);
nand U11013 (N_11013,N_7195,N_6203);
nor U11014 (N_11014,N_5899,N_5660);
nor U11015 (N_11015,N_8992,N_8504);
nand U11016 (N_11016,N_7377,N_8153);
and U11017 (N_11017,N_9226,N_8960);
nor U11018 (N_11018,N_8350,N_7853);
or U11019 (N_11019,N_6019,N_5764);
and U11020 (N_11020,N_5424,N_7605);
and U11021 (N_11021,N_7063,N_7979);
nor U11022 (N_11022,N_9105,N_7745);
and U11023 (N_11023,N_5414,N_9143);
or U11024 (N_11024,N_7152,N_5516);
and U11025 (N_11025,N_8684,N_5941);
nand U11026 (N_11026,N_7771,N_5847);
nand U11027 (N_11027,N_8461,N_8070);
nand U11028 (N_11028,N_8659,N_9293);
nor U11029 (N_11029,N_8371,N_6040);
nand U11030 (N_11030,N_5750,N_8310);
nand U11031 (N_11031,N_9178,N_6891);
nand U11032 (N_11032,N_9059,N_7736);
nor U11033 (N_11033,N_9964,N_9676);
nand U11034 (N_11034,N_9596,N_5702);
and U11035 (N_11035,N_7289,N_5485);
nand U11036 (N_11036,N_9109,N_8305);
xor U11037 (N_11037,N_6764,N_9792);
and U11038 (N_11038,N_7765,N_5681);
or U11039 (N_11039,N_7837,N_6797);
nor U11040 (N_11040,N_5824,N_9381);
nor U11041 (N_11041,N_8799,N_7113);
nand U11042 (N_11042,N_7211,N_8039);
xor U11043 (N_11043,N_7267,N_8165);
nor U11044 (N_11044,N_7209,N_8724);
xnor U11045 (N_11045,N_6426,N_9256);
nand U11046 (N_11046,N_5680,N_9621);
or U11047 (N_11047,N_9776,N_6644);
xor U11048 (N_11048,N_5927,N_8972);
or U11049 (N_11049,N_6608,N_7306);
xnor U11050 (N_11050,N_6873,N_8076);
and U11051 (N_11051,N_7661,N_9040);
and U11052 (N_11052,N_9795,N_5909);
nor U11053 (N_11053,N_9007,N_5676);
xor U11054 (N_11054,N_7355,N_9386);
and U11055 (N_11055,N_7915,N_7687);
or U11056 (N_11056,N_5951,N_6150);
nor U11057 (N_11057,N_9962,N_7189);
xor U11058 (N_11058,N_9028,N_8824);
or U11059 (N_11059,N_7185,N_9622);
nor U11060 (N_11060,N_9172,N_5151);
or U11061 (N_11061,N_8489,N_9785);
and U11062 (N_11062,N_9388,N_6996);
nor U11063 (N_11063,N_7740,N_8405);
nand U11064 (N_11064,N_7482,N_6802);
nand U11065 (N_11065,N_8718,N_7487);
nand U11066 (N_11066,N_8150,N_9920);
nor U11067 (N_11067,N_7548,N_5064);
nand U11068 (N_11068,N_9482,N_8510);
and U11069 (N_11069,N_7266,N_6587);
nand U11070 (N_11070,N_5021,N_6920);
and U11071 (N_11071,N_6949,N_7849);
nor U11072 (N_11072,N_7870,N_5789);
nor U11073 (N_11073,N_8537,N_8251);
xnor U11074 (N_11074,N_9778,N_6227);
and U11075 (N_11075,N_9135,N_9236);
nor U11076 (N_11076,N_6259,N_8826);
nor U11077 (N_11077,N_9680,N_8040);
and U11078 (N_11078,N_6977,N_7460);
nor U11079 (N_11079,N_6196,N_7250);
and U11080 (N_11080,N_6583,N_6480);
and U11081 (N_11081,N_6056,N_8920);
and U11082 (N_11082,N_9076,N_8368);
nand U11083 (N_11083,N_8253,N_7247);
nand U11084 (N_11084,N_6895,N_6380);
or U11085 (N_11085,N_8268,N_7562);
or U11086 (N_11086,N_6034,N_6954);
or U11087 (N_11087,N_8008,N_8032);
nand U11088 (N_11088,N_5382,N_8466);
nor U11089 (N_11089,N_7233,N_6302);
nand U11090 (N_11090,N_5332,N_9330);
or U11091 (N_11091,N_7090,N_9262);
nor U11092 (N_11092,N_7132,N_5482);
nand U11093 (N_11093,N_7417,N_9103);
nor U11094 (N_11094,N_5001,N_6000);
nand U11095 (N_11095,N_5753,N_7940);
or U11096 (N_11096,N_5141,N_8864);
nor U11097 (N_11097,N_6287,N_5148);
nand U11098 (N_11098,N_9845,N_9836);
nand U11099 (N_11099,N_9276,N_8094);
xnor U11100 (N_11100,N_7821,N_9073);
xor U11101 (N_11101,N_6147,N_8518);
nor U11102 (N_11102,N_6969,N_9230);
or U11103 (N_11103,N_5486,N_5757);
or U11104 (N_11104,N_7317,N_5348);
or U11105 (N_11105,N_7141,N_6871);
and U11106 (N_11106,N_8055,N_6047);
xor U11107 (N_11107,N_8190,N_7335);
or U11108 (N_11108,N_5915,N_8811);
nor U11109 (N_11109,N_9852,N_9803);
nand U11110 (N_11110,N_5866,N_8676);
or U11111 (N_11111,N_9851,N_8663);
or U11112 (N_11112,N_5099,N_9586);
nand U11113 (N_11113,N_5288,N_6562);
and U11114 (N_11114,N_8022,N_7354);
nor U11115 (N_11115,N_8939,N_8780);
or U11116 (N_11116,N_7958,N_7297);
or U11117 (N_11117,N_9942,N_8192);
nand U11118 (N_11118,N_6377,N_8440);
or U11119 (N_11119,N_8810,N_9505);
nor U11120 (N_11120,N_5731,N_5039);
and U11121 (N_11121,N_8819,N_6329);
or U11122 (N_11122,N_9297,N_8410);
and U11123 (N_11123,N_8672,N_8449);
or U11124 (N_11124,N_9006,N_6096);
xor U11125 (N_11125,N_6614,N_5125);
and U11126 (N_11126,N_5894,N_9923);
nand U11127 (N_11127,N_6700,N_7388);
or U11128 (N_11128,N_7885,N_5609);
nand U11129 (N_11129,N_9760,N_6558);
nor U11130 (N_11130,N_6507,N_8156);
and U11131 (N_11131,N_5111,N_7954);
or U11132 (N_11132,N_9764,N_6195);
nor U11133 (N_11133,N_9170,N_5574);
xor U11134 (N_11134,N_6432,N_8553);
nor U11135 (N_11135,N_5374,N_8912);
and U11136 (N_11136,N_5575,N_8787);
or U11137 (N_11137,N_6154,N_6032);
nand U11138 (N_11138,N_8998,N_6888);
xor U11139 (N_11139,N_5744,N_5377);
and U11140 (N_11140,N_8127,N_7789);
and U11141 (N_11141,N_7061,N_5173);
nand U11142 (N_11142,N_8719,N_5497);
nand U11143 (N_11143,N_5127,N_5161);
or U11144 (N_11144,N_8749,N_6533);
nand U11145 (N_11145,N_7032,N_6786);
nand U11146 (N_11146,N_8185,N_7976);
nand U11147 (N_11147,N_6767,N_5768);
nand U11148 (N_11148,N_5720,N_7718);
or U11149 (N_11149,N_8346,N_8467);
nor U11150 (N_11150,N_8687,N_6393);
or U11151 (N_11151,N_8195,N_6177);
xor U11152 (N_11152,N_5793,N_7791);
xor U11153 (N_11153,N_7538,N_6942);
nand U11154 (N_11154,N_8336,N_9683);
nand U11155 (N_11155,N_7071,N_6261);
nor U11156 (N_11156,N_6271,N_9113);
and U11157 (N_11157,N_6398,N_7327);
nor U11158 (N_11158,N_5245,N_8680);
and U11159 (N_11159,N_7018,N_9730);
nor U11160 (N_11160,N_6210,N_5083);
and U11161 (N_11161,N_6916,N_5420);
nand U11162 (N_11162,N_5770,N_5644);
xor U11163 (N_11163,N_7467,N_9518);
nor U11164 (N_11164,N_6543,N_8436);
nand U11165 (N_11165,N_7001,N_5839);
xnor U11166 (N_11166,N_8004,N_9604);
or U11167 (N_11167,N_6306,N_5878);
or U11168 (N_11168,N_5769,N_5693);
xnor U11169 (N_11169,N_7812,N_5395);
and U11170 (N_11170,N_9477,N_8399);
and U11171 (N_11171,N_5310,N_8117);
or U11172 (N_11172,N_7326,N_6039);
nor U11173 (N_11173,N_5462,N_6151);
nor U11174 (N_11174,N_8332,N_8850);
or U11175 (N_11175,N_7657,N_8932);
and U11176 (N_11176,N_7658,N_5895);
nor U11177 (N_11177,N_9376,N_7416);
nor U11178 (N_11178,N_9635,N_6588);
and U11179 (N_11179,N_7041,N_7148);
and U11180 (N_11180,N_5057,N_6506);
and U11181 (N_11181,N_5763,N_9008);
and U11182 (N_11182,N_5926,N_9944);
and U11183 (N_11183,N_5829,N_9713);
nand U11184 (N_11184,N_9758,N_9508);
nand U11185 (N_11185,N_6130,N_8633);
and U11186 (N_11186,N_5647,N_9950);
or U11187 (N_11187,N_7397,N_7608);
or U11188 (N_11188,N_6750,N_5727);
and U11189 (N_11189,N_7056,N_7519);
xnor U11190 (N_11190,N_7525,N_9576);
nand U11191 (N_11191,N_9250,N_7881);
or U11192 (N_11192,N_8808,N_6980);
or U11193 (N_11193,N_8258,N_9759);
nand U11194 (N_11194,N_7797,N_5570);
or U11195 (N_11195,N_6551,N_8829);
nand U11196 (N_11196,N_8917,N_9260);
and U11197 (N_11197,N_8091,N_7437);
and U11198 (N_11198,N_7333,N_7632);
or U11199 (N_11199,N_8564,N_6171);
xnor U11200 (N_11200,N_7439,N_6193);
or U11201 (N_11201,N_5249,N_6038);
nor U11202 (N_11202,N_8726,N_7726);
xnor U11203 (N_11203,N_8182,N_8318);
and U11204 (N_11204,N_9249,N_9550);
nand U11205 (N_11205,N_5108,N_5551);
nor U11206 (N_11206,N_7550,N_7288);
and U11207 (N_11207,N_5804,N_5595);
nor U11208 (N_11208,N_7117,N_5116);
xor U11209 (N_11209,N_8411,N_5580);
nand U11210 (N_11210,N_7652,N_7813);
and U11211 (N_11211,N_9411,N_5047);
nand U11212 (N_11212,N_7855,N_9865);
nor U11213 (N_11213,N_7081,N_7284);
nand U11214 (N_11214,N_5935,N_8186);
xor U11215 (N_11215,N_7938,N_8915);
nand U11216 (N_11216,N_6866,N_5944);
or U11217 (N_11217,N_6118,N_5439);
and U11218 (N_11218,N_8652,N_8342);
xnor U11219 (N_11219,N_6379,N_7356);
nand U11220 (N_11220,N_9831,N_8747);
or U11221 (N_11221,N_6215,N_6544);
nor U11222 (N_11222,N_6804,N_8419);
and U11223 (N_11223,N_9321,N_7751);
nand U11224 (N_11224,N_7631,N_8037);
nand U11225 (N_11225,N_9811,N_6176);
and U11226 (N_11226,N_7854,N_5671);
and U11227 (N_11227,N_7970,N_8500);
and U11228 (N_11228,N_8590,N_7479);
and U11229 (N_11229,N_5674,N_5373);
and U11230 (N_11230,N_6887,N_5767);
nor U11231 (N_11231,N_9735,N_9274);
nor U11232 (N_11232,N_9131,N_6276);
nand U11233 (N_11233,N_6719,N_8794);
or U11234 (N_11234,N_8283,N_9149);
or U11235 (N_11235,N_8382,N_6449);
and U11236 (N_11236,N_9506,N_9602);
xor U11237 (N_11237,N_8226,N_6813);
nor U11238 (N_11238,N_6712,N_6301);
and U11239 (N_11239,N_8409,N_9905);
or U11240 (N_11240,N_8525,N_9138);
nand U11241 (N_11241,N_7127,N_7624);
or U11242 (N_11242,N_7180,N_5102);
nand U11243 (N_11243,N_6991,N_7234);
nand U11244 (N_11244,N_8005,N_5985);
or U11245 (N_11245,N_9173,N_5196);
and U11246 (N_11246,N_7828,N_5231);
nand U11247 (N_11247,N_5699,N_7296);
nand U11248 (N_11248,N_7775,N_9100);
nand U11249 (N_11249,N_9877,N_7877);
nor U11250 (N_11250,N_6869,N_9961);
nand U11251 (N_11251,N_6072,N_6368);
or U11252 (N_11252,N_5542,N_7095);
xor U11253 (N_11253,N_5271,N_8948);
and U11254 (N_11254,N_6598,N_8454);
nor U11255 (N_11255,N_9981,N_9242);
nand U11256 (N_11256,N_5019,N_6652);
or U11257 (N_11257,N_8485,N_9120);
nand U11258 (N_11258,N_8793,N_6404);
xnor U11259 (N_11259,N_8072,N_5223);
or U11260 (N_11260,N_8204,N_5918);
nor U11261 (N_11261,N_9027,N_9355);
and U11262 (N_11262,N_8838,N_6944);
and U11263 (N_11263,N_7182,N_6243);
nor U11264 (N_11264,N_7809,N_9041);
nand U11265 (N_11265,N_5272,N_7008);
nand U11266 (N_11266,N_6616,N_7783);
or U11267 (N_11267,N_6629,N_5247);
nand U11268 (N_11268,N_6337,N_7974);
and U11269 (N_11269,N_9917,N_7805);
nand U11270 (N_11270,N_5266,N_9424);
and U11271 (N_11271,N_8249,N_7223);
nand U11272 (N_11272,N_9316,N_9441);
and U11273 (N_11273,N_5519,N_9042);
nand U11274 (N_11274,N_7432,N_8624);
nor U11275 (N_11275,N_9642,N_5274);
nor U11276 (N_11276,N_7888,N_7827);
nor U11277 (N_11277,N_6091,N_7131);
nor U11278 (N_11278,N_8376,N_8800);
or U11279 (N_11279,N_9664,N_9114);
and U11280 (N_11280,N_7531,N_7713);
and U11281 (N_11281,N_9466,N_8844);
and U11282 (N_11282,N_5422,N_6254);
nand U11283 (N_11283,N_6416,N_7691);
xor U11284 (N_11284,N_7561,N_5649);
or U11285 (N_11285,N_6355,N_5883);
nand U11286 (N_11286,N_8583,N_9102);
nand U11287 (N_11287,N_8790,N_6647);
nand U11288 (N_11288,N_8448,N_9259);
or U11289 (N_11289,N_9370,N_9417);
nor U11290 (N_11290,N_7607,N_5850);
xnor U11291 (N_11291,N_9081,N_5556);
nor U11292 (N_11292,N_7516,N_7414);
nand U11293 (N_11293,N_6429,N_6043);
nand U11294 (N_11294,N_8125,N_8773);
xor U11295 (N_11295,N_5330,N_8770);
nor U11296 (N_11296,N_7873,N_5642);
or U11297 (N_11297,N_7810,N_7134);
xnor U11298 (N_11298,N_5638,N_8388);
xnor U11299 (N_11299,N_5730,N_6492);
nand U11300 (N_11300,N_5976,N_5765);
nand U11301 (N_11301,N_9408,N_5472);
nor U11302 (N_11302,N_6417,N_5298);
nand U11303 (N_11303,N_9847,N_7689);
and U11304 (N_11304,N_7404,N_7492);
nand U11305 (N_11305,N_7065,N_9866);
nor U11306 (N_11306,N_9435,N_7339);
nand U11307 (N_11307,N_8512,N_6428);
or U11308 (N_11308,N_7279,N_8804);
or U11309 (N_11309,N_8660,N_6159);
nor U11310 (N_11310,N_5037,N_5107);
nand U11311 (N_11311,N_9229,N_7801);
nor U11312 (N_11312,N_8609,N_6762);
nor U11313 (N_11313,N_9044,N_8444);
xor U11314 (N_11314,N_6918,N_5596);
nor U11315 (N_11315,N_9052,N_5094);
nand U11316 (N_11316,N_9740,N_8413);
nand U11317 (N_11317,N_8866,N_8180);
or U11318 (N_11318,N_8297,N_7665);
nor U11319 (N_11319,N_8307,N_5197);
nand U11320 (N_11320,N_5664,N_8570);
xnor U11321 (N_11321,N_8468,N_5276);
nor U11322 (N_11322,N_8049,N_5799);
xnor U11323 (N_11323,N_6317,N_8894);
xor U11324 (N_11324,N_9808,N_6251);
and U11325 (N_11325,N_7901,N_9887);
or U11326 (N_11326,N_5312,N_7541);
nand U11327 (N_11327,N_5898,N_9142);
or U11328 (N_11328,N_7393,N_7370);
and U11329 (N_11329,N_8791,N_6297);
or U11330 (N_11330,N_6055,N_5737);
xnor U11331 (N_11331,N_6075,N_5017);
nand U11332 (N_11332,N_9495,N_6219);
or U11333 (N_11333,N_9169,N_5009);
and U11334 (N_11334,N_9751,N_8931);
nor U11335 (N_11335,N_8469,N_9013);
and U11336 (N_11336,N_8344,N_6191);
and U11337 (N_11337,N_6517,N_8035);
xnor U11338 (N_11338,N_5412,N_8031);
nand U11339 (N_11339,N_8777,N_9584);
and U11340 (N_11340,N_7030,N_5135);
and U11341 (N_11341,N_9716,N_8882);
or U11342 (N_11342,N_8028,N_8158);
nand U11343 (N_11343,N_5518,N_9755);
nand U11344 (N_11344,N_9492,N_9154);
nor U11345 (N_11345,N_6720,N_8762);
nand U11346 (N_11346,N_7836,N_7826);
nor U11347 (N_11347,N_9257,N_8597);
nor U11348 (N_11348,N_7491,N_5068);
nor U11349 (N_11349,N_6609,N_5499);
or U11350 (N_11350,N_7342,N_7027);
and U11351 (N_11351,N_9834,N_9022);
or U11352 (N_11352,N_7456,N_5957);
or U11353 (N_11353,N_5242,N_8009);
nand U11354 (N_11354,N_9967,N_5875);
nand U11355 (N_11355,N_8952,N_6618);
xnor U11356 (N_11356,N_9938,N_6841);
nor U11357 (N_11357,N_8327,N_9475);
nor U11358 (N_11358,N_5701,N_7999);
nor U11359 (N_11359,N_5687,N_6654);
or U11360 (N_11360,N_5721,N_9245);
or U11361 (N_11361,N_9841,N_7727);
nand U11362 (N_11362,N_5491,N_5815);
and U11363 (N_11363,N_6345,N_6765);
or U11364 (N_11364,N_6120,N_8495);
or U11365 (N_11365,N_7930,N_7238);
or U11366 (N_11366,N_7077,N_7380);
nand U11367 (N_11367,N_5316,N_9419);
nor U11368 (N_11368,N_7528,N_8923);
and U11369 (N_11369,N_6939,N_6861);
and U11370 (N_11370,N_6574,N_5071);
nor U11371 (N_11371,N_6729,N_6152);
nor U11372 (N_11372,N_8383,N_8476);
and U11373 (N_11373,N_7629,N_7839);
xor U11374 (N_11374,N_7281,N_9314);
or U11375 (N_11375,N_7513,N_9480);
nor U11376 (N_11376,N_5907,N_6746);
xnor U11377 (N_11377,N_8513,N_8353);
nor U11378 (N_11378,N_9913,N_6951);
nor U11379 (N_11379,N_7678,N_7066);
nor U11380 (N_11380,N_7966,N_6548);
nor U11381 (N_11381,N_6894,N_6205);
and U11382 (N_11382,N_7832,N_7330);
nor U11383 (N_11383,N_6410,N_5483);
xnor U11384 (N_11384,N_6604,N_9999);
or U11385 (N_11385,N_7709,N_8571);
nand U11386 (N_11386,N_8646,N_9165);
and U11387 (N_11387,N_9083,N_7031);
or U11388 (N_11388,N_8968,N_5581);
nor U11389 (N_11389,N_6467,N_7639);
and U11390 (N_11390,N_9496,N_7443);
nor U11391 (N_11391,N_7046,N_6922);
and U11392 (N_11392,N_6270,N_6325);
nand U11393 (N_11393,N_8976,N_8568);
nand U11394 (N_11394,N_6934,N_5171);
nor U11395 (N_11395,N_5739,N_6535);
xnor U11396 (N_11396,N_8748,N_7707);
nor U11397 (N_11397,N_5736,N_5117);
nor U11398 (N_11398,N_7603,N_6170);
nand U11399 (N_11399,N_8395,N_7649);
nor U11400 (N_11400,N_9956,N_5974);
or U11401 (N_11401,N_7278,N_5156);
nor U11402 (N_11402,N_5990,N_7627);
and U11403 (N_11403,N_6630,N_5304);
and U11404 (N_11404,N_8598,N_6050);
nand U11405 (N_11405,N_5323,N_9869);
nor U11406 (N_11406,N_7496,N_5539);
or U11407 (N_11407,N_7136,N_7741);
nand U11408 (N_11408,N_6791,N_5279);
and U11409 (N_11409,N_9430,N_5157);
and U11410 (N_11410,N_9977,N_8074);
or U11411 (N_11411,N_8325,N_7315);
nor U11412 (N_11412,N_9731,N_8164);
and U11413 (N_11413,N_6051,N_9728);
nor U11414 (N_11414,N_5797,N_7656);
nor U11415 (N_11415,N_9675,N_5814);
xor U11416 (N_11416,N_9587,N_5407);
nand U11417 (N_11417,N_9784,N_6648);
nor U11418 (N_11418,N_8820,N_8102);
nor U11419 (N_11419,N_5656,N_9098);
nand U11420 (N_11420,N_6183,N_9069);
nor U11421 (N_11421,N_7529,N_7305);
or U11422 (N_11422,N_6623,N_5262);
or U11423 (N_11423,N_8942,N_9684);
nor U11424 (N_11424,N_8151,N_9774);
xnor U11425 (N_11425,N_9941,N_7571);
xor U11426 (N_11426,N_5544,N_9467);
and U11427 (N_11427,N_7874,N_9543);
and U11428 (N_11428,N_9318,N_5065);
nor U11429 (N_11429,N_7213,N_7676);
xnor U11430 (N_11430,N_7196,N_8958);
nand U11431 (N_11431,N_7286,N_9166);
nand U11432 (N_11432,N_5128,N_7232);
or U11433 (N_11433,N_5444,N_7753);
and U11434 (N_11434,N_5713,N_7523);
and U11435 (N_11435,N_5020,N_6356);
nor U11436 (N_11436,N_8935,N_7876);
nor U11437 (N_11437,N_8152,N_5093);
or U11438 (N_11438,N_9782,N_5597);
and U11439 (N_11439,N_9722,N_8661);
nor U11440 (N_11440,N_8809,N_9812);
or U11441 (N_11441,N_6706,N_5854);
and U11442 (N_11442,N_7149,N_6422);
or U11443 (N_11443,N_6589,N_6148);
and U11444 (N_11444,N_8771,N_7536);
nand U11445 (N_11445,N_7673,N_7621);
or U11446 (N_11446,N_9225,N_6620);
nor U11447 (N_11447,N_5745,N_9360);
nor U11448 (N_11448,N_6026,N_7651);
or U11449 (N_11449,N_5650,N_7300);
nor U11450 (N_11450,N_9849,N_5146);
nand U11451 (N_11451,N_8752,N_8728);
or U11452 (N_11452,N_8539,N_7361);
nand U11453 (N_11453,N_5906,N_9134);
nor U11454 (N_11454,N_9464,N_9244);
nand U11455 (N_11455,N_6565,N_8089);
nand U11456 (N_11456,N_9415,N_5966);
xor U11457 (N_11457,N_8365,N_6086);
nor U11458 (N_11458,N_8832,N_6768);
xnor U11459 (N_11459,N_9671,N_6882);
nor U11460 (N_11460,N_5707,N_8259);
or U11461 (N_11461,N_6178,N_5987);
nand U11462 (N_11462,N_9539,N_5179);
or U11463 (N_11463,N_7610,N_8366);
or U11464 (N_11464,N_6443,N_5525);
nor U11465 (N_11465,N_5147,N_7205);
nand U11466 (N_11466,N_8021,N_7160);
nor U11467 (N_11467,N_7154,N_6724);
and U11468 (N_11468,N_8390,N_7696);
nor U11469 (N_11469,N_6298,N_5113);
nor U11470 (N_11470,N_6992,N_8611);
and U11471 (N_11471,N_5812,N_5756);
xor U11472 (N_11472,N_7702,N_9246);
or U11473 (N_11473,N_9512,N_7038);
nand U11474 (N_11474,N_9872,N_6189);
nand U11475 (N_11475,N_9350,N_9546);
nand U11476 (N_11476,N_6119,N_8560);
nor U11477 (N_11477,N_7021,N_6925);
nor U11478 (N_11478,N_6439,N_7480);
nand U11479 (N_11479,N_5306,N_9359);
nor U11480 (N_11480,N_8559,N_8282);
or U11481 (N_11481,N_8176,N_6115);
xor U11482 (N_11482,N_8105,N_9132);
and U11483 (N_11483,N_9661,N_5458);
nor U11484 (N_11484,N_8591,N_6400);
nand U11485 (N_11485,N_8919,N_5722);
nor U11486 (N_11486,N_8046,N_8596);
and U11487 (N_11487,N_6174,N_8367);
or U11488 (N_11488,N_7577,N_9552);
and U11489 (N_11489,N_5187,N_7107);
and U11490 (N_11490,N_5115,N_7217);
nand U11491 (N_11491,N_5734,N_8015);
nor U11492 (N_11492,N_8579,N_8375);
and U11493 (N_11493,N_9179,N_5916);
and U11494 (N_11494,N_9598,N_8123);
and U11495 (N_11495,N_6462,N_7952);
nor U11496 (N_11496,N_6622,N_5994);
and U11497 (N_11497,N_9174,N_8404);
nand U11498 (N_11498,N_9485,N_8487);
or U11499 (N_11499,N_6161,N_8841);
nor U11500 (N_11500,N_7052,N_8128);
and U11501 (N_11501,N_6626,N_8144);
and U11502 (N_11502,N_8551,N_7803);
and U11503 (N_11503,N_7780,N_5531);
or U11504 (N_11504,N_7844,N_6472);
nand U11505 (N_11505,N_8427,N_5321);
nand U11506 (N_11506,N_6153,N_6494);
nand U11507 (N_11507,N_6823,N_8517);
and U11508 (N_11508,N_6246,N_6245);
nand U11509 (N_11509,N_8860,N_9397);
nor U11510 (N_11510,N_7641,N_8746);
nand U11511 (N_11511,N_5455,N_7622);
nor U11512 (N_11512,N_9971,N_9186);
xnor U11513 (N_11513,N_6007,N_8193);
nor U11514 (N_11514,N_8434,N_6656);
nor U11515 (N_11515,N_9404,N_9853);
xor U11516 (N_11516,N_5774,N_6591);
or U11517 (N_11517,N_8768,N_8095);
nand U11518 (N_11518,N_8909,N_7650);
nand U11519 (N_11519,N_9819,N_8481);
and U11520 (N_11520,N_7385,N_5980);
and U11521 (N_11521,N_9571,N_5828);
or U11522 (N_11522,N_6566,N_7732);
and U11523 (N_11523,N_9358,N_5466);
and U11524 (N_11524,N_8422,N_7563);
nand U11525 (N_11525,N_8823,N_6525);
or U11526 (N_11526,N_6362,N_5036);
nand U11527 (N_11527,N_5970,N_8802);
xor U11528 (N_11528,N_5145,N_8502);
and U11529 (N_11529,N_5696,N_5121);
nand U11530 (N_11530,N_7900,N_9659);
nor U11531 (N_11531,N_8608,N_9241);
xor U11532 (N_11532,N_6973,N_6670);
nor U11533 (N_11533,N_7929,N_5426);
nand U11534 (N_11534,N_8971,N_9555);
nand U11535 (N_11535,N_8545,N_6485);
nand U11536 (N_11536,N_9488,N_8993);
xnor U11537 (N_11537,N_6836,N_9313);
and U11538 (N_11538,N_8855,N_9793);
xnor U11539 (N_11539,N_8373,N_8106);
or U11540 (N_11540,N_6433,N_5760);
and U11541 (N_11541,N_7483,N_6957);
nor U11542 (N_11542,N_9459,N_6226);
and U11543 (N_11543,N_5158,N_8082);
nand U11544 (N_11544,N_7729,N_5033);
nor U11545 (N_11545,N_5761,N_9072);
or U11546 (N_11546,N_9608,N_5511);
nor U11547 (N_11547,N_9311,N_8536);
nor U11548 (N_11548,N_9644,N_6773);
and U11549 (N_11549,N_8431,N_8477);
nor U11550 (N_11550,N_9227,N_7353);
nand U11551 (N_11551,N_7814,N_7159);
nand U11552 (N_11552,N_5050,N_6381);
or U11553 (N_11553,N_9348,N_6902);
and U11554 (N_11554,N_9278,N_5216);
nor U11555 (N_11555,N_5110,N_9544);
nor U11556 (N_11556,N_8109,N_9507);
and U11557 (N_11557,N_9788,N_8418);
nor U11558 (N_11558,N_5295,N_5174);
nor U11559 (N_11559,N_5752,N_6761);
nor U11560 (N_11560,N_8441,N_7965);
or U11561 (N_11561,N_9378,N_6136);
nand U11562 (N_11562,N_7193,N_7386);
nor U11563 (N_11563,N_9075,N_6632);
or U11564 (N_11564,N_5259,N_5999);
nor U11565 (N_11565,N_7565,N_8087);
and U11566 (N_11566,N_9636,N_8406);
or U11567 (N_11567,N_8528,N_9176);
or U11568 (N_11568,N_8991,N_5154);
and U11569 (N_11569,N_7969,N_6853);
xnor U11570 (N_11570,N_6044,N_7229);
and U11571 (N_11571,N_7169,N_7941);
or U11572 (N_11572,N_5257,N_8149);
nor U11573 (N_11573,N_7880,N_5832);
nor U11574 (N_11574,N_8896,N_6639);
and U11575 (N_11575,N_9323,N_6870);
or U11576 (N_11576,N_9861,N_8006);
nor U11577 (N_11577,N_7364,N_5543);
nor U11578 (N_11578,N_7993,N_8738);
or U11579 (N_11579,N_5776,N_7909);
or U11580 (N_11580,N_6235,N_7706);
nor U11581 (N_11581,N_6446,N_5221);
nor U11582 (N_11582,N_5404,N_7944);
or U11583 (N_11583,N_9373,N_7913);
nand U11584 (N_11584,N_5501,N_8017);
xnor U11585 (N_11585,N_5344,N_5843);
or U11586 (N_11586,N_7125,N_9055);
nor U11587 (N_11587,N_6388,N_7493);
nor U11588 (N_11588,N_9678,N_8104);
nand U11589 (N_11589,N_7926,N_9504);
or U11590 (N_11590,N_8298,N_9338);
and U11591 (N_11591,N_7578,N_9897);
nand U11592 (N_11592,N_7301,N_8781);
nand U11593 (N_11593,N_6213,N_9181);
nor U11594 (N_11594,N_8238,N_9390);
and U11595 (N_11595,N_5624,N_5398);
nand U11596 (N_11596,N_5872,N_7161);
nand U11597 (N_11597,N_9294,N_6460);
nand U11598 (N_11598,N_6285,N_6617);
nor U11599 (N_11599,N_6917,N_8831);
xnor U11600 (N_11600,N_9096,N_7879);
and U11601 (N_11601,N_8224,N_7768);
or U11602 (N_11602,N_5396,N_9595);
and U11603 (N_11603,N_7190,N_8228);
xor U11604 (N_11604,N_7587,N_5949);
nand U11605 (N_11605,N_5096,N_9195);
nand U11606 (N_11606,N_8212,N_5495);
and U11607 (N_11607,N_8402,N_6976);
nand U11608 (N_11608,N_8638,N_5827);
or U11609 (N_11609,N_9324,N_5626);
and U11610 (N_11610,N_5984,N_6122);
xnor U11611 (N_11611,N_5532,N_7770);
or U11612 (N_11612,N_9911,N_9693);
or U11613 (N_11613,N_9770,N_5661);
or U11614 (N_11614,N_8816,N_6216);
or U11615 (N_11615,N_5849,N_7507);
xor U11616 (N_11616,N_5322,N_7645);
nand U11617 (N_11617,N_5289,N_9585);
and U11618 (N_11618,N_9914,N_6365);
nor U11619 (N_11619,N_7012,N_9447);
or U11620 (N_11620,N_9298,N_9036);
and U11621 (N_11621,N_8985,N_5683);
or U11622 (N_11622,N_8223,N_9520);
and U11623 (N_11623,N_7616,N_5007);
and U11624 (N_11624,N_9736,N_7685);
nand U11625 (N_11625,N_7829,N_9185);
nand U11626 (N_11626,N_6262,N_7323);
or U11627 (N_11627,N_7458,N_6522);
xnor U11628 (N_11628,N_6093,N_8879);
nand U11629 (N_11629,N_6843,N_8695);
nor U11630 (N_11630,N_7526,N_7530);
nor U11631 (N_11631,N_7784,N_6790);
nand U11632 (N_11632,N_7471,N_6437);
nand U11633 (N_11633,N_7668,N_5371);
nand U11634 (N_11634,N_8331,N_7017);
nand U11635 (N_11635,N_6158,N_6772);
or U11636 (N_11636,N_6615,N_9665);
xnor U11637 (N_11637,N_9346,N_8867);
or U11638 (N_11638,N_9379,N_9356);
xnor U11639 (N_11639,N_9045,N_6714);
or U11640 (N_11640,N_5562,N_5489);
xnor U11641 (N_11641,N_9842,N_6269);
and U11642 (N_11642,N_6127,N_5090);
nand U11643 (N_11643,N_7759,N_6847);
or U11644 (N_11644,N_8966,N_5087);
nor U11645 (N_11645,N_7002,N_8792);
xnor U11646 (N_11646,N_8263,N_9453);
nor U11647 (N_11647,N_5630,N_9091);
nor U11648 (N_11648,N_5802,N_6930);
or U11649 (N_11649,N_7322,N_8873);
nand U11650 (N_11650,N_5002,N_6640);
or U11651 (N_11651,N_5946,N_9410);
or U11652 (N_11652,N_8730,N_8296);
nor U11653 (N_11653,N_6781,N_7635);
or U11654 (N_11654,N_7150,N_5484);
nor U11655 (N_11655,N_9698,N_7007);
nand U11656 (N_11656,N_7336,N_8727);
and U11657 (N_11657,N_5564,N_6084);
and U11658 (N_11658,N_9802,N_9899);
nand U11659 (N_11659,N_8098,N_6967);
nand U11660 (N_11660,N_5446,N_7405);
nor U11661 (N_11661,N_8042,N_6530);
nand U11662 (N_11662,N_5457,N_8235);
or U11663 (N_11663,N_7082,N_6008);
or U11664 (N_11664,N_5986,N_7916);
nor U11665 (N_11665,N_9216,N_5783);
xnor U11666 (N_11666,N_8758,N_5704);
nor U11667 (N_11667,N_8507,N_9614);
nand U11668 (N_11668,N_6137,N_5195);
nand U11669 (N_11669,N_5868,N_7088);
nor U11670 (N_11670,N_6534,N_8863);
or U11671 (N_11671,N_6997,N_6694);
or U11672 (N_11672,N_8847,N_9933);
nor U11673 (N_11673,N_9606,N_8172);
or U11674 (N_11674,N_8392,N_5136);
or U11675 (N_11675,N_7725,N_9652);
nor U11676 (N_11676,N_9915,N_8601);
or U11677 (N_11677,N_5967,N_7478);
xnor U11678 (N_11678,N_5860,N_7455);
or U11679 (N_11679,N_6214,N_8414);
or U11680 (N_11680,N_7440,N_5277);
nor U11681 (N_11681,N_6481,N_6296);
or U11682 (N_11682,N_5937,N_8876);
and U11683 (N_11683,N_5268,N_7984);
nand U11684 (N_11684,N_8034,N_7547);
nor U11685 (N_11685,N_7100,N_6128);
and U11686 (N_11686,N_7747,N_9701);
nand U11687 (N_11687,N_8905,N_8721);
nand U11688 (N_11688,N_8301,N_7179);
nor U11689 (N_11689,N_7039,N_5026);
xor U11690 (N_11690,N_5545,N_5013);
nand U11691 (N_11691,N_5662,N_7378);
nor U11692 (N_11692,N_6921,N_9239);
or U11693 (N_11693,N_8013,N_8043);
and U11694 (N_11694,N_8688,N_8666);
nor U11695 (N_11695,N_8474,N_8615);
xor U11696 (N_11696,N_6661,N_7997);
nor U11697 (N_11697,N_6468,N_5386);
nand U11698 (N_11698,N_9337,N_8891);
nor U11699 (N_11699,N_7951,N_9115);
nand U11700 (N_11700,N_8269,N_8407);
and U11701 (N_11701,N_9486,N_5604);
and U11702 (N_11702,N_8933,N_8788);
or U11703 (N_11703,N_5400,N_5358);
and U11704 (N_11704,N_5445,N_8702);
and U11705 (N_11705,N_6448,N_6131);
nand U11706 (N_11706,N_9422,N_9384);
or U11707 (N_11707,N_5751,N_7101);
and U11708 (N_11708,N_5493,N_7990);
nor U11709 (N_11709,N_5526,N_7677);
and U11710 (N_11710,N_6139,N_9279);
nor U11711 (N_11711,N_6914,N_9112);
or U11712 (N_11712,N_7786,N_5175);
or U11713 (N_11713,N_5968,N_9369);
nor U11714 (N_11714,N_7474,N_6815);
nand U11715 (N_11715,N_5351,N_8705);
and U11716 (N_11716,N_6496,N_5778);
nand U11717 (N_11717,N_5379,N_7743);
nand U11718 (N_11718,N_5206,N_9118);
and U11719 (N_11719,N_8085,N_5855);
or U11720 (N_11720,N_6371,N_6476);
nand U11721 (N_11721,N_6883,N_6307);
or U11722 (N_11722,N_6856,N_6451);
and U11723 (N_11723,N_9304,N_5548);
nand U11724 (N_11724,N_5023,N_5943);
nor U11725 (N_11725,N_6288,N_5338);
and U11726 (N_11726,N_8300,N_5628);
nand U11727 (N_11727,N_6612,N_6402);
nand U11728 (N_11728,N_8603,N_6082);
nor U11729 (N_11729,N_5193,N_6165);
xnor U11730 (N_11730,N_7462,N_5517);
and U11731 (N_11731,N_6438,N_9046);
nand U11732 (N_11732,N_9513,N_5410);
and U11733 (N_11733,N_9943,N_9739);
nand U11734 (N_11734,N_8612,N_9054);
or U11735 (N_11735,N_7375,N_8464);
nor U11736 (N_11736,N_5328,N_7614);
and U11737 (N_11737,N_9023,N_6450);
xnor U11738 (N_11738,N_6359,N_9306);
nand U11739 (N_11739,N_8445,N_6204);
nand U11740 (N_11740,N_6667,N_9128);
and U11741 (N_11741,N_7570,N_7793);
or U11742 (N_11742,N_9645,N_6845);
or U11743 (N_11743,N_8874,N_8851);
nand U11744 (N_11744,N_6844,N_5964);
nor U11745 (N_11745,N_7501,N_6827);
or U11746 (N_11746,N_6718,N_8940);
nor U11747 (N_11747,N_7572,N_7138);
or U11748 (N_11748,N_5337,N_9493);
xor U11749 (N_11749,N_9786,N_5461);
nand U11750 (N_11750,N_5082,N_5308);
nor U11751 (N_11751,N_5027,N_9763);
or U11752 (N_11752,N_5982,N_7868);
nand U11753 (N_11753,N_8052,N_5670);
xnor U11754 (N_11754,N_6642,N_8019);
nor U11755 (N_11755,N_7442,N_6206);
xnor U11756 (N_11756,N_9948,N_5390);
nor U11757 (N_11757,N_9667,N_7484);
or U11758 (N_11758,N_7351,N_6376);
nand U11759 (N_11759,N_5258,N_5712);
nor U11760 (N_11760,N_8516,N_7348);
or U11761 (N_11761,N_6123,N_8602);
nand U11762 (N_11762,N_7834,N_8145);
xor U11763 (N_11763,N_5820,N_8011);
nor U11764 (N_11764,N_8207,N_5048);
and U11765 (N_11765,N_8575,N_8892);
nor U11766 (N_11766,N_6807,N_6763);
nand U11767 (N_11767,N_8644,N_9200);
and U11768 (N_11768,N_5637,N_5521);
and U11769 (N_11769,N_7521,N_9035);
and U11770 (N_11770,N_6370,N_7511);
nand U11771 (N_11771,N_5385,N_7118);
nor U11772 (N_11772,N_7429,N_7441);
xnor U11773 (N_11773,N_5678,N_5120);
nand U11774 (N_11774,N_9015,N_6290);
nand U11775 (N_11775,N_9018,N_7928);
nand U11776 (N_11776,N_8556,N_8555);
or U11777 (N_11777,N_6730,N_5339);
or U11778 (N_11778,N_6482,N_6657);
or U11779 (N_11779,N_8558,N_6795);
nor U11780 (N_11780,N_5923,N_5189);
or U11781 (N_11781,N_7549,N_7520);
nand U11782 (N_11782,N_5425,N_6469);
nor U11783 (N_11783,N_6256,N_5648);
or U11784 (N_11784,N_5622,N_9394);
and U11785 (N_11785,N_9843,N_5663);
or U11786 (N_11786,N_9434,N_8003);
nor U11787 (N_11787,N_8668,N_5781);
and U11788 (N_11788,N_5255,N_6088);
nor U11789 (N_11789,N_8814,N_8634);
and U11790 (N_11790,N_9299,N_9617);
or U11791 (N_11791,N_8693,N_8979);
and U11792 (N_11792,N_9280,N_8071);
nor U11793 (N_11793,N_5035,N_8432);
or U11794 (N_11794,N_9556,N_9816);
and U11795 (N_11795,N_7846,N_5972);
and U11796 (N_11796,N_5694,N_7173);
and U11797 (N_11797,N_7158,N_8050);
and U11798 (N_11798,N_9218,N_9037);
and U11799 (N_11799,N_5238,N_5494);
nand U11800 (N_11800,N_9212,N_6406);
and U11801 (N_11801,N_6837,N_8122);
and U11802 (N_11802,N_7398,N_8341);
nor U11803 (N_11803,N_5269,N_6770);
nand U11804 (N_11804,N_7730,N_9868);
nor U11805 (N_11805,N_7103,N_8287);
nor U11806 (N_11806,N_8654,N_8716);
nand U11807 (N_11807,N_6293,N_9777);
nor U11808 (N_11808,N_7807,N_6228);
and U11809 (N_11809,N_9732,N_5415);
or U11810 (N_11810,N_7750,N_5114);
and U11811 (N_11811,N_9193,N_8063);
and U11812 (N_11812,N_6755,N_6909);
xnor U11813 (N_11813,N_8048,N_8970);
nor U11814 (N_11814,N_6028,N_7698);
nand U11815 (N_11815,N_9547,N_5131);
nor U11816 (N_11816,N_6988,N_8605);
or U11817 (N_11817,N_8997,N_6435);
nand U11818 (N_11818,N_9708,N_8999);
nand U11819 (N_11819,N_5641,N_5862);
and U11820 (N_11820,N_5073,N_5530);
nor U11821 (N_11821,N_9669,N_9024);
and U11822 (N_11822,N_5356,N_9523);
nand U11823 (N_11823,N_5056,N_6489);
xor U11824 (N_11824,N_8625,N_6445);
nand U11825 (N_11825,N_9265,N_5554);
or U11826 (N_11826,N_7269,N_9860);
nand U11827 (N_11827,N_5049,N_6956);
nand U11828 (N_11828,N_7749,N_8047);
xor U11829 (N_11829,N_8206,N_9498);
nand U11830 (N_11830,N_5726,N_8191);
nor U11831 (N_11831,N_5354,N_9787);
and U11832 (N_11832,N_5211,N_8016);
and U11833 (N_11833,N_5372,N_9753);
nand U11834 (N_11834,N_8077,N_6850);
or U11835 (N_11835,N_6985,N_9827);
or U11836 (N_11836,N_8755,N_6281);
nor U11837 (N_11837,N_5884,N_6753);
and U11838 (N_11838,N_5565,N_5507);
or U11839 (N_11839,N_8064,N_5522);
xor U11840 (N_11840,N_9231,N_7053);
or U11841 (N_11841,N_5549,N_7882);
or U11842 (N_11842,N_6611,N_9451);
nand U11843 (N_11843,N_8267,N_6573);
and U11844 (N_11844,N_7774,N_6633);
and U11845 (N_11845,N_9979,N_5209);
or U11846 (N_11846,N_5821,N_6800);
nor U11847 (N_11847,N_5573,N_7776);
nand U11848 (N_11848,N_8732,N_9070);
xor U11849 (N_11849,N_5958,N_8099);
nand U11850 (N_11850,N_6064,N_6805);
and U11851 (N_11851,N_8797,N_5315);
xor U11852 (N_11852,N_5840,N_9125);
and U11853 (N_11853,N_7359,N_5905);
nand U11854 (N_11854,N_8202,N_6372);
and U11855 (N_11855,N_8503,N_8902);
or U11856 (N_11856,N_5796,N_6569);
or U11857 (N_11857,N_5391,N_7542);
and U11858 (N_11858,N_7128,N_9820);
or U11859 (N_11859,N_5088,N_8957);
and U11860 (N_11860,N_9640,N_8714);
or U11861 (N_11861,N_5877,N_6239);
xor U11862 (N_11862,N_6751,N_7978);
and U11863 (N_11863,N_6194,N_7447);
nand U11864 (N_11864,N_6273,N_6913);
nor U11865 (N_11865,N_7060,N_9626);
and U11866 (N_11866,N_5475,N_9005);
nand U11867 (N_11867,N_5806,N_5465);
nand U11868 (N_11868,N_8967,N_9519);
or U11869 (N_11869,N_6567,N_5709);
and U11870 (N_11870,N_7428,N_5467);
xnor U11871 (N_11871,N_8822,N_9864);
or U11872 (N_11872,N_9322,N_6961);
and U11873 (N_11873,N_7421,N_7465);
nand U11874 (N_11874,N_8372,N_7155);
nor U11875 (N_11875,N_9591,N_8170);
or U11876 (N_11876,N_8614,N_7856);
nand U11877 (N_11877,N_6248,N_7352);
nand U11878 (N_11878,N_9781,N_9445);
nand U11879 (N_11879,N_6716,N_7708);
nand U11880 (N_11880,N_5889,N_6501);
or U11881 (N_11881,N_5614,N_8051);
nand U11882 (N_11882,N_7275,N_8766);
or U11883 (N_11883,N_8875,N_5403);
or U11884 (N_11884,N_6294,N_7446);
or U11885 (N_11885,N_5601,N_7074);
nor U11886 (N_11886,N_6783,N_5933);
or U11887 (N_11887,N_6006,N_9162);
nand U11888 (N_11888,N_7367,N_6005);
xor U11889 (N_11889,N_5303,N_8769);
nor U11890 (N_11890,N_8588,N_8796);
and U11891 (N_11891,N_9963,N_9053);
nor U11892 (N_11892,N_5237,N_6223);
and U11893 (N_11893,N_5629,N_7029);
nand U11894 (N_11894,N_7692,N_6974);
and U11895 (N_11895,N_6926,N_9383);
xor U11896 (N_11896,N_9692,N_7045);
nor U11897 (N_11897,N_7172,N_5229);
nand U11898 (N_11898,N_5932,N_7244);
nand U11899 (N_11899,N_5500,N_8586);
nor U11900 (N_11900,N_9829,N_6156);
nand U11901 (N_11901,N_7274,N_7950);
nand U11902 (N_11902,N_5627,N_5608);
or U11903 (N_11903,N_6140,N_7156);
and U11904 (N_11904,N_9533,N_6175);
nor U11905 (N_11905,N_5897,N_7518);
and U11906 (N_11906,N_7303,N_7062);
and U11907 (N_11907,N_9973,N_9065);
nand U11908 (N_11908,N_8607,N_5327);
nor U11909 (N_11909,N_5886,N_7609);
nor U11910 (N_11910,N_9272,N_8980);
and U11911 (N_11911,N_5585,N_5067);
nor U11912 (N_11912,N_9549,N_5773);
xor U11913 (N_11913,N_8394,N_8246);
nand U11914 (N_11914,N_6098,N_7435);
nand U11915 (N_11915,N_9421,N_7980);
nor U11916 (N_11916,N_7907,N_6466);
nand U11917 (N_11917,N_7737,N_9951);
nor U11918 (N_11918,N_6542,N_7091);
and U11919 (N_11919,N_7848,N_7047);
or U11920 (N_11920,N_6503,N_7972);
nor U11921 (N_11921,N_9922,N_9064);
nand U11922 (N_11922,N_9161,N_5301);
or U11923 (N_11923,N_6601,N_9454);
and U11924 (N_11924,N_5365,N_8675);
nor U11925 (N_11925,N_5346,N_8385);
or U11926 (N_11926,N_6110,N_7920);
nor U11927 (N_11927,N_8335,N_5488);
and U11928 (N_11928,N_7618,N_5890);
nand U11929 (N_11929,N_7630,N_5772);
nand U11930 (N_11930,N_8273,N_7710);
nand U11931 (N_11931,N_5540,N_7871);
and U11932 (N_11932,N_7625,N_8245);
or U11933 (N_11933,N_6068,N_9818);
or U11934 (N_11934,N_8265,N_6252);
or U11935 (N_11935,N_7260,N_9757);
xnor U11936 (N_11936,N_6928,N_6950);
nand U11937 (N_11937,N_7960,N_7408);
nand U11938 (N_11938,N_9302,N_6046);
nand U11939 (N_11939,N_6188,N_8628);
nor U11940 (N_11940,N_6389,N_9515);
xnor U11941 (N_11941,N_5950,N_9765);
nand U11942 (N_11942,N_6814,N_8348);
nor U11943 (N_11943,N_9937,N_7898);
nand U11944 (N_11944,N_6382,N_8211);
nand U11945 (N_11945,N_5011,N_8623);
or U11946 (N_11946,N_7316,N_9039);
or U11947 (N_11947,N_6935,N_6830);
or U11948 (N_11948,N_8700,N_9578);
and U11949 (N_11949,N_7451,N_6708);
or U11950 (N_11950,N_6164,N_6042);
xor U11951 (N_11951,N_7971,N_5865);
or U11952 (N_11952,N_9638,N_5192);
nand U11953 (N_11953,N_9630,N_5858);
or U11954 (N_11954,N_7738,N_8187);
or U11955 (N_11955,N_7290,N_8131);
and U11956 (N_11956,N_8456,N_6017);
nand U11957 (N_11957,N_7878,N_5015);
or U11958 (N_11958,N_9377,N_5867);
and U11959 (N_11959,N_6078,N_8739);
or U11960 (N_11960,N_7028,N_5253);
nand U11961 (N_11961,N_7943,N_9772);
or U11962 (N_11962,N_5996,N_7311);
or U11963 (N_11963,N_6735,N_5803);
nand U11964 (N_11964,N_7291,N_5044);
or U11965 (N_11965,N_8083,N_9449);
nand U11966 (N_11966,N_8116,N_6665);
nand U11967 (N_11967,N_8509,N_7896);
nand U11968 (N_11968,N_9969,N_5822);
and U11969 (N_11969,N_6263,N_9300);
and U11970 (N_11970,N_7240,N_5919);
xnor U11971 (N_11971,N_9637,N_6079);
nor U11972 (N_11972,N_6680,N_5902);
xnor U11973 (N_11973,N_6272,N_8229);
nor U11974 (N_11974,N_9395,N_5165);
and U11975 (N_11975,N_7033,N_9308);
or U11976 (N_11976,N_6707,N_7392);
nand U11977 (N_11977,N_8574,N_6267);
nor U11978 (N_11978,N_5440,N_9489);
and U11979 (N_11979,N_7083,N_6594);
nand U11980 (N_11980,N_6941,N_9393);
nor U11981 (N_11981,N_6577,N_9500);
xnor U11982 (N_11982,N_7660,N_9972);
or U11983 (N_11983,N_7895,N_6258);
and U11984 (N_11984,N_7162,N_9725);
nor U11985 (N_11985,N_6946,N_9334);
xor U11986 (N_11986,N_8442,N_9779);
xnor U11987 (N_11987,N_5920,N_6590);
or U11988 (N_11988,N_5076,N_8927);
or U11989 (N_11989,N_7551,N_6475);
or U11990 (N_11990,N_8674,N_6268);
or U11991 (N_11991,N_5317,N_6257);
nor U11992 (N_11992,N_8922,N_9752);
or U11993 (N_11993,N_7858,N_6892);
nor U11994 (N_11994,N_7403,N_6519);
nand U11995 (N_11995,N_7225,N_9838);
nand U11996 (N_11996,N_8849,N_8080);
nand U11997 (N_11997,N_5924,N_5290);
or U11998 (N_11998,N_7226,N_6754);
nor U11999 (N_11999,N_8492,N_7379);
nand U12000 (N_12000,N_8813,N_8240);
or U12001 (N_12001,N_9326,N_7961);
nor U12002 (N_12002,N_9674,N_7419);
and U12003 (N_12003,N_8148,N_7701);
or U12004 (N_12004,N_8054,N_7412);
nor U12005 (N_12005,N_5433,N_6948);
and U12006 (N_12006,N_5602,N_8722);
and U12007 (N_12007,N_8210,N_9600);
nor U12008 (N_12008,N_9858,N_6828);
nand U12009 (N_12009,N_9615,N_6994);
nor U12010 (N_12010,N_8642,N_5451);
nand U12011 (N_12011,N_8639,N_7647);
nor U12012 (N_12012,N_6554,N_6982);
nand U12013 (N_12013,N_9157,N_8965);
or U12014 (N_12014,N_6725,N_7872);
nand U12015 (N_12015,N_5089,N_5535);
nor U12016 (N_12016,N_6483,N_6582);
nor U12017 (N_12017,N_5502,N_6274);
or U12018 (N_12018,N_8397,N_5818);
or U12019 (N_12019,N_8521,N_8146);
and U12020 (N_12020,N_6114,N_8538);
xor U12021 (N_12021,N_8349,N_9030);
nand U12022 (N_12022,N_5069,N_7123);
or U12023 (N_12023,N_5042,N_7366);
xnor U12024 (N_12024,N_8292,N_8443);
nor U12025 (N_12025,N_9002,N_9958);
nand U12026 (N_12026,N_7598,N_5388);
or U12027 (N_12027,N_5176,N_9855);
nand U12028 (N_12028,N_8776,N_9891);
or U12029 (N_12029,N_5101,N_5881);
or U12030 (N_12030,N_9364,N_8581);
and U12031 (N_12031,N_7016,N_5945);
and U12032 (N_12032,N_5740,N_6277);
nor U12033 (N_12033,N_8262,N_9222);
and U12034 (N_12034,N_9767,N_5213);
nand U12035 (N_12035,N_6774,N_5000);
and U12036 (N_12036,N_9190,N_6286);
nand U12037 (N_12037,N_8622,N_6780);
or U12038 (N_12038,N_6339,N_5307);
and U12039 (N_12039,N_6486,N_9284);
and U12040 (N_12040,N_6796,N_5318);
nand U12041 (N_12041,N_9476,N_8743);
xnor U12042 (N_12042,N_5988,N_8401);
nand U12043 (N_12043,N_8658,N_7640);
nor U12044 (N_12044,N_5045,N_7568);
nor U12045 (N_12045,N_9724,N_6679);
nor U12046 (N_12046,N_7611,N_5555);
and U12047 (N_12047,N_5456,N_7025);
or U12048 (N_12048,N_7374,N_9372);
or U12049 (N_12049,N_5914,N_6782);
and U12050 (N_12050,N_8025,N_7596);
nand U12051 (N_12051,N_5450,N_5060);
nor U12052 (N_12052,N_7115,N_7270);
or U12053 (N_12053,N_8281,N_6125);
and U12054 (N_12054,N_8275,N_6312);
xor U12055 (N_12055,N_8709,N_9032);
nor U12056 (N_12056,N_5155,N_8027);
and U12057 (N_12057,N_9281,N_8843);
nor U12058 (N_12058,N_5870,N_5791);
xnor U12059 (N_12059,N_6593,N_5383);
nor U12060 (N_12060,N_8784,N_7255);
nand U12061 (N_12061,N_6571,N_8859);
xnor U12062 (N_12062,N_8491,N_8110);
nand U12063 (N_12063,N_6060,N_6233);
nand U12064 (N_12064,N_9879,N_8886);
and U12065 (N_12065,N_8501,N_6668);
and U12066 (N_12066,N_9412,N_9538);
nor U12067 (N_12067,N_6488,N_9806);
nor U12068 (N_12068,N_9220,N_5520);
nor U12069 (N_12069,N_7485,N_7936);
nand U12070 (N_12070,N_8936,N_8059);
nand U12071 (N_12071,N_5138,N_8314);
and U12072 (N_12072,N_7604,N_9714);
or U12073 (N_12073,N_6613,N_6915);
or U12074 (N_12074,N_5061,N_5682);
and U12075 (N_12075,N_7802,N_7494);
and U12076 (N_12076,N_9158,N_7762);
and U12077 (N_12077,N_6033,N_5431);
or U12078 (N_12078,N_6264,N_8827);
and U12079 (N_12079,N_8610,N_5441);
nor U12080 (N_12080,N_8546,N_8669);
and U12081 (N_12081,N_9483,N_6801);
nand U12082 (N_12082,N_7902,N_7010);
nor U12083 (N_12083,N_5921,N_8961);
nand U12084 (N_12084,N_7717,N_5998);
or U12085 (N_12085,N_7129,N_6599);
nor U12086 (N_12086,N_6367,N_5139);
and U12087 (N_12087,N_8041,N_5505);
and U12088 (N_12088,N_9089,N_7325);
and U12089 (N_12089,N_6414,N_7475);
nand U12090 (N_12090,N_6041,N_9746);
or U12091 (N_12091,N_9881,N_9420);
or U12092 (N_12092,N_6349,N_5278);
nor U12093 (N_12093,N_9857,N_9527);
nand U12094 (N_12094,N_6829,N_6334);
and U12095 (N_12095,N_7799,N_8508);
nand U12096 (N_12096,N_8254,N_7203);
and U12097 (N_12097,N_8641,N_7192);
xor U12098 (N_12098,N_8925,N_6728);
nor U12099 (N_12099,N_9848,N_8910);
or U12100 (N_12100,N_9711,N_7415);
nor U12101 (N_12101,N_9211,N_8978);
nor U12102 (N_12102,N_7142,N_9025);
or U12103 (N_12103,N_5126,N_5331);
and U12104 (N_12104,N_7022,N_7146);
and U12105 (N_12105,N_9940,N_7075);
and U12106 (N_12106,N_9884,N_6908);
nand U12107 (N_12107,N_6378,N_6070);
or U12108 (N_12108,N_5234,N_5782);
nor U12109 (N_12109,N_6637,N_9084);
nor U12110 (N_12110,N_9574,N_5912);
xor U12111 (N_12111,N_6666,N_7332);
and U12112 (N_12112,N_7712,N_9188);
and U12113 (N_12113,N_8067,N_8239);
and U12114 (N_12114,N_6244,N_6395);
and U12115 (N_12115,N_7436,N_7911);
nor U12116 (N_12116,N_9982,N_9264);
nand U12117 (N_12117,N_9192,N_9718);
or U12118 (N_12118,N_5034,N_5689);
or U12119 (N_12119,N_7532,N_7787);
nand U12120 (N_12120,N_6849,N_8386);
nand U12121 (N_12121,N_6848,N_7833);
and U12122 (N_12122,N_7242,N_9253);
nand U12123 (N_12123,N_8225,N_6692);
and U12124 (N_12124,N_8471,N_5243);
nor U12125 (N_12125,N_7466,N_9672);
or U12126 (N_12126,N_7390,N_8543);
nand U12127 (N_12127,N_7094,N_5749);
nand U12128 (N_12128,N_7994,N_8854);
nor U12129 (N_12129,N_8437,N_9048);
nand U12130 (N_12130,N_7124,N_5092);
nand U12131 (N_12131,N_7796,N_6561);
xnor U12132 (N_12132,N_5725,N_9090);
and U12133 (N_12133,N_6947,N_9289);
or U12134 (N_12134,N_5159,N_9685);
xnor U12135 (N_12135,N_5152,N_5359);
nor U12136 (N_12136,N_7042,N_7579);
nand U12137 (N_12137,N_9894,N_6532);
or U12138 (N_12138,N_7555,N_7830);
and U12139 (N_12139,N_9727,N_8426);
or U12140 (N_12140,N_7302,N_6324);
and U12141 (N_12141,N_7219,N_8653);
nand U12142 (N_12142,N_8097,N_6310);
and U12143 (N_12143,N_8786,N_6420);
or U12144 (N_12144,N_6218,N_5471);
nor U12145 (N_12145,N_5688,N_8308);
or U12146 (N_12146,N_8877,N_6049);
xnor U12147 (N_12147,N_9494,N_7144);
nand U12148 (N_12148,N_6461,N_7586);
or U12149 (N_12149,N_8470,N_8355);
nor U12150 (N_12150,N_7249,N_7294);
nand U12151 (N_12151,N_5992,N_8209);
or U12152 (N_12152,N_5098,N_5971);
nand U12153 (N_12153,N_6013,N_5362);
nand U12154 (N_12154,N_9603,N_8519);
or U12155 (N_12155,N_5227,N_9491);
nand U12156 (N_12156,N_8133,N_5684);
nand U12157 (N_12157,N_6097,N_5771);
nand U12158 (N_12158,N_8723,N_8938);
and U12159 (N_12159,N_9986,N_5214);
nor U12160 (N_12160,N_9352,N_8377);
nand U12161 (N_12161,N_7764,N_8682);
xnor U12162 (N_12162,N_7363,N_8242);
or U12163 (N_12163,N_6905,N_5748);
or U12164 (N_12164,N_8328,N_9206);
nor U12165 (N_12165,N_8880,N_7517);
nand U12166 (N_12166,N_5008,N_5533);
nor U12167 (N_12167,N_9892,N_7145);
nand U12168 (N_12168,N_6808,N_5724);
nor U12169 (N_12169,N_8277,N_8161);
nor U12170 (N_12170,N_6412,N_5137);
and U12171 (N_12171,N_9014,N_8357);
or U12172 (N_12172,N_6989,N_6409);
nor U12173 (N_12173,N_6874,N_8201);
and U12174 (N_12174,N_7564,N_6208);
nand U12175 (N_12175,N_5787,N_7613);
or U12176 (N_12176,N_9396,N_6658);
xor U12177 (N_12177,N_9605,N_5030);
and U12178 (N_12178,N_6490,N_7174);
or U12179 (N_12179,N_5464,N_7383);
xor U12180 (N_12180,N_8134,N_5217);
nor U12181 (N_12181,N_6758,N_7059);
or U12182 (N_12182,N_7382,N_7697);
nand U12183 (N_12183,N_7464,N_5177);
and U12184 (N_12184,N_8934,N_5953);
nor U12185 (N_12185,N_7643,N_8214);
or U12186 (N_12186,N_5571,N_5954);
nand U12187 (N_12187,N_8154,N_8701);
and U12188 (N_12188,N_9754,N_8828);
or U12189 (N_12189,N_5118,N_6628);
or U12190 (N_12190,N_5347,N_7044);
nand U12191 (N_12191,N_5320,N_8096);
and U12192 (N_12192,N_6904,N_7490);
or U12193 (N_12193,N_8835,N_5590);
nor U12194 (N_12194,N_8627,N_5063);
nand U12195 (N_12195,N_5547,N_5246);
or U12196 (N_12196,N_7344,N_9368);
nand U12197 (N_12197,N_9761,N_7919);
xnor U12198 (N_12198,N_8499,N_7096);
and U12199 (N_12199,N_7845,N_6009);
and U12200 (N_12200,N_5352,N_9945);
nand U12201 (N_12201,N_7166,N_6778);
nor U12202 (N_12202,N_7612,N_7026);
nor U12203 (N_12203,N_5130,N_8996);
or U12204 (N_12204,N_7258,N_8260);
and U12205 (N_12205,N_9079,N_6723);
or U12206 (N_12206,N_5232,N_6327);
nor U12207 (N_12207,N_7299,N_7515);
or U12208 (N_12208,N_7591,N_9965);
nand U12209 (N_12209,N_7675,N_9889);
or U12210 (N_12210,N_6142,N_9080);
or U12211 (N_12211,N_5550,N_6247);
nor U12212 (N_12212,N_6002,N_9261);
or U12213 (N_12213,N_8465,N_5955);
nor U12214 (N_12214,N_6709,N_7224);
nand U12215 (N_12215,N_5432,N_8903);
or U12216 (N_12216,N_8084,N_6431);
or U12217 (N_12217,N_6478,N_7318);
nor U12218 (N_12218,N_7654,N_6691);
nor U12219 (N_12219,N_6526,N_5845);
or U12220 (N_12220,N_6596,N_7206);
and U12221 (N_12221,N_7395,N_6166);
nand U12222 (N_12222,N_5965,N_7469);
or U12223 (N_12223,N_7772,N_9825);
xor U12224 (N_12224,N_6775,N_6529);
or U12225 (N_12225,N_5978,N_5376);
nor U12226 (N_12226,N_5340,N_9707);
nand U12227 (N_12227,N_5225,N_7251);
nor U12228 (N_12228,N_6671,N_5202);
or U12229 (N_12229,N_7575,N_5326);
nand U12230 (N_12230,N_5438,N_5336);
nor U12231 (N_12231,N_8101,N_5679);
nor U12232 (N_12232,N_5086,N_7569);
nand U12233 (N_12233,N_9566,N_7218);
nand U12234 (N_12234,N_8572,N_7023);
and U12235 (N_12235,N_6441,N_8438);
nor U12236 (N_12236,N_7221,N_8498);
and U12237 (N_12237,N_5329,N_8494);
nand U12238 (N_12238,N_7537,N_8430);
nand U12239 (N_12239,N_5654,N_9051);
and U12240 (N_12240,N_5492,N_8179);
nand U12241 (N_12241,N_6509,N_9634);
xnor U12242 (N_12242,N_7329,N_5447);
and U12243 (N_12243,N_5882,N_8731);
and U12244 (N_12244,N_5283,N_9452);
nand U12245 (N_12245,N_6197,N_6011);
nor U12246 (N_12246,N_6960,N_7287);
xor U12247 (N_12247,N_6859,N_5333);
or U12248 (N_12248,N_8062,N_7597);
nor U12249 (N_12249,N_8289,N_5479);
nand U12250 (N_12250,N_7188,N_9646);
nand U12251 (N_12251,N_8002,N_7757);
or U12252 (N_12252,N_6004,N_7139);
or U12253 (N_12253,N_7695,N_8733);
and U12254 (N_12254,N_8475,N_7268);
nand U12255 (N_12255,N_5006,N_9929);
nand U12256 (N_12256,N_6852,N_6619);
and U12257 (N_12257,N_9643,N_8248);
or U12258 (N_12258,N_7157,N_9474);
and U12259 (N_12259,N_5558,N_6464);
and U12260 (N_12260,N_8136,N_7975);
or U12261 (N_12261,N_6326,N_9536);
xnor U12262 (N_12262,N_6912,N_6341);
nand U12263 (N_12263,N_9570,N_8760);
nor U12264 (N_12264,N_8861,N_6016);
and U12265 (N_12265,N_9859,N_8600);
nor U12266 (N_12266,N_7931,N_5106);
nor U12267 (N_12267,N_8696,N_9291);
nor U12268 (N_12268,N_9541,N_5448);
nor U12269 (N_12269,N_9344,N_8656);
nand U12270 (N_12270,N_6133,N_7731);
xnor U12271 (N_12271,N_9481,N_6053);
or U12272 (N_12272,N_7313,N_6240);
nand U12273 (N_12273,N_5038,N_8578);
nor U12274 (N_12274,N_8169,N_8479);
or U12275 (N_12275,N_9823,N_9540);
and U12276 (N_12276,N_7752,N_8834);
and U12277 (N_12277,N_5349,N_8685);
xnor U12278 (N_12278,N_9010,N_5273);
nor U12279 (N_12279,N_6955,N_8462);
nand U12280 (N_12280,N_5293,N_7167);
or U12281 (N_12281,N_6641,N_9720);
nor U12282 (N_12282,N_5578,N_5798);
nor U12283 (N_12283,N_9484,N_9003);
nand U12284 (N_12284,N_8417,N_5018);
nand U12285 (N_12285,N_8421,N_9710);
or U12286 (N_12286,N_9068,N_9478);
and U12287 (N_12287,N_9903,N_7767);
nor U12288 (N_12288,N_7835,N_8266);
xnor U12289 (N_12289,N_5264,N_8763);
nor U12290 (N_12290,N_8463,N_6968);
xnor U12291 (N_12291,N_6527,N_7619);
and U12292 (N_12292,N_5353,N_8455);
or U12293 (N_12293,N_5513,N_6162);
nor U12294 (N_12294,N_8177,N_8715);
and U12295 (N_12295,N_9275,N_5075);
nor U12296 (N_12296,N_7099,N_7988);
nor U12297 (N_12297,N_8818,N_9433);
and U12298 (N_12298,N_9116,N_8272);
or U12299 (N_12299,N_6121,N_9340);
and U12300 (N_12300,N_7402,N_7314);
and U12301 (N_12301,N_8616,N_6553);
and U12302 (N_12302,N_7337,N_6167);
or U12303 (N_12303,N_8291,N_8450);
or U12304 (N_12304,N_9461,N_7681);
and U12305 (N_12305,N_8326,N_5948);
and U12306 (N_12306,N_5132,N_7477);
nand U12307 (N_12307,N_9521,N_5046);
nand U12308 (N_12308,N_8425,N_7599);
nand U12309 (N_12309,N_6077,N_7343);
xor U12310 (N_12310,N_7933,N_8533);
nand U12311 (N_12311,N_5122,N_5577);
nand U12312 (N_12312,N_8640,N_7688);
or U12313 (N_12313,N_7554,N_8690);
nand U12314 (N_12314,N_7079,N_8557);
and U12315 (N_12315,N_9957,N_6896);
xor U12316 (N_12316,N_5738,N_7199);
nor U12317 (N_12317,N_8565,N_6168);
nand U12318 (N_12318,N_8703,N_6885);
and U12319 (N_12319,N_5010,N_8315);
nand U12320 (N_12320,N_9597,N_7724);
and U12321 (N_12321,N_9164,N_5270);
nand U12322 (N_12322,N_7679,N_7043);
nand U12323 (N_12323,N_7927,N_8698);
and U12324 (N_12324,N_6080,N_8483);
or U12325 (N_12325,N_9522,N_5729);
and U12326 (N_12326,N_6363,N_6109);
nand U12327 (N_12327,N_7504,N_7371);
and U12328 (N_12328,N_9525,N_8689);
nor U12329 (N_12329,N_8001,N_5402);
nand U12330 (N_12330,N_9343,N_8921);
or U12331 (N_12331,N_8387,N_6071);
nor U12332 (N_12332,N_9095,N_6224);
and U12333 (N_12333,N_7822,N_8737);
nand U12334 (N_12334,N_7114,N_9088);
or U12335 (N_12335,N_7671,N_5419);
xor U12336 (N_12336,N_5646,N_9301);
nor U12337 (N_12337,N_8271,N_7522);
xor U12338 (N_12338,N_7573,N_5741);
nor U12339 (N_12339,N_5546,N_6061);
nor U12340 (N_12340,N_5405,N_6440);
or U12341 (N_12341,N_6144,N_7457);
and U12342 (N_12342,N_9462,N_9327);
nor U12343 (N_12343,N_9567,N_9254);
nor U12344 (N_12344,N_9935,N_9335);
nand U12345 (N_12345,N_9875,N_7133);
nand U12346 (N_12346,N_5449,N_5230);
nand U12347 (N_12347,N_5335,N_9150);
nand U12348 (N_12348,N_6320,N_9717);
nor U12349 (N_12349,N_9282,N_9733);
and U12350 (N_12350,N_9224,N_6549);
xnor U12351 (N_12351,N_8370,N_9062);
nor U12352 (N_12352,N_5169,N_5583);
and U12353 (N_12353,N_7264,N_8295);
and U12354 (N_12354,N_5896,N_7899);
xor U12355 (N_12355,N_7766,N_9994);
nor U12356 (N_12356,N_5239,N_7200);
nand U12357 (N_12357,N_9469,N_9908);
or U12358 (N_12358,N_7662,N_6890);
and U12359 (N_12359,N_5144,N_5861);
or U12360 (N_12360,N_5029,N_7983);
nand U12361 (N_12361,N_7177,N_5341);
nor U12362 (N_12362,N_9009,N_7261);
nor U12363 (N_12363,N_6932,N_5653);
nor U12364 (N_12364,N_6427,N_8550);
or U12365 (N_12365,N_9532,N_9425);
or U12366 (N_12366,N_9440,N_5536);
nand U12367 (N_12367,N_5149,N_7409);
or U12368 (N_12368,N_6063,N_8045);
nor U12369 (N_12369,N_5510,N_8789);
nand U12370 (N_12370,N_5473,N_9248);
nor U12371 (N_12371,N_6742,N_9805);
or U12372 (N_12372,N_8126,N_7924);
and U12373 (N_12373,N_6073,N_6157);
or U12374 (N_12374,N_6747,N_8750);
nand U12375 (N_12375,N_5166,N_7006);
nand U12376 (N_12376,N_8691,N_9607);
and U12377 (N_12377,N_5260,N_5956);
nand U12378 (N_12378,N_6903,N_8167);
nand U12379 (N_12379,N_7216,N_8817);
nor U12380 (N_12380,N_5095,N_5842);
and U12381 (N_12381,N_9564,N_6662);
or U12382 (N_12382,N_9663,N_8446);
nand U12383 (N_12383,N_6831,N_7423);
nor U12384 (N_12384,N_6603,N_9159);
nor U12385 (N_12385,N_9078,N_7758);
or U12386 (N_12386,N_7186,N_9252);
nor U12387 (N_12387,N_8108,N_6421);
nor U12388 (N_12388,N_9796,N_9810);
nand U12389 (N_12389,N_8805,N_8412);
and U12390 (N_12390,N_8286,N_6736);
xor U12391 (N_12391,N_8339,N_9882);
or U12392 (N_12392,N_8264,N_5250);
and U12393 (N_12393,N_5190,N_9450);
or U12394 (N_12394,N_9553,N_7559);
nand U12395 (N_12395,N_9993,N_8107);
nor U12396 (N_12396,N_8740,N_7906);
nand U12397 (N_12397,N_6555,N_7165);
or U12398 (N_12398,N_6190,N_7252);
nor U12399 (N_12399,N_6394,N_6076);
nor U12400 (N_12400,N_8734,N_7682);
or U12401 (N_12401,N_6545,N_8589);
nand U12402 (N_12402,N_5856,N_9240);
or U12403 (N_12403,N_9148,N_9551);
nor U12404 (N_12404,N_6354,N_6963);
nand U12405 (N_12405,N_7721,N_6546);
or U12406 (N_12406,N_6351,N_7438);
or U12407 (N_12407,N_5134,N_8075);
nor U12408 (N_12408,N_9341,N_9926);
and U12409 (N_12409,N_6832,N_7093);
xnor U12410 (N_12410,N_7280,N_9562);
or U12411 (N_12411,N_5275,N_5182);
nand U12412 (N_12412,N_5366,N_9800);
or U12413 (N_12413,N_8563,N_8036);
or U12414 (N_12414,N_7227,N_7600);
nor U12415 (N_12415,N_9931,N_5292);
nor U12416 (N_12416,N_8825,N_9534);
and U12417 (N_12417,N_5368,N_6134);
nand U12418 (N_12418,N_8785,N_8807);
or U12419 (N_12419,N_9679,N_7746);
xor U12420 (N_12420,N_8914,N_5324);
nand U12421 (N_12421,N_5031,N_7748);
nand U12422 (N_12422,N_9916,N_9057);
and U12423 (N_12423,N_5586,N_7013);
or U12424 (N_12424,N_9406,N_5908);
or U12425 (N_12425,N_6855,N_5233);
nor U12426 (N_12426,N_6048,N_9565);
or U12427 (N_12427,N_6528,N_8213);
and U12428 (N_12428,N_5218,N_8868);
and U12429 (N_12429,N_6025,N_7505);
nand U12430 (N_12430,N_6538,N_9524);
nand U12431 (N_12431,N_6595,N_9471);
nand U12432 (N_12432,N_9695,N_9690);
nor U12433 (N_12433,N_7992,N_8135);
xnor U12434 (N_12434,N_9171,N_6321);
nand U12435 (N_12435,N_6966,N_9649);
and U12436 (N_12436,N_7566,N_5054);
or U12437 (N_12437,N_6491,N_9124);
nor U12438 (N_12438,N_5715,N_9560);
nand U12439 (N_12439,N_8643,N_9529);
nand U12440 (N_12440,N_7328,N_9807);
and U12441 (N_12441,N_6851,N_9756);
and U12442 (N_12442,N_9487,N_7476);
nand U12443 (N_12443,N_9696,N_9503);
and U12444 (N_12444,N_7256,N_9203);
nand U12445 (N_12445,N_5515,N_6411);
and U12446 (N_12446,N_7595,N_5668);
xnor U12447 (N_12447,N_7867,N_6350);
nor U12448 (N_12448,N_6184,N_9966);
nor U12449 (N_12449,N_5163,N_8369);
nand U12450 (N_12450,N_8086,N_9175);
and U12451 (N_12451,N_7669,N_9409);
or U12452 (N_12452,N_8712,N_5800);
xor U12453 (N_12453,N_7470,N_5645);
or U12454 (N_12454,N_7963,N_9799);
nand U12455 (N_12455,N_6323,N_9251);
nand U12456 (N_12456,N_6284,N_6430);
and U12457 (N_12457,N_7859,N_6838);
nor U12458 (N_12458,N_8352,N_6881);
or U12459 (N_12459,N_8506,N_7331);
xnor U12460 (N_12460,N_7540,N_8415);
xor U12461 (N_12461,N_5810,N_8237);
nand U12462 (N_12462,N_8189,N_5263);
nor U12463 (N_12463,N_8140,N_8363);
and U12464 (N_12464,N_6557,N_9992);
and U12465 (N_12465,N_8782,N_9094);
nor U12466 (N_12466,N_9392,N_8362);
or U12467 (N_12467,N_8678,N_8573);
and U12468 (N_12468,N_5394,N_6413);
or U12469 (N_12469,N_7628,N_8707);
or U12470 (N_12470,N_5807,N_9670);
nand U12471 (N_12471,N_7852,N_8111);
xnor U12472 (N_12472,N_5808,N_6972);
xnor U12473 (N_12473,N_9873,N_8488);
or U12474 (N_12474,N_6634,N_8020);
nor U12475 (N_12475,N_5153,N_9953);
xnor U12476 (N_12476,N_6627,N_9263);
and U12477 (N_12477,N_8381,N_8256);
nor U12478 (N_12478,N_6695,N_7623);
or U12479 (N_12479,N_8400,N_8694);
and U12480 (N_12480,N_6717,N_5743);
nand U12481 (N_12481,N_5819,N_5853);
or U12482 (N_12482,N_5841,N_6523);
or U12483 (N_12483,N_7842,N_5809);
or U12484 (N_12484,N_7427,N_7080);
and U12485 (N_12485,N_6045,N_9559);
nor U12486 (N_12486,N_9673,N_5496);
or U12487 (N_12487,N_9361,N_7009);
and U12488 (N_12488,N_8486,N_5364);
nor U12489 (N_12489,N_6876,N_7508);
nor U12490 (N_12490,N_5621,N_8184);
or U12491 (N_12491,N_8890,N_6981);
or U12492 (N_12492,N_5487,N_8141);
and U12493 (N_12493,N_5284,N_9909);
and U12494 (N_12494,N_8231,N_6135);
or U12495 (N_12495,N_6880,N_9863);
or U12496 (N_12496,N_9402,N_6999);
nand U12497 (N_12497,N_9058,N_7384);
nand U12498 (N_12498,N_5700,N_8621);
nor U12499 (N_12499,N_9366,N_9004);
nand U12500 (N_12500,N_5021,N_9683);
xnor U12501 (N_12501,N_6980,N_9481);
nand U12502 (N_12502,N_6655,N_6447);
or U12503 (N_12503,N_5186,N_8319);
or U12504 (N_12504,N_5461,N_5336);
nor U12505 (N_12505,N_8439,N_6069);
nor U12506 (N_12506,N_8471,N_5980);
nor U12507 (N_12507,N_9378,N_7210);
nor U12508 (N_12508,N_6596,N_5089);
nand U12509 (N_12509,N_5517,N_7336);
nand U12510 (N_12510,N_5129,N_8234);
nor U12511 (N_12511,N_5211,N_6181);
and U12512 (N_12512,N_9431,N_9251);
nor U12513 (N_12513,N_8668,N_9074);
nor U12514 (N_12514,N_5947,N_6546);
and U12515 (N_12515,N_7887,N_5767);
and U12516 (N_12516,N_8903,N_6594);
or U12517 (N_12517,N_9290,N_8933);
or U12518 (N_12518,N_7250,N_6401);
or U12519 (N_12519,N_7223,N_9926);
nand U12520 (N_12520,N_8451,N_6170);
and U12521 (N_12521,N_9164,N_9224);
or U12522 (N_12522,N_5636,N_6777);
xnor U12523 (N_12523,N_9082,N_6950);
nor U12524 (N_12524,N_6062,N_8770);
nor U12525 (N_12525,N_5928,N_7061);
and U12526 (N_12526,N_7644,N_9170);
or U12527 (N_12527,N_5062,N_6072);
or U12528 (N_12528,N_7801,N_7107);
nor U12529 (N_12529,N_9590,N_9341);
xor U12530 (N_12530,N_6159,N_5020);
nor U12531 (N_12531,N_6988,N_7700);
xnor U12532 (N_12532,N_9058,N_6158);
nand U12533 (N_12533,N_8906,N_7836);
nor U12534 (N_12534,N_5167,N_7901);
and U12535 (N_12535,N_6077,N_6654);
and U12536 (N_12536,N_8486,N_7943);
nor U12537 (N_12537,N_8622,N_7100);
and U12538 (N_12538,N_9437,N_9290);
nor U12539 (N_12539,N_9611,N_6585);
and U12540 (N_12540,N_7927,N_5253);
xnor U12541 (N_12541,N_5719,N_9395);
or U12542 (N_12542,N_9349,N_7883);
nor U12543 (N_12543,N_7569,N_9197);
and U12544 (N_12544,N_7119,N_6954);
and U12545 (N_12545,N_7067,N_5033);
xor U12546 (N_12546,N_6620,N_5515);
or U12547 (N_12547,N_9707,N_8051);
or U12548 (N_12548,N_9869,N_6831);
and U12549 (N_12549,N_9773,N_8245);
nor U12550 (N_12550,N_7878,N_5543);
or U12551 (N_12551,N_5616,N_9246);
nor U12552 (N_12552,N_5239,N_8402);
nand U12553 (N_12553,N_8723,N_9938);
or U12554 (N_12554,N_7975,N_6611);
nor U12555 (N_12555,N_6454,N_9631);
or U12556 (N_12556,N_5473,N_6166);
nor U12557 (N_12557,N_8900,N_8871);
nor U12558 (N_12558,N_9693,N_8825);
or U12559 (N_12559,N_9621,N_5058);
and U12560 (N_12560,N_6228,N_9875);
or U12561 (N_12561,N_6623,N_8075);
or U12562 (N_12562,N_6496,N_9577);
or U12563 (N_12563,N_7265,N_7138);
nor U12564 (N_12564,N_7609,N_7426);
nor U12565 (N_12565,N_9271,N_6514);
and U12566 (N_12566,N_6891,N_6633);
nand U12567 (N_12567,N_9686,N_8848);
nand U12568 (N_12568,N_6411,N_8834);
nor U12569 (N_12569,N_5258,N_9160);
or U12570 (N_12570,N_8682,N_9839);
nand U12571 (N_12571,N_6532,N_5956);
or U12572 (N_12572,N_7420,N_6783);
or U12573 (N_12573,N_7670,N_5718);
nor U12574 (N_12574,N_6208,N_5339);
xor U12575 (N_12575,N_6159,N_9259);
or U12576 (N_12576,N_6219,N_6455);
or U12577 (N_12577,N_8121,N_8694);
nor U12578 (N_12578,N_7990,N_6413);
and U12579 (N_12579,N_8402,N_5074);
nand U12580 (N_12580,N_6221,N_7283);
or U12581 (N_12581,N_5370,N_5084);
or U12582 (N_12582,N_9318,N_9699);
nor U12583 (N_12583,N_8402,N_8946);
nor U12584 (N_12584,N_6775,N_8390);
nor U12585 (N_12585,N_7707,N_7337);
nor U12586 (N_12586,N_6836,N_7258);
nand U12587 (N_12587,N_9102,N_6721);
nor U12588 (N_12588,N_5282,N_6916);
nand U12589 (N_12589,N_5573,N_7871);
or U12590 (N_12590,N_7210,N_7335);
nand U12591 (N_12591,N_8799,N_8613);
and U12592 (N_12592,N_5032,N_7891);
nand U12593 (N_12593,N_5134,N_7589);
and U12594 (N_12594,N_9525,N_8387);
nor U12595 (N_12595,N_5677,N_6283);
nand U12596 (N_12596,N_5309,N_9298);
nor U12597 (N_12597,N_8437,N_9570);
nand U12598 (N_12598,N_6252,N_7041);
or U12599 (N_12599,N_7062,N_8003);
nor U12600 (N_12600,N_7266,N_9367);
nor U12601 (N_12601,N_5079,N_5049);
or U12602 (N_12602,N_7633,N_8879);
and U12603 (N_12603,N_7180,N_7545);
and U12604 (N_12604,N_6850,N_6232);
nand U12605 (N_12605,N_8340,N_5612);
nand U12606 (N_12606,N_7513,N_5298);
nand U12607 (N_12607,N_5664,N_7503);
nor U12608 (N_12608,N_7926,N_8905);
nand U12609 (N_12609,N_7488,N_9683);
or U12610 (N_12610,N_7205,N_6542);
nor U12611 (N_12611,N_9159,N_6887);
and U12612 (N_12612,N_9329,N_6970);
nor U12613 (N_12613,N_8891,N_7266);
or U12614 (N_12614,N_8202,N_7361);
nand U12615 (N_12615,N_8001,N_8560);
nor U12616 (N_12616,N_6974,N_7803);
nor U12617 (N_12617,N_6716,N_9449);
and U12618 (N_12618,N_7689,N_9014);
xor U12619 (N_12619,N_9025,N_9284);
and U12620 (N_12620,N_8204,N_9242);
or U12621 (N_12621,N_8368,N_7503);
nor U12622 (N_12622,N_7631,N_8417);
or U12623 (N_12623,N_7632,N_6076);
nor U12624 (N_12624,N_6295,N_8493);
nand U12625 (N_12625,N_6940,N_8348);
or U12626 (N_12626,N_9834,N_7315);
nand U12627 (N_12627,N_7727,N_7460);
nor U12628 (N_12628,N_5835,N_8616);
xnor U12629 (N_12629,N_5364,N_7836);
nand U12630 (N_12630,N_8802,N_7330);
xor U12631 (N_12631,N_5234,N_5181);
nor U12632 (N_12632,N_8068,N_9938);
xnor U12633 (N_12633,N_7575,N_9755);
nand U12634 (N_12634,N_5818,N_5833);
nor U12635 (N_12635,N_5027,N_8723);
nor U12636 (N_12636,N_7175,N_5682);
nor U12637 (N_12637,N_5480,N_8423);
or U12638 (N_12638,N_6245,N_8448);
or U12639 (N_12639,N_5913,N_8471);
nand U12640 (N_12640,N_6080,N_9114);
nand U12641 (N_12641,N_8661,N_6257);
nor U12642 (N_12642,N_6224,N_7194);
or U12643 (N_12643,N_7919,N_9373);
xor U12644 (N_12644,N_5191,N_8335);
nand U12645 (N_12645,N_7443,N_6172);
nand U12646 (N_12646,N_8621,N_6334);
or U12647 (N_12647,N_9154,N_6979);
nor U12648 (N_12648,N_7099,N_6029);
xor U12649 (N_12649,N_6775,N_5050);
nand U12650 (N_12650,N_5930,N_8182);
nor U12651 (N_12651,N_8861,N_9671);
or U12652 (N_12652,N_6248,N_6604);
or U12653 (N_12653,N_7081,N_5079);
and U12654 (N_12654,N_5154,N_9050);
and U12655 (N_12655,N_8870,N_7117);
nor U12656 (N_12656,N_9691,N_6258);
nor U12657 (N_12657,N_9104,N_9618);
nand U12658 (N_12658,N_5852,N_5409);
or U12659 (N_12659,N_7183,N_5639);
and U12660 (N_12660,N_9704,N_7908);
or U12661 (N_12661,N_8699,N_9698);
or U12662 (N_12662,N_6964,N_5331);
nand U12663 (N_12663,N_6013,N_8681);
nor U12664 (N_12664,N_9084,N_8230);
or U12665 (N_12665,N_7042,N_9736);
nor U12666 (N_12666,N_7920,N_9131);
and U12667 (N_12667,N_7940,N_7722);
and U12668 (N_12668,N_9402,N_6033);
or U12669 (N_12669,N_5533,N_8634);
xor U12670 (N_12670,N_8454,N_6937);
and U12671 (N_12671,N_7860,N_5928);
and U12672 (N_12672,N_6147,N_6924);
nor U12673 (N_12673,N_9463,N_6269);
nor U12674 (N_12674,N_9575,N_9232);
nor U12675 (N_12675,N_7466,N_6016);
and U12676 (N_12676,N_6983,N_5697);
nand U12677 (N_12677,N_9157,N_7678);
or U12678 (N_12678,N_5076,N_8643);
and U12679 (N_12679,N_7276,N_9206);
nand U12680 (N_12680,N_8429,N_6257);
and U12681 (N_12681,N_6270,N_8581);
and U12682 (N_12682,N_5284,N_8963);
or U12683 (N_12683,N_5357,N_7385);
or U12684 (N_12684,N_6857,N_9915);
or U12685 (N_12685,N_6976,N_6079);
and U12686 (N_12686,N_9914,N_9983);
or U12687 (N_12687,N_8425,N_6345);
nand U12688 (N_12688,N_6918,N_6633);
or U12689 (N_12689,N_8115,N_8062);
nor U12690 (N_12690,N_9177,N_8703);
nand U12691 (N_12691,N_5617,N_7192);
nor U12692 (N_12692,N_7490,N_5086);
xnor U12693 (N_12693,N_8138,N_6994);
xor U12694 (N_12694,N_8760,N_7579);
nand U12695 (N_12695,N_9309,N_9316);
nand U12696 (N_12696,N_7876,N_6910);
or U12697 (N_12697,N_7136,N_5759);
nor U12698 (N_12698,N_6831,N_8856);
nor U12699 (N_12699,N_9575,N_9098);
nand U12700 (N_12700,N_7692,N_5043);
or U12701 (N_12701,N_5913,N_7381);
or U12702 (N_12702,N_7174,N_5930);
and U12703 (N_12703,N_7696,N_9244);
xnor U12704 (N_12704,N_5169,N_5048);
and U12705 (N_12705,N_5639,N_7125);
or U12706 (N_12706,N_9469,N_6451);
or U12707 (N_12707,N_8639,N_8137);
and U12708 (N_12708,N_7306,N_8971);
nor U12709 (N_12709,N_5225,N_6935);
xnor U12710 (N_12710,N_6501,N_8672);
or U12711 (N_12711,N_5057,N_9730);
xor U12712 (N_12712,N_8191,N_6930);
xnor U12713 (N_12713,N_5488,N_7781);
or U12714 (N_12714,N_8538,N_9924);
nand U12715 (N_12715,N_6737,N_9520);
or U12716 (N_12716,N_7136,N_6635);
xor U12717 (N_12717,N_6228,N_6048);
and U12718 (N_12718,N_5355,N_8865);
xor U12719 (N_12719,N_5300,N_9234);
nand U12720 (N_12720,N_7454,N_9699);
and U12721 (N_12721,N_6179,N_7865);
xnor U12722 (N_12722,N_9067,N_5071);
nand U12723 (N_12723,N_7894,N_6475);
nor U12724 (N_12724,N_8430,N_7630);
xor U12725 (N_12725,N_9141,N_6162);
and U12726 (N_12726,N_7217,N_8901);
nand U12727 (N_12727,N_6086,N_7812);
nand U12728 (N_12728,N_7643,N_9409);
nor U12729 (N_12729,N_8285,N_5370);
nand U12730 (N_12730,N_5329,N_8387);
or U12731 (N_12731,N_7438,N_5833);
or U12732 (N_12732,N_8031,N_9900);
or U12733 (N_12733,N_7432,N_8958);
nand U12734 (N_12734,N_7381,N_7455);
nand U12735 (N_12735,N_5502,N_8363);
or U12736 (N_12736,N_6769,N_7726);
and U12737 (N_12737,N_9753,N_8232);
nand U12738 (N_12738,N_9256,N_6601);
and U12739 (N_12739,N_8261,N_9879);
xnor U12740 (N_12740,N_7738,N_7971);
or U12741 (N_12741,N_8506,N_6637);
nor U12742 (N_12742,N_5704,N_7075);
or U12743 (N_12743,N_8410,N_8673);
and U12744 (N_12744,N_5387,N_7617);
and U12745 (N_12745,N_6608,N_8549);
nor U12746 (N_12746,N_6018,N_9215);
nor U12747 (N_12747,N_7494,N_6696);
nor U12748 (N_12748,N_6070,N_7102);
nor U12749 (N_12749,N_9418,N_9155);
or U12750 (N_12750,N_6448,N_6903);
nand U12751 (N_12751,N_9353,N_5271);
or U12752 (N_12752,N_8130,N_9503);
nand U12753 (N_12753,N_5270,N_5486);
or U12754 (N_12754,N_9935,N_7796);
nand U12755 (N_12755,N_5958,N_6113);
nand U12756 (N_12756,N_7971,N_9252);
and U12757 (N_12757,N_5057,N_7396);
nand U12758 (N_12758,N_7266,N_6327);
and U12759 (N_12759,N_9855,N_8575);
nor U12760 (N_12760,N_8164,N_5484);
xnor U12761 (N_12761,N_8395,N_6161);
nand U12762 (N_12762,N_9186,N_8923);
and U12763 (N_12763,N_5507,N_5061);
xor U12764 (N_12764,N_9032,N_9033);
nand U12765 (N_12765,N_5736,N_8283);
or U12766 (N_12766,N_5627,N_6828);
nor U12767 (N_12767,N_8523,N_9285);
nor U12768 (N_12768,N_7392,N_6693);
nor U12769 (N_12769,N_5309,N_7687);
or U12770 (N_12770,N_6713,N_6421);
nor U12771 (N_12771,N_5659,N_5930);
nor U12772 (N_12772,N_8183,N_5716);
xnor U12773 (N_12773,N_8625,N_6529);
nand U12774 (N_12774,N_8776,N_7065);
nor U12775 (N_12775,N_9259,N_8072);
nand U12776 (N_12776,N_8474,N_5716);
and U12777 (N_12777,N_6098,N_6839);
and U12778 (N_12778,N_8013,N_6774);
or U12779 (N_12779,N_7222,N_5693);
nand U12780 (N_12780,N_5780,N_8068);
or U12781 (N_12781,N_7820,N_8597);
and U12782 (N_12782,N_5063,N_8811);
or U12783 (N_12783,N_8110,N_5538);
and U12784 (N_12784,N_8659,N_8729);
nor U12785 (N_12785,N_6506,N_7321);
nand U12786 (N_12786,N_6753,N_9351);
nor U12787 (N_12787,N_6201,N_5142);
nor U12788 (N_12788,N_8220,N_7653);
xor U12789 (N_12789,N_5669,N_6745);
nor U12790 (N_12790,N_7805,N_5879);
xor U12791 (N_12791,N_7682,N_5239);
nor U12792 (N_12792,N_7472,N_8383);
nand U12793 (N_12793,N_5942,N_7263);
or U12794 (N_12794,N_9101,N_7289);
nor U12795 (N_12795,N_5878,N_8818);
nand U12796 (N_12796,N_8333,N_6677);
xor U12797 (N_12797,N_8377,N_6217);
and U12798 (N_12798,N_9100,N_9638);
and U12799 (N_12799,N_8800,N_6377);
nand U12800 (N_12800,N_7705,N_7903);
nor U12801 (N_12801,N_9250,N_9053);
nor U12802 (N_12802,N_7513,N_6525);
and U12803 (N_12803,N_9735,N_5563);
nor U12804 (N_12804,N_7208,N_8861);
or U12805 (N_12805,N_7991,N_5456);
or U12806 (N_12806,N_6324,N_8788);
nor U12807 (N_12807,N_8149,N_5003);
nor U12808 (N_12808,N_9123,N_9438);
nand U12809 (N_12809,N_7035,N_7788);
nand U12810 (N_12810,N_6061,N_9674);
nand U12811 (N_12811,N_5061,N_7737);
xnor U12812 (N_12812,N_6995,N_5999);
nand U12813 (N_12813,N_6084,N_6793);
and U12814 (N_12814,N_8182,N_9329);
xor U12815 (N_12815,N_6185,N_8061);
or U12816 (N_12816,N_7763,N_5945);
nor U12817 (N_12817,N_6453,N_6769);
or U12818 (N_12818,N_6507,N_7484);
and U12819 (N_12819,N_8388,N_8900);
nand U12820 (N_12820,N_5966,N_8927);
nand U12821 (N_12821,N_9499,N_6247);
xnor U12822 (N_12822,N_8133,N_9346);
xor U12823 (N_12823,N_6410,N_8983);
or U12824 (N_12824,N_5803,N_8195);
nand U12825 (N_12825,N_6073,N_9873);
nand U12826 (N_12826,N_8226,N_8189);
and U12827 (N_12827,N_6212,N_9444);
and U12828 (N_12828,N_9935,N_8048);
or U12829 (N_12829,N_8352,N_6624);
nand U12830 (N_12830,N_6332,N_6059);
nor U12831 (N_12831,N_9773,N_6619);
nand U12832 (N_12832,N_7598,N_9280);
nor U12833 (N_12833,N_5427,N_8635);
xor U12834 (N_12834,N_9874,N_9619);
nor U12835 (N_12835,N_9633,N_9738);
nor U12836 (N_12836,N_5972,N_9535);
and U12837 (N_12837,N_7635,N_6811);
nor U12838 (N_12838,N_9468,N_5999);
nor U12839 (N_12839,N_9545,N_9712);
nand U12840 (N_12840,N_6508,N_9641);
nor U12841 (N_12841,N_9711,N_9940);
and U12842 (N_12842,N_6830,N_6142);
or U12843 (N_12843,N_8711,N_8149);
nor U12844 (N_12844,N_6615,N_7462);
nand U12845 (N_12845,N_9332,N_7733);
nor U12846 (N_12846,N_6974,N_8026);
nor U12847 (N_12847,N_7757,N_7726);
or U12848 (N_12848,N_5910,N_9944);
xor U12849 (N_12849,N_9231,N_6077);
nand U12850 (N_12850,N_8314,N_7300);
nand U12851 (N_12851,N_9020,N_5591);
and U12852 (N_12852,N_8655,N_7928);
nand U12853 (N_12853,N_9851,N_5730);
nand U12854 (N_12854,N_7669,N_8890);
or U12855 (N_12855,N_8856,N_6869);
and U12856 (N_12856,N_5073,N_8814);
or U12857 (N_12857,N_8885,N_7333);
or U12858 (N_12858,N_7980,N_8359);
xor U12859 (N_12859,N_5894,N_5012);
nor U12860 (N_12860,N_9270,N_7769);
nor U12861 (N_12861,N_7586,N_9963);
nand U12862 (N_12862,N_5097,N_9462);
and U12863 (N_12863,N_7464,N_5316);
xor U12864 (N_12864,N_5187,N_6479);
or U12865 (N_12865,N_8751,N_5064);
and U12866 (N_12866,N_9789,N_7382);
nor U12867 (N_12867,N_8264,N_5395);
and U12868 (N_12868,N_5553,N_5295);
or U12869 (N_12869,N_8950,N_7883);
nor U12870 (N_12870,N_6869,N_7741);
nor U12871 (N_12871,N_5639,N_7720);
nor U12872 (N_12872,N_9458,N_8440);
nand U12873 (N_12873,N_9819,N_7380);
and U12874 (N_12874,N_6979,N_9826);
nand U12875 (N_12875,N_5731,N_7519);
xnor U12876 (N_12876,N_6074,N_6692);
or U12877 (N_12877,N_8631,N_7788);
xnor U12878 (N_12878,N_7378,N_9735);
nor U12879 (N_12879,N_5701,N_5569);
nor U12880 (N_12880,N_7516,N_9758);
nand U12881 (N_12881,N_5820,N_6852);
nor U12882 (N_12882,N_8661,N_8295);
xor U12883 (N_12883,N_8615,N_8581);
and U12884 (N_12884,N_8800,N_9669);
nand U12885 (N_12885,N_8877,N_5585);
or U12886 (N_12886,N_9590,N_8866);
and U12887 (N_12887,N_7935,N_6861);
or U12888 (N_12888,N_9159,N_6486);
or U12889 (N_12889,N_9920,N_9877);
and U12890 (N_12890,N_7138,N_5183);
nand U12891 (N_12891,N_7232,N_9850);
and U12892 (N_12892,N_6039,N_9394);
and U12893 (N_12893,N_6756,N_8044);
or U12894 (N_12894,N_5099,N_7691);
nor U12895 (N_12895,N_9851,N_6548);
and U12896 (N_12896,N_5114,N_6751);
nor U12897 (N_12897,N_8918,N_7510);
or U12898 (N_12898,N_6466,N_5828);
xnor U12899 (N_12899,N_9327,N_9721);
nor U12900 (N_12900,N_6365,N_6780);
or U12901 (N_12901,N_9503,N_9276);
nand U12902 (N_12902,N_7477,N_8088);
or U12903 (N_12903,N_5078,N_5617);
nand U12904 (N_12904,N_5118,N_5332);
nor U12905 (N_12905,N_8475,N_8819);
nor U12906 (N_12906,N_7585,N_9322);
xor U12907 (N_12907,N_6566,N_7931);
nor U12908 (N_12908,N_6438,N_7965);
or U12909 (N_12909,N_6199,N_9250);
or U12910 (N_12910,N_6544,N_5895);
nand U12911 (N_12911,N_6859,N_8218);
or U12912 (N_12912,N_6446,N_6637);
nor U12913 (N_12913,N_7232,N_7429);
nand U12914 (N_12914,N_8846,N_9019);
and U12915 (N_12915,N_7873,N_6647);
and U12916 (N_12916,N_8926,N_7315);
nor U12917 (N_12917,N_6975,N_9809);
nor U12918 (N_12918,N_6376,N_9805);
nor U12919 (N_12919,N_7584,N_5946);
nor U12920 (N_12920,N_5283,N_5259);
or U12921 (N_12921,N_6657,N_7972);
nor U12922 (N_12922,N_8374,N_5971);
and U12923 (N_12923,N_8706,N_5968);
nand U12924 (N_12924,N_8867,N_7757);
and U12925 (N_12925,N_6407,N_6301);
nand U12926 (N_12926,N_6155,N_8595);
nand U12927 (N_12927,N_7834,N_8521);
and U12928 (N_12928,N_9171,N_8732);
or U12929 (N_12929,N_8214,N_6561);
and U12930 (N_12930,N_7130,N_7325);
nor U12931 (N_12931,N_6532,N_8421);
and U12932 (N_12932,N_5529,N_8450);
or U12933 (N_12933,N_9651,N_5288);
nand U12934 (N_12934,N_5203,N_6276);
or U12935 (N_12935,N_7854,N_8803);
nor U12936 (N_12936,N_9867,N_9475);
nand U12937 (N_12937,N_5021,N_5442);
nor U12938 (N_12938,N_8883,N_6141);
nor U12939 (N_12939,N_9822,N_5602);
and U12940 (N_12940,N_5091,N_6379);
or U12941 (N_12941,N_9389,N_9082);
nor U12942 (N_12942,N_7321,N_7060);
nor U12943 (N_12943,N_6632,N_6681);
and U12944 (N_12944,N_7066,N_8804);
nand U12945 (N_12945,N_7441,N_6921);
and U12946 (N_12946,N_8422,N_5407);
nand U12947 (N_12947,N_6531,N_5194);
and U12948 (N_12948,N_6311,N_5926);
and U12949 (N_12949,N_8889,N_9453);
xnor U12950 (N_12950,N_9721,N_5283);
nand U12951 (N_12951,N_8451,N_5011);
nor U12952 (N_12952,N_9515,N_9343);
or U12953 (N_12953,N_9075,N_8433);
nor U12954 (N_12954,N_7905,N_9020);
nor U12955 (N_12955,N_9307,N_9456);
nand U12956 (N_12956,N_9209,N_6685);
nand U12957 (N_12957,N_6854,N_6687);
or U12958 (N_12958,N_6134,N_7475);
nand U12959 (N_12959,N_5714,N_5282);
and U12960 (N_12960,N_6393,N_5701);
xnor U12961 (N_12961,N_8930,N_5613);
nor U12962 (N_12962,N_6789,N_6651);
or U12963 (N_12963,N_6166,N_5067);
xor U12964 (N_12964,N_7040,N_5939);
or U12965 (N_12965,N_8916,N_6136);
and U12966 (N_12966,N_8097,N_6058);
nand U12967 (N_12967,N_8237,N_5437);
nand U12968 (N_12968,N_8540,N_5472);
nand U12969 (N_12969,N_8844,N_8008);
nor U12970 (N_12970,N_7407,N_9493);
or U12971 (N_12971,N_7795,N_6247);
or U12972 (N_12972,N_8679,N_9773);
or U12973 (N_12973,N_8615,N_9461);
nor U12974 (N_12974,N_6288,N_5445);
nor U12975 (N_12975,N_7870,N_5358);
xor U12976 (N_12976,N_8174,N_8237);
or U12977 (N_12977,N_7445,N_9145);
nand U12978 (N_12978,N_7072,N_9999);
nor U12979 (N_12979,N_8986,N_5967);
and U12980 (N_12980,N_5561,N_9485);
nand U12981 (N_12981,N_8865,N_7175);
nor U12982 (N_12982,N_5499,N_7805);
nor U12983 (N_12983,N_9907,N_9604);
and U12984 (N_12984,N_7099,N_5406);
and U12985 (N_12985,N_5099,N_7548);
nor U12986 (N_12986,N_8157,N_8924);
nand U12987 (N_12987,N_7592,N_5506);
and U12988 (N_12988,N_5376,N_9881);
nand U12989 (N_12989,N_6598,N_6697);
or U12990 (N_12990,N_9365,N_6492);
nand U12991 (N_12991,N_6194,N_6292);
or U12992 (N_12992,N_8536,N_5979);
and U12993 (N_12993,N_8383,N_8977);
and U12994 (N_12994,N_5820,N_6841);
or U12995 (N_12995,N_8751,N_6376);
nand U12996 (N_12996,N_7785,N_8409);
nor U12997 (N_12997,N_8373,N_8516);
xnor U12998 (N_12998,N_6911,N_5169);
and U12999 (N_12999,N_8462,N_9923);
or U13000 (N_13000,N_6640,N_7712);
nor U13001 (N_13001,N_9999,N_6443);
nand U13002 (N_13002,N_7483,N_9688);
nor U13003 (N_13003,N_9614,N_5910);
and U13004 (N_13004,N_7468,N_6391);
and U13005 (N_13005,N_7006,N_6785);
or U13006 (N_13006,N_6697,N_7920);
nand U13007 (N_13007,N_9203,N_8111);
or U13008 (N_13008,N_6888,N_8242);
and U13009 (N_13009,N_7915,N_8165);
xor U13010 (N_13010,N_9081,N_6018);
nand U13011 (N_13011,N_9684,N_6362);
or U13012 (N_13012,N_5368,N_9657);
or U13013 (N_13013,N_6889,N_7412);
nand U13014 (N_13014,N_5109,N_6558);
and U13015 (N_13015,N_7880,N_8102);
and U13016 (N_13016,N_8760,N_6008);
nor U13017 (N_13017,N_7186,N_7145);
nor U13018 (N_13018,N_9598,N_9013);
and U13019 (N_13019,N_8014,N_9985);
xor U13020 (N_13020,N_8989,N_6869);
or U13021 (N_13021,N_5955,N_5028);
or U13022 (N_13022,N_6900,N_6016);
or U13023 (N_13023,N_5051,N_9538);
nor U13024 (N_13024,N_9861,N_8542);
or U13025 (N_13025,N_7167,N_9843);
xor U13026 (N_13026,N_7019,N_7040);
or U13027 (N_13027,N_6404,N_7762);
or U13028 (N_13028,N_6270,N_7298);
or U13029 (N_13029,N_6546,N_8800);
and U13030 (N_13030,N_5346,N_5672);
or U13031 (N_13031,N_5690,N_7527);
xnor U13032 (N_13032,N_6411,N_9390);
or U13033 (N_13033,N_9842,N_8583);
nand U13034 (N_13034,N_9799,N_6553);
and U13035 (N_13035,N_6512,N_8892);
nor U13036 (N_13036,N_7440,N_7150);
nand U13037 (N_13037,N_9921,N_8954);
nor U13038 (N_13038,N_9674,N_6408);
nand U13039 (N_13039,N_6142,N_8318);
and U13040 (N_13040,N_5515,N_6914);
xor U13041 (N_13041,N_8298,N_8648);
nor U13042 (N_13042,N_7640,N_8159);
or U13043 (N_13043,N_5932,N_6520);
and U13044 (N_13044,N_5040,N_6213);
nand U13045 (N_13045,N_5163,N_7321);
and U13046 (N_13046,N_5721,N_8485);
nand U13047 (N_13047,N_6151,N_8906);
nor U13048 (N_13048,N_5143,N_6131);
nand U13049 (N_13049,N_9123,N_6280);
nor U13050 (N_13050,N_9144,N_8065);
and U13051 (N_13051,N_8454,N_6199);
or U13052 (N_13052,N_7528,N_5235);
nand U13053 (N_13053,N_9013,N_9561);
nand U13054 (N_13054,N_9353,N_5283);
or U13055 (N_13055,N_6049,N_9683);
xnor U13056 (N_13056,N_5830,N_8426);
or U13057 (N_13057,N_7158,N_9638);
and U13058 (N_13058,N_9032,N_9620);
and U13059 (N_13059,N_5630,N_6686);
nand U13060 (N_13060,N_5357,N_6716);
and U13061 (N_13061,N_8470,N_8204);
or U13062 (N_13062,N_8728,N_8997);
or U13063 (N_13063,N_7962,N_9911);
or U13064 (N_13064,N_5708,N_8703);
xor U13065 (N_13065,N_9196,N_5709);
nand U13066 (N_13066,N_9223,N_5366);
xnor U13067 (N_13067,N_9053,N_9543);
xor U13068 (N_13068,N_9897,N_9106);
nand U13069 (N_13069,N_9842,N_6216);
and U13070 (N_13070,N_9686,N_5883);
and U13071 (N_13071,N_6981,N_5695);
xnor U13072 (N_13072,N_9113,N_9529);
and U13073 (N_13073,N_5382,N_8935);
nand U13074 (N_13074,N_9736,N_7171);
nor U13075 (N_13075,N_7535,N_9214);
nand U13076 (N_13076,N_7710,N_5879);
nor U13077 (N_13077,N_8755,N_8300);
or U13078 (N_13078,N_8062,N_9331);
or U13079 (N_13079,N_6913,N_8421);
nand U13080 (N_13080,N_7814,N_6977);
or U13081 (N_13081,N_5332,N_5537);
xor U13082 (N_13082,N_6184,N_7487);
nor U13083 (N_13083,N_6750,N_7263);
nor U13084 (N_13084,N_7382,N_5465);
nor U13085 (N_13085,N_6490,N_7666);
nor U13086 (N_13086,N_8008,N_9010);
nand U13087 (N_13087,N_9603,N_5339);
nand U13088 (N_13088,N_9032,N_7126);
or U13089 (N_13089,N_7366,N_5786);
nand U13090 (N_13090,N_9771,N_9285);
nand U13091 (N_13091,N_8594,N_6603);
and U13092 (N_13092,N_6437,N_5136);
and U13093 (N_13093,N_6386,N_6753);
nor U13094 (N_13094,N_6888,N_7908);
and U13095 (N_13095,N_8337,N_9173);
nand U13096 (N_13096,N_8963,N_7498);
xnor U13097 (N_13097,N_7258,N_5518);
or U13098 (N_13098,N_7480,N_7721);
and U13099 (N_13099,N_5872,N_7548);
nand U13100 (N_13100,N_6500,N_8775);
nor U13101 (N_13101,N_6170,N_8363);
nand U13102 (N_13102,N_7661,N_9311);
and U13103 (N_13103,N_5211,N_9345);
or U13104 (N_13104,N_5071,N_7581);
and U13105 (N_13105,N_5271,N_7856);
xnor U13106 (N_13106,N_5711,N_8813);
and U13107 (N_13107,N_8808,N_9528);
and U13108 (N_13108,N_6375,N_6685);
or U13109 (N_13109,N_8108,N_7305);
nor U13110 (N_13110,N_8197,N_8730);
xnor U13111 (N_13111,N_9138,N_8367);
or U13112 (N_13112,N_6342,N_7497);
nand U13113 (N_13113,N_9207,N_6644);
or U13114 (N_13114,N_8957,N_7706);
xnor U13115 (N_13115,N_8720,N_6728);
or U13116 (N_13116,N_5385,N_7826);
nor U13117 (N_13117,N_7326,N_8650);
and U13118 (N_13118,N_9851,N_9424);
nand U13119 (N_13119,N_6359,N_6445);
or U13120 (N_13120,N_6465,N_6766);
or U13121 (N_13121,N_7388,N_6220);
or U13122 (N_13122,N_8367,N_9194);
nor U13123 (N_13123,N_9234,N_7285);
nor U13124 (N_13124,N_6203,N_9203);
or U13125 (N_13125,N_9783,N_5187);
nor U13126 (N_13126,N_8595,N_6005);
or U13127 (N_13127,N_9299,N_7540);
xnor U13128 (N_13128,N_9933,N_9559);
or U13129 (N_13129,N_7939,N_7336);
xor U13130 (N_13130,N_6518,N_6138);
xnor U13131 (N_13131,N_6557,N_5901);
nor U13132 (N_13132,N_7637,N_9431);
nand U13133 (N_13133,N_9326,N_5462);
nand U13134 (N_13134,N_9136,N_5771);
and U13135 (N_13135,N_5271,N_6083);
or U13136 (N_13136,N_8723,N_5611);
and U13137 (N_13137,N_5761,N_9497);
xor U13138 (N_13138,N_5879,N_7240);
or U13139 (N_13139,N_7268,N_6664);
and U13140 (N_13140,N_6747,N_7410);
nor U13141 (N_13141,N_8286,N_6190);
or U13142 (N_13142,N_6908,N_6966);
xor U13143 (N_13143,N_6814,N_9499);
and U13144 (N_13144,N_9621,N_8057);
or U13145 (N_13145,N_5486,N_8073);
nand U13146 (N_13146,N_6668,N_7857);
nand U13147 (N_13147,N_6127,N_5606);
nand U13148 (N_13148,N_7123,N_5345);
and U13149 (N_13149,N_5386,N_8419);
nand U13150 (N_13150,N_5936,N_9745);
nand U13151 (N_13151,N_9405,N_8065);
nand U13152 (N_13152,N_7115,N_9311);
and U13153 (N_13153,N_7689,N_7493);
and U13154 (N_13154,N_5443,N_6633);
or U13155 (N_13155,N_8831,N_8111);
or U13156 (N_13156,N_7589,N_6408);
nor U13157 (N_13157,N_9456,N_6925);
nand U13158 (N_13158,N_9386,N_7798);
nand U13159 (N_13159,N_9811,N_5240);
nor U13160 (N_13160,N_6525,N_6900);
nor U13161 (N_13161,N_8850,N_6737);
or U13162 (N_13162,N_7746,N_8179);
nand U13163 (N_13163,N_6004,N_9209);
nor U13164 (N_13164,N_6353,N_9470);
nand U13165 (N_13165,N_6059,N_8441);
nor U13166 (N_13166,N_7037,N_6215);
nand U13167 (N_13167,N_5030,N_8474);
and U13168 (N_13168,N_5185,N_7088);
nand U13169 (N_13169,N_5475,N_7388);
or U13170 (N_13170,N_7224,N_6099);
or U13171 (N_13171,N_9635,N_9986);
or U13172 (N_13172,N_8642,N_8731);
nor U13173 (N_13173,N_7147,N_5481);
nand U13174 (N_13174,N_9905,N_8184);
nor U13175 (N_13175,N_5484,N_7853);
and U13176 (N_13176,N_8966,N_8249);
or U13177 (N_13177,N_8727,N_9029);
and U13178 (N_13178,N_6144,N_8509);
nand U13179 (N_13179,N_7352,N_7599);
and U13180 (N_13180,N_6041,N_8966);
xnor U13181 (N_13181,N_5400,N_8897);
or U13182 (N_13182,N_5989,N_8075);
nor U13183 (N_13183,N_6977,N_5275);
and U13184 (N_13184,N_7060,N_9748);
nor U13185 (N_13185,N_9436,N_9182);
and U13186 (N_13186,N_6240,N_8516);
nor U13187 (N_13187,N_7466,N_5618);
and U13188 (N_13188,N_8942,N_9554);
nand U13189 (N_13189,N_8040,N_9027);
xnor U13190 (N_13190,N_7864,N_8180);
nand U13191 (N_13191,N_7276,N_9181);
or U13192 (N_13192,N_7488,N_9802);
and U13193 (N_13193,N_9246,N_6200);
and U13194 (N_13194,N_5093,N_8682);
nand U13195 (N_13195,N_6620,N_5291);
or U13196 (N_13196,N_9471,N_9845);
nor U13197 (N_13197,N_7763,N_9076);
nand U13198 (N_13198,N_5041,N_5948);
and U13199 (N_13199,N_5562,N_8077);
and U13200 (N_13200,N_8890,N_5685);
nand U13201 (N_13201,N_6142,N_7692);
and U13202 (N_13202,N_6904,N_7293);
nor U13203 (N_13203,N_6071,N_9122);
xnor U13204 (N_13204,N_5398,N_6994);
nand U13205 (N_13205,N_6959,N_5878);
or U13206 (N_13206,N_6912,N_7247);
or U13207 (N_13207,N_8491,N_7864);
or U13208 (N_13208,N_6793,N_7168);
and U13209 (N_13209,N_8146,N_8607);
nor U13210 (N_13210,N_7382,N_5677);
and U13211 (N_13211,N_8836,N_9300);
nor U13212 (N_13212,N_8794,N_9422);
nand U13213 (N_13213,N_7986,N_6190);
nand U13214 (N_13214,N_7391,N_7229);
or U13215 (N_13215,N_9262,N_6677);
or U13216 (N_13216,N_5358,N_7981);
and U13217 (N_13217,N_8899,N_8662);
and U13218 (N_13218,N_9008,N_6002);
and U13219 (N_13219,N_9387,N_9610);
nor U13220 (N_13220,N_6932,N_9443);
and U13221 (N_13221,N_5818,N_9261);
nor U13222 (N_13222,N_5092,N_6671);
and U13223 (N_13223,N_6462,N_6484);
nor U13224 (N_13224,N_9146,N_8296);
and U13225 (N_13225,N_7396,N_6935);
nand U13226 (N_13226,N_8721,N_5640);
and U13227 (N_13227,N_5806,N_8333);
nand U13228 (N_13228,N_6471,N_8619);
nand U13229 (N_13229,N_5595,N_7503);
and U13230 (N_13230,N_6993,N_8909);
and U13231 (N_13231,N_5662,N_6216);
and U13232 (N_13232,N_9128,N_7594);
nor U13233 (N_13233,N_6914,N_7491);
and U13234 (N_13234,N_6767,N_8591);
nand U13235 (N_13235,N_9155,N_7008);
nand U13236 (N_13236,N_8417,N_6364);
and U13237 (N_13237,N_8072,N_5467);
xor U13238 (N_13238,N_8312,N_6687);
and U13239 (N_13239,N_7650,N_7553);
xor U13240 (N_13240,N_8698,N_7210);
or U13241 (N_13241,N_5379,N_6228);
nor U13242 (N_13242,N_5494,N_6936);
nand U13243 (N_13243,N_8265,N_8145);
nand U13244 (N_13244,N_6629,N_5328);
and U13245 (N_13245,N_7802,N_9227);
or U13246 (N_13246,N_8631,N_5513);
or U13247 (N_13247,N_5866,N_5852);
nor U13248 (N_13248,N_7147,N_9189);
xnor U13249 (N_13249,N_7993,N_7444);
or U13250 (N_13250,N_5034,N_6341);
nor U13251 (N_13251,N_5030,N_7550);
nor U13252 (N_13252,N_7606,N_5554);
and U13253 (N_13253,N_5709,N_7054);
nand U13254 (N_13254,N_9601,N_5350);
nor U13255 (N_13255,N_9426,N_9504);
and U13256 (N_13256,N_8424,N_7473);
and U13257 (N_13257,N_6467,N_6545);
nor U13258 (N_13258,N_9223,N_8638);
nor U13259 (N_13259,N_6791,N_6505);
nor U13260 (N_13260,N_6524,N_6959);
nand U13261 (N_13261,N_7439,N_7077);
or U13262 (N_13262,N_5434,N_8507);
nor U13263 (N_13263,N_8551,N_7672);
and U13264 (N_13264,N_9521,N_7034);
nand U13265 (N_13265,N_8435,N_5962);
or U13266 (N_13266,N_6132,N_7566);
nor U13267 (N_13267,N_9674,N_8347);
or U13268 (N_13268,N_9873,N_7342);
or U13269 (N_13269,N_5515,N_7426);
and U13270 (N_13270,N_9875,N_5019);
nor U13271 (N_13271,N_6982,N_5387);
nor U13272 (N_13272,N_6769,N_6930);
nor U13273 (N_13273,N_7045,N_5251);
nand U13274 (N_13274,N_8455,N_8229);
or U13275 (N_13275,N_7014,N_8647);
and U13276 (N_13276,N_9205,N_5400);
and U13277 (N_13277,N_9648,N_5821);
or U13278 (N_13278,N_7042,N_7991);
and U13279 (N_13279,N_8158,N_9991);
xor U13280 (N_13280,N_9044,N_6879);
nand U13281 (N_13281,N_8071,N_8292);
nor U13282 (N_13282,N_7024,N_8398);
and U13283 (N_13283,N_7753,N_5402);
nor U13284 (N_13284,N_8552,N_9464);
nor U13285 (N_13285,N_6580,N_8230);
and U13286 (N_13286,N_6274,N_7424);
and U13287 (N_13287,N_6998,N_9182);
nor U13288 (N_13288,N_6790,N_9769);
nor U13289 (N_13289,N_5256,N_5476);
and U13290 (N_13290,N_5429,N_5484);
nor U13291 (N_13291,N_8640,N_7692);
nor U13292 (N_13292,N_8432,N_9125);
nand U13293 (N_13293,N_6498,N_6521);
xor U13294 (N_13294,N_5377,N_7841);
or U13295 (N_13295,N_7175,N_7771);
nor U13296 (N_13296,N_6995,N_6069);
or U13297 (N_13297,N_6652,N_6394);
nor U13298 (N_13298,N_6586,N_5674);
nor U13299 (N_13299,N_7332,N_5152);
and U13300 (N_13300,N_8938,N_5207);
or U13301 (N_13301,N_9993,N_5669);
or U13302 (N_13302,N_9049,N_5598);
and U13303 (N_13303,N_6413,N_7316);
nand U13304 (N_13304,N_5454,N_6599);
nand U13305 (N_13305,N_6004,N_8518);
and U13306 (N_13306,N_9554,N_9288);
and U13307 (N_13307,N_9918,N_7549);
and U13308 (N_13308,N_6152,N_7004);
nor U13309 (N_13309,N_9387,N_6372);
xnor U13310 (N_13310,N_8314,N_9513);
or U13311 (N_13311,N_9832,N_5687);
nor U13312 (N_13312,N_7974,N_9331);
nor U13313 (N_13313,N_7582,N_8743);
and U13314 (N_13314,N_5994,N_5287);
or U13315 (N_13315,N_6292,N_5104);
or U13316 (N_13316,N_9257,N_9733);
nor U13317 (N_13317,N_5951,N_5701);
nand U13318 (N_13318,N_5620,N_8372);
or U13319 (N_13319,N_5029,N_6484);
and U13320 (N_13320,N_7907,N_8382);
nand U13321 (N_13321,N_5525,N_5265);
nand U13322 (N_13322,N_8254,N_8463);
xor U13323 (N_13323,N_6309,N_5272);
or U13324 (N_13324,N_6500,N_6818);
nand U13325 (N_13325,N_6619,N_8917);
nor U13326 (N_13326,N_9015,N_8052);
and U13327 (N_13327,N_7845,N_7084);
xnor U13328 (N_13328,N_8938,N_7659);
nand U13329 (N_13329,N_5050,N_6275);
or U13330 (N_13330,N_8521,N_7252);
and U13331 (N_13331,N_5052,N_9622);
nor U13332 (N_13332,N_8532,N_9998);
nor U13333 (N_13333,N_5495,N_8719);
nand U13334 (N_13334,N_6340,N_7020);
xnor U13335 (N_13335,N_6568,N_6818);
and U13336 (N_13336,N_6924,N_8766);
or U13337 (N_13337,N_6324,N_8984);
nor U13338 (N_13338,N_8142,N_8083);
nand U13339 (N_13339,N_5133,N_9820);
or U13340 (N_13340,N_5919,N_7139);
and U13341 (N_13341,N_6324,N_7845);
nor U13342 (N_13342,N_9080,N_6636);
and U13343 (N_13343,N_9874,N_5698);
or U13344 (N_13344,N_9254,N_5801);
nor U13345 (N_13345,N_6621,N_9833);
nand U13346 (N_13346,N_7129,N_5776);
xnor U13347 (N_13347,N_9377,N_6539);
and U13348 (N_13348,N_8163,N_6416);
nand U13349 (N_13349,N_5126,N_9912);
and U13350 (N_13350,N_7640,N_9196);
nand U13351 (N_13351,N_9241,N_9731);
nor U13352 (N_13352,N_9203,N_5388);
nand U13353 (N_13353,N_5052,N_9143);
nand U13354 (N_13354,N_5113,N_8611);
and U13355 (N_13355,N_9968,N_5597);
xor U13356 (N_13356,N_5875,N_8640);
xnor U13357 (N_13357,N_5463,N_8886);
nor U13358 (N_13358,N_8198,N_8808);
or U13359 (N_13359,N_6485,N_9902);
and U13360 (N_13360,N_7365,N_5267);
or U13361 (N_13361,N_6659,N_7991);
xor U13362 (N_13362,N_9088,N_5665);
nor U13363 (N_13363,N_7743,N_9067);
and U13364 (N_13364,N_6316,N_7382);
xor U13365 (N_13365,N_8007,N_6386);
nand U13366 (N_13366,N_6959,N_9960);
xor U13367 (N_13367,N_6178,N_8339);
or U13368 (N_13368,N_9633,N_5782);
and U13369 (N_13369,N_9814,N_9569);
or U13370 (N_13370,N_6759,N_5952);
nor U13371 (N_13371,N_6152,N_9571);
nor U13372 (N_13372,N_7161,N_5756);
nand U13373 (N_13373,N_9378,N_5593);
nand U13374 (N_13374,N_6309,N_8175);
nand U13375 (N_13375,N_9535,N_5249);
and U13376 (N_13376,N_5723,N_6278);
and U13377 (N_13377,N_6624,N_8003);
nor U13378 (N_13378,N_7877,N_6518);
xor U13379 (N_13379,N_7911,N_6363);
nand U13380 (N_13380,N_9625,N_7734);
or U13381 (N_13381,N_7319,N_6032);
nand U13382 (N_13382,N_6017,N_5417);
nor U13383 (N_13383,N_6160,N_8212);
or U13384 (N_13384,N_6396,N_9949);
nand U13385 (N_13385,N_7981,N_7100);
nand U13386 (N_13386,N_8932,N_9362);
xor U13387 (N_13387,N_6993,N_9960);
xor U13388 (N_13388,N_5602,N_5979);
and U13389 (N_13389,N_8829,N_5157);
or U13390 (N_13390,N_8307,N_9854);
and U13391 (N_13391,N_8458,N_9462);
and U13392 (N_13392,N_9630,N_5552);
nor U13393 (N_13393,N_7844,N_9088);
xor U13394 (N_13394,N_7972,N_7931);
nand U13395 (N_13395,N_5988,N_6563);
nand U13396 (N_13396,N_6402,N_7465);
nor U13397 (N_13397,N_6613,N_9500);
nand U13398 (N_13398,N_6718,N_5715);
xnor U13399 (N_13399,N_8912,N_5599);
nor U13400 (N_13400,N_9990,N_7721);
and U13401 (N_13401,N_9428,N_9775);
and U13402 (N_13402,N_5357,N_8799);
and U13403 (N_13403,N_6111,N_9189);
or U13404 (N_13404,N_8491,N_9283);
nor U13405 (N_13405,N_8988,N_9222);
nor U13406 (N_13406,N_8876,N_8370);
or U13407 (N_13407,N_5072,N_6455);
nor U13408 (N_13408,N_7098,N_6042);
and U13409 (N_13409,N_9838,N_5060);
nor U13410 (N_13410,N_9449,N_5376);
nor U13411 (N_13411,N_7183,N_9874);
and U13412 (N_13412,N_6074,N_8839);
nand U13413 (N_13413,N_7421,N_7414);
xor U13414 (N_13414,N_8141,N_7543);
and U13415 (N_13415,N_5157,N_6321);
and U13416 (N_13416,N_7291,N_7859);
or U13417 (N_13417,N_9024,N_6583);
and U13418 (N_13418,N_8801,N_9624);
and U13419 (N_13419,N_9521,N_8765);
nand U13420 (N_13420,N_7890,N_5883);
and U13421 (N_13421,N_9539,N_7587);
nand U13422 (N_13422,N_6750,N_7945);
and U13423 (N_13423,N_8585,N_7438);
or U13424 (N_13424,N_6626,N_5927);
nand U13425 (N_13425,N_7613,N_7376);
or U13426 (N_13426,N_5568,N_9286);
and U13427 (N_13427,N_8626,N_5132);
xnor U13428 (N_13428,N_7021,N_6027);
xnor U13429 (N_13429,N_9352,N_9314);
or U13430 (N_13430,N_5911,N_8699);
nor U13431 (N_13431,N_6210,N_6339);
and U13432 (N_13432,N_7361,N_7834);
nor U13433 (N_13433,N_8058,N_7827);
and U13434 (N_13434,N_8771,N_6290);
and U13435 (N_13435,N_8740,N_9610);
nand U13436 (N_13436,N_9303,N_5400);
nor U13437 (N_13437,N_5489,N_5411);
nand U13438 (N_13438,N_8131,N_5698);
nand U13439 (N_13439,N_5662,N_9942);
or U13440 (N_13440,N_8432,N_7512);
and U13441 (N_13441,N_8876,N_9747);
or U13442 (N_13442,N_7217,N_6794);
nor U13443 (N_13443,N_8088,N_8343);
nor U13444 (N_13444,N_5161,N_9668);
and U13445 (N_13445,N_8139,N_8719);
nor U13446 (N_13446,N_9825,N_8435);
or U13447 (N_13447,N_6556,N_8869);
and U13448 (N_13448,N_8057,N_6586);
or U13449 (N_13449,N_6529,N_9939);
or U13450 (N_13450,N_5415,N_8807);
and U13451 (N_13451,N_7919,N_7723);
and U13452 (N_13452,N_8338,N_7601);
nand U13453 (N_13453,N_8306,N_7728);
nand U13454 (N_13454,N_5027,N_9810);
xor U13455 (N_13455,N_9314,N_7286);
nand U13456 (N_13456,N_9994,N_9464);
xnor U13457 (N_13457,N_5592,N_7029);
xnor U13458 (N_13458,N_9978,N_7426);
and U13459 (N_13459,N_7981,N_7029);
nor U13460 (N_13460,N_9565,N_8838);
nor U13461 (N_13461,N_9659,N_8809);
and U13462 (N_13462,N_9406,N_6837);
nor U13463 (N_13463,N_9278,N_6907);
nor U13464 (N_13464,N_6421,N_7425);
and U13465 (N_13465,N_6012,N_5877);
nand U13466 (N_13466,N_9126,N_6647);
nand U13467 (N_13467,N_5970,N_9827);
nor U13468 (N_13468,N_7892,N_6892);
nor U13469 (N_13469,N_5215,N_9676);
and U13470 (N_13470,N_6238,N_6597);
nor U13471 (N_13471,N_5586,N_6343);
or U13472 (N_13472,N_8497,N_6800);
nand U13473 (N_13473,N_6450,N_9946);
and U13474 (N_13474,N_5186,N_5979);
and U13475 (N_13475,N_6356,N_7366);
nor U13476 (N_13476,N_9265,N_8704);
nand U13477 (N_13477,N_9011,N_6618);
or U13478 (N_13478,N_8970,N_9274);
nand U13479 (N_13479,N_6074,N_8491);
nor U13480 (N_13480,N_9060,N_7954);
nand U13481 (N_13481,N_5352,N_5773);
and U13482 (N_13482,N_6430,N_6353);
and U13483 (N_13483,N_5525,N_9288);
and U13484 (N_13484,N_7449,N_5177);
nand U13485 (N_13485,N_5399,N_6970);
or U13486 (N_13486,N_6551,N_5709);
and U13487 (N_13487,N_6358,N_9307);
and U13488 (N_13488,N_7569,N_9527);
nor U13489 (N_13489,N_8675,N_9605);
nand U13490 (N_13490,N_6771,N_6367);
xnor U13491 (N_13491,N_9617,N_7010);
nor U13492 (N_13492,N_7696,N_9324);
nor U13493 (N_13493,N_9563,N_8278);
or U13494 (N_13494,N_7691,N_7599);
nor U13495 (N_13495,N_9387,N_8850);
or U13496 (N_13496,N_7329,N_8889);
or U13497 (N_13497,N_8396,N_6632);
nor U13498 (N_13498,N_9482,N_5797);
nor U13499 (N_13499,N_5714,N_7135);
nor U13500 (N_13500,N_6596,N_8862);
and U13501 (N_13501,N_7657,N_5167);
nand U13502 (N_13502,N_6667,N_9144);
nor U13503 (N_13503,N_9722,N_9046);
nand U13504 (N_13504,N_8960,N_8817);
xnor U13505 (N_13505,N_6020,N_7290);
nand U13506 (N_13506,N_6968,N_5854);
and U13507 (N_13507,N_8950,N_8549);
or U13508 (N_13508,N_7529,N_8454);
nand U13509 (N_13509,N_5418,N_9497);
nand U13510 (N_13510,N_5995,N_9142);
nor U13511 (N_13511,N_7214,N_6977);
nand U13512 (N_13512,N_9595,N_6233);
and U13513 (N_13513,N_6284,N_9872);
nand U13514 (N_13514,N_7521,N_5991);
or U13515 (N_13515,N_5395,N_6130);
and U13516 (N_13516,N_9799,N_8915);
and U13517 (N_13517,N_9724,N_9711);
and U13518 (N_13518,N_6912,N_8854);
nor U13519 (N_13519,N_8607,N_7870);
and U13520 (N_13520,N_9039,N_8149);
nor U13521 (N_13521,N_5328,N_9641);
nor U13522 (N_13522,N_9457,N_8941);
nand U13523 (N_13523,N_9331,N_5215);
nor U13524 (N_13524,N_5990,N_6692);
nor U13525 (N_13525,N_5610,N_5612);
and U13526 (N_13526,N_6047,N_6355);
xor U13527 (N_13527,N_9585,N_7834);
and U13528 (N_13528,N_5655,N_6284);
xor U13529 (N_13529,N_7958,N_9442);
nand U13530 (N_13530,N_5065,N_8683);
and U13531 (N_13531,N_7910,N_6944);
nor U13532 (N_13532,N_6105,N_7170);
nand U13533 (N_13533,N_9532,N_8088);
or U13534 (N_13534,N_5160,N_7287);
nor U13535 (N_13535,N_8311,N_7316);
or U13536 (N_13536,N_5099,N_9276);
nor U13537 (N_13537,N_5043,N_9334);
or U13538 (N_13538,N_7255,N_7445);
nand U13539 (N_13539,N_7852,N_5577);
or U13540 (N_13540,N_6423,N_5400);
nand U13541 (N_13541,N_7423,N_8113);
and U13542 (N_13542,N_6540,N_6254);
nor U13543 (N_13543,N_5351,N_8379);
nor U13544 (N_13544,N_7696,N_7664);
nand U13545 (N_13545,N_9412,N_9268);
nor U13546 (N_13546,N_6210,N_7273);
or U13547 (N_13547,N_6712,N_9972);
nand U13548 (N_13548,N_5392,N_6002);
nor U13549 (N_13549,N_7385,N_5133);
or U13550 (N_13550,N_7783,N_6565);
and U13551 (N_13551,N_6495,N_8728);
or U13552 (N_13552,N_6482,N_6941);
nor U13553 (N_13553,N_8641,N_9020);
xnor U13554 (N_13554,N_9809,N_9477);
or U13555 (N_13555,N_9887,N_5386);
nand U13556 (N_13556,N_7068,N_5738);
nand U13557 (N_13557,N_9638,N_7723);
or U13558 (N_13558,N_9459,N_7611);
nor U13559 (N_13559,N_9822,N_6209);
or U13560 (N_13560,N_6507,N_9388);
and U13561 (N_13561,N_6918,N_7810);
or U13562 (N_13562,N_7117,N_9022);
or U13563 (N_13563,N_7524,N_5607);
nor U13564 (N_13564,N_7745,N_6643);
nor U13565 (N_13565,N_5456,N_5854);
nor U13566 (N_13566,N_6025,N_7741);
nor U13567 (N_13567,N_6221,N_9024);
nand U13568 (N_13568,N_8687,N_6414);
and U13569 (N_13569,N_9515,N_7443);
nand U13570 (N_13570,N_8782,N_6326);
nand U13571 (N_13571,N_6706,N_8924);
xnor U13572 (N_13572,N_8019,N_8053);
xor U13573 (N_13573,N_5150,N_5062);
nand U13574 (N_13574,N_8728,N_8705);
xor U13575 (N_13575,N_5696,N_6760);
nand U13576 (N_13576,N_9551,N_9909);
nand U13577 (N_13577,N_8289,N_9126);
and U13578 (N_13578,N_6855,N_5024);
nor U13579 (N_13579,N_8895,N_7432);
and U13580 (N_13580,N_8088,N_6001);
nor U13581 (N_13581,N_6294,N_6191);
nor U13582 (N_13582,N_8134,N_6478);
nand U13583 (N_13583,N_5674,N_9546);
or U13584 (N_13584,N_8825,N_7901);
nor U13585 (N_13585,N_8602,N_9892);
nor U13586 (N_13586,N_6324,N_9582);
nand U13587 (N_13587,N_8599,N_7526);
and U13588 (N_13588,N_8760,N_9901);
nor U13589 (N_13589,N_9173,N_5822);
and U13590 (N_13590,N_6689,N_6272);
xor U13591 (N_13591,N_6912,N_8255);
and U13592 (N_13592,N_7659,N_7465);
nand U13593 (N_13593,N_5614,N_9390);
nor U13594 (N_13594,N_9538,N_7489);
and U13595 (N_13595,N_5808,N_6440);
nand U13596 (N_13596,N_6741,N_5009);
nor U13597 (N_13597,N_6063,N_8868);
nand U13598 (N_13598,N_9647,N_5446);
and U13599 (N_13599,N_6597,N_5892);
nand U13600 (N_13600,N_8158,N_7947);
nor U13601 (N_13601,N_5335,N_7340);
and U13602 (N_13602,N_6078,N_9023);
or U13603 (N_13603,N_7653,N_9622);
xor U13604 (N_13604,N_6561,N_5300);
nor U13605 (N_13605,N_8496,N_9011);
nor U13606 (N_13606,N_5852,N_6689);
nand U13607 (N_13607,N_9622,N_9839);
and U13608 (N_13608,N_9209,N_7660);
or U13609 (N_13609,N_9836,N_9538);
nand U13610 (N_13610,N_8418,N_6360);
nor U13611 (N_13611,N_8790,N_8077);
nor U13612 (N_13612,N_9423,N_9640);
xor U13613 (N_13613,N_6918,N_6546);
nor U13614 (N_13614,N_7182,N_5981);
nand U13615 (N_13615,N_6312,N_7486);
nor U13616 (N_13616,N_6711,N_6937);
or U13617 (N_13617,N_7510,N_9390);
nand U13618 (N_13618,N_5281,N_8379);
nor U13619 (N_13619,N_8601,N_7456);
or U13620 (N_13620,N_5753,N_8119);
nor U13621 (N_13621,N_8818,N_8413);
nand U13622 (N_13622,N_6452,N_5339);
nor U13623 (N_13623,N_8856,N_5102);
and U13624 (N_13624,N_5869,N_7770);
or U13625 (N_13625,N_9054,N_8267);
or U13626 (N_13626,N_6225,N_9281);
nand U13627 (N_13627,N_9357,N_7385);
xor U13628 (N_13628,N_6037,N_9665);
or U13629 (N_13629,N_7996,N_8399);
xnor U13630 (N_13630,N_7056,N_9098);
and U13631 (N_13631,N_8599,N_6126);
nor U13632 (N_13632,N_6437,N_9161);
or U13633 (N_13633,N_6308,N_5237);
or U13634 (N_13634,N_8258,N_8659);
nor U13635 (N_13635,N_6715,N_5011);
and U13636 (N_13636,N_6461,N_5273);
and U13637 (N_13637,N_8883,N_7407);
and U13638 (N_13638,N_5924,N_6342);
and U13639 (N_13639,N_9702,N_9446);
or U13640 (N_13640,N_9448,N_6576);
or U13641 (N_13641,N_9888,N_8161);
xor U13642 (N_13642,N_6108,N_7016);
xnor U13643 (N_13643,N_7093,N_8557);
nor U13644 (N_13644,N_9173,N_6910);
or U13645 (N_13645,N_5352,N_6338);
nand U13646 (N_13646,N_8212,N_9994);
or U13647 (N_13647,N_7018,N_5985);
or U13648 (N_13648,N_6027,N_9018);
nor U13649 (N_13649,N_6628,N_8169);
or U13650 (N_13650,N_5952,N_6104);
nand U13651 (N_13651,N_6159,N_6166);
nor U13652 (N_13652,N_5382,N_9677);
xnor U13653 (N_13653,N_6035,N_7385);
and U13654 (N_13654,N_9048,N_7781);
and U13655 (N_13655,N_9707,N_7725);
nor U13656 (N_13656,N_6636,N_6352);
and U13657 (N_13657,N_8829,N_6723);
or U13658 (N_13658,N_7662,N_6129);
nand U13659 (N_13659,N_6925,N_8464);
xor U13660 (N_13660,N_5008,N_8428);
nand U13661 (N_13661,N_6964,N_9457);
nor U13662 (N_13662,N_6821,N_7387);
nor U13663 (N_13663,N_6579,N_9963);
or U13664 (N_13664,N_9509,N_9604);
nand U13665 (N_13665,N_9737,N_7308);
xor U13666 (N_13666,N_7127,N_7476);
nand U13667 (N_13667,N_7684,N_5475);
and U13668 (N_13668,N_6123,N_7940);
xor U13669 (N_13669,N_7962,N_8387);
and U13670 (N_13670,N_7473,N_5433);
and U13671 (N_13671,N_5801,N_8216);
or U13672 (N_13672,N_8522,N_9962);
and U13673 (N_13673,N_7808,N_7771);
nor U13674 (N_13674,N_5509,N_8454);
nor U13675 (N_13675,N_9615,N_9713);
and U13676 (N_13676,N_9572,N_5626);
or U13677 (N_13677,N_7669,N_8354);
nor U13678 (N_13678,N_6579,N_6978);
nand U13679 (N_13679,N_5263,N_7521);
nor U13680 (N_13680,N_7908,N_7844);
and U13681 (N_13681,N_7945,N_6464);
or U13682 (N_13682,N_9138,N_8549);
or U13683 (N_13683,N_9515,N_7107);
xor U13684 (N_13684,N_5965,N_5894);
or U13685 (N_13685,N_8215,N_9716);
and U13686 (N_13686,N_9055,N_7811);
and U13687 (N_13687,N_5105,N_7303);
nor U13688 (N_13688,N_9063,N_5434);
and U13689 (N_13689,N_6521,N_6254);
nand U13690 (N_13690,N_9930,N_5358);
nor U13691 (N_13691,N_5998,N_5678);
nand U13692 (N_13692,N_6671,N_9849);
nor U13693 (N_13693,N_9202,N_6182);
nor U13694 (N_13694,N_6427,N_8396);
nor U13695 (N_13695,N_8883,N_6382);
nand U13696 (N_13696,N_8386,N_7684);
nand U13697 (N_13697,N_5544,N_9208);
xor U13698 (N_13698,N_6077,N_7245);
nand U13699 (N_13699,N_5266,N_5693);
and U13700 (N_13700,N_9105,N_8679);
nor U13701 (N_13701,N_7275,N_6003);
nor U13702 (N_13702,N_8027,N_5931);
and U13703 (N_13703,N_9120,N_5432);
or U13704 (N_13704,N_6510,N_5792);
xnor U13705 (N_13705,N_9498,N_6373);
nor U13706 (N_13706,N_7298,N_9127);
nor U13707 (N_13707,N_6495,N_6472);
or U13708 (N_13708,N_6560,N_9680);
nor U13709 (N_13709,N_9037,N_5618);
or U13710 (N_13710,N_5449,N_7658);
xnor U13711 (N_13711,N_7621,N_8789);
or U13712 (N_13712,N_8046,N_5203);
nand U13713 (N_13713,N_7509,N_8726);
nand U13714 (N_13714,N_6272,N_6056);
and U13715 (N_13715,N_7440,N_9682);
xnor U13716 (N_13716,N_7787,N_5958);
or U13717 (N_13717,N_9195,N_5689);
xor U13718 (N_13718,N_8636,N_5684);
and U13719 (N_13719,N_8463,N_8925);
nand U13720 (N_13720,N_6069,N_7372);
and U13721 (N_13721,N_6035,N_5467);
or U13722 (N_13722,N_8969,N_8236);
or U13723 (N_13723,N_7234,N_7096);
xor U13724 (N_13724,N_5059,N_8646);
nor U13725 (N_13725,N_6727,N_5372);
nor U13726 (N_13726,N_7857,N_8924);
or U13727 (N_13727,N_6679,N_6392);
or U13728 (N_13728,N_7947,N_8862);
nand U13729 (N_13729,N_8343,N_8852);
and U13730 (N_13730,N_5716,N_5399);
xor U13731 (N_13731,N_5250,N_7841);
nand U13732 (N_13732,N_7950,N_8687);
nand U13733 (N_13733,N_5468,N_5018);
nand U13734 (N_13734,N_7937,N_6909);
nor U13735 (N_13735,N_5742,N_6751);
or U13736 (N_13736,N_9129,N_9680);
nand U13737 (N_13737,N_9943,N_6313);
or U13738 (N_13738,N_8683,N_8000);
nand U13739 (N_13739,N_9013,N_5979);
nand U13740 (N_13740,N_7788,N_5447);
xnor U13741 (N_13741,N_9709,N_6074);
nor U13742 (N_13742,N_9886,N_7050);
nor U13743 (N_13743,N_5680,N_9960);
nand U13744 (N_13744,N_5079,N_8587);
and U13745 (N_13745,N_8350,N_7815);
nand U13746 (N_13746,N_9897,N_6394);
or U13747 (N_13747,N_6732,N_6770);
and U13748 (N_13748,N_9338,N_6042);
xor U13749 (N_13749,N_9300,N_5107);
nand U13750 (N_13750,N_8622,N_9847);
and U13751 (N_13751,N_5929,N_6121);
nand U13752 (N_13752,N_6698,N_5841);
nor U13753 (N_13753,N_6945,N_8064);
nand U13754 (N_13754,N_9612,N_6063);
nand U13755 (N_13755,N_9503,N_9084);
and U13756 (N_13756,N_7428,N_9355);
or U13757 (N_13757,N_5761,N_8547);
nor U13758 (N_13758,N_9661,N_7928);
nand U13759 (N_13759,N_6798,N_7841);
nand U13760 (N_13760,N_7838,N_5326);
or U13761 (N_13761,N_7561,N_6672);
and U13762 (N_13762,N_7296,N_6942);
or U13763 (N_13763,N_9051,N_8202);
or U13764 (N_13764,N_5055,N_9430);
or U13765 (N_13765,N_8734,N_8695);
and U13766 (N_13766,N_8234,N_9502);
nor U13767 (N_13767,N_6621,N_7857);
nor U13768 (N_13768,N_6995,N_6806);
nand U13769 (N_13769,N_6072,N_8059);
nor U13770 (N_13770,N_5965,N_9822);
nor U13771 (N_13771,N_6659,N_8726);
nor U13772 (N_13772,N_9331,N_7637);
or U13773 (N_13773,N_8878,N_8421);
or U13774 (N_13774,N_8387,N_9777);
nand U13775 (N_13775,N_5871,N_5203);
nor U13776 (N_13776,N_6476,N_9588);
nor U13777 (N_13777,N_5688,N_5344);
nand U13778 (N_13778,N_5749,N_5398);
and U13779 (N_13779,N_5280,N_7520);
nor U13780 (N_13780,N_8874,N_5322);
or U13781 (N_13781,N_8815,N_5089);
xnor U13782 (N_13782,N_5744,N_7708);
and U13783 (N_13783,N_8477,N_5904);
and U13784 (N_13784,N_9927,N_7909);
nor U13785 (N_13785,N_7773,N_6160);
nand U13786 (N_13786,N_6106,N_6467);
or U13787 (N_13787,N_6660,N_5369);
nand U13788 (N_13788,N_7571,N_9381);
and U13789 (N_13789,N_9261,N_8087);
nor U13790 (N_13790,N_5608,N_8364);
or U13791 (N_13791,N_6836,N_9354);
nand U13792 (N_13792,N_5738,N_5747);
and U13793 (N_13793,N_6878,N_6403);
or U13794 (N_13794,N_9271,N_5250);
or U13795 (N_13795,N_6387,N_7270);
xor U13796 (N_13796,N_5758,N_5494);
nand U13797 (N_13797,N_6341,N_9575);
nor U13798 (N_13798,N_7459,N_5753);
nand U13799 (N_13799,N_9710,N_9886);
xor U13800 (N_13800,N_8626,N_6746);
nor U13801 (N_13801,N_5436,N_5255);
nor U13802 (N_13802,N_7660,N_9677);
and U13803 (N_13803,N_5437,N_6488);
nand U13804 (N_13804,N_6952,N_7616);
and U13805 (N_13805,N_6485,N_7135);
xnor U13806 (N_13806,N_7744,N_8743);
xnor U13807 (N_13807,N_9129,N_8066);
or U13808 (N_13808,N_9905,N_9822);
and U13809 (N_13809,N_6827,N_7861);
xnor U13810 (N_13810,N_7449,N_5899);
and U13811 (N_13811,N_9514,N_5120);
xnor U13812 (N_13812,N_7311,N_6718);
nand U13813 (N_13813,N_7393,N_5606);
nand U13814 (N_13814,N_6593,N_5544);
xnor U13815 (N_13815,N_7599,N_7296);
xnor U13816 (N_13816,N_8608,N_8610);
nand U13817 (N_13817,N_5750,N_5729);
or U13818 (N_13818,N_6960,N_7013);
or U13819 (N_13819,N_8243,N_7195);
nand U13820 (N_13820,N_8245,N_5098);
nand U13821 (N_13821,N_8636,N_7985);
nor U13822 (N_13822,N_9098,N_7403);
nor U13823 (N_13823,N_9143,N_8611);
nor U13824 (N_13824,N_5284,N_5135);
nor U13825 (N_13825,N_5814,N_7977);
nor U13826 (N_13826,N_9235,N_8888);
or U13827 (N_13827,N_6427,N_7058);
and U13828 (N_13828,N_9295,N_8384);
nand U13829 (N_13829,N_5007,N_7373);
or U13830 (N_13830,N_7203,N_7027);
nand U13831 (N_13831,N_9116,N_7345);
nor U13832 (N_13832,N_6172,N_8146);
and U13833 (N_13833,N_9381,N_6742);
nor U13834 (N_13834,N_8105,N_9417);
nand U13835 (N_13835,N_8206,N_5222);
and U13836 (N_13836,N_9966,N_5417);
or U13837 (N_13837,N_7326,N_6252);
and U13838 (N_13838,N_9101,N_6053);
xnor U13839 (N_13839,N_6785,N_7628);
or U13840 (N_13840,N_8933,N_5119);
nand U13841 (N_13841,N_6091,N_8947);
nor U13842 (N_13842,N_9862,N_8946);
xnor U13843 (N_13843,N_8209,N_7900);
nand U13844 (N_13844,N_7685,N_9337);
nor U13845 (N_13845,N_6853,N_5747);
nand U13846 (N_13846,N_6045,N_7309);
or U13847 (N_13847,N_6495,N_6742);
or U13848 (N_13848,N_5526,N_8818);
and U13849 (N_13849,N_6697,N_9649);
nand U13850 (N_13850,N_8121,N_7369);
or U13851 (N_13851,N_7164,N_5408);
nand U13852 (N_13852,N_6773,N_5075);
and U13853 (N_13853,N_5804,N_8485);
nor U13854 (N_13854,N_5945,N_7536);
nand U13855 (N_13855,N_8352,N_5527);
and U13856 (N_13856,N_9348,N_5309);
or U13857 (N_13857,N_5667,N_9303);
nand U13858 (N_13858,N_6653,N_7361);
nor U13859 (N_13859,N_9590,N_9207);
or U13860 (N_13860,N_9949,N_8037);
or U13861 (N_13861,N_8042,N_8276);
and U13862 (N_13862,N_6794,N_6000);
and U13863 (N_13863,N_9367,N_9089);
nand U13864 (N_13864,N_5143,N_5471);
or U13865 (N_13865,N_9843,N_6497);
nor U13866 (N_13866,N_8516,N_5170);
and U13867 (N_13867,N_7274,N_9335);
or U13868 (N_13868,N_5247,N_7214);
nor U13869 (N_13869,N_6590,N_7914);
and U13870 (N_13870,N_6679,N_5157);
xnor U13871 (N_13871,N_9098,N_9883);
nand U13872 (N_13872,N_8771,N_9993);
or U13873 (N_13873,N_7941,N_8660);
and U13874 (N_13874,N_9064,N_9506);
and U13875 (N_13875,N_7730,N_8670);
nand U13876 (N_13876,N_5263,N_5713);
nor U13877 (N_13877,N_6949,N_5674);
or U13878 (N_13878,N_7926,N_8103);
nor U13879 (N_13879,N_9486,N_6030);
nand U13880 (N_13880,N_5798,N_9046);
nor U13881 (N_13881,N_8711,N_8255);
nor U13882 (N_13882,N_7170,N_7177);
and U13883 (N_13883,N_9219,N_9290);
nor U13884 (N_13884,N_6674,N_5227);
and U13885 (N_13885,N_7914,N_5972);
and U13886 (N_13886,N_5572,N_5317);
or U13887 (N_13887,N_5985,N_8417);
nor U13888 (N_13888,N_6020,N_8047);
and U13889 (N_13889,N_5004,N_8331);
or U13890 (N_13890,N_9479,N_7280);
or U13891 (N_13891,N_9609,N_7440);
nor U13892 (N_13892,N_5355,N_5816);
xnor U13893 (N_13893,N_9952,N_8020);
or U13894 (N_13894,N_5226,N_9536);
or U13895 (N_13895,N_9968,N_7777);
nor U13896 (N_13896,N_6820,N_8684);
xor U13897 (N_13897,N_6085,N_7766);
and U13898 (N_13898,N_9112,N_5154);
and U13899 (N_13899,N_6037,N_6283);
or U13900 (N_13900,N_7768,N_9901);
xor U13901 (N_13901,N_8413,N_9822);
or U13902 (N_13902,N_7776,N_9091);
or U13903 (N_13903,N_9828,N_8757);
nand U13904 (N_13904,N_6263,N_9784);
nand U13905 (N_13905,N_8420,N_8456);
xnor U13906 (N_13906,N_9702,N_5780);
nor U13907 (N_13907,N_6259,N_9688);
or U13908 (N_13908,N_5553,N_5671);
nor U13909 (N_13909,N_9838,N_9898);
or U13910 (N_13910,N_5254,N_9146);
or U13911 (N_13911,N_9829,N_8916);
nor U13912 (N_13912,N_9804,N_6658);
or U13913 (N_13913,N_8380,N_9097);
and U13914 (N_13914,N_8051,N_8921);
and U13915 (N_13915,N_9284,N_5897);
nand U13916 (N_13916,N_9797,N_7796);
nor U13917 (N_13917,N_7989,N_8657);
and U13918 (N_13918,N_8929,N_7578);
or U13919 (N_13919,N_9937,N_8662);
nand U13920 (N_13920,N_5123,N_6143);
nand U13921 (N_13921,N_5612,N_5248);
nand U13922 (N_13922,N_9730,N_6097);
nand U13923 (N_13923,N_7588,N_8450);
and U13924 (N_13924,N_8985,N_7156);
or U13925 (N_13925,N_8555,N_7477);
or U13926 (N_13926,N_9335,N_6564);
nand U13927 (N_13927,N_7824,N_7109);
xnor U13928 (N_13928,N_5233,N_7476);
nand U13929 (N_13929,N_9947,N_8338);
nor U13930 (N_13930,N_7694,N_9970);
or U13931 (N_13931,N_8080,N_7660);
nand U13932 (N_13932,N_7371,N_8201);
nand U13933 (N_13933,N_5520,N_6740);
nor U13934 (N_13934,N_9669,N_6227);
or U13935 (N_13935,N_7627,N_7834);
nor U13936 (N_13936,N_6855,N_8051);
nor U13937 (N_13937,N_8954,N_5036);
nand U13938 (N_13938,N_7488,N_9442);
nand U13939 (N_13939,N_9191,N_7131);
nor U13940 (N_13940,N_7741,N_9930);
and U13941 (N_13941,N_6781,N_6619);
nor U13942 (N_13942,N_9605,N_5839);
nand U13943 (N_13943,N_8801,N_8847);
or U13944 (N_13944,N_9062,N_7646);
nand U13945 (N_13945,N_9800,N_7935);
or U13946 (N_13946,N_8167,N_7170);
nand U13947 (N_13947,N_9891,N_8946);
xor U13948 (N_13948,N_9301,N_5640);
nor U13949 (N_13949,N_6820,N_7571);
nand U13950 (N_13950,N_7217,N_7488);
nand U13951 (N_13951,N_7144,N_7892);
and U13952 (N_13952,N_6898,N_5907);
xnor U13953 (N_13953,N_5534,N_7016);
nor U13954 (N_13954,N_7935,N_8066);
nand U13955 (N_13955,N_9765,N_9986);
and U13956 (N_13956,N_6629,N_5093);
and U13957 (N_13957,N_8787,N_7488);
and U13958 (N_13958,N_9870,N_8896);
and U13959 (N_13959,N_9585,N_9597);
and U13960 (N_13960,N_6656,N_9099);
xnor U13961 (N_13961,N_8873,N_5690);
nor U13962 (N_13962,N_6492,N_8997);
or U13963 (N_13963,N_5682,N_7008);
nand U13964 (N_13964,N_5383,N_6146);
and U13965 (N_13965,N_7349,N_5205);
nand U13966 (N_13966,N_9561,N_9002);
nor U13967 (N_13967,N_8893,N_6967);
nor U13968 (N_13968,N_9575,N_8759);
or U13969 (N_13969,N_5953,N_8706);
nand U13970 (N_13970,N_7727,N_6908);
or U13971 (N_13971,N_7102,N_5411);
nor U13972 (N_13972,N_5693,N_7341);
and U13973 (N_13973,N_7986,N_8805);
and U13974 (N_13974,N_9325,N_6722);
or U13975 (N_13975,N_6218,N_5042);
and U13976 (N_13976,N_5619,N_8419);
nand U13977 (N_13977,N_5958,N_8191);
nand U13978 (N_13978,N_6026,N_8984);
nor U13979 (N_13979,N_8419,N_8978);
nand U13980 (N_13980,N_9477,N_9980);
or U13981 (N_13981,N_8328,N_8247);
nor U13982 (N_13982,N_5469,N_5863);
nand U13983 (N_13983,N_9461,N_5653);
nor U13984 (N_13984,N_8997,N_7862);
nor U13985 (N_13985,N_7531,N_9403);
and U13986 (N_13986,N_9766,N_5681);
nor U13987 (N_13987,N_5318,N_9056);
nand U13988 (N_13988,N_6668,N_7463);
nor U13989 (N_13989,N_9703,N_6546);
xor U13990 (N_13990,N_8950,N_6060);
or U13991 (N_13991,N_8237,N_8052);
and U13992 (N_13992,N_6113,N_5915);
nand U13993 (N_13993,N_7071,N_7358);
nand U13994 (N_13994,N_9436,N_5861);
nand U13995 (N_13995,N_5052,N_6669);
or U13996 (N_13996,N_9673,N_8811);
or U13997 (N_13997,N_5611,N_8405);
or U13998 (N_13998,N_7986,N_7914);
or U13999 (N_13999,N_5467,N_5469);
and U14000 (N_14000,N_5764,N_6768);
and U14001 (N_14001,N_8658,N_9283);
and U14002 (N_14002,N_9614,N_9879);
xnor U14003 (N_14003,N_9002,N_7313);
or U14004 (N_14004,N_7739,N_8740);
and U14005 (N_14005,N_8360,N_5776);
and U14006 (N_14006,N_6664,N_6661);
or U14007 (N_14007,N_9498,N_5286);
and U14008 (N_14008,N_7822,N_7453);
and U14009 (N_14009,N_5337,N_6411);
or U14010 (N_14010,N_5338,N_8399);
or U14011 (N_14011,N_8053,N_7551);
nor U14012 (N_14012,N_5734,N_7869);
nand U14013 (N_14013,N_5209,N_9933);
nor U14014 (N_14014,N_6094,N_6003);
xor U14015 (N_14015,N_7995,N_8127);
nor U14016 (N_14016,N_8207,N_7069);
nor U14017 (N_14017,N_6262,N_8871);
nand U14018 (N_14018,N_9861,N_7198);
nor U14019 (N_14019,N_6094,N_7647);
or U14020 (N_14020,N_8808,N_7563);
or U14021 (N_14021,N_5041,N_9325);
nor U14022 (N_14022,N_6359,N_5031);
nor U14023 (N_14023,N_5221,N_9312);
nor U14024 (N_14024,N_8206,N_9057);
or U14025 (N_14025,N_6404,N_9064);
nand U14026 (N_14026,N_9014,N_5230);
and U14027 (N_14027,N_9484,N_8830);
xnor U14028 (N_14028,N_6447,N_7979);
or U14029 (N_14029,N_9339,N_8725);
nand U14030 (N_14030,N_9394,N_5070);
or U14031 (N_14031,N_8698,N_8565);
nor U14032 (N_14032,N_5810,N_5920);
nand U14033 (N_14033,N_8423,N_9219);
nor U14034 (N_14034,N_8468,N_5862);
or U14035 (N_14035,N_5585,N_5253);
nor U14036 (N_14036,N_8912,N_7884);
nand U14037 (N_14037,N_6250,N_9542);
or U14038 (N_14038,N_5631,N_7006);
nand U14039 (N_14039,N_5177,N_9013);
nor U14040 (N_14040,N_5489,N_6763);
nor U14041 (N_14041,N_7904,N_5735);
nand U14042 (N_14042,N_5861,N_7869);
or U14043 (N_14043,N_7166,N_5860);
or U14044 (N_14044,N_8891,N_6621);
and U14045 (N_14045,N_8462,N_9560);
nor U14046 (N_14046,N_5336,N_5662);
or U14047 (N_14047,N_7962,N_7015);
or U14048 (N_14048,N_9154,N_7243);
or U14049 (N_14049,N_5713,N_6539);
or U14050 (N_14050,N_9577,N_8814);
or U14051 (N_14051,N_7945,N_5719);
and U14052 (N_14052,N_5372,N_9891);
and U14053 (N_14053,N_8882,N_8158);
or U14054 (N_14054,N_7404,N_7833);
and U14055 (N_14055,N_9993,N_6339);
nand U14056 (N_14056,N_8929,N_5176);
nand U14057 (N_14057,N_5081,N_8883);
or U14058 (N_14058,N_5371,N_5934);
nor U14059 (N_14059,N_8290,N_9783);
nand U14060 (N_14060,N_6478,N_7539);
and U14061 (N_14061,N_9623,N_9169);
nor U14062 (N_14062,N_7438,N_7778);
nor U14063 (N_14063,N_9518,N_6265);
nand U14064 (N_14064,N_5302,N_8704);
nor U14065 (N_14065,N_5650,N_8640);
and U14066 (N_14066,N_9355,N_7953);
nor U14067 (N_14067,N_8387,N_9076);
nand U14068 (N_14068,N_8022,N_8784);
or U14069 (N_14069,N_8891,N_5518);
nand U14070 (N_14070,N_7288,N_8092);
nor U14071 (N_14071,N_9268,N_6360);
nand U14072 (N_14072,N_9964,N_5052);
nor U14073 (N_14073,N_8604,N_9782);
or U14074 (N_14074,N_8645,N_7826);
and U14075 (N_14075,N_8895,N_6155);
nand U14076 (N_14076,N_7312,N_9903);
or U14077 (N_14077,N_9503,N_7029);
or U14078 (N_14078,N_7589,N_5186);
nor U14079 (N_14079,N_7900,N_6291);
nand U14080 (N_14080,N_9663,N_7113);
and U14081 (N_14081,N_5056,N_7982);
or U14082 (N_14082,N_5428,N_6316);
nor U14083 (N_14083,N_9365,N_5276);
nand U14084 (N_14084,N_8514,N_5789);
or U14085 (N_14085,N_8854,N_9539);
nand U14086 (N_14086,N_9525,N_9376);
nor U14087 (N_14087,N_5477,N_6990);
or U14088 (N_14088,N_8658,N_7160);
nand U14089 (N_14089,N_9848,N_5147);
nand U14090 (N_14090,N_6071,N_6925);
nor U14091 (N_14091,N_5639,N_9476);
or U14092 (N_14092,N_7083,N_7106);
or U14093 (N_14093,N_9529,N_6644);
and U14094 (N_14094,N_8209,N_7664);
and U14095 (N_14095,N_6983,N_6908);
nor U14096 (N_14096,N_6668,N_8133);
nor U14097 (N_14097,N_6708,N_8600);
nor U14098 (N_14098,N_6793,N_8986);
or U14099 (N_14099,N_9634,N_7455);
and U14100 (N_14100,N_9491,N_7630);
or U14101 (N_14101,N_7392,N_9004);
nand U14102 (N_14102,N_6702,N_9254);
nor U14103 (N_14103,N_7437,N_7558);
or U14104 (N_14104,N_8309,N_7727);
and U14105 (N_14105,N_8642,N_5247);
nand U14106 (N_14106,N_5172,N_6857);
and U14107 (N_14107,N_9297,N_9405);
nor U14108 (N_14108,N_5803,N_6664);
and U14109 (N_14109,N_9229,N_8307);
nand U14110 (N_14110,N_7078,N_8864);
or U14111 (N_14111,N_9912,N_6067);
nor U14112 (N_14112,N_6026,N_7194);
or U14113 (N_14113,N_7250,N_5322);
nand U14114 (N_14114,N_7183,N_8693);
nand U14115 (N_14115,N_6673,N_7794);
nand U14116 (N_14116,N_8597,N_6312);
and U14117 (N_14117,N_7625,N_8106);
nor U14118 (N_14118,N_6641,N_8640);
xnor U14119 (N_14119,N_8331,N_9146);
nor U14120 (N_14120,N_8126,N_8081);
nand U14121 (N_14121,N_7015,N_8493);
nand U14122 (N_14122,N_9726,N_5593);
nor U14123 (N_14123,N_5922,N_5796);
and U14124 (N_14124,N_7761,N_8677);
or U14125 (N_14125,N_6072,N_5021);
nand U14126 (N_14126,N_9330,N_9367);
or U14127 (N_14127,N_7444,N_9812);
nand U14128 (N_14128,N_8877,N_8110);
or U14129 (N_14129,N_7012,N_5539);
nand U14130 (N_14130,N_6235,N_7797);
nor U14131 (N_14131,N_9765,N_5158);
nor U14132 (N_14132,N_7845,N_9688);
nand U14133 (N_14133,N_8892,N_7282);
and U14134 (N_14134,N_5230,N_5802);
or U14135 (N_14135,N_7110,N_6788);
or U14136 (N_14136,N_8797,N_9181);
xor U14137 (N_14137,N_8054,N_9072);
or U14138 (N_14138,N_5351,N_6200);
nand U14139 (N_14139,N_5981,N_5765);
nand U14140 (N_14140,N_6798,N_6029);
and U14141 (N_14141,N_9959,N_7691);
xor U14142 (N_14142,N_8983,N_7201);
nand U14143 (N_14143,N_7685,N_9501);
nor U14144 (N_14144,N_6124,N_9190);
or U14145 (N_14145,N_5687,N_7178);
nor U14146 (N_14146,N_7759,N_5263);
and U14147 (N_14147,N_6208,N_6011);
and U14148 (N_14148,N_7095,N_5526);
nor U14149 (N_14149,N_9306,N_8159);
nor U14150 (N_14150,N_8977,N_6941);
and U14151 (N_14151,N_5127,N_6170);
or U14152 (N_14152,N_7937,N_8609);
nor U14153 (N_14153,N_5407,N_9877);
or U14154 (N_14154,N_6977,N_7847);
nor U14155 (N_14155,N_8213,N_6887);
or U14156 (N_14156,N_7913,N_7168);
or U14157 (N_14157,N_8740,N_7460);
nor U14158 (N_14158,N_7931,N_9574);
or U14159 (N_14159,N_7087,N_8565);
or U14160 (N_14160,N_9410,N_5306);
nor U14161 (N_14161,N_9160,N_6054);
nor U14162 (N_14162,N_7920,N_5041);
nor U14163 (N_14163,N_9639,N_6169);
and U14164 (N_14164,N_6617,N_6502);
or U14165 (N_14165,N_5449,N_6486);
nor U14166 (N_14166,N_6178,N_6763);
xnor U14167 (N_14167,N_7289,N_5011);
and U14168 (N_14168,N_8136,N_7382);
xor U14169 (N_14169,N_8465,N_8175);
nor U14170 (N_14170,N_8757,N_7249);
and U14171 (N_14171,N_8084,N_8355);
and U14172 (N_14172,N_6217,N_9267);
or U14173 (N_14173,N_9423,N_6842);
nor U14174 (N_14174,N_6224,N_5715);
and U14175 (N_14175,N_5954,N_7586);
and U14176 (N_14176,N_9685,N_8936);
and U14177 (N_14177,N_6769,N_7981);
nor U14178 (N_14178,N_5847,N_7783);
and U14179 (N_14179,N_6561,N_5586);
or U14180 (N_14180,N_8772,N_5027);
or U14181 (N_14181,N_7408,N_8091);
nand U14182 (N_14182,N_7606,N_7764);
nand U14183 (N_14183,N_7670,N_6825);
nor U14184 (N_14184,N_9360,N_9730);
or U14185 (N_14185,N_5486,N_9822);
nand U14186 (N_14186,N_7758,N_9551);
and U14187 (N_14187,N_6375,N_5451);
or U14188 (N_14188,N_6830,N_5889);
xnor U14189 (N_14189,N_8255,N_5418);
or U14190 (N_14190,N_8023,N_8545);
and U14191 (N_14191,N_9450,N_5499);
or U14192 (N_14192,N_6876,N_5023);
and U14193 (N_14193,N_8891,N_5528);
nor U14194 (N_14194,N_7288,N_8104);
nor U14195 (N_14195,N_9622,N_7915);
nand U14196 (N_14196,N_6069,N_8377);
nand U14197 (N_14197,N_5430,N_6508);
nor U14198 (N_14198,N_9213,N_7884);
nor U14199 (N_14199,N_8464,N_8986);
nor U14200 (N_14200,N_8496,N_7095);
and U14201 (N_14201,N_9571,N_8344);
and U14202 (N_14202,N_7375,N_6566);
or U14203 (N_14203,N_6872,N_5977);
nor U14204 (N_14204,N_9087,N_6407);
and U14205 (N_14205,N_5912,N_5620);
nand U14206 (N_14206,N_8325,N_9939);
nand U14207 (N_14207,N_7454,N_5748);
nand U14208 (N_14208,N_7924,N_6640);
nor U14209 (N_14209,N_9206,N_7014);
or U14210 (N_14210,N_8314,N_9175);
nand U14211 (N_14211,N_5483,N_9255);
and U14212 (N_14212,N_6645,N_5607);
nand U14213 (N_14213,N_5959,N_6856);
or U14214 (N_14214,N_9529,N_5460);
xnor U14215 (N_14215,N_7323,N_6235);
nand U14216 (N_14216,N_5894,N_8386);
or U14217 (N_14217,N_5067,N_8678);
and U14218 (N_14218,N_8172,N_5463);
nor U14219 (N_14219,N_5009,N_8173);
nor U14220 (N_14220,N_7456,N_6781);
nand U14221 (N_14221,N_9547,N_8351);
or U14222 (N_14222,N_9331,N_7658);
or U14223 (N_14223,N_9652,N_9286);
xnor U14224 (N_14224,N_9671,N_9378);
nor U14225 (N_14225,N_7195,N_7827);
nor U14226 (N_14226,N_9474,N_7545);
xor U14227 (N_14227,N_8492,N_5450);
xnor U14228 (N_14228,N_9494,N_8856);
nor U14229 (N_14229,N_6637,N_5976);
and U14230 (N_14230,N_9226,N_6485);
and U14231 (N_14231,N_7000,N_5415);
nor U14232 (N_14232,N_9470,N_5818);
or U14233 (N_14233,N_7840,N_7010);
xnor U14234 (N_14234,N_9630,N_7998);
nand U14235 (N_14235,N_7177,N_5684);
nand U14236 (N_14236,N_6350,N_7704);
or U14237 (N_14237,N_6728,N_9748);
or U14238 (N_14238,N_5443,N_5700);
xor U14239 (N_14239,N_7266,N_6507);
xnor U14240 (N_14240,N_5702,N_8432);
nor U14241 (N_14241,N_8789,N_9195);
nor U14242 (N_14242,N_6080,N_6660);
or U14243 (N_14243,N_6023,N_7639);
or U14244 (N_14244,N_5872,N_8242);
nand U14245 (N_14245,N_9824,N_5196);
and U14246 (N_14246,N_8327,N_8971);
and U14247 (N_14247,N_9955,N_5895);
nand U14248 (N_14248,N_5558,N_6160);
or U14249 (N_14249,N_6986,N_6794);
nand U14250 (N_14250,N_7898,N_7747);
or U14251 (N_14251,N_6723,N_8610);
xor U14252 (N_14252,N_8266,N_9195);
xnor U14253 (N_14253,N_9341,N_8702);
nor U14254 (N_14254,N_9681,N_7374);
nor U14255 (N_14255,N_5663,N_9490);
and U14256 (N_14256,N_9183,N_7865);
nand U14257 (N_14257,N_8548,N_9587);
xnor U14258 (N_14258,N_9383,N_7535);
or U14259 (N_14259,N_8686,N_6322);
nor U14260 (N_14260,N_8411,N_6753);
or U14261 (N_14261,N_6004,N_9250);
nand U14262 (N_14262,N_5644,N_8856);
or U14263 (N_14263,N_6533,N_9470);
nor U14264 (N_14264,N_7104,N_7347);
and U14265 (N_14265,N_5204,N_7975);
xnor U14266 (N_14266,N_7098,N_8464);
nand U14267 (N_14267,N_6029,N_7967);
xnor U14268 (N_14268,N_8245,N_9929);
and U14269 (N_14269,N_5092,N_5770);
nand U14270 (N_14270,N_6606,N_7335);
nand U14271 (N_14271,N_5633,N_5406);
nor U14272 (N_14272,N_8459,N_7645);
and U14273 (N_14273,N_7420,N_6312);
and U14274 (N_14274,N_7513,N_9273);
or U14275 (N_14275,N_5061,N_7504);
nor U14276 (N_14276,N_7337,N_9014);
xnor U14277 (N_14277,N_9411,N_7142);
nor U14278 (N_14278,N_9961,N_5787);
or U14279 (N_14279,N_9425,N_6539);
or U14280 (N_14280,N_8401,N_7450);
and U14281 (N_14281,N_9734,N_9338);
and U14282 (N_14282,N_7176,N_6126);
xnor U14283 (N_14283,N_9333,N_9962);
nand U14284 (N_14284,N_5150,N_7530);
nor U14285 (N_14285,N_7343,N_8297);
and U14286 (N_14286,N_6079,N_5706);
nor U14287 (N_14287,N_9000,N_5488);
nand U14288 (N_14288,N_5368,N_5064);
nor U14289 (N_14289,N_7490,N_9483);
nand U14290 (N_14290,N_7445,N_6548);
nor U14291 (N_14291,N_5389,N_7554);
nor U14292 (N_14292,N_6406,N_7014);
and U14293 (N_14293,N_6887,N_9063);
and U14294 (N_14294,N_7882,N_6527);
nor U14295 (N_14295,N_8545,N_8196);
or U14296 (N_14296,N_5457,N_5645);
nor U14297 (N_14297,N_6141,N_9812);
nor U14298 (N_14298,N_7760,N_9278);
nor U14299 (N_14299,N_7170,N_9930);
nor U14300 (N_14300,N_9682,N_6578);
nor U14301 (N_14301,N_5147,N_7566);
nor U14302 (N_14302,N_7644,N_8960);
xnor U14303 (N_14303,N_9841,N_9602);
and U14304 (N_14304,N_6662,N_9798);
nor U14305 (N_14305,N_7174,N_9133);
or U14306 (N_14306,N_9518,N_8857);
and U14307 (N_14307,N_6010,N_8124);
nor U14308 (N_14308,N_6491,N_9411);
nor U14309 (N_14309,N_6484,N_8700);
nand U14310 (N_14310,N_7922,N_6544);
or U14311 (N_14311,N_9689,N_8260);
xor U14312 (N_14312,N_9596,N_6361);
or U14313 (N_14313,N_8200,N_5293);
and U14314 (N_14314,N_6387,N_7030);
nand U14315 (N_14315,N_8104,N_9711);
or U14316 (N_14316,N_7237,N_7650);
xnor U14317 (N_14317,N_8593,N_5562);
xor U14318 (N_14318,N_9732,N_5254);
nand U14319 (N_14319,N_7948,N_6356);
nor U14320 (N_14320,N_6389,N_9934);
nand U14321 (N_14321,N_7540,N_7357);
or U14322 (N_14322,N_9298,N_5429);
and U14323 (N_14323,N_6997,N_7887);
nand U14324 (N_14324,N_8809,N_8422);
and U14325 (N_14325,N_9571,N_6938);
nand U14326 (N_14326,N_9459,N_5212);
and U14327 (N_14327,N_9162,N_7422);
nand U14328 (N_14328,N_9879,N_6836);
nand U14329 (N_14329,N_5772,N_8453);
nand U14330 (N_14330,N_6814,N_9698);
nor U14331 (N_14331,N_6669,N_6280);
nor U14332 (N_14332,N_5164,N_5212);
nand U14333 (N_14333,N_9174,N_7642);
or U14334 (N_14334,N_7970,N_7575);
or U14335 (N_14335,N_7733,N_8516);
or U14336 (N_14336,N_7523,N_7110);
or U14337 (N_14337,N_7131,N_5842);
and U14338 (N_14338,N_5848,N_6230);
nand U14339 (N_14339,N_8454,N_9166);
xnor U14340 (N_14340,N_6546,N_6967);
or U14341 (N_14341,N_9782,N_5759);
or U14342 (N_14342,N_8657,N_9340);
nand U14343 (N_14343,N_5745,N_8934);
nor U14344 (N_14344,N_8307,N_7418);
and U14345 (N_14345,N_7874,N_8253);
nand U14346 (N_14346,N_8933,N_6014);
or U14347 (N_14347,N_9870,N_8850);
or U14348 (N_14348,N_7456,N_6469);
nor U14349 (N_14349,N_9127,N_7068);
nor U14350 (N_14350,N_7289,N_9133);
nor U14351 (N_14351,N_9573,N_6073);
nor U14352 (N_14352,N_5919,N_9690);
or U14353 (N_14353,N_5498,N_6540);
nand U14354 (N_14354,N_5624,N_9424);
or U14355 (N_14355,N_5390,N_8412);
nand U14356 (N_14356,N_8443,N_7904);
and U14357 (N_14357,N_7686,N_6799);
nor U14358 (N_14358,N_9069,N_5037);
nor U14359 (N_14359,N_6170,N_7401);
nand U14360 (N_14360,N_8280,N_5655);
nand U14361 (N_14361,N_5920,N_7747);
nand U14362 (N_14362,N_9856,N_8194);
or U14363 (N_14363,N_5665,N_9940);
xor U14364 (N_14364,N_6415,N_5067);
nor U14365 (N_14365,N_8970,N_6914);
and U14366 (N_14366,N_7815,N_9771);
or U14367 (N_14367,N_5555,N_7285);
nand U14368 (N_14368,N_9963,N_8377);
or U14369 (N_14369,N_8896,N_7223);
nor U14370 (N_14370,N_7571,N_9214);
and U14371 (N_14371,N_7057,N_9306);
nor U14372 (N_14372,N_6029,N_8358);
nand U14373 (N_14373,N_5513,N_5246);
and U14374 (N_14374,N_6539,N_7533);
xor U14375 (N_14375,N_5197,N_9912);
nor U14376 (N_14376,N_6938,N_5834);
or U14377 (N_14377,N_8929,N_8544);
or U14378 (N_14378,N_7207,N_9149);
nor U14379 (N_14379,N_8050,N_9974);
nor U14380 (N_14380,N_6194,N_8296);
xnor U14381 (N_14381,N_6120,N_8999);
nand U14382 (N_14382,N_9996,N_6552);
and U14383 (N_14383,N_7666,N_8668);
and U14384 (N_14384,N_5995,N_8102);
and U14385 (N_14385,N_8786,N_6436);
nor U14386 (N_14386,N_9479,N_7019);
or U14387 (N_14387,N_8541,N_9213);
and U14388 (N_14388,N_8655,N_5308);
and U14389 (N_14389,N_6536,N_6185);
xnor U14390 (N_14390,N_8188,N_6735);
nand U14391 (N_14391,N_8925,N_9217);
xor U14392 (N_14392,N_5985,N_8427);
or U14393 (N_14393,N_9244,N_9456);
and U14394 (N_14394,N_6161,N_5737);
nor U14395 (N_14395,N_9415,N_5538);
and U14396 (N_14396,N_8612,N_5222);
and U14397 (N_14397,N_5359,N_6503);
or U14398 (N_14398,N_6164,N_9238);
nor U14399 (N_14399,N_6712,N_7824);
nor U14400 (N_14400,N_7890,N_9250);
or U14401 (N_14401,N_7473,N_6069);
nand U14402 (N_14402,N_5014,N_5766);
nor U14403 (N_14403,N_7880,N_8158);
xnor U14404 (N_14404,N_6001,N_5165);
or U14405 (N_14405,N_9645,N_7057);
nand U14406 (N_14406,N_9596,N_9493);
nor U14407 (N_14407,N_9993,N_7931);
and U14408 (N_14408,N_6908,N_5305);
nor U14409 (N_14409,N_9733,N_9932);
nand U14410 (N_14410,N_5135,N_8028);
and U14411 (N_14411,N_6369,N_5913);
nor U14412 (N_14412,N_5377,N_9166);
nand U14413 (N_14413,N_9284,N_6590);
nand U14414 (N_14414,N_7294,N_5974);
nor U14415 (N_14415,N_7576,N_9781);
nand U14416 (N_14416,N_6421,N_9469);
nand U14417 (N_14417,N_8985,N_5564);
and U14418 (N_14418,N_5243,N_9460);
or U14419 (N_14419,N_8371,N_8102);
nor U14420 (N_14420,N_9880,N_6227);
nand U14421 (N_14421,N_5041,N_7828);
nor U14422 (N_14422,N_6781,N_8445);
nand U14423 (N_14423,N_6390,N_8413);
nand U14424 (N_14424,N_7696,N_7147);
xor U14425 (N_14425,N_6988,N_8578);
nand U14426 (N_14426,N_5236,N_9827);
or U14427 (N_14427,N_9203,N_9765);
nor U14428 (N_14428,N_8636,N_8998);
and U14429 (N_14429,N_7645,N_7433);
nand U14430 (N_14430,N_9567,N_7942);
or U14431 (N_14431,N_6712,N_5657);
and U14432 (N_14432,N_6947,N_6859);
nor U14433 (N_14433,N_8993,N_8726);
nand U14434 (N_14434,N_9873,N_5607);
or U14435 (N_14435,N_5706,N_7155);
and U14436 (N_14436,N_6835,N_9745);
or U14437 (N_14437,N_5215,N_8469);
nor U14438 (N_14438,N_9506,N_7751);
xor U14439 (N_14439,N_8085,N_6349);
nor U14440 (N_14440,N_5438,N_8113);
or U14441 (N_14441,N_5156,N_9782);
nor U14442 (N_14442,N_7125,N_7867);
nor U14443 (N_14443,N_6105,N_8359);
nor U14444 (N_14444,N_5724,N_5393);
and U14445 (N_14445,N_6719,N_5448);
and U14446 (N_14446,N_6584,N_5091);
and U14447 (N_14447,N_5941,N_6311);
nor U14448 (N_14448,N_6089,N_8094);
nor U14449 (N_14449,N_6541,N_5478);
and U14450 (N_14450,N_6576,N_9588);
nand U14451 (N_14451,N_5416,N_5765);
nand U14452 (N_14452,N_8920,N_6434);
nand U14453 (N_14453,N_6972,N_9930);
nor U14454 (N_14454,N_8617,N_8080);
nor U14455 (N_14455,N_8498,N_5883);
or U14456 (N_14456,N_7670,N_8538);
nand U14457 (N_14457,N_9582,N_5967);
xnor U14458 (N_14458,N_6844,N_7023);
xnor U14459 (N_14459,N_6397,N_8905);
nor U14460 (N_14460,N_8181,N_6905);
nand U14461 (N_14461,N_5918,N_9801);
nand U14462 (N_14462,N_6397,N_8303);
nor U14463 (N_14463,N_9790,N_8391);
nor U14464 (N_14464,N_5042,N_8871);
or U14465 (N_14465,N_8937,N_6844);
nor U14466 (N_14466,N_9116,N_7167);
and U14467 (N_14467,N_8349,N_9216);
nor U14468 (N_14468,N_9331,N_7462);
or U14469 (N_14469,N_7648,N_7654);
nand U14470 (N_14470,N_6311,N_6885);
nor U14471 (N_14471,N_6987,N_6626);
nor U14472 (N_14472,N_8607,N_5029);
nand U14473 (N_14473,N_6321,N_5561);
or U14474 (N_14474,N_6741,N_8265);
or U14475 (N_14475,N_6348,N_8776);
nor U14476 (N_14476,N_9840,N_5651);
nor U14477 (N_14477,N_8690,N_9255);
and U14478 (N_14478,N_6206,N_7045);
and U14479 (N_14479,N_5443,N_6802);
nor U14480 (N_14480,N_6030,N_9392);
and U14481 (N_14481,N_8490,N_6880);
xor U14482 (N_14482,N_5211,N_5592);
nand U14483 (N_14483,N_5269,N_7626);
nor U14484 (N_14484,N_7600,N_7563);
nor U14485 (N_14485,N_7012,N_5735);
or U14486 (N_14486,N_6039,N_6527);
nor U14487 (N_14487,N_5568,N_7229);
or U14488 (N_14488,N_8128,N_5798);
or U14489 (N_14489,N_8248,N_8153);
xnor U14490 (N_14490,N_7990,N_5842);
and U14491 (N_14491,N_9462,N_5160);
nor U14492 (N_14492,N_7672,N_9979);
xnor U14493 (N_14493,N_6388,N_6585);
xnor U14494 (N_14494,N_5274,N_7516);
or U14495 (N_14495,N_7466,N_9028);
nor U14496 (N_14496,N_8601,N_6054);
nand U14497 (N_14497,N_8187,N_8621);
nor U14498 (N_14498,N_8843,N_8119);
nor U14499 (N_14499,N_5152,N_6396);
nor U14500 (N_14500,N_8892,N_7232);
nand U14501 (N_14501,N_8830,N_8900);
or U14502 (N_14502,N_5577,N_8084);
or U14503 (N_14503,N_6252,N_6006);
nor U14504 (N_14504,N_6399,N_6763);
nor U14505 (N_14505,N_8809,N_8358);
nand U14506 (N_14506,N_9285,N_8300);
and U14507 (N_14507,N_8636,N_5530);
or U14508 (N_14508,N_9750,N_9036);
or U14509 (N_14509,N_8697,N_7816);
and U14510 (N_14510,N_7742,N_8740);
nor U14511 (N_14511,N_6479,N_9346);
nor U14512 (N_14512,N_8087,N_6722);
or U14513 (N_14513,N_6628,N_6862);
nor U14514 (N_14514,N_9995,N_5987);
nor U14515 (N_14515,N_9856,N_7402);
nor U14516 (N_14516,N_9838,N_8729);
xnor U14517 (N_14517,N_9323,N_7715);
nand U14518 (N_14518,N_9864,N_9769);
xnor U14519 (N_14519,N_8507,N_6137);
nand U14520 (N_14520,N_8430,N_9704);
nand U14521 (N_14521,N_8545,N_7954);
nand U14522 (N_14522,N_8261,N_6490);
nand U14523 (N_14523,N_5230,N_7923);
or U14524 (N_14524,N_6362,N_7460);
nand U14525 (N_14525,N_6974,N_6540);
or U14526 (N_14526,N_7708,N_7193);
and U14527 (N_14527,N_6650,N_6854);
nand U14528 (N_14528,N_5159,N_5179);
nand U14529 (N_14529,N_5185,N_6528);
nand U14530 (N_14530,N_9849,N_5982);
xnor U14531 (N_14531,N_6495,N_7727);
xnor U14532 (N_14532,N_7895,N_6434);
and U14533 (N_14533,N_5170,N_7611);
nor U14534 (N_14534,N_7934,N_5464);
or U14535 (N_14535,N_9530,N_7788);
and U14536 (N_14536,N_8517,N_8574);
nand U14537 (N_14537,N_8867,N_6027);
nand U14538 (N_14538,N_5609,N_9831);
nor U14539 (N_14539,N_9162,N_9568);
or U14540 (N_14540,N_6412,N_7107);
or U14541 (N_14541,N_9744,N_5481);
nor U14542 (N_14542,N_8990,N_5299);
nor U14543 (N_14543,N_8392,N_6552);
nand U14544 (N_14544,N_5942,N_9424);
and U14545 (N_14545,N_5361,N_7920);
nand U14546 (N_14546,N_9945,N_7615);
and U14547 (N_14547,N_5757,N_7523);
or U14548 (N_14548,N_9204,N_8235);
and U14549 (N_14549,N_5867,N_8574);
xnor U14550 (N_14550,N_6272,N_9820);
and U14551 (N_14551,N_6575,N_6915);
nand U14552 (N_14552,N_5051,N_6454);
nand U14553 (N_14553,N_5148,N_6592);
nor U14554 (N_14554,N_7565,N_5967);
nor U14555 (N_14555,N_6066,N_5413);
xor U14556 (N_14556,N_6589,N_6708);
or U14557 (N_14557,N_7722,N_7413);
or U14558 (N_14558,N_9582,N_7261);
nor U14559 (N_14559,N_7320,N_6472);
nor U14560 (N_14560,N_6035,N_9007);
nand U14561 (N_14561,N_7014,N_5824);
nand U14562 (N_14562,N_7998,N_6301);
nand U14563 (N_14563,N_7273,N_6500);
or U14564 (N_14564,N_9831,N_8467);
or U14565 (N_14565,N_5065,N_8500);
and U14566 (N_14566,N_6930,N_9722);
nor U14567 (N_14567,N_9313,N_5883);
or U14568 (N_14568,N_9075,N_6846);
or U14569 (N_14569,N_5469,N_9522);
and U14570 (N_14570,N_7507,N_5902);
and U14571 (N_14571,N_6077,N_7692);
nor U14572 (N_14572,N_5330,N_6555);
and U14573 (N_14573,N_7762,N_8628);
and U14574 (N_14574,N_5616,N_7710);
xnor U14575 (N_14575,N_6137,N_8322);
nor U14576 (N_14576,N_9591,N_7942);
nand U14577 (N_14577,N_9275,N_9921);
or U14578 (N_14578,N_9921,N_7138);
or U14579 (N_14579,N_9638,N_6164);
or U14580 (N_14580,N_7882,N_6063);
or U14581 (N_14581,N_7356,N_8282);
nand U14582 (N_14582,N_5724,N_8134);
nor U14583 (N_14583,N_9233,N_9248);
or U14584 (N_14584,N_7251,N_9140);
or U14585 (N_14585,N_9936,N_5167);
nor U14586 (N_14586,N_6045,N_6600);
nor U14587 (N_14587,N_5761,N_5642);
nand U14588 (N_14588,N_5665,N_7597);
xor U14589 (N_14589,N_7647,N_7207);
nand U14590 (N_14590,N_5347,N_5125);
and U14591 (N_14591,N_6569,N_5733);
and U14592 (N_14592,N_9069,N_8268);
xnor U14593 (N_14593,N_6010,N_9621);
and U14594 (N_14594,N_9038,N_9571);
and U14595 (N_14595,N_7125,N_8287);
nand U14596 (N_14596,N_7654,N_9954);
or U14597 (N_14597,N_7111,N_9563);
nor U14598 (N_14598,N_6880,N_7118);
and U14599 (N_14599,N_6941,N_9292);
nor U14600 (N_14600,N_5726,N_8447);
and U14601 (N_14601,N_7833,N_7033);
nand U14602 (N_14602,N_5019,N_7814);
and U14603 (N_14603,N_6831,N_7680);
xnor U14604 (N_14604,N_6818,N_7145);
and U14605 (N_14605,N_8110,N_8967);
nor U14606 (N_14606,N_9698,N_9257);
nand U14607 (N_14607,N_7787,N_7810);
or U14608 (N_14608,N_6875,N_6158);
xnor U14609 (N_14609,N_9971,N_9900);
nor U14610 (N_14610,N_8983,N_7394);
nand U14611 (N_14611,N_6102,N_7300);
and U14612 (N_14612,N_9062,N_9784);
or U14613 (N_14613,N_7001,N_5594);
and U14614 (N_14614,N_7480,N_5878);
xnor U14615 (N_14615,N_7098,N_5505);
nor U14616 (N_14616,N_7289,N_8265);
or U14617 (N_14617,N_5108,N_6780);
and U14618 (N_14618,N_6484,N_5143);
nor U14619 (N_14619,N_7183,N_8573);
nor U14620 (N_14620,N_7521,N_6849);
or U14621 (N_14621,N_5832,N_6818);
and U14622 (N_14622,N_6053,N_5944);
nor U14623 (N_14623,N_7940,N_9977);
nand U14624 (N_14624,N_6443,N_6591);
or U14625 (N_14625,N_6863,N_6549);
nor U14626 (N_14626,N_8524,N_5073);
xnor U14627 (N_14627,N_6553,N_9654);
nor U14628 (N_14628,N_9421,N_6488);
and U14629 (N_14629,N_5478,N_8059);
nor U14630 (N_14630,N_7973,N_6545);
or U14631 (N_14631,N_6649,N_8960);
nand U14632 (N_14632,N_9761,N_8444);
or U14633 (N_14633,N_6529,N_6691);
nand U14634 (N_14634,N_7555,N_9758);
nand U14635 (N_14635,N_9836,N_8225);
or U14636 (N_14636,N_7307,N_5609);
or U14637 (N_14637,N_7936,N_5261);
nor U14638 (N_14638,N_6513,N_5928);
or U14639 (N_14639,N_7204,N_5461);
or U14640 (N_14640,N_7640,N_6653);
xnor U14641 (N_14641,N_6293,N_7060);
nand U14642 (N_14642,N_6241,N_7869);
xnor U14643 (N_14643,N_6936,N_8298);
or U14644 (N_14644,N_6915,N_9332);
or U14645 (N_14645,N_6479,N_9644);
or U14646 (N_14646,N_8208,N_6930);
xor U14647 (N_14647,N_8585,N_9628);
or U14648 (N_14648,N_9339,N_6137);
or U14649 (N_14649,N_7620,N_5330);
or U14650 (N_14650,N_8571,N_7258);
nand U14651 (N_14651,N_8279,N_9874);
nor U14652 (N_14652,N_8177,N_9461);
nor U14653 (N_14653,N_8852,N_9403);
xnor U14654 (N_14654,N_9709,N_9058);
nand U14655 (N_14655,N_5938,N_6111);
and U14656 (N_14656,N_7417,N_5291);
or U14657 (N_14657,N_7227,N_5777);
nor U14658 (N_14658,N_7919,N_7443);
and U14659 (N_14659,N_9147,N_9261);
or U14660 (N_14660,N_8746,N_7610);
nand U14661 (N_14661,N_5929,N_9127);
or U14662 (N_14662,N_5097,N_7502);
nand U14663 (N_14663,N_9704,N_5527);
nand U14664 (N_14664,N_9457,N_8119);
xor U14665 (N_14665,N_5135,N_7559);
or U14666 (N_14666,N_6681,N_6462);
nand U14667 (N_14667,N_8488,N_8777);
nor U14668 (N_14668,N_8419,N_7037);
and U14669 (N_14669,N_9904,N_5260);
nand U14670 (N_14670,N_6863,N_8976);
nor U14671 (N_14671,N_7831,N_9088);
or U14672 (N_14672,N_7471,N_9747);
or U14673 (N_14673,N_5944,N_9217);
nor U14674 (N_14674,N_6278,N_6320);
or U14675 (N_14675,N_8624,N_7971);
nand U14676 (N_14676,N_8126,N_6636);
xnor U14677 (N_14677,N_7213,N_5118);
and U14678 (N_14678,N_9420,N_5419);
and U14679 (N_14679,N_8744,N_7199);
nor U14680 (N_14680,N_9081,N_8806);
nand U14681 (N_14681,N_6048,N_9202);
or U14682 (N_14682,N_5326,N_6733);
xor U14683 (N_14683,N_8706,N_6862);
nand U14684 (N_14684,N_6462,N_9682);
and U14685 (N_14685,N_6575,N_6571);
nand U14686 (N_14686,N_9803,N_8093);
or U14687 (N_14687,N_6540,N_6457);
nor U14688 (N_14688,N_8051,N_7574);
and U14689 (N_14689,N_9284,N_6284);
nor U14690 (N_14690,N_9586,N_7001);
or U14691 (N_14691,N_8263,N_9826);
nor U14692 (N_14692,N_8327,N_8225);
or U14693 (N_14693,N_5524,N_8477);
or U14694 (N_14694,N_9057,N_8871);
and U14695 (N_14695,N_7002,N_5222);
xor U14696 (N_14696,N_9729,N_7120);
or U14697 (N_14697,N_8994,N_6603);
nor U14698 (N_14698,N_9303,N_5552);
nand U14699 (N_14699,N_9388,N_5798);
and U14700 (N_14700,N_7322,N_6261);
xnor U14701 (N_14701,N_5697,N_5811);
nor U14702 (N_14702,N_5675,N_5754);
nor U14703 (N_14703,N_9855,N_9774);
nor U14704 (N_14704,N_6636,N_9843);
nand U14705 (N_14705,N_8753,N_8629);
xor U14706 (N_14706,N_9101,N_6192);
nor U14707 (N_14707,N_7312,N_9194);
or U14708 (N_14708,N_6409,N_6350);
nor U14709 (N_14709,N_6323,N_8936);
or U14710 (N_14710,N_6659,N_8848);
or U14711 (N_14711,N_7706,N_8543);
and U14712 (N_14712,N_7377,N_7264);
or U14713 (N_14713,N_6725,N_7690);
and U14714 (N_14714,N_7283,N_7785);
nand U14715 (N_14715,N_8551,N_5318);
nor U14716 (N_14716,N_9532,N_6016);
nor U14717 (N_14717,N_6468,N_6063);
nor U14718 (N_14718,N_9658,N_9101);
xor U14719 (N_14719,N_7757,N_5932);
nand U14720 (N_14720,N_9884,N_5589);
nand U14721 (N_14721,N_5880,N_6481);
or U14722 (N_14722,N_5432,N_5573);
nor U14723 (N_14723,N_7377,N_6662);
nand U14724 (N_14724,N_6107,N_9197);
or U14725 (N_14725,N_6239,N_7258);
and U14726 (N_14726,N_7997,N_5060);
nor U14727 (N_14727,N_9537,N_7591);
or U14728 (N_14728,N_8352,N_8722);
nand U14729 (N_14729,N_5521,N_5978);
xnor U14730 (N_14730,N_7433,N_6075);
nand U14731 (N_14731,N_7272,N_8547);
nand U14732 (N_14732,N_8346,N_5034);
or U14733 (N_14733,N_5295,N_5077);
nand U14734 (N_14734,N_9113,N_8491);
or U14735 (N_14735,N_5211,N_6480);
and U14736 (N_14736,N_9510,N_7717);
nand U14737 (N_14737,N_8758,N_6245);
or U14738 (N_14738,N_9228,N_7237);
nand U14739 (N_14739,N_6037,N_5523);
and U14740 (N_14740,N_6558,N_6332);
nand U14741 (N_14741,N_9411,N_5606);
nor U14742 (N_14742,N_6987,N_6177);
nor U14743 (N_14743,N_5640,N_9585);
nor U14744 (N_14744,N_5451,N_7204);
xor U14745 (N_14745,N_5769,N_6049);
nand U14746 (N_14746,N_7085,N_9257);
and U14747 (N_14747,N_8399,N_5252);
nor U14748 (N_14748,N_6390,N_5678);
nor U14749 (N_14749,N_6681,N_9464);
nor U14750 (N_14750,N_6357,N_9759);
xor U14751 (N_14751,N_9792,N_9032);
or U14752 (N_14752,N_6524,N_9021);
nor U14753 (N_14753,N_8394,N_9688);
nand U14754 (N_14754,N_6055,N_8351);
nor U14755 (N_14755,N_6932,N_5157);
or U14756 (N_14756,N_8597,N_9200);
xor U14757 (N_14757,N_7131,N_5296);
and U14758 (N_14758,N_9232,N_9827);
nor U14759 (N_14759,N_9437,N_5778);
or U14760 (N_14760,N_9986,N_5575);
nand U14761 (N_14761,N_7706,N_7031);
or U14762 (N_14762,N_8350,N_9972);
nand U14763 (N_14763,N_6855,N_8476);
or U14764 (N_14764,N_6685,N_5493);
nor U14765 (N_14765,N_6729,N_9513);
nand U14766 (N_14766,N_6687,N_7868);
xnor U14767 (N_14767,N_9012,N_7371);
nand U14768 (N_14768,N_5076,N_7503);
nand U14769 (N_14769,N_7121,N_9096);
nand U14770 (N_14770,N_5203,N_6175);
nand U14771 (N_14771,N_5997,N_9543);
or U14772 (N_14772,N_6468,N_8011);
and U14773 (N_14773,N_8124,N_7495);
or U14774 (N_14774,N_5588,N_9120);
and U14775 (N_14775,N_5427,N_7669);
nand U14776 (N_14776,N_9928,N_9538);
nand U14777 (N_14777,N_5419,N_8271);
or U14778 (N_14778,N_7365,N_7573);
nor U14779 (N_14779,N_6165,N_6560);
and U14780 (N_14780,N_8242,N_9011);
xor U14781 (N_14781,N_8666,N_6232);
and U14782 (N_14782,N_5592,N_5964);
and U14783 (N_14783,N_9692,N_6559);
nor U14784 (N_14784,N_7717,N_6361);
nor U14785 (N_14785,N_9821,N_7764);
nand U14786 (N_14786,N_6267,N_9985);
or U14787 (N_14787,N_7903,N_5616);
or U14788 (N_14788,N_5802,N_6028);
xnor U14789 (N_14789,N_9294,N_5717);
or U14790 (N_14790,N_5491,N_7626);
and U14791 (N_14791,N_6841,N_8122);
or U14792 (N_14792,N_9134,N_8289);
and U14793 (N_14793,N_6528,N_8638);
or U14794 (N_14794,N_9869,N_9398);
and U14795 (N_14795,N_9913,N_6297);
nor U14796 (N_14796,N_6038,N_5687);
nand U14797 (N_14797,N_5079,N_5800);
nand U14798 (N_14798,N_9913,N_5034);
and U14799 (N_14799,N_9272,N_5721);
or U14800 (N_14800,N_6862,N_7669);
nor U14801 (N_14801,N_9242,N_7637);
nand U14802 (N_14802,N_5094,N_8843);
or U14803 (N_14803,N_5193,N_8942);
nor U14804 (N_14804,N_7251,N_7324);
and U14805 (N_14805,N_9806,N_7924);
nor U14806 (N_14806,N_9183,N_7496);
nand U14807 (N_14807,N_8868,N_7774);
xor U14808 (N_14808,N_6071,N_9823);
or U14809 (N_14809,N_9956,N_9672);
nor U14810 (N_14810,N_7035,N_7218);
and U14811 (N_14811,N_8480,N_8664);
and U14812 (N_14812,N_8877,N_9926);
and U14813 (N_14813,N_8136,N_8031);
nand U14814 (N_14814,N_6557,N_9661);
nor U14815 (N_14815,N_7817,N_5923);
nor U14816 (N_14816,N_5499,N_5662);
and U14817 (N_14817,N_6885,N_8262);
nor U14818 (N_14818,N_7757,N_7658);
or U14819 (N_14819,N_8666,N_6450);
nand U14820 (N_14820,N_8121,N_8331);
xor U14821 (N_14821,N_6183,N_6475);
nor U14822 (N_14822,N_5792,N_7797);
nor U14823 (N_14823,N_6938,N_8482);
nor U14824 (N_14824,N_8639,N_8396);
and U14825 (N_14825,N_6381,N_5254);
nand U14826 (N_14826,N_7071,N_5881);
nor U14827 (N_14827,N_6814,N_8602);
nand U14828 (N_14828,N_8354,N_9270);
nor U14829 (N_14829,N_5242,N_5945);
nor U14830 (N_14830,N_8914,N_8683);
and U14831 (N_14831,N_9138,N_8535);
nor U14832 (N_14832,N_7210,N_9303);
or U14833 (N_14833,N_6036,N_8410);
nand U14834 (N_14834,N_9830,N_6250);
nand U14835 (N_14835,N_8102,N_6919);
nand U14836 (N_14836,N_6574,N_9551);
xnor U14837 (N_14837,N_7990,N_8772);
nand U14838 (N_14838,N_5876,N_7121);
and U14839 (N_14839,N_9880,N_9795);
xor U14840 (N_14840,N_5033,N_9655);
nor U14841 (N_14841,N_6878,N_6880);
nand U14842 (N_14842,N_7275,N_9997);
or U14843 (N_14843,N_6496,N_7330);
or U14844 (N_14844,N_7298,N_8616);
or U14845 (N_14845,N_9160,N_7605);
xor U14846 (N_14846,N_7740,N_7699);
and U14847 (N_14847,N_6337,N_5157);
nor U14848 (N_14848,N_8112,N_9317);
or U14849 (N_14849,N_9005,N_9909);
nand U14850 (N_14850,N_6413,N_7442);
xor U14851 (N_14851,N_7762,N_5767);
nand U14852 (N_14852,N_5243,N_5844);
nand U14853 (N_14853,N_8269,N_6867);
and U14854 (N_14854,N_7535,N_9308);
xor U14855 (N_14855,N_7520,N_9007);
or U14856 (N_14856,N_8354,N_6205);
nor U14857 (N_14857,N_6726,N_5834);
and U14858 (N_14858,N_7951,N_8487);
xor U14859 (N_14859,N_8458,N_8049);
and U14860 (N_14860,N_8668,N_8320);
and U14861 (N_14861,N_8592,N_5881);
xnor U14862 (N_14862,N_5931,N_7717);
nor U14863 (N_14863,N_6188,N_8719);
xnor U14864 (N_14864,N_5569,N_5113);
or U14865 (N_14865,N_7868,N_8746);
and U14866 (N_14866,N_7942,N_5110);
nand U14867 (N_14867,N_9426,N_5231);
nand U14868 (N_14868,N_8484,N_6769);
nor U14869 (N_14869,N_8970,N_9088);
or U14870 (N_14870,N_7543,N_7691);
nor U14871 (N_14871,N_5583,N_6027);
nand U14872 (N_14872,N_8051,N_7347);
nor U14873 (N_14873,N_6205,N_8492);
nor U14874 (N_14874,N_5105,N_7599);
or U14875 (N_14875,N_7353,N_5192);
and U14876 (N_14876,N_9614,N_7013);
xor U14877 (N_14877,N_7186,N_9772);
or U14878 (N_14878,N_9976,N_9639);
and U14879 (N_14879,N_9382,N_7457);
nor U14880 (N_14880,N_9937,N_9310);
nand U14881 (N_14881,N_5162,N_5710);
or U14882 (N_14882,N_7974,N_8856);
nor U14883 (N_14883,N_5825,N_6024);
and U14884 (N_14884,N_6306,N_6605);
nand U14885 (N_14885,N_7860,N_7011);
and U14886 (N_14886,N_7071,N_7032);
nand U14887 (N_14887,N_6985,N_5516);
nand U14888 (N_14888,N_5748,N_7347);
nand U14889 (N_14889,N_6426,N_9501);
xor U14890 (N_14890,N_8589,N_8666);
nand U14891 (N_14891,N_7670,N_9195);
nor U14892 (N_14892,N_8413,N_7926);
nand U14893 (N_14893,N_8294,N_9603);
xnor U14894 (N_14894,N_5866,N_9250);
xor U14895 (N_14895,N_5074,N_7346);
nor U14896 (N_14896,N_7144,N_7146);
or U14897 (N_14897,N_8094,N_9442);
and U14898 (N_14898,N_9692,N_8440);
xnor U14899 (N_14899,N_5290,N_9981);
or U14900 (N_14900,N_6703,N_5177);
or U14901 (N_14901,N_8844,N_6298);
xnor U14902 (N_14902,N_5669,N_5748);
or U14903 (N_14903,N_7111,N_7055);
nand U14904 (N_14904,N_5563,N_8206);
nand U14905 (N_14905,N_5842,N_5635);
nand U14906 (N_14906,N_5286,N_6135);
or U14907 (N_14907,N_7782,N_9686);
and U14908 (N_14908,N_9824,N_6729);
nand U14909 (N_14909,N_9631,N_6569);
nand U14910 (N_14910,N_8581,N_7191);
or U14911 (N_14911,N_8469,N_5370);
or U14912 (N_14912,N_5285,N_7990);
nand U14913 (N_14913,N_7356,N_8925);
and U14914 (N_14914,N_7480,N_8659);
nand U14915 (N_14915,N_5418,N_8861);
nand U14916 (N_14916,N_7442,N_7575);
or U14917 (N_14917,N_9168,N_9316);
nand U14918 (N_14918,N_8197,N_8800);
nor U14919 (N_14919,N_9220,N_9855);
or U14920 (N_14920,N_8800,N_5496);
nand U14921 (N_14921,N_9151,N_7883);
nand U14922 (N_14922,N_7612,N_7937);
nor U14923 (N_14923,N_5033,N_7480);
nor U14924 (N_14924,N_8138,N_8909);
nand U14925 (N_14925,N_8843,N_5660);
nand U14926 (N_14926,N_5341,N_8218);
and U14927 (N_14927,N_6854,N_9953);
and U14928 (N_14928,N_9790,N_5750);
xnor U14929 (N_14929,N_8692,N_8305);
xnor U14930 (N_14930,N_6781,N_7582);
nor U14931 (N_14931,N_6748,N_6998);
or U14932 (N_14932,N_9911,N_6602);
or U14933 (N_14933,N_7221,N_8908);
and U14934 (N_14934,N_6662,N_9555);
nand U14935 (N_14935,N_6215,N_5432);
and U14936 (N_14936,N_6992,N_6129);
and U14937 (N_14937,N_5557,N_9181);
nand U14938 (N_14938,N_9909,N_7458);
or U14939 (N_14939,N_5263,N_9006);
or U14940 (N_14940,N_7220,N_6203);
xor U14941 (N_14941,N_9345,N_7658);
xor U14942 (N_14942,N_8547,N_5358);
nand U14943 (N_14943,N_5216,N_7699);
or U14944 (N_14944,N_9888,N_7232);
or U14945 (N_14945,N_7571,N_7702);
xnor U14946 (N_14946,N_5699,N_9909);
nand U14947 (N_14947,N_5480,N_5917);
nor U14948 (N_14948,N_6392,N_8686);
and U14949 (N_14949,N_7588,N_7787);
nor U14950 (N_14950,N_9500,N_7425);
nor U14951 (N_14951,N_6110,N_8800);
xor U14952 (N_14952,N_9938,N_6944);
nand U14953 (N_14953,N_9666,N_8862);
xnor U14954 (N_14954,N_6203,N_8907);
nand U14955 (N_14955,N_7800,N_9514);
or U14956 (N_14956,N_8727,N_8718);
nor U14957 (N_14957,N_8778,N_8897);
or U14958 (N_14958,N_7920,N_6400);
or U14959 (N_14959,N_7090,N_8363);
or U14960 (N_14960,N_5298,N_6662);
nor U14961 (N_14961,N_9064,N_5067);
nand U14962 (N_14962,N_7924,N_8779);
nor U14963 (N_14963,N_9730,N_6751);
nand U14964 (N_14964,N_9170,N_9980);
and U14965 (N_14965,N_9982,N_8451);
and U14966 (N_14966,N_7396,N_7648);
and U14967 (N_14967,N_7395,N_8520);
nor U14968 (N_14968,N_5430,N_9125);
and U14969 (N_14969,N_7520,N_7809);
nor U14970 (N_14970,N_7294,N_5164);
nand U14971 (N_14971,N_8196,N_6916);
nand U14972 (N_14972,N_6719,N_6247);
nand U14973 (N_14973,N_9293,N_7718);
and U14974 (N_14974,N_7833,N_7001);
and U14975 (N_14975,N_6997,N_9881);
or U14976 (N_14976,N_6266,N_6476);
and U14977 (N_14977,N_9133,N_5990);
and U14978 (N_14978,N_9268,N_8544);
or U14979 (N_14979,N_5002,N_5566);
xnor U14980 (N_14980,N_6238,N_8556);
xnor U14981 (N_14981,N_6733,N_5345);
nor U14982 (N_14982,N_9647,N_9566);
nor U14983 (N_14983,N_7395,N_8252);
or U14984 (N_14984,N_6938,N_8668);
nand U14985 (N_14985,N_9236,N_8447);
or U14986 (N_14986,N_8464,N_6722);
nand U14987 (N_14987,N_9218,N_7791);
nor U14988 (N_14988,N_5471,N_8577);
or U14989 (N_14989,N_5284,N_9001);
nand U14990 (N_14990,N_7946,N_6310);
nor U14991 (N_14991,N_8259,N_8195);
or U14992 (N_14992,N_8950,N_7838);
and U14993 (N_14993,N_7379,N_9678);
nand U14994 (N_14994,N_5512,N_9985);
xor U14995 (N_14995,N_8090,N_7399);
or U14996 (N_14996,N_8388,N_6085);
and U14997 (N_14997,N_7478,N_9488);
and U14998 (N_14998,N_9787,N_7488);
or U14999 (N_14999,N_8406,N_9858);
nand UO_0 (O_0,N_11938,N_13133);
and UO_1 (O_1,N_10124,N_10029);
nand UO_2 (O_2,N_10201,N_12926);
nor UO_3 (O_3,N_10241,N_12083);
or UO_4 (O_4,N_11559,N_13071);
or UO_5 (O_5,N_11979,N_11891);
and UO_6 (O_6,N_14935,N_11416);
xor UO_7 (O_7,N_13452,N_13809);
nor UO_8 (O_8,N_10839,N_10525);
nand UO_9 (O_9,N_13019,N_11266);
nor UO_10 (O_10,N_14793,N_10361);
and UO_11 (O_11,N_13598,N_11111);
nor UO_12 (O_12,N_10588,N_11787);
nand UO_13 (O_13,N_10375,N_13514);
and UO_14 (O_14,N_11428,N_14806);
xor UO_15 (O_15,N_12437,N_10501);
nor UO_16 (O_16,N_11620,N_14158);
or UO_17 (O_17,N_11810,N_11526);
or UO_18 (O_18,N_11451,N_14223);
or UO_19 (O_19,N_14985,N_14212);
and UO_20 (O_20,N_14361,N_13747);
nor UO_21 (O_21,N_12917,N_11060);
nor UO_22 (O_22,N_12744,N_13474);
and UO_23 (O_23,N_13880,N_13265);
or UO_24 (O_24,N_13412,N_11755);
and UO_25 (O_25,N_13640,N_13571);
nand UO_26 (O_26,N_11418,N_13688);
and UO_27 (O_27,N_11550,N_14026);
nand UO_28 (O_28,N_10044,N_13009);
nand UO_29 (O_29,N_11320,N_12497);
nor UO_30 (O_30,N_14242,N_11676);
nand UO_31 (O_31,N_10846,N_13173);
nor UO_32 (O_32,N_13006,N_14017);
nand UO_33 (O_33,N_11095,N_10554);
and UO_34 (O_34,N_14251,N_11900);
nor UO_35 (O_35,N_12305,N_13738);
or UO_36 (O_36,N_13287,N_12820);
nor UO_37 (O_37,N_12873,N_14481);
nand UO_38 (O_38,N_10366,N_12197);
nand UO_39 (O_39,N_13953,N_10833);
nor UO_40 (O_40,N_13303,N_12043);
nor UO_41 (O_41,N_10317,N_11818);
and UO_42 (O_42,N_14829,N_12075);
xnor UO_43 (O_43,N_13084,N_10357);
or UO_44 (O_44,N_11823,N_10632);
or UO_45 (O_45,N_14079,N_12021);
or UO_46 (O_46,N_14678,N_11785);
or UO_47 (O_47,N_11606,N_11403);
and UO_48 (O_48,N_14204,N_10172);
nor UO_49 (O_49,N_13035,N_14392);
nor UO_50 (O_50,N_14743,N_13448);
nand UO_51 (O_51,N_11975,N_11086);
or UO_52 (O_52,N_13352,N_10113);
xor UO_53 (O_53,N_13537,N_12832);
or UO_54 (O_54,N_13965,N_14731);
nand UO_55 (O_55,N_14000,N_10011);
or UO_56 (O_56,N_13915,N_11328);
and UO_57 (O_57,N_10030,N_13193);
nor UO_58 (O_58,N_13120,N_10774);
or UO_59 (O_59,N_10580,N_11674);
nand UO_60 (O_60,N_10252,N_10021);
nor UO_61 (O_61,N_10876,N_11410);
nand UO_62 (O_62,N_14162,N_13758);
or UO_63 (O_63,N_11472,N_12470);
or UO_64 (O_64,N_10305,N_10165);
and UO_65 (O_65,N_13468,N_11064);
nor UO_66 (O_66,N_14578,N_10147);
or UO_67 (O_67,N_14009,N_13842);
or UO_68 (O_68,N_13430,N_10890);
nor UO_69 (O_69,N_12971,N_10077);
or UO_70 (O_70,N_11133,N_12833);
and UO_71 (O_71,N_13914,N_14813);
xnor UO_72 (O_72,N_14291,N_14659);
and UO_73 (O_73,N_14488,N_12204);
xnor UO_74 (O_74,N_12830,N_10692);
or UO_75 (O_75,N_11523,N_11276);
nor UO_76 (O_76,N_14238,N_13581);
nand UO_77 (O_77,N_12297,N_13821);
or UO_78 (O_78,N_11866,N_10962);
nor UO_79 (O_79,N_13093,N_11951);
or UO_80 (O_80,N_10001,N_12367);
xnor UO_81 (O_81,N_13671,N_12855);
nand UO_82 (O_82,N_12153,N_14496);
xnor UO_83 (O_83,N_13388,N_13270);
nand UO_84 (O_84,N_10797,N_10205);
or UO_85 (O_85,N_10488,N_13941);
or UO_86 (O_86,N_12239,N_14747);
nor UO_87 (O_87,N_13852,N_11300);
and UO_88 (O_88,N_14343,N_12062);
xnor UO_89 (O_89,N_14145,N_13207);
and UO_90 (O_90,N_11074,N_12532);
or UO_91 (O_91,N_12656,N_12608);
nor UO_92 (O_92,N_13716,N_14202);
nand UO_93 (O_93,N_14833,N_13470);
or UO_94 (O_94,N_11983,N_10384);
nand UO_95 (O_95,N_14548,N_11008);
nand UO_96 (O_96,N_11994,N_12945);
nand UO_97 (O_97,N_10593,N_14781);
and UO_98 (O_98,N_11654,N_13000);
nor UO_99 (O_99,N_12427,N_12277);
or UO_100 (O_100,N_14575,N_10302);
nand UO_101 (O_101,N_14058,N_13961);
nor UO_102 (O_102,N_12316,N_14825);
nor UO_103 (O_103,N_11119,N_12911);
nand UO_104 (O_104,N_11690,N_14459);
or UO_105 (O_105,N_12867,N_14433);
nand UO_106 (O_106,N_12835,N_11644);
and UO_107 (O_107,N_13551,N_10489);
nor UO_108 (O_108,N_11597,N_14429);
nor UO_109 (O_109,N_14537,N_12963);
and UO_110 (O_110,N_11360,N_12184);
and UO_111 (O_111,N_12872,N_13310);
or UO_112 (O_112,N_13808,N_12604);
nand UO_113 (O_113,N_13580,N_11520);
nor UO_114 (O_114,N_11100,N_12482);
or UO_115 (O_115,N_11960,N_11429);
nand UO_116 (O_116,N_14556,N_14335);
and UO_117 (O_117,N_12851,N_13724);
nand UO_118 (O_118,N_14258,N_12233);
and UO_119 (O_119,N_13905,N_10997);
and UO_120 (O_120,N_12560,N_12008);
or UO_121 (O_121,N_10280,N_11933);
and UO_122 (O_122,N_12568,N_10415);
and UO_123 (O_123,N_10903,N_14667);
nand UO_124 (O_124,N_12457,N_10943);
and UO_125 (O_125,N_10281,N_10836);
or UO_126 (O_126,N_12077,N_10119);
nor UO_127 (O_127,N_10288,N_11725);
nor UO_128 (O_128,N_10822,N_10636);
or UO_129 (O_129,N_13423,N_14783);
or UO_130 (O_130,N_14755,N_12230);
and UO_131 (O_131,N_10518,N_14155);
nand UO_132 (O_132,N_12397,N_14854);
and UO_133 (O_133,N_11030,N_12773);
or UO_134 (O_134,N_12871,N_14601);
nand UO_135 (O_135,N_13204,N_13404);
nand UO_136 (O_136,N_12190,N_11660);
and UO_137 (O_137,N_12319,N_11368);
nor UO_138 (O_138,N_14734,N_10958);
nor UO_139 (O_139,N_12035,N_10996);
nand UO_140 (O_140,N_12157,N_13554);
or UO_141 (O_141,N_11105,N_14776);
nor UO_142 (O_142,N_12399,N_13179);
nand UO_143 (O_143,N_12813,N_11208);
and UO_144 (O_144,N_10671,N_12811);
and UO_145 (O_145,N_10637,N_14549);
nand UO_146 (O_146,N_10666,N_14246);
nand UO_147 (O_147,N_13160,N_13703);
xnor UO_148 (O_148,N_13261,N_10910);
nand UO_149 (O_149,N_14053,N_11804);
nor UO_150 (O_150,N_11342,N_12022);
and UO_151 (O_151,N_13523,N_13393);
and UO_152 (O_152,N_13814,N_14217);
xnor UO_153 (O_153,N_13075,N_14638);
nand UO_154 (O_154,N_11466,N_11189);
and UO_155 (O_155,N_13651,N_10279);
and UO_156 (O_156,N_11009,N_11640);
nand UO_157 (O_157,N_12671,N_12693);
xor UO_158 (O_158,N_14919,N_13024);
or UO_159 (O_159,N_14722,N_14338);
or UO_160 (O_160,N_11110,N_14860);
and UO_161 (O_161,N_12617,N_11781);
nor UO_162 (O_162,N_12267,N_14619);
or UO_163 (O_163,N_12764,N_11291);
nor UO_164 (O_164,N_10649,N_11565);
nor UO_165 (O_165,N_13951,N_14893);
or UO_166 (O_166,N_12439,N_12025);
nand UO_167 (O_167,N_11683,N_10176);
nand UO_168 (O_168,N_13039,N_11691);
nor UO_169 (O_169,N_11874,N_14666);
and UO_170 (O_170,N_10466,N_10523);
nor UO_171 (O_171,N_14405,N_13123);
nor UO_172 (O_172,N_10059,N_13807);
or UO_173 (O_173,N_13685,N_12026);
nand UO_174 (O_174,N_12189,N_11831);
or UO_175 (O_175,N_11058,N_13455);
and UO_176 (O_176,N_13140,N_12970);
or UO_177 (O_177,N_14080,N_10827);
and UO_178 (O_178,N_13232,N_12335);
nand UO_179 (O_179,N_14802,N_14931);
nor UO_180 (O_180,N_12440,N_11098);
or UO_181 (O_181,N_14224,N_10834);
and UO_182 (O_182,N_14800,N_13426);
nand UO_183 (O_183,N_14305,N_14206);
nand UO_184 (O_184,N_11706,N_11446);
and UO_185 (O_185,N_10605,N_14400);
nand UO_186 (O_186,N_10633,N_14271);
nand UO_187 (O_187,N_11404,N_13519);
and UO_188 (O_188,N_14452,N_13712);
or UO_189 (O_189,N_14623,N_12716);
or UO_190 (O_190,N_10584,N_10849);
or UO_191 (O_191,N_10283,N_11204);
nor UO_192 (O_192,N_14780,N_13366);
nor UO_193 (O_193,N_14140,N_12962);
and UO_194 (O_194,N_13332,N_12674);
nand UO_195 (O_195,N_12048,N_12868);
xor UO_196 (O_196,N_14131,N_12073);
or UO_197 (O_197,N_12850,N_11921);
or UO_198 (O_198,N_14352,N_13679);
nand UO_199 (O_199,N_10611,N_14418);
nor UO_200 (O_200,N_14877,N_11247);
nor UO_201 (O_201,N_12332,N_14236);
xor UO_202 (O_202,N_14989,N_10899);
nand UO_203 (O_203,N_12139,N_10779);
nor UO_204 (O_204,N_14292,N_13141);
nor UO_205 (O_205,N_12389,N_10679);
or UO_206 (O_206,N_13048,N_10186);
nand UO_207 (O_207,N_14089,N_12195);
nor UO_208 (O_208,N_14968,N_12169);
or UO_209 (O_209,N_13343,N_11528);
nand UO_210 (O_210,N_13175,N_12713);
or UO_211 (O_211,N_13734,N_10703);
and UO_212 (O_212,N_10957,N_10093);
or UO_213 (O_213,N_13478,N_14501);
nand UO_214 (O_214,N_12018,N_11500);
nand UO_215 (O_215,N_14830,N_11414);
xor UO_216 (O_216,N_14748,N_14999);
or UO_217 (O_217,N_14336,N_10456);
or UO_218 (O_218,N_13198,N_11199);
or UO_219 (O_219,N_11799,N_12187);
or UO_220 (O_220,N_14859,N_11575);
or UO_221 (O_221,N_10723,N_10018);
nor UO_222 (O_222,N_14589,N_10801);
nand UO_223 (O_223,N_10949,N_14113);
or UO_224 (O_224,N_13991,N_12802);
or UO_225 (O_225,N_12033,N_13907);
xor UO_226 (O_226,N_14446,N_11758);
and UO_227 (O_227,N_10669,N_14998);
or UO_228 (O_228,N_10812,N_11637);
nor UO_229 (O_229,N_10835,N_11426);
or UO_230 (O_230,N_11635,N_12434);
or UO_231 (O_231,N_12063,N_14043);
or UO_232 (O_232,N_11335,N_11498);
and UO_233 (O_233,N_14333,N_14592);
and UO_234 (O_234,N_14035,N_14144);
and UO_235 (O_235,N_14448,N_14901);
nor UO_236 (O_236,N_11778,N_13078);
or UO_237 (O_237,N_14094,N_12141);
nand UO_238 (O_238,N_10054,N_13859);
and UO_239 (O_239,N_11570,N_12113);
and UO_240 (O_240,N_11090,N_10098);
nand UO_241 (O_241,N_14492,N_13956);
nor UO_242 (O_242,N_11892,N_11936);
nor UO_243 (O_243,N_14453,N_12624);
or UO_244 (O_244,N_14346,N_10096);
nand UO_245 (O_245,N_14234,N_14288);
and UO_246 (O_246,N_10739,N_10749);
or UO_247 (O_247,N_14134,N_14318);
nor UO_248 (O_248,N_13829,N_13566);
xor UO_249 (O_249,N_10751,N_11152);
or UO_250 (O_250,N_13913,N_11883);
or UO_251 (O_251,N_13759,N_11494);
or UO_252 (O_252,N_10852,N_10531);
and UO_253 (O_253,N_13999,N_10437);
nor UO_254 (O_254,N_12422,N_13016);
nand UO_255 (O_255,N_14777,N_12742);
and UO_256 (O_256,N_14220,N_11529);
or UO_257 (O_257,N_12535,N_13674);
nor UO_258 (O_258,N_12552,N_12756);
or UO_259 (O_259,N_13678,N_12780);
and UO_260 (O_260,N_13320,N_11041);
xor UO_261 (O_261,N_13329,N_14386);
and UO_262 (O_262,N_13378,N_13397);
and UO_263 (O_263,N_10148,N_10304);
or UO_264 (O_264,N_11470,N_12673);
nand UO_265 (O_265,N_11474,N_10537);
or UO_266 (O_266,N_14827,N_10952);
and UO_267 (O_267,N_13459,N_13108);
nor UO_268 (O_268,N_14595,N_10706);
nand UO_269 (O_269,N_11516,N_12613);
or UO_270 (O_270,N_10869,N_11845);
or UO_271 (O_271,N_14583,N_13288);
and UO_272 (O_272,N_12899,N_14172);
or UO_273 (O_273,N_13544,N_12585);
nand UO_274 (O_274,N_11696,N_11768);
xor UO_275 (O_275,N_11720,N_13973);
nand UO_276 (O_276,N_10575,N_11519);
or UO_277 (O_277,N_14821,N_11774);
nand UO_278 (O_278,N_13063,N_14653);
nand UO_279 (O_279,N_11971,N_11742);
nand UO_280 (O_280,N_10735,N_12089);
xor UO_281 (O_281,N_11760,N_12969);
nor UO_282 (O_282,N_11407,N_13543);
and UO_283 (O_283,N_13906,N_12255);
xor UO_284 (O_284,N_13153,N_11260);
and UO_285 (O_285,N_12291,N_14628);
or UO_286 (O_286,N_12584,N_11135);
and UO_287 (O_287,N_12100,N_11566);
nand UO_288 (O_288,N_12738,N_13233);
or UO_289 (O_289,N_11532,N_13978);
and UO_290 (O_290,N_10911,N_12056);
xor UO_291 (O_291,N_10259,N_12896);
or UO_292 (O_292,N_12476,N_14873);
nand UO_293 (O_293,N_11980,N_10106);
nor UO_294 (O_294,N_11997,N_12375);
or UO_295 (O_295,N_14772,N_12629);
and UO_296 (O_296,N_13383,N_12946);
and UO_297 (O_297,N_10771,N_11383);
or UO_298 (O_298,N_11314,N_13838);
nor UO_299 (O_299,N_13803,N_11744);
nand UO_300 (O_300,N_14988,N_14347);
nand UO_301 (O_301,N_12317,N_13341);
nor UO_302 (O_302,N_12829,N_13846);
and UO_303 (O_303,N_10121,N_14315);
xnor UO_304 (O_304,N_12420,N_10604);
nor UO_305 (O_305,N_14792,N_12270);
xor UO_306 (O_306,N_11370,N_13602);
nand UO_307 (O_307,N_13300,N_14366);
and UO_308 (O_308,N_10495,N_14752);
nand UO_309 (O_309,N_14099,N_13825);
and UO_310 (O_310,N_12014,N_12898);
nor UO_311 (O_311,N_10104,N_14624);
and UO_312 (O_312,N_14164,N_10837);
nor UO_313 (O_313,N_13305,N_10556);
nor UO_314 (O_314,N_13606,N_10482);
or UO_315 (O_315,N_14816,N_13656);
and UO_316 (O_316,N_14281,N_12009);
xnor UO_317 (O_317,N_13599,N_14329);
xnor UO_318 (O_318,N_10975,N_10491);
nor UO_319 (O_319,N_12134,N_14279);
nor UO_320 (O_320,N_11684,N_14907);
nand UO_321 (O_321,N_14963,N_14439);
nor UO_322 (O_322,N_10236,N_10700);
and UO_323 (O_323,N_14550,N_12181);
and UO_324 (O_324,N_13542,N_10450);
xnor UO_325 (O_325,N_13345,N_13782);
nand UO_326 (O_326,N_13684,N_14194);
and UO_327 (O_327,N_11766,N_13466);
nand UO_328 (O_328,N_12264,N_14528);
nand UO_329 (O_329,N_10233,N_12750);
nor UO_330 (O_330,N_12555,N_14904);
nand UO_331 (O_331,N_10057,N_13159);
nor UO_332 (O_332,N_10813,N_14403);
nor UO_333 (O_333,N_10691,N_14729);
and UO_334 (O_334,N_13647,N_13109);
nand UO_335 (O_335,N_11540,N_11968);
or UO_336 (O_336,N_14739,N_11844);
nand UO_337 (O_337,N_10938,N_14141);
nand UO_338 (O_338,N_11857,N_11029);
and UO_339 (O_339,N_14953,N_10820);
xor UO_340 (O_340,N_14690,N_14054);
nor UO_341 (O_341,N_14148,N_10453);
nor UO_342 (O_342,N_12236,N_11107);
and UO_343 (O_343,N_12357,N_11807);
nor UO_344 (O_344,N_11382,N_13411);
xor UO_345 (O_345,N_14074,N_11927);
xnor UO_346 (O_346,N_10253,N_12206);
xnor UO_347 (O_347,N_12921,N_10896);
or UO_348 (O_348,N_14178,N_11339);
and UO_349 (O_349,N_11033,N_11480);
nor UO_350 (O_350,N_10931,N_12124);
and UO_351 (O_351,N_11607,N_10320);
nor UO_352 (O_352,N_14375,N_11609);
nand UO_353 (O_353,N_14709,N_14925);
nor UO_354 (O_354,N_13046,N_13550);
or UO_355 (O_355,N_13711,N_10239);
or UO_356 (O_356,N_10249,N_14817);
nor UO_357 (O_357,N_10509,N_11424);
or UO_358 (O_358,N_12681,N_12976);
or UO_359 (O_359,N_14264,N_13218);
xnor UO_360 (O_360,N_12350,N_12165);
xor UO_361 (O_361,N_14196,N_12462);
nand UO_362 (O_362,N_14645,N_14487);
nor UO_363 (O_363,N_13936,N_14654);
or UO_364 (O_364,N_12531,N_14368);
nand UO_365 (O_365,N_10055,N_12133);
or UO_366 (O_366,N_10514,N_14055);
nor UO_367 (O_367,N_12839,N_11154);
nand UO_368 (O_368,N_12289,N_12732);
or UO_369 (O_369,N_11859,N_13802);
and UO_370 (O_370,N_10309,N_10325);
and UO_371 (O_371,N_12965,N_12513);
or UO_372 (O_372,N_11993,N_10327);
xnor UO_373 (O_373,N_13146,N_12372);
and UO_374 (O_374,N_14317,N_13137);
and UO_375 (O_375,N_10994,N_12566);
and UO_376 (O_376,N_14658,N_13178);
nor UO_377 (O_377,N_12620,N_11765);
nor UO_378 (O_378,N_10326,N_10108);
nand UO_379 (O_379,N_10284,N_11651);
and UO_380 (O_380,N_13603,N_13805);
and UO_381 (O_381,N_14489,N_10944);
xor UO_382 (O_382,N_14930,N_14351);
or UO_383 (O_383,N_10356,N_14419);
xor UO_384 (O_384,N_11602,N_13768);
or UO_385 (O_385,N_12046,N_12477);
and UO_386 (O_386,N_11294,N_13186);
and UO_387 (O_387,N_10404,N_11564);
nor UO_388 (O_388,N_12808,N_12699);
xnor UO_389 (O_389,N_14805,N_14615);
nor UO_390 (O_390,N_12246,N_11121);
and UO_391 (O_391,N_10369,N_14661);
or UO_392 (O_392,N_14215,N_10647);
nor UO_393 (O_393,N_12524,N_11037);
nand UO_394 (O_394,N_12545,N_11327);
and UO_395 (O_395,N_14233,N_12171);
and UO_396 (O_396,N_11379,N_10673);
or UO_397 (O_397,N_10906,N_12985);
nor UO_398 (O_398,N_10135,N_13552);
nor UO_399 (O_399,N_12663,N_13811);
and UO_400 (O_400,N_11759,N_13988);
xnor UO_401 (O_401,N_10208,N_11272);
nand UO_402 (O_402,N_13432,N_14334);
nand UO_403 (O_403,N_11485,N_14852);
or UO_404 (O_404,N_11065,N_11228);
xnor UO_405 (O_405,N_12792,N_13481);
nor UO_406 (O_406,N_13385,N_11202);
nand UO_407 (O_407,N_13219,N_13769);
xor UO_408 (O_408,N_10376,N_12458);
and UO_409 (O_409,N_14296,N_13401);
nand UO_410 (O_410,N_12052,N_11603);
and UO_411 (O_411,N_13083,N_13832);
nor UO_412 (O_412,N_12842,N_11045);
and UO_413 (O_413,N_13636,N_14869);
xnor UO_414 (O_414,N_13056,N_11371);
and UO_415 (O_415,N_12146,N_13621);
nand UO_416 (O_416,N_11307,N_14557);
nand UO_417 (O_417,N_10885,N_13793);
nand UO_418 (O_418,N_13624,N_14253);
xor UO_419 (O_419,N_12130,N_14521);
or UO_420 (O_420,N_11180,N_10040);
nand UO_421 (O_421,N_12569,N_11634);
or UO_422 (O_422,N_11506,N_13834);
and UO_423 (O_423,N_12910,N_12484);
nand UO_424 (O_424,N_14129,N_12064);
and UO_425 (O_425,N_10503,N_13041);
and UO_426 (O_426,N_11162,N_12161);
nand UO_427 (O_427,N_14710,N_13997);
and UO_428 (O_428,N_10550,N_14715);
nand UO_429 (O_429,N_13791,N_13979);
xnor UO_430 (O_430,N_12730,N_11944);
nand UO_431 (O_431,N_14834,N_10155);
and UO_432 (O_432,N_10053,N_12004);
or UO_433 (O_433,N_12186,N_13344);
xnor UO_434 (O_434,N_10478,N_13148);
and UO_435 (O_435,N_13276,N_11636);
or UO_436 (O_436,N_12346,N_13515);
xnor UO_437 (O_437,N_11286,N_14200);
nand UO_438 (O_438,N_11776,N_13528);
xnor UO_439 (O_439,N_11226,N_13823);
nor UO_440 (O_440,N_12991,N_14276);
and UO_441 (O_441,N_13620,N_12232);
or UO_442 (O_442,N_12456,N_14316);
nand UO_443 (O_443,N_13086,N_13097);
nand UO_444 (O_444,N_11326,N_11297);
nor UO_445 (O_445,N_11561,N_10821);
xor UO_446 (O_446,N_11109,N_14727);
nand UO_447 (O_447,N_11793,N_14498);
and UO_448 (O_448,N_10222,N_12968);
nand UO_449 (O_449,N_12554,N_13949);
nand UO_450 (O_450,N_12770,N_10661);
or UO_451 (O_451,N_11806,N_11200);
nand UO_452 (O_452,N_10504,N_12448);
or UO_453 (O_453,N_11377,N_11843);
and UO_454 (O_454,N_12743,N_10371);
xor UO_455 (O_455,N_10672,N_11643);
or UO_456 (O_456,N_10736,N_11885);
nand UO_457 (O_457,N_11471,N_11157);
nor UO_458 (O_458,N_10829,N_12015);
nand UO_459 (O_459,N_13280,N_11233);
nand UO_460 (O_460,N_13837,N_13082);
and UO_461 (O_461,N_12809,N_11128);
nor UO_462 (O_462,N_13057,N_12374);
and UO_463 (O_463,N_12559,N_14533);
nor UO_464 (O_464,N_12818,N_10347);
or UO_465 (O_465,N_11458,N_10122);
or UO_466 (O_466,N_12402,N_10577);
and UO_467 (O_467,N_14568,N_14637);
xor UO_468 (O_468,N_14245,N_13313);
nand UO_469 (O_469,N_13434,N_10825);
nand UO_470 (O_470,N_12522,N_14044);
and UO_471 (O_471,N_10085,N_14294);
or UO_472 (O_472,N_12533,N_11417);
or UO_473 (O_473,N_13536,N_13336);
and UO_474 (O_474,N_13861,N_13594);
nand UO_475 (O_475,N_11860,N_13980);
and UO_476 (O_476,N_13080,N_14938);
nand UO_477 (O_477,N_12953,N_14010);
or UO_478 (O_478,N_10877,N_11647);
nand UO_479 (O_479,N_12769,N_11246);
xnor UO_480 (O_480,N_11223,N_13690);
nand UO_481 (O_481,N_11423,N_11488);
or UO_482 (O_482,N_14552,N_12979);
nand UO_483 (O_483,N_14289,N_12074);
xnor UO_484 (O_484,N_10479,N_11349);
xor UO_485 (O_485,N_12821,N_14273);
and UO_486 (O_486,N_10436,N_14714);
and UO_487 (O_487,N_10770,N_11605);
nor UO_488 (O_488,N_12478,N_13185);
nor UO_489 (O_489,N_10712,N_13076);
and UO_490 (O_490,N_14219,N_11836);
nor UO_491 (O_491,N_13167,N_14304);
nand UO_492 (O_492,N_11131,N_12084);
nor UO_493 (O_493,N_13909,N_13069);
xnor UO_494 (O_494,N_14889,N_11555);
nand UO_495 (O_495,N_10791,N_11315);
xor UO_496 (O_496,N_12589,N_12473);
nand UO_497 (O_497,N_10526,N_10291);
nand UO_498 (O_498,N_14840,N_13492);
and UO_499 (O_499,N_11650,N_13587);
xor UO_500 (O_500,N_14390,N_14861);
nor UO_501 (O_501,N_11478,N_12231);
or UO_502 (O_502,N_13694,N_13822);
nand UO_503 (O_503,N_11415,N_12597);
nand UO_504 (O_504,N_10354,N_13529);
nor UO_505 (O_505,N_12208,N_11489);
nand UO_506 (O_506,N_13673,N_10684);
nor UO_507 (O_507,N_12712,N_12602);
and UO_508 (O_508,N_11576,N_10146);
nor UO_509 (O_509,N_13943,N_14365);
xnor UO_510 (O_510,N_10854,N_12329);
and UO_511 (O_511,N_14339,N_12237);
nand UO_512 (O_512,N_12327,N_12574);
nand UO_513 (O_513,N_12326,N_11973);
or UO_514 (O_514,N_11206,N_14341);
nor UO_515 (O_515,N_11491,N_14187);
and UO_516 (O_516,N_13263,N_11829);
or UO_517 (O_517,N_13067,N_12283);
or UO_518 (O_518,N_10708,N_13172);
nand UO_519 (O_519,N_13004,N_10111);
and UO_520 (O_520,N_13256,N_12626);
nor UO_521 (O_521,N_14451,N_12942);
nor UO_522 (O_522,N_10151,N_14263);
and UO_523 (O_523,N_13142,N_12651);
nor UO_524 (O_524,N_10467,N_14928);
nand UO_525 (O_525,N_14767,N_13894);
nor UO_526 (O_526,N_11612,N_10432);
nor UO_527 (O_527,N_14945,N_10138);
nor UO_528 (O_528,N_10271,N_14763);
or UO_529 (O_529,N_13743,N_14944);
and UO_530 (O_530,N_10941,N_12262);
xnor UO_531 (O_531,N_13015,N_12708);
and UO_532 (O_532,N_14048,N_13446);
and UO_533 (O_533,N_11256,N_14555);
and UO_534 (O_534,N_14216,N_10710);
nor UO_535 (O_535,N_12772,N_10099);
xor UO_536 (O_536,N_11723,N_12040);
or UO_537 (O_537,N_10228,N_10103);
nand UO_538 (O_538,N_10884,N_13563);
nand UO_539 (O_539,N_13469,N_12486);
nor UO_540 (O_540,N_11782,N_10315);
or UO_541 (O_541,N_11868,N_13221);
or UO_542 (O_542,N_10844,N_14894);
nand UO_543 (O_543,N_11147,N_13972);
xor UO_544 (O_544,N_14167,N_12810);
nand UO_545 (O_545,N_14331,N_14831);
nand UO_546 (O_546,N_12118,N_12775);
or UO_547 (O_547,N_13777,N_13224);
nand UO_548 (O_548,N_11117,N_10999);
nor UO_549 (O_549,N_12313,N_13740);
xnor UO_550 (O_550,N_13760,N_10069);
or UO_551 (O_551,N_12205,N_11897);
or UO_552 (O_552,N_10757,N_14847);
or UO_553 (O_553,N_13477,N_13876);
nand UO_554 (O_554,N_12692,N_14337);
nand UO_555 (O_555,N_11299,N_14559);
or UO_556 (O_556,N_11321,N_13228);
nor UO_557 (O_557,N_11132,N_13693);
or UO_558 (O_558,N_13525,N_11185);
or UO_559 (O_559,N_14116,N_13670);
nor UO_560 (O_560,N_10777,N_14038);
nor UO_561 (O_561,N_14593,N_14128);
or UO_562 (O_562,N_11739,N_10902);
nand UO_563 (O_563,N_14076,N_11225);
nor UO_564 (O_564,N_10071,N_10979);
xor UO_565 (O_565,N_12664,N_10359);
nand UO_566 (O_566,N_13170,N_13463);
and UO_567 (O_567,N_11499,N_11882);
and UO_568 (O_568,N_10330,N_11187);
nand UO_569 (O_569,N_14648,N_14891);
nand UO_570 (O_570,N_12644,N_11655);
nor UO_571 (O_571,N_12031,N_11067);
nor UO_572 (O_572,N_11412,N_14540);
and UO_573 (O_573,N_10628,N_11275);
nand UO_574 (O_574,N_13903,N_12481);
nor UO_575 (O_575,N_12902,N_10221);
nand UO_576 (O_576,N_14240,N_11497);
and UO_577 (O_577,N_12616,N_11894);
nand UO_578 (O_578,N_14256,N_13169);
nor UO_579 (O_579,N_10709,N_13735);
nand UO_580 (O_580,N_12480,N_14340);
nor UO_581 (O_581,N_11948,N_12269);
nor UO_582 (O_582,N_11369,N_12178);
or UO_583 (O_583,N_12284,N_14031);
and UO_584 (O_584,N_14929,N_11167);
and UO_585 (O_585,N_10007,N_13974);
nor UO_586 (O_586,N_14406,N_13072);
nand UO_587 (O_587,N_14049,N_10272);
or UO_588 (O_588,N_14912,N_10412);
nand UO_589 (O_589,N_10303,N_11183);
or UO_590 (O_590,N_14151,N_12786);
nand UO_591 (O_591,N_13127,N_10769);
nand UO_592 (O_592,N_11939,N_12342);
nor UO_593 (O_593,N_12132,N_11838);
nand UO_594 (O_594,N_14896,N_10349);
nor UO_595 (O_595,N_13722,N_10483);
nor UO_596 (O_596,N_11141,N_10244);
or UO_597 (O_597,N_12224,N_13707);
or UO_598 (O_598,N_13509,N_13297);
nor UO_599 (O_599,N_14958,N_12330);
and UO_600 (O_600,N_10145,N_12200);
nand UO_601 (O_601,N_13680,N_14464);
nor UO_602 (O_602,N_12121,N_14431);
or UO_603 (O_603,N_14310,N_11702);
nand UO_604 (O_604,N_14460,N_13683);
or UO_605 (O_605,N_10275,N_12667);
nand UO_606 (O_606,N_14632,N_13454);
nor UO_607 (O_607,N_11815,N_14278);
or UO_608 (O_608,N_12304,N_13848);
and UO_609 (O_609,N_11018,N_10982);
or UO_610 (O_610,N_11083,N_14190);
and UO_611 (O_611,N_11005,N_12956);
nand UO_612 (O_612,N_13933,N_14819);
nor UO_613 (O_613,N_14878,N_12210);
nor UO_614 (O_614,N_11261,N_11905);
nor UO_615 (O_615,N_14975,N_10718);
or UO_616 (O_616,N_13853,N_13723);
and UO_617 (O_617,N_11981,N_11234);
nand UO_618 (O_618,N_14790,N_12272);
nor UO_619 (O_619,N_12883,N_13847);
or UO_620 (O_620,N_10298,N_11062);
or UO_621 (O_621,N_13149,N_11704);
nor UO_622 (O_622,N_13900,N_10819);
and UO_623 (O_623,N_14588,N_13435);
and UO_624 (O_624,N_10072,N_11068);
nand UO_625 (O_625,N_14036,N_11169);
nor UO_626 (O_626,N_14574,N_11669);
nor UO_627 (O_627,N_13761,N_11752);
or UO_628 (O_628,N_11194,N_12551);
nand UO_629 (O_629,N_13418,N_11950);
xor UO_630 (O_630,N_14319,N_10548);
or UO_631 (O_631,N_14458,N_13666);
nand UO_632 (O_632,N_11646,N_11854);
and UO_633 (O_633,N_13151,N_12594);
nand UO_634 (O_634,N_10032,N_11337);
or UO_635 (O_635,N_13596,N_13574);
nand UO_636 (O_636,N_10864,N_10573);
and UO_637 (O_637,N_14964,N_10170);
nand UO_638 (O_638,N_12907,N_13471);
or UO_639 (O_639,N_14378,N_11826);
or UO_640 (O_640,N_13567,N_14539);
or UO_641 (O_641,N_11732,N_12405);
and UO_642 (O_642,N_13538,N_14135);
or UO_643 (O_643,N_13349,N_10560);
or UO_644 (O_644,N_13714,N_13251);
xnor UO_645 (O_645,N_10845,N_12977);
nor UO_646 (O_646,N_10793,N_13533);
nand UO_647 (O_647,N_14222,N_12690);
xnor UO_648 (O_648,N_11663,N_13362);
and UO_649 (O_649,N_10150,N_11136);
nor UO_650 (O_650,N_12752,N_10727);
or UO_651 (O_651,N_13145,N_14607);
and UO_652 (O_652,N_11237,N_14669);
or UO_653 (O_653,N_12142,N_13330);
and UO_654 (O_654,N_13517,N_14411);
nand UO_655 (O_655,N_13260,N_12331);
or UO_656 (O_656,N_10760,N_11440);
or UO_657 (O_657,N_10363,N_13271);
nand UO_658 (O_658,N_12918,N_11244);
nor UO_659 (O_659,N_12353,N_12155);
nand UO_660 (O_660,N_10031,N_10024);
or UO_661 (O_661,N_13867,N_10973);
or UO_662 (O_662,N_11639,N_12085);
nand UO_663 (O_663,N_10395,N_12846);
nor UO_664 (O_664,N_10675,N_10392);
or UO_665 (O_665,N_14857,N_10986);
nor UO_666 (O_666,N_11552,N_12650);
nand UO_667 (O_667,N_13014,N_13302);
nand UO_668 (O_668,N_14456,N_13750);
or UO_669 (O_669,N_10956,N_11192);
or UO_670 (O_670,N_11087,N_12392);
nor UO_671 (O_671,N_11503,N_12930);
nand UO_672 (O_672,N_10566,N_11775);
nor UO_673 (O_673,N_10694,N_14454);
and UO_674 (O_674,N_14387,N_14171);
nand UO_675 (O_675,N_14905,N_13025);
or UO_676 (O_676,N_12993,N_12365);
nor UO_677 (O_677,N_13018,N_12665);
nor UO_678 (O_678,N_13431,N_12707);
or UO_679 (O_679,N_13700,N_11103);
or UO_680 (O_680,N_10179,N_12220);
nand UO_681 (O_681,N_11205,N_11372);
xnor UO_682 (O_682,N_14479,N_12463);
or UO_683 (O_683,N_11301,N_10803);
nand UO_684 (O_684,N_13012,N_12094);
nand UO_685 (O_685,N_10762,N_11140);
or UO_686 (O_686,N_11746,N_14656);
nand UO_687 (O_687,N_11513,N_11317);
and UO_688 (O_688,N_14868,N_11071);
or UO_689 (O_689,N_14703,N_14413);
xnor UO_690 (O_690,N_13922,N_13795);
or UO_691 (O_691,N_12779,N_12527);
nor UO_692 (O_692,N_14573,N_12279);
nor UO_693 (O_693,N_12998,N_10458);
nor UO_694 (O_694,N_12514,N_13495);
nand UO_695 (O_695,N_13994,N_14770);
and UO_696 (O_696,N_14762,N_11391);
nand UO_697 (O_697,N_14922,N_11539);
or UO_698 (O_698,N_12000,N_12906);
or UO_699 (O_699,N_10160,N_14828);
nor UO_700 (O_700,N_11687,N_11334);
nand UO_701 (O_701,N_14143,N_10895);
or UO_702 (O_702,N_10017,N_13629);
nand UO_703 (O_703,N_13781,N_12192);
nor UO_704 (O_704,N_11361,N_12599);
nor UO_705 (O_705,N_14969,N_11069);
and UO_706 (O_706,N_11544,N_13618);
and UO_707 (O_707,N_12097,N_13187);
or UO_708 (O_708,N_14494,N_13575);
xnor UO_709 (O_709,N_12523,N_10781);
and UO_710 (O_710,N_13225,N_11043);
or UO_711 (O_711,N_11231,N_14478);
or UO_712 (O_712,N_14435,N_14095);
and UO_713 (O_713,N_11073,N_13830);
xor UO_714 (O_714,N_12468,N_13013);
and UO_715 (O_715,N_13840,N_10650);
or UO_716 (O_716,N_14257,N_12381);
nor UO_717 (O_717,N_10009,N_12557);
nor UO_718 (O_718,N_14142,N_14499);
nor UO_719 (O_719,N_14161,N_14150);
nor UO_720 (O_720,N_12250,N_11254);
and UO_721 (O_721,N_12934,N_13503);
or UO_722 (O_722,N_13995,N_14088);
nor UO_723 (O_723,N_13885,N_10659);
nor UO_724 (O_724,N_11982,N_13889);
nand UO_725 (O_725,N_12546,N_13414);
or UO_726 (O_726,N_11998,N_12955);
nor UO_727 (O_727,N_12737,N_12687);
and UO_728 (O_728,N_10502,N_10292);
nand UO_729 (O_729,N_14662,N_14376);
or UO_730 (O_730,N_10004,N_13534);
and UO_731 (O_731,N_13630,N_11197);
and UO_732 (O_732,N_11102,N_14473);
nor UO_733 (O_733,N_14810,N_11926);
xnor UO_734 (O_734,N_13844,N_10642);
xor UO_735 (O_735,N_10570,N_14417);
or UO_736 (O_736,N_12489,N_11740);
nand UO_737 (O_737,N_11163,N_10492);
and UO_738 (O_738,N_11712,N_11356);
xnor UO_739 (O_739,N_13736,N_10614);
or UO_740 (O_740,N_11419,N_12337);
or UO_741 (O_741,N_10216,N_13878);
and UO_742 (O_742,N_14735,N_14543);
nand UO_743 (O_743,N_10610,N_14198);
nor UO_744 (O_744,N_10619,N_14622);
or UO_745 (O_745,N_14103,N_10977);
nor UO_746 (O_746,N_12705,N_14814);
nand UO_747 (O_747,N_10913,N_13129);
and UO_748 (O_748,N_10506,N_11257);
nand UO_749 (O_749,N_10547,N_12718);
nand UO_750 (O_750,N_11924,N_10037);
nor UO_751 (O_751,N_13223,N_12460);
xor UO_752 (O_752,N_11625,N_10522);
nand UO_753 (O_753,N_11293,N_11101);
nand UO_754 (O_754,N_14455,N_10223);
xor UO_755 (O_755,N_12028,N_12424);
nand UO_756 (O_756,N_13548,N_11879);
or UO_757 (O_757,N_14916,N_14426);
nand UO_758 (O_758,N_11718,N_13184);
nor UO_759 (O_759,N_12341,N_13111);
and UO_760 (O_760,N_14290,N_13122);
nand UO_761 (O_761,N_10595,N_12032);
nor UO_762 (O_762,N_13387,N_12815);
and UO_763 (O_763,N_14966,N_12079);
nand UO_764 (O_764,N_12238,N_14836);
nor UO_765 (O_765,N_10726,N_10293);
xnor UO_766 (O_766,N_12636,N_10961);
nor UO_767 (O_767,N_14004,N_11137);
and UO_768 (O_768,N_14372,N_10741);
nand UO_769 (O_769,N_13188,N_14684);
nand UO_770 (O_770,N_12092,N_14751);
nand UO_771 (O_771,N_13920,N_13569);
or UO_772 (O_772,N_12662,N_13721);
or UO_773 (O_773,N_11461,N_14758);
or UO_774 (O_774,N_11456,N_12499);
nand UO_775 (O_775,N_10582,N_10971);
nor UO_776 (O_776,N_10970,N_10722);
nand UO_777 (O_777,N_10164,N_12104);
nor UO_778 (O_778,N_14915,N_10116);
nor UO_779 (O_779,N_12879,N_12386);
and UO_780 (O_780,N_10196,N_10766);
and UO_781 (O_781,N_11824,N_10250);
and UO_782 (O_782,N_12549,N_12771);
xor UO_783 (O_783,N_13938,N_12234);
or UO_784 (O_784,N_13952,N_14354);
nand UO_785 (O_785,N_11518,N_10189);
xor UO_786 (O_786,N_14108,N_12428);
nand UO_787 (O_787,N_11613,N_10914);
nor UO_788 (O_788,N_10796,N_12201);
or UO_789 (O_789,N_13546,N_11693);
and UO_790 (O_790,N_11310,N_12050);
or UO_791 (O_791,N_11701,N_13739);
nor UO_792 (O_792,N_13719,N_14025);
nor UO_793 (O_793,N_12696,N_10715);
or UO_794 (O_794,N_10080,N_14990);
or UO_795 (O_795,N_12455,N_12782);
nand UO_796 (O_796,N_11604,N_14696);
nor UO_797 (O_797,N_10546,N_14522);
or UO_798 (O_798,N_11642,N_13916);
nor UO_799 (O_799,N_14702,N_11425);
or UO_800 (O_800,N_10645,N_10752);
nand UO_801 (O_801,N_14740,N_13928);
and UO_802 (O_802,N_11218,N_12798);
nand UO_803 (O_803,N_10394,N_10112);
xnor UO_804 (O_804,N_13318,N_14582);
or UO_805 (O_805,N_12814,N_14766);
nand UO_806 (O_806,N_13322,N_14646);
or UO_807 (O_807,N_13077,N_10088);
and UO_808 (O_808,N_11623,N_12512);
or UO_809 (O_809,N_10486,N_13835);
nor UO_810 (O_810,N_13730,N_12804);
or UO_811 (O_811,N_14796,N_11511);
and UO_812 (O_812,N_12490,N_10377);
or UO_813 (O_813,N_12404,N_13564);
nor UO_814 (O_814,N_10603,N_11574);
and UO_815 (O_815,N_13976,N_13634);
xor UO_816 (O_816,N_14986,N_13589);
or UO_817 (O_817,N_13810,N_12994);
nor UO_818 (O_818,N_10873,N_14123);
nand UO_819 (O_819,N_12578,N_11277);
nor UO_820 (O_820,N_12385,N_13869);
and UO_821 (O_821,N_12950,N_12041);
and UO_822 (O_822,N_11089,N_11048);
nand UO_823 (O_823,N_11709,N_12973);
nor UO_824 (O_824,N_10400,N_11991);
and UO_825 (O_825,N_12831,N_12044);
nand UO_826 (O_826,N_12253,N_14357);
xor UO_827 (O_827,N_13030,N_12363);
nand UO_828 (O_828,N_11274,N_11972);
nand UO_829 (O_829,N_13797,N_12450);
nand UO_830 (O_830,N_12078,N_13246);
and UO_831 (O_831,N_13945,N_11134);
and UO_832 (O_832,N_11630,N_10945);
nand UO_833 (O_833,N_12054,N_11193);
nand UO_834 (O_834,N_12459,N_11333);
or UO_835 (O_835,N_10598,N_10078);
nor UO_836 (O_836,N_11259,N_11593);
nand UO_837 (O_837,N_14726,N_14467);
xor UO_838 (O_838,N_10863,N_12098);
and UO_839 (O_839,N_11568,N_14226);
nand UO_840 (O_840,N_13704,N_11961);
nand UO_841 (O_841,N_12494,N_13214);
nor UO_842 (O_842,N_12869,N_14514);
and UO_843 (O_843,N_12382,N_14614);
nor UO_844 (O_844,N_14284,N_12507);
nor UO_845 (O_845,N_12495,N_14482);
nand UO_846 (O_846,N_11345,N_12660);
nor UO_847 (O_847,N_12975,N_14313);
nand UO_848 (O_848,N_14408,N_12572);
or UO_849 (O_849,N_10197,N_10447);
and UO_850 (O_850,N_13396,N_12120);
nand UO_851 (O_851,N_11928,N_12658);
and UO_852 (O_852,N_10714,N_13354);
and UO_853 (O_853,N_14393,N_12496);
or UO_854 (O_854,N_12426,N_13649);
and UO_855 (O_855,N_13325,N_14287);
nand UO_856 (O_856,N_12728,N_14071);
xnor UO_857 (O_857,N_10612,N_13237);
xor UO_858 (O_858,N_10600,N_11330);
or UO_859 (O_859,N_14626,N_13710);
or UO_860 (O_860,N_14856,N_11177);
or UO_861 (O_861,N_12340,N_13475);
or UO_862 (O_862,N_10405,N_11940);
xor UO_863 (O_863,N_12525,N_14064);
nand UO_864 (O_864,N_12465,N_13570);
xnor UO_865 (O_865,N_14850,N_14476);
xnor UO_866 (O_866,N_11380,N_13406);
and UO_867 (O_867,N_10569,N_10321);
and UO_868 (O_868,N_12302,N_11408);
xor UO_869 (O_869,N_13588,N_10033);
or UO_870 (O_870,N_12593,N_13865);
and UO_871 (O_871,N_12252,N_10912);
or UO_872 (O_872,N_11573,N_10786);
nor UO_873 (O_873,N_10061,N_12150);
nand UO_874 (O_874,N_12958,N_13742);
nor UO_875 (O_875,N_14087,N_11878);
nor UO_876 (O_876,N_14997,N_11322);
nand UO_877 (O_877,N_13307,N_14039);
nand UO_878 (O_878,N_11455,N_10980);
or UO_879 (O_879,N_10372,N_11287);
xor UO_880 (O_880,N_11852,N_14724);
and UO_881 (O_881,N_10981,N_13757);
nor UO_882 (O_882,N_11316,N_11338);
and UO_883 (O_883,N_12143,N_14532);
or UO_884 (O_884,N_14490,N_14991);
nor UO_885 (O_885,N_11682,N_14349);
nor UO_886 (O_886,N_11011,N_12029);
or UO_887 (O_887,N_12894,N_14059);
nand UO_888 (O_888,N_12012,N_12689);
nand UO_889 (O_889,N_13190,N_14385);
nand UO_890 (O_890,N_13003,N_11324);
and UO_891 (O_891,N_13156,N_13783);
and UO_892 (O_892,N_11689,N_14152);
nand UO_893 (O_893,N_13641,N_12735);
nand UO_894 (O_894,N_10535,N_11190);
and UO_895 (O_895,N_10640,N_10345);
or UO_896 (O_896,N_13460,N_10780);
nand UO_897 (O_897,N_12371,N_12023);
nand UO_898 (O_898,N_13627,N_14261);
xor UO_899 (O_899,N_10860,N_13254);
xor UO_900 (O_900,N_11106,N_10159);
nor UO_901 (O_901,N_10025,N_11512);
nor UO_902 (O_902,N_10676,N_12294);
nor UO_903 (O_903,N_13150,N_14719);
and UO_904 (O_904,N_11588,N_14504);
and UO_905 (O_905,N_10618,N_11395);
or UO_906 (O_906,N_13166,N_10107);
nor UO_907 (O_907,N_11149,N_12710);
nor UO_908 (O_908,N_10027,N_10396);
xnor UO_909 (O_909,N_14047,N_10505);
nor UO_910 (O_910,N_12300,N_11127);
xor UO_911 (O_911,N_10274,N_11918);
or UO_912 (O_912,N_14042,N_12126);
and UO_913 (O_913,N_13511,N_11238);
and UO_914 (O_914,N_11487,N_13960);
nand UO_915 (O_915,N_12927,N_14937);
and UO_916 (O_916,N_13899,N_13944);
and UO_917 (O_917,N_14229,N_10734);
nor UO_918 (O_918,N_11955,N_14949);
or UO_919 (O_919,N_13066,N_10094);
xor UO_920 (O_920,N_13094,N_10229);
and UO_921 (O_921,N_14547,N_14069);
and UO_922 (O_922,N_10109,N_12816);
or UO_923 (O_923,N_14785,N_12194);
nor UO_924 (O_924,N_13060,N_11241);
or UO_925 (O_925,N_12556,N_10125);
or UO_926 (O_926,N_14468,N_13068);
or UO_927 (O_927,N_14272,N_11763);
or UO_928 (O_928,N_11945,N_13592);
xor UO_929 (O_929,N_13124,N_10792);
nand UO_930 (O_930,N_11340,N_14753);
and UO_931 (O_931,N_11546,N_14118);
or UO_932 (O_932,N_12919,N_14110);
nand UO_933 (O_933,N_13632,N_14672);
nor UO_934 (O_934,N_10323,N_14993);
or UO_935 (O_935,N_14693,N_13021);
and UO_936 (O_936,N_10698,N_13578);
or UO_937 (O_937,N_11336,N_12498);
xnor UO_938 (O_938,N_12265,N_12986);
xor UO_939 (O_939,N_13539,N_14644);
or UO_940 (O_940,N_11929,N_13518);
nand UO_941 (O_941,N_14849,N_14946);
and UO_942 (O_942,N_10680,N_13790);
xnor UO_943 (O_943,N_14629,N_10815);
and UO_944 (O_944,N_10576,N_14608);
nor UO_945 (O_945,N_11145,N_11627);
nand UO_946 (O_946,N_11413,N_11931);
nor UO_947 (O_947,N_14839,N_13650);
nand UO_948 (O_948,N_11173,N_10449);
or UO_949 (O_949,N_13801,N_10264);
nor UO_950 (O_950,N_14663,N_13987);
nand UO_951 (O_951,N_12506,N_13873);
nor UO_952 (O_952,N_10294,N_12227);
xnor UO_953 (O_953,N_10539,N_10188);
nor UO_954 (O_954,N_11726,N_10050);
and UO_955 (O_955,N_13464,N_10788);
nor UO_956 (O_956,N_14173,N_11406);
and UO_957 (O_957,N_11084,N_10872);
nand UO_958 (O_958,N_14068,N_13762);
and UO_959 (O_959,N_12235,N_10974);
nor UO_960 (O_960,N_12885,N_12241);
nor UO_961 (O_961,N_14900,N_13792);
nor UO_962 (O_962,N_13764,N_10180);
or UO_963 (O_963,N_14191,N_14185);
or UO_964 (O_964,N_12430,N_14362);
nor UO_965 (O_965,N_13766,N_13752);
or UO_966 (O_966,N_11024,N_10586);
xnor UO_967 (O_967,N_14105,N_11366);
nand UO_968 (O_968,N_14812,N_10520);
xor UO_969 (O_969,N_13607,N_10946);
or UO_970 (O_970,N_11665,N_11970);
and UO_971 (O_971,N_14465,N_10049);
nand UO_972 (O_972,N_13353,N_11447);
or UO_973 (O_973,N_10187,N_10260);
or UO_974 (O_974,N_12020,N_11010);
nor UO_975 (O_975,N_13351,N_13697);
and UO_976 (O_976,N_14630,N_14611);
nand UO_977 (O_977,N_14824,N_14235);
xnor UO_978 (O_978,N_12292,N_11738);
nand UO_979 (O_979,N_11172,N_14477);
nor UO_980 (O_980,N_11354,N_10631);
xor UO_981 (O_981,N_11401,N_14121);
and UO_982 (O_982,N_13451,N_11248);
nand UO_983 (O_983,N_11329,N_11475);
xor UO_984 (O_984,N_14799,N_13191);
nor UO_985 (O_985,N_10340,N_10551);
nand UO_986 (O_986,N_12932,N_11473);
or UO_987 (O_987,N_11698,N_14895);
and UO_988 (O_988,N_11359,N_13202);
nor UO_989 (O_989,N_12027,N_11070);
or UO_990 (O_990,N_14940,N_11243);
nand UO_991 (O_991,N_11253,N_10324);
or UO_992 (O_992,N_11917,N_10203);
nor UO_993 (O_993,N_10701,N_10382);
nand UO_994 (O_994,N_13020,N_13501);
nor UO_995 (O_995,N_14742,N_10657);
and UO_996 (O_996,N_12003,N_14111);
and UO_997 (O_997,N_11126,N_12347);
nor UO_998 (O_998,N_11700,N_10311);
and UO_999 (O_999,N_12339,N_13892);
or UO_1000 (O_1000,N_13695,N_14704);
and UO_1001 (O_1001,N_11901,N_14728);
or UO_1002 (O_1002,N_11278,N_12072);
and UO_1003 (O_1003,N_14911,N_13767);
nand UO_1004 (O_1004,N_12725,N_14415);
or UO_1005 (O_1005,N_10529,N_12066);
nand UO_1006 (O_1006,N_13487,N_10262);
or UO_1007 (O_1007,N_13441,N_13211);
nor UO_1008 (O_1008,N_14422,N_14466);
or UO_1009 (O_1009,N_10297,N_12614);
or UO_1010 (O_1010,N_10157,N_10805);
nand UO_1011 (O_1011,N_11436,N_11967);
nand UO_1012 (O_1012,N_10861,N_12333);
nand UO_1013 (O_1013,N_13252,N_14193);
or UO_1014 (O_1014,N_14061,N_12011);
and UO_1015 (O_1015,N_12933,N_11794);
or UO_1016 (O_1016,N_11848,N_11082);
xor UO_1017 (O_1017,N_11553,N_11454);
nor UO_1018 (O_1018,N_13317,N_12677);
nand UO_1019 (O_1019,N_10181,N_12837);
and UO_1020 (O_1020,N_11821,N_14618);
nor UO_1021 (O_1021,N_11099,N_11268);
xor UO_1022 (O_1022,N_13130,N_11510);
and UO_1023 (O_1023,N_10014,N_14218);
nand UO_1024 (O_1024,N_11538,N_13106);
xor UO_1025 (O_1025,N_10198,N_10089);
or UO_1026 (O_1026,N_11517,N_10387);
nor UO_1027 (O_1027,N_10959,N_11995);
nor UO_1028 (O_1028,N_10567,N_11168);
and UO_1029 (O_1029,N_13549,N_11795);
or UO_1030 (O_1030,N_12774,N_11949);
nand UO_1031 (O_1031,N_11645,N_11042);
or UO_1032 (O_1032,N_13398,N_12889);
nand UO_1033 (O_1033,N_12632,N_13091);
and UO_1034 (O_1034,N_10927,N_12564);
or UO_1035 (O_1035,N_14228,N_13858);
xnor UO_1036 (O_1036,N_12793,N_14590);
or UO_1037 (O_1037,N_12645,N_13741);
and UO_1038 (O_1038,N_10587,N_10210);
and UO_1039 (O_1039,N_13833,N_14784);
and UO_1040 (O_1040,N_14950,N_13334);
and UO_1041 (O_1041,N_12138,N_12882);
xnor UO_1042 (O_1042,N_12951,N_10579);
or UO_1043 (O_1043,N_10128,N_13854);
nor UO_1044 (O_1044,N_13485,N_13194);
nand UO_1045 (O_1045,N_10474,N_10355);
and UO_1046 (O_1046,N_11589,N_12923);
or UO_1047 (O_1047,N_10076,N_14677);
xor UO_1048 (O_1048,N_12179,N_14117);
or UO_1049 (O_1049,N_13644,N_13698);
and UO_1050 (O_1050,N_12794,N_14028);
or UO_1051 (O_1051,N_14685,N_14884);
and UO_1052 (O_1052,N_13610,N_10048);
and UO_1053 (O_1053,N_10544,N_12836);
or UO_1054 (O_1054,N_11865,N_11734);
nor UO_1055 (O_1055,N_12288,N_10225);
and UO_1056 (O_1056,N_13011,N_13749);
nor UO_1057 (O_1057,N_12358,N_10020);
and UO_1058 (O_1058,N_10925,N_12007);
nand UO_1059 (O_1059,N_12803,N_12108);
or UO_1060 (O_1060,N_10397,N_10572);
or UO_1061 (O_1061,N_13365,N_10102);
nand UO_1062 (O_1062,N_11847,N_12324);
nor UO_1063 (O_1063,N_12722,N_12445);
nor UO_1064 (O_1064,N_14697,N_14567);
nand UO_1065 (O_1065,N_11055,N_12384);
or UO_1066 (O_1066,N_13827,N_10802);
nand UO_1067 (O_1067,N_12081,N_14332);
nand UO_1068 (O_1068,N_13008,N_11695);
and UO_1069 (O_1069,N_13051,N_12619);
and UO_1070 (O_1070,N_12591,N_12149);
nor UO_1071 (O_1071,N_14119,N_14052);
nor UO_1072 (O_1072,N_11433,N_13410);
nand UO_1073 (O_1073,N_11468,N_13209);
nor UO_1074 (O_1074,N_13050,N_12396);
and UO_1075 (O_1075,N_10866,N_12753);
nor UO_1076 (O_1076,N_11056,N_12824);
xor UO_1077 (O_1077,N_12412,N_14436);
nor UO_1078 (O_1078,N_14692,N_11227);
nor UO_1079 (O_1079,N_14538,N_10616);
or UO_1080 (O_1080,N_10270,N_13472);
or UO_1081 (O_1081,N_14262,N_12167);
and UO_1082 (O_1082,N_13107,N_13992);
nor UO_1083 (O_1083,N_10175,N_12096);
or UO_1084 (O_1084,N_12226,N_10880);
nor UO_1085 (O_1085,N_12761,N_14848);
or UO_1086 (O_1086,N_14109,N_11459);
nor UO_1087 (O_1087,N_13284,N_11594);
nor UO_1088 (O_1088,N_11153,N_11964);
nand UO_1089 (O_1089,N_12493,N_10393);
or UO_1090 (O_1090,N_14461,N_11432);
nand UO_1091 (O_1091,N_12418,N_10035);
and UO_1092 (O_1092,N_11805,N_14432);
or UO_1093 (O_1093,N_11942,N_10373);
and UO_1094 (O_1094,N_13845,N_13340);
nand UO_1095 (O_1095,N_11014,N_13090);
or UO_1096 (O_1096,N_11713,N_14032);
nand UO_1097 (O_1097,N_10534,N_13877);
or UO_1098 (O_1098,N_13613,N_13235);
nand UO_1099 (O_1099,N_13702,N_14438);
and UO_1100 (O_1100,N_12790,N_11209);
and UO_1101 (O_1101,N_11822,N_11367);
nor UO_1102 (O_1102,N_13560,N_14718);
and UO_1103 (O_1103,N_10152,N_14801);
nor UO_1104 (O_1104,N_11809,N_13059);
nor UO_1105 (O_1105,N_14749,N_14096);
nor UO_1106 (O_1106,N_14227,N_13279);
nand UO_1107 (O_1107,N_11263,N_11943);
nor UO_1108 (O_1108,N_10527,N_10732);
and UO_1109 (O_1109,N_12800,N_12937);
nand UO_1110 (O_1110,N_10824,N_12685);
nor UO_1111 (O_1111,N_10917,N_12152);
xnor UO_1112 (O_1112,N_11108,N_12351);
nand UO_1113 (O_1113,N_10563,N_13819);
xnor UO_1114 (O_1114,N_10200,N_11444);
or UO_1115 (O_1115,N_14474,N_13243);
or UO_1116 (O_1116,N_13245,N_10485);
nor UO_1117 (O_1117,N_14687,N_13486);
and UO_1118 (O_1118,N_13870,N_14525);
nand UO_1119 (O_1119,N_10455,N_14297);
or UO_1120 (O_1120,N_13189,N_13206);
nand UO_1121 (O_1121,N_11989,N_10886);
and UO_1122 (O_1122,N_13681,N_11756);
and UO_1123 (O_1123,N_14424,N_14005);
or UO_1124 (O_1124,N_12368,N_12603);
xor UO_1125 (O_1125,N_12378,N_14942);
xor UO_1126 (O_1126,N_12954,N_11230);
or UO_1127 (O_1127,N_14327,N_14170);
or UO_1128 (O_1128,N_10784,N_12325);
and UO_1129 (O_1129,N_11524,N_12702);
xnor UO_1130 (O_1130,N_14434,N_13508);
nor UO_1131 (O_1131,N_10454,N_14270);
or UO_1132 (O_1132,N_11834,N_11522);
or UO_1133 (O_1133,N_11661,N_12148);
or UO_1134 (O_1134,N_13196,N_12627);
nor UO_1135 (O_1135,N_10916,N_11150);
and UO_1136 (O_1136,N_13643,N_10193);
nand UO_1137 (O_1137,N_10988,N_11769);
nor UO_1138 (O_1138,N_10583,N_14399);
nand UO_1139 (O_1139,N_13637,N_14104);
or UO_1140 (O_1140,N_12214,N_11492);
and UO_1141 (O_1141,N_13085,N_14682);
and UO_1142 (O_1142,N_12765,N_11049);
or UO_1143 (O_1143,N_11464,N_12067);
xnor UO_1144 (O_1144,N_13784,N_12659);
nor UO_1145 (O_1145,N_14665,N_13138);
xor UO_1146 (O_1146,N_14516,N_12542);
nand UO_1147 (O_1147,N_11598,N_12483);
or UO_1148 (O_1148,N_11236,N_13301);
or UO_1149 (O_1149,N_10707,N_12622);
xnor UO_1150 (O_1150,N_14382,N_14867);
and UO_1151 (O_1151,N_10806,N_10848);
nor UO_1152 (O_1152,N_11536,N_12682);
nand UO_1153 (O_1153,N_13664,N_10858);
and UO_1154 (O_1154,N_12596,N_14612);
and UO_1155 (O_1155,N_14898,N_10841);
nor UO_1156 (O_1156,N_13429,N_10565);
or UO_1157 (O_1157,N_12999,N_14771);
nand UO_1158 (O_1158,N_12362,N_10634);
nand UO_1159 (O_1159,N_14423,N_12983);
or UO_1160 (O_1160,N_13849,N_14932);
nor UO_1161 (O_1161,N_13281,N_11362);
and UO_1162 (O_1162,N_10473,N_11502);
and UO_1163 (O_1163,N_10549,N_13327);
or UO_1164 (O_1164,N_11914,N_14561);
nand UO_1165 (O_1165,N_14586,N_11164);
nand UO_1166 (O_1166,N_12567,N_10730);
nand UO_1167 (O_1167,N_11767,N_11910);
nand UO_1168 (O_1168,N_13047,N_10137);
and UO_1169 (O_1169,N_11811,N_10826);
and UO_1170 (O_1170,N_10042,N_14698);
nor UO_1171 (O_1171,N_13079,N_12042);
and UO_1172 (O_1172,N_13062,N_14314);
nand UO_1173 (O_1173,N_11912,N_10117);
nor UO_1174 (O_1174,N_10742,N_13990);
nor UO_1175 (O_1175,N_14380,N_12454);
and UO_1176 (O_1176,N_11721,N_11697);
or UO_1177 (O_1177,N_11849,N_11394);
and UO_1178 (O_1178,N_11469,N_13614);
nor UO_1179 (O_1179,N_10095,N_10702);
nor UO_1180 (O_1180,N_10144,N_13851);
nand UO_1181 (O_1181,N_11828,N_11282);
xor UO_1182 (O_1182,N_11434,N_11923);
nand UO_1183 (O_1183,N_11560,N_11670);
nor UO_1184 (O_1184,N_12633,N_13939);
xnor UO_1185 (O_1185,N_10282,N_10379);
nand UO_1186 (O_1186,N_10517,N_10028);
nor UO_1187 (O_1187,N_11129,N_11580);
or UO_1188 (O_1188,N_14199,N_11827);
and UO_1189 (O_1189,N_14254,N_13428);
nand UO_1190 (O_1190,N_13326,N_11858);
nand UO_1191 (O_1191,N_14006,N_12306);
nor UO_1192 (O_1192,N_10853,N_12400);
and UO_1193 (O_1193,N_13895,N_10073);
nor UO_1194 (O_1194,N_11869,N_12890);
or UO_1195 (O_1195,N_11873,N_11727);
or UO_1196 (O_1196,N_11533,N_10019);
nand UO_1197 (O_1197,N_10772,N_14283);
xnor UO_1198 (O_1198,N_14165,N_14450);
nand UO_1199 (O_1199,N_10207,N_10838);
nor UO_1200 (O_1200,N_10728,N_14344);
nor UO_1201 (O_1201,N_12309,N_11207);
or UO_1202 (O_1202,N_12034,N_10515);
or UO_1203 (O_1203,N_13682,N_13375);
nor UO_1204 (O_1204,N_14136,N_12168);
and UO_1205 (O_1205,N_11063,N_13420);
nand UO_1206 (O_1206,N_14569,N_11906);
xor UO_1207 (O_1207,N_11963,N_13765);
xor UO_1208 (O_1208,N_12909,N_11686);
nand UO_1209 (O_1209,N_14587,N_11431);
or UO_1210 (O_1210,N_12049,N_12796);
nand UO_1211 (O_1211,N_14513,N_13500);
nand UO_1212 (O_1212,N_14570,N_11543);
nor UO_1213 (O_1213,N_11728,N_13176);
or UO_1214 (O_1214,N_11210,N_12715);
and UO_1215 (O_1215,N_13726,N_14732);
nor UO_1216 (O_1216,N_14789,N_13864);
and UO_1217 (O_1217,N_10843,N_12844);
nor UO_1218 (O_1218,N_11384,N_10038);
xor UO_1219 (O_1219,N_12822,N_14960);
and UO_1220 (O_1220,N_11066,N_11618);
and UO_1221 (O_1221,N_11638,N_12182);
nor UO_1222 (O_1222,N_10430,N_10754);
or UO_1223 (O_1223,N_13579,N_13102);
or UO_1224 (O_1224,N_11052,N_13982);
or UO_1225 (O_1225,N_13227,N_12307);
nor UO_1226 (O_1226,N_10883,N_14737);
and UO_1227 (O_1227,N_12213,N_11020);
and UO_1228 (O_1228,N_13989,N_11664);
nor UO_1229 (O_1229,N_10892,N_14050);
or UO_1230 (O_1230,N_10558,N_10620);
nand UO_1231 (O_1231,N_12807,N_13597);
and UO_1232 (O_1232,N_12526,N_11614);
nor UO_1233 (O_1233,N_14649,N_14409);
and UO_1234 (O_1234,N_13010,N_10758);
and UO_1235 (O_1235,N_13274,N_10591);
and UO_1236 (O_1236,N_14782,N_14040);
nor UO_1237 (O_1237,N_10613,N_10763);
or UO_1238 (O_1238,N_10939,N_12299);
and UO_1239 (O_1239,N_10194,N_14689);
nand UO_1240 (O_1240,N_14208,N_13161);
and UO_1241 (O_1241,N_13372,N_10115);
and UO_1242 (O_1242,N_14787,N_10799);
and UO_1243 (O_1243,N_12391,N_13121);
nand UO_1244 (O_1244,N_14720,N_10585);
or UO_1245 (O_1245,N_12819,N_11851);
or UO_1246 (O_1246,N_13946,N_12854);
nand UO_1247 (O_1247,N_11061,N_12643);
nand UO_1248 (O_1248,N_13234,N_12727);
or UO_1249 (O_1249,N_10574,N_14597);
and UO_1250 (O_1250,N_11477,N_14823);
or UO_1251 (O_1251,N_12904,N_13862);
nor UO_1252 (O_1252,N_14512,N_10278);
and UO_1253 (O_1253,N_14759,N_11358);
nand UO_1254 (O_1254,N_10635,N_14086);
nand UO_1255 (O_1255,N_12948,N_12887);
nand UO_1256 (O_1256,N_13557,N_14520);
nor UO_1257 (O_1257,N_12071,N_11930);
or UO_1258 (O_1258,N_14300,N_13386);
or UO_1259 (O_1259,N_10606,N_14920);
and UO_1260 (O_1260,N_14838,N_14673);
nor UO_1261 (O_1261,N_14779,N_12485);
or UO_1262 (O_1262,N_12768,N_12045);
or UO_1263 (O_1263,N_10704,N_13512);
and UO_1264 (O_1264,N_11788,N_14153);
and UO_1265 (O_1265,N_10985,N_12925);
nor UO_1266 (O_1266,N_11656,N_14410);
or UO_1267 (O_1267,N_14106,N_11747);
nand UO_1268 (O_1268,N_12641,N_12211);
nand UO_1269 (O_1269,N_11313,N_10627);
nand UO_1270 (O_1270,N_13993,N_11420);
nand UO_1271 (O_1271,N_14939,N_11038);
nand UO_1272 (O_1272,N_13165,N_13522);
nor UO_1273 (O_1273,N_13026,N_14397);
and UO_1274 (O_1274,N_13112,N_12863);
xor UO_1275 (O_1275,N_14954,N_11054);
and UO_1276 (O_1276,N_12492,N_10168);
and UO_1277 (O_1277,N_11671,N_13174);
nor UO_1278 (O_1278,N_11028,N_12369);
or UO_1279 (O_1279,N_14756,N_11445);
and UO_1280 (O_1280,N_13812,N_10850);
nand UO_1281 (O_1281,N_10421,N_14530);
nand UO_1282 (O_1282,N_13886,N_10365);
or UO_1283 (O_1283,N_12892,N_10015);
nand UO_1284 (O_1284,N_13498,N_14970);
or UO_1285 (O_1285,N_11579,N_14707);
nand UO_1286 (O_1286,N_13147,N_14175);
nand UO_1287 (O_1287,N_12366,N_12908);
or UO_1288 (O_1288,N_14778,N_14959);
and UO_1289 (O_1289,N_10063,N_13342);
and UO_1290 (O_1290,N_13022,N_12321);
xor UO_1291 (O_1291,N_11381,N_14122);
nor UO_1292 (O_1292,N_14457,N_14244);
nand UO_1293 (O_1293,N_11703,N_13890);
nor UO_1294 (O_1294,N_14842,N_10118);
or UO_1295 (O_1295,N_11467,N_12571);
and UO_1296 (O_1296,N_12528,N_14671);
xor UO_1297 (O_1297,N_12287,N_10964);
or UO_1298 (O_1298,N_12082,N_14515);
nor UO_1299 (O_1299,N_14804,N_12268);
or UO_1300 (O_1300,N_10462,N_10494);
or UO_1301 (O_1301,N_10273,N_14757);
nand UO_1302 (O_1302,N_11375,N_11040);
or UO_1303 (O_1303,N_11791,N_10156);
and UO_1304 (O_1304,N_11026,N_11761);
or UO_1305 (O_1305,N_11214,N_11279);
xnor UO_1306 (O_1306,N_13754,N_10407);
nand UO_1307 (O_1307,N_11959,N_10438);
or UO_1308 (O_1308,N_12491,N_14822);
nor UO_1309 (O_1309,N_10434,N_13785);
and UO_1310 (O_1310,N_11021,N_11495);
nor UO_1311 (O_1311,N_10953,N_10154);
and UO_1312 (O_1312,N_13582,N_10868);
or UO_1313 (O_1313,N_14560,N_10257);
xor UO_1314 (O_1314,N_10626,N_11076);
nand UO_1315 (O_1315,N_12295,N_11735);
nand UO_1316 (O_1316,N_11178,N_11622);
nand UO_1317 (O_1317,N_12095,N_10695);
nor UO_1318 (O_1318,N_12751,N_10423);
nor UO_1319 (O_1319,N_12501,N_11350);
nor UO_1320 (O_1320,N_11780,N_11999);
or UO_1321 (O_1321,N_10738,N_12789);
nand UO_1322 (O_1322,N_14524,N_14367);
nor UO_1323 (O_1323,N_10341,N_12941);
or UO_1324 (O_1324,N_14982,N_11764);
and UO_1325 (O_1325,N_10937,N_11798);
and UO_1326 (O_1326,N_11582,N_11587);
and UO_1327 (O_1327,N_11548,N_10255);
or UO_1328 (O_1328,N_13818,N_14154);
nand UO_1329 (O_1329,N_11352,N_13872);
nor UO_1330 (O_1330,N_14359,N_11965);
and UO_1331 (O_1331,N_10410,N_10123);
or UO_1332 (O_1332,N_11673,N_12859);
and UO_1333 (O_1333,N_10243,N_10247);
nor UO_1334 (O_1334,N_13192,N_12510);
nor UO_1335 (O_1335,N_11800,N_14853);
xnor UO_1336 (O_1336,N_11479,N_13255);
xnor UO_1337 (O_1337,N_10905,N_14926);
and UO_1338 (O_1338,N_12379,N_10867);
nand UO_1339 (O_1339,N_14265,N_12261);
and UO_1340 (O_1340,N_14360,N_10232);
nor UO_1341 (O_1341,N_14602,N_10951);
and UO_1342 (O_1342,N_14531,N_12960);
or UO_1343 (O_1343,N_14321,N_14576);
nor UO_1344 (O_1344,N_14201,N_10656);
nand UO_1345 (O_1345,N_12310,N_10746);
and UO_1346 (O_1346,N_14342,N_14738);
xnor UO_1347 (O_1347,N_14903,N_10132);
nand UO_1348 (O_1348,N_10006,N_10003);
or UO_1349 (O_1349,N_10510,N_13268);
nor UO_1350 (O_1350,N_13308,N_14765);
and UO_1351 (O_1351,N_11186,N_10870);
and UO_1352 (O_1352,N_12720,N_11124);
nor UO_1353 (O_1353,N_13884,N_10562);
or UO_1354 (O_1354,N_13238,N_11872);
or UO_1355 (O_1355,N_14500,N_13950);
nor UO_1356 (O_1356,N_10218,N_10008);
or UO_1357 (O_1357,N_11685,N_10056);
xnor UO_1358 (O_1358,N_10468,N_14965);
nand UO_1359 (O_1359,N_13917,N_10333);
nand UO_1360 (O_1360,N_12997,N_12242);
nor UO_1361 (O_1361,N_12672,N_10857);
nor UO_1362 (O_1362,N_13180,N_10795);
nor UO_1363 (O_1363,N_11584,N_13244);
nand UO_1364 (O_1364,N_11165,N_14034);
or UO_1365 (O_1365,N_11355,N_10184);
nand UO_1366 (O_1366,N_10545,N_14599);
nand UO_1367 (O_1367,N_12640,N_11952);
or UO_1368 (O_1368,N_12219,N_14631);
xor UO_1369 (O_1369,N_14609,N_13732);
nor UO_1370 (O_1370,N_13052,N_12913);
nand UO_1371 (O_1371,N_11016,N_13358);
xnor UO_1372 (O_1372,N_13443,N_13881);
nand UO_1373 (O_1373,N_12920,N_11653);
nand UO_1374 (O_1374,N_11430,N_11863);
nand UO_1375 (O_1375,N_13098,N_12880);
and UO_1376 (O_1376,N_13737,N_10646);
nor UO_1377 (O_1377,N_11629,N_11590);
xor UO_1378 (O_1378,N_10245,N_10991);
nand UO_1379 (O_1379,N_10785,N_12929);
nor UO_1380 (O_1380,N_12561,N_13648);
nor UO_1381 (O_1381,N_11657,N_10261);
or UO_1382 (O_1382,N_14956,N_14843);
or UO_1383 (O_1383,N_10664,N_12534);
nor UO_1384 (O_1384,N_11378,N_13753);
and UO_1385 (O_1385,N_11269,N_10789);
xnor UO_1386 (O_1386,N_13437,N_12117);
nand UO_1387 (O_1387,N_14120,N_10185);
and UO_1388 (O_1388,N_14416,N_13045);
or UO_1389 (O_1389,N_13789,N_13970);
and UO_1390 (O_1390,N_12163,N_14437);
nand UO_1391 (O_1391,N_13277,N_13521);
or UO_1392 (O_1392,N_14020,N_12776);
or UO_1393 (O_1393,N_14023,N_11893);
or UO_1394 (O_1394,N_13363,N_13718);
or UO_1395 (O_1395,N_11978,N_12903);
and UO_1396 (O_1396,N_14716,N_11932);
nand UO_1397 (O_1397,N_14370,N_11146);
or UO_1398 (O_1398,N_10367,N_14484);
and UO_1399 (O_1399,N_10484,N_14660);
or UO_1400 (O_1400,N_13626,N_13215);
and UO_1401 (O_1401,N_14694,N_14163);
xor UO_1402 (O_1402,N_10602,N_13335);
and UO_1403 (O_1403,N_11104,N_14174);
nand UO_1404 (O_1404,N_14887,N_11962);
nand UO_1405 (O_1405,N_13292,N_12409);
or UO_1406 (O_1406,N_13333,N_14014);
nor UO_1407 (O_1407,N_10731,N_14885);
and UO_1408 (O_1408,N_10887,N_10064);
nand UO_1409 (O_1409,N_10158,N_13360);
nor UO_1410 (O_1410,N_10276,N_14768);
nand UO_1411 (O_1411,N_12888,N_12905);
nand UO_1412 (O_1412,N_10954,N_14864);
or UO_1413 (O_1413,N_11779,N_13787);
xor UO_1414 (O_1414,N_10705,N_11711);
or UO_1415 (O_1415,N_10969,N_11213);
nor UO_1416 (O_1416,N_13065,N_14398);
nand UO_1417 (O_1417,N_12719,N_12207);
or UO_1418 (O_1418,N_10380,N_10524);
nor UO_1419 (O_1419,N_12278,N_10269);
and UO_1420 (O_1420,N_12410,N_13181);
nand UO_1421 (O_1421,N_12502,N_10212);
and UO_1422 (O_1422,N_13482,N_12503);
nor UO_1423 (O_1423,N_12668,N_13315);
xor UO_1424 (O_1424,N_14977,N_13369);
or UO_1425 (O_1425,N_12519,N_12849);
and UO_1426 (O_1426,N_13491,N_11915);
and UO_1427 (O_1427,N_11699,N_11182);
and UO_1428 (O_1428,N_14414,N_12175);
or UO_1429 (O_1429,N_13113,N_11249);
nand UO_1430 (O_1430,N_12442,N_13350);
and UO_1431 (O_1431,N_11280,N_10465);
nor UO_1432 (O_1432,N_11988,N_10469);
nand UO_1433 (O_1433,N_12576,N_10130);
nand UO_1434 (O_1434,N_12102,N_13311);
nor UO_1435 (O_1435,N_10855,N_11443);
nand UO_1436 (O_1436,N_10052,N_10590);
nor UO_1437 (O_1437,N_13037,N_10211);
or UO_1438 (O_1438,N_11839,N_11862);
nand UO_1439 (O_1439,N_13773,N_10173);
and UO_1440 (O_1440,N_13110,N_10740);
nand UO_1441 (O_1441,N_13584,N_13376);
or UO_1442 (O_1442,N_13672,N_13442);
and UO_1443 (O_1443,N_10817,N_12541);
and UO_1444 (O_1444,N_10167,N_12393);
and UO_1445 (O_1445,N_10926,N_13499);
nor UO_1446 (O_1446,N_10555,N_12258);
nand UO_1447 (O_1447,N_12511,N_14892);
nor UO_1448 (O_1448,N_14691,N_12812);
or UO_1449 (O_1449,N_13658,N_13828);
nand UO_1450 (O_1450,N_10215,N_13831);
nor UO_1451 (O_1451,N_13390,N_11789);
nand UO_1452 (O_1452,N_10989,N_12609);
and UO_1453 (O_1453,N_14606,N_13296);
or UO_1454 (O_1454,N_11875,N_12657);
xnor UO_1455 (O_1455,N_14301,N_12474);
nor UO_1456 (O_1456,N_12354,N_10778);
nor UO_1457 (O_1457,N_10428,N_12172);
and UO_1458 (O_1458,N_12334,N_13416);
and UO_1459 (O_1459,N_13918,N_12886);
nor UO_1460 (O_1460,N_11508,N_11181);
nand UO_1461 (O_1461,N_10775,N_12303);
and UO_1462 (O_1462,N_13669,N_12550);
xnor UO_1463 (O_1463,N_14239,N_11790);
or UO_1464 (O_1464,N_14491,N_11745);
and UO_1465 (O_1465,N_13898,N_11486);
nor UO_1466 (O_1466,N_14875,N_11641);
nand UO_1467 (O_1467,N_11953,N_10596);
and UO_1468 (O_1468,N_12577,N_13339);
or UO_1469 (O_1469,N_13053,N_11319);
nor UO_1470 (O_1470,N_14923,N_14412);
nand UO_1471 (O_1471,N_10729,N_12441);
nor UO_1472 (O_1472,N_11392,N_13659);
nand UO_1473 (O_1473,N_11387,N_14846);
and UO_1474 (O_1474,N_14462,N_10755);
or UO_1475 (O_1475,N_12729,N_13558);
nand UO_1476 (O_1476,N_12055,N_11130);
nor UO_1477 (O_1477,N_12928,N_11422);
or UO_1478 (O_1478,N_12039,N_12655);
and UO_1479 (O_1479,N_11710,N_11318);
and UO_1480 (O_1480,N_14311,N_12615);
nor UO_1481 (O_1481,N_10332,N_10617);
nor UO_1482 (O_1482,N_10920,N_11977);
xor UO_1483 (O_1483,N_12345,N_13299);
and UO_1484 (O_1484,N_12580,N_13295);
or UO_1485 (O_1485,N_12959,N_10328);
and UO_1486 (O_1486,N_10768,N_10907);
nand UO_1487 (O_1487,N_11631,N_12516);
nand UO_1488 (O_1488,N_11112,N_11397);
xnor UO_1489 (O_1489,N_10419,N_11398);
nor UO_1490 (O_1490,N_12487,N_10690);
nor UO_1491 (O_1491,N_12714,N_12154);
nor UO_1492 (O_1492,N_12106,N_11442);
and UO_1493 (O_1493,N_13389,N_12558);
nor UO_1494 (O_1494,N_10075,N_14642);
nand UO_1495 (O_1495,N_11890,N_11596);
nand UO_1496 (O_1496,N_12974,N_12562);
or UO_1497 (O_1497,N_11840,N_13893);
nor UO_1498 (O_1498,N_10713,N_10629);
or UO_1499 (O_1499,N_10950,N_13359);
or UO_1500 (O_1500,N_11937,N_10389);
or UO_1501 (O_1501,N_13465,N_11448);
and UO_1502 (O_1502,N_13210,N_14820);
nor UO_1503 (O_1503,N_13405,N_14803);
or UO_1504 (O_1504,N_11224,N_10177);
nand UO_1505 (O_1505,N_14541,N_14274);
xnor UO_1506 (O_1506,N_10149,N_14021);
or UO_1507 (O_1507,N_10536,N_10960);
nand UO_1508 (O_1508,N_14636,N_13457);
or UO_1509 (O_1509,N_14363,N_14137);
and UO_1510 (O_1510,N_10670,N_10541);
nor UO_1511 (O_1511,N_12217,N_13384);
nor UO_1512 (O_1512,N_11816,N_12711);
xnor UO_1513 (O_1513,N_12359,N_11390);
nand UO_1514 (O_1514,N_14003,N_10067);
and UO_1515 (O_1515,N_13266,N_12010);
nand UO_1516 (O_1516,N_11306,N_10832);
nand UO_1517 (O_1517,N_13368,N_13912);
nand UO_1518 (O_1518,N_11679,N_10133);
xnor UO_1519 (O_1519,N_10609,N_13115);
and UO_1520 (O_1520,N_13654,N_11549);
nand UO_1521 (O_1521,N_10398,N_14146);
nor UO_1522 (O_1522,N_11271,N_10471);
nand UO_1523 (O_1523,N_10652,N_13049);
or UO_1524 (O_1524,N_14307,N_12639);
nand UO_1525 (O_1525,N_10480,N_14835);
nand UO_1526 (O_1526,N_13963,N_12646);
nor UO_1527 (O_1527,N_13250,N_14951);
nand UO_1528 (O_1528,N_12992,N_13042);
nand UO_1529 (O_1529,N_13786,N_10807);
or UO_1530 (O_1530,N_12539,N_14471);
or UO_1531 (O_1531,N_11871,N_13417);
xor UO_1532 (O_1532,N_10139,N_11017);
and UO_1533 (O_1533,N_13652,N_14420);
or UO_1534 (O_1534,N_14961,N_10678);
and UO_1535 (O_1535,N_13400,N_10242);
xnor UO_1536 (O_1536,N_13269,N_11039);
nand UO_1537 (O_1537,N_11265,N_10688);
and UO_1538 (O_1538,N_11986,N_11303);
or UO_1539 (O_1539,N_12653,N_14973);
nor UO_1540 (O_1540,N_10561,N_11537);
or UO_1541 (O_1541,N_13715,N_11023);
or UO_1542 (O_1542,N_12308,N_14225);
or UO_1543 (O_1543,N_11925,N_12421);
or UO_1544 (O_1544,N_14326,N_11895);
nand UO_1545 (O_1545,N_11341,N_12691);
nor UO_1546 (O_1546,N_13285,N_12679);
xor UO_1547 (O_1547,N_14139,N_10043);
or UO_1548 (O_1548,N_14511,N_12741);
nor UO_1549 (O_1549,N_11325,N_12529);
and UO_1550 (O_1550,N_12649,N_12103);
and UO_1551 (O_1551,N_12989,N_13504);
nand UO_1552 (O_1552,N_13622,N_11820);
and UO_1553 (O_1553,N_13240,N_11648);
and UO_1554 (O_1554,N_11958,N_14180);
or UO_1555 (O_1555,N_12360,N_13239);
or UO_1556 (O_1556,N_12107,N_13073);
and UO_1557 (O_1557,N_11463,N_14379);
nand UO_1558 (O_1558,N_11610,N_14268);
nor UO_1559 (O_1559,N_13969,N_13510);
nand UO_1560 (O_1560,N_13619,N_14081);
or UO_1561 (O_1561,N_12508,N_14066);
and UO_1562 (O_1562,N_13253,N_13208);
and UO_1563 (O_1563,N_10251,N_10079);
xor UO_1564 (O_1564,N_13220,N_12795);
and UO_1565 (O_1565,N_13314,N_13323);
nor UO_1566 (O_1566,N_12280,N_10231);
and UO_1567 (O_1567,N_14070,N_12444);
nand UO_1568 (O_1568,N_13117,N_14248);
or UO_1569 (O_1569,N_12697,N_11814);
nor UO_1570 (O_1570,N_10329,N_10411);
nand UO_1571 (O_1571,N_13955,N_14130);
xor UO_1572 (O_1572,N_12413,N_10874);
and UO_1573 (O_1573,N_13668,N_12051);
nor UO_1574 (O_1574,N_11714,N_10919);
nor UO_1575 (O_1575,N_10904,N_11484);
xor UO_1576 (O_1576,N_14237,N_10265);
and UO_1577 (O_1577,N_13799,N_14746);
nand UO_1578 (O_1578,N_14469,N_10443);
or UO_1579 (O_1579,N_13447,N_12706);
and UO_1580 (O_1580,N_10644,N_13230);
or UO_1581 (O_1581,N_10891,N_13222);
or UO_1582 (O_1582,N_12312,N_13572);
and UO_1583 (O_1583,N_11750,N_13655);
or UO_1584 (O_1584,N_10651,N_10638);
or UO_1585 (O_1585,N_13975,N_13116);
nor UO_1586 (O_1586,N_13713,N_10351);
and UO_1587 (O_1587,N_11332,N_14717);
or UO_1588 (O_1588,N_10448,N_12686);
or UO_1589 (O_1589,N_11514,N_11666);
nor UO_1590 (O_1590,N_12964,N_14883);
nand UO_1591 (O_1591,N_12053,N_14497);
nand UO_1592 (O_1592,N_14635,N_12988);
or UO_1593 (O_1593,N_13772,N_12019);
or UO_1594 (O_1594,N_14921,N_10783);
nor UO_1595 (O_1595,N_13164,N_13921);
and UO_1596 (O_1596,N_12834,N_13653);
nand UO_1597 (O_1597,N_12766,N_13604);
nand UO_1598 (O_1598,N_13605,N_14328);
nand UO_1599 (O_1599,N_14183,N_13565);
and UO_1600 (O_1600,N_12296,N_12274);
and UO_1601 (O_1601,N_12446,N_14924);
and UO_1602 (O_1602,N_11143,N_11521);
xor UO_1603 (O_1603,N_14862,N_14323);
nand UO_1604 (O_1604,N_10787,N_11675);
or UO_1605 (O_1605,N_14177,N_14441);
and UO_1606 (O_1606,N_10601,N_10358);
or UO_1607 (O_1607,N_13576,N_11976);
nand UO_1608 (O_1608,N_12225,N_14396);
nand UO_1609 (O_1609,N_10685,N_11221);
and UO_1610 (O_1610,N_14427,N_14181);
and UO_1611 (O_1611,N_13379,N_12006);
nor UO_1612 (O_1612,N_11717,N_14761);
nand UO_1613 (O_1613,N_13125,N_10083);
or UO_1614 (O_1614,N_10068,N_10552);
xnor UO_1615 (O_1615,N_11569,N_10416);
nand UO_1616 (O_1616,N_12757,N_12912);
and UO_1617 (O_1617,N_14995,N_11819);
nor UO_1618 (O_1618,N_13850,N_12336);
nand UO_1619 (O_1619,N_11184,N_14668);
nor UO_1620 (O_1620,N_10623,N_11753);
or UO_1621 (O_1621,N_10592,N_11876);
nor UO_1622 (O_1622,N_13687,N_10862);
nor UO_1623 (O_1623,N_13374,N_10070);
or UO_1624 (O_1624,N_12036,N_12395);
nand UO_1625 (O_1625,N_12416,N_12471);
and UO_1626 (O_1626,N_12156,N_11438);
xor UO_1627 (O_1627,N_14978,N_10743);
and UO_1628 (O_1628,N_11496,N_11934);
nor UO_1629 (O_1629,N_10878,N_13033);
xor UO_1630 (O_1630,N_13729,N_13696);
nand UO_1631 (O_1631,N_12001,N_11081);
nand UO_1632 (O_1632,N_10334,N_14166);
or UO_1633 (O_1633,N_14974,N_14700);
and UO_1634 (O_1634,N_13983,N_14299);
nor UO_1635 (O_1635,N_10370,N_10446);
or UO_1636 (O_1636,N_10767,N_10888);
and UO_1637 (O_1637,N_13415,N_13985);
or UO_1638 (O_1638,N_11019,N_11196);
nand UO_1639 (O_1639,N_12618,N_11771);
and UO_1640 (O_1640,N_13545,N_11051);
xor UO_1641 (O_1641,N_11093,N_13788);
nand UO_1642 (O_1642,N_14594,N_11724);
nor UO_1643 (O_1643,N_13927,N_13887);
and UO_1644 (O_1644,N_10060,N_11365);
nor UO_1645 (O_1645,N_13967,N_13381);
xor UO_1646 (O_1646,N_10818,N_14401);
or UO_1647 (O_1647,N_11311,N_13038);
nor UO_1648 (O_1648,N_11504,N_11344);
nor UO_1649 (O_1649,N_12709,N_13774);
or UO_1650 (O_1650,N_11437,N_11662);
and UO_1651 (O_1651,N_14870,N_12698);
nand UO_1652 (O_1652,N_12093,N_11122);
nor UO_1653 (O_1653,N_10865,N_10289);
or UO_1654 (O_1654,N_13450,N_13273);
nand UO_1655 (O_1655,N_10022,N_12588);
nand UO_1656 (O_1656,N_10442,N_12061);
nand UO_1657 (O_1657,N_11094,N_13901);
and UO_1658 (O_1658,N_13199,N_11283);
nor UO_1659 (O_1659,N_11572,N_14112);
nand UO_1660 (O_1660,N_11737,N_13306);
and UO_1661 (O_1661,N_12281,N_13357);
nor UO_1662 (O_1662,N_12924,N_12451);
and UO_1663 (O_1663,N_10900,N_14097);
nor UO_1664 (O_1664,N_12952,N_14030);
and UO_1665 (O_1665,N_13321,N_13023);
nand UO_1666 (O_1666,N_10790,N_14518);
nor UO_1667 (O_1667,N_13158,N_11002);
nor UO_1668 (O_1668,N_12086,N_10516);
nor UO_1669 (O_1669,N_11842,N_12436);
nand UO_1670 (O_1670,N_10759,N_13183);
nand UO_1671 (O_1671,N_12721,N_14844);
or UO_1672 (O_1672,N_13691,N_12731);
xnor UO_1673 (O_1673,N_13908,N_10451);
or UO_1674 (O_1674,N_10922,N_13816);
xor UO_1675 (O_1675,N_13248,N_12322);
nand UO_1676 (O_1676,N_11595,N_13731);
nand UO_1677 (O_1677,N_13407,N_14633);
nor UO_1678 (O_1678,N_14470,N_12469);
nand UO_1679 (O_1679,N_12748,N_11373);
xor UO_1680 (O_1680,N_13462,N_11902);
and UO_1681 (O_1681,N_12675,N_12069);
nor UO_1682 (O_1682,N_12575,N_11562);
or UO_1683 (O_1683,N_13502,N_14312);
nor UO_1684 (O_1684,N_13520,N_10810);
and UO_1685 (O_1685,N_14046,N_10719);
and UO_1686 (O_1686,N_10016,N_14971);
or UO_1687 (O_1687,N_10460,N_11171);
nor UO_1688 (O_1688,N_14641,N_13633);
nor UO_1689 (O_1689,N_10498,N_14502);
or UO_1690 (O_1690,N_11786,N_13663);
xor UO_1691 (O_1691,N_11773,N_12826);
and UO_1692 (O_1692,N_10161,N_12057);
nand UO_1693 (O_1693,N_10086,N_12290);
nor UO_1694 (O_1694,N_13272,N_11889);
xnor UO_1695 (O_1695,N_13935,N_13677);
and UO_1696 (O_1696,N_11161,N_11053);
or UO_1697 (O_1697,N_14686,N_12112);
nand UO_1698 (O_1698,N_13445,N_11031);
nand UO_1699 (O_1699,N_12538,N_10339);
xor UO_1700 (O_1700,N_11731,N_14754);
nor UO_1701 (O_1701,N_13755,N_13135);
or UO_1702 (O_1702,N_11585,N_10162);
and UO_1703 (O_1703,N_12841,N_11754);
or UO_1704 (O_1704,N_11748,N_12475);
nand UO_1705 (O_1705,N_13925,N_13919);
nand UO_1706 (O_1706,N_10599,N_12990);
or UO_1707 (O_1707,N_14345,N_13531);
or UO_1708 (O_1708,N_11861,N_14655);
nor UO_1709 (O_1709,N_12099,N_14078);
or UO_1710 (O_1710,N_14277,N_13436);
or UO_1711 (O_1711,N_13962,N_10246);
and UO_1712 (O_1712,N_13824,N_11601);
nor UO_1713 (O_1713,N_13940,N_10716);
and UO_1714 (O_1714,N_13119,N_12318);
and UO_1715 (O_1715,N_13433,N_12543);
nand UO_1716 (O_1716,N_12218,N_10499);
xor UO_1717 (O_1717,N_11556,N_10041);
or UO_1718 (O_1718,N_11957,N_10564);
and UO_1719 (O_1719,N_14584,N_12949);
or UO_1720 (O_1720,N_11435,N_12784);
xor UO_1721 (O_1721,N_14572,N_14688);
and UO_1722 (O_1722,N_10882,N_10893);
nand UO_1723 (O_1723,N_10814,N_10429);
xor UO_1724 (O_1724,N_13264,N_14169);
or UO_1725 (O_1725,N_13748,N_14383);
nand UO_1726 (O_1726,N_14675,N_10051);
nand UO_1727 (O_1727,N_10219,N_12805);
nand UO_1728 (O_1728,N_14324,N_11796);
or UO_1729 (O_1729,N_14421,N_11285);
xor UO_1730 (O_1730,N_10439,N_14865);
nor UO_1731 (O_1731,N_14994,N_12940);
or UO_1732 (O_1732,N_10065,N_11855);
xor UO_1733 (O_1733,N_11619,N_14943);
xor UO_1734 (O_1734,N_14996,N_11577);
nor UO_1735 (O_1735,N_11091,N_12582);
nand UO_1736 (O_1736,N_10528,N_12874);
or UO_1737 (O_1737,N_10532,N_12517);
nor UO_1738 (O_1738,N_11343,N_12967);
nand UO_1739 (O_1739,N_10811,N_12972);
nand UO_1740 (O_1740,N_11501,N_14647);
and UO_1741 (O_1741,N_11762,N_12944);
or UO_1742 (O_1742,N_13820,N_13017);
nor UO_1743 (O_1743,N_12209,N_13841);
and UO_1744 (O_1744,N_13236,N_12701);
and UO_1745 (O_1745,N_14210,N_14018);
or UO_1746 (O_1746,N_13427,N_14529);
nand UO_1747 (O_1747,N_14325,N_11708);
or UO_1748 (O_1748,N_10266,N_12723);
nor UO_1749 (O_1749,N_10178,N_12828);
nor UO_1750 (O_1750,N_10667,N_14723);
nand UO_1751 (O_1751,N_12038,N_12587);
nor UO_1752 (O_1752,N_13328,N_12387);
nor UO_1753 (O_1753,N_12222,N_13883);
and UO_1754 (O_1754,N_13002,N_10374);
nand UO_1755 (O_1755,N_10990,N_13657);
or UO_1756 (O_1756,N_13733,N_13195);
nor UO_1757 (O_1757,N_13286,N_12419);
nand UO_1758 (O_1758,N_12915,N_13689);
nor UO_1759 (O_1759,N_11079,N_13971);
nand UO_1760 (O_1760,N_13001,N_14795);
xnor UO_1761 (O_1761,N_11035,N_11158);
and UO_1762 (O_1762,N_12961,N_14826);
and UO_1763 (O_1763,N_11116,N_13055);
nand UO_1764 (O_1764,N_14214,N_10463);
nor UO_1765 (O_1765,N_14188,N_14683);
or UO_1766 (O_1766,N_10100,N_10624);
or UO_1767 (O_1767,N_13346,N_11250);
nor UO_1768 (O_1768,N_10487,N_14024);
nor UO_1769 (O_1769,N_14189,N_13902);
xnor UO_1770 (O_1770,N_12202,N_14480);
xor UO_1771 (O_1771,N_11867,N_13267);
nor UO_1772 (O_1772,N_12996,N_14243);
or UO_1773 (O_1773,N_14192,N_14107);
nor UO_1774 (O_1774,N_14984,N_10924);
nand UO_1775 (O_1775,N_14085,N_12853);
nand UO_1776 (O_1776,N_10571,N_14389);
xnor UO_1777 (O_1777,N_11916,N_14505);
nand UO_1778 (O_1778,N_10312,N_10540);
and UO_1779 (O_1779,N_14563,N_13675);
and UO_1780 (O_1780,N_13958,N_12606);
nand UO_1781 (O_1781,N_13699,N_12311);
nor UO_1782 (O_1782,N_11835,N_10000);
and UO_1783 (O_1783,N_12754,N_13241);
nand UO_1784 (O_1784,N_12286,N_13421);
nor UO_1785 (O_1785,N_13131,N_12878);
nor UO_1786 (O_1786,N_14509,N_13728);
or UO_1787 (O_1787,N_10352,N_14444);
or UO_1788 (O_1788,N_10697,N_11075);
nand UO_1789 (O_1789,N_10005,N_10856);
or UO_1790 (O_1790,N_14286,N_12479);
xor UO_1791 (O_1791,N_10681,N_10084);
xnor UO_1792 (O_1792,N_14564,N_13275);
nor UO_1793 (O_1793,N_13031,N_11216);
nor UO_1794 (O_1794,N_10654,N_11626);
nand UO_1795 (O_1795,N_11057,N_14610);
and UO_1796 (O_1796,N_10840,N_10513);
or UO_1797 (O_1797,N_12203,N_12314);
nand UO_1798 (O_1798,N_12881,N_13054);
nand UO_1799 (O_1799,N_12388,N_13490);
nand UO_1800 (O_1800,N_13934,N_14797);
nand UO_1801 (O_1801,N_10967,N_13660);
and UO_1802 (O_1802,N_11608,N_14269);
or UO_1803 (O_1803,N_14791,N_10081);
or UO_1804 (O_1804,N_14062,N_12136);
nand UO_1805 (O_1805,N_14394,N_10337);
xnor UO_1806 (O_1806,N_14440,N_10010);
nor UO_1807 (O_1807,N_14866,N_10747);
nand UO_1808 (O_1808,N_11571,N_12005);
nor UO_1809 (O_1809,N_14084,N_13424);
or UO_1810 (O_1810,N_13930,N_12791);
or UO_1811 (O_1811,N_12553,N_12600);
nor UO_1812 (O_1812,N_12740,N_12895);
nand UO_1813 (O_1813,N_11097,N_11599);
or UO_1814 (O_1814,N_10682,N_11044);
and UO_1815 (O_1815,N_10240,N_10409);
or UO_1816 (O_1816,N_11586,N_14625);
or UO_1817 (O_1817,N_12151,N_11770);
xnor UO_1818 (O_1818,N_13104,N_10972);
nand UO_1819 (O_1819,N_13203,N_13911);
nor UO_1820 (O_1820,N_13535,N_13294);
nor UO_1821 (O_1821,N_10933,N_14508);
and UO_1822 (O_1822,N_14616,N_10047);
or UO_1823 (O_1823,N_13293,N_10090);
or UO_1824 (O_1824,N_11551,N_14674);
or UO_1825 (O_1825,N_11490,N_12037);
nor UO_1826 (O_1826,N_14002,N_11482);
or UO_1827 (O_1827,N_14160,N_12401);
nand UO_1828 (O_1828,N_14546,N_12158);
nor UO_1829 (O_1829,N_11624,N_12758);
nand UO_1830 (O_1830,N_14643,N_13439);
nand UO_1831 (O_1831,N_12257,N_10782);
nor UO_1832 (O_1832,N_10847,N_10256);
nand UO_1833 (O_1833,N_10660,N_11450);
or UO_1834 (O_1834,N_11396,N_12090);
nor UO_1835 (O_1835,N_12338,N_14855);
or UO_1836 (O_1836,N_12900,N_11155);
and UO_1837 (O_1837,N_13559,N_12183);
and UO_1838 (O_1838,N_13213,N_10045);
or UO_1839 (O_1839,N_14241,N_13312);
and UO_1840 (O_1840,N_10511,N_10313);
nand UO_1841 (O_1841,N_14544,N_11405);
nor UO_1842 (O_1842,N_11542,N_14934);
nor UO_1843 (O_1843,N_11308,N_11252);
nand UO_1844 (O_1844,N_11211,N_13319);
xor UO_1845 (O_1845,N_13128,N_12411);
or UO_1846 (O_1846,N_13291,N_13776);
or UO_1847 (O_1847,N_11922,N_12244);
xor UO_1848 (O_1848,N_10182,N_12781);
xnor UO_1849 (O_1849,N_14430,N_13937);
and UO_1850 (O_1850,N_12843,N_10140);
nor UO_1851 (O_1851,N_10721,N_12398);
nand UO_1852 (O_1852,N_10909,N_10386);
nand UO_1853 (O_1853,N_14063,N_14880);
or UO_1854 (O_1854,N_10508,N_11125);
nand UO_1855 (O_1855,N_10581,N_10687);
or UO_1856 (O_1856,N_13126,N_13815);
or UO_1857 (O_1857,N_11114,N_14733);
or UO_1858 (O_1858,N_13625,N_10114);
and UO_1859 (O_1859,N_11175,N_11990);
nand UO_1860 (O_1860,N_12703,N_12373);
nand UO_1861 (O_1861,N_10717,N_13796);
nand UO_1862 (O_1862,N_14051,N_10750);
and UO_1863 (O_1863,N_10163,N_14348);
and UO_1864 (O_1864,N_12013,N_13720);
nor UO_1865 (O_1865,N_14056,N_14127);
nor UO_1866 (O_1866,N_12349,N_14957);
and UO_1867 (O_1867,N_13298,N_13081);
or UO_1868 (O_1868,N_13600,N_13488);
and UO_1869 (O_1869,N_11115,N_12676);
or UO_1870 (O_1870,N_13612,N_11262);
xor UO_1871 (O_1871,N_13399,N_14012);
or UO_1872 (O_1872,N_14176,N_10699);
or UO_1873 (O_1873,N_14837,N_11881);
or UO_1874 (O_1874,N_10622,N_12065);
nand UO_1875 (O_1875,N_12724,N_11312);
nor UO_1876 (O_1876,N_11388,N_10668);
or UO_1877 (O_1877,N_14721,N_10507);
and UO_1878 (O_1878,N_11449,N_13556);
or UO_1879 (O_1879,N_14979,N_12666);
nand UO_1880 (O_1880,N_12581,N_13177);
or UO_1881 (O_1881,N_11908,N_12628);
xnor UO_1882 (O_1882,N_12131,N_10519);
nand UO_1883 (O_1883,N_13984,N_12893);
and UO_1884 (O_1884,N_10362,N_13751);
nand UO_1885 (O_1885,N_11452,N_13530);
and UO_1886 (O_1886,N_10464,N_10493);
or UO_1887 (O_1887,N_12343,N_13034);
xnor UO_1888 (O_1888,N_14967,N_11877);
nor UO_1889 (O_1889,N_11547,N_14906);
nor UO_1890 (O_1890,N_10306,N_14364);
and UO_1891 (O_1891,N_12109,N_13043);
and UO_1892 (O_1892,N_12590,N_10290);
nor UO_1893 (O_1893,N_11505,N_13981);
or UO_1894 (O_1894,N_13029,N_11113);
xor UO_1895 (O_1895,N_12030,N_14298);
or UO_1896 (O_1896,N_14384,N_11032);
nor UO_1897 (O_1897,N_14057,N_14156);
nand UO_1898 (O_1898,N_11688,N_12788);
nand UO_1899 (O_1899,N_14902,N_10928);
nor UO_1900 (O_1900,N_10921,N_12860);
or UO_1901 (O_1901,N_11558,N_10828);
nand UO_1902 (O_1902,N_11617,N_12128);
nand UO_1903 (O_1903,N_11460,N_11188);
nand UO_1904 (O_1904,N_14259,N_13996);
or UO_1905 (O_1905,N_11733,N_13337);
and UO_1906 (O_1906,N_12114,N_13118);
or UO_1907 (O_1907,N_12101,N_14863);
nand UO_1908 (O_1908,N_12140,N_10204);
nand UO_1909 (O_1909,N_11427,N_10023);
and UO_1910 (O_1910,N_11841,N_12901);
and UO_1911 (O_1911,N_10318,N_10533);
or UO_1912 (O_1912,N_14350,N_10142);
and UO_1913 (O_1913,N_14293,N_14517);
nor UO_1914 (O_1914,N_13948,N_10748);
and UO_1915 (O_1915,N_14947,N_14634);
or UO_1916 (O_1916,N_10490,N_14736);
nor UO_1917 (O_1917,N_13904,N_11302);
nor UO_1918 (O_1918,N_13608,N_14519);
xor UO_1919 (O_1919,N_11047,N_14090);
nand UO_1920 (O_1920,N_12870,N_13661);
nor UO_1921 (O_1921,N_13857,N_10500);
nor UO_1922 (O_1922,N_13154,N_13717);
and UO_1923 (O_1923,N_10066,N_14132);
nand UO_1924 (O_1924,N_11476,N_11123);
or UO_1925 (O_1925,N_14807,N_13027);
nand UO_1926 (O_1926,N_13609,N_14933);
nand UO_1927 (O_1927,N_14881,N_11667);
nor UO_1928 (O_1928,N_11668,N_12845);
nor UO_1929 (O_1929,N_12621,N_10459);
nand UO_1930 (O_1930,N_12638,N_10677);
or UO_1931 (O_1931,N_11996,N_10002);
or UO_1932 (O_1932,N_12647,N_13601);
or UO_1933 (O_1933,N_14580,N_14485);
or UO_1934 (O_1934,N_11899,N_11707);
nand UO_1935 (O_1935,N_14065,N_11245);
and UO_1936 (O_1936,N_10689,N_14007);
xor UO_1937 (O_1937,N_10992,N_10908);
and UO_1938 (O_1938,N_12777,N_13701);
and UO_1939 (O_1939,N_11072,N_12579);
nor UO_1940 (O_1940,N_13775,N_10174);
nand UO_1941 (O_1941,N_14917,N_14115);
nand UO_1942 (O_1942,N_12223,N_11232);
and UO_1943 (O_1943,N_13364,N_13007);
nor UO_1944 (O_1944,N_14981,N_12488);
nor UO_1945 (O_1945,N_12344,N_10773);
or UO_1946 (O_1946,N_12348,N_12273);
nand UO_1947 (O_1947,N_12212,N_11974);
or UO_1948 (O_1948,N_12745,N_12135);
nand UO_1949 (O_1949,N_13309,N_12680);
or UO_1950 (O_1950,N_10578,N_14402);
nand UO_1951 (O_1951,N_14231,N_10589);
or UO_1952 (O_1952,N_13114,N_10214);
nor UO_1953 (O_1953,N_10166,N_14045);
nor UO_1954 (O_1954,N_14126,N_13800);
or UO_1955 (O_1955,N_13476,N_12068);
nor UO_1956 (O_1956,N_12547,N_10227);
or UO_1957 (O_1957,N_10761,N_12431);
xor UO_1958 (O_1958,N_10808,N_14551);
and UO_1959 (O_1959,N_12504,N_12978);
xnor UO_1960 (O_1960,N_10696,N_14527);
nor UO_1961 (O_1961,N_14871,N_11003);
or UO_1962 (O_1962,N_10383,N_13756);
xor UO_1963 (O_1963,N_11239,N_11219);
nor UO_1964 (O_1964,N_10543,N_12254);
nand UO_1965 (O_1965,N_14428,N_14603);
or UO_1966 (O_1966,N_14060,N_11364);
xor UO_1967 (O_1967,N_12605,N_13061);
xnor UO_1968 (O_1968,N_12916,N_10521);
xnor UO_1969 (O_1969,N_14353,N_13526);
or UO_1970 (O_1970,N_12838,N_11258);
or UO_1971 (O_1971,N_10403,N_14100);
or UO_1972 (O_1972,N_14019,N_13282);
nand UO_1973 (O_1973,N_14075,N_13088);
nand UO_1974 (O_1974,N_13577,N_12080);
or UO_1975 (O_1975,N_13136,N_12377);
nor UO_1976 (O_1976,N_13216,N_12981);
or UO_1977 (O_1977,N_14888,N_12858);
nand UO_1978 (O_1978,N_12726,N_13456);
or UO_1979 (O_1979,N_11677,N_13044);
nor UO_1980 (O_1980,N_12247,N_13705);
and UO_1981 (O_1981,N_14832,N_14914);
or UO_1982 (O_1982,N_14211,N_10307);
xnor UO_1983 (O_1983,N_11402,N_13897);
or UO_1984 (O_1984,N_14358,N_11832);
nor UO_1985 (O_1985,N_11837,N_11808);
nand UO_1986 (O_1986,N_12017,N_13947);
nor UO_1987 (O_1987,N_13513,N_11592);
and UO_1988 (O_1988,N_10422,N_13377);
or UO_1989 (O_1989,N_12823,N_13868);
xnor UO_1990 (O_1990,N_11088,N_12875);
nand UO_1991 (O_1991,N_12634,N_11678);
nor UO_1992 (O_1992,N_14680,N_13449);
nand UO_1993 (O_1993,N_11909,N_11658);
nand UO_1994 (O_1994,N_11217,N_10391);
nor UO_1995 (O_1995,N_14197,N_13665);
xor UO_1996 (O_1996,N_12631,N_12298);
nor UO_1997 (O_1997,N_13070,N_11139);
and UO_1998 (O_1998,N_10424,N_13744);
nand UO_1999 (O_1999,N_10418,N_14308);
endmodule