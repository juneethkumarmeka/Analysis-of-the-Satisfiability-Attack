module basic_5000_50000_5000_20_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
xor U0 (N_0,In_1700,In_561);
and U1 (N_1,In_2626,In_1766);
or U2 (N_2,In_4492,In_4199);
or U3 (N_3,In_489,In_3166);
or U4 (N_4,In_4298,In_1007);
nor U5 (N_5,In_4488,In_4621);
nand U6 (N_6,In_1373,In_1817);
or U7 (N_7,In_4242,In_2292);
nand U8 (N_8,In_3232,In_1089);
and U9 (N_9,In_2997,In_2212);
and U10 (N_10,In_4524,In_4062);
nand U11 (N_11,In_3975,In_2296);
xnor U12 (N_12,In_3840,In_2681);
xnor U13 (N_13,In_4831,In_1831);
nand U14 (N_14,In_1711,In_3401);
and U15 (N_15,In_3842,In_2052);
xor U16 (N_16,In_501,In_4160);
and U17 (N_17,In_2353,In_3866);
xnor U18 (N_18,In_4181,In_4750);
nor U19 (N_19,In_3294,In_1465);
or U20 (N_20,In_3947,In_1548);
nor U21 (N_21,In_3884,In_4201);
and U22 (N_22,In_3501,In_4216);
nor U23 (N_23,In_3107,In_2173);
or U24 (N_24,In_941,In_3353);
nor U25 (N_25,In_2555,In_3986);
nand U26 (N_26,In_1922,In_2197);
or U27 (N_27,In_4941,In_1463);
nor U28 (N_28,In_642,In_3678);
nor U29 (N_29,In_3769,In_4790);
or U30 (N_30,In_4183,In_3360);
and U31 (N_31,In_3637,In_2265);
and U32 (N_32,In_953,In_4195);
and U33 (N_33,In_388,In_3803);
nor U34 (N_34,In_4102,In_848);
or U35 (N_35,In_2479,In_4397);
and U36 (N_36,In_267,In_4832);
or U37 (N_37,In_2911,In_4047);
or U38 (N_38,In_4811,In_1311);
or U39 (N_39,In_4786,In_1347);
or U40 (N_40,In_4755,In_3454);
or U41 (N_41,In_3466,In_4280);
nand U42 (N_42,In_422,In_2102);
xnor U43 (N_43,In_4079,In_3811);
and U44 (N_44,In_4198,In_400);
and U45 (N_45,In_627,In_236);
or U46 (N_46,In_2427,In_620);
or U47 (N_47,In_3080,In_4515);
xnor U48 (N_48,In_453,In_1083);
or U49 (N_49,In_377,In_1818);
or U50 (N_50,In_1540,In_3263);
nand U51 (N_51,In_3764,In_262);
and U52 (N_52,In_4539,In_793);
xor U53 (N_53,In_1858,In_3922);
nand U54 (N_54,In_3389,In_630);
and U55 (N_55,In_4628,In_1549);
nand U56 (N_56,In_3442,In_314);
and U57 (N_57,In_307,In_3517);
xor U58 (N_58,In_1014,In_2431);
xnor U59 (N_59,In_2940,In_4306);
xnor U60 (N_60,In_49,In_2299);
xor U61 (N_61,In_2652,In_4262);
xnor U62 (N_62,In_4632,In_3753);
or U63 (N_63,In_2313,In_329);
and U64 (N_64,In_2340,In_185);
nor U65 (N_65,In_2915,In_4050);
and U66 (N_66,In_2149,In_4999);
xnor U67 (N_67,In_799,In_3857);
nor U68 (N_68,In_4871,In_302);
or U69 (N_69,In_3139,In_27);
or U70 (N_70,In_2241,In_2395);
nor U71 (N_71,In_1130,In_4029);
or U72 (N_72,In_3807,In_2795);
nor U73 (N_73,In_2889,In_4646);
or U74 (N_74,In_3689,In_3621);
and U75 (N_75,In_474,In_1026);
and U76 (N_76,In_2247,In_4509);
xor U77 (N_77,In_4133,In_1341);
or U78 (N_78,In_2415,In_2642);
and U79 (N_79,In_2097,In_2971);
nor U80 (N_80,In_3130,In_1087);
xor U81 (N_81,In_2138,In_3108);
xor U82 (N_82,In_4481,In_749);
nor U83 (N_83,In_2633,In_4144);
and U84 (N_84,In_1616,In_4041);
xnor U85 (N_85,In_2569,In_3687);
nand U86 (N_86,In_356,In_4208);
and U87 (N_87,In_2288,In_2957);
nor U88 (N_88,In_3437,In_4318);
nand U89 (N_89,In_733,In_4876);
nor U90 (N_90,In_1919,In_3522);
nand U91 (N_91,In_4446,In_3252);
nand U92 (N_92,In_615,In_4759);
and U93 (N_93,In_1173,In_2846);
xnor U94 (N_94,In_1245,In_1969);
xor U95 (N_95,In_891,In_3780);
nor U96 (N_96,In_2743,In_831);
nor U97 (N_97,In_2105,In_2703);
or U98 (N_98,In_4223,In_1501);
xnor U99 (N_99,In_160,In_3830);
and U100 (N_100,In_3644,In_3729);
or U101 (N_101,In_4954,In_732);
nor U102 (N_102,In_4091,In_881);
nand U103 (N_103,In_766,In_3336);
nand U104 (N_104,In_3077,In_2770);
xnor U105 (N_105,In_3709,In_3755);
nand U106 (N_106,In_4374,In_2949);
nand U107 (N_107,In_762,In_463);
nor U108 (N_108,In_3193,In_1231);
nand U109 (N_109,In_1637,In_1183);
and U110 (N_110,In_2399,In_2028);
nand U111 (N_111,In_4417,In_3276);
xnor U112 (N_112,In_450,In_3874);
xor U113 (N_113,In_317,In_40);
xnor U114 (N_114,In_297,In_3520);
xnor U115 (N_115,In_445,In_2482);
and U116 (N_116,In_1170,In_604);
nor U117 (N_117,In_4136,In_1495);
nand U118 (N_118,In_4219,In_2640);
and U119 (N_119,In_2628,In_2794);
nand U120 (N_120,In_504,In_3950);
nor U121 (N_121,In_1342,In_3296);
and U122 (N_122,In_1984,In_1456);
xnor U123 (N_123,In_4114,In_3714);
xnor U124 (N_124,In_1684,In_3576);
nand U125 (N_125,In_696,In_2434);
and U126 (N_126,In_4415,In_1203);
and U127 (N_127,In_4897,In_2538);
nor U128 (N_128,In_2301,In_2203);
xor U129 (N_129,In_4536,In_4347);
or U130 (N_130,In_3225,In_2043);
nand U131 (N_131,In_3660,In_2358);
or U132 (N_132,In_2025,In_4159);
nand U133 (N_133,In_4889,In_3904);
and U134 (N_134,In_82,In_715);
or U135 (N_135,In_1195,In_2455);
nor U136 (N_136,In_3335,In_917);
xnor U137 (N_137,In_2049,In_992);
xnor U138 (N_138,In_2179,In_1079);
nand U139 (N_139,In_181,In_2088);
or U140 (N_140,In_2541,In_3777);
nor U141 (N_141,In_477,In_381);
nor U142 (N_142,In_10,In_3916);
nor U143 (N_143,In_3743,In_3487);
xnor U144 (N_144,In_3284,In_791);
nand U145 (N_145,In_4233,In_745);
and U146 (N_146,In_4443,In_3843);
nand U147 (N_147,In_2848,In_4361);
nand U148 (N_148,In_190,In_4908);
and U149 (N_149,In_1846,In_1849);
xor U150 (N_150,In_2896,In_89);
nor U151 (N_151,In_4752,In_2876);
or U152 (N_152,In_4020,In_901);
nand U153 (N_153,In_2375,In_3515);
nand U154 (N_154,In_4192,In_2214);
xor U155 (N_155,In_4804,In_940);
and U156 (N_156,In_4528,In_134);
xnor U157 (N_157,In_4513,In_2542);
or U158 (N_158,In_1688,In_786);
xnor U159 (N_159,In_3577,In_908);
and U160 (N_160,In_2035,In_2412);
xnor U161 (N_161,In_3929,In_214);
xnor U162 (N_162,In_3741,In_2580);
or U163 (N_163,In_3834,In_2689);
xor U164 (N_164,In_4141,In_610);
xor U165 (N_165,In_4931,In_122);
or U166 (N_166,In_380,In_1242);
or U167 (N_167,In_800,In_2958);
nand U168 (N_168,In_1571,In_3779);
xor U169 (N_169,In_11,In_2788);
nand U170 (N_170,In_2638,In_3949);
nand U171 (N_171,In_1981,In_4266);
and U172 (N_172,In_2967,In_3273);
nand U173 (N_173,In_3901,In_4578);
nand U174 (N_174,In_1980,In_2491);
nor U175 (N_175,In_492,In_2665);
xor U176 (N_176,In_187,In_3176);
nor U177 (N_177,In_470,In_4211);
xor U178 (N_178,In_4964,In_2091);
or U179 (N_179,In_2120,In_622);
and U180 (N_180,In_3398,In_1398);
nor U181 (N_181,In_1836,In_2079);
nor U182 (N_182,In_3253,In_2366);
nand U183 (N_183,In_2547,In_631);
nand U184 (N_184,In_1985,In_4658);
nand U185 (N_185,In_3793,In_6);
and U186 (N_186,In_4129,In_3763);
xor U187 (N_187,In_867,In_1277);
nand U188 (N_188,In_3892,In_4953);
nand U189 (N_189,In_4801,In_687);
or U190 (N_190,In_4324,In_2089);
xnor U191 (N_191,In_3008,In_2956);
or U192 (N_192,In_4344,In_163);
or U193 (N_193,In_3505,In_807);
nor U194 (N_194,In_3756,In_1955);
and U195 (N_195,In_4231,In_2080);
and U196 (N_196,In_943,In_1075);
nor U197 (N_197,In_2895,In_2706);
nor U198 (N_198,In_781,In_3732);
nand U199 (N_199,In_3765,In_3485);
and U200 (N_200,In_4793,In_3731);
and U201 (N_201,In_4603,In_4264);
nor U202 (N_202,In_1214,In_741);
or U203 (N_203,In_3509,In_1826);
and U204 (N_204,In_430,In_2112);
and U205 (N_205,In_1941,In_1620);
or U206 (N_206,In_3425,In_4990);
or U207 (N_207,In_3733,In_70);
nor U208 (N_208,In_2015,In_1359);
or U209 (N_209,In_3532,In_4044);
nand U210 (N_210,In_3529,In_4402);
nor U211 (N_211,In_554,In_363);
or U212 (N_212,In_1496,In_227);
nor U213 (N_213,In_2072,In_3103);
and U214 (N_214,In_3980,In_4304);
xor U215 (N_215,In_3951,In_462);
and U216 (N_216,In_1161,In_997);
and U217 (N_217,In_4084,In_3625);
xor U218 (N_218,In_3792,In_1899);
nand U219 (N_219,In_280,In_3898);
or U220 (N_220,In_4377,In_2466);
nor U221 (N_221,In_544,In_4185);
nor U222 (N_222,In_1845,In_1679);
or U223 (N_223,In_4436,In_4637);
nand U224 (N_224,In_1215,In_3664);
or U225 (N_225,In_1697,In_1597);
nand U226 (N_226,In_413,In_958);
nor U227 (N_227,In_1361,In_2832);
xor U228 (N_228,In_3682,In_3183);
xor U229 (N_229,In_4860,In_2501);
or U230 (N_230,In_2209,In_3169);
nand U231 (N_231,In_678,In_2118);
nand U232 (N_232,In_3340,In_735);
nor U233 (N_233,In_4093,In_4367);
nand U234 (N_234,In_2732,In_2239);
xnor U235 (N_235,In_2750,In_4497);
and U236 (N_236,In_3343,In_312);
xnor U237 (N_237,In_2014,In_4314);
or U238 (N_238,In_3945,In_3323);
and U239 (N_239,In_1656,In_1712);
nor U240 (N_240,In_3527,In_4935);
xnor U241 (N_241,In_4085,In_3146);
or U242 (N_242,In_4799,In_487);
and U243 (N_243,In_728,In_3278);
or U244 (N_244,In_2483,In_2158);
and U245 (N_245,In_140,In_2230);
nor U246 (N_246,In_4498,In_1614);
or U247 (N_247,In_4457,In_4918);
nand U248 (N_248,In_2568,In_2755);
xnor U249 (N_249,In_3698,In_2615);
xor U250 (N_250,In_63,In_3988);
nor U251 (N_251,In_3317,In_330);
and U252 (N_252,In_4901,In_4857);
nor U253 (N_253,In_399,In_4239);
and U254 (N_254,In_3405,In_811);
or U255 (N_255,In_361,In_3414);
or U256 (N_256,In_1200,In_3470);
nor U257 (N_257,In_2669,In_4945);
xnor U258 (N_258,In_551,In_3472);
xnor U259 (N_259,In_2360,In_577);
and U260 (N_260,In_1728,In_659);
xor U261 (N_261,In_3014,In_1362);
and U262 (N_262,In_1098,In_661);
or U263 (N_263,In_2053,In_2180);
nor U264 (N_264,In_2887,In_4355);
nor U265 (N_265,In_1393,In_2965);
xor U266 (N_266,In_1041,In_4977);
and U267 (N_267,In_3806,In_524);
or U268 (N_268,In_3519,In_1360);
nand U269 (N_269,In_3966,In_3381);
nor U270 (N_270,In_4994,In_2013);
or U271 (N_271,In_4618,In_4516);
xor U272 (N_272,In_3248,In_1392);
or U273 (N_273,In_1211,In_4422);
or U274 (N_274,In_537,In_2700);
xnor U275 (N_275,In_1686,In_407);
xor U276 (N_276,In_198,In_195);
or U277 (N_277,In_4914,In_4021);
xnor U278 (N_278,In_2040,In_419);
xor U279 (N_279,In_3967,In_465);
or U280 (N_280,In_1583,In_3067);
nor U281 (N_281,In_1879,In_4012);
xor U282 (N_282,In_1598,In_2338);
nand U283 (N_283,In_2246,In_2060);
and U284 (N_284,In_3750,In_1366);
nand U285 (N_285,In_532,In_981);
or U286 (N_286,In_3586,In_75);
xor U287 (N_287,In_3566,In_1269);
and U288 (N_288,In_1542,In_904);
or U289 (N_289,In_1971,In_3483);
xor U290 (N_290,In_4451,In_1988);
nor U291 (N_291,In_1233,In_3942);
and U292 (N_292,In_1666,In_736);
xnor U293 (N_293,In_2909,In_3770);
or U294 (N_294,In_2469,In_3100);
or U295 (N_295,In_4385,In_3259);
xor U296 (N_296,In_2756,In_1085);
nand U297 (N_297,In_268,In_2557);
xor U298 (N_298,In_2121,In_3507);
nand U299 (N_299,In_1380,In_2018);
nand U300 (N_300,In_1774,In_2565);
nor U301 (N_301,In_4569,In_3998);
nand U302 (N_302,In_1049,In_1555);
nand U303 (N_303,In_1144,In_3106);
and U304 (N_304,In_2521,In_2868);
and U305 (N_305,In_2090,In_116);
nor U306 (N_306,In_1272,In_4576);
nand U307 (N_307,In_1088,In_1095);
xnor U308 (N_308,In_3616,In_4106);
nand U309 (N_309,In_2923,In_1478);
and U310 (N_310,In_1934,In_779);
nor U311 (N_311,In_4297,In_798);
or U312 (N_312,In_1338,In_4372);
and U313 (N_313,In_841,In_4137);
nor U314 (N_314,In_115,In_1454);
xnor U315 (N_315,In_3025,In_2444);
nand U316 (N_316,In_744,In_2720);
nor U317 (N_317,In_3555,In_1678);
nor U318 (N_318,In_318,In_4709);
nand U319 (N_319,In_3627,In_4157);
nor U320 (N_320,In_2948,In_2471);
nand U321 (N_321,In_3020,In_4563);
or U322 (N_322,In_747,In_1396);
nor U323 (N_323,In_3290,In_2405);
or U324 (N_324,In_1662,In_4321);
or U325 (N_325,In_3283,In_2352);
xnor U326 (N_326,In_3222,In_4890);
nand U327 (N_327,In_2477,In_3663);
nand U328 (N_328,In_3933,In_2063);
nor U329 (N_329,In_566,In_4295);
nand U330 (N_330,In_2506,In_1695);
nor U331 (N_331,In_4476,In_2524);
and U332 (N_332,In_4676,In_442);
and U333 (N_333,In_4340,In_510);
nor U334 (N_334,In_259,In_16);
and U335 (N_335,In_3861,In_1512);
nor U336 (N_336,In_3081,In_990);
or U337 (N_337,In_2485,In_816);
xor U338 (N_338,In_3113,In_1343);
nand U339 (N_339,In_1869,In_2082);
and U340 (N_340,In_2251,In_2882);
and U341 (N_341,In_258,In_3172);
or U342 (N_342,In_2242,In_3280);
xnor U343 (N_343,In_2027,In_1125);
and U344 (N_344,In_1467,In_4325);
nor U345 (N_345,In_506,In_241);
nand U346 (N_346,In_3603,In_4026);
and U347 (N_347,In_2746,In_797);
nor U348 (N_348,In_3416,In_2658);
and U349 (N_349,In_4859,In_1994);
and U350 (N_350,In_4835,In_1682);
or U351 (N_351,In_2019,In_217);
or U352 (N_352,In_906,In_4809);
or U353 (N_353,In_3030,In_2843);
nand U354 (N_354,In_4405,In_4473);
nand U355 (N_355,In_2294,In_1237);
and U356 (N_356,In_1880,In_125);
and U357 (N_357,In_2,In_1395);
and U358 (N_358,In_345,In_3123);
nor U359 (N_359,In_1166,In_3821);
and U360 (N_360,In_4822,In_730);
or U361 (N_361,In_4568,In_662);
xor U362 (N_362,In_2677,In_4130);
or U363 (N_363,In_3590,In_3269);
or U364 (N_364,In_3299,In_3907);
or U365 (N_365,In_4139,In_271);
and U366 (N_366,In_4903,In_4283);
or U367 (N_367,In_4919,In_2614);
nand U368 (N_368,In_651,In_2048);
or U369 (N_369,In_4033,In_4693);
xnor U370 (N_370,In_3395,In_580);
nand U371 (N_371,In_2883,In_1931);
nand U372 (N_372,In_15,In_682);
and U373 (N_373,In_151,In_505);
nor U374 (N_374,In_3746,In_2183);
nand U375 (N_375,In_3924,In_2199);
nand U376 (N_376,In_3881,In_3011);
or U377 (N_377,In_669,In_3339);
nand U378 (N_378,In_2588,In_3013);
nor U379 (N_379,In_1607,In_2920);
xor U380 (N_380,In_4191,In_4595);
xor U381 (N_381,In_437,In_4175);
or U382 (N_382,In_2596,In_2168);
and U383 (N_383,In_677,In_548);
nor U384 (N_384,In_438,In_2100);
xnor U385 (N_385,In_4128,In_495);
nor U386 (N_386,In_288,In_1596);
nor U387 (N_387,In_1929,In_974);
and U388 (N_388,In_640,In_1693);
nand U389 (N_389,In_2221,In_2969);
nor U390 (N_390,In_3496,In_595);
xor U391 (N_391,In_1725,In_2845);
nor U392 (N_392,In_1767,In_3363);
xnor U393 (N_393,In_1406,In_1517);
xnor U394 (N_394,In_859,In_3265);
nor U395 (N_395,In_2440,In_4588);
and U396 (N_396,In_3293,In_3835);
nand U397 (N_397,In_664,In_4644);
and U398 (N_398,In_4712,In_1781);
and U399 (N_399,In_1107,In_1574);
nand U400 (N_400,In_4484,In_1802);
nor U401 (N_401,In_4565,In_2675);
and U402 (N_402,In_2618,In_230);
or U403 (N_403,In_371,In_309);
xnor U404 (N_404,In_1726,In_1350);
nor U405 (N_405,In_2092,In_2961);
nand U406 (N_406,In_603,In_2085);
xnor U407 (N_407,In_1627,In_468);
nand U408 (N_408,In_3128,In_4757);
xor U409 (N_409,In_4928,In_4572);
or U410 (N_410,In_4459,In_1553);
xor U411 (N_411,In_1696,In_2438);
nand U412 (N_412,In_713,In_3592);
xnor U413 (N_413,In_59,In_1405);
nor U414 (N_414,In_3480,In_3179);
nand U415 (N_415,In_4881,In_2315);
xor U416 (N_416,In_1873,In_4791);
or U417 (N_417,In_3112,In_4710);
nand U418 (N_418,In_3258,In_2106);
and U419 (N_419,In_4504,In_1485);
xor U420 (N_420,In_2844,In_1308);
or U421 (N_421,In_4132,In_3665);
and U422 (N_422,In_1992,In_201);
nor U423 (N_423,In_2371,In_3332);
and U424 (N_424,In_1212,In_1068);
xor U425 (N_425,In_26,In_1702);
and U426 (N_426,In_2222,In_4827);
nor U427 (N_427,In_4071,In_2680);
or U428 (N_428,In_2935,In_2817);
and U429 (N_429,In_2684,In_1073);
or U430 (N_430,In_2777,In_2177);
and U431 (N_431,In_2321,In_2289);
and U432 (N_432,In_39,In_1246);
nand U433 (N_433,In_2074,In_4046);
xnor U434 (N_434,In_61,In_4877);
nor U435 (N_435,In_3745,In_4165);
xnor U436 (N_436,In_1012,In_2649);
nand U437 (N_437,In_4329,In_4200);
nand U438 (N_438,In_2779,In_562);
nand U439 (N_439,In_4022,In_7);
nand U440 (N_440,In_3187,In_2824);
nor U441 (N_441,In_3679,In_606);
and U442 (N_442,In_4169,In_2853);
nor U443 (N_443,In_2164,In_4917);
nand U444 (N_444,In_4898,In_4075);
xnor U445 (N_445,In_1851,In_2548);
and U446 (N_446,In_4925,In_359);
nand U447 (N_447,In_4483,In_355);
xnor U448 (N_448,In_1008,In_1481);
nand U449 (N_449,In_2486,In_4273);
nand U450 (N_450,In_3328,In_3799);
and U451 (N_451,In_2211,In_4713);
or U452 (N_452,In_1050,In_1243);
nand U453 (N_453,In_4956,In_4474);
xnor U454 (N_454,In_1102,In_3262);
xor U455 (N_455,In_4055,In_3148);
nor U456 (N_456,In_691,In_2855);
xor U457 (N_457,In_480,In_4888);
nand U458 (N_458,In_1652,In_2503);
nand U459 (N_459,In_2809,In_2009);
nor U460 (N_460,In_3870,In_4230);
xor U461 (N_461,In_2269,In_2724);
and U462 (N_462,In_2616,In_3662);
and U463 (N_463,In_4444,In_349);
nand U464 (N_464,In_3019,In_3184);
nand U465 (N_465,In_3740,In_1151);
or U466 (N_466,In_725,In_4867);
or U467 (N_467,In_4270,In_498);
nand U468 (N_468,In_2805,In_2229);
and U469 (N_469,In_4048,In_714);
nand U470 (N_470,In_4196,In_1755);
nor U471 (N_471,In_789,In_738);
xnor U472 (N_472,In_4096,In_210);
or U473 (N_473,In_3261,In_1643);
nand U474 (N_474,In_1986,In_3138);
nor U475 (N_475,In_3917,In_1256);
and U476 (N_476,In_1967,In_4217);
and U477 (N_477,In_3046,In_1262);
xnor U478 (N_478,In_1156,In_81);
nor U479 (N_479,In_1197,In_4316);
and U480 (N_480,In_826,In_3221);
or U481 (N_481,In_1670,In_3506);
xor U482 (N_482,In_3704,In_4627);
xnor U483 (N_483,In_724,In_3127);
xnor U484 (N_484,In_1267,In_2166);
and U485 (N_485,In_3692,In_1832);
nor U486 (N_486,In_3026,In_3147);
or U487 (N_487,In_256,In_3475);
and U488 (N_488,In_539,In_790);
xor U489 (N_489,In_3070,In_4927);
xnor U490 (N_490,In_3612,In_3163);
and U491 (N_491,In_3045,In_1641);
xor U492 (N_492,In_4651,In_4054);
or U493 (N_493,In_3552,In_1149);
nor U494 (N_494,In_1152,In_885);
nor U495 (N_495,In_2813,In_2862);
or U496 (N_496,In_3034,In_3498);
and U497 (N_497,In_4471,In_2828);
nor U498 (N_498,In_4662,In_1539);
or U499 (N_499,In_3648,In_576);
nand U500 (N_500,In_1743,In_1825);
xor U501 (N_501,In_1524,In_85);
xnor U502 (N_502,In_2760,In_1507);
nor U503 (N_503,In_2627,In_3432);
and U504 (N_504,In_1282,In_4687);
nand U505 (N_505,In_1676,In_1569);
nand U506 (N_506,In_3926,In_1636);
nand U507 (N_507,In_2637,In_2916);
and U508 (N_508,In_1490,In_2898);
nor U509 (N_509,In_3076,In_3645);
nand U510 (N_510,In_4031,In_2372);
nor U511 (N_511,In_2578,In_4425);
nor U512 (N_512,In_285,In_4380);
nand U513 (N_513,In_466,In_530);
nand U514 (N_514,In_846,In_609);
nand U515 (N_515,In_761,In_3934);
and U516 (N_516,In_1281,In_666);
nand U517 (N_517,In_31,In_1091);
nor U518 (N_518,In_1615,In_2749);
or U519 (N_519,In_2624,In_2530);
and U520 (N_520,In_2235,In_2467);
nor U521 (N_521,In_2492,In_835);
nor U522 (N_522,In_3906,In_396);
nor U523 (N_523,In_4767,In_815);
nor U524 (N_524,In_3611,In_2807);
and U525 (N_525,In_2202,In_896);
nand U526 (N_526,In_4741,In_2531);
nor U527 (N_527,In_3229,In_3905);
nor U528 (N_528,In_344,In_1045);
and U529 (N_529,In_3715,In_4970);
and U530 (N_530,In_2396,In_3444);
xor U531 (N_531,In_2661,In_3383);
nand U532 (N_532,In_2701,In_2586);
nand U533 (N_533,In_2870,In_4580);
or U534 (N_534,In_4313,In_2116);
nor U535 (N_535,In_1017,In_2122);
nor U536 (N_536,In_2816,In_3460);
and U537 (N_537,In_2219,In_2857);
or U538 (N_538,In_1097,In_4345);
and U539 (N_539,In_4490,In_2157);
nand U540 (N_540,In_601,In_2767);
or U541 (N_541,In_431,In_4486);
or U542 (N_542,In_808,In_2990);
xnor U543 (N_543,In_686,In_771);
or U544 (N_544,In_1074,In_4787);
xnor U545 (N_545,In_3914,In_2488);
xnor U546 (N_546,In_1179,In_4449);
or U547 (N_547,In_868,In_4838);
nand U548 (N_548,In_4996,In_257);
and U549 (N_549,In_1672,In_3990);
or U550 (N_550,In_265,In_240);
and U551 (N_551,In_4697,In_4496);
xor U552 (N_552,In_2291,In_4802);
and U553 (N_553,In_1915,In_932);
or U554 (N_554,In_22,In_2858);
nor U555 (N_555,In_2549,In_2449);
and U556 (N_556,In_586,In_3632);
and U557 (N_557,In_4749,In_2610);
or U558 (N_558,In_4991,In_3808);
nand U559 (N_559,In_2348,In_4535);
xnor U560 (N_560,In_3338,In_2917);
and U561 (N_561,In_2475,In_2678);
nor U562 (N_562,In_4883,In_2963);
xor U563 (N_563,In_4064,In_4816);
or U564 (N_564,In_649,In_571);
xor U565 (N_565,In_3826,In_1909);
xor U566 (N_566,In_2020,In_1119);
xnor U567 (N_567,In_2005,In_3385);
and U568 (N_568,In_3408,In_2207);
nand U569 (N_569,In_2243,In_861);
xor U570 (N_570,In_4162,In_538);
nor U571 (N_571,In_2583,In_4783);
and U572 (N_572,In_3004,In_2416);
xnor U573 (N_573,In_1724,In_3782);
and U574 (N_574,In_1186,In_21);
and U575 (N_575,In_4218,In_3996);
or U576 (N_576,In_4577,In_4258);
and U577 (N_577,In_1358,In_563);
nand U578 (N_578,In_531,In_2389);
nand U579 (N_579,In_369,In_4943);
xor U580 (N_580,In_2368,In_353);
nand U581 (N_581,In_1514,In_2146);
nor U582 (N_582,In_938,In_2993);
nand U583 (N_583,In_608,In_4711);
or U584 (N_584,In_4681,In_1004);
and U585 (N_585,In_2127,In_3346);
or U586 (N_586,In_2249,In_3144);
nor U587 (N_587,In_801,In_3155);
xnor U588 (N_588,In_1177,In_3370);
nor U589 (N_589,In_889,In_3309);
xor U590 (N_590,In_2317,In_4598);
xnor U591 (N_591,In_3838,In_1618);
nand U592 (N_592,In_4445,In_1978);
nand U593 (N_593,In_3114,In_3886);
xor U594 (N_594,In_985,In_4777);
nor U595 (N_595,In_2899,In_1723);
or U596 (N_596,In_2754,In_111);
nand U597 (N_597,In_2603,In_753);
nand U598 (N_598,In_3300,In_4909);
nand U599 (N_599,In_888,In_4267);
and U600 (N_600,In_1911,In_1400);
and U601 (N_601,In_2996,In_3235);
nand U602 (N_602,In_4635,In_1735);
xor U603 (N_603,In_1390,In_1661);
nor U604 (N_604,In_433,In_1213);
nor U605 (N_605,In_101,In_2901);
and U606 (N_606,In_1357,In_2790);
xor U607 (N_607,In_4862,In_4666);
and U608 (N_608,In_4865,In_1715);
xnor U609 (N_609,In_3448,In_3463);
xor U610 (N_610,In_4561,In_1913);
or U611 (N_611,In_3940,In_866);
nor U612 (N_612,In_1563,In_545);
nor U613 (N_613,In_3912,In_4466);
and U614 (N_614,In_2631,In_1556);
and U615 (N_615,In_3364,In_964);
xnor U616 (N_616,In_1047,In_3499);
nand U617 (N_617,In_1547,In_587);
xnor U618 (N_618,In_998,In_4602);
and U619 (N_619,In_2162,In_2108);
nor U620 (N_620,In_2954,In_1896);
xor U621 (N_621,In_883,In_3009);
nand U622 (N_622,In_914,In_3458);
or U623 (N_623,In_565,In_2682);
nand U624 (N_624,In_3938,In_857);
and U625 (N_625,In_1751,In_4640);
nand U626 (N_626,In_402,In_4452);
nor U627 (N_627,In_130,In_1863);
or U628 (N_628,In_2579,In_4829);
and U629 (N_629,In_535,In_35);
nand U630 (N_630,In_192,In_1906);
xnor U631 (N_631,In_1055,In_1286);
nor U632 (N_632,In_269,In_174);
or U633 (N_633,In_968,In_3575);
xor U634 (N_634,In_3952,In_2041);
nor U635 (N_635,In_1603,In_2987);
nor U636 (N_636,In_2008,In_3289);
nand U637 (N_637,In_2439,In_4570);
nor U638 (N_638,In_4573,In_1842);
and U639 (N_639,In_4213,In_23);
and U640 (N_640,In_1760,In_2671);
xor U641 (N_641,In_2031,In_293);
and U642 (N_642,In_279,In_3140);
or U643 (N_643,In_4946,In_444);
xnor U644 (N_644,In_3647,In_3802);
nand U645 (N_645,In_2840,In_2406);
or U646 (N_646,In_2984,In_907);
nor U647 (N_647,In_3473,In_1783);
nor U648 (N_648,In_605,In_3044);
nand U649 (N_649,In_3305,In_3142);
xor U650 (N_650,In_1609,In_1993);
and U651 (N_651,In_51,In_4148);
xor U652 (N_652,In_41,In_4030);
xnor U653 (N_653,In_2699,In_3890);
nor U654 (N_654,In_884,In_806);
and U655 (N_655,In_1184,In_754);
and U656 (N_656,In_1837,In_2657);
and U657 (N_657,In_3712,In_308);
xnor U658 (N_658,In_1519,In_1477);
nand U659 (N_659,In_4728,In_1946);
xor U660 (N_660,In_4269,In_3413);
nand U661 (N_661,In_584,In_3141);
and U662 (N_662,In_2740,In_1290);
nor U663 (N_663,In_2913,In_1129);
nor U664 (N_664,In_4013,In_4981);
and U665 (N_665,In_3378,In_819);
or U666 (N_666,In_3523,In_922);
or U667 (N_667,In_654,In_387);
or U668 (N_668,In_3686,In_4756);
nand U669 (N_669,In_2184,In_3504);
and U670 (N_670,In_3530,In_2812);
nand U671 (N_671,In_4215,In_3968);
nor U672 (N_672,In_1455,In_1475);
or U673 (N_673,In_46,In_4432);
nand U674 (N_674,In_28,In_1572);
or U675 (N_675,In_644,In_4526);
and U676 (N_676,In_3115,In_3614);
nor U677 (N_677,In_2381,In_4461);
xnor U678 (N_678,In_4673,In_1115);
xor U679 (N_679,In_3035,In_4506);
and U680 (N_680,In_4652,In_2526);
and U681 (N_681,In_4179,In_1632);
nand U682 (N_682,In_597,In_4057);
nand U683 (N_683,In_4197,In_3367);
xor U684 (N_684,In_3957,In_4396);
xnor U685 (N_685,In_936,In_1807);
xnor U686 (N_686,In_4407,In_1313);
and U687 (N_687,In_3972,In_459);
xnor U688 (N_688,In_3292,In_366);
nand U689 (N_689,In_4411,In_4782);
and U690 (N_690,In_3931,In_813);
and U691 (N_691,In_4512,In_3810);
nor U692 (N_692,In_4235,In_2859);
and U693 (N_693,In_3913,In_432);
and U694 (N_694,In_3436,In_684);
and U695 (N_695,In_3595,In_3921);
nor U696 (N_696,In_3919,In_2139);
nand U697 (N_697,In_4118,In_2611);
xor U698 (N_698,In_32,In_378);
or U699 (N_699,In_978,In_2476);
and U700 (N_700,In_517,In_1599);
and U701 (N_701,In_2714,In_4985);
and U702 (N_702,In_1298,In_3272);
nor U703 (N_703,In_66,In_795);
nand U704 (N_704,In_2339,In_339);
nor U705 (N_705,In_3479,In_92);
nor U706 (N_706,In_4667,In_956);
xnor U707 (N_707,In_4107,In_3719);
nand U708 (N_708,In_2973,In_1419);
or U709 (N_709,In_660,In_4660);
or U710 (N_710,In_3455,In_2598);
nor U711 (N_711,In_2551,In_2621);
nor U712 (N_712,In_1487,In_3609);
nand U713 (N_713,In_3684,In_4533);
nor U714 (N_714,In_4035,In_1031);
xnor U715 (N_715,In_4720,In_3757);
nor U716 (N_716,In_2535,In_3528);
xor U717 (N_717,In_2729,In_4337);
nor U718 (N_718,In_1325,In_4625);
nand U719 (N_719,In_1740,In_4854);
and U720 (N_720,In_3431,In_2793);
and U721 (N_721,In_823,In_3173);
and U722 (N_722,In_2653,In_4292);
nand U723 (N_723,In_1296,In_1099);
nor U724 (N_724,In_2111,In_1503);
nor U725 (N_725,In_1796,In_3214);
or U726 (N_726,In_3599,In_1123);
nand U727 (N_727,In_4289,In_3776);
and U728 (N_728,In_132,In_2245);
nand U729 (N_729,In_2705,In_4167);
nor U730 (N_730,In_2231,In_1585);
xor U731 (N_731,In_4088,In_129);
xnor U732 (N_732,In_4849,In_3989);
nand U733 (N_733,In_239,In_1413);
nand U734 (N_734,In_4684,In_221);
nor U735 (N_735,In_2309,In_1792);
nor U736 (N_736,In_3579,In_4188);
and U737 (N_737,In_4338,In_485);
or U738 (N_738,In_2944,In_3211);
and U739 (N_739,In_3074,In_1464);
nand U740 (N_740,In_1742,In_1575);
nand U741 (N_741,In_3823,In_2520);
nand U742 (N_742,In_2156,In_3);
xor U743 (N_743,In_3321,In_2386);
and U744 (N_744,In_3794,In_2939);
or U745 (N_745,In_4855,In_2410);
nand U746 (N_746,In_643,In_136);
and U747 (N_747,In_2781,In_1157);
nand U748 (N_748,In_476,In_2190);
or U749 (N_749,In_1363,In_2103);
nor U750 (N_750,In_4210,In_1060);
and U751 (N_751,In_4073,In_2495);
or U752 (N_752,In_763,In_219);
or U753 (N_753,In_1354,In_2263);
nand U754 (N_754,In_4979,In_1527);
or U755 (N_755,In_1928,In_4810);
xnor U756 (N_756,In_3478,In_2575);
nor U757 (N_757,In_2470,In_2272);
xnor U758 (N_758,In_856,In_3301);
nand U759 (N_759,In_4416,In_1729);
and U760 (N_760,In_3622,In_2165);
and U761 (N_761,In_558,In_2260);
or U762 (N_762,In_3832,In_1531);
nand U763 (N_763,In_2233,In_2201);
or U764 (N_764,In_4654,In_1494);
nor U765 (N_765,In_782,In_3241);
and U766 (N_766,In_4679,In_4024);
nor U767 (N_767,In_2968,In_1447);
xnor U768 (N_768,In_2433,In_1147);
nor U769 (N_769,In_3594,In_4462);
xnor U770 (N_770,In_4170,In_3227);
or U771 (N_771,In_123,In_1710);
and U772 (N_772,In_261,In_390);
xnor U773 (N_773,In_4376,In_3178);
nor U774 (N_774,In_2950,In_2236);
xor U775 (N_775,In_709,In_3578);
nand U776 (N_776,In_2278,In_1168);
or U777 (N_777,In_2039,In_3958);
nor U778 (N_778,In_3524,In_1968);
xnor U779 (N_779,In_4704,In_340);
or U780 (N_780,In_1263,In_723);
or U781 (N_781,In_1683,In_2145);
and U782 (N_782,In_4284,In_3981);
and U783 (N_783,In_331,In_616);
and U784 (N_784,In_350,In_3617);
and U785 (N_785,In_4,In_4694);
xnor U786 (N_786,In_1977,In_2709);
and U787 (N_787,In_4571,In_2354);
nor U788 (N_788,In_2474,In_2441);
nand U789 (N_789,In_4967,In_3541);
xor U790 (N_790,In_4691,In_1866);
nand U791 (N_791,In_3844,In_2099);
xor U792 (N_792,In_336,In_154);
xnor U793 (N_793,In_2584,In_977);
nand U794 (N_794,In_2763,In_4730);
and U795 (N_795,In_2880,In_2591);
nand U796 (N_796,In_4121,In_3429);
xnor U797 (N_797,In_2776,In_2985);
xnor U798 (N_798,In_1330,In_4880);
xor U799 (N_799,In_3868,In_3192);
and U800 (N_800,In_2998,In_4548);
nand U801 (N_801,In_191,In_635);
and U802 (N_802,In_1247,In_1878);
nor U803 (N_803,In_4537,In_3911);
nand U804 (N_804,In_497,In_1223);
nor U805 (N_805,In_849,In_2811);
nand U806 (N_806,In_1128,In_4294);
nand U807 (N_807,In_3131,In_1016);
nor U808 (N_808,In_4633,In_1720);
nand U809 (N_809,In_1086,In_1417);
nand U810 (N_810,In_2937,In_646);
or U811 (N_811,In_3234,In_1009);
xnor U812 (N_812,In_72,In_2255);
or U813 (N_813,In_1989,In_1506);
nor U814 (N_814,In_4051,In_4659);
nand U815 (N_815,In_4523,In_4517);
or U816 (N_816,In_3251,In_3316);
and U817 (N_817,In_676,In_2558);
nand U818 (N_818,In_611,In_2071);
and U819 (N_819,In_872,In_4480);
nand U820 (N_820,In_1857,In_3539);
nand U821 (N_821,In_1523,In_1916);
nand U822 (N_822,In_3203,In_512);
and U823 (N_823,In_4017,In_375);
xnor U824 (N_824,In_4665,In_1346);
xor U825 (N_825,In_4904,In_4623);
and U826 (N_826,In_207,In_4986);
and U827 (N_827,In_1737,In_4525);
nor U828 (N_828,In_2347,In_1813);
xnor U829 (N_829,In_30,In_2837);
and U830 (N_830,In_2510,In_855);
nand U831 (N_831,In_3634,In_3331);
or U832 (N_832,In_4869,In_4921);
or U833 (N_833,In_1424,In_3982);
and U834 (N_834,In_4905,In_3027);
and U835 (N_835,In_3271,In_1535);
nand U836 (N_836,In_3282,In_493);
xor U837 (N_837,In_2608,In_2820);
nand U838 (N_838,In_4373,In_994);
nor U839 (N_839,In_623,In_636);
or U840 (N_840,In_3356,In_4145);
nand U841 (N_841,In_650,In_4655);
or U842 (N_842,In_4450,In_2098);
nand U843 (N_843,In_1516,In_1537);
nand U844 (N_844,In_3867,In_607);
nand U845 (N_845,In_3492,In_4645);
nand U846 (N_846,In_2980,In_58);
nor U847 (N_847,In_391,In_3785);
nor U848 (N_848,In_1418,In_3706);
or U849 (N_849,In_710,In_1002);
nor U850 (N_850,In_523,In_2425);
or U851 (N_851,In_3503,In_1960);
nand U852 (N_852,In_3915,In_3700);
xor U853 (N_853,In_954,In_2442);
nor U854 (N_854,In_2273,In_97);
nor U855 (N_855,In_3001,In_1425);
and U856 (N_856,In_2719,In_3897);
xnor U857 (N_857,In_3693,In_3347);
nand U858 (N_858,In_2227,In_3571);
or U859 (N_859,In_2457,In_4875);
and U860 (N_860,In_4779,In_2195);
nand U861 (N_861,In_4400,In_440);
or U862 (N_862,In_1821,In_3849);
and U863 (N_863,In_1040,In_4575);
nor U864 (N_864,In_4257,In_921);
nor U865 (N_865,In_1384,In_1108);
nand U866 (N_866,In_1367,In_1132);
nor U867 (N_867,In_3358,In_3992);
nand U868 (N_868,In_3848,In_2632);
xor U869 (N_869,In_2311,In_4155);
nor U870 (N_870,In_3060,In_4070);
xor U871 (N_871,In_109,In_3032);
nor U872 (N_872,In_1326,In_980);
and U873 (N_873,In_1453,In_2625);
nand U874 (N_874,In_2952,In_900);
nor U875 (N_875,In_1940,In_1790);
or U876 (N_876,In_1024,In_4934);
nor U877 (N_877,In_428,In_1870);
or U878 (N_878,In_3287,In_1394);
and U879 (N_879,In_4232,In_3885);
and U880 (N_880,In_1379,In_4113);
nor U881 (N_881,In_4980,In_384);
or U882 (N_882,In_995,In_335);
or U883 (N_883,In_913,In_1333);
nand U884 (N_884,In_556,In_4590);
nor U885 (N_885,In_1990,In_4358);
or U886 (N_886,In_2765,In_1759);
or U887 (N_887,In_4604,In_4716);
xor U888 (N_888,In_4275,In_3279);
or U889 (N_889,In_4699,In_2059);
xnor U890 (N_890,In_1847,In_4955);
xor U891 (N_891,In_1003,In_3433);
nand U892 (N_892,In_4527,In_4805);
nor U893 (N_893,In_3091,In_3888);
nor U894 (N_894,In_4836,In_2343);
and U895 (N_895,In_4762,In_4522);
xnor U896 (N_896,In_2589,In_2147);
or U897 (N_897,In_688,In_2513);
or U898 (N_898,In_2026,In_4770);
or U899 (N_899,In_3677,In_2411);
nor U900 (N_900,In_1376,In_4748);
xor U901 (N_901,In_882,In_4156);
or U902 (N_902,In_4301,In_4882);
nand U903 (N_903,In_3591,In_596);
nor U904 (N_904,In_4310,In_962);
nand U905 (N_905,In_2369,In_3661);
nor U906 (N_906,In_2494,In_957);
nand U907 (N_907,In_88,In_1169);
nand U908 (N_908,In_2382,In_3876);
nand U909 (N_909,In_814,In_48);
nor U910 (N_910,In_4647,In_3366);
and U911 (N_911,In_4992,In_1306);
or U912 (N_912,In_2349,In_3690);
nor U913 (N_913,In_1404,In_2017);
xnor U914 (N_914,In_4995,In_2907);
nand U915 (N_915,In_4205,In_3544);
or U916 (N_916,In_4222,In_2666);
and U917 (N_917,In_168,In_2659);
xor U918 (N_918,In_1996,In_2124);
nand U919 (N_919,In_4014,In_3307);
nor U920 (N_920,In_1582,In_397);
or U921 (N_921,In_996,In_1348);
nand U922 (N_922,In_4557,In_2908);
or U923 (N_923,In_1730,In_2046);
and U924 (N_924,In_178,In_3036);
nand U925 (N_925,In_4419,In_2738);
and U926 (N_926,In_1680,In_829);
nor U927 (N_927,In_1544,In_1139);
xor U928 (N_928,In_3963,In_4926);
xor U929 (N_929,In_598,In_4116);
xnor U930 (N_930,In_2841,In_126);
xnor U931 (N_931,In_443,In_4989);
xnor U932 (N_932,In_2620,In_2078);
nand U933 (N_933,In_4562,In_67);
xnor U934 (N_934,In_1888,In_3457);
xor U935 (N_935,In_4501,In_2553);
nor U936 (N_936,In_1900,In_4912);
or U937 (N_937,In_4817,In_3180);
nand U938 (N_938,In_582,In_4101);
xnor U939 (N_939,In_4738,In_1897);
nor U940 (N_940,In_639,In_161);
nor U941 (N_941,In_4363,In_3859);
nor U942 (N_942,In_3415,In_3633);
nand U943 (N_943,In_1638,In_173);
nand U944 (N_944,In_76,In_2722);
xnor U945 (N_945,In_1613,In_3553);
or U946 (N_946,In_581,In_481);
xnor U947 (N_947,In_1789,In_645);
or U948 (N_948,In_4638,In_1226);
and U949 (N_949,In_57,In_1707);
xnor U950 (N_950,In_1657,In_275);
and U951 (N_951,In_4983,In_3895);
nor U952 (N_952,In_43,In_4226);
and U953 (N_953,In_2397,In_3230);
xnor U954 (N_954,In_3820,In_3006);
nor U955 (N_955,In_425,In_4558);
or U956 (N_956,In_2393,In_295);
and U957 (N_957,In_796,In_1794);
nor U958 (N_958,In_4606,In_707);
xnor U959 (N_959,In_1639,In_4308);
nor U960 (N_960,In_1103,In_2891);
and U961 (N_961,In_4393,In_1834);
and U962 (N_962,In_4290,In_689);
and U963 (N_963,In_1191,In_3188);
or U964 (N_964,In_4765,In_2955);
nand U965 (N_965,In_4248,In_2561);
nor U966 (N_966,In_156,In_1208);
nor U967 (N_967,In_4872,In_4027);
nand U968 (N_968,In_987,In_3624);
and U969 (N_969,In_3043,In_902);
or U970 (N_970,In_1852,In_228);
nand U971 (N_971,In_3676,In_4803);
and U972 (N_972,In_890,In_1844);
nor U973 (N_973,In_3082,In_251);
or U974 (N_974,In_479,In_3111);
nor U975 (N_975,In_3749,In_755);
and U976 (N_976,In_1397,In_3548);
xor U977 (N_977,In_95,In_1473);
and U978 (N_978,In_4874,In_4916);
nand U979 (N_979,In_1278,In_1244);
xor U980 (N_980,In_1520,In_1032);
nand U981 (N_981,In_4605,In_424);
nor U982 (N_982,In_2737,In_4680);
nor U983 (N_983,In_2148,In_3809);
xnor U984 (N_984,In_2161,In_4936);
or U985 (N_985,In_887,In_455);
xor U986 (N_986,In_3285,In_1309);
nor U987 (N_987,In_2413,In_3207);
or U988 (N_988,In_4394,In_892);
nand U989 (N_989,In_1328,In_1285);
and U990 (N_990,In_4566,In_2650);
nand U991 (N_991,In_3497,In_2708);
nand U992 (N_992,In_423,In_4682);
and U993 (N_993,In_2037,In_4065);
nor U994 (N_994,In_152,In_3083);
xnor U995 (N_995,In_1221,In_4785);
xnor U996 (N_996,In_1033,In_933);
nor U997 (N_997,In_1081,In_2261);
nand U998 (N_998,In_304,In_2516);
and U999 (N_999,In_4371,In_321);
and U1000 (N_1000,In_2223,In_3124);
or U1001 (N_1001,In_4006,In_4502);
or U1002 (N_1002,In_105,In_4334);
nor U1003 (N_1003,In_3122,In_4962);
or U1004 (N_1004,In_2061,In_2892);
xnor U1005 (N_1005,In_663,In_1035);
and U1006 (N_1006,In_1633,In_1736);
or U1007 (N_1007,In_949,In_1066);
nor U1008 (N_1008,In_3979,In_1578);
xor U1009 (N_1009,In_2822,In_383);
xnor U1010 (N_1010,In_1833,In_4154);
and U1011 (N_1011,In_4620,In_2711);
xor U1012 (N_1012,In_1861,In_2066);
nor U1013 (N_1013,In_4000,In_1140);
nor U1014 (N_1014,In_4172,In_4381);
xor U1015 (N_1015,In_1261,In_233);
and U1016 (N_1016,In_3508,In_1387);
nor U1017 (N_1017,In_1964,In_334);
xnor U1018 (N_1018,In_993,In_1491);
nand U1019 (N_1019,In_1719,In_3329);
nor U1020 (N_1020,In_984,In_1052);
nor U1021 (N_1021,In_415,In_1521);
xor U1022 (N_1022,In_172,In_64);
nor U1023 (N_1023,In_3017,In_827);
nand U1024 (N_1024,In_3620,In_2619);
or U1025 (N_1025,In_2056,In_4599);
and U1026 (N_1026,In_897,In_1080);
and U1027 (N_1027,In_2137,In_4761);
nand U1028 (N_1028,In_2376,In_193);
nand U1029 (N_1029,In_148,In_2143);
and U1030 (N_1030,In_785,In_2772);
xor U1031 (N_1031,In_4545,In_4388);
nand U1032 (N_1032,In_4797,In_2721);
nand U1033 (N_1033,In_4161,In_3291);
or U1034 (N_1034,In_2690,In_3400);
xor U1035 (N_1035,In_469,In_975);
nor U1036 (N_1036,In_3350,In_4193);
and U1037 (N_1037,In_365,In_3593);
xnor U1038 (N_1038,In_3643,In_1294);
and U1039 (N_1039,In_4326,In_3402);
nand U1040 (N_1040,In_175,In_3016);
or U1041 (N_1041,In_170,In_2300);
and U1042 (N_1042,In_1864,In_3117);
xnor U1043 (N_1043,In_1626,In_65);
xnor U1044 (N_1044,In_3159,In_1167);
nor U1045 (N_1045,In_4286,In_2597);
nand U1046 (N_1046,In_1145,In_3930);
xor U1047 (N_1047,In_171,In_1932);
and U1048 (N_1048,In_3572,In_3908);
or U1049 (N_1049,In_4884,In_3602);
and U1050 (N_1050,In_2402,In_4847);
nand U1051 (N_1051,In_3333,In_1997);
or U1052 (N_1052,In_4853,In_4596);
and U1053 (N_1053,In_1293,In_107);
and U1054 (N_1054,In_559,In_3318);
nand U1055 (N_1055,In_3129,In_3228);
nand U1056 (N_1056,In_1444,In_4858);
or U1057 (N_1057,In_1258,In_3196);
xor U1058 (N_1058,In_478,In_2914);
or U1059 (N_1059,In_206,In_1289);
and U1060 (N_1060,In_2835,In_1270);
nand U1061 (N_1061,In_4463,In_4932);
xor U1062 (N_1062,In_1687,In_1987);
or U1063 (N_1063,In_543,In_4142);
xor U1064 (N_1064,In_3411,In_1505);
nor U1065 (N_1065,In_4707,In_3467);
nor U1066 (N_1066,In_3825,In_2030);
nand U1067 (N_1067,In_4634,In_2808);
or U1068 (N_1068,In_2453,In_4153);
and U1069 (N_1069,In_726,In_2966);
and U1070 (N_1070,In_1340,In_4987);
nand U1071 (N_1071,In_4390,In_1830);
nand U1072 (N_1072,In_2713,In_184);
nor U1073 (N_1073,In_4468,In_1698);
and U1074 (N_1074,In_1440,In_1619);
nand U1075 (N_1075,In_333,In_1756);
nor U1076 (N_1076,In_4094,In_4614);
xor U1077 (N_1077,In_1973,In_2437);
nand U1078 (N_1078,In_270,In_683);
nor U1079 (N_1079,In_1364,In_944);
nor U1080 (N_1080,In_1942,In_3355);
xnor U1081 (N_1081,In_2819,In_3220);
nor U1082 (N_1082,In_1368,In_3557);
nor U1083 (N_1083,In_2716,In_4317);
xnor U1084 (N_1084,In_342,In_1194);
and U1085 (N_1085,In_3828,In_4398);
nor U1086 (N_1086,In_3094,In_1608);
xnor U1087 (N_1087,In_2215,In_3481);
and U1088 (N_1088,In_983,In_2387);
nor U1089 (N_1089,In_1647,In_4742);
xor U1090 (N_1090,In_3875,In_4842);
xnor U1091 (N_1091,In_743,In_2874);
or U1092 (N_1092,In_3369,In_2093);
or U1093 (N_1093,In_2975,In_773);
nor U1094 (N_1094,In_4686,In_4773);
or U1095 (N_1095,In_3991,In_2999);
and U1096 (N_1096,In_2324,In_591);
or U1097 (N_1097,In_3817,In_1579);
nor U1098 (N_1098,In_166,In_1975);
and U1099 (N_1099,In_2029,In_792);
and U1100 (N_1100,In_3896,In_2428);
nand U1101 (N_1101,In_4045,In_4339);
xor U1102 (N_1102,In_873,In_1738);
nor U1103 (N_1103,In_180,In_3237);
nand U1104 (N_1104,In_911,In_2672);
xnor U1105 (N_1105,In_2268,In_991);
nor U1106 (N_1106,In_1895,In_1071);
nand U1107 (N_1107,In_1101,In_362);
and U1108 (N_1108,In_4894,In_3158);
nand U1109 (N_1109,In_4042,In_2730);
xnor U1110 (N_1110,In_212,In_2151);
nand U1111 (N_1111,In_2210,In_1814);
xnor U1112 (N_1112,In_4800,In_2083);
or U1113 (N_1113,In_3659,In_4110);
and U1114 (N_1114,In_1229,In_1560);
or U1115 (N_1115,In_2306,In_3250);
xnor U1116 (N_1116,In_3422,In_4538);
nor U1117 (N_1117,In_844,In_1526);
or U1118 (N_1118,In_1908,In_4058);
and U1119 (N_1119,In_4807,In_3465);
xor U1120 (N_1120,In_1658,In_613);
nor U1121 (N_1121,In_2942,In_3049);
nand U1122 (N_1122,In_971,In_4721);
nor U1123 (N_1123,In_4601,In_3439);
xor U1124 (N_1124,In_4610,In_2670);
or U1125 (N_1125,In_1791,In_915);
and U1126 (N_1126,In_1757,In_2725);
xnor U1127 (N_1127,In_301,In_93);
or U1128 (N_1128,In_3542,In_1264);
nand U1129 (N_1129,In_4670,In_2119);
or U1130 (N_1130,In_2926,In_4723);
nor U1131 (N_1131,In_4470,In_2036);
nor U1132 (N_1132,In_1664,In_1155);
and U1133 (N_1133,In_4090,In_4961);
xnor U1134 (N_1134,In_243,In_1492);
xor U1135 (N_1135,In_1528,In_3388);
and U1136 (N_1136,In_4109,In_4383);
or U1137 (N_1137,In_1611,In_1077);
nand U1138 (N_1138,In_4221,In_3018);
nand U1139 (N_1139,In_332,In_594);
nor U1140 (N_1140,In_4546,In_3393);
or U1141 (N_1141,In_1862,In_4902);
nand U1142 (N_1142,In_2378,In_4238);
or U1143 (N_1143,In_4103,In_4152);
xnor U1144 (N_1144,In_4007,In_4774);
nand U1145 (N_1145,In_254,In_3090);
nor U1146 (N_1146,In_1912,In_3918);
xnor U1147 (N_1147,In_2000,In_3833);
nand U1148 (N_1148,In_2302,In_1877);
nand U1149 (N_1149,In_2791,In_4690);
nand U1150 (N_1150,In_2612,In_4039);
and U1151 (N_1151,In_1116,In_53);
xnor U1152 (N_1152,In_780,In_386);
nor U1153 (N_1153,In_3790,In_1232);
xor U1154 (N_1154,In_2866,In_3526);
and U1155 (N_1155,In_3003,In_513);
or U1156 (N_1156,In_2331,In_1644);
nor U1157 (N_1157,In_3041,In_1799);
or U1158 (N_1158,In_549,In_4746);
nor U1159 (N_1159,In_4893,In_590);
nor U1160 (N_1160,In_633,In_3322);
or U1161 (N_1161,In_1782,In_3474);
or U1162 (N_1162,In_1853,In_508);
xor U1163 (N_1163,In_2517,In_4937);
and U1164 (N_1164,In_457,In_1894);
nand U1165 (N_1165,In_2938,In_4784);
nand U1166 (N_1166,In_3977,In_1174);
nor U1167 (N_1167,In_2379,In_3126);
xnor U1168 (N_1168,In_1780,In_560);
xnor U1169 (N_1169,In_20,In_1339);
nand U1170 (N_1170,In_215,In_4702);
or U1171 (N_1171,In_1557,In_4433);
nor U1172 (N_1172,In_2602,In_832);
or U1173 (N_1173,In_1648,In_934);
nor U1174 (N_1174,In_395,In_3310);
and U1175 (N_1175,In_90,In_2766);
and U1176 (N_1176,In_1630,In_2408);
nand U1177 (N_1177,In_2062,In_149);
and U1178 (N_1178,In_2136,In_3680);
nand U1179 (N_1179,In_4249,In_3315);
or U1180 (N_1180,In_2974,In_2075);
nor U1181 (N_1181,In_3748,In_2067);
xor U1182 (N_1182,In_965,In_3939);
xnor U1183 (N_1183,In_1642,In_1651);
and U1184 (N_1184,In_2068,In_417);
or U1185 (N_1185,In_4734,In_4487);
nand U1186 (N_1186,In_3337,In_128);
and U1187 (N_1187,In_1776,In_1472);
or U1188 (N_1188,In_2218,In_1429);
nand U1189 (N_1189,In_2003,In_1754);
nand U1190 (N_1190,In_2496,In_1409);
xor U1191 (N_1191,In_4263,In_1601);
or U1192 (N_1192,In_675,In_4319);
nor U1193 (N_1193,In_189,In_1255);
nor U1194 (N_1194,In_700,In_1266);
and U1195 (N_1195,In_4378,In_1329);
or U1196 (N_1196,In_2783,In_3894);
and U1197 (N_1197,In_4583,In_579);
or U1198 (N_1198,In_542,In_850);
or U1199 (N_1199,In_657,In_229);
xor U1200 (N_1200,In_246,In_1470);
and U1201 (N_1201,In_281,In_1515);
xnor U1202 (N_1202,In_865,In_1439);
and U1203 (N_1203,In_4973,In_3846);
xnor U1204 (N_1204,In_1056,In_1317);
or U1205 (N_1205,In_555,In_104);
and U1206 (N_1206,In_2128,In_3718);
xnor U1207 (N_1207,In_2254,In_2133);
and U1208 (N_1208,In_2910,In_739);
xor U1209 (N_1209,In_4099,In_719);
nand U1210 (N_1210,In_323,In_2947);
or U1211 (N_1211,In_4305,In_2511);
xor U1212 (N_1212,In_238,In_903);
xor U1213 (N_1213,In_86,In_3198);
nand U1214 (N_1214,In_2757,In_3827);
nand U1215 (N_1215,In_414,In_1391);
nor U1216 (N_1216,In_4900,In_536);
nor U1217 (N_1217,In_3775,In_74);
xor U1218 (N_1218,In_2117,In_2925);
and U1219 (N_1219,In_1204,In_3449);
nand U1220 (N_1220,In_2919,In_385);
and U1221 (N_1221,In_3000,In_1192);
nor U1222 (N_1222,In_1399,In_2515);
nand U1223 (N_1223,In_2897,In_1466);
nand U1224 (N_1224,In_717,In_4386);
nor U1225 (N_1225,In_3720,In_4104);
or U1226 (N_1226,In_54,In_3238);
xnor U1227 (N_1227,In_1320,In_29);
nor U1228 (N_1228,In_570,In_3889);
nor U1229 (N_1229,In_3694,In_1787);
nand U1230 (N_1230,In_1268,In_1543);
nand U1231 (N_1231,In_1336,In_833);
nor U1232 (N_1232,In_2768,In_752);
or U1233 (N_1233,In_94,In_2450);
or U1234 (N_1234,In_4543,In_1949);
xnor U1235 (N_1235,In_4458,In_2744);
nor U1236 (N_1236,In_1434,In_2323);
xor U1237 (N_1237,In_1323,In_3002);
nand U1238 (N_1238,In_4236,In_3953);
nand U1239 (N_1239,In_3226,In_3650);
or U1240 (N_1240,In_1706,In_1022);
or U1241 (N_1241,In_1025,In_1565);
nor U1242 (N_1242,In_484,In_1019);
and U1243 (N_1243,In_1190,In_925);
and U1244 (N_1244,In_1316,In_3382);
and U1245 (N_1245,In_1120,In_1612);
or U1246 (N_1246,In_4553,In_3215);
and U1247 (N_1247,In_3853,In_2787);
xnor U1248 (N_1248,In_2635,In_4948);
and U1249 (N_1249,In_2654,In_1421);
and U1250 (N_1250,In_820,In_1044);
or U1251 (N_1251,In_2641,In_4442);
nand U1252 (N_1252,In_810,In_4843);
nand U1253 (N_1253,In_3653,In_2284);
nand U1254 (N_1254,In_4174,In_3266);
nand U1255 (N_1255,In_3688,In_2487);
nor U1256 (N_1256,In_4089,In_4040);
nand U1257 (N_1257,In_1474,In_1892);
xor U1258 (N_1258,In_4138,In_4629);
xnor U1259 (N_1259,In_2109,In_2660);
xnor U1260 (N_1260,In_4619,In_2800);
or U1261 (N_1261,In_3302,In_3969);
nand U1262 (N_1262,In_3088,In_4066);
and U1263 (N_1263,In_2622,In_1999);
and U1264 (N_1264,In_4341,In_3095);
or U1265 (N_1265,In_2417,In_2651);
or U1266 (N_1266,In_3354,In_1645);
nor U1267 (N_1267,In_2044,In_3878);
xor U1268 (N_1268,In_3961,In_1764);
and U1269 (N_1269,In_2664,In_2826);
xor U1270 (N_1270,In_708,In_3314);
nor U1271 (N_1271,In_3270,In_3673);
and U1272 (N_1272,In_14,In_853);
and U1273 (N_1273,In_4957,In_2810);
and U1274 (N_1274,In_1772,In_1570);
nand U1275 (N_1275,In_3295,In_794);
nor U1276 (N_1276,In_3119,In_4806);
xnor U1277 (N_1277,In_1322,In_2991);
nand U1278 (N_1278,In_1353,In_3531);
nand U1279 (N_1279,In_877,In_4661);
nand U1280 (N_1280,In_4725,In_1146);
nor U1281 (N_1281,In_1459,In_272);
nand U1282 (N_1282,In_2132,In_4824);
nand U1283 (N_1283,In_2893,In_3954);
or U1284 (N_1284,In_3087,In_138);
and U1285 (N_1285,In_3937,In_3691);
or U1286 (N_1286,In_3877,In_3038);
nand U1287 (N_1287,In_2497,In_4246);
nand U1288 (N_1288,In_3640,In_2786);
nor U1289 (N_1289,In_2629,In_2663);
nor U1290 (N_1290,In_1769,In_3767);
or U1291 (N_1291,In_2505,In_837);
and U1292 (N_1292,In_3089,In_4186);
nand U1293 (N_1293,In_100,In_290);
xor U1294 (N_1294,In_4769,In_1302);
nor U1295 (N_1295,In_3063,In_3851);
or U1296 (N_1296,In_1674,In_4331);
nor U1297 (N_1297,In_3404,In_1731);
nor U1298 (N_1298,In_638,In_2206);
nand U1299 (N_1299,In_3628,In_1704);
or U1300 (N_1300,In_1758,In_3754);
nand U1301 (N_1301,In_731,In_2856);
nor U1302 (N_1302,In_1124,In_483);
or U1303 (N_1303,In_3189,In_783);
nand U1304 (N_1304,In_3075,In_3569);
xor U1305 (N_1305,In_772,In_1761);
or U1306 (N_1306,In_768,In_165);
nand U1307 (N_1307,In_3288,In_2345);
nor U1308 (N_1308,In_2022,In_1546);
xor U1309 (N_1309,In_1038,In_234);
nor U1310 (N_1310,In_950,In_2581);
nand U1311 (N_1311,In_1835,In_3319);
and U1312 (N_1312,In_2885,In_298);
nor U1313 (N_1313,In_96,In_2900);
xor U1314 (N_1314,In_1291,In_237);
and U1315 (N_1315,In_3469,In_3583);
xnor U1316 (N_1316,In_845,In_3242);
and U1317 (N_1317,In_1804,In_4929);
and U1318 (N_1318,In_1875,In_1747);
xor U1319 (N_1319,In_102,In_2863);
nand U1320 (N_1320,In_412,In_1798);
and U1321 (N_1321,In_392,In_629);
nand U1322 (N_1322,In_5,In_2319);
and U1323 (N_1323,In_3443,In_1172);
and U1324 (N_1324,In_4851,In_78);
or U1325 (N_1325,In_1937,In_4234);
nand U1326 (N_1326,In_3170,In_4550);
and U1327 (N_1327,In_557,In_4354);
and U1328 (N_1328,In_287,In_4131);
nand U1329 (N_1329,In_3537,In_2295);
and U1330 (N_1330,In_1646,In_4140);
nor U1331 (N_1331,In_4285,In_4798);
or U1332 (N_1332,In_2443,In_4387);
xnor U1333 (N_1333,In_2130,In_368);
xnor U1334 (N_1334,In_4332,In_3927);
and U1335 (N_1335,In_3641,In_716);
nor U1336 (N_1336,In_98,In_4714);
and U1337 (N_1337,In_880,In_4441);
or U1338 (N_1338,In_1668,In_4384);
or U1339 (N_1339,In_572,In_17);
or U1340 (N_1340,In_2461,In_137);
nor U1341 (N_1341,In_4178,In_862);
xnor U1342 (N_1342,In_3202,In_1905);
or U1343 (N_1343,In_1722,In_1430);
or U1344 (N_1344,In_2552,In_634);
or U1345 (N_1345,In_3722,In_1460);
nor U1346 (N_1346,In_4731,In_2839);
nand U1347 (N_1347,In_4455,In_1370);
nand U1348 (N_1348,In_3376,In_1558);
nand U1349 (N_1349,In_2992,In_4726);
and U1350 (N_1350,In_2527,In_1051);
or U1351 (N_1351,In_2803,In_475);
or U1352 (N_1352,In_2016,In_4622);
nor U1353 (N_1353,In_1872,In_839);
xor U1354 (N_1354,In_3655,In_3120);
xor U1355 (N_1355,In_712,In_24);
nand U1356 (N_1356,In_1271,In_2356);
and U1357 (N_1357,In_4352,In_4034);
nor U1358 (N_1358,In_2414,In_1469);
nand U1359 (N_1359,In_3055,In_1659);
nor U1360 (N_1360,In_1288,In_656);
nor U1361 (N_1361,In_4567,In_4958);
nor U1362 (N_1362,In_1513,In_1576);
and U1363 (N_1363,In_45,In_2057);
nand U1364 (N_1364,In_4664,In_1739);
xnor U1365 (N_1365,In_1819,In_496);
or U1366 (N_1366,In_2424,In_2385);
or U1367 (N_1367,In_4771,In_389);
xnor U1368 (N_1368,In_1741,In_2884);
or U1369 (N_1369,In_4878,In_2290);
nor U1370 (N_1370,In_1381,In_3816);
nand U1371 (N_1371,In_3670,In_2838);
and U1372 (N_1372,In_4814,In_2498);
and U1373 (N_1373,In_648,In_4820);
nor U1374 (N_1374,In_4019,In_4542);
and U1375 (N_1375,In_303,In_540);
or U1376 (N_1376,In_706,In_4514);
xor U1377 (N_1377,In_3223,In_99);
xor U1378 (N_1378,In_4819,In_2734);
nand U1379 (N_1379,In_1265,In_435);
nand U1380 (N_1380,In_4631,In_1327);
or U1381 (N_1381,In_1377,In_2801);
nand U1382 (N_1382,In_3277,In_3656);
xnor U1383 (N_1383,In_3056,In_4541);
nand U1384 (N_1384,In_434,In_3236);
and U1385 (N_1385,In_2293,In_3856);
nor U1386 (N_1386,In_3510,In_112);
nand U1387 (N_1387,In_942,In_1567);
nor U1388 (N_1388,In_4312,In_804);
xor U1389 (N_1389,In_3987,In_2707);
or U1390 (N_1390,In_158,In_73);
nand U1391 (N_1391,In_2752,In_3909);
and U1392 (N_1392,In_4753,In_114);
xnor U1393 (N_1393,In_1827,In_379);
or U1394 (N_1394,In_142,In_4225);
nor U1395 (N_1395,In_401,In_2362);
nand U1396 (N_1396,In_3149,In_3651);
and U1397 (N_1397,In_2188,In_50);
xnor U1398 (N_1398,In_2086,In_1423);
or U1399 (N_1399,In_1234,In_2673);
or U1400 (N_1400,In_533,In_3362);
xnor U1401 (N_1401,In_1240,In_4500);
and U1402 (N_1402,In_249,In_4343);
nand U1403 (N_1403,In_2478,In_625);
xor U1404 (N_1404,In_418,In_4669);
nand U1405 (N_1405,In_951,In_188);
xor U1406 (N_1406,In_3774,In_4342);
nor U1407 (N_1407,In_2131,In_1100);
xnor U1408 (N_1408,In_2861,In_1770);
nand U1409 (N_1409,In_1592,In_4892);
xnor U1410 (N_1410,In_3330,In_3050);
nand U1411 (N_1411,In_658,In_3286);
and U1412 (N_1412,In_4891,In_3701);
nand U1413 (N_1413,In_2002,In_1868);
nor U1414 (N_1414,In_4863,In_2906);
xor U1415 (N_1415,In_1048,In_4998);
xnor U1416 (N_1416,In_4607,In_52);
nand U1417 (N_1417,In_1930,In_4465);
nand U1418 (N_1418,In_1283,In_1777);
xnor U1419 (N_1419,In_2751,In_211);
xor U1420 (N_1420,In_2459,In_451);
nor U1421 (N_1421,In_3771,In_695);
nor U1422 (N_1422,In_3375,In_441);
or U1423 (N_1423,In_3587,In_2865);
xor U1424 (N_1424,In_3654,In_4796);
or U1425 (N_1425,In_526,In_247);
xor U1426 (N_1426,In_2656,In_3154);
nor U1427 (N_1427,In_2304,In_3652);
and U1428 (N_1428,In_3359,In_926);
and U1429 (N_1429,In_1793,In_4780);
or U1430 (N_1430,In_999,In_961);
xnor U1431 (N_1431,In_2771,In_3102);
nor U1432 (N_1432,In_701,In_1497);
and U1433 (N_1433,In_179,In_2687);
nand U1434 (N_1434,In_1691,In_3994);
and U1435 (N_1435,In_3450,In_4511);
nand U1436 (N_1436,In_4764,In_4938);
xor U1437 (N_1437,In_1903,In_1305);
xnor U1438 (N_1438,In_2715,In_3403);
or U1439 (N_1439,In_4187,In_1595);
nand U1440 (N_1440,In_2782,In_2644);
and U1441 (N_1441,In_3464,In_2995);
and U1442 (N_1442,In_2055,In_3209);
or U1443 (N_1443,In_2875,In_1709);
nor U1444 (N_1444,In_196,In_1865);
nand U1445 (N_1445,In_315,In_2220);
nand U1446 (N_1446,In_4410,In_2287);
or U1447 (N_1447,In_1748,In_1721);
nor U1448 (N_1448,In_1279,In_1259);
or U1449 (N_1449,In_2959,In_1580);
and U1450 (N_1450,In_614,In_4259);
or U1451 (N_1451,In_673,In_1945);
nand U1452 (N_1452,In_3910,In_3345);
nor U1453 (N_1453,In_4025,In_898);
or U1454 (N_1454,In_183,In_1902);
and U1455 (N_1455,In_1665,In_2344);
nor U1456 (N_1456,In_1113,In_205);
xnor U1457 (N_1457,In_2432,In_4224);
nor U1458 (N_1458,In_2606,In_2544);
and U1459 (N_1459,In_1775,In_1884);
and U1460 (N_1460,In_218,In_2423);
xnor U1461 (N_1461,In_4600,In_2367);
xnor U1462 (N_1462,In_4692,In_3588);
or U1463 (N_1463,In_343,In_360);
xor U1464 (N_1464,In_1753,In_3900);
and U1465 (N_1465,In_2332,In_4933);
and U1466 (N_1466,In_3860,In_1530);
or U1467 (N_1467,In_4074,In_982);
xor U1468 (N_1468,In_436,In_4163);
xor U1469 (N_1469,In_600,In_1175);
and U1470 (N_1470,In_1649,In_1062);
xor U1471 (N_1471,In_1142,In_4508);
xor U1472 (N_1472,In_4069,In_4813);
xor U1473 (N_1473,In_1778,In_4251);
or U1474 (N_1474,In_4011,In_1749);
and U1475 (N_1475,In_2630,In_1924);
nand U1476 (N_1476,In_3024,In_1251);
or U1477 (N_1477,In_2945,In_2518);
nor U1478 (N_1478,In_734,In_3452);
nand U1479 (N_1479,In_4947,In_3097);
nor U1480 (N_1480,In_4794,In_778);
or U1481 (N_1481,In_4485,In_4540);
nand U1482 (N_1482,In_824,In_4924);
xnor U1483 (N_1483,In_3925,In_3039);
xnor U1484 (N_1484,In_1628,In_3995);
nand U1485 (N_1485,In_1445,In_200);
nand U1486 (N_1486,In_2904,In_2590);
or U1487 (N_1487,In_575,In_2623);
xnor U1488 (N_1488,In_3407,In_2463);
and U1489 (N_1489,In_1907,In_4302);
nor U1490 (N_1490,In_3135,In_1134);
and U1491 (N_1491,In_1917,In_2592);
xor U1492 (N_1492,In_199,In_3549);
nor U1493 (N_1493,In_4789,In_2228);
xnor U1494 (N_1494,In_3642,In_2694);
nand U1495 (N_1495,In_1001,In_3072);
and U1496 (N_1496,In_3268,In_4503);
and U1497 (N_1497,In_1933,In_164);
xor U1498 (N_1498,In_2986,In_703);
nand U1499 (N_1499,In_2401,In_2081);
nor U1500 (N_1500,In_208,In_534);
and U1501 (N_1501,In_2941,In_4521);
nor U1502 (N_1502,In_3760,In_4435);
nand U1503 (N_1503,In_507,In_2333);
nor U1504 (N_1504,In_3219,In_2601);
nor U1505 (N_1505,In_2226,In_1677);
nor U1506 (N_1506,In_4642,In_1065);
and U1507 (N_1507,In_3697,In_2609);
nand U1508 (N_1508,In_3902,In_1708);
and U1509 (N_1509,In_1805,In_411);
and U1510 (N_1510,In_2456,In_373);
xor U1511 (N_1511,In_1923,In_1159);
or U1512 (N_1512,In_2934,In_4472);
nor U1513 (N_1513,In_502,In_3459);
nand U1514 (N_1514,In_1401,In_3511);
and U1515 (N_1515,In_133,In_912);
and U1516 (N_1516,In_2960,In_9);
xnor U1517 (N_1517,In_1411,In_1188);
and U1518 (N_1518,In_3964,In_1590);
and U1519 (N_1519,In_4015,In_2753);
or U1520 (N_1520,In_4053,In_2182);
or U1521 (N_1521,In_4499,In_3563);
and U1522 (N_1522,In_2696,In_2087);
and U1523 (N_1523,In_1046,In_2308);
or U1524 (N_1524,In_2679,In_3758);
xor U1525 (N_1525,In_1484,In_931);
nand U1526 (N_1526,In_847,In_4585);
nand U1527 (N_1527,In_157,In_764);
nand U1528 (N_1528,In_3256,In_3186);
nand U1529 (N_1529,In_3361,In_3568);
nand U1530 (N_1530,In_1744,In_3513);
nor U1531 (N_1531,In_2012,In_748);
xor U1532 (N_1532,In_3880,In_1750);
nor U1533 (N_1533,In_3558,In_3033);
or U1534 (N_1534,In_2676,In_1970);
and U1535 (N_1535,In_4127,In_2577);
nor U1536 (N_1536,In_2747,In_283);
or U1537 (N_1537,In_124,In_3518);
and U1538 (N_1538,In_1957,In_945);
xor U1539 (N_1539,In_509,In_2639);
nor U1540 (N_1540,In_2556,In_1058);
nor U1541 (N_1541,In_989,In_1010);
and U1542 (N_1542,In_1552,In_2225);
or U1543 (N_1543,In_822,In_4615);
and U1544 (N_1544,In_3412,In_817);
nor U1545 (N_1545,In_4437,In_2686);
nor U1546 (N_1546,In_1448,In_2134);
or U1547 (N_1547,In_3125,In_36);
nor U1548 (N_1548,In_296,In_4194);
nor U1549 (N_1549,In_4108,In_337);
or U1550 (N_1550,In_3297,In_628);
nand U1551 (N_1551,In_3324,In_2238);
nand U1552 (N_1552,In_4309,In_1388);
nor U1553 (N_1553,In_4840,In_2007);
nand U1554 (N_1554,In_3887,In_2739);
xor U1555 (N_1555,In_2604,In_3093);
nor U1556 (N_1556,In_1319,In_1412);
nand U1557 (N_1557,In_3836,In_1669);
and U1558 (N_1558,In_56,In_2283);
and U1559 (N_1559,In_4038,In_2545);
nor U1560 (N_1560,In_1187,In_4656);
xnor U1561 (N_1561,In_4560,In_1254);
and U1562 (N_1562,In_3742,In_1498);
xor U1563 (N_1563,In_3231,In_225);
or U1564 (N_1564,In_4866,In_4389);
or U1565 (N_1565,In_3352,In_1227);
nor U1566 (N_1566,In_2836,In_274);
and U1567 (N_1567,In_3772,In_4003);
and U1568 (N_1568,In_4362,In_3705);
xnor U1569 (N_1569,In_3213,In_3983);
or U1570 (N_1570,In_2773,In_1104);
xor U1571 (N_1571,In_1006,In_3387);
xnor U1572 (N_1572,In_2129,In_2933);
and U1573 (N_1573,In_3883,In_960);
xor U1574 (N_1574,In_711,In_3798);
xor U1575 (N_1575,In_2454,In_3441);
nor U1576 (N_1576,In_2823,In_4778);
and U1577 (N_1577,In_1141,In_4061);
xor U1578 (N_1578,In_4974,In_4293);
and U1579 (N_1579,In_2429,In_2034);
xnor U1580 (N_1580,In_3818,In_77);
and U1581 (N_1581,In_2351,In_4582);
xor U1582 (N_1582,In_2600,In_2125);
and U1583 (N_1583,In_1441,In_3096);
and U1584 (N_1584,In_893,In_899);
nand U1585 (N_1585,In_2473,In_3618);
or U1586 (N_1586,In_1703,In_2712);
nor U1587 (N_1587,In_1382,In_2234);
or U1588 (N_1588,In_553,In_177);
nor U1589 (N_1589,In_4426,In_144);
or U1590 (N_1590,In_2888,In_2519);
nor U1591 (N_1591,In_4717,In_4479);
nand U1592 (N_1592,In_746,In_347);
xor U1593 (N_1593,In_4382,In_4250);
xnor U1594 (N_1594,In_3311,In_1511);
nor U1595 (N_1595,In_3716,In_3545);
and U1596 (N_1596,In_2528,In_923);
nor U1597 (N_1597,In_3766,In_4004);
xor U1598 (N_1598,In_2514,In_4718);
or U1599 (N_1599,In_685,In_3136);
or U1600 (N_1600,In_3424,In_1586);
nand U1601 (N_1601,In_3177,In_2170);
nand U1602 (N_1602,In_1816,In_2932);
and U1603 (N_1603,In_446,In_3804);
nand U1604 (N_1604,In_1180,In_44);
nand U1605 (N_1605,In_3841,In_3217);
and U1606 (N_1606,In_2979,In_3639);
xnor U1607 (N_1607,In_2187,In_514);
or U1608 (N_1608,In_244,In_4812);
nand U1609 (N_1609,In_1667,In_3725);
xor U1610 (N_1610,In_511,In_1995);
and U1611 (N_1611,In_1407,In_1389);
and U1612 (N_1612,In_4959,In_3536);
nand U1613 (N_1613,In_223,In_3784);
xor U1614 (N_1614,In_2276,In_2636);
xor U1615 (N_1615,In_42,In_197);
nor U1616 (N_1616,In_4530,In_520);
nor U1617 (N_1617,In_860,In_759);
or U1618 (N_1618,In_2391,In_277);
or U1619 (N_1619,In_3695,In_4335);
xnor U1620 (N_1620,In_4885,In_472);
nand U1621 (N_1621,In_1634,In_4430);
nor U1622 (N_1622,In_4555,In_2499);
or U1623 (N_1623,In_1956,In_870);
nor U1624 (N_1624,In_1812,In_3863);
nand U1625 (N_1625,In_599,In_2559);
or U1626 (N_1626,In_409,In_273);
or U1627 (N_1627,In_1561,In_2512);
or U1628 (N_1628,In_3872,In_1961);
xor U1629 (N_1629,In_1982,In_3751);
and U1630 (N_1630,In_3786,In_4584);
and U1631 (N_1631,In_2240,In_3105);
and U1632 (N_1632,In_2748,In_1673);
or U1633 (N_1633,In_2370,In_1551);
nor U1634 (N_1634,In_1078,In_894);
nand U1635 (N_1635,In_4653,In_4037);
nand U1636 (N_1636,In_1090,In_370);
or U1637 (N_1637,In_3428,In_3574);
and U1638 (N_1638,In_4613,In_1230);
and U1639 (N_1639,In_1137,In_4507);
nor U1640 (N_1640,In_2326,In_1806);
nand U1641 (N_1641,In_4190,In_3891);
nand U1642 (N_1642,In_2104,In_802);
and U1643 (N_1643,In_2981,In_4532);
nand U1644 (N_1644,In_3484,In_2259);
nor U1645 (N_1645,In_529,In_322);
or U1646 (N_1646,In_4056,In_2780);
xor U1647 (N_1647,In_1594,In_1117);
and U1648 (N_1648,In_248,In_2742);
or U1649 (N_1649,In_4189,In_2796);
and U1650 (N_1650,In_222,In_4278);
xnor U1651 (N_1651,In_3048,In_3085);
nor U1652 (N_1652,In_784,In_2196);
nand U1653 (N_1653,In_3516,In_2702);
or U1654 (N_1654,In_4212,In_405);
nand U1655 (N_1655,In_2646,In_4288);
nor U1656 (N_1656,In_680,In_720);
xor U1657 (N_1657,In_3681,In_2350);
xor U1658 (N_1658,In_2877,In_4950);
nand U1659 (N_1659,In_1650,In_2983);
xor U1660 (N_1660,In_828,In_1797);
and U1661 (N_1661,In_1587,In_3249);
xnor U1662 (N_1662,In_3879,In_2400);
nand U1663 (N_1663,In_2563,In_3137);
xnor U1664 (N_1664,In_1321,In_2258);
and U1665 (N_1665,In_4126,In_4379);
or U1666 (N_1666,In_3047,In_879);
and U1667 (N_1667,In_2774,In_1030);
and U1668 (N_1668,In_1433,In_1675);
xnor U1669 (N_1669,In_4164,In_2286);
nor U1670 (N_1670,In_1209,In_1248);
nand U1671 (N_1671,In_4624,In_1332);
and U1672 (N_1672,In_1292,In_4124);
xnor U1673 (N_1673,In_4737,In_3053);
or U1674 (N_1674,In_569,In_4825);
and U1675 (N_1675,In_2829,In_2745);
and U1676 (N_1676,In_4643,In_585);
nor U1677 (N_1677,In_4510,In_2761);
or U1678 (N_1678,In_619,In_2152);
nand U1679 (N_1679,In_4151,In_3605);
and U1680 (N_1680,In_3121,In_4460);
nand U1681 (N_1681,In_2298,In_1823);
xor U1682 (N_1682,In_2595,In_2509);
and U1683 (N_1683,In_1034,In_1337);
or U1684 (N_1684,In_1610,In_2867);
nand U1685 (N_1685,In_3133,In_729);
xnor U1686 (N_1686,In_3596,In_2570);
nor U1687 (N_1687,In_4564,In_3391);
nand U1688 (N_1688,In_1883,In_2890);
nand U1689 (N_1689,In_3165,In_0);
or U1690 (N_1690,In_4323,In_2574);
xnor U1691 (N_1691,In_1023,In_4245);
nand U1692 (N_1692,In_3959,In_2084);
nor U1693 (N_1693,In_2186,In_4001);
or U1694 (N_1694,In_4864,In_4975);
xor U1695 (N_1695,In_4636,In_4168);
xnor U1696 (N_1696,In_652,In_3062);
nor U1697 (N_1697,In_1717,In_2335);
and U1698 (N_1698,In_4237,In_970);
nand U1699 (N_1699,In_3281,In_4176);
or U1700 (N_1700,In_979,In_3197);
xor U1701 (N_1701,In_1252,In_121);
or U1702 (N_1702,In_1355,In_2113);
or U1703 (N_1703,In_3160,In_2878);
xor U1704 (N_1704,In_2328,In_4736);
xnor U1705 (N_1705,In_1525,In_952);
nand U1706 (N_1706,In_4781,In_3410);
xor U1707 (N_1707,In_3533,In_1402);
xnor U1708 (N_1708,In_311,In_4649);
or U1709 (N_1709,In_2736,In_4792);
xnor U1710 (N_1710,In_2804,In_2927);
nor U1711 (N_1711,In_1027,In_3143);
nand U1712 (N_1712,In_1143,In_1640);
xor U1713 (N_1713,In_3386,In_1216);
nand U1714 (N_1714,In_2827,In_3254);
nor U1715 (N_1715,In_2536,In_3824);
nor U1716 (N_1716,In_3976,In_3313);
and U1717 (N_1717,In_1694,In_3427);
or U1718 (N_1718,In_186,In_461);
or U1719 (N_1719,In_4272,In_1504);
xnor U1720 (N_1720,In_357,In_3312);
nor U1721 (N_1721,In_2264,In_1);
nor U1722 (N_1722,In_1076,In_1843);
nor U1723 (N_1723,In_3858,In_306);
xnor U1724 (N_1724,In_3190,In_4579);
nor U1725 (N_1725,In_3073,In_4009);
or U1726 (N_1726,In_4972,In_4043);
nor U1727 (N_1727,In_4268,In_840);
xor U1728 (N_1728,In_4589,In_4839);
nand U1729 (N_1729,In_3965,In_3796);
or U1730 (N_1730,In_2390,In_310);
xnor U1731 (N_1731,In_4993,In_1959);
nand U1732 (N_1732,In_2436,In_4930);
nor U1733 (N_1733,In_3495,In_3946);
xnor U1734 (N_1734,In_1820,In_2972);
xnor U1735 (N_1735,In_2153,In_4551);
or U1736 (N_1736,In_976,In_2566);
or U1737 (N_1737,In_3233,In_2447);
xor U1738 (N_1738,In_2421,In_3066);
nor U1739 (N_1739,In_2420,In_895);
nand U1740 (N_1740,In_4758,In_4392);
nand U1741 (N_1741,In_55,In_573);
or U1742 (N_1742,In_1625,In_2930);
nor U1743 (N_1743,In_1029,In_2193);
xnor U1744 (N_1744,In_2281,In_3397);
or U1745 (N_1745,In_1356,In_568);
or U1746 (N_1746,In_1811,In_2407);
or U1747 (N_1747,In_812,In_2181);
and U1748 (N_1748,In_1136,In_1428);
nand U1749 (N_1749,In_255,In_2204);
nand U1750 (N_1750,In_1534,In_2849);
xnor U1751 (N_1751,In_4244,In_697);
and U1752 (N_1752,In_624,In_886);
nand U1753 (N_1753,In_3167,In_2797);
xor U1754 (N_1754,In_3373,In_653);
nand U1755 (N_1755,In_1926,In_3257);
xnor U1756 (N_1756,In_3168,In_3550);
or U1757 (N_1757,In_2359,In_3051);
xnor U1758 (N_1758,In_4418,In_2599);
nand U1759 (N_1759,In_2252,In_4678);
xor U1760 (N_1760,In_2873,In_2799);
or U1761 (N_1761,In_2346,In_3717);
and U1762 (N_1762,In_3928,In_3646);
and U1763 (N_1763,In_2275,In_521);
nor U1764 (N_1764,In_4351,In_679);
or U1765 (N_1765,In_1809,In_4271);
and U1766 (N_1766,In_612,In_4592);
xor U1767 (N_1767,In_1371,In_1185);
xnor U1768 (N_1768,In_1732,In_2216);
and U1769 (N_1769,In_2693,In_4823);
nor U1770 (N_1770,In_1943,In_4907);
xnor U1771 (N_1771,In_2546,In_4454);
xor U1772 (N_1772,In_324,In_4120);
and U1773 (N_1773,In_491,In_2262);
and U1774 (N_1774,In_3344,In_3377);
nand U1775 (N_1775,In_4456,In_2613);
and U1776 (N_1776,In_1176,In_4696);
and U1777 (N_1777,In_4008,In_3744);
or U1778 (N_1778,In_3788,In_876);
or U1779 (N_1779,In_4612,In_4910);
nand U1780 (N_1780,In_1111,In_2784);
nor U1781 (N_1781,In_973,In_4067);
and U1782 (N_1782,In_4406,In_1476);
nor U1783 (N_1783,In_1318,In_3069);
xor U1784 (N_1784,In_4320,In_3819);
nand U1785 (N_1785,In_871,In_1351);
or U1786 (N_1786,In_2329,In_2918);
or U1787 (N_1787,In_1378,In_1965);
xnor U1788 (N_1788,In_467,In_1280);
nand U1789 (N_1789,In_1274,In_776);
nand U1790 (N_1790,In_2821,In_2305);
nor U1791 (N_1791,In_2905,In_4735);
or U1792 (N_1792,In_1617,In_3005);
xnor U1793 (N_1793,In_1559,In_4534);
or U1794 (N_1794,In_1699,In_2154);
nor U1795 (N_1795,In_2135,In_3065);
and U1796 (N_1796,In_203,In_1573);
nand U1797 (N_1797,In_2540,In_3010);
and U1798 (N_1798,In_1158,In_3873);
and U1799 (N_1799,In_694,In_3419);
nor U1800 (N_1800,In_1219,In_1972);
xor U1801 (N_1801,In_2872,In_1408);
nor U1802 (N_1802,In_1624,In_4346);
xor U1803 (N_1803,In_325,In_1225);
xnor U1804 (N_1804,In_3623,In_1217);
or U1805 (N_1805,In_458,In_3562);
nand U1806 (N_1806,In_1228,In_2011);
nand U1807 (N_1807,In_1891,In_1631);
xor U1808 (N_1808,In_2312,In_4068);
and U1809 (N_1809,In_2365,In_4146);
xnor U1810 (N_1810,In_1072,In_4963);
xnor U1811 (N_1811,In_681,In_416);
nand U1812 (N_1812,In_946,In_1480);
nor U1813 (N_1813,In_4018,In_3635);
and U1814 (N_1814,In_1164,In_1718);
xor U1815 (N_1815,In_2380,In_351);
nand U1816 (N_1816,In_1039,In_3671);
and U1817 (N_1817,In_4965,In_1260);
nand U1818 (N_1818,In_1938,In_3260);
xnor U1819 (N_1819,In_3850,In_12);
xnor U1820 (N_1820,In_4002,In_641);
xnor U1821 (N_1821,In_2605,In_4097);
and U1822 (N_1822,In_3201,In_698);
nand U1823 (N_1823,In_4747,In_2593);
or U1824 (N_1824,In_327,In_3462);
and U1825 (N_1825,In_3837,In_2879);
nand U1826 (N_1826,In_1577,In_4082);
nor U1827 (N_1827,In_2310,In_3675);
nand U1828 (N_1828,In_4253,In_1681);
nand U1829 (N_1829,In_787,In_1944);
and U1830 (N_1830,In_4077,In_3098);
nor U1831 (N_1831,In_1352,In_2502);
and U1832 (N_1832,In_3702,In_1457);
nor U1833 (N_1833,In_1064,In_3204);
xnor U1834 (N_1834,In_1458,In_750);
and U1835 (N_1835,In_4489,In_1069);
and U1836 (N_1836,In_3795,In_1199);
xor U1837 (N_1837,In_2010,In_1629);
and U1838 (N_1838,In_4276,In_167);
nor U1839 (N_1839,In_4078,In_1122);
nor U1840 (N_1840,In_3264,In_3728);
xnor U1841 (N_1841,In_986,In_2266);
xnor U1842 (N_1842,In_3791,In_2894);
and U1843 (N_1843,In_1182,In_145);
nand U1844 (N_1844,In_1822,In_3726);
xnor U1845 (N_1845,In_1803,In_2962);
nand U1846 (N_1846,In_2698,In_2662);
or U1847 (N_1847,In_1042,In_4556);
nand U1848 (N_1848,In_1762,In_4906);
and U1849 (N_1849,In_4830,In_3773);
or U1850 (N_1850,In_4845,In_4243);
xnor U1851 (N_1851,In_3584,In_3099);
nor U1852 (N_1852,In_4265,In_1349);
and U1853 (N_1853,In_84,In_3327);
or U1854 (N_1854,In_3723,In_1036);
xnor U1855 (N_1855,In_4409,In_4952);
nand U1856 (N_1856,In_3730,In_4063);
and U1857 (N_1857,In_3956,In_3512);
or U1858 (N_1858,In_4095,In_1502);
or U1859 (N_1859,In_3847,In_2825);
nor U1860 (N_1860,In_1692,In_3372);
nand U1861 (N_1861,In_313,In_4733);
or U1862 (N_1862,In_4886,In_869);
nor U1863 (N_1863,In_488,In_1096);
nand U1864 (N_1864,In_4100,In_3581);
nand U1865 (N_1865,In_547,In_3368);
nor U1866 (N_1866,In_4671,In_2562);
and U1867 (N_1867,In_4359,In_1005);
and U1868 (N_1868,In_4135,In_2484);
nand U1869 (N_1869,In_3935,In_62);
and U1870 (N_1870,In_3157,In_1206);
nor U1871 (N_1871,In_449,In_4732);
and U1872 (N_1872,In_4705,In_3423);
nor U1873 (N_1873,In_354,In_3932);
and U1874 (N_1874,In_4766,In_1701);
and U1875 (N_1875,In_4311,In_159);
and U1876 (N_1876,In_2462,In_2274);
or U1877 (N_1877,In_4870,In_2191);
or U1878 (N_1878,In_2472,In_1420);
or U1879 (N_1879,In_3456,In_3488);
or U1880 (N_1880,In_1979,In_2834);
nor U1881 (N_1881,In_3737,In_1914);
xor U1882 (N_1882,In_621,In_1015);
nand U1883 (N_1883,In_3348,In_2069);
nand U1884 (N_1884,In_2970,In_2718);
nand U1885 (N_1885,In_2560,In_266);
nand U1886 (N_1886,In_3805,In_875);
and U1887 (N_1887,In_874,In_2785);
xnor U1888 (N_1888,In_2789,In_2585);
nand U1889 (N_1889,In_3490,In_2902);
nand U1890 (N_1890,In_1013,In_4180);
or U1891 (N_1891,In_213,In_4059);
xor U1892 (N_1892,In_4447,In_4184);
xnor U1893 (N_1893,In_4650,In_1196);
xnor U1894 (N_1894,In_3829,In_4287);
nand U1895 (N_1895,In_3626,In_988);
and U1896 (N_1896,In_1588,In_4491);
or U1897 (N_1897,In_3086,In_769);
xnor U1898 (N_1898,In_2977,In_2213);
nand U1899 (N_1899,In_2964,In_4915);
and U1900 (N_1900,In_3275,In_3304);
nand U1901 (N_1901,In_4404,In_1733);
nand U1902 (N_1902,In_1532,In_1591);
nor U1903 (N_1903,In_3708,In_4300);
nor U1904 (N_1904,In_2115,In_863);
xnor U1905 (N_1905,In_4322,In_3985);
xor U1906 (N_1906,In_2798,In_1310);
and U1907 (N_1907,In_4395,In_2192);
xor U1908 (N_1908,In_583,In_4818);
xor U1909 (N_1909,In_2042,In_1403);
nor U1910 (N_1910,In_131,In_3205);
nand U1911 (N_1911,In_1257,In_2050);
or U1912 (N_1912,In_328,In_1593);
xor U1913 (N_1913,In_2464,In_4518);
and U1914 (N_1914,In_4616,In_3920);
xor U1915 (N_1915,In_2953,In_1150);
and U1916 (N_1916,In_382,In_3224);
and U1917 (N_1917,In_420,In_2769);
nor U1918 (N_1918,In_3713,In_1936);
and U1919 (N_1919,In_1784,In_284);
nand U1920 (N_1920,In_216,In_1000);
nand U1921 (N_1921,In_2537,In_2307);
xor U1922 (N_1922,In_2634,In_1315);
or U1923 (N_1923,In_3357,In_4617);
and U1924 (N_1924,In_4147,In_4403);
and U1925 (N_1925,In_2617,In_1773);
and U1926 (N_1926,In_1427,In_3551);
nand U1927 (N_1927,In_905,In_37);
nand U1928 (N_1928,In_2422,In_1127);
xor U1929 (N_1929,In_253,In_1859);
nor U1930 (N_1930,In_2006,In_1499);
nor U1931 (N_1931,In_2185,In_1685);
nor U1932 (N_1932,In_1839,In_4122);
or U1933 (N_1933,In_3556,In_4722);
nand U1934 (N_1934,In_2257,In_4369);
nor U1935 (N_1935,In_2123,In_169);
or U1936 (N_1936,In_2988,In_2704);
and U1937 (N_1937,In_364,In_2073);
and U1938 (N_1938,In_4399,In_2045);
nand U1939 (N_1939,In_316,In_578);
nor U1940 (N_1940,In_767,In_25);
nand U1941 (N_1941,In_3162,In_2383);
and U1942 (N_1942,In_3610,In_935);
nor U1943 (N_1943,In_2946,In_34);
and U1944 (N_1944,In_1871,In_2095);
nor U1945 (N_1945,In_2576,In_2297);
nand U1946 (N_1946,In_2172,In_4639);
xor U1947 (N_1947,In_692,In_1606);
nor U1948 (N_1948,In_1133,In_3012);
xnor U1949 (N_1949,In_4083,In_1824);
or U1950 (N_1950,In_3418,In_1297);
xor U1951 (N_1951,In_3440,In_2384);
and U1952 (N_1952,In_110,In_1522);
xor U1953 (N_1953,In_3104,In_2587);
nor U1954 (N_1954,In_4228,In_3546);
xor U1955 (N_1955,In_3057,In_3747);
xor U1956 (N_1956,In_3711,In_194);
and U1957 (N_1957,In_3658,In_4544);
nand U1958 (N_1958,In_3696,In_1201);
nor U1959 (N_1959,In_1881,In_2792);
or U1960 (N_1960,In_2564,In_2159);
nand U1961 (N_1961,In_4923,In_3783);
nor U1962 (N_1962,In_3078,In_4143);
nor U1963 (N_1963,In_2418,In_3597);
nor U1964 (N_1964,In_4708,In_1422);
and U1965 (N_1965,In_3175,In_4493);
nand U1966 (N_1966,In_821,In_231);
and U1967 (N_1967,In_4475,In_2330);
nand U1968 (N_1968,In_3298,In_2465);
xor U1969 (N_1969,In_3491,In_2806);
or U1970 (N_1970,In_4939,In_4081);
and U1971 (N_1971,In_1198,In_19);
xor U1972 (N_1972,In_3174,In_2731);
or U1973 (N_1973,In_2277,In_1904);
and U1974 (N_1974,In_647,In_426);
xnor U1975 (N_1975,In_3274,In_3669);
or U1976 (N_1976,In_3435,In_3152);
xor U1977 (N_1977,In_150,In_918);
nand U1978 (N_1978,In_3325,In_1654);
nor U1979 (N_1979,In_1848,In_1344);
nand U1980 (N_1980,In_242,In_3471);
nor U1981 (N_1981,In_2070,In_4260);
xnor U1982 (N_1982,In_1410,In_2409);
and U1983 (N_1983,In_1432,In_3738);
or U1984 (N_1984,In_119,In_486);
nor U1985 (N_1985,In_3984,In_4209);
nor U1986 (N_1986,In_3396,In_3540);
xnor U1987 (N_1987,In_948,In_2943);
and U1988 (N_1988,In_2285,In_4984);
nand U1989 (N_1989,In_3132,In_2217);
or U1990 (N_1990,In_1021,In_2847);
nor U1991 (N_1991,In_550,In_4942);
xnor U1992 (N_1992,In_4092,In_2250);
and U1993 (N_1993,In_3839,In_3525);
xnor U1994 (N_1994,In_454,In_473);
nor U1995 (N_1995,In_4150,In_13);
and U1996 (N_1996,In_3615,In_1193);
nand U1997 (N_1997,In_3015,In_4494);
nand U1998 (N_1998,In_878,In_2717);
nor U1999 (N_1999,In_4098,In_3601);
or U2000 (N_2000,In_4630,In_2248);
nand U2001 (N_2001,In_71,In_292);
xor U2002 (N_2002,In_775,In_2871);
or U2003 (N_2003,In_1566,In_4982);
nand U2004 (N_2004,In_1053,In_3210);
nand U2005 (N_2005,In_3349,In_2178);
xnor U2006 (N_2006,In_3735,In_147);
nor U2007 (N_2007,In_3923,In_1178);
and U2008 (N_2008,In_1856,In_3042);
xor U2009 (N_2009,In_4328,In_1584);
xor U2010 (N_2010,In_3392,In_2775);
and U2011 (N_2011,In_1876,In_245);
nor U2012 (N_2012,In_2854,In_291);
and U2013 (N_2013,In_4519,In_4559);
and U2014 (N_2014,In_4229,In_4279);
or U2015 (N_2015,In_2280,In_4856);
nand U2016 (N_2016,In_2430,In_2928);
xor U2017 (N_2017,In_2539,In_4282);
nor U2018 (N_2018,In_120,In_4366);
or U2019 (N_2019,In_1840,In_1037);
and U2020 (N_2020,In_2931,In_1126);
nor U2021 (N_2021,In_567,In_3970);
nand U2022 (N_2022,In_4672,In_1785);
or U2023 (N_2023,In_3852,In_3869);
nor U2024 (N_2024,In_4978,In_3936);
or U2025 (N_2025,In_3589,In_1705);
nand U2026 (N_2026,In_3064,In_2327);
nor U2027 (N_2027,In_3535,In_2802);
nand U2028 (N_2028,In_3134,In_4467);
or U2029 (N_2029,In_2270,In_4739);
or U2030 (N_2030,In_1898,In_1299);
nand U2031 (N_2031,In_3022,In_4428);
nand U2032 (N_2032,In_3240,In_2490);
xnor U2033 (N_2033,In_3759,In_232);
or U2034 (N_2034,In_1854,In_2727);
xor U2035 (N_2035,In_4336,In_289);
nor U2036 (N_2036,In_348,In_1841);
nor U2037 (N_2037,In_4695,In_838);
nor U2038 (N_2038,In_3489,In_2982);
and U2039 (N_2039,In_4349,In_4960);
nand U2040 (N_2040,In_4815,In_4241);
xor U2041 (N_2041,In_1713,In_2163);
nor U2042 (N_2042,In_2198,In_394);
nand U2043 (N_2043,In_3101,In_774);
xor U2044 (N_2044,In_2912,In_4674);
or U2045 (N_2045,In_3365,In_2094);
xor U2046 (N_2046,In_2728,In_2500);
or U2047 (N_2047,In_2648,In_1771);
or U2048 (N_2048,In_47,In_1622);
or U2049 (N_2049,In_4423,In_3409);
nand U2050 (N_2050,In_928,In_4353);
nor U2051 (N_2051,In_593,In_4431);
nand U2052 (N_2052,In_588,In_3334);
nand U2053 (N_2053,In_3606,In_1287);
nand U2054 (N_2054,In_1564,In_1238);
or U2055 (N_2055,In_393,In_4478);
nor U2056 (N_2056,In_4581,In_4587);
nor U2057 (N_2057,In_3303,In_2342);
or U2058 (N_2058,In_1808,In_4413);
xnor U2059 (N_2059,In_2692,In_263);
and U2060 (N_2060,In_1621,In_3638);
nand U2061 (N_2061,In_1655,In_3308);
nor U2062 (N_2062,In_2683,In_4112);
nand U2063 (N_2063,In_1947,In_3156);
and U2064 (N_2064,In_972,In_4846);
and U2065 (N_2065,In_1431,In_910);
or U2066 (N_2066,In_4495,In_319);
and U2067 (N_2067,In_1307,In_3109);
xor U2068 (N_2068,In_1284,In_4330);
or U2069 (N_2069,In_3865,In_1786);
nand U2070 (N_2070,In_2543,In_1885);
xor U2071 (N_2071,In_3801,In_4086);
nand U2072 (N_2072,In_439,In_4641);
nand U2073 (N_2073,In_4833,In_4391);
or U2074 (N_2074,In_851,In_2404);
nand U2075 (N_2075,In_546,In_2271);
xnor U2076 (N_2076,In_3164,In_3560);
or U2077 (N_2077,In_38,In_3781);
or U2078 (N_2078,In_3636,In_3037);
nand U2079 (N_2079,In_1779,In_4529);
or U2080 (N_2080,In_2607,In_3672);
nor U2081 (N_2081,In_2532,In_1890);
and U2082 (N_2082,In_376,In_1235);
nand U2083 (N_2083,In_4281,In_1752);
xnor U2084 (N_2084,In_4440,In_3685);
nor U2085 (N_2085,In_3667,In_3893);
xnor U2086 (N_2086,In_959,In_3944);
or U2087 (N_2087,In_3797,In_3208);
nand U2088 (N_2088,In_4204,In_4477);
nand U2089 (N_2089,In_338,In_3246);
or U2090 (N_2090,In_4887,In_447);
or U2091 (N_2091,In_3421,In_3420);
nor U2092 (N_2092,In_3787,In_2033);
nor U2093 (N_2093,In_818,In_406);
nand U2094 (N_2094,In_2921,In_4052);
xnor U2095 (N_2095,In_803,In_2224);
nor U2096 (N_2096,In_3390,In_4277);
and U2097 (N_2097,In_3118,In_4668);
or U2098 (N_2098,In_398,In_3021);
and U2099 (N_2099,In_3351,In_4240);
and U2100 (N_2100,In_4609,In_2758);
or U2101 (N_2101,In_1148,In_919);
or U2102 (N_2102,In_1509,In_3608);
and U2103 (N_2103,In_282,In_226);
xnor U2104 (N_2104,In_2647,In_202);
or U2105 (N_2105,In_3151,In_2695);
or U2106 (N_2106,In_4848,In_1974);
or U2107 (N_2107,In_4005,In_3707);
or U2108 (N_2108,In_1369,In_2032);
or U2109 (N_2109,In_1374,In_4023);
or U2110 (N_2110,In_3153,In_858);
nor U2111 (N_2111,In_4453,In_1301);
nand U2112 (N_2112,In_2361,In_1063);
nand U2113 (N_2113,In_1939,In_3607);
nor U2114 (N_2114,In_693,In_2508);
or U2115 (N_2115,In_4837,In_235);
and U2116 (N_2116,In_1768,In_2850);
nand U2117 (N_2117,In_3813,In_2723);
and U2118 (N_2118,In_1314,In_1901);
nand U2119 (N_2119,In_3882,In_3218);
nand U2120 (N_2120,In_1948,In_4076);
nor U2121 (N_2121,In_1312,In_4920);
xnor U2122 (N_2122,In_2051,In_1829);
and U2123 (N_2123,In_765,In_2279);
xnor U2124 (N_2124,In_3960,In_1568);
and U2125 (N_2125,In_4724,In_4424);
nor U2126 (N_2126,In_3374,In_2435);
and U2127 (N_2127,In_3040,In_4149);
or U2128 (N_2128,In_3438,In_1436);
xnor U2129 (N_2129,In_1018,In_2864);
and U2130 (N_2130,In_2363,In_4364);
nor U2131 (N_2131,In_3216,In_1153);
nor U2132 (N_2132,In_1810,In_500);
nor U2133 (N_2133,In_2171,In_1304);
xor U2134 (N_2134,In_2594,In_1886);
nand U2135 (N_2135,In_528,In_1893);
and U2136 (N_2136,In_204,In_3244);
and U2137 (N_2137,In_8,In_408);
and U2138 (N_2138,In_618,In_2314);
nor U2139 (N_2139,In_1489,In_300);
nand U2140 (N_2140,In_4922,In_4401);
or U2141 (N_2141,In_4727,In_1375);
xor U2142 (N_2142,In_1105,In_2522);
nor U2143 (N_2143,In_927,In_1070);
xnor U2144 (N_2144,In_3724,In_1663);
nor U2145 (N_2145,In_2571,In_2403);
xnor U2146 (N_2146,In_4951,In_1887);
or U2147 (N_2147,In_670,In_410);
or U2148 (N_2148,In_3561,In_2655);
or U2149 (N_2149,In_1253,In_4123);
or U2150 (N_2150,In_2200,In_2869);
xor U2151 (N_2151,In_3239,In_139);
nor U2152 (N_2152,In_3500,In_4834);
xor U2153 (N_2153,In_3116,In_3110);
nor U2154 (N_2154,In_929,In_4821);
or U2155 (N_2155,In_2886,In_4715);
nor U2156 (N_2156,In_3161,In_1518);
or U2157 (N_2157,In_2976,In_671);
or U2158 (N_2158,In_1765,In_305);
nand U2159 (N_2159,In_4357,In_1028);
or U2160 (N_2160,In_2392,In_4689);
nor U2161 (N_2161,In_127,In_4751);
and U2162 (N_2162,In_2814,In_1910);
nor U2163 (N_2163,In_2357,In_346);
nor U2164 (N_2164,In_1295,In_3800);
nand U2165 (N_2165,In_1536,In_3059);
xor U2166 (N_2166,In_2355,In_1927);
nand U2167 (N_2167,In_3417,In_3023);
nand U2168 (N_2168,In_1416,In_3629);
nor U2169 (N_2169,In_1882,In_705);
or U2170 (N_2170,In_4744,In_3306);
and U2171 (N_2171,In_153,In_3703);
or U2172 (N_2172,In_3054,In_3486);
nand U2173 (N_2173,In_4976,In_519);
nand U2174 (N_2174,In_3028,In_294);
nand U2175 (N_2175,In_3445,In_4119);
or U2176 (N_2176,In_2054,In_1450);
nand U2177 (N_2177,In_3029,In_4971);
nor U2178 (N_2178,In_2881,In_727);
xor U2179 (N_2179,In_4997,In_854);
nor U2180 (N_2180,In_1202,In_4028);
nor U2181 (N_2181,In_3598,In_4220);
nor U2182 (N_2182,In_4776,In_260);
nor U2183 (N_2183,In_4434,In_18);
xnor U2184 (N_2184,In_3446,In_4944);
nor U2185 (N_2185,In_1828,In_1918);
or U2186 (N_2186,In_1550,In_3185);
nand U2187 (N_2187,In_3243,In_2815);
or U2188 (N_2188,In_3948,In_4296);
nand U2189 (N_2189,In_3052,In_118);
nand U2190 (N_2190,In_471,In_2924);
and U2191 (N_2191,In_3200,In_602);
xnor U2192 (N_2192,In_2047,In_3573);
nor U2193 (N_2193,In_117,In_2141);
nand U2194 (N_2194,In_3451,In_4214);
or U2195 (N_2195,In_963,In_3061);
or U2196 (N_2196,In_3962,In_4429);
nor U2197 (N_2197,In_592,In_2852);
xor U2198 (N_2198,In_2445,In_4117);
xnor U2199 (N_2199,In_1092,In_4247);
and U2200 (N_2200,In_176,In_3434);
and U2201 (N_2201,In_1093,In_4368);
and U2202 (N_2202,In_3899,In_522);
nor U2203 (N_2203,In_864,In_3194);
nand U2204 (N_2204,In_1604,In_2169);
xnor U2205 (N_2205,In_1094,In_1061);
nand U2206 (N_2206,In_2697,In_2451);
xnor U2207 (N_2207,In_372,In_320);
or U2208 (N_2208,In_1365,In_4115);
xnor U2209 (N_2209,In_3182,In_3855);
xor U2210 (N_2210,In_1236,In_2110);
and U2211 (N_2211,In_87,In_1745);
or U2212 (N_2212,In_637,In_2065);
nand U2213 (N_2213,In_1224,In_699);
and U2214 (N_2214,In_2951,In_1468);
nor U2215 (N_2215,In_1954,In_2741);
nor U2216 (N_2216,In_966,In_2818);
or U2217 (N_2217,In_2126,In_770);
nand U2218 (N_2218,In_1815,In_1482);
nand U2219 (N_2219,In_4356,In_1950);
or U2220 (N_2220,In_1958,In_2833);
nor U2221 (N_2221,In_757,In_2989);
and U2222 (N_2222,In_552,In_1385);
or U2223 (N_2223,In_4182,In_525);
and U2224 (N_2224,In_4360,In_1275);
nor U2225 (N_2225,In_2523,In_135);
xor U2226 (N_2226,In_1345,In_3565);
and U2227 (N_2227,In_4745,In_2398);
nor U2228 (N_2228,In_4899,In_2643);
nand U2229 (N_2229,In_1442,In_4795);
or U2230 (N_2230,In_3613,In_3721);
xnor U2231 (N_2231,In_4291,In_4350);
xnor U2232 (N_2232,In_737,In_113);
nor U2233 (N_2233,In_404,In_1867);
or U2234 (N_2234,In_358,In_3993);
xor U2235 (N_2235,In_1746,In_3394);
and U2236 (N_2236,In_3666,In_1461);
nand U2237 (N_2237,In_3683,In_920);
or U2238 (N_2238,In_3538,In_2303);
xnor U2239 (N_2239,In_3079,In_4158);
xor U2240 (N_2240,In_108,In_1795);
nand U2241 (N_2241,In_2534,In_2529);
nor U2242 (N_2242,In_667,In_1118);
nor U2243 (N_2243,In_2493,In_2155);
xor U2244 (N_2244,In_4677,In_1171);
xnor U2245 (N_2245,In_1602,In_4861);
xnor U2246 (N_2246,In_967,In_2004);
xor U2247 (N_2247,In_3631,In_4427);
nor U2248 (N_2248,In_4706,In_518);
or U2249 (N_2249,In_1471,In_286);
xor U2250 (N_2250,In_3171,In_4032);
nor U2251 (N_2251,In_4060,In_4252);
or U2252 (N_2252,In_482,In_1763);
or U2253 (N_2253,In_3789,In_1250);
or U2254 (N_2254,In_3145,In_617);
and U2255 (N_2255,In_2710,In_2142);
nand U2256 (N_2256,In_3862,In_718);
nand U2257 (N_2257,In_3406,In_3199);
nand U2258 (N_2258,In_4348,In_2860);
xor U2259 (N_2259,In_3761,In_2341);
nand U2260 (N_2260,In_2458,In_1057);
or U2261 (N_2261,In_516,In_3543);
or U2262 (N_2262,In_103,In_955);
xnor U2263 (N_2263,In_4166,In_4608);
nand U2264 (N_2264,In_909,In_4370);
and U2265 (N_2265,In_3854,In_4760);
nand U2266 (N_2266,In_3007,In_3245);
nand U2267 (N_2267,In_374,In_2735);
or U2268 (N_2268,In_2726,In_4505);
and U2269 (N_2269,In_4408,In_1438);
nand U2270 (N_2270,In_722,In_1486);
xnor U2271 (N_2271,In_1324,In_69);
nand U2272 (N_2272,In_4202,In_589);
or U2273 (N_2273,In_1533,In_1110);
or U2274 (N_2274,In_1331,In_1160);
and U2275 (N_2275,In_2550,In_930);
nand U2276 (N_2276,In_3943,In_1043);
xnor U2277 (N_2277,In_427,In_1605);
nor U2278 (N_2278,In_690,In_527);
and U2279 (N_2279,In_665,In_1443);
and U2280 (N_2280,In_4648,In_1529);
and U2281 (N_2281,In_91,In_326);
and U2282 (N_2282,In_2325,In_4438);
nor U2283 (N_2283,In_4173,In_1635);
xnor U2284 (N_2284,In_4177,In_4087);
or U2285 (N_2285,In_1067,In_341);
nor U2286 (N_2286,In_1951,In_3727);
or U2287 (N_2287,In_3461,In_1727);
nand U2288 (N_2288,In_805,In_2468);
and U2289 (N_2289,In_3247,In_4719);
or U2290 (N_2290,In_4788,In_515);
or U2291 (N_2291,In_3514,In_224);
xnor U2292 (N_2292,In_3476,In_4203);
and U2293 (N_2293,In_3559,In_4549);
nand U2294 (N_2294,In_836,In_276);
and U2295 (N_2295,In_2038,In_830);
nand U2296 (N_2296,In_4207,In_2446);
nand U2297 (N_2297,In_3630,In_3150);
nand U2298 (N_2298,In_3739,In_3567);
or U2299 (N_2299,In_4464,In_1935);
nand U2300 (N_2300,In_2903,In_947);
and U2301 (N_2301,In_2267,In_1838);
or U2302 (N_2302,In_2831,In_4850);
nor U2303 (N_2303,In_2320,In_1801);
and U2304 (N_2304,In_2101,In_367);
and U2305 (N_2305,In_3092,In_4531);
nor U2306 (N_2306,In_2194,In_3477);
xor U2307 (N_2307,In_3482,In_1623);
or U2308 (N_2308,In_106,In_2688);
nand U2309 (N_2309,In_4125,In_4552);
nor U2310 (N_2310,In_3831,In_1500);
and U2311 (N_2311,In_1451,In_2336);
or U2312 (N_2312,In_1109,In_740);
xor U2313 (N_2313,In_3380,In_182);
nor U2314 (N_2314,In_1207,In_1545);
or U2315 (N_2315,In_3564,In_2674);
nor U2316 (N_2316,In_499,In_4421);
xor U2317 (N_2317,In_1508,In_2377);
nor U2318 (N_2318,In_2144,In_1983);
xnor U2319 (N_2319,In_1963,In_1414);
nor U2320 (N_2320,In_1181,In_2394);
xor U2321 (N_2321,In_2176,In_1446);
nor U2322 (N_2322,In_3997,In_2001);
nand U2323 (N_2323,In_4072,In_4315);
or U2324 (N_2324,In_2936,In_4365);
nor U2325 (N_2325,In_2096,In_2322);
and U2326 (N_2326,In_4969,In_2150);
nand U2327 (N_2327,In_220,In_494);
nor U2328 (N_2328,In_4700,In_4968);
xor U2329 (N_2329,In_2189,In_3326);
and U2330 (N_2330,In_4597,In_1222);
xor U2331 (N_2331,In_1449,In_4254);
nor U2332 (N_2332,In_4010,In_4611);
or U2333 (N_2333,In_4683,In_3212);
nand U2334 (N_2334,In_68,In_4763);
nor U2335 (N_2335,In_3031,In_4469);
or U2336 (N_2336,In_4591,In_2572);
or U2337 (N_2337,In_4016,In_2208);
and U2338 (N_2338,In_2733,In_1011);
xnor U2339 (N_2339,In_1671,In_2691);
nor U2340 (N_2340,In_4844,In_2778);
xnor U2341 (N_2341,In_4879,In_1998);
nand U2342 (N_2342,In_3822,In_1493);
xnor U2343 (N_2343,In_2388,In_4688);
xor U2344 (N_2344,In_3580,In_3657);
or U2345 (N_2345,In_2253,In_83);
and U2346 (N_2346,In_1426,In_4703);
nand U2347 (N_2347,In_809,In_3649);
nand U2348 (N_2348,In_4698,In_760);
or U2349 (N_2349,In_1084,In_4940);
or U2350 (N_2350,In_252,In_4171);
and U2351 (N_2351,In_3399,In_3768);
xnor U2352 (N_2352,In_758,In_4868);
or U2353 (N_2353,In_3971,In_4574);
nor U2354 (N_2354,In_4729,In_4520);
nor U2355 (N_2355,In_4375,In_3379);
and U2356 (N_2356,In_2504,In_299);
nand U2357 (N_2357,In_1689,In_937);
nand U2358 (N_2358,In_2232,In_4554);
nand U2359 (N_2359,In_4080,In_721);
nor U2360 (N_2360,In_1131,In_2489);
or U2361 (N_2361,In_4828,In_490);
or U2362 (N_2362,In_4895,In_674);
nand U2363 (N_2363,In_1437,In_1855);
and U2364 (N_2364,In_2994,In_4626);
nor U2365 (N_2365,In_1920,In_777);
and U2366 (N_2366,In_788,In_4826);
xnor U2367 (N_2367,In_1554,In_3752);
or U2368 (N_2368,In_3736,In_1483);
xnor U2369 (N_2369,In_3447,In_1452);
xor U2370 (N_2370,In_4303,In_2160);
nor U2371 (N_2371,In_2114,In_4913);
or U2372 (N_2372,In_4873,In_4049);
nand U2373 (N_2373,In_3453,In_460);
nor U2374 (N_2374,In_1860,In_452);
and U2375 (N_2375,In_3191,In_4663);
xor U2376 (N_2376,In_1220,In_4988);
or U2377 (N_2377,In_4657,In_1921);
and U2378 (N_2378,In_704,In_1239);
xnor U2379 (N_2379,In_4448,In_2525);
nor U2380 (N_2380,In_1538,In_4134);
nor U2381 (N_2381,In_2244,In_4586);
nor U2382 (N_2382,In_4772,In_1218);
and U2383 (N_2383,In_162,In_4841);
nor U2384 (N_2384,In_2830,In_503);
nor U2385 (N_2385,In_3468,In_3903);
nor U2386 (N_2386,In_4593,In_1510);
and U2387 (N_2387,In_2842,In_1334);
nand U2388 (N_2388,In_2645,In_1154);
and U2389 (N_2389,In_2533,In_1966);
nor U2390 (N_2390,In_626,In_3181);
and U2391 (N_2391,In_2058,In_1135);
or U2392 (N_2392,In_2480,In_278);
xor U2393 (N_2393,In_3814,In_3341);
nand U2394 (N_2394,In_1716,In_1189);
xnor U2395 (N_2395,In_4420,In_2373);
or U2396 (N_2396,In_2205,In_2507);
nor U2397 (N_2397,In_3710,In_1800);
nor U2398 (N_2398,In_1205,In_924);
nand U2399 (N_2399,In_1581,In_4896);
xor U2400 (N_2400,In_1415,In_4414);
and U2401 (N_2401,In_4911,In_4255);
nor U2402 (N_2402,In_3534,In_1114);
nand U2403 (N_2403,In_3521,In_3845);
xor U2404 (N_2404,In_403,In_1241);
and U2405 (N_2405,In_2460,In_33);
xnor U2406 (N_2406,In_1300,In_3547);
nand U2407 (N_2407,In_2282,In_4111);
or U2408 (N_2408,In_2929,In_209);
or U2409 (N_2409,In_4274,In_2759);
or U2410 (N_2410,In_3084,In_4775);
nor U2411 (N_2411,In_4675,In_852);
nand U2412 (N_2412,In_2334,In_1600);
and U2413 (N_2413,In_3674,In_2318);
or U2414 (N_2414,In_2167,In_4261);
nand U2415 (N_2415,In_3554,In_3493);
or U2416 (N_2416,In_4327,In_1435);
nand U2417 (N_2417,In_672,In_969);
or U2418 (N_2418,In_1976,In_250);
xnor U2419 (N_2419,In_1788,In_2567);
nand U2420 (N_2420,In_1690,In_4482);
nand U2421 (N_2421,In_1276,In_3585);
xor U2422 (N_2422,In_742,In_2077);
xnor U2423 (N_2423,In_1660,In_1020);
xor U2424 (N_2424,In_3384,In_842);
nand U2425 (N_2425,In_143,In_2024);
nand U2426 (N_2426,In_939,In_1850);
xnor U2427 (N_2427,In_1952,In_2374);
nor U2428 (N_2428,In_756,In_141);
and U2429 (N_2429,In_4740,In_1165);
xor U2430 (N_2430,In_1714,In_1138);
nor U2431 (N_2431,In_421,In_4594);
nand U2432 (N_2432,In_3502,In_702);
nand U2433 (N_2433,In_2922,In_4036);
or U2434 (N_2434,In_668,In_1303);
and U2435 (N_2435,In_1082,In_2667);
nand U2436 (N_2436,In_3955,In_2076);
and U2437 (N_2437,In_1210,In_2237);
nand U2438 (N_2438,In_155,In_2107);
xor U2439 (N_2439,In_2364,In_2481);
nor U2440 (N_2440,In_2668,In_834);
or U2441 (N_2441,In_2174,In_3871);
nand U2442 (N_2442,In_464,In_1112);
nand U2443 (N_2443,In_4852,In_456);
nand U2444 (N_2444,In_3342,In_4547);
and U2445 (N_2445,In_60,In_2452);
and U2446 (N_2446,In_4768,In_1874);
and U2447 (N_2447,In_2316,In_2023);
xor U2448 (N_2448,In_1059,In_1962);
nand U2449 (N_2449,In_80,In_3762);
xor U2450 (N_2450,In_3426,In_1163);
nand U2451 (N_2451,In_2021,In_1335);
and U2452 (N_2452,In_3668,In_4754);
or U2453 (N_2453,In_429,In_843);
or U2454 (N_2454,In_1386,In_2175);
or U2455 (N_2455,In_4439,In_352);
and U2456 (N_2456,In_2978,In_3974);
and U2457 (N_2457,In_2337,In_1383);
or U2458 (N_2458,In_1589,In_2764);
or U2459 (N_2459,In_3812,In_3699);
xor U2460 (N_2460,In_3267,In_4701);
or U2461 (N_2461,In_632,In_3582);
or U2462 (N_2462,In_1991,In_3604);
or U2463 (N_2463,In_3978,In_3815);
and U2464 (N_2464,In_1106,In_3371);
nor U2465 (N_2465,In_1653,In_4206);
xor U2466 (N_2466,In_4227,In_3619);
nor U2467 (N_2467,In_916,In_751);
or U2468 (N_2468,In_79,In_4412);
nor U2469 (N_2469,In_264,In_1953);
and U2470 (N_2470,In_4808,In_4685);
nor U2471 (N_2471,In_1054,In_3570);
nor U2472 (N_2472,In_3071,In_1273);
or U2473 (N_2473,In_825,In_564);
nor U2474 (N_2474,In_1488,In_2851);
nor U2475 (N_2475,In_2554,In_3195);
or U2476 (N_2476,In_4949,In_1162);
nor U2477 (N_2477,In_3778,In_1479);
nand U2478 (N_2478,In_3320,In_3973);
nor U2479 (N_2479,In_3864,In_4743);
and U2480 (N_2480,In_1889,In_1121);
nor U2481 (N_2481,In_3206,In_574);
and U2482 (N_2482,In_2582,In_2426);
nand U2483 (N_2483,In_2573,In_3494);
nand U2484 (N_2484,In_4966,In_2762);
nor U2485 (N_2485,In_3941,In_448);
and U2486 (N_2486,In_1541,In_4307);
nor U2487 (N_2487,In_3600,In_4333);
xor U2488 (N_2488,In_1734,In_541);
and U2489 (N_2489,In_4299,In_1562);
xnor U2490 (N_2490,In_655,In_3068);
or U2491 (N_2491,In_3430,In_1249);
or U2492 (N_2492,In_4256,In_1372);
xor U2493 (N_2493,In_146,In_4105);
and U2494 (N_2494,In_2419,In_2448);
or U2495 (N_2495,In_2256,In_2064);
nor U2496 (N_2496,In_2685,In_3999);
nand U2497 (N_2497,In_1925,In_3058);
nand U2498 (N_2498,In_2140,In_3734);
nand U2499 (N_2499,In_3255,In_1462);
xor U2500 (N_2500,N_1157,N_2476);
or U2501 (N_2501,N_1110,N_717);
or U2502 (N_2502,N_755,N_1699);
and U2503 (N_2503,N_2119,N_1341);
or U2504 (N_2504,N_871,N_154);
xnor U2505 (N_2505,N_610,N_2274);
and U2506 (N_2506,N_1993,N_1906);
and U2507 (N_2507,N_1589,N_253);
and U2508 (N_2508,N_1401,N_368);
and U2509 (N_2509,N_2068,N_2116);
xor U2510 (N_2510,N_1420,N_97);
nor U2511 (N_2511,N_2468,N_762);
xor U2512 (N_2512,N_967,N_1412);
nand U2513 (N_2513,N_2220,N_2249);
and U2514 (N_2514,N_1601,N_815);
xor U2515 (N_2515,N_2262,N_309);
and U2516 (N_2516,N_1124,N_988);
nor U2517 (N_2517,N_1723,N_2366);
nand U2518 (N_2518,N_2238,N_446);
or U2519 (N_2519,N_379,N_1178);
and U2520 (N_2520,N_2266,N_24);
nand U2521 (N_2521,N_1541,N_177);
xnor U2522 (N_2522,N_1977,N_506);
or U2523 (N_2523,N_655,N_573);
nand U2524 (N_2524,N_2372,N_1599);
and U2525 (N_2525,N_1812,N_2190);
or U2526 (N_2526,N_1400,N_1422);
and U2527 (N_2527,N_727,N_2030);
or U2528 (N_2528,N_1384,N_269);
nor U2529 (N_2529,N_1170,N_518);
or U2530 (N_2530,N_1956,N_541);
or U2531 (N_2531,N_2141,N_759);
and U2532 (N_2532,N_308,N_1509);
nand U2533 (N_2533,N_1221,N_1835);
nor U2534 (N_2534,N_262,N_1694);
nand U2535 (N_2535,N_882,N_942);
and U2536 (N_2536,N_1173,N_2046);
nand U2537 (N_2537,N_1647,N_2304);
xnor U2538 (N_2538,N_2165,N_2154);
xor U2539 (N_2539,N_367,N_965);
or U2540 (N_2540,N_462,N_658);
nand U2541 (N_2541,N_774,N_547);
and U2542 (N_2542,N_2383,N_472);
nor U2543 (N_2543,N_1714,N_2260);
xnor U2544 (N_2544,N_1641,N_1101);
or U2545 (N_2545,N_1482,N_1668);
and U2546 (N_2546,N_495,N_1710);
and U2547 (N_2547,N_1770,N_412);
nand U2548 (N_2548,N_587,N_2496);
nor U2549 (N_2549,N_685,N_635);
or U2550 (N_2550,N_2329,N_158);
nand U2551 (N_2551,N_1379,N_591);
nor U2552 (N_2552,N_519,N_350);
nand U2553 (N_2553,N_1343,N_1188);
nor U2554 (N_2554,N_66,N_1697);
or U2555 (N_2555,N_544,N_1167);
or U2556 (N_2556,N_2302,N_1480);
and U2557 (N_2557,N_829,N_789);
and U2558 (N_2558,N_1107,N_2074);
and U2559 (N_2559,N_665,N_1499);
or U2560 (N_2560,N_1204,N_1251);
or U2561 (N_2561,N_411,N_1455);
nand U2562 (N_2562,N_776,N_1963);
and U2563 (N_2563,N_1784,N_513);
nor U2564 (N_2564,N_1381,N_2129);
and U2565 (N_2565,N_819,N_950);
xor U2566 (N_2566,N_1155,N_2282);
or U2567 (N_2567,N_2297,N_732);
nand U2568 (N_2568,N_456,N_861);
and U2569 (N_2569,N_2354,N_1281);
nand U2570 (N_2570,N_1225,N_729);
or U2571 (N_2571,N_469,N_54);
and U2572 (N_2572,N_1100,N_981);
or U2573 (N_2573,N_2182,N_364);
xnor U2574 (N_2574,N_2093,N_466);
xnor U2575 (N_2575,N_1123,N_178);
and U2576 (N_2576,N_1563,N_1873);
nor U2577 (N_2577,N_468,N_1266);
or U2578 (N_2578,N_767,N_2479);
nand U2579 (N_2579,N_1255,N_1529);
xor U2580 (N_2580,N_1994,N_482);
or U2581 (N_2581,N_1539,N_1036);
xor U2582 (N_2582,N_1942,N_2015);
and U2583 (N_2583,N_1282,N_2237);
and U2584 (N_2584,N_1559,N_2127);
xor U2585 (N_2585,N_1201,N_1461);
or U2586 (N_2586,N_1958,N_1317);
or U2587 (N_2587,N_2310,N_1081);
or U2588 (N_2588,N_1274,N_169);
and U2589 (N_2589,N_1872,N_1339);
or U2590 (N_2590,N_2031,N_167);
or U2591 (N_2591,N_535,N_413);
nor U2592 (N_2592,N_1376,N_285);
or U2593 (N_2593,N_80,N_1314);
nor U2594 (N_2594,N_2184,N_1626);
and U2595 (N_2595,N_1236,N_372);
and U2596 (N_2596,N_1181,N_2273);
or U2597 (N_2597,N_838,N_422);
xor U2598 (N_2598,N_1202,N_71);
nor U2599 (N_2599,N_2392,N_991);
xnor U2600 (N_2600,N_927,N_2358);
nand U2601 (N_2601,N_576,N_686);
or U2602 (N_2602,N_1740,N_1351);
and U2603 (N_2603,N_969,N_1816);
nor U2604 (N_2604,N_1187,N_1088);
xnor U2605 (N_2605,N_1238,N_1260);
or U2606 (N_2606,N_1556,N_130);
and U2607 (N_2607,N_83,N_159);
nor U2608 (N_2608,N_1834,N_2123);
xnor U2609 (N_2609,N_1063,N_596);
nor U2610 (N_2610,N_2294,N_1295);
or U2611 (N_2611,N_1980,N_890);
or U2612 (N_2612,N_2363,N_1442);
nor U2613 (N_2613,N_1790,N_488);
nand U2614 (N_2614,N_2150,N_1961);
xnor U2615 (N_2615,N_444,N_438);
nand U2616 (N_2616,N_376,N_88);
xor U2617 (N_2617,N_28,N_624);
nand U2618 (N_2618,N_1566,N_2126);
or U2619 (N_2619,N_2198,N_1995);
or U2620 (N_2620,N_1015,N_94);
or U2621 (N_2621,N_876,N_1273);
xor U2622 (N_2622,N_1753,N_1917);
nand U2623 (N_2623,N_1334,N_1741);
or U2624 (N_2624,N_2443,N_440);
or U2625 (N_2625,N_1750,N_494);
or U2626 (N_2626,N_608,N_2491);
nand U2627 (N_2627,N_615,N_300);
xor U2628 (N_2628,N_640,N_1734);
or U2629 (N_2629,N_2436,N_1707);
or U2630 (N_2630,N_2364,N_1012);
xnor U2631 (N_2631,N_2120,N_246);
nor U2632 (N_2632,N_779,N_2477);
or U2633 (N_2633,N_2248,N_1335);
xnor U2634 (N_2634,N_20,N_923);
or U2635 (N_2635,N_770,N_2464);
nand U2636 (N_2636,N_389,N_143);
or U2637 (N_2637,N_1861,N_1452);
nand U2638 (N_2638,N_715,N_604);
nor U2639 (N_2639,N_2102,N_1465);
or U2640 (N_2640,N_237,N_1711);
nor U2641 (N_2641,N_445,N_1965);
nor U2642 (N_2642,N_943,N_135);
xnor U2643 (N_2643,N_1720,N_1520);
nor U2644 (N_2644,N_2080,N_2047);
and U2645 (N_2645,N_2332,N_1346);
or U2646 (N_2646,N_853,N_2385);
nor U2647 (N_2647,N_216,N_607);
nand U2648 (N_2648,N_252,N_419);
nand U2649 (N_2649,N_1754,N_1970);
nor U2650 (N_2650,N_1933,N_1922);
xnor U2651 (N_2651,N_410,N_378);
nor U2652 (N_2652,N_89,N_588);
nor U2653 (N_2653,N_1193,N_1329);
and U2654 (N_2654,N_2118,N_2255);
or U2655 (N_2655,N_2444,N_2267);
nor U2656 (N_2656,N_348,N_1133);
xnor U2657 (N_2657,N_1405,N_741);
xor U2658 (N_2658,N_2140,N_1706);
nor U2659 (N_2659,N_185,N_1732);
or U2660 (N_2660,N_1206,N_534);
nor U2661 (N_2661,N_2158,N_2278);
or U2662 (N_2662,N_2131,N_296);
or U2663 (N_2663,N_1066,N_572);
nor U2664 (N_2664,N_2315,N_1211);
and U2665 (N_2665,N_1948,N_811);
xor U2666 (N_2666,N_299,N_1879);
and U2667 (N_2667,N_1165,N_2054);
nand U2668 (N_2668,N_1747,N_1368);
and U2669 (N_2669,N_1569,N_680);
and U2670 (N_2670,N_1393,N_945);
nor U2671 (N_2671,N_60,N_2099);
or U2672 (N_2672,N_1827,N_814);
xor U2673 (N_2673,N_322,N_2271);
nand U2674 (N_2674,N_1474,N_131);
xnor U2675 (N_2675,N_2293,N_875);
and U2676 (N_2676,N_1654,N_1548);
or U2677 (N_2677,N_1809,N_1851);
nand U2678 (N_2678,N_2258,N_1111);
nand U2679 (N_2679,N_2388,N_1089);
and U2680 (N_2680,N_1567,N_1543);
and U2681 (N_2681,N_1357,N_1146);
nor U2682 (N_2682,N_224,N_1764);
xor U2683 (N_2683,N_1925,N_2334);
nand U2684 (N_2684,N_2064,N_2175);
xor U2685 (N_2685,N_1976,N_1028);
nor U2686 (N_2686,N_810,N_707);
or U2687 (N_2687,N_2454,N_1733);
nand U2688 (N_2688,N_1115,N_464);
nor U2689 (N_2689,N_1491,N_1250);
or U2690 (N_2690,N_2263,N_1693);
xor U2691 (N_2691,N_161,N_2359);
nor U2692 (N_2692,N_559,N_644);
nand U2693 (N_2693,N_90,N_2242);
nand U2694 (N_2694,N_293,N_1386);
and U2695 (N_2695,N_1148,N_1888);
xor U2696 (N_2696,N_2375,N_2097);
or U2697 (N_2697,N_1528,N_2484);
xor U2698 (N_2698,N_977,N_848);
nor U2699 (N_2699,N_515,N_647);
nand U2700 (N_2700,N_980,N_1447);
and U2701 (N_2701,N_2405,N_1056);
xor U2702 (N_2702,N_2403,N_643);
nand U2703 (N_2703,N_1313,N_1817);
nor U2704 (N_2704,N_1432,N_501);
or U2705 (N_2705,N_1007,N_713);
nor U2706 (N_2706,N_920,N_98);
nand U2707 (N_2707,N_651,N_1014);
nor U2708 (N_2708,N_406,N_1006);
nor U2709 (N_2709,N_1721,N_2396);
xor U2710 (N_2710,N_41,N_1848);
nand U2711 (N_2711,N_2090,N_1046);
or U2712 (N_2712,N_492,N_683);
or U2713 (N_2713,N_450,N_1826);
nand U2714 (N_2714,N_465,N_1672);
xnor U2715 (N_2715,N_1945,N_1813);
and U2716 (N_2716,N_577,N_805);
xor U2717 (N_2717,N_754,N_2394);
or U2718 (N_2718,N_405,N_1928);
xor U2719 (N_2719,N_286,N_1618);
nand U2720 (N_2720,N_1568,N_1793);
and U2721 (N_2721,N_2117,N_345);
xor U2722 (N_2722,N_653,N_1031);
and U2723 (N_2723,N_1365,N_2122);
xor U2724 (N_2724,N_297,N_2470);
xor U2725 (N_2725,N_1217,N_1798);
xor U2726 (N_2726,N_1907,N_863);
nor U2727 (N_2727,N_2077,N_1501);
nand U2728 (N_2728,N_2110,N_1644);
or U2729 (N_2729,N_2494,N_197);
xnor U2730 (N_2730,N_200,N_85);
nand U2731 (N_2731,N_1911,N_168);
xnor U2732 (N_2732,N_1129,N_2200);
xor U2733 (N_2733,N_2397,N_1145);
nand U2734 (N_2734,N_491,N_1463);
nor U2735 (N_2735,N_1633,N_1609);
or U2736 (N_2736,N_2040,N_1999);
xor U2737 (N_2737,N_26,N_726);
xor U2738 (N_2738,N_629,N_59);
nor U2739 (N_2739,N_219,N_101);
or U2740 (N_2740,N_48,N_118);
xnor U2741 (N_2741,N_2445,N_1268);
and U2742 (N_2742,N_2100,N_872);
or U2743 (N_2743,N_354,N_1240);
xnor U2744 (N_2744,N_1916,N_1280);
or U2745 (N_2745,N_1870,N_1985);
or U2746 (N_2746,N_793,N_151);
nand U2747 (N_2747,N_301,N_1389);
or U2748 (N_2748,N_1118,N_1426);
nor U2749 (N_2749,N_1199,N_1515);
or U2750 (N_2750,N_336,N_1921);
and U2751 (N_2751,N_321,N_477);
nand U2752 (N_2752,N_1064,N_2101);
xor U2753 (N_2753,N_1675,N_720);
or U2754 (N_2754,N_1554,N_899);
nor U2755 (N_2755,N_2025,N_1032);
and U2756 (N_2756,N_1600,N_1805);
or U2757 (N_2757,N_1586,N_149);
nand U2758 (N_2758,N_1375,N_2434);
nor U2759 (N_2759,N_1411,N_702);
nand U2760 (N_2760,N_1739,N_1839);
or U2761 (N_2761,N_2053,N_1900);
nor U2762 (N_2762,N_509,N_2211);
nor U2763 (N_2763,N_1470,N_2420);
nand U2764 (N_2764,N_256,N_649);
and U2765 (N_2765,N_260,N_999);
nor U2766 (N_2766,N_989,N_1846);
xor U2767 (N_2767,N_839,N_1781);
xnor U2768 (N_2768,N_1987,N_1409);
xor U2769 (N_2769,N_2395,N_1289);
nand U2770 (N_2770,N_1910,N_851);
nor U2771 (N_2771,N_855,N_1392);
or U2772 (N_2772,N_1356,N_986);
or U2773 (N_2773,N_985,N_1514);
nand U2774 (N_2774,N_1172,N_396);
xor U2775 (N_2775,N_1134,N_2071);
nand U2776 (N_2776,N_2422,N_40);
or U2777 (N_2777,N_2353,N_1516);
nor U2778 (N_2778,N_470,N_1850);
nand U2779 (N_2779,N_1751,N_2027);
or U2780 (N_2780,N_2192,N_1161);
xor U2781 (N_2781,N_2428,N_2291);
and U2782 (N_2782,N_387,N_783);
xnor U2783 (N_2783,N_1477,N_2034);
nand U2784 (N_2784,N_641,N_1086);
or U2785 (N_2785,N_127,N_639);
nand U2786 (N_2786,N_1444,N_1445);
or U2787 (N_2787,N_1642,N_327);
or U2788 (N_2788,N_995,N_670);
or U2789 (N_2789,N_276,N_1308);
nor U2790 (N_2790,N_837,N_1082);
xnor U2791 (N_2791,N_2414,N_187);
or U2792 (N_2792,N_1252,N_1150);
and U2793 (N_2793,N_1069,N_30);
nor U2794 (N_2794,N_1092,N_889);
or U2795 (N_2795,N_263,N_2433);
or U2796 (N_2796,N_399,N_81);
nor U2797 (N_2797,N_2384,N_928);
nor U2798 (N_2798,N_880,N_1655);
xnor U2799 (N_2799,N_339,N_1020);
nor U2800 (N_2800,N_341,N_1305);
nand U2801 (N_2801,N_1459,N_2152);
xnor U2802 (N_2802,N_2284,N_791);
nor U2803 (N_2803,N_994,N_1540);
nor U2804 (N_2804,N_1591,N_1180);
nor U2805 (N_2805,N_1508,N_773);
nand U2806 (N_2806,N_2333,N_424);
and U2807 (N_2807,N_2018,N_1439);
xnor U2808 (N_2808,N_1832,N_1561);
and U2809 (N_2809,N_1228,N_731);
and U2810 (N_2810,N_1914,N_2296);
and U2811 (N_2811,N_121,N_1902);
xor U2812 (N_2812,N_1363,N_1912);
or U2813 (N_2813,N_2145,N_1712);
nor U2814 (N_2814,N_613,N_2298);
nand U2815 (N_2815,N_2148,N_292);
or U2816 (N_2816,N_2438,N_245);
or U2817 (N_2817,N_2455,N_2199);
or U2818 (N_2818,N_1083,N_598);
xnor U2819 (N_2819,N_728,N_1617);
nand U2820 (N_2820,N_792,N_1865);
and U2821 (N_2821,N_674,N_2341);
and U2822 (N_2822,N_1468,N_264);
nand U2823 (N_2823,N_1004,N_1510);
and U2824 (N_2824,N_1628,N_184);
xnor U2825 (N_2825,N_932,N_497);
or U2826 (N_2826,N_1936,N_722);
or U2827 (N_2827,N_951,N_710);
nor U2828 (N_2828,N_2038,N_2151);
xnor U2829 (N_2829,N_1222,N_663);
nor U2830 (N_2830,N_2130,N_2060);
nor U2831 (N_2831,N_2239,N_857);
nand U2832 (N_2832,N_589,N_433);
nand U2833 (N_2833,N_146,N_1637);
and U2834 (N_2834,N_2221,N_2194);
and U2835 (N_2835,N_61,N_1768);
and U2836 (N_2836,N_2431,N_2275);
nor U2837 (N_2837,N_175,N_232);
xor U2838 (N_2838,N_304,N_997);
nand U2839 (N_2839,N_2390,N_134);
nand U2840 (N_2840,N_893,N_145);
or U2841 (N_2841,N_2169,N_599);
and U2842 (N_2842,N_694,N_673);
xnor U2843 (N_2843,N_1639,N_1243);
or U2844 (N_2844,N_590,N_895);
xor U2845 (N_2845,N_2168,N_105);
nand U2846 (N_2846,N_2014,N_1160);
nand U2847 (N_2847,N_1702,N_1512);
and U2848 (N_2848,N_677,N_16);
and U2849 (N_2849,N_171,N_2265);
or U2850 (N_2850,N_2104,N_1661);
nand U2851 (N_2851,N_1562,N_102);
xor U2852 (N_2852,N_229,N_1899);
nand U2853 (N_2853,N_250,N_956);
nor U2854 (N_2854,N_1858,N_402);
nand U2855 (N_2855,N_1483,N_2);
nor U2856 (N_2856,N_471,N_2082);
xor U2857 (N_2857,N_1823,N_1533);
nor U2858 (N_2858,N_822,N_361);
nor U2859 (N_2859,N_2475,N_57);
and U2860 (N_2860,N_705,N_667);
nand U2861 (N_2861,N_952,N_1881);
or U2862 (N_2862,N_257,N_681);
xnor U2863 (N_2863,N_1288,N_708);
and U2864 (N_2864,N_2224,N_343);
nor U2865 (N_2865,N_334,N_1819);
xor U2866 (N_2866,N_894,N_1478);
nand U2867 (N_2867,N_2300,N_21);
and U2868 (N_2868,N_679,N_2084);
and U2869 (N_2869,N_824,N_2020);
nor U2870 (N_2870,N_195,N_2268);
xnor U2871 (N_2871,N_1103,N_233);
or U2872 (N_2872,N_1208,N_1627);
or U2873 (N_2873,N_314,N_867);
or U2874 (N_2874,N_1342,N_2009);
nand U2875 (N_2875,N_1276,N_1472);
nor U2876 (N_2876,N_1698,N_2035);
xnor U2877 (N_2877,N_210,N_1467);
and U2878 (N_2878,N_128,N_2280);
nor U2879 (N_2879,N_2067,N_2462);
nor U2880 (N_2880,N_2234,N_983);
or U2881 (N_2881,N_1746,N_1350);
xnor U2882 (N_2882,N_2103,N_545);
or U2883 (N_2883,N_868,N_2085);
and U2884 (N_2884,N_2189,N_1538);
xor U2885 (N_2885,N_1149,N_542);
xor U2886 (N_2886,N_1203,N_916);
nand U2887 (N_2887,N_1953,N_1460);
and U2888 (N_2888,N_124,N_374);
or U2889 (N_2889,N_10,N_1291);
nor U2890 (N_2890,N_1679,N_1373);
nor U2891 (N_2891,N_2365,N_2223);
and U2892 (N_2892,N_2437,N_95);
xnor U2893 (N_2893,N_1275,N_371);
nand U2894 (N_2894,N_1079,N_1519);
nand U2895 (N_2895,N_1789,N_1978);
nand U2896 (N_2896,N_675,N_1717);
nand U2897 (N_2897,N_750,N_821);
nand U2898 (N_2898,N_2004,N_1352);
nand U2899 (N_2899,N_1169,N_548);
xor U2900 (N_2900,N_3,N_1254);
and U2901 (N_2901,N_921,N_574);
nor U2902 (N_2902,N_692,N_646);
nand U2903 (N_2903,N_108,N_777);
or U2904 (N_2904,N_196,N_1245);
xor U2905 (N_2905,N_583,N_1299);
nand U2906 (N_2906,N_1773,N_1132);
nand U2907 (N_2907,N_1546,N_568);
xor U2908 (N_2908,N_1836,N_2051);
xor U2909 (N_2909,N_597,N_254);
nand U2910 (N_2910,N_415,N_745);
nand U2911 (N_2911,N_1957,N_1545);
nand U2912 (N_2912,N_1494,N_1716);
nor U2913 (N_2913,N_520,N_1549);
xor U2914 (N_2914,N_2446,N_1037);
nor U2915 (N_2915,N_1828,N_1473);
or U2916 (N_2916,N_91,N_1128);
or U2917 (N_2917,N_704,N_2335);
xnor U2918 (N_2918,N_392,N_1537);
xnor U2919 (N_2919,N_2215,N_630);
or U2920 (N_2920,N_2324,N_813);
nor U2921 (N_2921,N_425,N_2073);
nand U2922 (N_2922,N_1755,N_2007);
and U2923 (N_2923,N_17,N_2303);
nor U2924 (N_2924,N_688,N_517);
and U2925 (N_2925,N_481,N_2180);
or U2926 (N_2926,N_189,N_258);
xnor U2927 (N_2927,N_1689,N_1233);
nand U2928 (N_2928,N_719,N_1200);
and U2929 (N_2929,N_1230,N_14);
nand U2930 (N_2930,N_214,N_2023);
xor U2931 (N_2931,N_230,N_2493);
nand U2932 (N_2932,N_375,N_633);
nand U2933 (N_2933,N_1045,N_1792);
nand U2934 (N_2934,N_1191,N_265);
nand U2935 (N_2935,N_1758,N_1080);
nor U2936 (N_2936,N_1575,N_2269);
nand U2937 (N_2937,N_2430,N_2241);
nor U2938 (N_2938,N_906,N_2351);
nor U2939 (N_2939,N_1429,N_1290);
and U2940 (N_2940,N_2217,N_2498);
xor U2941 (N_2941,N_564,N_947);
xnor U2942 (N_2942,N_1744,N_1403);
and U2943 (N_2943,N_1523,N_205);
xor U2944 (N_2944,N_836,N_459);
nor U2945 (N_2945,N_2250,N_2166);
nand U2946 (N_2946,N_329,N_738);
nor U2947 (N_2947,N_423,N_23);
nor U2948 (N_2948,N_666,N_2355);
xnor U2949 (N_2949,N_436,N_2426);
nand U2950 (N_2950,N_1634,N_1039);
and U2951 (N_2951,N_2473,N_1862);
xor U2952 (N_2952,N_812,N_1983);
xnor U2953 (N_2953,N_496,N_900);
or U2954 (N_2954,N_32,N_1492);
and U2955 (N_2955,N_1223,N_531);
and U2956 (N_2956,N_1000,N_1414);
xor U2957 (N_2957,N_148,N_2379);
xor U2958 (N_2958,N_2195,N_2465);
and U2959 (N_2959,N_2393,N_1960);
or U2960 (N_2960,N_2163,N_915);
nor U2961 (N_2961,N_58,N_2196);
nor U2962 (N_2962,N_771,N_2456);
nor U2963 (N_2963,N_12,N_1527);
nand U2964 (N_2964,N_2362,N_2256);
and U2965 (N_2965,N_2240,N_2164);
nor U2966 (N_2966,N_1786,N_866);
and U2967 (N_2967,N_2466,N_2049);
xnor U2968 (N_2968,N_213,N_2001);
nand U2969 (N_2969,N_614,N_846);
or U2970 (N_2970,N_804,N_1038);
nand U2971 (N_2971,N_1316,N_961);
nand U2972 (N_2972,N_2057,N_2019);
nor U2973 (N_2973,N_2457,N_1246);
nand U2974 (N_2974,N_2214,N_1822);
xor U2975 (N_2975,N_2346,N_856);
or U2976 (N_2976,N_1309,N_560);
nand U2977 (N_2977,N_1859,N_1638);
nand U2978 (N_2978,N_2218,N_1162);
nor U2979 (N_2979,N_173,N_602);
xor U2980 (N_2980,N_523,N_1635);
or U2981 (N_2981,N_2135,N_2092);
nand U2982 (N_2982,N_772,N_2376);
nand U2983 (N_2983,N_2156,N_6);
and U2984 (N_2984,N_1653,N_2316);
and U2985 (N_2985,N_2061,N_645);
or U2986 (N_2986,N_690,N_2338);
nor U2987 (N_2987,N_1500,N_803);
nand U2988 (N_2988,N_1319,N_242);
nor U2989 (N_2989,N_162,N_2226);
and U2990 (N_2990,N_2089,N_1497);
nor U2991 (N_2991,N_502,N_1924);
xor U2992 (N_2992,N_2094,N_382);
nand U2993 (N_2993,N_2069,N_1152);
and U2994 (N_2994,N_2228,N_429);
nand U2995 (N_2995,N_393,N_2421);
or U2996 (N_2996,N_611,N_295);
and U2997 (N_2997,N_1142,N_1560);
nor U2998 (N_2998,N_2339,N_2401);
xnor U2999 (N_2999,N_1380,N_1284);
nand U3000 (N_3000,N_1437,N_275);
xnor U3001 (N_3001,N_2413,N_2106);
nor U3002 (N_3002,N_1674,N_394);
nand U3003 (N_3003,N_623,N_2292);
xnor U3004 (N_3004,N_2086,N_122);
or U3005 (N_3005,N_199,N_592);
nand U3006 (N_3006,N_427,N_225);
nand U3007 (N_3007,N_1743,N_288);
nor U3008 (N_3008,N_570,N_1073);
nand U3009 (N_3009,N_1050,N_2459);
nand U3010 (N_3010,N_1863,N_1745);
nand U3011 (N_3011,N_1318,N_2277);
nand U3012 (N_3012,N_2139,N_1801);
or U3013 (N_3013,N_801,N_2318);
nor U3014 (N_3014,N_1364,N_353);
and U3015 (N_3015,N_1443,N_1913);
or U3016 (N_3016,N_1582,N_403);
xnor U3017 (N_3017,N_1019,N_43);
or U3018 (N_3018,N_1269,N_2216);
nor U3019 (N_3019,N_52,N_1778);
and U3020 (N_3020,N_1507,N_74);
or U3021 (N_3021,N_1771,N_2157);
nor U3022 (N_3022,N_1372,N_1757);
xor U3023 (N_3023,N_310,N_2486);
nor U3024 (N_3024,N_736,N_1190);
nand U3025 (N_3025,N_2006,N_211);
nand U3026 (N_3026,N_207,N_1196);
nand U3027 (N_3027,N_1571,N_1495);
nor U3028 (N_3028,N_552,N_1300);
xor U3029 (N_3029,N_1423,N_1896);
or U3030 (N_3030,N_2235,N_904);
or U3031 (N_3031,N_691,N_2251);
nor U3032 (N_3032,N_1737,N_2012);
nand U3033 (N_3033,N_1067,N_2399);
or U3034 (N_3034,N_1033,N_1462);
nand U3035 (N_3035,N_1883,N_706);
or U3036 (N_3036,N_1297,N_346);
xor U3037 (N_3037,N_553,N_1615);
or U3038 (N_3038,N_1302,N_2172);
or U3039 (N_3039,N_898,N_687);
and U3040 (N_3040,N_787,N_1466);
xor U3041 (N_3041,N_1029,N_979);
and U3042 (N_3042,N_2415,N_384);
nand U3043 (N_3043,N_318,N_1643);
xnor U3044 (N_3044,N_794,N_1068);
xor U3045 (N_3045,N_1756,N_968);
or U3046 (N_3046,N_557,N_1513);
xnor U3047 (N_3047,N_938,N_2325);
or U3048 (N_3048,N_1408,N_1441);
and U3049 (N_3049,N_176,N_458);
nor U3050 (N_3050,N_718,N_1293);
and U3051 (N_3051,N_2406,N_500);
xor U3052 (N_3052,N_996,N_742);
and U3053 (N_3053,N_1903,N_1469);
nor U3054 (N_3054,N_147,N_626);
nand U3055 (N_3055,N_693,N_1315);
nor U3056 (N_3056,N_539,N_2042);
and U3057 (N_3057,N_1889,N_1893);
xnor U3058 (N_3058,N_730,N_1894);
nand U3059 (N_3059,N_860,N_2429);
and U3060 (N_3060,N_1434,N_2337);
xor U3061 (N_3061,N_807,N_2153);
xnor U3062 (N_3062,N_238,N_2309);
nor U3063 (N_3063,N_709,N_1874);
and U3064 (N_3064,N_380,N_319);
and U3065 (N_3065,N_1532,N_948);
or U3066 (N_3066,N_1908,N_584);
nor U3067 (N_3067,N_1997,N_1010);
nor U3068 (N_3068,N_316,N_2369);
nand U3069 (N_3069,N_1915,N_2232);
or U3070 (N_3070,N_266,N_404);
nor U3071 (N_3071,N_42,N_571);
xnor U3072 (N_3072,N_1927,N_25);
nor U3073 (N_3073,N_2143,N_1909);
xor U3074 (N_3074,N_1814,N_910);
nand U3075 (N_3075,N_72,N_1059);
or U3076 (N_3076,N_1645,N_1060);
nand U3077 (N_3077,N_1324,N_711);
and U3078 (N_3078,N_931,N_919);
nand U3079 (N_3079,N_1136,N_1703);
and U3080 (N_3080,N_62,N_897);
or U3081 (N_3081,N_1799,N_2144);
nand U3082 (N_3082,N_2400,N_1534);
nor U3083 (N_3083,N_84,N_69);
nand U3084 (N_3084,N_2440,N_831);
nor U3085 (N_3085,N_827,N_49);
xor U3086 (N_3086,N_1241,N_1526);
nor U3087 (N_3087,N_1742,N_1209);
xor U3088 (N_3088,N_1666,N_2345);
xnor U3089 (N_3089,N_306,N_68);
or U3090 (N_3090,N_684,N_1967);
nor U3091 (N_3091,N_2404,N_1141);
or U3092 (N_3092,N_1062,N_1518);
or U3093 (N_3093,N_764,N_516);
nand U3094 (N_3094,N_2432,N_864);
nor U3095 (N_3095,N_281,N_1176);
nor U3096 (N_3096,N_1415,N_360);
nand U3097 (N_3097,N_1102,N_2243);
nand U3098 (N_3098,N_241,N_716);
xor U3099 (N_3099,N_1189,N_1340);
or U3100 (N_3100,N_2386,N_1855);
xor U3101 (N_3101,N_528,N_1325);
nand U3102 (N_3102,N_1052,N_757);
nand U3103 (N_3103,N_2409,N_1580);
nor U3104 (N_3104,N_1860,N_1624);
nand U3105 (N_3105,N_2417,N_1656);
nor U3106 (N_3106,N_2281,N_1803);
xnor U3107 (N_3107,N_619,N_1475);
nand U3108 (N_3108,N_2044,N_1244);
nand U3109 (N_3109,N_1937,N_273);
and U3110 (N_3110,N_1336,N_1005);
xor U3111 (N_3111,N_1602,N_2146);
nor U3112 (N_3112,N_2185,N_625);
xnor U3113 (N_3113,N_1824,N_409);
or U3114 (N_3114,N_1488,N_1671);
and U3115 (N_3115,N_1078,N_1684);
xor U3116 (N_3116,N_2083,N_2411);
or U3117 (N_3117,N_418,N_356);
nor U3118 (N_3118,N_756,N_1048);
xnor U3119 (N_3119,N_2453,N_1522);
nor U3120 (N_3120,N_1456,N_1802);
nor U3121 (N_3121,N_251,N_888);
xor U3122 (N_3122,N_2076,N_678);
or U3123 (N_3123,N_2408,N_2497);
and U3124 (N_3124,N_1349,N_859);
nor U3125 (N_3125,N_270,N_896);
or U3126 (N_3126,N_2016,N_747);
nand U3127 (N_3127,N_463,N_2114);
and U3128 (N_3128,N_926,N_1074);
or U3129 (N_3129,N_201,N_1121);
or U3130 (N_3130,N_1868,N_1640);
or U3131 (N_3131,N_543,N_486);
nor U3132 (N_3132,N_2155,N_2317);
nor U3133 (N_3133,N_1766,N_1505);
nand U3134 (N_3134,N_1117,N_291);
nand U3135 (N_3135,N_1194,N_1070);
or U3136 (N_3136,N_1875,N_1366);
nand U3137 (N_3137,N_386,N_1989);
and U3138 (N_3138,N_2380,N_2313);
and U3139 (N_3139,N_657,N_73);
or U3140 (N_3140,N_1748,N_150);
and U3141 (N_3141,N_2474,N_1407);
xor U3142 (N_3142,N_2170,N_2231);
nand U3143 (N_3143,N_1929,N_1797);
xnor U3144 (N_3144,N_737,N_1607);
nand U3145 (N_3145,N_1944,N_1841);
nand U3146 (N_3146,N_538,N_50);
nand U3147 (N_3147,N_8,N_2347);
nand U3148 (N_3148,N_1857,N_1620);
nand U3149 (N_3149,N_1182,N_426);
xnor U3150 (N_3150,N_1248,N_1804);
or U3151 (N_3151,N_2439,N_1776);
nand U3152 (N_3152,N_2173,N_2021);
nor U3153 (N_3153,N_35,N_1517);
or U3154 (N_3154,N_1986,N_2307);
nor U3155 (N_3155,N_1558,N_2205);
or U3156 (N_3156,N_1759,N_1390);
or U3157 (N_3157,N_474,N_1815);
or U3158 (N_3158,N_64,N_1428);
or U3159 (N_3159,N_569,N_1890);
xnor U3160 (N_3160,N_320,N_2452);
nor U3161 (N_3161,N_1761,N_326);
nor U3162 (N_3162,N_1030,N_1347);
xnor U3163 (N_3163,N_36,N_1159);
or U3164 (N_3164,N_152,N_2201);
nor U3165 (N_3165,N_1320,N_1213);
nand U3166 (N_3166,N_781,N_1511);
xnor U3167 (N_3167,N_1930,N_160);
nor U3168 (N_3168,N_2017,N_483);
xor U3169 (N_3169,N_1780,N_352);
nor U3170 (N_3170,N_723,N_96);
xor U3171 (N_3171,N_2373,N_1931);
and U3172 (N_3172,N_1762,N_2467);
or U3173 (N_3173,N_1657,N_1791);
nand U3174 (N_3174,N_498,N_970);
or U3175 (N_3175,N_578,N_1506);
nor U3176 (N_3176,N_1662,N_1330);
nor U3177 (N_3177,N_303,N_1119);
or U3178 (N_3178,N_561,N_489);
nor U3179 (N_3179,N_82,N_634);
xor U3180 (N_3180,N_1096,N_1713);
or U3181 (N_3181,N_475,N_138);
nor U3182 (N_3182,N_1310,N_656);
xor U3183 (N_3183,N_1332,N_2087);
and U3184 (N_3184,N_1087,N_1451);
or U3185 (N_3185,N_581,N_116);
and U3186 (N_3186,N_338,N_1370);
xnor U3187 (N_3187,N_701,N_1884);
xor U3188 (N_3188,N_841,N_1621);
nand U3189 (N_3189,N_854,N_2050);
xor U3190 (N_3190,N_315,N_698);
and U3191 (N_3191,N_982,N_2312);
nor U3192 (N_3192,N_1433,N_1821);
nor U3193 (N_3193,N_1728,N_700);
or U3194 (N_3194,N_1701,N_1287);
xor U3195 (N_3195,N_2111,N_1752);
xor U3196 (N_3196,N_1729,N_550);
nand U3197 (N_3197,N_1886,N_802);
nor U3198 (N_3198,N_990,N_473);
and U3199 (N_3199,N_222,N_826);
nand U3200 (N_3200,N_1453,N_2091);
nand U3201 (N_3201,N_1126,N_112);
and U3202 (N_3202,N_268,N_1438);
nor U3203 (N_3203,N_1227,N_511);
nor U3204 (N_3204,N_2246,N_289);
nor U3205 (N_3205,N_1726,N_1397);
or U3206 (N_3206,N_959,N_1962);
or U3207 (N_3207,N_1636,N_870);
nand U3208 (N_3208,N_881,N_1168);
nand U3209 (N_3209,N_734,N_714);
xor U3210 (N_3210,N_1677,N_2330);
xor U3211 (N_3211,N_1772,N_1592);
and U3212 (N_3212,N_1975,N_929);
xor U3213 (N_3213,N_946,N_1009);
or U3214 (N_3214,N_1003,N_2202);
nor U3215 (N_3215,N_18,N_2137);
nor U3216 (N_3216,N_2149,N_249);
and U3217 (N_3217,N_1610,N_586);
or U3218 (N_3218,N_1454,N_2010);
nand U3219 (N_3219,N_435,N_75);
and U3220 (N_3220,N_1611,N_259);
nor U3221 (N_3221,N_1680,N_5);
xnor U3222 (N_3222,N_2418,N_305);
nor U3223 (N_3223,N_780,N_1174);
and U3224 (N_3224,N_699,N_671);
xnor U3225 (N_3225,N_976,N_1226);
xor U3226 (N_3226,N_998,N_840);
nor U3227 (N_3227,N_2326,N_421);
nand U3228 (N_3228,N_530,N_1192);
and U3229 (N_3229,N_1810,N_987);
or U3230 (N_3230,N_775,N_689);
xor U3231 (N_3231,N_333,N_2340);
nand U3232 (N_3232,N_909,N_1137);
nor U3233 (N_3233,N_964,N_935);
or U3234 (N_3234,N_957,N_1247);
or U3235 (N_3235,N_2206,N_2279);
and U3236 (N_3236,N_29,N_843);
xnor U3237 (N_3237,N_2276,N_1185);
or U3238 (N_3238,N_2314,N_638);
or U3239 (N_3239,N_1705,N_865);
nor U3240 (N_3240,N_1198,N_672);
nand U3241 (N_3241,N_499,N_235);
or U3242 (N_3242,N_676,N_1984);
xnor U3243 (N_3243,N_1578,N_761);
nand U3244 (N_3244,N_1735,N_1767);
or U3245 (N_3245,N_180,N_417);
or U3246 (N_3246,N_172,N_579);
xor U3247 (N_3247,N_914,N_1440);
and U3248 (N_3248,N_2058,N_2081);
or U3249 (N_3249,N_954,N_11);
and U3250 (N_3250,N_510,N_1887);
or U3251 (N_3251,N_1550,N_1843);
nor U3252 (N_3252,N_283,N_992);
and U3253 (N_3253,N_391,N_1854);
or U3254 (N_3254,N_125,N_834);
nand U3255 (N_3255,N_1139,N_113);
xnor U3256 (N_3256,N_760,N_2381);
nor U3257 (N_3257,N_2203,N_782);
and U3258 (N_3258,N_2036,N_431);
nand U3259 (N_3259,N_63,N_87);
nand U3260 (N_3260,N_1114,N_1344);
and U3261 (N_3261,N_2002,N_2209);
or U3262 (N_3262,N_165,N_778);
xor U3263 (N_3263,N_437,N_2225);
nand U3264 (N_3264,N_1207,N_2264);
and U3265 (N_3265,N_1597,N_2387);
or U3266 (N_3266,N_1553,N_1493);
and U3267 (N_3267,N_1969,N_1988);
nor U3268 (N_3268,N_284,N_1934);
or U3269 (N_3269,N_2286,N_1120);
xor U3270 (N_3270,N_901,N_33);
nor U3271 (N_3271,N_434,N_79);
nor U3272 (N_3272,N_650,N_1261);
xnor U3273 (N_3273,N_1864,N_467);
or U3274 (N_3274,N_1171,N_1667);
or U3275 (N_3275,N_2159,N_1725);
nor U3276 (N_3276,N_664,N_1842);
nand U3277 (N_3277,N_370,N_377);
xor U3278 (N_3278,N_2109,N_849);
or U3279 (N_3279,N_170,N_1895);
nor U3280 (N_3280,N_605,N_1061);
xor U3281 (N_3281,N_1820,N_2254);
nor U3282 (N_3282,N_2483,N_763);
nor U3283 (N_3283,N_163,N_2062);
xor U3284 (N_3284,N_1581,N_820);
xor U3285 (N_3285,N_1450,N_2028);
xnor U3286 (N_3286,N_1326,N_1053);
nor U3287 (N_3287,N_2382,N_2096);
nor U3288 (N_3288,N_56,N_696);
or U3289 (N_3289,N_1590,N_1219);
and U3290 (N_3290,N_137,N_1664);
xor U3291 (N_3291,N_2322,N_78);
xor U3292 (N_3292,N_1606,N_1555);
nor U3293 (N_3293,N_2045,N_1551);
xor U3294 (N_3294,N_2197,N_1322);
nand U3295 (N_3295,N_1709,N_1570);
nand U3296 (N_3296,N_349,N_451);
and U3297 (N_3297,N_1949,N_885);
and U3298 (N_3298,N_695,N_844);
or U3299 (N_3299,N_912,N_1484);
nand U3300 (N_3300,N_1294,N_1271);
xor U3301 (N_3301,N_582,N_2253);
nand U3302 (N_3302,N_365,N_749);
and U3303 (N_3303,N_565,N_1277);
and U3304 (N_3304,N_558,N_2402);
nor U3305 (N_3305,N_1183,N_1321);
and U3306 (N_3306,N_2285,N_1557);
nor U3307 (N_3307,N_1788,N_1041);
nand U3308 (N_3308,N_1085,N_355);
nor U3309 (N_3309,N_1435,N_1008);
or U3310 (N_3310,N_290,N_966);
nor U3311 (N_3311,N_2343,N_15);
nor U3312 (N_3312,N_179,N_1625);
xor U3313 (N_3313,N_2252,N_1981);
nor U3314 (N_3314,N_2024,N_1090);
nor U3315 (N_3315,N_191,N_123);
and U3316 (N_3316,N_1113,N_2272);
nor U3317 (N_3317,N_1220,N_2391);
or U3318 (N_3318,N_107,N_1235);
or U3319 (N_3319,N_1765,N_231);
xor U3320 (N_3320,N_2070,N_1775);
nand U3321 (N_3321,N_1692,N_294);
nand U3322 (N_3322,N_323,N_2008);
and U3323 (N_3323,N_2488,N_2378);
nor U3324 (N_3324,N_2193,N_117);
nand U3325 (N_3325,N_1749,N_223);
xor U3326 (N_3326,N_1806,N_2244);
xnor U3327 (N_3327,N_1387,N_1175);
nand U3328 (N_3328,N_1943,N_1151);
or U3329 (N_3329,N_1966,N_796);
nand U3330 (N_3330,N_1877,N_949);
xor U3331 (N_3331,N_1552,N_1283);
nand U3332 (N_3332,N_508,N_648);
xor U3333 (N_3333,N_240,N_660);
nand U3334 (N_3334,N_1779,N_194);
xor U3335 (N_3335,N_1938,N_2368);
xor U3336 (N_3336,N_1278,N_622);
and U3337 (N_3337,N_1094,N_34);
and U3338 (N_3338,N_39,N_1871);
and U3339 (N_3339,N_1378,N_537);
nand U3340 (N_3340,N_1777,N_282);
and U3341 (N_3341,N_1304,N_1279);
nor U3342 (N_3342,N_1027,N_2183);
nor U3343 (N_3343,N_302,N_261);
xnor U3344 (N_3344,N_799,N_1307);
nor U3345 (N_3345,N_1218,N_1669);
and U3346 (N_3346,N_1731,N_271);
nand U3347 (N_3347,N_442,N_2013);
xor U3348 (N_3348,N_1622,N_453);
nand U3349 (N_3349,N_1853,N_661);
nand U3350 (N_3350,N_1603,N_1001);
xor U3351 (N_3351,N_1576,N_830);
nand U3352 (N_3352,N_1623,N_600);
and U3353 (N_3353,N_2210,N_1156);
and U3354 (N_3354,N_2398,N_1783);
xor U3355 (N_3355,N_2160,N_1130);
nand U3356 (N_3356,N_879,N_220);
xnor U3357 (N_3357,N_1446,N_1179);
xor U3358 (N_3358,N_457,N_751);
nand U3359 (N_3359,N_616,N_908);
and U3360 (N_3360,N_925,N_526);
xor U3361 (N_3361,N_2022,N_1982);
and U3362 (N_3362,N_2112,N_1479);
nor U3363 (N_3363,N_2233,N_842);
xor U3364 (N_3364,N_115,N_567);
nor U3365 (N_3365,N_1424,N_1234);
or U3366 (N_3366,N_1270,N_443);
or U3367 (N_3367,N_1021,N_522);
nand U3368 (N_3368,N_1681,N_603);
and U3369 (N_3369,N_390,N_1065);
xor U3370 (N_3370,N_978,N_2026);
or U3371 (N_3371,N_784,N_1481);
nor U3372 (N_3372,N_2075,N_712);
nor U3373 (N_3373,N_1024,N_215);
nor U3374 (N_3374,N_1091,N_1369);
nor U3375 (N_3375,N_924,N_1125);
nor U3376 (N_3376,N_930,N_2357);
xnor U3377 (N_3377,N_407,N_324);
or U3378 (N_3378,N_1584,N_55);
or U3379 (N_3379,N_918,N_67);
or U3380 (N_3380,N_2212,N_7);
xnor U3381 (N_3381,N_887,N_1328);
nand U3382 (N_3382,N_485,N_2011);
nor U3383 (N_3383,N_1116,N_984);
nor U3384 (N_3384,N_2492,N_1849);
or U3385 (N_3385,N_247,N_280);
nor U3386 (N_3386,N_1489,N_2481);
nor U3387 (N_3387,N_823,N_1700);
nand U3388 (N_3388,N_198,N_1498);
or U3389 (N_3389,N_1940,N_337);
nand U3390 (N_3390,N_2134,N_2186);
or U3391 (N_3391,N_1670,N_1013);
nand U3392 (N_3392,N_746,N_2472);
xnor U3393 (N_3393,N_1996,N_2308);
or U3394 (N_3394,N_236,N_2142);
xor U3395 (N_3395,N_1876,N_795);
nand U3396 (N_3396,N_1918,N_1629);
nor U3397 (N_3397,N_1394,N_2048);
or U3398 (N_3398,N_2136,N_104);
nor U3399 (N_3399,N_142,N_2261);
or U3400 (N_3400,N_1259,N_279);
xor U3401 (N_3401,N_1867,N_2124);
xor U3402 (N_3402,N_937,N_395);
nor U3403 (N_3403,N_1612,N_369);
nor U3404 (N_3404,N_1845,N_1919);
xor U3405 (N_3405,N_886,N_1954);
or U3406 (N_3406,N_381,N_311);
nor U3407 (N_3407,N_212,N_862);
and U3408 (N_3408,N_1044,N_342);
nor U3409 (N_3409,N_1047,N_1572);
and U3410 (N_3410,N_1991,N_1077);
and U3411 (N_3411,N_1388,N_164);
nor U3412 (N_3412,N_1521,N_917);
nor U3413 (N_3413,N_157,N_1109);
or U3414 (N_3414,N_1490,N_2133);
nand U3415 (N_3415,N_878,N_480);
nand U3416 (N_3416,N_1727,N_1237);
xnor U3417 (N_3417,N_1593,N_1730);
xnor U3418 (N_3418,N_2257,N_874);
nand U3419 (N_3419,N_2289,N_873);
nand U3420 (N_3420,N_1017,N_1311);
or U3421 (N_3421,N_2247,N_1127);
xnor U3422 (N_3422,N_1272,N_1547);
nand U3423 (N_3423,N_1417,N_2078);
and U3424 (N_3424,N_2177,N_110);
nand U3425 (N_3425,N_1099,N_1327);
or U3426 (N_3426,N_1410,N_47);
nor U3427 (N_3427,N_753,N_618);
and U3428 (N_3428,N_243,N_1598);
xor U3429 (N_3429,N_312,N_385);
xnor U3430 (N_3430,N_1676,N_153);
and U3431 (N_3431,N_109,N_1830);
nand U3432 (N_3432,N_1427,N_2041);
nand U3433 (N_3433,N_1338,N_2181);
and U3434 (N_3434,N_850,N_740);
or U3435 (N_3435,N_1418,N_2176);
xor U3436 (N_3436,N_575,N_77);
nand U3437 (N_3437,N_272,N_554);
xnor U3438 (N_3438,N_2108,N_697);
xnor U3439 (N_3439,N_325,N_227);
and U3440 (N_3440,N_2132,N_1258);
nor U3441 (N_3441,N_2208,N_744);
nand U3442 (N_3442,N_852,N_1782);
and U3443 (N_3443,N_1158,N_1496);
xnor U3444 (N_3444,N_2204,N_2336);
nand U3445 (N_3445,N_1257,N_940);
and U3446 (N_3446,N_769,N_86);
nand U3447 (N_3447,N_156,N_2072);
and U3448 (N_3448,N_1382,N_551);
or U3449 (N_3449,N_1323,N_2138);
or U3450 (N_3450,N_9,N_609);
nand U3451 (N_3451,N_546,N_317);
xor U3452 (N_3452,N_1840,N_621);
nand U3453 (N_3453,N_503,N_533);
nand U3454 (N_3454,N_2306,N_1108);
nand U3455 (N_3455,N_476,N_132);
or U3456 (N_3456,N_1040,N_2441);
xnor U3457 (N_3457,N_478,N_606);
or U3458 (N_3458,N_129,N_1663);
xnor U3459 (N_3459,N_1690,N_743);
and U3460 (N_3460,N_1458,N_892);
nand U3461 (N_3461,N_832,N_933);
or U3462 (N_3462,N_1574,N_654);
or U3463 (N_3463,N_1097,N_2461);
and U3464 (N_3464,N_1577,N_65);
nor U3465 (N_3465,N_351,N_1022);
nor U3466 (N_3466,N_1594,N_1652);
or U3467 (N_3467,N_1333,N_373);
nand U3468 (N_3468,N_1935,N_922);
and U3469 (N_3469,N_1106,N_913);
nand U3470 (N_3470,N_479,N_903);
and U3471 (N_3471,N_816,N_636);
or U3472 (N_3472,N_1616,N_208);
and U3473 (N_3473,N_141,N_397);
xor U3474 (N_3474,N_106,N_2356);
and U3475 (N_3475,N_1891,N_974);
xor U3476 (N_3476,N_2039,N_1054);
nor U3477 (N_3477,N_2447,N_1154);
or U3478 (N_3478,N_328,N_1147);
xnor U3479 (N_3479,N_4,N_1829);
nor U3480 (N_3480,N_1486,N_911);
nor U3481 (N_3481,N_493,N_1301);
and U3482 (N_3482,N_1055,N_1153);
xnor U3483 (N_3483,N_972,N_1449);
or U3484 (N_3484,N_939,N_100);
and U3485 (N_3485,N_448,N_357);
and U3486 (N_3486,N_1564,N_1947);
nor U3487 (N_3487,N_1998,N_1361);
nor U3488 (N_3488,N_1239,N_1253);
nand U3489 (N_3489,N_2328,N_1419);
and U3490 (N_3490,N_682,N_725);
or U3491 (N_3491,N_1436,N_934);
xnor U3492 (N_3492,N_1398,N_1002);
or U3493 (N_3493,N_1585,N_593);
xor U3494 (N_3494,N_1687,N_1358);
nor U3495 (N_3495,N_359,N_758);
and U3496 (N_3496,N_2412,N_1818);
xor U3497 (N_3497,N_2342,N_2179);
and U3498 (N_3498,N_439,N_1166);
nand U3499 (N_3499,N_1619,N_2311);
and U3500 (N_3500,N_1385,N_1416);
or U3501 (N_3501,N_1683,N_1964);
xor U3502 (N_3502,N_1897,N_1973);
nand U3503 (N_3503,N_733,N_1869);
and U3504 (N_3504,N_1262,N_1143);
nand U3505 (N_3505,N_366,N_884);
and U3506 (N_3506,N_1682,N_70);
or U3507 (N_3507,N_2449,N_1135);
xnor U3508 (N_3508,N_766,N_1098);
xor U3509 (N_3509,N_1787,N_1794);
and U3510 (N_3510,N_1901,N_2227);
nand U3511 (N_3511,N_1374,N_521);
or U3512 (N_3512,N_2105,N_2361);
or U3513 (N_3513,N_1691,N_752);
or U3514 (N_3514,N_344,N_2352);
and U3515 (N_3515,N_788,N_2370);
nor U3516 (N_3516,N_936,N_1504);
and U3517 (N_3517,N_2098,N_136);
and U3518 (N_3518,N_1476,N_2463);
xnor U3519 (N_3519,N_1708,N_809);
xnor U3520 (N_3520,N_1383,N_505);
nor U3521 (N_3521,N_53,N_2320);
nor U3522 (N_3522,N_1941,N_2331);
nand U3523 (N_3523,N_825,N_845);
or U3524 (N_3524,N_2187,N_958);
and U3525 (N_3525,N_2469,N_155);
and U3526 (N_3526,N_1951,N_1530);
nand U3527 (N_3527,N_447,N_1431);
nand U3528 (N_3528,N_869,N_1979);
nor U3529 (N_3529,N_1355,N_2230);
xnor U3530 (N_3530,N_27,N_642);
xor U3531 (N_3531,N_2213,N_1882);
nor U3532 (N_3532,N_2319,N_1);
and U3533 (N_3533,N_612,N_1396);
nor U3534 (N_3534,N_452,N_182);
nand U3535 (N_3535,N_206,N_883);
xnor U3536 (N_3536,N_193,N_1760);
and U3537 (N_3537,N_2115,N_858);
and U3538 (N_3538,N_1811,N_1838);
and U3539 (N_3539,N_668,N_2499);
xnor U3540 (N_3540,N_566,N_416);
nor U3541 (N_3541,N_1579,N_1144);
and U3542 (N_3542,N_529,N_414);
xor U3543 (N_3543,N_2052,N_441);
nand U3544 (N_3544,N_1448,N_1303);
xor U3545 (N_3545,N_330,N_1354);
or U3546 (N_3546,N_1093,N_962);
or U3547 (N_3547,N_1704,N_1404);
or U3548 (N_3548,N_19,N_1391);
nand U3549 (N_3549,N_188,N_2424);
xnor U3550 (N_3550,N_1395,N_1524);
nor U3551 (N_3551,N_1542,N_1425);
nand U3552 (N_3552,N_2121,N_1112);
nor U3553 (N_3553,N_111,N_1095);
or U3554 (N_3554,N_556,N_601);
nand U3555 (N_3555,N_2147,N_428);
or U3556 (N_3556,N_1774,N_2003);
and U3557 (N_3557,N_2056,N_2079);
nor U3558 (N_3558,N_313,N_620);
nand U3559 (N_3559,N_905,N_1430);
nor U3560 (N_3560,N_1898,N_632);
xor U3561 (N_3561,N_1353,N_487);
or U3562 (N_3562,N_1256,N_1825);
or U3563 (N_3563,N_204,N_1785);
nand U3564 (N_3564,N_190,N_1892);
xor U3565 (N_3565,N_907,N_1016);
and U3566 (N_3566,N_1215,N_2419);
nor U3567 (N_3567,N_806,N_1795);
xor U3568 (N_3568,N_203,N_430);
xnor U3569 (N_3569,N_2360,N_563);
or U3570 (N_3570,N_383,N_1738);
xor U3571 (N_3571,N_1632,N_2478);
nand U3572 (N_3572,N_1807,N_2374);
nor U3573 (N_3573,N_768,N_1312);
xnor U3574 (N_3574,N_2059,N_484);
and U3575 (N_3575,N_274,N_585);
and U3576 (N_3576,N_221,N_1880);
nor U3577 (N_3577,N_1084,N_1763);
nor U3578 (N_3578,N_580,N_1264);
nand U3579 (N_3579,N_808,N_1076);
and U3580 (N_3580,N_2367,N_1011);
and U3581 (N_3581,N_2425,N_631);
nand U3582 (N_3582,N_960,N_1296);
or U3583 (N_3583,N_46,N_1138);
or U3584 (N_3584,N_1715,N_2125);
xnor U3585 (N_3585,N_2480,N_955);
or U3586 (N_3586,N_2283,N_76);
nor U3587 (N_3587,N_724,N_1769);
nor U3588 (N_3588,N_1525,N_652);
and U3589 (N_3589,N_953,N_490);
xnor U3590 (N_3590,N_2174,N_1242);
and U3591 (N_3591,N_2442,N_2458);
nor U3592 (N_3592,N_347,N_877);
and U3593 (N_3593,N_1025,N_1485);
and U3594 (N_3594,N_186,N_45);
or U3595 (N_3595,N_255,N_1688);
or U3596 (N_3596,N_1831,N_1216);
xor U3597 (N_3597,N_2270,N_790);
xor U3598 (N_3598,N_1932,N_2043);
nor U3599 (N_3599,N_514,N_2236);
nor U3600 (N_3600,N_993,N_525);
and U3601 (N_3601,N_549,N_1608);
nor U3602 (N_3602,N_1195,N_51);
and U3603 (N_3603,N_454,N_119);
or U3604 (N_3604,N_192,N_144);
nor U3605 (N_3605,N_400,N_114);
or U3606 (N_3606,N_1249,N_358);
or U3607 (N_3607,N_2113,N_2188);
nand U3608 (N_3608,N_2063,N_1685);
or U3609 (N_3609,N_1658,N_2427);
and U3610 (N_3610,N_617,N_1075);
or U3611 (N_3611,N_1630,N_2451);
xnor U3612 (N_3612,N_1406,N_217);
or U3613 (N_3613,N_461,N_1837);
nor U3614 (N_3614,N_1923,N_1796);
nand U3615 (N_3615,N_2344,N_941);
nand U3616 (N_3616,N_1536,N_2128);
nor U3617 (N_3617,N_1337,N_2037);
or U3618 (N_3618,N_1026,N_2066);
nor U3619 (N_3619,N_594,N_1057);
nand U3620 (N_3620,N_1471,N_1565);
nand U3621 (N_3621,N_536,N_637);
nand U3622 (N_3622,N_244,N_1531);
xor U3623 (N_3623,N_2435,N_2207);
nor U3624 (N_3624,N_2416,N_1650);
nand U3625 (N_3625,N_267,N_2350);
nand U3626 (N_3626,N_1371,N_401);
nor U3627 (N_3627,N_1990,N_555);
nand U3628 (N_3628,N_1718,N_659);
or U3629 (N_3629,N_1659,N_2191);
xnor U3630 (N_3630,N_1267,N_449);
nand U3631 (N_3631,N_703,N_2321);
xnor U3632 (N_3632,N_1229,N_0);
xor U3633 (N_3633,N_1833,N_963);
and U3634 (N_3634,N_504,N_2371);
nor U3635 (N_3635,N_1678,N_1856);
nor U3636 (N_3636,N_2489,N_2088);
and U3637 (N_3637,N_218,N_797);
or U3638 (N_3638,N_278,N_1952);
xnor U3639 (N_3639,N_1631,N_1184);
nand U3640 (N_3640,N_2327,N_1946);
or U3641 (N_3641,N_1878,N_2167);
nand U3642 (N_3642,N_335,N_975);
and U3643 (N_3643,N_166,N_669);
xnor U3644 (N_3644,N_1402,N_2410);
xor U3645 (N_3645,N_786,N_1905);
or U3646 (N_3646,N_93,N_2305);
nand U3647 (N_3647,N_1377,N_739);
and U3648 (N_3648,N_31,N_2485);
and U3649 (N_3649,N_1197,N_248);
and U3650 (N_3650,N_1665,N_388);
nand U3651 (N_3651,N_828,N_1535);
or U3652 (N_3652,N_1348,N_202);
nand U3653 (N_3653,N_1205,N_2301);
nor U3654 (N_3654,N_1212,N_2029);
and U3655 (N_3655,N_662,N_524);
or U3656 (N_3656,N_595,N_1614);
xor U3657 (N_3657,N_1421,N_126);
nor U3658 (N_3658,N_748,N_1695);
and U3659 (N_3659,N_1186,N_1457);
nand U3660 (N_3660,N_2490,N_765);
xor U3661 (N_3661,N_532,N_2482);
and U3662 (N_3662,N_1950,N_1104);
nand U3663 (N_3663,N_133,N_2323);
xor U3664 (N_3664,N_22,N_1920);
nor U3665 (N_3665,N_1649,N_1722);
and U3666 (N_3666,N_1164,N_1808);
nand U3667 (N_3667,N_1359,N_38);
nor U3668 (N_3668,N_2290,N_1464);
xor U3669 (N_3669,N_226,N_2162);
and U3670 (N_3670,N_1331,N_1955);
or U3671 (N_3671,N_1844,N_1686);
or U3672 (N_3672,N_2423,N_1163);
nor U3673 (N_3673,N_2161,N_1214);
nand U3674 (N_3674,N_239,N_2032);
xor U3675 (N_3675,N_2495,N_277);
xnor U3676 (N_3676,N_891,N_1573);
or U3677 (N_3677,N_1719,N_1503);
nor U3678 (N_3678,N_1939,N_44);
nand U3679 (N_3679,N_340,N_140);
or U3680 (N_3680,N_1502,N_455);
and U3681 (N_3681,N_1042,N_735);
or U3682 (N_3682,N_2471,N_228);
nand U3683 (N_3683,N_835,N_1177);
nor U3684 (N_3684,N_971,N_902);
xnor U3685 (N_3685,N_944,N_1231);
or U3686 (N_3686,N_1360,N_307);
nand U3687 (N_3687,N_37,N_1613);
and U3688 (N_3688,N_1904,N_1210);
xnor U3689 (N_3689,N_331,N_332);
and U3690 (N_3690,N_2299,N_420);
nor U3691 (N_3691,N_1051,N_527);
nor U3692 (N_3692,N_398,N_181);
nand U3693 (N_3693,N_721,N_1131);
nor U3694 (N_3694,N_1847,N_1043);
nand U3695 (N_3695,N_512,N_1696);
xnor U3696 (N_3696,N_1049,N_1105);
and U3697 (N_3697,N_2349,N_234);
and U3698 (N_3698,N_2450,N_1224);
nor U3699 (N_3699,N_833,N_1071);
xor U3700 (N_3700,N_1122,N_2107);
or U3701 (N_3701,N_818,N_2348);
nand U3702 (N_3702,N_1959,N_1971);
nor U3703 (N_3703,N_2287,N_2295);
nor U3704 (N_3704,N_363,N_2288);
nand U3705 (N_3705,N_1035,N_1263);
nand U3706 (N_3706,N_2222,N_1926);
nor U3707 (N_3707,N_2065,N_1058);
nand U3708 (N_3708,N_1399,N_1367);
nor U3709 (N_3709,N_1023,N_2407);
nor U3710 (N_3710,N_1286,N_1968);
nand U3711 (N_3711,N_1673,N_1604);
or U3712 (N_3712,N_1583,N_628);
xnor U3713 (N_3713,N_1034,N_99);
and U3714 (N_3714,N_120,N_847);
nor U3715 (N_3715,N_540,N_817);
and U3716 (N_3716,N_460,N_1345);
nor U3717 (N_3717,N_798,N_1265);
or U3718 (N_3718,N_1306,N_183);
nand U3719 (N_3719,N_1992,N_2389);
nand U3720 (N_3720,N_1140,N_1544);
xnor U3721 (N_3721,N_103,N_1651);
or U3722 (N_3722,N_2487,N_562);
and U3723 (N_3723,N_1885,N_1852);
nand U3724 (N_3724,N_1072,N_1018);
xnor U3725 (N_3725,N_627,N_2005);
nor U3726 (N_3726,N_1605,N_1413);
xor U3727 (N_3727,N_298,N_92);
nor U3728 (N_3728,N_2000,N_2055);
nor U3729 (N_3729,N_2460,N_2377);
nand U3730 (N_3730,N_1232,N_1800);
and U3731 (N_3731,N_1724,N_408);
nor U3732 (N_3732,N_174,N_1285);
or U3733 (N_3733,N_507,N_13);
or U3734 (N_3734,N_2095,N_139);
or U3735 (N_3735,N_1974,N_1736);
and U3736 (N_3736,N_1595,N_2178);
and U3737 (N_3737,N_1596,N_209);
nand U3738 (N_3738,N_2259,N_2033);
nor U3739 (N_3739,N_1292,N_1866);
or U3740 (N_3740,N_362,N_1660);
or U3741 (N_3741,N_800,N_287);
nand U3742 (N_3742,N_432,N_2448);
nor U3743 (N_3743,N_1298,N_1362);
or U3744 (N_3744,N_2245,N_2229);
nor U3745 (N_3745,N_1646,N_1972);
and U3746 (N_3746,N_973,N_2171);
xnor U3747 (N_3747,N_1587,N_2219);
nand U3748 (N_3748,N_1588,N_785);
and U3749 (N_3749,N_1487,N_1648);
and U3750 (N_3750,N_1822,N_98);
xnor U3751 (N_3751,N_2135,N_479);
and U3752 (N_3752,N_252,N_870);
or U3753 (N_3753,N_278,N_581);
nand U3754 (N_3754,N_435,N_190);
nor U3755 (N_3755,N_1284,N_651);
or U3756 (N_3756,N_856,N_2138);
or U3757 (N_3757,N_446,N_2262);
and U3758 (N_3758,N_1772,N_1146);
xor U3759 (N_3759,N_183,N_1778);
and U3760 (N_3760,N_1017,N_2445);
nor U3761 (N_3761,N_519,N_1245);
or U3762 (N_3762,N_252,N_425);
and U3763 (N_3763,N_821,N_216);
or U3764 (N_3764,N_1673,N_109);
xor U3765 (N_3765,N_607,N_573);
xor U3766 (N_3766,N_1606,N_2405);
or U3767 (N_3767,N_1472,N_436);
and U3768 (N_3768,N_824,N_1428);
nor U3769 (N_3769,N_1956,N_1210);
nor U3770 (N_3770,N_2229,N_233);
nand U3771 (N_3771,N_187,N_916);
or U3772 (N_3772,N_2422,N_450);
nand U3773 (N_3773,N_450,N_456);
nor U3774 (N_3774,N_1831,N_259);
or U3775 (N_3775,N_1789,N_1477);
and U3776 (N_3776,N_1078,N_55);
nor U3777 (N_3777,N_2200,N_2196);
nand U3778 (N_3778,N_1194,N_1154);
nand U3779 (N_3779,N_1106,N_717);
and U3780 (N_3780,N_1753,N_388);
or U3781 (N_3781,N_565,N_1498);
or U3782 (N_3782,N_1467,N_2273);
nand U3783 (N_3783,N_933,N_2101);
or U3784 (N_3784,N_2003,N_479);
xor U3785 (N_3785,N_2264,N_2005);
nand U3786 (N_3786,N_1510,N_2342);
nand U3787 (N_3787,N_638,N_1518);
and U3788 (N_3788,N_1635,N_2244);
and U3789 (N_3789,N_1999,N_227);
nor U3790 (N_3790,N_1605,N_1807);
nand U3791 (N_3791,N_790,N_365);
xor U3792 (N_3792,N_1491,N_1509);
or U3793 (N_3793,N_1525,N_1402);
or U3794 (N_3794,N_41,N_364);
and U3795 (N_3795,N_460,N_1483);
or U3796 (N_3796,N_561,N_2292);
xnor U3797 (N_3797,N_745,N_1513);
nor U3798 (N_3798,N_2084,N_592);
and U3799 (N_3799,N_2224,N_202);
and U3800 (N_3800,N_1345,N_425);
and U3801 (N_3801,N_2031,N_301);
nand U3802 (N_3802,N_2193,N_192);
nand U3803 (N_3803,N_1719,N_1589);
nor U3804 (N_3804,N_873,N_1781);
or U3805 (N_3805,N_2147,N_140);
nor U3806 (N_3806,N_1574,N_1865);
nand U3807 (N_3807,N_2468,N_1607);
or U3808 (N_3808,N_322,N_501);
nor U3809 (N_3809,N_1840,N_14);
and U3810 (N_3810,N_361,N_1437);
nand U3811 (N_3811,N_1942,N_1746);
nand U3812 (N_3812,N_1593,N_1774);
nor U3813 (N_3813,N_2267,N_1791);
or U3814 (N_3814,N_1314,N_400);
nor U3815 (N_3815,N_792,N_868);
nand U3816 (N_3816,N_1358,N_1655);
nand U3817 (N_3817,N_1626,N_1656);
nand U3818 (N_3818,N_637,N_1280);
nor U3819 (N_3819,N_712,N_2326);
nand U3820 (N_3820,N_1968,N_1309);
nor U3821 (N_3821,N_1918,N_186);
and U3822 (N_3822,N_494,N_310);
and U3823 (N_3823,N_539,N_2005);
nand U3824 (N_3824,N_1390,N_245);
and U3825 (N_3825,N_714,N_2306);
xnor U3826 (N_3826,N_1413,N_2138);
nand U3827 (N_3827,N_1847,N_2049);
nand U3828 (N_3828,N_1419,N_772);
nand U3829 (N_3829,N_2187,N_1777);
nor U3830 (N_3830,N_2451,N_1937);
nor U3831 (N_3831,N_197,N_1241);
nand U3832 (N_3832,N_1101,N_1347);
or U3833 (N_3833,N_2428,N_650);
xnor U3834 (N_3834,N_1922,N_2108);
nor U3835 (N_3835,N_1805,N_283);
nand U3836 (N_3836,N_769,N_127);
or U3837 (N_3837,N_1112,N_795);
and U3838 (N_3838,N_1758,N_2123);
xor U3839 (N_3839,N_606,N_317);
or U3840 (N_3840,N_1062,N_2059);
nand U3841 (N_3841,N_2200,N_407);
nor U3842 (N_3842,N_598,N_2397);
nor U3843 (N_3843,N_398,N_169);
or U3844 (N_3844,N_2394,N_1207);
nand U3845 (N_3845,N_851,N_396);
nor U3846 (N_3846,N_325,N_2456);
nor U3847 (N_3847,N_455,N_447);
and U3848 (N_3848,N_2333,N_2437);
xor U3849 (N_3849,N_1197,N_938);
xor U3850 (N_3850,N_1243,N_1274);
or U3851 (N_3851,N_793,N_1547);
or U3852 (N_3852,N_1891,N_882);
or U3853 (N_3853,N_1958,N_2470);
and U3854 (N_3854,N_533,N_1991);
xnor U3855 (N_3855,N_482,N_1013);
xnor U3856 (N_3856,N_2197,N_739);
and U3857 (N_3857,N_1002,N_518);
and U3858 (N_3858,N_1562,N_388);
xor U3859 (N_3859,N_633,N_1599);
or U3860 (N_3860,N_1549,N_1317);
nor U3861 (N_3861,N_777,N_1340);
xor U3862 (N_3862,N_382,N_132);
or U3863 (N_3863,N_580,N_2032);
xor U3864 (N_3864,N_2479,N_1048);
nor U3865 (N_3865,N_971,N_613);
and U3866 (N_3866,N_1691,N_883);
and U3867 (N_3867,N_1314,N_1575);
nand U3868 (N_3868,N_699,N_2240);
and U3869 (N_3869,N_1315,N_1180);
xnor U3870 (N_3870,N_1796,N_1875);
xor U3871 (N_3871,N_583,N_396);
nand U3872 (N_3872,N_1679,N_2369);
or U3873 (N_3873,N_1961,N_1126);
nor U3874 (N_3874,N_701,N_721);
nor U3875 (N_3875,N_184,N_2370);
or U3876 (N_3876,N_1001,N_1595);
and U3877 (N_3877,N_2112,N_1230);
and U3878 (N_3878,N_1561,N_2073);
nand U3879 (N_3879,N_2208,N_1873);
nor U3880 (N_3880,N_739,N_2263);
nor U3881 (N_3881,N_78,N_462);
and U3882 (N_3882,N_1478,N_2337);
xnor U3883 (N_3883,N_870,N_1730);
and U3884 (N_3884,N_486,N_260);
nand U3885 (N_3885,N_1964,N_1653);
or U3886 (N_3886,N_1268,N_2216);
xnor U3887 (N_3887,N_795,N_406);
nor U3888 (N_3888,N_206,N_409);
nand U3889 (N_3889,N_1412,N_246);
xor U3890 (N_3890,N_198,N_2470);
and U3891 (N_3891,N_840,N_1748);
or U3892 (N_3892,N_1145,N_904);
nand U3893 (N_3893,N_1409,N_2336);
nor U3894 (N_3894,N_391,N_251);
nor U3895 (N_3895,N_1426,N_2272);
nand U3896 (N_3896,N_324,N_2184);
nand U3897 (N_3897,N_342,N_206);
nand U3898 (N_3898,N_1161,N_1449);
xor U3899 (N_3899,N_2199,N_1);
or U3900 (N_3900,N_1223,N_385);
nor U3901 (N_3901,N_1298,N_1991);
nand U3902 (N_3902,N_894,N_320);
nor U3903 (N_3903,N_1696,N_2189);
xnor U3904 (N_3904,N_2068,N_88);
nand U3905 (N_3905,N_909,N_1640);
and U3906 (N_3906,N_2049,N_2192);
or U3907 (N_3907,N_1524,N_1322);
nor U3908 (N_3908,N_1498,N_1999);
nand U3909 (N_3909,N_2251,N_1900);
and U3910 (N_3910,N_2190,N_1279);
or U3911 (N_3911,N_757,N_106);
nand U3912 (N_3912,N_280,N_2069);
nor U3913 (N_3913,N_1474,N_1273);
nand U3914 (N_3914,N_2447,N_2202);
xor U3915 (N_3915,N_1691,N_1672);
nor U3916 (N_3916,N_730,N_1870);
or U3917 (N_3917,N_2355,N_2157);
nor U3918 (N_3918,N_1724,N_1197);
nor U3919 (N_3919,N_807,N_921);
and U3920 (N_3920,N_1519,N_347);
and U3921 (N_3921,N_420,N_418);
or U3922 (N_3922,N_1020,N_489);
nand U3923 (N_3923,N_398,N_2355);
nor U3924 (N_3924,N_1016,N_2309);
nand U3925 (N_3925,N_1071,N_614);
nor U3926 (N_3926,N_2126,N_1455);
nand U3927 (N_3927,N_535,N_2414);
nor U3928 (N_3928,N_2059,N_1139);
xor U3929 (N_3929,N_2303,N_542);
nor U3930 (N_3930,N_1865,N_143);
nand U3931 (N_3931,N_2256,N_1601);
xor U3932 (N_3932,N_960,N_968);
nor U3933 (N_3933,N_1060,N_2086);
nor U3934 (N_3934,N_2272,N_1883);
and U3935 (N_3935,N_410,N_2448);
nand U3936 (N_3936,N_1633,N_650);
xnor U3937 (N_3937,N_556,N_1017);
and U3938 (N_3938,N_543,N_1959);
or U3939 (N_3939,N_728,N_199);
and U3940 (N_3940,N_369,N_1984);
xnor U3941 (N_3941,N_353,N_1135);
and U3942 (N_3942,N_1076,N_1340);
xor U3943 (N_3943,N_1296,N_2251);
or U3944 (N_3944,N_2025,N_142);
nand U3945 (N_3945,N_2470,N_2491);
or U3946 (N_3946,N_1976,N_310);
xor U3947 (N_3947,N_277,N_1899);
nand U3948 (N_3948,N_1288,N_1908);
xor U3949 (N_3949,N_436,N_1652);
nor U3950 (N_3950,N_1225,N_1728);
or U3951 (N_3951,N_182,N_1073);
xor U3952 (N_3952,N_926,N_1091);
xnor U3953 (N_3953,N_1307,N_1528);
xor U3954 (N_3954,N_1259,N_633);
nor U3955 (N_3955,N_2208,N_1667);
xnor U3956 (N_3956,N_1338,N_558);
nand U3957 (N_3957,N_1520,N_811);
and U3958 (N_3958,N_57,N_806);
nor U3959 (N_3959,N_1898,N_746);
or U3960 (N_3960,N_523,N_699);
or U3961 (N_3961,N_1940,N_569);
or U3962 (N_3962,N_195,N_735);
xnor U3963 (N_3963,N_1071,N_1816);
and U3964 (N_3964,N_406,N_1847);
nand U3965 (N_3965,N_532,N_59);
nor U3966 (N_3966,N_2486,N_868);
and U3967 (N_3967,N_1815,N_2274);
nand U3968 (N_3968,N_850,N_511);
xor U3969 (N_3969,N_1686,N_2439);
nor U3970 (N_3970,N_1,N_812);
xor U3971 (N_3971,N_660,N_1645);
nor U3972 (N_3972,N_468,N_2017);
xnor U3973 (N_3973,N_2380,N_1786);
nand U3974 (N_3974,N_1340,N_0);
nand U3975 (N_3975,N_805,N_1299);
and U3976 (N_3976,N_1448,N_1660);
or U3977 (N_3977,N_263,N_2112);
nor U3978 (N_3978,N_1896,N_1949);
nand U3979 (N_3979,N_264,N_1663);
nand U3980 (N_3980,N_2176,N_1037);
nand U3981 (N_3981,N_1245,N_2269);
xor U3982 (N_3982,N_2349,N_1722);
nand U3983 (N_3983,N_1569,N_1935);
and U3984 (N_3984,N_1991,N_1401);
and U3985 (N_3985,N_2260,N_296);
nor U3986 (N_3986,N_2023,N_316);
or U3987 (N_3987,N_1807,N_1226);
or U3988 (N_3988,N_1243,N_2020);
or U3989 (N_3989,N_2439,N_1718);
and U3990 (N_3990,N_2367,N_2234);
xnor U3991 (N_3991,N_825,N_668);
xor U3992 (N_3992,N_1204,N_1101);
nand U3993 (N_3993,N_2035,N_1399);
nand U3994 (N_3994,N_1155,N_2429);
xnor U3995 (N_3995,N_141,N_2323);
or U3996 (N_3996,N_1029,N_34);
xor U3997 (N_3997,N_1618,N_2040);
or U3998 (N_3998,N_276,N_2290);
nand U3999 (N_3999,N_1104,N_838);
and U4000 (N_4000,N_1159,N_1708);
and U4001 (N_4001,N_1818,N_1547);
xor U4002 (N_4002,N_723,N_1693);
or U4003 (N_4003,N_69,N_2039);
nand U4004 (N_4004,N_1936,N_816);
or U4005 (N_4005,N_1357,N_1852);
nand U4006 (N_4006,N_1074,N_1844);
nand U4007 (N_4007,N_1883,N_981);
xnor U4008 (N_4008,N_1135,N_1742);
nand U4009 (N_4009,N_302,N_274);
and U4010 (N_4010,N_396,N_1146);
nor U4011 (N_4011,N_414,N_947);
xor U4012 (N_4012,N_1487,N_700);
or U4013 (N_4013,N_954,N_1718);
or U4014 (N_4014,N_220,N_483);
nor U4015 (N_4015,N_1972,N_2280);
nand U4016 (N_4016,N_234,N_2306);
or U4017 (N_4017,N_1399,N_1455);
nor U4018 (N_4018,N_922,N_1092);
nor U4019 (N_4019,N_110,N_104);
nor U4020 (N_4020,N_106,N_288);
nand U4021 (N_4021,N_2448,N_1937);
or U4022 (N_4022,N_556,N_1808);
nand U4023 (N_4023,N_356,N_2173);
and U4024 (N_4024,N_934,N_194);
nand U4025 (N_4025,N_1549,N_909);
nand U4026 (N_4026,N_1661,N_387);
or U4027 (N_4027,N_103,N_33);
xnor U4028 (N_4028,N_449,N_1342);
nand U4029 (N_4029,N_1871,N_2169);
nand U4030 (N_4030,N_125,N_2208);
and U4031 (N_4031,N_1124,N_2332);
xnor U4032 (N_4032,N_2014,N_1056);
nand U4033 (N_4033,N_1593,N_960);
nand U4034 (N_4034,N_393,N_1785);
nor U4035 (N_4035,N_2249,N_824);
and U4036 (N_4036,N_774,N_1402);
and U4037 (N_4037,N_2045,N_699);
nand U4038 (N_4038,N_855,N_1598);
or U4039 (N_4039,N_2260,N_1404);
xor U4040 (N_4040,N_2240,N_1233);
and U4041 (N_4041,N_1666,N_2472);
and U4042 (N_4042,N_2271,N_1037);
and U4043 (N_4043,N_539,N_1381);
nor U4044 (N_4044,N_1082,N_1144);
and U4045 (N_4045,N_1048,N_144);
nand U4046 (N_4046,N_1994,N_2263);
xor U4047 (N_4047,N_1759,N_547);
nand U4048 (N_4048,N_86,N_2379);
xnor U4049 (N_4049,N_2141,N_1293);
nor U4050 (N_4050,N_2139,N_2054);
nor U4051 (N_4051,N_592,N_1094);
xor U4052 (N_4052,N_2032,N_2455);
nor U4053 (N_4053,N_2498,N_153);
xor U4054 (N_4054,N_2184,N_1298);
or U4055 (N_4055,N_499,N_1401);
xor U4056 (N_4056,N_273,N_1113);
or U4057 (N_4057,N_957,N_339);
or U4058 (N_4058,N_1323,N_1803);
xor U4059 (N_4059,N_1378,N_95);
or U4060 (N_4060,N_455,N_1735);
nor U4061 (N_4061,N_892,N_1746);
nor U4062 (N_4062,N_1177,N_1554);
and U4063 (N_4063,N_1804,N_2001);
or U4064 (N_4064,N_2305,N_300);
nand U4065 (N_4065,N_1651,N_867);
and U4066 (N_4066,N_955,N_484);
nand U4067 (N_4067,N_2464,N_2113);
xor U4068 (N_4068,N_565,N_2206);
and U4069 (N_4069,N_461,N_17);
nor U4070 (N_4070,N_2161,N_2261);
nor U4071 (N_4071,N_723,N_1676);
nand U4072 (N_4072,N_1085,N_77);
or U4073 (N_4073,N_560,N_1908);
xor U4074 (N_4074,N_8,N_1863);
xor U4075 (N_4075,N_2312,N_372);
and U4076 (N_4076,N_29,N_1855);
nand U4077 (N_4077,N_2326,N_588);
and U4078 (N_4078,N_226,N_404);
xnor U4079 (N_4079,N_1932,N_16);
and U4080 (N_4080,N_2011,N_1557);
or U4081 (N_4081,N_2088,N_2236);
nor U4082 (N_4082,N_1779,N_581);
nand U4083 (N_4083,N_2023,N_1951);
and U4084 (N_4084,N_1177,N_2393);
nand U4085 (N_4085,N_948,N_1144);
or U4086 (N_4086,N_392,N_1746);
nand U4087 (N_4087,N_1512,N_1777);
nor U4088 (N_4088,N_2024,N_298);
nor U4089 (N_4089,N_2231,N_1984);
or U4090 (N_4090,N_872,N_1378);
and U4091 (N_4091,N_358,N_2224);
nand U4092 (N_4092,N_2440,N_2310);
and U4093 (N_4093,N_2316,N_1655);
xor U4094 (N_4094,N_1053,N_1837);
nor U4095 (N_4095,N_2215,N_2365);
and U4096 (N_4096,N_156,N_2013);
or U4097 (N_4097,N_1387,N_256);
nor U4098 (N_4098,N_2487,N_2060);
xnor U4099 (N_4099,N_2098,N_350);
and U4100 (N_4100,N_2220,N_659);
nor U4101 (N_4101,N_261,N_1007);
nor U4102 (N_4102,N_1477,N_1813);
and U4103 (N_4103,N_66,N_180);
xnor U4104 (N_4104,N_2141,N_754);
nand U4105 (N_4105,N_1750,N_55);
nor U4106 (N_4106,N_2092,N_371);
xnor U4107 (N_4107,N_1290,N_2302);
or U4108 (N_4108,N_1565,N_1025);
nand U4109 (N_4109,N_2490,N_1438);
nand U4110 (N_4110,N_1002,N_844);
or U4111 (N_4111,N_1500,N_32);
and U4112 (N_4112,N_1961,N_810);
and U4113 (N_4113,N_60,N_2063);
and U4114 (N_4114,N_1751,N_67);
or U4115 (N_4115,N_2046,N_220);
nand U4116 (N_4116,N_1493,N_1882);
or U4117 (N_4117,N_1755,N_1314);
and U4118 (N_4118,N_1225,N_1382);
and U4119 (N_4119,N_2023,N_2448);
and U4120 (N_4120,N_1158,N_298);
or U4121 (N_4121,N_1744,N_1838);
and U4122 (N_4122,N_2073,N_307);
and U4123 (N_4123,N_1627,N_488);
or U4124 (N_4124,N_2456,N_1825);
and U4125 (N_4125,N_2459,N_914);
nand U4126 (N_4126,N_2357,N_608);
and U4127 (N_4127,N_1139,N_71);
nor U4128 (N_4128,N_1843,N_2183);
nand U4129 (N_4129,N_2414,N_1330);
and U4130 (N_4130,N_1298,N_1068);
xor U4131 (N_4131,N_1171,N_608);
nand U4132 (N_4132,N_16,N_506);
nor U4133 (N_4133,N_1050,N_2438);
xor U4134 (N_4134,N_1847,N_1163);
or U4135 (N_4135,N_1084,N_1456);
or U4136 (N_4136,N_1254,N_1415);
nand U4137 (N_4137,N_818,N_1959);
nor U4138 (N_4138,N_2241,N_1546);
nor U4139 (N_4139,N_732,N_1382);
or U4140 (N_4140,N_1385,N_1902);
nor U4141 (N_4141,N_1465,N_360);
xor U4142 (N_4142,N_1109,N_1657);
or U4143 (N_4143,N_1924,N_1956);
nor U4144 (N_4144,N_1296,N_1289);
nor U4145 (N_4145,N_1794,N_1439);
or U4146 (N_4146,N_2325,N_147);
and U4147 (N_4147,N_405,N_2114);
nand U4148 (N_4148,N_834,N_912);
xor U4149 (N_4149,N_416,N_2461);
nand U4150 (N_4150,N_1253,N_1979);
nor U4151 (N_4151,N_1960,N_1578);
nand U4152 (N_4152,N_2418,N_1290);
xor U4153 (N_4153,N_1940,N_1753);
xnor U4154 (N_4154,N_1003,N_2467);
nor U4155 (N_4155,N_282,N_517);
xnor U4156 (N_4156,N_2211,N_370);
nor U4157 (N_4157,N_1271,N_702);
and U4158 (N_4158,N_1381,N_1222);
or U4159 (N_4159,N_2380,N_580);
nor U4160 (N_4160,N_428,N_307);
nor U4161 (N_4161,N_21,N_1082);
nand U4162 (N_4162,N_2276,N_451);
or U4163 (N_4163,N_2388,N_475);
xnor U4164 (N_4164,N_2009,N_845);
xnor U4165 (N_4165,N_1913,N_2057);
nand U4166 (N_4166,N_40,N_2188);
nand U4167 (N_4167,N_2416,N_1050);
nand U4168 (N_4168,N_1613,N_414);
nor U4169 (N_4169,N_2374,N_91);
and U4170 (N_4170,N_2363,N_378);
and U4171 (N_4171,N_2494,N_779);
nand U4172 (N_4172,N_1927,N_1124);
and U4173 (N_4173,N_801,N_38);
nand U4174 (N_4174,N_734,N_2309);
nor U4175 (N_4175,N_1731,N_1969);
and U4176 (N_4176,N_1931,N_61);
xnor U4177 (N_4177,N_423,N_2344);
and U4178 (N_4178,N_2370,N_1421);
and U4179 (N_4179,N_2148,N_1041);
nor U4180 (N_4180,N_1962,N_2039);
and U4181 (N_4181,N_2392,N_937);
nand U4182 (N_4182,N_906,N_181);
and U4183 (N_4183,N_611,N_2009);
nor U4184 (N_4184,N_1470,N_401);
nand U4185 (N_4185,N_1933,N_1045);
nand U4186 (N_4186,N_1985,N_71);
nand U4187 (N_4187,N_1174,N_1411);
and U4188 (N_4188,N_955,N_814);
and U4189 (N_4189,N_1527,N_953);
nand U4190 (N_4190,N_2379,N_2399);
and U4191 (N_4191,N_766,N_88);
or U4192 (N_4192,N_1776,N_585);
and U4193 (N_4193,N_1948,N_1453);
or U4194 (N_4194,N_430,N_1933);
and U4195 (N_4195,N_2228,N_1765);
nor U4196 (N_4196,N_1595,N_17);
or U4197 (N_4197,N_69,N_657);
nand U4198 (N_4198,N_307,N_2278);
nand U4199 (N_4199,N_183,N_2485);
and U4200 (N_4200,N_1967,N_1386);
nand U4201 (N_4201,N_2092,N_764);
nand U4202 (N_4202,N_284,N_2224);
nand U4203 (N_4203,N_66,N_1872);
or U4204 (N_4204,N_2320,N_2106);
and U4205 (N_4205,N_198,N_2059);
nor U4206 (N_4206,N_2063,N_1396);
xnor U4207 (N_4207,N_1243,N_2271);
and U4208 (N_4208,N_2125,N_995);
nor U4209 (N_4209,N_1733,N_2384);
nor U4210 (N_4210,N_905,N_370);
and U4211 (N_4211,N_25,N_674);
nand U4212 (N_4212,N_358,N_2407);
nor U4213 (N_4213,N_428,N_316);
nor U4214 (N_4214,N_1861,N_1909);
and U4215 (N_4215,N_2217,N_1684);
nand U4216 (N_4216,N_1093,N_1480);
nand U4217 (N_4217,N_1416,N_698);
and U4218 (N_4218,N_2217,N_1345);
or U4219 (N_4219,N_1938,N_1820);
xnor U4220 (N_4220,N_937,N_2175);
and U4221 (N_4221,N_2149,N_828);
nand U4222 (N_4222,N_2221,N_2459);
nand U4223 (N_4223,N_1716,N_718);
and U4224 (N_4224,N_1698,N_1925);
or U4225 (N_4225,N_533,N_2092);
xnor U4226 (N_4226,N_703,N_1914);
nor U4227 (N_4227,N_1292,N_958);
or U4228 (N_4228,N_2473,N_564);
nand U4229 (N_4229,N_1398,N_238);
and U4230 (N_4230,N_749,N_1593);
or U4231 (N_4231,N_1711,N_2423);
nor U4232 (N_4232,N_949,N_1990);
and U4233 (N_4233,N_1196,N_1298);
and U4234 (N_4234,N_2196,N_755);
nand U4235 (N_4235,N_1578,N_819);
xor U4236 (N_4236,N_827,N_1887);
or U4237 (N_4237,N_1874,N_1923);
xor U4238 (N_4238,N_2060,N_1989);
nor U4239 (N_4239,N_2227,N_1120);
and U4240 (N_4240,N_249,N_503);
xor U4241 (N_4241,N_1513,N_2012);
xor U4242 (N_4242,N_568,N_1817);
xor U4243 (N_4243,N_1545,N_2214);
or U4244 (N_4244,N_1774,N_1577);
nand U4245 (N_4245,N_1873,N_705);
xnor U4246 (N_4246,N_1611,N_2325);
nor U4247 (N_4247,N_843,N_1275);
or U4248 (N_4248,N_2111,N_1033);
nor U4249 (N_4249,N_790,N_2294);
xnor U4250 (N_4250,N_977,N_1909);
nor U4251 (N_4251,N_1183,N_739);
nand U4252 (N_4252,N_917,N_1049);
or U4253 (N_4253,N_2088,N_1418);
and U4254 (N_4254,N_1933,N_541);
or U4255 (N_4255,N_1390,N_1542);
nand U4256 (N_4256,N_1072,N_1879);
nor U4257 (N_4257,N_704,N_1107);
nand U4258 (N_4258,N_1499,N_2018);
and U4259 (N_4259,N_1398,N_2192);
xor U4260 (N_4260,N_488,N_1296);
and U4261 (N_4261,N_2251,N_2012);
and U4262 (N_4262,N_1377,N_325);
xor U4263 (N_4263,N_2055,N_1729);
nor U4264 (N_4264,N_1377,N_498);
xor U4265 (N_4265,N_1570,N_1531);
nand U4266 (N_4266,N_1426,N_49);
nand U4267 (N_4267,N_149,N_250);
xnor U4268 (N_4268,N_1483,N_149);
or U4269 (N_4269,N_628,N_197);
or U4270 (N_4270,N_641,N_2129);
or U4271 (N_4271,N_2102,N_1785);
nand U4272 (N_4272,N_1733,N_164);
nand U4273 (N_4273,N_1248,N_1643);
and U4274 (N_4274,N_221,N_2318);
and U4275 (N_4275,N_1963,N_78);
xor U4276 (N_4276,N_131,N_2469);
xnor U4277 (N_4277,N_1637,N_1833);
or U4278 (N_4278,N_1848,N_1526);
or U4279 (N_4279,N_609,N_1509);
nor U4280 (N_4280,N_1780,N_484);
and U4281 (N_4281,N_219,N_577);
xnor U4282 (N_4282,N_895,N_479);
or U4283 (N_4283,N_186,N_202);
nor U4284 (N_4284,N_1732,N_151);
nand U4285 (N_4285,N_1488,N_1145);
xor U4286 (N_4286,N_25,N_1313);
or U4287 (N_4287,N_115,N_1812);
or U4288 (N_4288,N_1556,N_1586);
and U4289 (N_4289,N_346,N_133);
and U4290 (N_4290,N_2163,N_1690);
and U4291 (N_4291,N_665,N_478);
nor U4292 (N_4292,N_775,N_750);
xor U4293 (N_4293,N_169,N_620);
and U4294 (N_4294,N_1409,N_1961);
and U4295 (N_4295,N_2138,N_386);
or U4296 (N_4296,N_2399,N_293);
or U4297 (N_4297,N_1388,N_1343);
nor U4298 (N_4298,N_1759,N_1122);
nor U4299 (N_4299,N_439,N_2406);
nand U4300 (N_4300,N_2440,N_881);
xnor U4301 (N_4301,N_1473,N_1879);
or U4302 (N_4302,N_625,N_281);
xor U4303 (N_4303,N_2340,N_2404);
nand U4304 (N_4304,N_2085,N_512);
xnor U4305 (N_4305,N_675,N_1176);
xnor U4306 (N_4306,N_1838,N_1646);
and U4307 (N_4307,N_551,N_395);
and U4308 (N_4308,N_1787,N_2261);
or U4309 (N_4309,N_122,N_1536);
nor U4310 (N_4310,N_2498,N_1296);
xor U4311 (N_4311,N_142,N_2310);
and U4312 (N_4312,N_673,N_1879);
xor U4313 (N_4313,N_365,N_1820);
nor U4314 (N_4314,N_851,N_1746);
nand U4315 (N_4315,N_874,N_205);
xnor U4316 (N_4316,N_1377,N_2015);
nand U4317 (N_4317,N_736,N_2485);
nor U4318 (N_4318,N_302,N_916);
and U4319 (N_4319,N_781,N_2164);
nor U4320 (N_4320,N_2020,N_216);
nor U4321 (N_4321,N_654,N_168);
and U4322 (N_4322,N_1449,N_2243);
nor U4323 (N_4323,N_1617,N_926);
nand U4324 (N_4324,N_1234,N_1726);
and U4325 (N_4325,N_109,N_1153);
nor U4326 (N_4326,N_348,N_2184);
nor U4327 (N_4327,N_1467,N_2384);
or U4328 (N_4328,N_1744,N_592);
nand U4329 (N_4329,N_2189,N_1478);
nor U4330 (N_4330,N_2053,N_2407);
and U4331 (N_4331,N_1915,N_313);
and U4332 (N_4332,N_757,N_2033);
nor U4333 (N_4333,N_1827,N_1502);
or U4334 (N_4334,N_150,N_90);
nand U4335 (N_4335,N_1267,N_312);
or U4336 (N_4336,N_2169,N_2232);
or U4337 (N_4337,N_1306,N_1900);
and U4338 (N_4338,N_384,N_2395);
or U4339 (N_4339,N_1214,N_1431);
or U4340 (N_4340,N_713,N_1383);
nor U4341 (N_4341,N_2489,N_26);
nor U4342 (N_4342,N_1978,N_877);
and U4343 (N_4343,N_503,N_2221);
nand U4344 (N_4344,N_1019,N_2102);
or U4345 (N_4345,N_894,N_1740);
nor U4346 (N_4346,N_499,N_1486);
nand U4347 (N_4347,N_973,N_887);
nand U4348 (N_4348,N_410,N_654);
and U4349 (N_4349,N_1322,N_64);
or U4350 (N_4350,N_2225,N_1902);
xor U4351 (N_4351,N_328,N_304);
xnor U4352 (N_4352,N_1399,N_491);
nor U4353 (N_4353,N_561,N_2206);
xnor U4354 (N_4354,N_2306,N_2299);
or U4355 (N_4355,N_1024,N_910);
or U4356 (N_4356,N_2144,N_1809);
or U4357 (N_4357,N_1385,N_887);
nor U4358 (N_4358,N_1543,N_1736);
nand U4359 (N_4359,N_1938,N_746);
xnor U4360 (N_4360,N_243,N_1478);
xor U4361 (N_4361,N_2062,N_24);
or U4362 (N_4362,N_647,N_2090);
xor U4363 (N_4363,N_606,N_242);
or U4364 (N_4364,N_2379,N_561);
nand U4365 (N_4365,N_270,N_1037);
xnor U4366 (N_4366,N_937,N_1133);
and U4367 (N_4367,N_980,N_2180);
xor U4368 (N_4368,N_475,N_1594);
or U4369 (N_4369,N_1352,N_749);
xor U4370 (N_4370,N_1514,N_723);
xnor U4371 (N_4371,N_198,N_649);
nor U4372 (N_4372,N_754,N_2379);
and U4373 (N_4373,N_2410,N_1962);
and U4374 (N_4374,N_2363,N_837);
or U4375 (N_4375,N_1243,N_621);
nand U4376 (N_4376,N_1789,N_871);
or U4377 (N_4377,N_181,N_1848);
xor U4378 (N_4378,N_1374,N_903);
nor U4379 (N_4379,N_871,N_410);
nor U4380 (N_4380,N_2168,N_1910);
nor U4381 (N_4381,N_1037,N_285);
nand U4382 (N_4382,N_705,N_1354);
or U4383 (N_4383,N_2187,N_1446);
xor U4384 (N_4384,N_905,N_1648);
and U4385 (N_4385,N_1278,N_1435);
or U4386 (N_4386,N_1137,N_613);
and U4387 (N_4387,N_288,N_609);
xnor U4388 (N_4388,N_947,N_1184);
and U4389 (N_4389,N_114,N_44);
xor U4390 (N_4390,N_476,N_63);
xor U4391 (N_4391,N_679,N_443);
nor U4392 (N_4392,N_1074,N_2321);
or U4393 (N_4393,N_2024,N_1330);
or U4394 (N_4394,N_948,N_2314);
or U4395 (N_4395,N_2131,N_1471);
nand U4396 (N_4396,N_371,N_2264);
or U4397 (N_4397,N_1070,N_108);
xor U4398 (N_4398,N_87,N_2155);
or U4399 (N_4399,N_349,N_1563);
nand U4400 (N_4400,N_599,N_2127);
nor U4401 (N_4401,N_2092,N_2185);
nor U4402 (N_4402,N_2317,N_1341);
or U4403 (N_4403,N_578,N_281);
nor U4404 (N_4404,N_482,N_980);
and U4405 (N_4405,N_345,N_654);
xnor U4406 (N_4406,N_411,N_1940);
nor U4407 (N_4407,N_576,N_1347);
nand U4408 (N_4408,N_893,N_913);
xor U4409 (N_4409,N_1438,N_1371);
or U4410 (N_4410,N_2276,N_1128);
nand U4411 (N_4411,N_2101,N_2144);
or U4412 (N_4412,N_2216,N_515);
or U4413 (N_4413,N_942,N_1873);
and U4414 (N_4414,N_2074,N_846);
or U4415 (N_4415,N_1405,N_553);
nand U4416 (N_4416,N_78,N_1138);
nand U4417 (N_4417,N_118,N_7);
xnor U4418 (N_4418,N_1364,N_1225);
nor U4419 (N_4419,N_783,N_776);
xor U4420 (N_4420,N_2421,N_2121);
nor U4421 (N_4421,N_2496,N_1932);
and U4422 (N_4422,N_1710,N_911);
xnor U4423 (N_4423,N_1373,N_1402);
nand U4424 (N_4424,N_1717,N_981);
nand U4425 (N_4425,N_257,N_1178);
and U4426 (N_4426,N_1596,N_2320);
nor U4427 (N_4427,N_2433,N_336);
nor U4428 (N_4428,N_1591,N_2090);
nand U4429 (N_4429,N_937,N_2135);
and U4430 (N_4430,N_1804,N_135);
nand U4431 (N_4431,N_642,N_435);
nor U4432 (N_4432,N_999,N_1041);
nor U4433 (N_4433,N_1896,N_1363);
xnor U4434 (N_4434,N_1014,N_2200);
nor U4435 (N_4435,N_2171,N_2057);
and U4436 (N_4436,N_202,N_950);
or U4437 (N_4437,N_1859,N_651);
or U4438 (N_4438,N_2493,N_1346);
nor U4439 (N_4439,N_2011,N_475);
and U4440 (N_4440,N_1524,N_614);
or U4441 (N_4441,N_1755,N_545);
xor U4442 (N_4442,N_1107,N_1276);
nor U4443 (N_4443,N_2275,N_794);
nand U4444 (N_4444,N_761,N_2030);
nand U4445 (N_4445,N_724,N_814);
or U4446 (N_4446,N_1315,N_356);
nand U4447 (N_4447,N_1118,N_1763);
nor U4448 (N_4448,N_596,N_556);
and U4449 (N_4449,N_2454,N_1330);
and U4450 (N_4450,N_358,N_2010);
xor U4451 (N_4451,N_10,N_930);
nand U4452 (N_4452,N_723,N_2078);
xnor U4453 (N_4453,N_462,N_2100);
xnor U4454 (N_4454,N_337,N_1035);
nand U4455 (N_4455,N_1746,N_1779);
and U4456 (N_4456,N_1243,N_2315);
and U4457 (N_4457,N_1780,N_1021);
nand U4458 (N_4458,N_2074,N_2171);
nor U4459 (N_4459,N_477,N_1692);
or U4460 (N_4460,N_313,N_1325);
or U4461 (N_4461,N_221,N_1772);
nor U4462 (N_4462,N_1285,N_848);
nor U4463 (N_4463,N_203,N_2261);
and U4464 (N_4464,N_914,N_1706);
and U4465 (N_4465,N_420,N_1744);
nor U4466 (N_4466,N_1783,N_444);
xnor U4467 (N_4467,N_804,N_314);
and U4468 (N_4468,N_1055,N_277);
nor U4469 (N_4469,N_780,N_1541);
nand U4470 (N_4470,N_2344,N_1387);
or U4471 (N_4471,N_1902,N_723);
xor U4472 (N_4472,N_297,N_1735);
or U4473 (N_4473,N_1375,N_285);
or U4474 (N_4474,N_1278,N_99);
xor U4475 (N_4475,N_2262,N_218);
xnor U4476 (N_4476,N_1507,N_1982);
xor U4477 (N_4477,N_1775,N_535);
nand U4478 (N_4478,N_392,N_719);
and U4479 (N_4479,N_1763,N_2389);
nor U4480 (N_4480,N_151,N_1141);
xnor U4481 (N_4481,N_1088,N_1471);
or U4482 (N_4482,N_803,N_1450);
nand U4483 (N_4483,N_1413,N_1034);
xnor U4484 (N_4484,N_450,N_512);
and U4485 (N_4485,N_1526,N_11);
and U4486 (N_4486,N_996,N_1562);
xnor U4487 (N_4487,N_45,N_1895);
and U4488 (N_4488,N_1221,N_1825);
or U4489 (N_4489,N_1904,N_565);
or U4490 (N_4490,N_394,N_1092);
and U4491 (N_4491,N_2160,N_91);
nor U4492 (N_4492,N_887,N_1818);
xnor U4493 (N_4493,N_1740,N_1471);
and U4494 (N_4494,N_690,N_1302);
or U4495 (N_4495,N_324,N_2432);
or U4496 (N_4496,N_677,N_375);
and U4497 (N_4497,N_98,N_1513);
xnor U4498 (N_4498,N_1936,N_344);
or U4499 (N_4499,N_1775,N_359);
nand U4500 (N_4500,N_1084,N_2252);
nor U4501 (N_4501,N_1202,N_1061);
xor U4502 (N_4502,N_1824,N_1630);
nor U4503 (N_4503,N_1617,N_1303);
or U4504 (N_4504,N_1057,N_984);
xnor U4505 (N_4505,N_63,N_2338);
nor U4506 (N_4506,N_878,N_460);
and U4507 (N_4507,N_485,N_342);
or U4508 (N_4508,N_73,N_91);
xnor U4509 (N_4509,N_1117,N_2164);
nand U4510 (N_4510,N_2329,N_1111);
xor U4511 (N_4511,N_608,N_1127);
nand U4512 (N_4512,N_1264,N_541);
or U4513 (N_4513,N_2399,N_1055);
or U4514 (N_4514,N_175,N_2051);
nand U4515 (N_4515,N_1061,N_2039);
or U4516 (N_4516,N_395,N_705);
nor U4517 (N_4517,N_2355,N_180);
xor U4518 (N_4518,N_817,N_2464);
nand U4519 (N_4519,N_1541,N_772);
or U4520 (N_4520,N_518,N_1774);
or U4521 (N_4521,N_2212,N_620);
nor U4522 (N_4522,N_1102,N_1043);
nor U4523 (N_4523,N_483,N_800);
nor U4524 (N_4524,N_1500,N_2274);
nand U4525 (N_4525,N_1195,N_673);
and U4526 (N_4526,N_948,N_386);
nor U4527 (N_4527,N_2043,N_1570);
and U4528 (N_4528,N_1927,N_2311);
nand U4529 (N_4529,N_815,N_1965);
or U4530 (N_4530,N_1829,N_1051);
and U4531 (N_4531,N_2195,N_667);
nand U4532 (N_4532,N_2378,N_1720);
nand U4533 (N_4533,N_1084,N_643);
nor U4534 (N_4534,N_1400,N_1777);
xor U4535 (N_4535,N_319,N_200);
nand U4536 (N_4536,N_528,N_1142);
or U4537 (N_4537,N_2198,N_1713);
nor U4538 (N_4538,N_2312,N_1939);
or U4539 (N_4539,N_1899,N_1266);
or U4540 (N_4540,N_2119,N_2493);
xnor U4541 (N_4541,N_232,N_982);
or U4542 (N_4542,N_2281,N_1483);
xnor U4543 (N_4543,N_1899,N_2196);
nor U4544 (N_4544,N_1175,N_1902);
xor U4545 (N_4545,N_1351,N_417);
or U4546 (N_4546,N_310,N_1831);
nor U4547 (N_4547,N_250,N_1202);
nor U4548 (N_4548,N_1412,N_1190);
nor U4549 (N_4549,N_308,N_1919);
nand U4550 (N_4550,N_1896,N_49);
or U4551 (N_4551,N_1209,N_952);
nor U4552 (N_4552,N_1648,N_1973);
and U4553 (N_4553,N_2215,N_753);
nor U4554 (N_4554,N_2364,N_1973);
nand U4555 (N_4555,N_500,N_2295);
nor U4556 (N_4556,N_928,N_1771);
or U4557 (N_4557,N_317,N_694);
nor U4558 (N_4558,N_1382,N_5);
xor U4559 (N_4559,N_1201,N_59);
nand U4560 (N_4560,N_2287,N_1432);
and U4561 (N_4561,N_934,N_1790);
or U4562 (N_4562,N_760,N_1802);
xnor U4563 (N_4563,N_2298,N_2000);
or U4564 (N_4564,N_2167,N_981);
xor U4565 (N_4565,N_1474,N_831);
nor U4566 (N_4566,N_2080,N_740);
nor U4567 (N_4567,N_2238,N_1424);
and U4568 (N_4568,N_90,N_2338);
or U4569 (N_4569,N_294,N_92);
nor U4570 (N_4570,N_1775,N_2253);
and U4571 (N_4571,N_551,N_2035);
or U4572 (N_4572,N_2149,N_111);
nand U4573 (N_4573,N_1067,N_379);
or U4574 (N_4574,N_2294,N_706);
nand U4575 (N_4575,N_1758,N_223);
and U4576 (N_4576,N_534,N_2275);
or U4577 (N_4577,N_2256,N_2081);
and U4578 (N_4578,N_712,N_379);
nand U4579 (N_4579,N_605,N_1357);
or U4580 (N_4580,N_1773,N_1689);
or U4581 (N_4581,N_681,N_132);
or U4582 (N_4582,N_2196,N_2172);
nor U4583 (N_4583,N_1893,N_1055);
nand U4584 (N_4584,N_1062,N_1993);
xnor U4585 (N_4585,N_369,N_1624);
xor U4586 (N_4586,N_150,N_1870);
nor U4587 (N_4587,N_711,N_1051);
nand U4588 (N_4588,N_1605,N_1399);
nor U4589 (N_4589,N_1112,N_2156);
or U4590 (N_4590,N_1264,N_912);
and U4591 (N_4591,N_2471,N_25);
nor U4592 (N_4592,N_1552,N_163);
and U4593 (N_4593,N_944,N_1501);
xor U4594 (N_4594,N_2231,N_2047);
or U4595 (N_4595,N_587,N_450);
and U4596 (N_4596,N_1751,N_33);
nor U4597 (N_4597,N_1603,N_1403);
or U4598 (N_4598,N_1318,N_1827);
xnor U4599 (N_4599,N_2283,N_1615);
and U4600 (N_4600,N_1271,N_1876);
xor U4601 (N_4601,N_2170,N_1903);
nand U4602 (N_4602,N_1912,N_670);
and U4603 (N_4603,N_2319,N_2341);
and U4604 (N_4604,N_2395,N_1689);
nor U4605 (N_4605,N_2029,N_1452);
nor U4606 (N_4606,N_210,N_907);
or U4607 (N_4607,N_688,N_2458);
or U4608 (N_4608,N_1612,N_232);
xor U4609 (N_4609,N_731,N_1808);
nor U4610 (N_4610,N_495,N_1887);
nor U4611 (N_4611,N_1197,N_833);
or U4612 (N_4612,N_643,N_2292);
or U4613 (N_4613,N_2031,N_1222);
and U4614 (N_4614,N_1709,N_1022);
xor U4615 (N_4615,N_689,N_1057);
or U4616 (N_4616,N_1855,N_449);
nor U4617 (N_4617,N_2118,N_1414);
nand U4618 (N_4618,N_938,N_1072);
nor U4619 (N_4619,N_1714,N_2155);
nor U4620 (N_4620,N_2119,N_68);
nor U4621 (N_4621,N_314,N_1165);
nor U4622 (N_4622,N_1930,N_1115);
nand U4623 (N_4623,N_995,N_1996);
and U4624 (N_4624,N_443,N_1544);
nor U4625 (N_4625,N_89,N_1380);
nor U4626 (N_4626,N_208,N_1872);
nand U4627 (N_4627,N_2315,N_2074);
or U4628 (N_4628,N_354,N_743);
and U4629 (N_4629,N_1588,N_1971);
and U4630 (N_4630,N_1195,N_1645);
and U4631 (N_4631,N_1318,N_2329);
nand U4632 (N_4632,N_2478,N_22);
xor U4633 (N_4633,N_384,N_1135);
and U4634 (N_4634,N_2121,N_2159);
and U4635 (N_4635,N_1165,N_1036);
or U4636 (N_4636,N_1057,N_895);
and U4637 (N_4637,N_2312,N_2157);
nand U4638 (N_4638,N_997,N_1161);
or U4639 (N_4639,N_507,N_1850);
nand U4640 (N_4640,N_2166,N_459);
nor U4641 (N_4641,N_827,N_443);
nand U4642 (N_4642,N_1578,N_850);
or U4643 (N_4643,N_585,N_628);
xnor U4644 (N_4644,N_2436,N_1250);
xor U4645 (N_4645,N_1286,N_2354);
nor U4646 (N_4646,N_1201,N_892);
xnor U4647 (N_4647,N_806,N_981);
or U4648 (N_4648,N_1804,N_880);
and U4649 (N_4649,N_1259,N_1629);
nor U4650 (N_4650,N_1125,N_1940);
xnor U4651 (N_4651,N_1908,N_2278);
xor U4652 (N_4652,N_1479,N_2327);
or U4653 (N_4653,N_195,N_2290);
or U4654 (N_4654,N_1175,N_187);
and U4655 (N_4655,N_1243,N_698);
xor U4656 (N_4656,N_254,N_465);
xor U4657 (N_4657,N_784,N_1912);
and U4658 (N_4658,N_1920,N_718);
or U4659 (N_4659,N_1892,N_383);
or U4660 (N_4660,N_2252,N_2063);
nand U4661 (N_4661,N_1095,N_1622);
xnor U4662 (N_4662,N_262,N_2187);
nor U4663 (N_4663,N_680,N_385);
nor U4664 (N_4664,N_713,N_821);
nand U4665 (N_4665,N_170,N_691);
or U4666 (N_4666,N_1673,N_594);
or U4667 (N_4667,N_748,N_2390);
nor U4668 (N_4668,N_903,N_2197);
nand U4669 (N_4669,N_701,N_1259);
or U4670 (N_4670,N_705,N_1899);
and U4671 (N_4671,N_1742,N_923);
or U4672 (N_4672,N_1125,N_958);
xor U4673 (N_4673,N_858,N_1698);
nand U4674 (N_4674,N_371,N_2323);
xor U4675 (N_4675,N_389,N_894);
nor U4676 (N_4676,N_422,N_2434);
nor U4677 (N_4677,N_1711,N_1297);
nand U4678 (N_4678,N_183,N_2266);
and U4679 (N_4679,N_485,N_1804);
or U4680 (N_4680,N_450,N_1209);
xnor U4681 (N_4681,N_701,N_57);
xor U4682 (N_4682,N_1940,N_668);
nor U4683 (N_4683,N_426,N_2279);
or U4684 (N_4684,N_1637,N_2414);
xnor U4685 (N_4685,N_1368,N_2109);
nand U4686 (N_4686,N_62,N_1729);
and U4687 (N_4687,N_2261,N_990);
nand U4688 (N_4688,N_1957,N_877);
nor U4689 (N_4689,N_1222,N_383);
or U4690 (N_4690,N_861,N_1823);
and U4691 (N_4691,N_1114,N_1792);
and U4692 (N_4692,N_866,N_908);
nand U4693 (N_4693,N_835,N_1785);
or U4694 (N_4694,N_444,N_741);
nor U4695 (N_4695,N_1280,N_800);
nand U4696 (N_4696,N_902,N_656);
or U4697 (N_4697,N_1207,N_422);
nor U4698 (N_4698,N_1261,N_1017);
or U4699 (N_4699,N_1100,N_939);
and U4700 (N_4700,N_1796,N_1747);
nand U4701 (N_4701,N_1491,N_705);
and U4702 (N_4702,N_2055,N_2362);
or U4703 (N_4703,N_2461,N_2229);
xnor U4704 (N_4704,N_1675,N_2348);
nand U4705 (N_4705,N_1623,N_895);
nand U4706 (N_4706,N_1451,N_441);
xnor U4707 (N_4707,N_2373,N_1921);
or U4708 (N_4708,N_1290,N_1854);
nand U4709 (N_4709,N_1340,N_1411);
and U4710 (N_4710,N_1379,N_17);
nand U4711 (N_4711,N_1556,N_1091);
xor U4712 (N_4712,N_719,N_718);
nand U4713 (N_4713,N_777,N_1601);
and U4714 (N_4714,N_601,N_830);
nor U4715 (N_4715,N_1404,N_2160);
nor U4716 (N_4716,N_149,N_1374);
nor U4717 (N_4717,N_539,N_2348);
and U4718 (N_4718,N_1052,N_807);
and U4719 (N_4719,N_2302,N_2275);
nor U4720 (N_4720,N_2368,N_95);
xor U4721 (N_4721,N_2329,N_522);
and U4722 (N_4722,N_1160,N_1086);
nand U4723 (N_4723,N_2318,N_1871);
nor U4724 (N_4724,N_420,N_944);
nand U4725 (N_4725,N_1223,N_796);
nand U4726 (N_4726,N_248,N_1477);
or U4727 (N_4727,N_612,N_1554);
nand U4728 (N_4728,N_1543,N_1010);
or U4729 (N_4729,N_2011,N_2003);
nand U4730 (N_4730,N_1341,N_536);
nor U4731 (N_4731,N_1243,N_532);
xor U4732 (N_4732,N_221,N_1985);
and U4733 (N_4733,N_16,N_928);
nor U4734 (N_4734,N_900,N_2199);
or U4735 (N_4735,N_505,N_1856);
nor U4736 (N_4736,N_1493,N_2335);
nor U4737 (N_4737,N_2184,N_1859);
nand U4738 (N_4738,N_1248,N_1727);
nand U4739 (N_4739,N_1407,N_44);
and U4740 (N_4740,N_18,N_890);
nand U4741 (N_4741,N_635,N_1498);
and U4742 (N_4742,N_1212,N_2048);
or U4743 (N_4743,N_1497,N_1522);
and U4744 (N_4744,N_87,N_884);
nand U4745 (N_4745,N_278,N_1998);
nand U4746 (N_4746,N_1067,N_1793);
xor U4747 (N_4747,N_1579,N_1140);
nor U4748 (N_4748,N_1888,N_172);
nand U4749 (N_4749,N_2274,N_1697);
xor U4750 (N_4750,N_270,N_62);
nand U4751 (N_4751,N_1459,N_1290);
xor U4752 (N_4752,N_1483,N_2469);
and U4753 (N_4753,N_411,N_494);
or U4754 (N_4754,N_2043,N_49);
and U4755 (N_4755,N_1197,N_1814);
or U4756 (N_4756,N_1422,N_935);
xnor U4757 (N_4757,N_821,N_879);
nand U4758 (N_4758,N_1381,N_1112);
nand U4759 (N_4759,N_1997,N_1757);
or U4760 (N_4760,N_231,N_2063);
nor U4761 (N_4761,N_2449,N_1655);
and U4762 (N_4762,N_1916,N_1119);
or U4763 (N_4763,N_2447,N_2140);
and U4764 (N_4764,N_485,N_704);
nand U4765 (N_4765,N_425,N_2164);
xnor U4766 (N_4766,N_674,N_2428);
xor U4767 (N_4767,N_797,N_369);
nor U4768 (N_4768,N_131,N_108);
xor U4769 (N_4769,N_81,N_843);
and U4770 (N_4770,N_2262,N_1687);
nand U4771 (N_4771,N_2198,N_1614);
or U4772 (N_4772,N_2255,N_504);
or U4773 (N_4773,N_629,N_1685);
nand U4774 (N_4774,N_2423,N_611);
nor U4775 (N_4775,N_579,N_1414);
xor U4776 (N_4776,N_1069,N_2429);
or U4777 (N_4777,N_1076,N_1200);
and U4778 (N_4778,N_2422,N_10);
xnor U4779 (N_4779,N_711,N_1181);
nand U4780 (N_4780,N_1985,N_1627);
and U4781 (N_4781,N_2120,N_1654);
or U4782 (N_4782,N_429,N_1478);
nand U4783 (N_4783,N_932,N_1097);
or U4784 (N_4784,N_2121,N_141);
or U4785 (N_4785,N_1672,N_1115);
xnor U4786 (N_4786,N_2493,N_375);
or U4787 (N_4787,N_1040,N_904);
and U4788 (N_4788,N_1598,N_989);
or U4789 (N_4789,N_331,N_362);
and U4790 (N_4790,N_2355,N_2352);
nor U4791 (N_4791,N_460,N_725);
nand U4792 (N_4792,N_186,N_365);
or U4793 (N_4793,N_2497,N_1579);
and U4794 (N_4794,N_1580,N_1621);
xnor U4795 (N_4795,N_320,N_1576);
nor U4796 (N_4796,N_993,N_1045);
or U4797 (N_4797,N_2044,N_1426);
xor U4798 (N_4798,N_2459,N_143);
xnor U4799 (N_4799,N_1326,N_643);
or U4800 (N_4800,N_381,N_1794);
xnor U4801 (N_4801,N_2285,N_2324);
or U4802 (N_4802,N_1319,N_2133);
or U4803 (N_4803,N_476,N_1238);
xor U4804 (N_4804,N_2263,N_1649);
nand U4805 (N_4805,N_2045,N_2285);
nand U4806 (N_4806,N_2488,N_1049);
nand U4807 (N_4807,N_1121,N_786);
nand U4808 (N_4808,N_1893,N_127);
or U4809 (N_4809,N_1936,N_2223);
or U4810 (N_4810,N_250,N_544);
or U4811 (N_4811,N_258,N_1789);
or U4812 (N_4812,N_1491,N_462);
nor U4813 (N_4813,N_1176,N_563);
and U4814 (N_4814,N_1092,N_1785);
nand U4815 (N_4815,N_2115,N_2315);
nor U4816 (N_4816,N_2057,N_2010);
and U4817 (N_4817,N_2232,N_1917);
xor U4818 (N_4818,N_1109,N_1670);
xor U4819 (N_4819,N_175,N_1470);
or U4820 (N_4820,N_1295,N_1126);
nand U4821 (N_4821,N_925,N_1638);
nand U4822 (N_4822,N_989,N_1819);
and U4823 (N_4823,N_15,N_256);
nor U4824 (N_4824,N_2141,N_1522);
nor U4825 (N_4825,N_1530,N_2260);
and U4826 (N_4826,N_1771,N_2090);
xor U4827 (N_4827,N_2132,N_1915);
and U4828 (N_4828,N_1198,N_2192);
nor U4829 (N_4829,N_129,N_1777);
nor U4830 (N_4830,N_774,N_429);
and U4831 (N_4831,N_1276,N_612);
nor U4832 (N_4832,N_2405,N_846);
or U4833 (N_4833,N_1200,N_901);
or U4834 (N_4834,N_1045,N_300);
nand U4835 (N_4835,N_948,N_2486);
nor U4836 (N_4836,N_603,N_1196);
and U4837 (N_4837,N_1319,N_2482);
or U4838 (N_4838,N_2326,N_1677);
nand U4839 (N_4839,N_47,N_847);
xnor U4840 (N_4840,N_584,N_2086);
nand U4841 (N_4841,N_1930,N_1233);
nor U4842 (N_4842,N_97,N_435);
and U4843 (N_4843,N_1954,N_168);
and U4844 (N_4844,N_1370,N_307);
and U4845 (N_4845,N_1211,N_1170);
xor U4846 (N_4846,N_2383,N_1624);
nand U4847 (N_4847,N_1480,N_2276);
and U4848 (N_4848,N_1541,N_56);
nor U4849 (N_4849,N_2192,N_1353);
and U4850 (N_4850,N_539,N_46);
or U4851 (N_4851,N_1067,N_475);
nand U4852 (N_4852,N_2434,N_691);
and U4853 (N_4853,N_2079,N_1018);
nor U4854 (N_4854,N_1921,N_675);
nor U4855 (N_4855,N_1138,N_224);
xnor U4856 (N_4856,N_219,N_2077);
or U4857 (N_4857,N_102,N_832);
and U4858 (N_4858,N_1926,N_164);
nor U4859 (N_4859,N_1304,N_1435);
nand U4860 (N_4860,N_1297,N_1903);
and U4861 (N_4861,N_1817,N_1991);
or U4862 (N_4862,N_510,N_1843);
xnor U4863 (N_4863,N_1202,N_2317);
xor U4864 (N_4864,N_1694,N_83);
and U4865 (N_4865,N_1612,N_1279);
xnor U4866 (N_4866,N_1369,N_607);
or U4867 (N_4867,N_347,N_1354);
and U4868 (N_4868,N_65,N_307);
and U4869 (N_4869,N_1805,N_268);
xnor U4870 (N_4870,N_1389,N_1221);
xor U4871 (N_4871,N_2403,N_895);
xor U4872 (N_4872,N_679,N_1780);
nor U4873 (N_4873,N_1310,N_115);
xnor U4874 (N_4874,N_306,N_870);
and U4875 (N_4875,N_2269,N_1706);
xor U4876 (N_4876,N_1127,N_2299);
and U4877 (N_4877,N_584,N_1977);
nand U4878 (N_4878,N_418,N_1202);
xnor U4879 (N_4879,N_1384,N_791);
xnor U4880 (N_4880,N_80,N_2227);
xor U4881 (N_4881,N_817,N_1620);
nand U4882 (N_4882,N_2222,N_1726);
nor U4883 (N_4883,N_1787,N_1634);
xnor U4884 (N_4884,N_1351,N_2260);
and U4885 (N_4885,N_1521,N_1434);
xor U4886 (N_4886,N_1277,N_70);
nor U4887 (N_4887,N_1427,N_1471);
or U4888 (N_4888,N_1527,N_1457);
xnor U4889 (N_4889,N_63,N_591);
nor U4890 (N_4890,N_469,N_2417);
nand U4891 (N_4891,N_1882,N_401);
and U4892 (N_4892,N_466,N_593);
or U4893 (N_4893,N_2389,N_986);
or U4894 (N_4894,N_55,N_746);
xnor U4895 (N_4895,N_1287,N_1841);
and U4896 (N_4896,N_2263,N_1519);
or U4897 (N_4897,N_242,N_2486);
nand U4898 (N_4898,N_142,N_331);
or U4899 (N_4899,N_370,N_2241);
xor U4900 (N_4900,N_867,N_2095);
or U4901 (N_4901,N_1701,N_1569);
xnor U4902 (N_4902,N_2056,N_1094);
nor U4903 (N_4903,N_2203,N_1683);
and U4904 (N_4904,N_972,N_11);
nand U4905 (N_4905,N_2365,N_36);
and U4906 (N_4906,N_559,N_258);
or U4907 (N_4907,N_2053,N_2149);
xnor U4908 (N_4908,N_1924,N_1794);
xnor U4909 (N_4909,N_154,N_839);
and U4910 (N_4910,N_331,N_45);
or U4911 (N_4911,N_520,N_2365);
xor U4912 (N_4912,N_2344,N_1463);
and U4913 (N_4913,N_1877,N_1611);
or U4914 (N_4914,N_1028,N_2321);
nand U4915 (N_4915,N_968,N_864);
xor U4916 (N_4916,N_138,N_1191);
and U4917 (N_4917,N_2222,N_2290);
nor U4918 (N_4918,N_1454,N_2396);
nor U4919 (N_4919,N_637,N_1920);
xnor U4920 (N_4920,N_1854,N_142);
nand U4921 (N_4921,N_1694,N_2249);
or U4922 (N_4922,N_1404,N_1141);
and U4923 (N_4923,N_1229,N_600);
nand U4924 (N_4924,N_1879,N_964);
nor U4925 (N_4925,N_2424,N_957);
xnor U4926 (N_4926,N_2057,N_965);
and U4927 (N_4927,N_1965,N_1454);
nand U4928 (N_4928,N_2079,N_444);
nor U4929 (N_4929,N_1820,N_1044);
xnor U4930 (N_4930,N_2270,N_1976);
nand U4931 (N_4931,N_1379,N_1481);
xnor U4932 (N_4932,N_2429,N_828);
nor U4933 (N_4933,N_65,N_1949);
xnor U4934 (N_4934,N_1539,N_2184);
and U4935 (N_4935,N_1788,N_1672);
xor U4936 (N_4936,N_1538,N_400);
nand U4937 (N_4937,N_1056,N_2441);
nor U4938 (N_4938,N_1985,N_1133);
and U4939 (N_4939,N_163,N_1902);
xor U4940 (N_4940,N_2392,N_2292);
nor U4941 (N_4941,N_865,N_1275);
or U4942 (N_4942,N_1522,N_1001);
or U4943 (N_4943,N_1472,N_967);
and U4944 (N_4944,N_587,N_1123);
or U4945 (N_4945,N_2111,N_324);
nand U4946 (N_4946,N_147,N_162);
nand U4947 (N_4947,N_2332,N_2263);
and U4948 (N_4948,N_1742,N_853);
and U4949 (N_4949,N_1783,N_838);
or U4950 (N_4950,N_745,N_421);
and U4951 (N_4951,N_731,N_2067);
and U4952 (N_4952,N_463,N_732);
nand U4953 (N_4953,N_1542,N_1889);
nand U4954 (N_4954,N_1479,N_635);
nor U4955 (N_4955,N_1281,N_1994);
and U4956 (N_4956,N_260,N_1424);
xnor U4957 (N_4957,N_277,N_1439);
or U4958 (N_4958,N_1242,N_1652);
nor U4959 (N_4959,N_284,N_1391);
or U4960 (N_4960,N_445,N_1026);
xnor U4961 (N_4961,N_1538,N_2406);
nand U4962 (N_4962,N_1671,N_880);
xnor U4963 (N_4963,N_978,N_1983);
nor U4964 (N_4964,N_2498,N_1598);
nor U4965 (N_4965,N_1744,N_1776);
and U4966 (N_4966,N_356,N_2042);
nand U4967 (N_4967,N_749,N_267);
nor U4968 (N_4968,N_160,N_1707);
or U4969 (N_4969,N_579,N_2264);
nand U4970 (N_4970,N_1915,N_1509);
xnor U4971 (N_4971,N_832,N_2147);
and U4972 (N_4972,N_2059,N_253);
nand U4973 (N_4973,N_186,N_747);
xnor U4974 (N_4974,N_273,N_1785);
and U4975 (N_4975,N_1720,N_603);
nand U4976 (N_4976,N_217,N_119);
xnor U4977 (N_4977,N_645,N_2480);
xor U4978 (N_4978,N_298,N_371);
or U4979 (N_4979,N_2223,N_1051);
nand U4980 (N_4980,N_2220,N_740);
and U4981 (N_4981,N_937,N_374);
and U4982 (N_4982,N_1179,N_1816);
or U4983 (N_4983,N_396,N_2429);
xor U4984 (N_4984,N_598,N_36);
or U4985 (N_4985,N_124,N_1276);
or U4986 (N_4986,N_2246,N_358);
xnor U4987 (N_4987,N_34,N_77);
nor U4988 (N_4988,N_657,N_71);
and U4989 (N_4989,N_1864,N_1961);
xnor U4990 (N_4990,N_971,N_1355);
xor U4991 (N_4991,N_961,N_440);
xor U4992 (N_4992,N_2261,N_1118);
nand U4993 (N_4993,N_1346,N_323);
nand U4994 (N_4994,N_813,N_2387);
nor U4995 (N_4995,N_368,N_1781);
or U4996 (N_4996,N_2210,N_1245);
nor U4997 (N_4997,N_1412,N_1789);
nor U4998 (N_4998,N_95,N_1922);
and U4999 (N_4999,N_2466,N_820);
nand U5000 (N_5000,N_4141,N_2849);
or U5001 (N_5001,N_4598,N_4686);
or U5002 (N_5002,N_4450,N_4860);
xnor U5003 (N_5003,N_2877,N_4461);
and U5004 (N_5004,N_2547,N_3707);
or U5005 (N_5005,N_3458,N_4837);
nor U5006 (N_5006,N_4884,N_4424);
and U5007 (N_5007,N_4490,N_4983);
nor U5008 (N_5008,N_4687,N_3105);
nor U5009 (N_5009,N_4236,N_2764);
nor U5010 (N_5010,N_2776,N_3510);
and U5011 (N_5011,N_3949,N_4906);
and U5012 (N_5012,N_4868,N_2845);
nand U5013 (N_5013,N_4846,N_4858);
nand U5014 (N_5014,N_2783,N_2625);
or U5015 (N_5015,N_4955,N_3104);
nor U5016 (N_5016,N_2627,N_3820);
and U5017 (N_5017,N_3073,N_4965);
xor U5018 (N_5018,N_4932,N_3403);
nand U5019 (N_5019,N_2553,N_3290);
or U5020 (N_5020,N_3401,N_4668);
and U5021 (N_5021,N_3211,N_4621);
xnor U5022 (N_5022,N_3460,N_4558);
or U5023 (N_5023,N_4250,N_3503);
or U5024 (N_5024,N_4924,N_4227);
nor U5025 (N_5025,N_2773,N_3415);
xor U5026 (N_5026,N_2980,N_3123);
nor U5027 (N_5027,N_2653,N_3421);
and U5028 (N_5028,N_3232,N_4468);
nor U5029 (N_5029,N_3739,N_3579);
and U5030 (N_5030,N_4184,N_4277);
nor U5031 (N_5031,N_3940,N_4781);
nand U5032 (N_5032,N_3295,N_3916);
nand U5033 (N_5033,N_4644,N_4909);
and U5034 (N_5034,N_4084,N_4625);
or U5035 (N_5035,N_4859,N_3167);
nand U5036 (N_5036,N_3067,N_2780);
nor U5037 (N_5037,N_4109,N_2957);
nand U5038 (N_5038,N_3423,N_3692);
nand U5039 (N_5039,N_3191,N_3530);
xor U5040 (N_5040,N_3077,N_3994);
nand U5041 (N_5041,N_3584,N_4241);
nor U5042 (N_5042,N_2556,N_3734);
nor U5043 (N_5043,N_4413,N_3651);
and U5044 (N_5044,N_4376,N_3800);
or U5045 (N_5045,N_2614,N_3494);
nand U5046 (N_5046,N_2648,N_3576);
and U5047 (N_5047,N_3449,N_3010);
xnor U5048 (N_5048,N_4820,N_4667);
nor U5049 (N_5049,N_3022,N_2623);
and U5050 (N_5050,N_3902,N_4824);
nor U5051 (N_5051,N_3234,N_2812);
or U5052 (N_5052,N_3374,N_4723);
xnor U5053 (N_5053,N_4029,N_2528);
xor U5054 (N_5054,N_3122,N_4460);
and U5055 (N_5055,N_2684,N_4519);
and U5056 (N_5056,N_4513,N_4321);
nand U5057 (N_5057,N_4193,N_3453);
nand U5058 (N_5058,N_3454,N_4721);
or U5059 (N_5059,N_3544,N_2637);
nand U5060 (N_5060,N_4582,N_3223);
nand U5061 (N_5061,N_4606,N_4019);
nor U5062 (N_5062,N_2620,N_2523);
nand U5063 (N_5063,N_2792,N_3407);
nand U5064 (N_5064,N_2633,N_3144);
xor U5065 (N_5065,N_4384,N_3642);
or U5066 (N_5066,N_3773,N_3682);
and U5067 (N_5067,N_4192,N_3942);
xnor U5068 (N_5068,N_4295,N_3496);
and U5069 (N_5069,N_4744,N_4794);
or U5070 (N_5070,N_3293,N_2664);
and U5071 (N_5071,N_4374,N_4529);
xor U5072 (N_5072,N_2722,N_3023);
xnor U5073 (N_5073,N_2994,N_3359);
nand U5074 (N_5074,N_4684,N_4467);
xor U5075 (N_5075,N_4394,N_2679);
and U5076 (N_5076,N_3491,N_2751);
xor U5077 (N_5077,N_3370,N_4850);
nor U5078 (N_5078,N_3649,N_3975);
xor U5079 (N_5079,N_4616,N_3622);
nor U5080 (N_5080,N_4849,N_3200);
or U5081 (N_5081,N_4525,N_2631);
xor U5082 (N_5082,N_3516,N_4627);
or U5083 (N_5083,N_3482,N_3178);
and U5084 (N_5084,N_3981,N_2605);
nor U5085 (N_5085,N_3891,N_3957);
nor U5086 (N_5086,N_3656,N_3101);
nor U5087 (N_5087,N_4808,N_3390);
xnor U5088 (N_5088,N_4202,N_3065);
and U5089 (N_5089,N_4501,N_4695);
xnor U5090 (N_5090,N_3896,N_3645);
nor U5091 (N_5091,N_3470,N_3464);
nor U5092 (N_5092,N_4987,N_2928);
xnor U5093 (N_5093,N_4007,N_2870);
or U5094 (N_5094,N_4156,N_3671);
or U5095 (N_5095,N_3059,N_2744);
xor U5096 (N_5096,N_3786,N_3261);
nand U5097 (N_5097,N_2883,N_4379);
nand U5098 (N_5098,N_4206,N_3974);
nand U5099 (N_5099,N_3589,N_4425);
nor U5100 (N_5100,N_3680,N_4713);
or U5101 (N_5101,N_3898,N_3970);
or U5102 (N_5102,N_4654,N_3157);
and U5103 (N_5103,N_3054,N_3485);
nand U5104 (N_5104,N_3131,N_3623);
and U5105 (N_5105,N_3695,N_4431);
nand U5106 (N_5106,N_4343,N_3979);
or U5107 (N_5107,N_3219,N_4632);
and U5108 (N_5108,N_4171,N_4998);
or U5109 (N_5109,N_4039,N_3409);
nor U5110 (N_5110,N_4051,N_3932);
or U5111 (N_5111,N_3360,N_4871);
xor U5112 (N_5112,N_3352,N_2854);
nor U5113 (N_5113,N_4328,N_4053);
nand U5114 (N_5114,N_4506,N_2887);
nor U5115 (N_5115,N_3260,N_4068);
nand U5116 (N_5116,N_2896,N_4726);
nor U5117 (N_5117,N_4026,N_2910);
or U5118 (N_5118,N_4257,N_4892);
nand U5119 (N_5119,N_4040,N_4307);
and U5120 (N_5120,N_4327,N_4420);
xor U5121 (N_5121,N_3930,N_3712);
nand U5122 (N_5122,N_3484,N_3110);
nand U5123 (N_5123,N_4989,N_3309);
nand U5124 (N_5124,N_3967,N_3334);
nor U5125 (N_5125,N_2800,N_3526);
nor U5126 (N_5126,N_4309,N_4521);
xor U5127 (N_5127,N_3426,N_3667);
nand U5128 (N_5128,N_4159,N_3330);
and U5129 (N_5129,N_2732,N_3286);
nor U5130 (N_5130,N_3189,N_3431);
nor U5131 (N_5131,N_3722,N_2789);
nor U5132 (N_5132,N_3808,N_3356);
nand U5133 (N_5133,N_3850,N_3049);
or U5134 (N_5134,N_4674,N_3305);
nand U5135 (N_5135,N_3117,N_2612);
xnor U5136 (N_5136,N_2685,N_3111);
nand U5137 (N_5137,N_3673,N_3338);
nor U5138 (N_5138,N_4825,N_3171);
xnor U5139 (N_5139,N_3648,N_3794);
xor U5140 (N_5140,N_4483,N_2639);
nor U5141 (N_5141,N_3302,N_4653);
and U5142 (N_5142,N_3128,N_4323);
and U5143 (N_5143,N_4404,N_4391);
nor U5144 (N_5144,N_3999,N_4382);
xnor U5145 (N_5145,N_4365,N_3976);
and U5146 (N_5146,N_4008,N_3133);
nor U5147 (N_5147,N_4408,N_2798);
xnor U5148 (N_5148,N_3728,N_2716);
nand U5149 (N_5149,N_2651,N_3418);
nand U5150 (N_5150,N_4560,N_3230);
nand U5151 (N_5151,N_3969,N_3795);
and U5152 (N_5152,N_4663,N_3253);
xnor U5153 (N_5153,N_4620,N_4023);
and U5154 (N_5154,N_4244,N_2766);
xor U5155 (N_5155,N_2532,N_3964);
or U5156 (N_5156,N_4724,N_4389);
nor U5157 (N_5157,N_2559,N_4622);
and U5158 (N_5158,N_2943,N_2743);
and U5159 (N_5159,N_3212,N_4759);
nand U5160 (N_5160,N_4796,N_3229);
xor U5161 (N_5161,N_2891,N_4304);
or U5162 (N_5162,N_3706,N_3531);
nand U5163 (N_5163,N_3790,N_3408);
nor U5164 (N_5164,N_2865,N_4199);
and U5165 (N_5165,N_4821,N_4981);
or U5166 (N_5166,N_4613,N_4269);
nand U5167 (N_5167,N_4847,N_4968);
and U5168 (N_5168,N_2861,N_2701);
nand U5169 (N_5169,N_4077,N_2586);
nand U5170 (N_5170,N_2831,N_4094);
and U5171 (N_5171,N_3939,N_2986);
or U5172 (N_5172,N_2977,N_3152);
nor U5173 (N_5173,N_2760,N_4243);
xor U5174 (N_5174,N_4528,N_3186);
nand U5175 (N_5175,N_3900,N_3590);
or U5176 (N_5176,N_3558,N_3775);
nand U5177 (N_5177,N_4226,N_2719);
nand U5178 (N_5178,N_3063,N_4362);
nand U5179 (N_5179,N_3277,N_4355);
or U5180 (N_5180,N_4615,N_4028);
and U5181 (N_5181,N_3249,N_4915);
nand U5182 (N_5182,N_3515,N_4055);
xnor U5183 (N_5183,N_4749,N_3050);
xnor U5184 (N_5184,N_2799,N_3816);
and U5185 (N_5185,N_4877,N_4364);
and U5186 (N_5186,N_3248,N_4419);
nand U5187 (N_5187,N_4802,N_2976);
xnor U5188 (N_5188,N_4381,N_3155);
or U5189 (N_5189,N_4401,N_3270);
nand U5190 (N_5190,N_3221,N_3265);
and U5191 (N_5191,N_3678,N_3165);
nor U5192 (N_5192,N_4888,N_3202);
xnor U5193 (N_5193,N_3910,N_3700);
and U5194 (N_5194,N_4511,N_3958);
nand U5195 (N_5195,N_4386,N_3581);
or U5196 (N_5196,N_3620,N_4918);
and U5197 (N_5197,N_4826,N_4913);
nand U5198 (N_5198,N_4089,N_4263);
xor U5199 (N_5199,N_4114,N_4046);
or U5200 (N_5200,N_4050,N_4747);
nor U5201 (N_5201,N_4251,N_4584);
xnor U5202 (N_5202,N_3318,N_4339);
xor U5203 (N_5203,N_2996,N_4000);
nand U5204 (N_5204,N_4861,N_2650);
xor U5205 (N_5205,N_4964,N_4075);
nor U5206 (N_5206,N_2611,N_3857);
or U5207 (N_5207,N_4363,N_3538);
nand U5208 (N_5208,N_4405,N_3220);
nand U5209 (N_5209,N_3345,N_2752);
nor U5210 (N_5210,N_3371,N_4372);
and U5211 (N_5211,N_2712,N_3708);
xor U5212 (N_5212,N_4149,N_3160);
nand U5213 (N_5213,N_3904,N_3084);
or U5214 (N_5214,N_3224,N_3320);
xor U5215 (N_5215,N_2787,N_4638);
nor U5216 (N_5216,N_3373,N_3114);
and U5217 (N_5217,N_4415,N_3029);
xnor U5218 (N_5218,N_4059,N_3086);
and U5219 (N_5219,N_3977,N_3859);
or U5220 (N_5220,N_3183,N_2671);
and U5221 (N_5221,N_3724,N_4880);
xnor U5222 (N_5222,N_4954,N_4911);
nor U5223 (N_5223,N_2654,N_3288);
xnor U5224 (N_5224,N_4676,N_2797);
nand U5225 (N_5225,N_3391,N_4882);
nand U5226 (N_5226,N_3846,N_3497);
or U5227 (N_5227,N_2552,N_4812);
nor U5228 (N_5228,N_3537,N_2715);
xor U5229 (N_5229,N_3750,N_3801);
and U5230 (N_5230,N_2568,N_4845);
xor U5231 (N_5231,N_3829,N_2932);
nor U5232 (N_5232,N_4478,N_4599);
and U5233 (N_5233,N_4716,N_4118);
nor U5234 (N_5234,N_3483,N_3276);
or U5235 (N_5235,N_4660,N_4991);
xor U5236 (N_5236,N_3313,N_4048);
nand U5237 (N_5237,N_4626,N_2515);
nand U5238 (N_5238,N_3612,N_2886);
and U5239 (N_5239,N_3254,N_4573);
nand U5240 (N_5240,N_4392,N_4217);
or U5241 (N_5241,N_4838,N_2500);
nor U5242 (N_5242,N_4898,N_4696);
nor U5243 (N_5243,N_4731,N_3019);
nand U5244 (N_5244,N_4298,N_2934);
nor U5245 (N_5245,N_4570,N_2714);
xnor U5246 (N_5246,N_2531,N_3412);
nand U5247 (N_5247,N_2579,N_3142);
xnor U5248 (N_5248,N_3000,N_4791);
nor U5249 (N_5249,N_4350,N_4755);
nand U5250 (N_5250,N_4196,N_4935);
and U5251 (N_5251,N_3299,N_2703);
nor U5252 (N_5252,N_2727,N_4894);
and U5253 (N_5253,N_4879,N_3210);
nand U5254 (N_5254,N_2692,N_3071);
or U5255 (N_5255,N_3582,N_4294);
and U5256 (N_5256,N_3560,N_3867);
and U5257 (N_5257,N_2666,N_2879);
xor U5258 (N_5258,N_4703,N_4941);
nand U5259 (N_5259,N_4066,N_4056);
or U5260 (N_5260,N_2900,N_4383);
nand U5261 (N_5261,N_3364,N_2520);
and U5262 (N_5262,N_3807,N_4139);
xnor U5263 (N_5263,N_3652,N_4130);
nand U5264 (N_5264,N_3135,N_4540);
nand U5265 (N_5265,N_3647,N_4578);
or U5266 (N_5266,N_4524,N_3832);
or U5267 (N_5267,N_4934,N_2768);
and U5268 (N_5268,N_3090,N_3246);
and U5269 (N_5269,N_3591,N_2991);
and U5270 (N_5270,N_4922,N_2670);
xnor U5271 (N_5271,N_4832,N_4268);
xnor U5272 (N_5272,N_3751,N_3550);
and U5273 (N_5273,N_2649,N_2643);
nor U5274 (N_5274,N_4612,N_3781);
nand U5275 (N_5275,N_3823,N_4623);
or U5276 (N_5276,N_2507,N_2504);
nand U5277 (N_5277,N_4673,N_3266);
and U5278 (N_5278,N_4980,N_4272);
nor U5279 (N_5279,N_2924,N_2616);
xnor U5280 (N_5280,N_4186,N_4016);
xor U5281 (N_5281,N_4788,N_4629);
xor U5282 (N_5282,N_3955,N_2518);
and U5283 (N_5283,N_2585,N_3727);
and U5284 (N_5284,N_2530,N_4969);
nand U5285 (N_5285,N_3243,N_2913);
and U5286 (N_5286,N_2882,N_4546);
or U5287 (N_5287,N_2624,N_4897);
or U5288 (N_5288,N_4448,N_2660);
xnor U5289 (N_5289,N_3319,N_2863);
or U5290 (N_5290,N_3132,N_3182);
nor U5291 (N_5291,N_2978,N_3919);
and U5292 (N_5292,N_3362,N_4591);
and U5293 (N_5293,N_4730,N_3517);
and U5294 (N_5294,N_3140,N_3765);
nor U5295 (N_5295,N_4722,N_4221);
nor U5296 (N_5296,N_3764,N_3961);
nor U5297 (N_5297,N_2810,N_4767);
xnor U5298 (N_5298,N_3281,N_2730);
nand U5299 (N_5299,N_4927,N_4471);
nor U5300 (N_5300,N_3956,N_3488);
nor U5301 (N_5301,N_3145,N_4571);
xnor U5302 (N_5302,N_4235,N_4018);
or U5303 (N_5303,N_4544,N_2794);
nand U5304 (N_5304,N_4958,N_2626);
or U5305 (N_5305,N_2808,N_4818);
xnor U5306 (N_5306,N_4736,N_3089);
nand U5307 (N_5307,N_3361,N_3709);
and U5308 (N_5308,N_4655,N_4495);
and U5309 (N_5309,N_3638,N_4204);
nand U5310 (N_5310,N_3689,N_2560);
or U5311 (N_5311,N_3987,N_4451);
nor U5312 (N_5312,N_3702,N_3520);
and U5313 (N_5313,N_3358,N_3197);
nor U5314 (N_5314,N_3736,N_3098);
nand U5315 (N_5315,N_3854,N_3255);
xnor U5316 (N_5316,N_3163,N_3830);
nand U5317 (N_5317,N_4387,N_2961);
nor U5318 (N_5318,N_3457,N_3081);
xnor U5319 (N_5319,N_2506,N_3038);
nand U5320 (N_5320,N_3476,N_4397);
xnor U5321 (N_5321,N_4764,N_4937);
nand U5322 (N_5322,N_3818,N_3321);
xnor U5323 (N_5323,N_3397,N_4208);
or U5324 (N_5324,N_3274,N_4956);
nor U5325 (N_5325,N_4423,N_3725);
xor U5326 (N_5326,N_3730,N_2689);
nand U5327 (N_5327,N_3100,N_4188);
or U5328 (N_5328,N_4943,N_2655);
or U5329 (N_5329,N_4010,N_3129);
nor U5330 (N_5330,N_2750,N_4301);
or U5331 (N_5331,N_3269,N_3162);
or U5332 (N_5332,N_3398,N_3913);
and U5333 (N_5333,N_4201,N_2584);
or U5334 (N_5334,N_3598,N_3027);
nand U5335 (N_5335,N_2514,N_4907);
xnor U5336 (N_5336,N_3635,N_2988);
and U5337 (N_5337,N_3267,N_4498);
or U5338 (N_5338,N_3597,N_4762);
nand U5339 (N_5339,N_4657,N_4293);
or U5340 (N_5340,N_3020,N_4848);
or U5341 (N_5341,N_2708,N_2704);
nand U5342 (N_5342,N_3676,N_4005);
nand U5343 (N_5343,N_4012,N_2509);
nand U5344 (N_5344,N_4097,N_4773);
nand U5345 (N_5345,N_4135,N_4532);
nand U5346 (N_5346,N_3005,N_2609);
and U5347 (N_5347,N_3174,N_2645);
nand U5348 (N_5348,N_3666,N_3012);
and U5349 (N_5349,N_3889,N_4705);
and U5350 (N_5350,N_4155,N_3720);
or U5351 (N_5351,N_3632,N_4311);
xor U5352 (N_5352,N_4500,N_4332);
nor U5353 (N_5353,N_4148,N_4265);
xnor U5354 (N_5354,N_3487,N_4462);
xor U5355 (N_5355,N_2821,N_4331);
nand U5356 (N_5356,N_2823,N_4190);
nand U5357 (N_5357,N_3514,N_4930);
or U5358 (N_5358,N_3438,N_3473);
nor U5359 (N_5359,N_4436,N_3331);
nand U5360 (N_5360,N_4480,N_3726);
nor U5361 (N_5361,N_3399,N_3437);
nor U5362 (N_5362,N_3381,N_3335);
or U5363 (N_5363,N_2904,N_3769);
xnor U5364 (N_5364,N_4275,N_3784);
and U5365 (N_5365,N_3585,N_3306);
nor U5366 (N_5366,N_2964,N_3450);
nor U5367 (N_5367,N_4729,N_4179);
and U5368 (N_5368,N_3699,N_4595);
nand U5369 (N_5369,N_4783,N_4926);
nand U5370 (N_5370,N_3744,N_3501);
nand U5371 (N_5371,N_4276,N_3732);
xor U5372 (N_5372,N_3568,N_3625);
nor U5373 (N_5373,N_4256,N_3349);
and U5374 (N_5374,N_4326,N_3116);
nor U5375 (N_5375,N_2925,N_4609);
xnor U5376 (N_5376,N_4957,N_4534);
nor U5377 (N_5377,N_3435,N_3203);
and U5378 (N_5378,N_4375,N_3353);
xor U5379 (N_5379,N_4670,N_4107);
or U5380 (N_5380,N_2930,N_4248);
nor U5381 (N_5381,N_2902,N_4414);
xnor U5382 (N_5382,N_4485,N_3687);
or U5383 (N_5383,N_3834,N_4766);
and U5384 (N_5384,N_3031,N_4640);
xnor U5385 (N_5385,N_2610,N_3018);
nor U5386 (N_5386,N_3646,N_3933);
or U5387 (N_5387,N_4588,N_4219);
nor U5388 (N_5388,N_4264,N_3559);
xor U5389 (N_5389,N_2950,N_3170);
or U5390 (N_5390,N_4806,N_4237);
or U5391 (N_5391,N_2982,N_2607);
nand U5392 (N_5392,N_4611,N_3095);
nand U5393 (N_5393,N_3989,N_4449);
nor U5394 (N_5394,N_3244,N_2889);
nand U5395 (N_5395,N_2756,N_4514);
nand U5396 (N_5396,N_4030,N_3561);
and U5397 (N_5397,N_3159,N_3528);
or U5398 (N_5398,N_2944,N_4765);
xor U5399 (N_5399,N_3139,N_4409);
xor U5400 (N_5400,N_3653,N_3870);
nand U5401 (N_5401,N_4651,N_2868);
nor U5402 (N_5402,N_3924,N_4662);
or U5403 (N_5403,N_4242,N_3684);
and U5404 (N_5404,N_4123,N_4049);
nor U5405 (N_5405,N_3701,N_4817);
nor U5406 (N_5406,N_3721,N_3766);
and U5407 (N_5407,N_4597,N_4677);
or U5408 (N_5408,N_4944,N_4688);
nor U5409 (N_5409,N_4580,N_4516);
nor U5410 (N_5410,N_4058,N_4711);
and U5411 (N_5411,N_2956,N_3273);
or U5412 (N_5412,N_2634,N_4999);
or U5413 (N_5413,N_3146,N_3665);
and U5414 (N_5414,N_4168,N_3149);
nand U5415 (N_5415,N_2574,N_4876);
and U5416 (N_5416,N_2517,N_2717);
xor U5417 (N_5417,N_4792,N_3475);
and U5418 (N_5418,N_3192,N_4337);
xnor U5419 (N_5419,N_3604,N_4508);
nor U5420 (N_5420,N_4177,N_3908);
nor U5421 (N_5421,N_2580,N_4738);
and U5422 (N_5422,N_3396,N_4349);
or U5423 (N_5423,N_3845,N_4176);
and U5424 (N_5424,N_2674,N_3588);
or U5425 (N_5425,N_2647,N_3452);
xor U5426 (N_5426,N_4851,N_3417);
nand U5427 (N_5427,N_3912,N_4671);
xor U5428 (N_5428,N_3057,N_2576);
nand U5429 (N_5429,N_4283,N_4554);
or U5430 (N_5430,N_3562,N_4921);
xnor U5431 (N_5431,N_4784,N_2818);
and U5432 (N_5432,N_2765,N_2851);
and U5433 (N_5433,N_2641,N_2613);
or U5434 (N_5434,N_4108,N_4220);
nor U5435 (N_5435,N_2640,N_4608);
nand U5436 (N_5436,N_3849,N_2842);
and U5437 (N_5437,N_2522,N_2562);
nor U5438 (N_5438,N_2505,N_4105);
xnor U5439 (N_5439,N_4754,N_3677);
and U5440 (N_5440,N_3905,N_3176);
or U5441 (N_5441,N_4195,N_4833);
xor U5442 (N_5442,N_2524,N_2774);
nand U5443 (N_5443,N_4704,N_3102);
nand U5444 (N_5444,N_3006,N_3606);
nand U5445 (N_5445,N_2916,N_4442);
xnor U5446 (N_5446,N_3885,N_2696);
nand U5447 (N_5447,N_4316,N_4564);
and U5448 (N_5448,N_4253,N_3378);
nand U5449 (N_5449,N_3740,N_3634);
and U5450 (N_5450,N_4706,N_3662);
and U5451 (N_5451,N_2816,N_3066);
and U5452 (N_5452,N_2577,N_4682);
and U5453 (N_5453,N_4473,N_3997);
nor U5454 (N_5454,N_3555,N_2917);
and U5455 (N_5455,N_2566,N_3040);
nor U5456 (N_5456,N_4052,N_2521);
or U5457 (N_5457,N_3541,N_3138);
nor U5458 (N_5458,N_3099,N_4280);
nor U5459 (N_5459,N_4403,N_3251);
xor U5460 (N_5460,N_3868,N_3400);
xor U5461 (N_5461,N_4230,N_4854);
or U5462 (N_5462,N_4134,N_4446);
nor U5463 (N_5463,N_3257,N_4970);
nand U5464 (N_5464,N_2602,N_4065);
xnor U5465 (N_5465,N_2694,N_4649);
nor U5466 (N_5466,N_4082,N_2815);
or U5467 (N_5467,N_3204,N_4798);
nand U5468 (N_5468,N_4659,N_3573);
nand U5469 (N_5469,N_4819,N_3445);
nor U5470 (N_5470,N_4537,N_3072);
xnor U5471 (N_5471,N_3119,N_3745);
xnor U5472 (N_5472,N_3941,N_4153);
xor U5473 (N_5473,N_3154,N_2652);
or U5474 (N_5474,N_3366,N_4656);
and U5475 (N_5475,N_4015,N_4240);
nor U5476 (N_5476,N_4189,N_3068);
nor U5477 (N_5477,N_2608,N_3172);
nand U5478 (N_5478,N_2646,N_4575);
or U5479 (N_5479,N_3236,N_4940);
and U5480 (N_5480,N_3636,N_3292);
or U5481 (N_5481,N_4557,N_3394);
xor U5482 (N_5482,N_3519,N_3540);
xnor U5483 (N_5483,N_4122,N_4101);
nor U5484 (N_5484,N_3860,N_3015);
nand U5485 (N_5485,N_3498,N_2931);
xor U5486 (N_5486,N_3828,N_2575);
nor U5487 (N_5487,N_3595,N_3026);
xor U5488 (N_5488,N_3075,N_4856);
nor U5489 (N_5489,N_3432,N_3906);
xnor U5490 (N_5490,N_3770,N_2909);
and U5491 (N_5491,N_4795,N_4840);
and U5492 (N_5492,N_2665,N_4691);
xor U5493 (N_5493,N_2600,N_3078);
nand U5494 (N_5494,N_3518,N_3754);
nand U5495 (N_5495,N_2711,N_4175);
or U5496 (N_5496,N_4062,N_4333);
and U5497 (N_5497,N_2663,N_4535);
xnor U5498 (N_5498,N_2728,N_3064);
or U5499 (N_5499,N_3499,N_4324);
nor U5500 (N_5500,N_4126,N_3694);
or U5501 (N_5501,N_4689,N_3205);
and U5502 (N_5502,N_3982,N_4665);
or U5503 (N_5503,N_3351,N_2839);
xor U5504 (N_5504,N_4239,N_3472);
nand U5505 (N_5505,N_2721,N_3053);
nor U5506 (N_5506,N_3434,N_2793);
or U5507 (N_5507,N_4022,N_3570);
nand U5508 (N_5508,N_3670,N_3307);
nand U5509 (N_5509,N_4931,N_2806);
nor U5510 (N_5510,N_4561,N_3045);
nand U5511 (N_5511,N_3546,N_3180);
and U5512 (N_5512,N_2967,N_3271);
nand U5513 (N_5513,N_3263,N_4367);
xor U5514 (N_5514,N_2918,N_3168);
nand U5515 (N_5515,N_3864,N_2805);
xnor U5516 (N_5516,N_4447,N_4757);
nor U5517 (N_5517,N_3629,N_3521);
nor U5518 (N_5518,N_4685,N_2829);
nor U5519 (N_5519,N_3978,N_3505);
nor U5520 (N_5520,N_3003,N_4305);
xor U5521 (N_5521,N_3793,N_3685);
and U5522 (N_5522,N_3136,N_3664);
nand U5523 (N_5523,N_3308,N_4600);
nand U5524 (N_5524,N_4421,N_2673);
or U5525 (N_5525,N_4972,N_4063);
xor U5526 (N_5526,N_3548,N_3596);
xor U5527 (N_5527,N_4746,N_4216);
nand U5528 (N_5528,N_3663,N_2948);
nor U5529 (N_5529,N_3363,N_2588);
or U5530 (N_5530,N_4912,N_3014);
and U5531 (N_5531,N_4828,N_2878);
nand U5532 (N_5532,N_4996,N_2820);
nand U5533 (N_5533,N_3847,N_3094);
xnor U5534 (N_5534,N_2817,N_4959);
xor U5535 (N_5535,N_3150,N_3324);
or U5536 (N_5536,N_3863,N_3480);
xnor U5537 (N_5537,N_3618,N_4618);
and U5538 (N_5538,N_4562,N_3347);
nand U5539 (N_5539,N_4070,N_2847);
nor U5540 (N_5540,N_4131,N_3675);
xnor U5541 (N_5541,N_4115,N_4034);
nor U5542 (N_5542,N_3763,N_4025);
xor U5543 (N_5543,N_4831,N_3315);
xnor U5544 (N_5544,N_4306,N_2619);
and U5545 (N_5545,N_4503,N_4300);
or U5546 (N_5546,N_4110,N_3580);
nor U5547 (N_5547,N_4088,N_4120);
or U5548 (N_5548,N_4371,N_4290);
or U5549 (N_5549,N_4281,N_4112);
nand U5550 (N_5550,N_3252,N_4661);
and U5551 (N_5551,N_3477,N_3039);
and U5552 (N_5552,N_4042,N_4901);
or U5553 (N_5553,N_4890,N_4510);
xor U5554 (N_5554,N_4047,N_3798);
xor U5555 (N_5555,N_3028,N_3346);
and U5556 (N_5556,N_4061,N_4254);
or U5557 (N_5557,N_4329,N_4533);
or U5558 (N_5558,N_4553,N_4072);
nand U5559 (N_5559,N_4287,N_3333);
nor U5560 (N_5560,N_2875,N_3876);
or U5561 (N_5561,N_4642,N_3681);
or U5562 (N_5562,N_3869,N_4357);
or U5563 (N_5563,N_4418,N_4003);
and U5564 (N_5564,N_3525,N_2551);
or U5565 (N_5565,N_4464,N_4238);
xnor U5566 (N_5566,N_2993,N_3231);
nand U5567 (N_5567,N_2937,N_4466);
xnor U5568 (N_5568,N_4267,N_3446);
or U5569 (N_5569,N_3564,N_3865);
nor U5570 (N_5570,N_4151,N_3718);
and U5571 (N_5571,N_4774,N_3046);
or U5572 (N_5572,N_3280,N_3545);
and U5573 (N_5573,N_3283,N_4487);
or U5574 (N_5574,N_3387,N_4270);
and U5575 (N_5575,N_4631,N_4430);
or U5576 (N_5576,N_2606,N_4645);
nand U5577 (N_5577,N_3384,N_2858);
xor U5578 (N_5578,N_3565,N_3690);
nand U5579 (N_5579,N_3741,N_2603);
nand U5580 (N_5580,N_3256,N_3194);
and U5581 (N_5581,N_4872,N_4214);
nand U5582 (N_5582,N_4865,N_3619);
nor U5583 (N_5583,N_4914,N_3388);
nand U5584 (N_5584,N_3310,N_3866);
or U5585 (N_5585,N_3772,N_4407);
nand U5586 (N_5586,N_2777,N_3443);
or U5587 (N_5587,N_2519,N_2748);
nor U5588 (N_5588,N_4908,N_4497);
or U5589 (N_5589,N_4282,N_2561);
nand U5590 (N_5590,N_4929,N_3536);
nor U5591 (N_5591,N_3926,N_4881);
and U5592 (N_5592,N_4111,N_3376);
and U5593 (N_5593,N_4804,N_2947);
nor U5594 (N_5594,N_3164,N_3493);
nand U5595 (N_5595,N_3106,N_4949);
nand U5596 (N_5596,N_3083,N_4024);
nor U5597 (N_5597,N_4157,N_3787);
or U5598 (N_5598,N_4603,N_2940);
xor U5599 (N_5599,N_3056,N_2734);
nand U5600 (N_5600,N_3237,N_4950);
and U5601 (N_5601,N_4545,N_3882);
and U5602 (N_5602,N_3593,N_4370);
and U5603 (N_5603,N_4694,N_2995);
or U5604 (N_5604,N_4786,N_3757);
xor U5605 (N_5605,N_3626,N_3217);
nor U5606 (N_5606,N_2677,N_4093);
or U5607 (N_5607,N_3242,N_4982);
xnor U5608 (N_5608,N_2843,N_4875);
xor U5609 (N_5609,N_4539,N_3713);
and U5610 (N_5610,N_3342,N_4810);
xor U5611 (N_5611,N_4031,N_2786);
nor U5612 (N_5612,N_3788,N_4325);
and U5613 (N_5613,N_3502,N_3339);
and U5614 (N_5614,N_2804,N_2958);
nor U5615 (N_5615,N_4225,N_4292);
xor U5616 (N_5616,N_3547,N_3756);
nand U5617 (N_5617,N_2959,N_3268);
xor U5618 (N_5618,N_3586,N_4079);
xor U5619 (N_5619,N_3747,N_2901);
nor U5620 (N_5620,N_2601,N_4493);
nor U5621 (N_5621,N_4099,N_3753);
nand U5622 (N_5622,N_2581,N_4132);
and U5623 (N_5623,N_4919,N_2512);
or U5624 (N_5624,N_3780,N_3322);
nand U5625 (N_5625,N_3609,N_2919);
and U5626 (N_5626,N_3911,N_4021);
or U5627 (N_5627,N_3973,N_2563);
or U5628 (N_5628,N_4038,N_4548);
nand U5629 (N_5629,N_3907,N_4013);
nor U5630 (N_5630,N_3851,N_3717);
nand U5631 (N_5631,N_4484,N_2687);
or U5632 (N_5632,N_3264,N_2658);
and U5633 (N_5633,N_2557,N_4576);
and U5634 (N_5634,N_2604,N_2775);
xor U5635 (N_5635,N_3848,N_3213);
xor U5636 (N_5636,N_2702,N_4100);
and U5637 (N_5637,N_4527,N_3447);
xnor U5638 (N_5638,N_4587,N_4037);
nand U5639 (N_5639,N_3841,N_4910);
nand U5640 (N_5640,N_3552,N_4259);
nor U5641 (N_5641,N_4102,N_3527);
and U5642 (N_5642,N_4946,N_2541);
nand U5643 (N_5643,N_3103,N_4181);
and U5644 (N_5644,N_2642,N_2632);
xnor U5645 (N_5645,N_2565,N_2644);
nand U5646 (N_5646,N_4162,N_4947);
or U5647 (N_5647,N_3729,N_3760);
xnor U5648 (N_5648,N_2824,N_4222);
and U5649 (N_5649,N_4076,N_4129);
or U5650 (N_5650,N_4338,N_3644);
nand U5651 (N_5651,N_4435,N_3465);
nor U5652 (N_5652,N_4207,N_4127);
xnor U5653 (N_5653,N_3971,N_3572);
xnor U5654 (N_5654,N_2622,N_3052);
and U5655 (N_5655,N_4807,N_3413);
nand U5656 (N_5656,N_4771,N_4017);
xnor U5657 (N_5657,N_3921,N_3556);
nor U5658 (N_5658,N_2598,N_3783);
and U5659 (N_5659,N_3522,N_3372);
xnor U5660 (N_5660,N_3508,N_3986);
and U5661 (N_5661,N_2567,N_2618);
nor U5662 (N_5662,N_2587,N_4180);
nor U5663 (N_5663,N_3992,N_3861);
or U5664 (N_5664,N_2899,N_3120);
nor U5665 (N_5665,N_3785,N_2782);
xnor U5666 (N_5666,N_4710,N_3909);
nand U5667 (N_5667,N_3074,N_4057);
and U5668 (N_5668,N_4945,N_3425);
nand U5669 (N_5669,N_4650,N_3036);
or U5670 (N_5670,N_4352,N_3683);
nor U5671 (N_5671,N_4809,N_2933);
nor U5672 (N_5672,N_2596,N_4517);
nor U5673 (N_5673,N_3298,N_2962);
and U5674 (N_5674,N_3965,N_3478);
and U5675 (N_5675,N_3507,N_4785);
or U5676 (N_5676,N_4133,N_3884);
nand U5677 (N_5677,N_3668,N_4823);
or U5678 (N_5678,N_2526,N_4942);
xnor U5679 (N_5679,N_3406,N_4143);
nand U5680 (N_5680,N_3778,N_2753);
or U5681 (N_5681,N_2848,N_3567);
or U5682 (N_5682,N_3044,N_2630);
xnor U5683 (N_5683,N_3890,N_3385);
nand U5684 (N_5684,N_4748,N_3831);
or U5685 (N_5685,N_3196,N_2735);
nand U5686 (N_5686,N_3946,N_4092);
or U5687 (N_5687,N_4334,N_3943);
xnor U5688 (N_5688,N_4170,N_3025);
and U5689 (N_5689,N_4218,N_3762);
nor U5690 (N_5690,N_4310,N_3688);
or U5691 (N_5691,N_3087,N_3738);
nor U5692 (N_5692,N_3962,N_4614);
nor U5693 (N_5693,N_4728,N_4583);
xnor U5694 (N_5694,N_2942,N_3972);
xnor U5695 (N_5695,N_4952,N_3633);
or U5696 (N_5696,N_4652,N_3948);
nand U5697 (N_5697,N_3672,N_3177);
and U5698 (N_5698,N_4278,N_4753);
xor U5699 (N_5699,N_3047,N_3055);
and U5700 (N_5700,N_3658,N_4249);
nor U5701 (N_5701,N_4636,N_3357);
and U5702 (N_5702,N_4646,N_4574);
or U5703 (N_5703,N_2617,N_4678);
xor U5704 (N_5704,N_4827,N_3809);
xnor U5705 (N_5705,N_4633,N_4707);
nand U5706 (N_5706,N_3228,N_3934);
nor U5707 (N_5707,N_3037,N_4158);
and U5708 (N_5708,N_3862,N_4224);
or U5709 (N_5709,N_4522,N_4160);
xnor U5710 (N_5710,N_4006,N_4427);
xnor U5711 (N_5711,N_4836,N_4715);
nand U5712 (N_5712,N_4002,N_2593);
and U5713 (N_5713,N_4318,N_3466);
or U5714 (N_5714,N_2540,N_3069);
and U5715 (N_5715,N_2972,N_4979);
nand U5716 (N_5716,N_2740,N_3563);
nand U5717 (N_5717,N_4011,N_3316);
or U5718 (N_5718,N_2809,N_4758);
or U5719 (N_5719,N_3314,N_4455);
nand U5720 (N_5720,N_3815,N_2814);
nor U5721 (N_5721,N_3839,N_3840);
nor U5722 (N_5722,N_4406,N_4549);
nor U5723 (N_5723,N_4104,N_3950);
or U5724 (N_5724,N_3737,N_3615);
and U5725 (N_5725,N_2915,N_4335);
nand U5726 (N_5726,N_4069,N_3016);
nor U5727 (N_5727,N_3894,N_4700);
xnor U5728 (N_5728,N_3628,N_3600);
xnor U5729 (N_5729,N_4739,N_4844);
nor U5730 (N_5730,N_4752,N_4014);
nand U5731 (N_5731,N_3287,N_3080);
nand U5732 (N_5732,N_4988,N_3082);
or U5733 (N_5733,N_2758,N_2914);
xor U5734 (N_5734,N_3878,N_3474);
and U5735 (N_5735,N_4161,N_4607);
nor U5736 (N_5736,N_4117,N_2893);
xor U5737 (N_5737,N_3805,N_3455);
or U5738 (N_5738,N_3463,N_4727);
and U5739 (N_5739,N_3833,N_4610);
xnor U5740 (N_5740,N_3858,N_4183);
xnor U5741 (N_5741,N_2569,N_3822);
or U5742 (N_5742,N_4951,N_3566);
or U5743 (N_5743,N_3272,N_3991);
nor U5744 (N_5744,N_2939,N_3603);
xor U5745 (N_5745,N_3416,N_3542);
xor U5746 (N_5746,N_3856,N_2558);
or U5747 (N_5747,N_4813,N_2846);
nor U5748 (N_5748,N_3963,N_2983);
nand U5749 (N_5749,N_3735,N_3746);
xor U5750 (N_5750,N_2906,N_4874);
nand U5751 (N_5751,N_4479,N_4630);
nor U5752 (N_5752,N_4916,N_2657);
or U5753 (N_5753,N_2871,N_3693);
or U5754 (N_5754,N_3070,N_4289);
nor U5755 (N_5755,N_4761,N_4074);
nor U5756 (N_5756,N_3420,N_4518);
and U5757 (N_5757,N_4044,N_3021);
nor U5758 (N_5758,N_4086,N_4852);
or U5759 (N_5759,N_3917,N_3960);
or U5760 (N_5760,N_4596,N_3813);
or U5761 (N_5761,N_4743,N_3569);
and U5762 (N_5762,N_2725,N_3091);
or U5763 (N_5763,N_4428,N_4273);
and U5764 (N_5764,N_3076,N_4816);
or U5765 (N_5765,N_4027,N_3886);
or U5766 (N_5766,N_2923,N_3605);
and U5767 (N_5767,N_3427,N_4393);
and U5768 (N_5768,N_3088,N_4445);
and U5769 (N_5769,N_4174,N_2767);
nor U5770 (N_5770,N_3184,N_4602);
xnor U5771 (N_5771,N_4429,N_3424);
nor U5772 (N_5772,N_3985,N_4441);
and U5773 (N_5773,N_4453,N_4211);
xor U5774 (N_5774,N_4869,N_4271);
nand U5775 (N_5775,N_4974,N_4463);
and U5776 (N_5776,N_3326,N_2825);
xor U5777 (N_5777,N_4091,N_2785);
xor U5778 (N_5778,N_4474,N_4672);
nand U5779 (N_5779,N_3395,N_4443);
nand U5780 (N_5780,N_2761,N_4643);
xnor U5781 (N_5781,N_3215,N_3641);
xor U5782 (N_5782,N_2869,N_2975);
and U5783 (N_5783,N_3291,N_3711);
xnor U5784 (N_5784,N_4863,N_4904);
xnor U5785 (N_5785,N_2867,N_3440);
and U5786 (N_5786,N_2973,N_4492);
or U5787 (N_5787,N_3631,N_4841);
or U5788 (N_5788,N_4203,N_3959);
or U5789 (N_5789,N_4344,N_3549);
xor U5790 (N_5790,N_3928,N_3195);
or U5791 (N_5791,N_4358,N_4878);
nor U5792 (N_5792,N_3377,N_4060);
nor U5793 (N_5793,N_2739,N_4080);
nor U5794 (N_5794,N_4531,N_2897);
nand U5795 (N_5795,N_4145,N_2686);
nor U5796 (N_5796,N_3679,N_4470);
nor U5797 (N_5797,N_4402,N_2710);
or U5798 (N_5798,N_4928,N_2790);
xnor U5799 (N_5799,N_4399,N_3835);
and U5800 (N_5800,N_4246,N_2720);
and U5801 (N_5801,N_2826,N_3187);
nand U5802 (N_5802,N_2583,N_3655);
nand U5803 (N_5803,N_3947,N_3723);
nor U5804 (N_5804,N_4041,N_2929);
nand U5805 (N_5805,N_3367,N_2907);
or U5806 (N_5806,N_4469,N_4735);
nor U5807 (N_5807,N_4889,N_2690);
and U5808 (N_5808,N_2688,N_2890);
xnor U5809 (N_5809,N_4348,N_4067);
nor U5810 (N_5810,N_4740,N_4228);
nor U5811 (N_5811,N_4563,N_2838);
nand U5812 (N_5812,N_4489,N_4920);
xor U5813 (N_5813,N_4147,N_2718);
and U5814 (N_5814,N_4345,N_3214);
nand U5815 (N_5815,N_2908,N_3650);
and U5816 (N_5816,N_3748,N_3574);
or U5817 (N_5817,N_3262,N_4347);
or U5818 (N_5818,N_2628,N_3578);
or U5819 (N_5819,N_3639,N_3422);
and U5820 (N_5820,N_2954,N_4683);
xnor U5821 (N_5821,N_2534,N_3459);
and U5822 (N_5822,N_3009,N_3587);
xor U5823 (N_5823,N_2691,N_4033);
nand U5824 (N_5824,N_4566,N_4185);
or U5825 (N_5825,N_2527,N_2669);
and U5826 (N_5826,N_3222,N_2638);
or U5827 (N_5827,N_3096,N_3017);
xor U5828 (N_5828,N_4103,N_4734);
nor U5829 (N_5829,N_3880,N_2672);
and U5830 (N_5830,N_4984,N_3410);
or U5831 (N_5831,N_4541,N_4439);
and U5832 (N_5832,N_2802,N_2757);
and U5833 (N_5833,N_4977,N_4150);
nand U5834 (N_5834,N_3444,N_4262);
or U5835 (N_5835,N_4396,N_3279);
or U5836 (N_5836,N_4975,N_3624);
and U5837 (N_5837,N_3393,N_2992);
and U5838 (N_5838,N_4020,N_3008);
nor U5839 (N_5839,N_4760,N_2985);
and U5840 (N_5840,N_3227,N_4223);
nor U5841 (N_5841,N_3853,N_3509);
or U5842 (N_5842,N_2864,N_3660);
nand U5843 (N_5843,N_3143,N_2796);
nand U5844 (N_5844,N_2892,N_4789);
nand U5845 (N_5845,N_4043,N_4353);
or U5846 (N_5846,N_3125,N_2737);
nor U5847 (N_5847,N_4895,N_3336);
xnor U5848 (N_5848,N_2564,N_4592);
and U5849 (N_5849,N_4322,N_3952);
nor U5850 (N_5850,N_4862,N_4045);
nor U5851 (N_5851,N_4504,N_4756);
xnor U5852 (N_5852,N_3804,N_4658);
and U5853 (N_5853,N_3993,N_2905);
or U5854 (N_5854,N_4398,N_4366);
and U5855 (N_5855,N_4004,N_4116);
nor U5856 (N_5856,N_3611,N_4547);
nor U5857 (N_5857,N_2571,N_4231);
and U5858 (N_5858,N_3436,N_3289);
or U5859 (N_5859,N_4330,N_3539);
or U5860 (N_5860,N_4779,N_3042);
or U5861 (N_5861,N_4083,N_3553);
xor U5862 (N_5862,N_3776,N_4559);
nand U5863 (N_5863,N_4702,N_4855);
or U5864 (N_5864,N_2597,N_4459);
nand U5865 (N_5865,N_3109,N_3686);
or U5866 (N_5866,N_4647,N_4274);
xor U5867 (N_5867,N_4742,N_4725);
and U5868 (N_5868,N_2555,N_4719);
nand U5869 (N_5869,N_4834,N_2920);
or U5870 (N_5870,N_2599,N_4717);
nand U5871 (N_5871,N_2676,N_2741);
nor U5872 (N_5872,N_4708,N_4590);
nand U5873 (N_5873,N_2781,N_2911);
xor U5874 (N_5874,N_3523,N_4302);
or U5875 (N_5875,N_4509,N_2661);
nor U5876 (N_5876,N_4472,N_4701);
nor U5877 (N_5877,N_3442,N_2834);
nor U5878 (N_5878,N_2549,N_2859);
or U5879 (N_5879,N_3414,N_3439);
nor U5880 (N_5880,N_4842,N_3337);
and U5881 (N_5881,N_3535,N_4679);
nand U5882 (N_5882,N_3996,N_3118);
xor U5883 (N_5883,N_3127,N_2749);
xor U5884 (N_5884,N_3529,N_2938);
nor U5885 (N_5885,N_3233,N_3481);
and U5886 (N_5886,N_3239,N_4291);
or U5887 (N_5887,N_4605,N_3661);
nand U5888 (N_5888,N_2738,N_3714);
and U5889 (N_5889,N_3380,N_2881);
and U5890 (N_5890,N_3797,N_4790);
nor U5891 (N_5891,N_4843,N_4637);
nand U5892 (N_5892,N_3657,N_4178);
nor U5893 (N_5893,N_3329,N_4870);
nand U5894 (N_5894,N_4299,N_2662);
xnor U5895 (N_5895,N_3193,N_3627);
nor U5896 (N_5896,N_4377,N_4312);
or U5897 (N_5897,N_4737,N_2966);
xnor U5898 (N_5898,N_3033,N_3383);
or U5899 (N_5899,N_4507,N_4720);
and U5900 (N_5900,N_3931,N_3207);
and U5901 (N_5901,N_4775,N_3179);
and U5902 (N_5902,N_4279,N_2747);
nor U5903 (N_5903,N_4732,N_3297);
nor U5904 (N_5904,N_4799,N_2898);
nor U5905 (N_5905,N_4594,N_3386);
nor U5906 (N_5906,N_4432,N_4903);
xnor U5907 (N_5907,N_4681,N_3843);
and U5908 (N_5908,N_2755,N_3206);
xnor U5909 (N_5909,N_4751,N_3035);
nor U5910 (N_5910,N_4090,N_4938);
xnor U5911 (N_5911,N_3317,N_2912);
xnor U5912 (N_5912,N_3312,N_2836);
or U5913 (N_5913,N_2529,N_3613);
and U5914 (N_5914,N_4936,N_4961);
xor U5915 (N_5915,N_3836,N_4628);
nand U5916 (N_5916,N_3871,N_4543);
nand U5917 (N_5917,N_4154,N_4288);
nand U5918 (N_5918,N_2827,N_2840);
nor U5919 (N_5919,N_4209,N_3350);
nand U5920 (N_5920,N_4939,N_2855);
xor U5921 (N_5921,N_3328,N_2866);
nor U5922 (N_5922,N_4198,N_3284);
xnor U5923 (N_5923,N_4457,N_3719);
or U5924 (N_5924,N_3225,N_2926);
and U5925 (N_5925,N_4585,N_4669);
nor U5926 (N_5926,N_2927,N_3285);
and U5927 (N_5927,N_3241,N_4835);
nor U5928 (N_5928,N_3806,N_3238);
nor U5929 (N_5929,N_4314,N_2884);
nor U5930 (N_5930,N_2578,N_4361);
and U5931 (N_5931,N_3936,N_3643);
nor U5932 (N_5932,N_4512,N_4001);
nand U5933 (N_5933,N_3311,N_3218);
nor U5934 (N_5934,N_2990,N_3247);
nor U5935 (N_5935,N_4925,N_4745);
and U5936 (N_5936,N_3630,N_2546);
or U5937 (N_5937,N_3108,N_3811);
and U5938 (N_5938,N_2535,N_3777);
xor U5939 (N_5939,N_3226,N_4163);
and U5940 (N_5940,N_3892,N_2860);
nor U5941 (N_5941,N_3872,N_3147);
nor U5942 (N_5942,N_2951,N_4285);
nand U5943 (N_5943,N_3208,N_4635);
and U5944 (N_5944,N_4948,N_4581);
xor U5945 (N_5945,N_4187,N_4354);
or U5946 (N_5946,N_3875,N_4883);
and U5947 (N_5947,N_4369,N_4675);
nor U5948 (N_5948,N_2678,N_4073);
xor U5949 (N_5949,N_2963,N_4800);
xor U5950 (N_5950,N_4128,N_4395);
nand U5951 (N_5951,N_3124,N_2791);
nand U5952 (N_5952,N_4258,N_4787);
nor U5953 (N_5953,N_3825,N_4604);
xnor U5954 (N_5954,N_4542,N_3901);
and U5955 (N_5955,N_3061,N_3323);
or U5956 (N_5956,N_3258,N_2998);
and U5957 (N_5957,N_2516,N_3161);
nand U5958 (N_5958,N_2706,N_3448);
and U5959 (N_5959,N_4718,N_4191);
nand U5960 (N_5960,N_2682,N_4194);
or U5961 (N_5961,N_4973,N_4985);
or U5962 (N_5962,N_3789,N_2589);
or U5963 (N_5963,N_4714,N_4071);
and U5964 (N_5964,N_4805,N_3697);
or U5965 (N_5965,N_4515,N_2837);
nor U5966 (N_5966,N_2501,N_2819);
nor U5967 (N_5967,N_3888,N_4106);
nand U5968 (N_5968,N_4245,N_3802);
nand U5969 (N_5969,N_3278,N_3874);
nor U5970 (N_5970,N_4617,N_2778);
and U5971 (N_5971,N_2856,N_2698);
nor U5972 (N_5972,N_3235,N_2615);
and U5973 (N_5973,N_2675,N_3504);
nor U5974 (N_5974,N_4589,N_2876);
xnor U5975 (N_5975,N_4822,N_4586);
or U5976 (N_5976,N_2724,N_4550);
or U5977 (N_5977,N_2592,N_4741);
and U5978 (N_5978,N_3173,N_4286);
nand U5979 (N_5979,N_2538,N_3300);
nor U5980 (N_5980,N_4565,N_3599);
nand U5981 (N_5981,N_3774,N_2709);
xnor U5982 (N_5982,N_2668,N_3348);
or U5983 (N_5983,N_4801,N_3153);
xor U5984 (N_5984,N_4966,N_3489);
xnor U5985 (N_5985,N_4692,N_4526);
nand U5986 (N_5986,N_4962,N_3392);
and U5987 (N_5987,N_3935,N_3827);
or U5988 (N_5988,N_4054,N_3355);
xor U5989 (N_5989,N_4412,N_4440);
xnor U5990 (N_5990,N_3404,N_3543);
xor U5991 (N_5991,N_4750,N_4095);
xnor U5992 (N_5992,N_4438,N_3467);
and U5993 (N_5993,N_2885,N_3121);
and U5994 (N_5994,N_4351,N_4297);
nor U5995 (N_5995,N_2707,N_4693);
xnor U5996 (N_5996,N_3013,N_4465);
nand U5997 (N_5997,N_3092,N_3855);
and U5998 (N_5998,N_2763,N_3844);
nand U5999 (N_5999,N_3601,N_3259);
or U6000 (N_6000,N_3137,N_3468);
nor U6001 (N_6001,N_3966,N_4811);
xnor U6002 (N_6002,N_4976,N_2700);
or U6003 (N_6003,N_4867,N_4712);
nand U6004 (N_6004,N_2874,N_4697);
or U6005 (N_6005,N_4036,N_4426);
and U6006 (N_6006,N_2813,N_2533);
xor U6007 (N_6007,N_4776,N_3428);
or U6008 (N_6008,N_4411,N_3998);
nand U6009 (N_6009,N_3768,N_3698);
nor U6010 (N_6010,N_2987,N_4172);
nand U6011 (N_6011,N_4530,N_3500);
xnor U6012 (N_6012,N_2946,N_3918);
nor U6013 (N_6013,N_4140,N_3097);
nand U6014 (N_6014,N_2945,N_4499);
or U6015 (N_6015,N_2545,N_2841);
xnor U6016 (N_6016,N_3341,N_3557);
nor U6017 (N_6017,N_4814,N_4680);
or U6018 (N_6018,N_4830,N_3691);
and U6019 (N_6019,N_3938,N_3616);
or U6020 (N_6020,N_4260,N_3703);
nand U6021 (N_6021,N_2949,N_2503);
nor U6022 (N_6022,N_4551,N_3303);
and U6023 (N_6023,N_4772,N_3742);
xnor U6024 (N_6024,N_4770,N_3877);
and U6025 (N_6025,N_4152,N_4803);
nand U6026 (N_6026,N_3301,N_3166);
or U6027 (N_6027,N_3980,N_3937);
nand U6028 (N_6028,N_2970,N_4990);
or U6029 (N_6029,N_3030,N_3524);
nand U6030 (N_6030,N_3511,N_4313);
nor U6031 (N_6031,N_2629,N_4698);
nand U6032 (N_6032,N_4373,N_4978);
or U6033 (N_6033,N_4136,N_4205);
xnor U6034 (N_6034,N_3001,N_3158);
xnor U6035 (N_6035,N_3093,N_2736);
nand U6036 (N_6036,N_4960,N_4648);
nand U6037 (N_6037,N_2683,N_4893);
nand U6038 (N_6038,N_4520,N_4993);
xor U6039 (N_6039,N_4873,N_2936);
xnor U6040 (N_6040,N_3883,N_3637);
and U6041 (N_6041,N_4142,N_2921);
xnor U6042 (N_6042,N_3513,N_2822);
nand U6043 (N_6043,N_4124,N_4359);
nor U6044 (N_6044,N_3617,N_3716);
xor U6045 (N_6045,N_4829,N_4619);
nand U6046 (N_6046,N_3988,N_4213);
and U6047 (N_6047,N_3669,N_4763);
nor U6048 (N_6048,N_4064,N_2759);
nand U6049 (N_6049,N_2852,N_3533);
and U6050 (N_6050,N_4579,N_4113);
or U6051 (N_6051,N_4641,N_3571);
nor U6052 (N_6052,N_4853,N_3275);
and U6053 (N_6053,N_2989,N_4009);
and U6054 (N_6054,N_2880,N_2779);
nor U6055 (N_6055,N_3199,N_2771);
or U6056 (N_6056,N_3914,N_3577);
nor U6057 (N_6057,N_3107,N_3043);
nor U6058 (N_6058,N_4266,N_4137);
or U6059 (N_6059,N_3842,N_3506);
xnor U6060 (N_6060,N_3837,N_4494);
xor U6061 (N_6061,N_3659,N_2894);
and U6062 (N_6062,N_4502,N_2525);
nand U6063 (N_6063,N_2769,N_3344);
nand U6064 (N_6064,N_4422,N_3903);
nand U6065 (N_6065,N_4096,N_2681);
nor U6066 (N_6066,N_4505,N_4336);
xnor U6067 (N_6067,N_4793,N_2570);
or U6068 (N_6068,N_4146,N_2746);
or U6069 (N_6069,N_3141,N_3608);
xor U6070 (N_6070,N_2984,N_2572);
nor U6071 (N_6071,N_2971,N_3156);
nor U6072 (N_6072,N_2801,N_2830);
nand U6073 (N_6073,N_4733,N_4971);
or U6074 (N_6074,N_3469,N_4899);
or U6075 (N_6075,N_2960,N_4639);
nand U6076 (N_6076,N_2828,N_4664);
xnor U6077 (N_6077,N_4797,N_4200);
and U6078 (N_6078,N_2835,N_3201);
nor U6079 (N_6079,N_3004,N_2726);
nor U6080 (N_6080,N_4308,N_4437);
nor U6081 (N_6081,N_3532,N_3113);
and U6082 (N_6082,N_2693,N_3873);
and U6083 (N_6083,N_3819,N_3951);
nand U6084 (N_6084,N_4032,N_3821);
nor U6085 (N_6085,N_3814,N_4992);
or U6086 (N_6086,N_4410,N_4780);
nor U6087 (N_6087,N_3879,N_2539);
xor U6088 (N_6088,N_3419,N_2590);
nor U6089 (N_6089,N_3058,N_2968);
xnor U6090 (N_6090,N_3190,N_3953);
xor U6091 (N_6091,N_4385,N_3929);
and U6092 (N_6092,N_4986,N_3731);
nand U6093 (N_6093,N_3944,N_3755);
nor U6094 (N_6094,N_4496,N_4121);
nand U6095 (N_6095,N_4923,N_2935);
or U6096 (N_6096,N_3433,N_4768);
or U6097 (N_6097,N_3826,N_2873);
nand U6098 (N_6098,N_3983,N_4577);
nor U6099 (N_6099,N_3803,N_4567);
xor U6100 (N_6100,N_4634,N_2997);
nor U6101 (N_6101,N_2788,N_4699);
nand U6102 (N_6102,N_3151,N_2922);
nand U6103 (N_6103,N_2595,N_4197);
or U6104 (N_6104,N_4164,N_4690);
and U6105 (N_6105,N_3327,N_4296);
xor U6106 (N_6106,N_3512,N_3752);
nand U6107 (N_6107,N_4444,N_4476);
xnor U6108 (N_6108,N_4360,N_2502);
xor U6109 (N_6109,N_4555,N_3799);
xor U6110 (N_6110,N_4319,N_3610);
xor U6111 (N_6111,N_2941,N_4568);
nand U6112 (N_6112,N_3479,N_4486);
nand U6113 (N_6113,N_3704,N_4341);
and U6114 (N_6114,N_3920,N_3810);
or U6115 (N_6115,N_4536,N_2811);
nand U6116 (N_6116,N_4488,N_3852);
nand U6117 (N_6117,N_4340,N_3282);
nand U6118 (N_6118,N_4261,N_2965);
and U6119 (N_6119,N_2850,N_2844);
and U6120 (N_6120,N_4905,N_3486);
nand U6121 (N_6121,N_3188,N_3575);
nor U6122 (N_6122,N_2695,N_3389);
or U6123 (N_6123,N_2656,N_3554);
xnor U6124 (N_6124,N_4255,N_2548);
nand U6125 (N_6125,N_2543,N_4356);
xnor U6126 (N_6126,N_4896,N_4252);
nand U6127 (N_6127,N_2729,N_2723);
or U6128 (N_6128,N_4247,N_2536);
nor U6129 (N_6129,N_2784,N_2544);
and U6130 (N_6130,N_3340,N_3715);
xnor U6131 (N_6131,N_4169,N_3365);
or U6132 (N_6132,N_2888,N_2733);
xor U6133 (N_6133,N_2862,N_4891);
and U6134 (N_6134,N_2667,N_4098);
nand U6135 (N_6135,N_2772,N_3175);
xor U6136 (N_6136,N_4433,N_4087);
xnor U6137 (N_6137,N_2754,N_3062);
and U6138 (N_6138,N_4997,N_3024);
and U6139 (N_6139,N_4138,N_4777);
xor U6140 (N_6140,N_3743,N_4994);
xnor U6141 (N_6141,N_3490,N_3369);
or U6142 (N_6142,N_3112,N_4458);
or U6143 (N_6143,N_2659,N_4624);
nand U6144 (N_6144,N_4995,N_3817);
xnor U6145 (N_6145,N_3441,N_3492);
nor U6146 (N_6146,N_2832,N_4900);
nand U6147 (N_6147,N_4569,N_3430);
nand U6148 (N_6148,N_3079,N_3968);
and U6149 (N_6149,N_4232,N_4165);
nor U6150 (N_6150,N_4233,N_2742);
xnor U6151 (N_6151,N_3034,N_4182);
nor U6152 (N_6152,N_3759,N_2853);
and U6153 (N_6153,N_3181,N_3354);
xnor U6154 (N_6154,N_4866,N_4346);
and U6155 (N_6155,N_3696,N_3583);
xnor U6156 (N_6156,N_4885,N_4782);
nand U6157 (N_6157,N_2953,N_3402);
or U6158 (N_6158,N_3060,N_4125);
or U6159 (N_6159,N_4552,N_3368);
nor U6160 (N_6160,N_2537,N_3897);
or U6161 (N_6161,N_2731,N_2713);
nand U6162 (N_6162,N_2635,N_4085);
or U6163 (N_6163,N_3767,N_4452);
nor U6164 (N_6164,N_2699,N_3990);
and U6165 (N_6165,N_3895,N_2511);
and U6166 (N_6166,N_4317,N_4709);
xor U6167 (N_6167,N_3607,N_3925);
nor U6168 (N_6168,N_4434,N_3594);
and U6169 (N_6169,N_3945,N_2999);
nand U6170 (N_6170,N_4173,N_3325);
nor U6171 (N_6171,N_4303,N_3995);
and U6172 (N_6172,N_4416,N_3812);
and U6173 (N_6173,N_4933,N_4417);
nand U6174 (N_6174,N_2795,N_3007);
nor U6175 (N_6175,N_4035,N_4556);
nand U6176 (N_6176,N_2872,N_3838);
xnor U6177 (N_6177,N_2594,N_4378);
nor U6178 (N_6178,N_3761,N_3332);
xor U6179 (N_6179,N_3881,N_2981);
and U6180 (N_6180,N_4229,N_4368);
xnor U6181 (N_6181,N_4119,N_2762);
and U6182 (N_6182,N_3011,N_3602);
and U6183 (N_6183,N_3771,N_4917);
nor U6184 (N_6184,N_4388,N_4886);
or U6185 (N_6185,N_3915,N_4167);
nand U6186 (N_6186,N_3621,N_4477);
xor U6187 (N_6187,N_2974,N_3927);
and U6188 (N_6188,N_3382,N_2573);
and U6189 (N_6189,N_4967,N_4778);
and U6190 (N_6190,N_3296,N_3758);
or U6191 (N_6191,N_2550,N_3534);
nand U6192 (N_6192,N_2510,N_2857);
xor U6193 (N_6193,N_2803,N_4215);
xnor U6194 (N_6194,N_2621,N_2955);
or U6195 (N_6195,N_3032,N_2745);
xor U6196 (N_6196,N_3551,N_2895);
and U6197 (N_6197,N_4857,N_3405);
and U6198 (N_6198,N_2952,N_2636);
nor U6199 (N_6199,N_4081,N_4166);
xor U6200 (N_6200,N_4210,N_3592);
xor U6201 (N_6201,N_4342,N_2508);
nor U6202 (N_6202,N_2680,N_4572);
nor U6203 (N_6203,N_3169,N_3245);
nand U6204 (N_6204,N_3954,N_3216);
xor U6205 (N_6205,N_4963,N_3640);
nand U6206 (N_6206,N_3887,N_2697);
xnor U6207 (N_6207,N_4390,N_3471);
nor U6208 (N_6208,N_4144,N_2582);
nor U6209 (N_6209,N_4815,N_3130);
nand U6210 (N_6210,N_3185,N_3674);
xor U6211 (N_6211,N_2705,N_3048);
nand U6212 (N_6212,N_2969,N_4601);
nor U6213 (N_6213,N_3343,N_2770);
xor U6214 (N_6214,N_2979,N_3654);
xnor U6215 (N_6215,N_4538,N_4400);
and U6216 (N_6216,N_3792,N_2542);
and U6217 (N_6217,N_4212,N_4315);
nor U6218 (N_6218,N_3126,N_3984);
and U6219 (N_6219,N_4078,N_3733);
or U6220 (N_6220,N_3375,N_2903);
nand U6221 (N_6221,N_3294,N_4380);
nor U6222 (N_6222,N_3379,N_2833);
nor U6223 (N_6223,N_4666,N_4839);
nand U6224 (N_6224,N_3710,N_3304);
or U6225 (N_6225,N_3495,N_3411);
and U6226 (N_6226,N_3429,N_4482);
nor U6227 (N_6227,N_4953,N_3115);
nand U6228 (N_6228,N_4320,N_2591);
nor U6229 (N_6229,N_3779,N_3002);
xor U6230 (N_6230,N_4902,N_3923);
and U6231 (N_6231,N_3893,N_4284);
nor U6232 (N_6232,N_3749,N_4769);
nor U6233 (N_6233,N_3791,N_3922);
or U6234 (N_6234,N_4481,N_3134);
and U6235 (N_6235,N_4234,N_4864);
and U6236 (N_6236,N_4454,N_3148);
or U6237 (N_6237,N_3051,N_3085);
nand U6238 (N_6238,N_3705,N_3782);
nor U6239 (N_6239,N_4491,N_3824);
or U6240 (N_6240,N_3461,N_3250);
nand U6241 (N_6241,N_3041,N_4456);
xnor U6242 (N_6242,N_3456,N_4475);
xnor U6243 (N_6243,N_4887,N_3899);
nor U6244 (N_6244,N_2554,N_2807);
nand U6245 (N_6245,N_3198,N_3451);
xnor U6246 (N_6246,N_3796,N_2513);
nand U6247 (N_6247,N_3240,N_4593);
xor U6248 (N_6248,N_3209,N_3462);
or U6249 (N_6249,N_4523,N_3614);
xnor U6250 (N_6250,N_2852,N_3418);
xor U6251 (N_6251,N_4972,N_3602);
nor U6252 (N_6252,N_4336,N_3905);
or U6253 (N_6253,N_3201,N_2829);
xor U6254 (N_6254,N_4823,N_3098);
nor U6255 (N_6255,N_4417,N_4446);
and U6256 (N_6256,N_4378,N_4407);
nor U6257 (N_6257,N_4800,N_3044);
nor U6258 (N_6258,N_4819,N_3561);
or U6259 (N_6259,N_3946,N_2572);
and U6260 (N_6260,N_4549,N_4604);
or U6261 (N_6261,N_4170,N_4851);
xor U6262 (N_6262,N_4447,N_3886);
xnor U6263 (N_6263,N_3654,N_4880);
xor U6264 (N_6264,N_4444,N_3982);
xnor U6265 (N_6265,N_3382,N_4806);
nor U6266 (N_6266,N_3423,N_2896);
nor U6267 (N_6267,N_4906,N_3393);
xor U6268 (N_6268,N_4629,N_4911);
xor U6269 (N_6269,N_2558,N_3788);
and U6270 (N_6270,N_4786,N_3297);
nor U6271 (N_6271,N_3901,N_2841);
and U6272 (N_6272,N_3809,N_4622);
nor U6273 (N_6273,N_3505,N_2625);
nand U6274 (N_6274,N_4646,N_2733);
or U6275 (N_6275,N_4436,N_4963);
and U6276 (N_6276,N_4982,N_4703);
nor U6277 (N_6277,N_3872,N_4880);
nor U6278 (N_6278,N_4406,N_3374);
or U6279 (N_6279,N_4867,N_3521);
nor U6280 (N_6280,N_4137,N_3717);
and U6281 (N_6281,N_4898,N_4110);
and U6282 (N_6282,N_3072,N_4936);
nand U6283 (N_6283,N_2562,N_4548);
nor U6284 (N_6284,N_2590,N_4038);
nor U6285 (N_6285,N_3240,N_4796);
nand U6286 (N_6286,N_3441,N_4330);
or U6287 (N_6287,N_4788,N_4713);
nand U6288 (N_6288,N_3335,N_3638);
nand U6289 (N_6289,N_2543,N_4778);
xnor U6290 (N_6290,N_3437,N_4841);
nand U6291 (N_6291,N_3975,N_3992);
nand U6292 (N_6292,N_3544,N_3892);
and U6293 (N_6293,N_4036,N_2757);
nand U6294 (N_6294,N_3112,N_4477);
and U6295 (N_6295,N_3860,N_3139);
and U6296 (N_6296,N_4490,N_3877);
xnor U6297 (N_6297,N_2993,N_3363);
and U6298 (N_6298,N_4309,N_2755);
xor U6299 (N_6299,N_3367,N_3366);
xor U6300 (N_6300,N_3850,N_3871);
or U6301 (N_6301,N_4866,N_4607);
or U6302 (N_6302,N_4696,N_3528);
xor U6303 (N_6303,N_4155,N_3962);
and U6304 (N_6304,N_4419,N_2658);
nor U6305 (N_6305,N_3415,N_3035);
nor U6306 (N_6306,N_4955,N_3843);
or U6307 (N_6307,N_4834,N_4672);
or U6308 (N_6308,N_3690,N_3418);
nand U6309 (N_6309,N_4619,N_2731);
xor U6310 (N_6310,N_3483,N_3742);
nor U6311 (N_6311,N_4209,N_3679);
xnor U6312 (N_6312,N_3586,N_3611);
nor U6313 (N_6313,N_2816,N_3526);
or U6314 (N_6314,N_2993,N_4039);
and U6315 (N_6315,N_3334,N_4587);
or U6316 (N_6316,N_3223,N_3107);
or U6317 (N_6317,N_2635,N_3530);
nand U6318 (N_6318,N_4032,N_3214);
xor U6319 (N_6319,N_4719,N_2544);
and U6320 (N_6320,N_4436,N_3347);
nand U6321 (N_6321,N_3681,N_4769);
nand U6322 (N_6322,N_2787,N_3053);
nor U6323 (N_6323,N_4837,N_4666);
or U6324 (N_6324,N_2824,N_2958);
nor U6325 (N_6325,N_2965,N_4687);
nor U6326 (N_6326,N_4324,N_2781);
nand U6327 (N_6327,N_4871,N_2557);
or U6328 (N_6328,N_2960,N_3828);
and U6329 (N_6329,N_3095,N_4088);
nor U6330 (N_6330,N_3845,N_3294);
nand U6331 (N_6331,N_3574,N_4304);
or U6332 (N_6332,N_4035,N_3277);
xor U6333 (N_6333,N_4526,N_4806);
or U6334 (N_6334,N_3122,N_4483);
and U6335 (N_6335,N_4024,N_3174);
nor U6336 (N_6336,N_3886,N_4314);
nor U6337 (N_6337,N_3877,N_4655);
nand U6338 (N_6338,N_2807,N_2751);
or U6339 (N_6339,N_3822,N_3574);
and U6340 (N_6340,N_2734,N_4848);
and U6341 (N_6341,N_3988,N_3864);
nor U6342 (N_6342,N_2757,N_4024);
or U6343 (N_6343,N_4409,N_4046);
or U6344 (N_6344,N_2531,N_4660);
xnor U6345 (N_6345,N_2555,N_3922);
nor U6346 (N_6346,N_3982,N_3360);
or U6347 (N_6347,N_3673,N_3978);
and U6348 (N_6348,N_4112,N_3978);
nand U6349 (N_6349,N_3490,N_3738);
and U6350 (N_6350,N_3683,N_2895);
and U6351 (N_6351,N_4696,N_2884);
xor U6352 (N_6352,N_4023,N_3889);
xnor U6353 (N_6353,N_3254,N_3659);
or U6354 (N_6354,N_4454,N_3425);
or U6355 (N_6355,N_4032,N_3631);
xor U6356 (N_6356,N_2546,N_4462);
nor U6357 (N_6357,N_3754,N_4099);
nor U6358 (N_6358,N_2586,N_2986);
and U6359 (N_6359,N_4384,N_4403);
nor U6360 (N_6360,N_4766,N_3654);
nand U6361 (N_6361,N_4732,N_3998);
nor U6362 (N_6362,N_2614,N_4898);
nand U6363 (N_6363,N_2750,N_3727);
and U6364 (N_6364,N_3254,N_3692);
and U6365 (N_6365,N_3635,N_2655);
or U6366 (N_6366,N_3336,N_2824);
xor U6367 (N_6367,N_4374,N_4470);
or U6368 (N_6368,N_2871,N_4545);
and U6369 (N_6369,N_3802,N_4057);
or U6370 (N_6370,N_4958,N_4111);
nand U6371 (N_6371,N_3479,N_2692);
and U6372 (N_6372,N_2966,N_4286);
nor U6373 (N_6373,N_4458,N_4205);
or U6374 (N_6374,N_4499,N_3536);
nand U6375 (N_6375,N_3610,N_3041);
or U6376 (N_6376,N_4689,N_4356);
or U6377 (N_6377,N_4578,N_2911);
and U6378 (N_6378,N_4421,N_4272);
or U6379 (N_6379,N_4916,N_3455);
and U6380 (N_6380,N_4688,N_4288);
xnor U6381 (N_6381,N_3337,N_4458);
nor U6382 (N_6382,N_2640,N_2999);
or U6383 (N_6383,N_4088,N_4903);
xnor U6384 (N_6384,N_4251,N_3851);
nand U6385 (N_6385,N_4542,N_3453);
or U6386 (N_6386,N_4100,N_3665);
or U6387 (N_6387,N_4080,N_4930);
or U6388 (N_6388,N_2501,N_4320);
nor U6389 (N_6389,N_3177,N_4263);
xor U6390 (N_6390,N_4210,N_3499);
and U6391 (N_6391,N_3285,N_2798);
and U6392 (N_6392,N_4074,N_2572);
xor U6393 (N_6393,N_3961,N_2646);
nor U6394 (N_6394,N_3015,N_2670);
nor U6395 (N_6395,N_3317,N_3835);
nor U6396 (N_6396,N_3819,N_3468);
xnor U6397 (N_6397,N_3458,N_3340);
or U6398 (N_6398,N_3356,N_4176);
xor U6399 (N_6399,N_2663,N_2835);
xnor U6400 (N_6400,N_2566,N_3829);
xnor U6401 (N_6401,N_4746,N_4523);
and U6402 (N_6402,N_3672,N_4770);
nor U6403 (N_6403,N_3458,N_2515);
nor U6404 (N_6404,N_2544,N_3539);
or U6405 (N_6405,N_3381,N_4842);
nor U6406 (N_6406,N_4471,N_3440);
or U6407 (N_6407,N_4949,N_2775);
and U6408 (N_6408,N_4443,N_4868);
nor U6409 (N_6409,N_4116,N_4770);
and U6410 (N_6410,N_4996,N_3556);
nor U6411 (N_6411,N_2897,N_3350);
or U6412 (N_6412,N_4268,N_3807);
xnor U6413 (N_6413,N_3813,N_2929);
and U6414 (N_6414,N_3416,N_4373);
or U6415 (N_6415,N_3622,N_4165);
xnor U6416 (N_6416,N_4053,N_2893);
xnor U6417 (N_6417,N_4724,N_4361);
xnor U6418 (N_6418,N_3227,N_4252);
nor U6419 (N_6419,N_2905,N_2763);
and U6420 (N_6420,N_3235,N_3752);
and U6421 (N_6421,N_2640,N_3956);
nand U6422 (N_6422,N_2830,N_3734);
nand U6423 (N_6423,N_2892,N_3681);
xnor U6424 (N_6424,N_4004,N_2799);
nor U6425 (N_6425,N_3426,N_2783);
or U6426 (N_6426,N_3369,N_4550);
xnor U6427 (N_6427,N_4313,N_4614);
xor U6428 (N_6428,N_3274,N_2937);
nor U6429 (N_6429,N_3983,N_4992);
or U6430 (N_6430,N_2881,N_3632);
and U6431 (N_6431,N_4246,N_4904);
or U6432 (N_6432,N_3235,N_3252);
or U6433 (N_6433,N_2746,N_4163);
and U6434 (N_6434,N_3948,N_4927);
nor U6435 (N_6435,N_3162,N_3829);
nor U6436 (N_6436,N_4951,N_4420);
nor U6437 (N_6437,N_4643,N_2656);
nor U6438 (N_6438,N_2667,N_3491);
nor U6439 (N_6439,N_3013,N_3791);
and U6440 (N_6440,N_3083,N_3277);
nand U6441 (N_6441,N_3718,N_3347);
nand U6442 (N_6442,N_2576,N_4743);
and U6443 (N_6443,N_2602,N_2726);
nand U6444 (N_6444,N_4168,N_3358);
or U6445 (N_6445,N_4189,N_3666);
nand U6446 (N_6446,N_3455,N_3260);
xor U6447 (N_6447,N_4221,N_2692);
or U6448 (N_6448,N_3730,N_3315);
xnor U6449 (N_6449,N_4104,N_3637);
nand U6450 (N_6450,N_4745,N_4616);
nand U6451 (N_6451,N_4407,N_3102);
and U6452 (N_6452,N_4193,N_3118);
xnor U6453 (N_6453,N_3863,N_4807);
and U6454 (N_6454,N_3393,N_4324);
or U6455 (N_6455,N_4136,N_4826);
xnor U6456 (N_6456,N_4261,N_4228);
or U6457 (N_6457,N_3317,N_4126);
and U6458 (N_6458,N_4727,N_3353);
or U6459 (N_6459,N_2875,N_4668);
and U6460 (N_6460,N_2733,N_3767);
nor U6461 (N_6461,N_3309,N_3786);
nor U6462 (N_6462,N_3764,N_2894);
xnor U6463 (N_6463,N_3937,N_4024);
or U6464 (N_6464,N_3406,N_2854);
and U6465 (N_6465,N_4612,N_4588);
nor U6466 (N_6466,N_4755,N_4628);
nand U6467 (N_6467,N_3383,N_3718);
or U6468 (N_6468,N_3284,N_3268);
nor U6469 (N_6469,N_2577,N_4941);
xnor U6470 (N_6470,N_3600,N_4192);
and U6471 (N_6471,N_3600,N_4737);
xor U6472 (N_6472,N_4387,N_3582);
or U6473 (N_6473,N_4920,N_2649);
nor U6474 (N_6474,N_2794,N_3921);
or U6475 (N_6475,N_4793,N_4267);
nand U6476 (N_6476,N_4100,N_3424);
nor U6477 (N_6477,N_4976,N_2579);
nor U6478 (N_6478,N_2526,N_4276);
xnor U6479 (N_6479,N_3794,N_4200);
nand U6480 (N_6480,N_2859,N_3000);
nor U6481 (N_6481,N_3657,N_4880);
and U6482 (N_6482,N_4246,N_2735);
xnor U6483 (N_6483,N_4210,N_2814);
nor U6484 (N_6484,N_3294,N_4663);
or U6485 (N_6485,N_3527,N_4634);
or U6486 (N_6486,N_4363,N_4707);
nor U6487 (N_6487,N_4750,N_4349);
and U6488 (N_6488,N_4151,N_4884);
nor U6489 (N_6489,N_2570,N_2948);
nor U6490 (N_6490,N_2970,N_4605);
nor U6491 (N_6491,N_4142,N_3866);
or U6492 (N_6492,N_2832,N_2615);
or U6493 (N_6493,N_4123,N_2723);
and U6494 (N_6494,N_4973,N_4170);
or U6495 (N_6495,N_4097,N_4384);
nand U6496 (N_6496,N_2615,N_4226);
nor U6497 (N_6497,N_4428,N_3932);
or U6498 (N_6498,N_3344,N_3173);
nand U6499 (N_6499,N_4649,N_2839);
nand U6500 (N_6500,N_4760,N_4873);
nor U6501 (N_6501,N_4080,N_4355);
nand U6502 (N_6502,N_3687,N_4289);
nor U6503 (N_6503,N_3780,N_2682);
xnor U6504 (N_6504,N_4685,N_3440);
xor U6505 (N_6505,N_2773,N_4585);
xnor U6506 (N_6506,N_3941,N_3537);
xor U6507 (N_6507,N_3206,N_4062);
xor U6508 (N_6508,N_3989,N_4078);
or U6509 (N_6509,N_2605,N_4498);
nand U6510 (N_6510,N_3212,N_4196);
nor U6511 (N_6511,N_4386,N_3217);
and U6512 (N_6512,N_2923,N_3344);
nor U6513 (N_6513,N_4156,N_4733);
xor U6514 (N_6514,N_3095,N_2582);
xnor U6515 (N_6515,N_3418,N_4059);
xnor U6516 (N_6516,N_3445,N_2666);
and U6517 (N_6517,N_4358,N_4585);
nand U6518 (N_6518,N_2753,N_4500);
nor U6519 (N_6519,N_4078,N_3797);
nor U6520 (N_6520,N_4593,N_4620);
nand U6521 (N_6521,N_4003,N_3520);
nand U6522 (N_6522,N_3974,N_3473);
or U6523 (N_6523,N_4471,N_3653);
nand U6524 (N_6524,N_4356,N_3333);
or U6525 (N_6525,N_3469,N_2951);
nand U6526 (N_6526,N_4398,N_2721);
or U6527 (N_6527,N_2593,N_4817);
xnor U6528 (N_6528,N_4839,N_2600);
nand U6529 (N_6529,N_3530,N_4643);
nor U6530 (N_6530,N_4054,N_3473);
and U6531 (N_6531,N_3806,N_3529);
or U6532 (N_6532,N_3333,N_4121);
nand U6533 (N_6533,N_3746,N_4834);
xnor U6534 (N_6534,N_4309,N_2996);
and U6535 (N_6535,N_4098,N_3857);
and U6536 (N_6536,N_4202,N_4205);
or U6537 (N_6537,N_4387,N_4746);
nor U6538 (N_6538,N_3625,N_2975);
nor U6539 (N_6539,N_3121,N_2933);
xnor U6540 (N_6540,N_3472,N_3724);
and U6541 (N_6541,N_4498,N_4819);
and U6542 (N_6542,N_3698,N_2578);
nand U6543 (N_6543,N_4758,N_4464);
nor U6544 (N_6544,N_4327,N_2856);
xor U6545 (N_6545,N_3425,N_4240);
or U6546 (N_6546,N_4626,N_3247);
or U6547 (N_6547,N_2637,N_4669);
or U6548 (N_6548,N_2632,N_4853);
or U6549 (N_6549,N_3534,N_3695);
and U6550 (N_6550,N_3798,N_4820);
xnor U6551 (N_6551,N_2886,N_4961);
nand U6552 (N_6552,N_4184,N_3246);
xnor U6553 (N_6553,N_3094,N_3519);
or U6554 (N_6554,N_3622,N_3950);
nor U6555 (N_6555,N_3606,N_2929);
or U6556 (N_6556,N_3798,N_2973);
nand U6557 (N_6557,N_2715,N_3465);
nor U6558 (N_6558,N_4510,N_4378);
xnor U6559 (N_6559,N_3427,N_3704);
xnor U6560 (N_6560,N_4352,N_3415);
xnor U6561 (N_6561,N_4523,N_4430);
nand U6562 (N_6562,N_4352,N_2755);
nand U6563 (N_6563,N_4287,N_4910);
or U6564 (N_6564,N_4997,N_4669);
xor U6565 (N_6565,N_3166,N_3076);
nor U6566 (N_6566,N_4721,N_3854);
xnor U6567 (N_6567,N_3210,N_3633);
nand U6568 (N_6568,N_4680,N_2909);
nor U6569 (N_6569,N_4894,N_4598);
or U6570 (N_6570,N_3210,N_3115);
and U6571 (N_6571,N_2767,N_3502);
or U6572 (N_6572,N_3725,N_2741);
or U6573 (N_6573,N_3610,N_4076);
nand U6574 (N_6574,N_3179,N_3981);
and U6575 (N_6575,N_4794,N_2753);
xor U6576 (N_6576,N_3426,N_4371);
nor U6577 (N_6577,N_4758,N_4718);
xor U6578 (N_6578,N_4398,N_4113);
and U6579 (N_6579,N_4411,N_4247);
nand U6580 (N_6580,N_4582,N_2759);
or U6581 (N_6581,N_3016,N_2525);
or U6582 (N_6582,N_3420,N_4665);
nand U6583 (N_6583,N_3287,N_4925);
nand U6584 (N_6584,N_4421,N_3951);
xor U6585 (N_6585,N_4127,N_4491);
and U6586 (N_6586,N_4156,N_3113);
nand U6587 (N_6587,N_3306,N_3789);
nand U6588 (N_6588,N_4071,N_2858);
or U6589 (N_6589,N_3701,N_3353);
nand U6590 (N_6590,N_4680,N_2607);
or U6591 (N_6591,N_3817,N_3081);
nand U6592 (N_6592,N_2974,N_3025);
or U6593 (N_6593,N_3055,N_4395);
and U6594 (N_6594,N_3527,N_4691);
and U6595 (N_6595,N_4552,N_3500);
or U6596 (N_6596,N_2761,N_3000);
and U6597 (N_6597,N_3058,N_4185);
nand U6598 (N_6598,N_3659,N_3237);
and U6599 (N_6599,N_2768,N_4443);
nand U6600 (N_6600,N_3148,N_4923);
nor U6601 (N_6601,N_3256,N_2773);
xnor U6602 (N_6602,N_4813,N_2527);
xor U6603 (N_6603,N_2586,N_4413);
nor U6604 (N_6604,N_2652,N_3153);
xor U6605 (N_6605,N_3417,N_3398);
xnor U6606 (N_6606,N_3285,N_4428);
xnor U6607 (N_6607,N_3220,N_3057);
xor U6608 (N_6608,N_4447,N_2975);
or U6609 (N_6609,N_4616,N_4017);
nor U6610 (N_6610,N_4533,N_4018);
and U6611 (N_6611,N_4626,N_4765);
nand U6612 (N_6612,N_3126,N_3084);
nand U6613 (N_6613,N_3899,N_4722);
and U6614 (N_6614,N_4036,N_4074);
nand U6615 (N_6615,N_3886,N_2837);
or U6616 (N_6616,N_3390,N_4528);
or U6617 (N_6617,N_3541,N_3176);
nand U6618 (N_6618,N_2705,N_3368);
or U6619 (N_6619,N_3364,N_4037);
and U6620 (N_6620,N_4841,N_3092);
or U6621 (N_6621,N_4069,N_2586);
nand U6622 (N_6622,N_4342,N_3265);
nor U6623 (N_6623,N_2599,N_2669);
nor U6624 (N_6624,N_3271,N_3616);
nand U6625 (N_6625,N_3372,N_3102);
nand U6626 (N_6626,N_3301,N_3576);
nand U6627 (N_6627,N_2558,N_3347);
and U6628 (N_6628,N_4425,N_3479);
and U6629 (N_6629,N_4610,N_2897);
nor U6630 (N_6630,N_2884,N_4449);
nor U6631 (N_6631,N_3200,N_2965);
nand U6632 (N_6632,N_4181,N_4533);
and U6633 (N_6633,N_2634,N_4965);
and U6634 (N_6634,N_4090,N_2551);
or U6635 (N_6635,N_2543,N_2888);
nor U6636 (N_6636,N_4233,N_3205);
nand U6637 (N_6637,N_4747,N_3287);
nand U6638 (N_6638,N_2620,N_3389);
nor U6639 (N_6639,N_4532,N_4982);
xor U6640 (N_6640,N_4748,N_2931);
nand U6641 (N_6641,N_3853,N_4775);
or U6642 (N_6642,N_4661,N_3928);
or U6643 (N_6643,N_4112,N_3251);
xnor U6644 (N_6644,N_3554,N_4174);
xor U6645 (N_6645,N_4949,N_4322);
nand U6646 (N_6646,N_3321,N_2979);
nor U6647 (N_6647,N_3311,N_4703);
xor U6648 (N_6648,N_2828,N_2974);
and U6649 (N_6649,N_3416,N_4456);
nor U6650 (N_6650,N_4630,N_2674);
xnor U6651 (N_6651,N_4103,N_4483);
nor U6652 (N_6652,N_4465,N_2910);
and U6653 (N_6653,N_3373,N_2754);
and U6654 (N_6654,N_3349,N_4663);
nor U6655 (N_6655,N_4741,N_2708);
nor U6656 (N_6656,N_4166,N_4311);
nand U6657 (N_6657,N_3323,N_3941);
or U6658 (N_6658,N_4672,N_4621);
xnor U6659 (N_6659,N_4947,N_2543);
nand U6660 (N_6660,N_4468,N_4224);
nand U6661 (N_6661,N_2650,N_4489);
nor U6662 (N_6662,N_3805,N_3321);
xnor U6663 (N_6663,N_4513,N_3941);
nand U6664 (N_6664,N_2888,N_4031);
nand U6665 (N_6665,N_2635,N_4044);
nor U6666 (N_6666,N_3590,N_3626);
or U6667 (N_6667,N_2623,N_4218);
nand U6668 (N_6668,N_3259,N_4076);
or U6669 (N_6669,N_4075,N_2902);
nor U6670 (N_6670,N_3593,N_3489);
or U6671 (N_6671,N_3447,N_4650);
xor U6672 (N_6672,N_3264,N_3784);
or U6673 (N_6673,N_2966,N_4806);
or U6674 (N_6674,N_2935,N_2554);
nand U6675 (N_6675,N_3449,N_3600);
or U6676 (N_6676,N_2601,N_3094);
and U6677 (N_6677,N_3166,N_3775);
or U6678 (N_6678,N_2524,N_4947);
nor U6679 (N_6679,N_3906,N_3378);
and U6680 (N_6680,N_2927,N_4775);
nor U6681 (N_6681,N_4908,N_4219);
and U6682 (N_6682,N_4931,N_4484);
or U6683 (N_6683,N_3522,N_3795);
nor U6684 (N_6684,N_3582,N_3517);
xnor U6685 (N_6685,N_3364,N_4997);
and U6686 (N_6686,N_3114,N_3428);
or U6687 (N_6687,N_4776,N_3919);
nand U6688 (N_6688,N_4854,N_3732);
or U6689 (N_6689,N_4197,N_3925);
and U6690 (N_6690,N_3852,N_2565);
and U6691 (N_6691,N_4138,N_4210);
nand U6692 (N_6692,N_3013,N_2980);
nand U6693 (N_6693,N_4603,N_3075);
and U6694 (N_6694,N_2877,N_4371);
nor U6695 (N_6695,N_4539,N_2679);
and U6696 (N_6696,N_3166,N_3279);
xnor U6697 (N_6697,N_4647,N_3200);
nand U6698 (N_6698,N_3780,N_4552);
nor U6699 (N_6699,N_3645,N_3431);
or U6700 (N_6700,N_4704,N_4798);
and U6701 (N_6701,N_4145,N_2871);
and U6702 (N_6702,N_3050,N_4740);
nand U6703 (N_6703,N_3726,N_3247);
xor U6704 (N_6704,N_4931,N_4158);
nor U6705 (N_6705,N_4760,N_3754);
nand U6706 (N_6706,N_2568,N_3129);
xor U6707 (N_6707,N_3845,N_4132);
xor U6708 (N_6708,N_4225,N_3564);
or U6709 (N_6709,N_3073,N_3725);
and U6710 (N_6710,N_2652,N_2708);
or U6711 (N_6711,N_4271,N_3622);
nor U6712 (N_6712,N_3855,N_3340);
or U6713 (N_6713,N_2654,N_4490);
or U6714 (N_6714,N_4264,N_2954);
nor U6715 (N_6715,N_4255,N_3016);
nor U6716 (N_6716,N_3084,N_2832);
xor U6717 (N_6717,N_3800,N_3261);
or U6718 (N_6718,N_3966,N_3050);
and U6719 (N_6719,N_2749,N_3856);
xor U6720 (N_6720,N_3139,N_4617);
nand U6721 (N_6721,N_3388,N_2987);
and U6722 (N_6722,N_3792,N_2563);
nor U6723 (N_6723,N_4970,N_3708);
xor U6724 (N_6724,N_4743,N_4235);
nor U6725 (N_6725,N_2651,N_4680);
or U6726 (N_6726,N_4048,N_4064);
and U6727 (N_6727,N_3771,N_4501);
nor U6728 (N_6728,N_3620,N_3997);
nor U6729 (N_6729,N_3838,N_3090);
and U6730 (N_6730,N_4595,N_3039);
nor U6731 (N_6731,N_4996,N_3282);
nor U6732 (N_6732,N_4006,N_2737);
nor U6733 (N_6733,N_3440,N_3518);
nor U6734 (N_6734,N_4756,N_4651);
nor U6735 (N_6735,N_3850,N_3906);
or U6736 (N_6736,N_3182,N_2660);
xnor U6737 (N_6737,N_3749,N_4382);
nand U6738 (N_6738,N_3471,N_4952);
nand U6739 (N_6739,N_3621,N_3646);
xnor U6740 (N_6740,N_4433,N_2791);
nand U6741 (N_6741,N_3667,N_2957);
or U6742 (N_6742,N_3249,N_4275);
nand U6743 (N_6743,N_4500,N_3138);
or U6744 (N_6744,N_3199,N_3826);
xnor U6745 (N_6745,N_2874,N_3097);
nor U6746 (N_6746,N_3273,N_2543);
xnor U6747 (N_6747,N_2954,N_3503);
nand U6748 (N_6748,N_2803,N_2918);
nand U6749 (N_6749,N_4213,N_4732);
nor U6750 (N_6750,N_3617,N_3889);
nor U6751 (N_6751,N_3375,N_4997);
and U6752 (N_6752,N_3239,N_4922);
nor U6753 (N_6753,N_4344,N_2983);
nand U6754 (N_6754,N_3357,N_3059);
nand U6755 (N_6755,N_2772,N_4269);
xor U6756 (N_6756,N_4599,N_4862);
nor U6757 (N_6757,N_3884,N_3422);
nor U6758 (N_6758,N_2610,N_4782);
nand U6759 (N_6759,N_3139,N_3593);
xnor U6760 (N_6760,N_2501,N_4829);
nand U6761 (N_6761,N_4441,N_2862);
nand U6762 (N_6762,N_3768,N_3598);
or U6763 (N_6763,N_4895,N_3436);
nor U6764 (N_6764,N_2556,N_3313);
xnor U6765 (N_6765,N_3403,N_2771);
or U6766 (N_6766,N_3147,N_3671);
and U6767 (N_6767,N_3551,N_2805);
or U6768 (N_6768,N_4366,N_4206);
xnor U6769 (N_6769,N_4028,N_3648);
nand U6770 (N_6770,N_2879,N_4414);
and U6771 (N_6771,N_4087,N_3467);
xor U6772 (N_6772,N_3382,N_4094);
xor U6773 (N_6773,N_4994,N_2688);
nor U6774 (N_6774,N_3274,N_4932);
nor U6775 (N_6775,N_4425,N_3027);
nand U6776 (N_6776,N_2822,N_3742);
nand U6777 (N_6777,N_4706,N_2822);
and U6778 (N_6778,N_3062,N_4848);
xor U6779 (N_6779,N_3339,N_3824);
nand U6780 (N_6780,N_4674,N_3285);
and U6781 (N_6781,N_4640,N_3391);
or U6782 (N_6782,N_2576,N_4297);
nand U6783 (N_6783,N_4274,N_3620);
and U6784 (N_6784,N_4019,N_3493);
and U6785 (N_6785,N_4373,N_3202);
or U6786 (N_6786,N_3787,N_2916);
and U6787 (N_6787,N_3096,N_4638);
nor U6788 (N_6788,N_3446,N_3217);
xor U6789 (N_6789,N_2692,N_2628);
and U6790 (N_6790,N_4691,N_3504);
or U6791 (N_6791,N_4992,N_2797);
and U6792 (N_6792,N_4652,N_3059);
or U6793 (N_6793,N_4736,N_2949);
or U6794 (N_6794,N_2538,N_2612);
xnor U6795 (N_6795,N_4848,N_3434);
or U6796 (N_6796,N_4035,N_2669);
nand U6797 (N_6797,N_3194,N_4437);
nand U6798 (N_6798,N_2896,N_4191);
and U6799 (N_6799,N_4851,N_3569);
nor U6800 (N_6800,N_2956,N_4415);
xnor U6801 (N_6801,N_4998,N_4271);
nor U6802 (N_6802,N_3859,N_3354);
xnor U6803 (N_6803,N_4600,N_3558);
nor U6804 (N_6804,N_2682,N_3072);
or U6805 (N_6805,N_3304,N_3399);
or U6806 (N_6806,N_4705,N_3166);
xor U6807 (N_6807,N_4096,N_3295);
and U6808 (N_6808,N_2636,N_3461);
nor U6809 (N_6809,N_3571,N_3984);
nand U6810 (N_6810,N_3199,N_4749);
nand U6811 (N_6811,N_4321,N_4888);
nand U6812 (N_6812,N_4210,N_3764);
xnor U6813 (N_6813,N_4807,N_3926);
xor U6814 (N_6814,N_4963,N_2540);
nor U6815 (N_6815,N_4046,N_3009);
or U6816 (N_6816,N_3224,N_2761);
nand U6817 (N_6817,N_3136,N_4059);
xnor U6818 (N_6818,N_2831,N_2677);
or U6819 (N_6819,N_3813,N_4193);
or U6820 (N_6820,N_3385,N_4054);
and U6821 (N_6821,N_3972,N_4238);
or U6822 (N_6822,N_3203,N_4715);
nand U6823 (N_6823,N_3613,N_4324);
nand U6824 (N_6824,N_4089,N_2770);
nand U6825 (N_6825,N_4579,N_2976);
nand U6826 (N_6826,N_2724,N_3175);
nor U6827 (N_6827,N_3543,N_4817);
or U6828 (N_6828,N_4927,N_2586);
nand U6829 (N_6829,N_3732,N_2767);
or U6830 (N_6830,N_4884,N_4468);
nand U6831 (N_6831,N_4167,N_4276);
or U6832 (N_6832,N_3503,N_2711);
nor U6833 (N_6833,N_4001,N_4253);
and U6834 (N_6834,N_4935,N_4201);
nor U6835 (N_6835,N_4742,N_4056);
xor U6836 (N_6836,N_4525,N_3574);
nor U6837 (N_6837,N_3345,N_2759);
or U6838 (N_6838,N_4321,N_4360);
nor U6839 (N_6839,N_4100,N_4284);
nor U6840 (N_6840,N_2628,N_3447);
or U6841 (N_6841,N_3019,N_2503);
nand U6842 (N_6842,N_4727,N_3327);
xor U6843 (N_6843,N_2945,N_4602);
or U6844 (N_6844,N_4727,N_3272);
xnor U6845 (N_6845,N_2981,N_2779);
and U6846 (N_6846,N_4272,N_3949);
nor U6847 (N_6847,N_3374,N_2990);
and U6848 (N_6848,N_2842,N_3973);
xor U6849 (N_6849,N_4233,N_4519);
nand U6850 (N_6850,N_4050,N_3486);
nor U6851 (N_6851,N_2524,N_3051);
nand U6852 (N_6852,N_3531,N_3428);
nor U6853 (N_6853,N_3518,N_2775);
xnor U6854 (N_6854,N_4220,N_4431);
and U6855 (N_6855,N_4316,N_3205);
and U6856 (N_6856,N_3196,N_3297);
nand U6857 (N_6857,N_3767,N_4800);
xnor U6858 (N_6858,N_2737,N_2833);
xnor U6859 (N_6859,N_3091,N_3730);
and U6860 (N_6860,N_4984,N_4547);
nor U6861 (N_6861,N_4863,N_4082);
nor U6862 (N_6862,N_2653,N_4585);
and U6863 (N_6863,N_4843,N_2797);
and U6864 (N_6864,N_4933,N_4115);
nand U6865 (N_6865,N_3128,N_3398);
or U6866 (N_6866,N_4400,N_3627);
nand U6867 (N_6867,N_4230,N_4153);
xor U6868 (N_6868,N_4379,N_3401);
nor U6869 (N_6869,N_3920,N_3405);
xnor U6870 (N_6870,N_3179,N_4262);
or U6871 (N_6871,N_4203,N_3933);
and U6872 (N_6872,N_2726,N_2999);
nand U6873 (N_6873,N_4567,N_4007);
nand U6874 (N_6874,N_3711,N_2956);
or U6875 (N_6875,N_3838,N_3900);
and U6876 (N_6876,N_4846,N_2974);
and U6877 (N_6877,N_4269,N_3130);
and U6878 (N_6878,N_3904,N_3758);
nor U6879 (N_6879,N_3648,N_4301);
and U6880 (N_6880,N_4916,N_2975);
xor U6881 (N_6881,N_3103,N_2605);
and U6882 (N_6882,N_3774,N_4077);
and U6883 (N_6883,N_2930,N_4314);
nor U6884 (N_6884,N_3472,N_2944);
and U6885 (N_6885,N_2929,N_4889);
and U6886 (N_6886,N_2863,N_3393);
nor U6887 (N_6887,N_3552,N_3462);
and U6888 (N_6888,N_3525,N_2760);
or U6889 (N_6889,N_4459,N_2706);
nor U6890 (N_6890,N_3896,N_3816);
xor U6891 (N_6891,N_4410,N_4303);
nand U6892 (N_6892,N_2799,N_4010);
xnor U6893 (N_6893,N_3733,N_4454);
nor U6894 (N_6894,N_3341,N_2696);
or U6895 (N_6895,N_3813,N_4345);
nor U6896 (N_6896,N_2693,N_3871);
nand U6897 (N_6897,N_4508,N_2798);
or U6898 (N_6898,N_2771,N_3911);
nor U6899 (N_6899,N_4271,N_4823);
nand U6900 (N_6900,N_4521,N_2696);
nor U6901 (N_6901,N_2819,N_4766);
xor U6902 (N_6902,N_4283,N_2565);
nor U6903 (N_6903,N_4266,N_3527);
nand U6904 (N_6904,N_4281,N_4168);
nor U6905 (N_6905,N_3436,N_3693);
and U6906 (N_6906,N_4805,N_3860);
nor U6907 (N_6907,N_2964,N_3871);
nand U6908 (N_6908,N_2767,N_3268);
nand U6909 (N_6909,N_4201,N_2817);
and U6910 (N_6910,N_4698,N_2612);
or U6911 (N_6911,N_2592,N_3516);
nor U6912 (N_6912,N_2588,N_3564);
or U6913 (N_6913,N_2529,N_2747);
and U6914 (N_6914,N_4042,N_4041);
nor U6915 (N_6915,N_3350,N_2772);
nor U6916 (N_6916,N_4097,N_3406);
and U6917 (N_6917,N_2887,N_3029);
or U6918 (N_6918,N_3277,N_4935);
nor U6919 (N_6919,N_4011,N_2648);
and U6920 (N_6920,N_2558,N_3980);
or U6921 (N_6921,N_2711,N_3192);
nand U6922 (N_6922,N_3335,N_2956);
or U6923 (N_6923,N_2869,N_4077);
nor U6924 (N_6924,N_4253,N_3651);
nand U6925 (N_6925,N_3762,N_3919);
xor U6926 (N_6926,N_3464,N_4469);
nand U6927 (N_6927,N_2507,N_4600);
nor U6928 (N_6928,N_3114,N_3104);
nand U6929 (N_6929,N_3198,N_3187);
and U6930 (N_6930,N_4178,N_3749);
nor U6931 (N_6931,N_2844,N_2654);
and U6932 (N_6932,N_4612,N_2938);
nor U6933 (N_6933,N_4946,N_3173);
xor U6934 (N_6934,N_3792,N_3406);
or U6935 (N_6935,N_2774,N_3553);
or U6936 (N_6936,N_4120,N_2968);
and U6937 (N_6937,N_2968,N_3561);
nand U6938 (N_6938,N_3905,N_3267);
or U6939 (N_6939,N_2779,N_4624);
and U6940 (N_6940,N_3445,N_3459);
or U6941 (N_6941,N_4453,N_3630);
xor U6942 (N_6942,N_4873,N_4982);
xnor U6943 (N_6943,N_4079,N_3307);
xnor U6944 (N_6944,N_2732,N_2590);
xor U6945 (N_6945,N_3200,N_2563);
and U6946 (N_6946,N_4616,N_3366);
nand U6947 (N_6947,N_3183,N_4009);
nor U6948 (N_6948,N_3983,N_4449);
xnor U6949 (N_6949,N_2858,N_4243);
nor U6950 (N_6950,N_4857,N_3742);
xor U6951 (N_6951,N_3283,N_2635);
or U6952 (N_6952,N_2585,N_4574);
or U6953 (N_6953,N_4992,N_2525);
nand U6954 (N_6954,N_3076,N_2750);
or U6955 (N_6955,N_4349,N_4125);
or U6956 (N_6956,N_4449,N_4142);
or U6957 (N_6957,N_3668,N_3921);
nand U6958 (N_6958,N_4785,N_2969);
and U6959 (N_6959,N_4761,N_3537);
xnor U6960 (N_6960,N_3349,N_3640);
nor U6961 (N_6961,N_2523,N_4989);
or U6962 (N_6962,N_2719,N_3660);
nand U6963 (N_6963,N_3491,N_2652);
or U6964 (N_6964,N_4043,N_2600);
or U6965 (N_6965,N_3569,N_3173);
and U6966 (N_6966,N_4004,N_4920);
nor U6967 (N_6967,N_4710,N_2762);
nand U6968 (N_6968,N_4711,N_4343);
nor U6969 (N_6969,N_3843,N_4901);
nor U6970 (N_6970,N_2943,N_4120);
nor U6971 (N_6971,N_4118,N_3581);
nor U6972 (N_6972,N_4945,N_2886);
xor U6973 (N_6973,N_4722,N_4548);
xnor U6974 (N_6974,N_4259,N_2665);
nand U6975 (N_6975,N_3293,N_4264);
or U6976 (N_6976,N_4945,N_2901);
and U6977 (N_6977,N_3589,N_4156);
nor U6978 (N_6978,N_4223,N_2535);
nor U6979 (N_6979,N_2639,N_4308);
nand U6980 (N_6980,N_2916,N_4375);
nand U6981 (N_6981,N_2645,N_3305);
xor U6982 (N_6982,N_3270,N_3375);
xnor U6983 (N_6983,N_2835,N_3083);
xnor U6984 (N_6984,N_4624,N_4896);
nor U6985 (N_6985,N_2875,N_3103);
nand U6986 (N_6986,N_4758,N_3328);
or U6987 (N_6987,N_4277,N_3486);
and U6988 (N_6988,N_3195,N_3971);
nand U6989 (N_6989,N_3109,N_3533);
or U6990 (N_6990,N_2514,N_3943);
or U6991 (N_6991,N_4697,N_4017);
nand U6992 (N_6992,N_3393,N_3363);
and U6993 (N_6993,N_2871,N_2814);
and U6994 (N_6994,N_4720,N_4497);
nand U6995 (N_6995,N_3859,N_2610);
nor U6996 (N_6996,N_3243,N_4549);
xnor U6997 (N_6997,N_4343,N_4786);
nor U6998 (N_6998,N_2920,N_2577);
nor U6999 (N_6999,N_3889,N_4268);
and U7000 (N_7000,N_3603,N_2999);
nor U7001 (N_7001,N_4001,N_2820);
and U7002 (N_7002,N_4630,N_3854);
or U7003 (N_7003,N_2855,N_3096);
xnor U7004 (N_7004,N_4179,N_4607);
xor U7005 (N_7005,N_3846,N_4967);
or U7006 (N_7006,N_3382,N_2851);
and U7007 (N_7007,N_2892,N_3116);
and U7008 (N_7008,N_4448,N_2707);
and U7009 (N_7009,N_2547,N_3729);
nand U7010 (N_7010,N_3564,N_2923);
and U7011 (N_7011,N_4319,N_4798);
xor U7012 (N_7012,N_2705,N_4799);
and U7013 (N_7013,N_4870,N_3407);
nand U7014 (N_7014,N_4289,N_3497);
nor U7015 (N_7015,N_3139,N_4874);
and U7016 (N_7016,N_4947,N_3868);
or U7017 (N_7017,N_2537,N_4703);
and U7018 (N_7018,N_3163,N_4980);
xnor U7019 (N_7019,N_4516,N_3845);
xnor U7020 (N_7020,N_3015,N_2755);
nor U7021 (N_7021,N_3549,N_3575);
nand U7022 (N_7022,N_3737,N_4987);
nor U7023 (N_7023,N_2570,N_4285);
or U7024 (N_7024,N_3887,N_4046);
nand U7025 (N_7025,N_2665,N_3661);
nand U7026 (N_7026,N_2789,N_3747);
or U7027 (N_7027,N_4288,N_3282);
xnor U7028 (N_7028,N_4450,N_3717);
nor U7029 (N_7029,N_2866,N_4169);
xnor U7030 (N_7030,N_4577,N_2725);
nor U7031 (N_7031,N_2803,N_3939);
and U7032 (N_7032,N_4818,N_4195);
or U7033 (N_7033,N_3549,N_4810);
nor U7034 (N_7034,N_4423,N_3116);
or U7035 (N_7035,N_3334,N_3590);
xor U7036 (N_7036,N_3384,N_4245);
and U7037 (N_7037,N_4160,N_4491);
nand U7038 (N_7038,N_4495,N_3642);
and U7039 (N_7039,N_3200,N_3568);
nand U7040 (N_7040,N_2651,N_4206);
or U7041 (N_7041,N_2941,N_4428);
nand U7042 (N_7042,N_2828,N_4143);
xor U7043 (N_7043,N_4819,N_4291);
xor U7044 (N_7044,N_4787,N_3630);
nand U7045 (N_7045,N_4846,N_3878);
and U7046 (N_7046,N_3441,N_4252);
nor U7047 (N_7047,N_2739,N_3919);
xnor U7048 (N_7048,N_4643,N_4942);
or U7049 (N_7049,N_3929,N_2759);
nand U7050 (N_7050,N_3609,N_3910);
or U7051 (N_7051,N_4009,N_3677);
xor U7052 (N_7052,N_4698,N_4363);
nor U7053 (N_7053,N_2728,N_2847);
xnor U7054 (N_7054,N_3064,N_2531);
nor U7055 (N_7055,N_3654,N_4507);
nand U7056 (N_7056,N_2537,N_4888);
nand U7057 (N_7057,N_4103,N_3629);
nand U7058 (N_7058,N_2510,N_4327);
xor U7059 (N_7059,N_4596,N_2764);
nand U7060 (N_7060,N_4452,N_3792);
xor U7061 (N_7061,N_4383,N_3228);
and U7062 (N_7062,N_4371,N_2533);
xnor U7063 (N_7063,N_2939,N_4929);
nor U7064 (N_7064,N_3355,N_4997);
or U7065 (N_7065,N_3994,N_4252);
and U7066 (N_7066,N_2787,N_2798);
nor U7067 (N_7067,N_4173,N_4923);
or U7068 (N_7068,N_3684,N_3231);
nor U7069 (N_7069,N_4701,N_4901);
xor U7070 (N_7070,N_3410,N_2629);
nor U7071 (N_7071,N_3458,N_2739);
and U7072 (N_7072,N_4540,N_3532);
and U7073 (N_7073,N_4511,N_2957);
or U7074 (N_7074,N_4345,N_3062);
xnor U7075 (N_7075,N_2718,N_4645);
nand U7076 (N_7076,N_4551,N_4734);
and U7077 (N_7077,N_2722,N_4781);
xor U7078 (N_7078,N_4644,N_3901);
nor U7079 (N_7079,N_4961,N_2942);
nand U7080 (N_7080,N_3162,N_4913);
or U7081 (N_7081,N_4583,N_3047);
xor U7082 (N_7082,N_4483,N_2607);
nand U7083 (N_7083,N_4001,N_2827);
and U7084 (N_7084,N_4964,N_4480);
nand U7085 (N_7085,N_3426,N_4412);
and U7086 (N_7086,N_3824,N_3787);
or U7087 (N_7087,N_4246,N_4510);
and U7088 (N_7088,N_4023,N_3387);
nor U7089 (N_7089,N_4122,N_4678);
and U7090 (N_7090,N_4259,N_3031);
nand U7091 (N_7091,N_3701,N_4234);
or U7092 (N_7092,N_3891,N_4719);
xnor U7093 (N_7093,N_4362,N_4194);
nor U7094 (N_7094,N_3980,N_3941);
nand U7095 (N_7095,N_4200,N_2923);
nor U7096 (N_7096,N_4061,N_3009);
or U7097 (N_7097,N_2942,N_3177);
nor U7098 (N_7098,N_4071,N_3806);
or U7099 (N_7099,N_4592,N_3331);
nand U7100 (N_7100,N_4492,N_4246);
xor U7101 (N_7101,N_4842,N_3448);
nand U7102 (N_7102,N_4139,N_3682);
or U7103 (N_7103,N_4436,N_3924);
and U7104 (N_7104,N_3909,N_3457);
and U7105 (N_7105,N_3149,N_4457);
nand U7106 (N_7106,N_3614,N_2535);
or U7107 (N_7107,N_4747,N_3664);
or U7108 (N_7108,N_3541,N_3925);
nor U7109 (N_7109,N_4204,N_3400);
xor U7110 (N_7110,N_2591,N_3630);
and U7111 (N_7111,N_3828,N_3673);
and U7112 (N_7112,N_3898,N_4585);
and U7113 (N_7113,N_2531,N_3684);
nor U7114 (N_7114,N_2896,N_3580);
nand U7115 (N_7115,N_3587,N_4533);
and U7116 (N_7116,N_4245,N_4351);
nand U7117 (N_7117,N_3261,N_3732);
and U7118 (N_7118,N_4364,N_3286);
xor U7119 (N_7119,N_2980,N_3425);
nand U7120 (N_7120,N_3288,N_4782);
nand U7121 (N_7121,N_4786,N_3222);
nor U7122 (N_7122,N_2524,N_2983);
nor U7123 (N_7123,N_4244,N_2568);
and U7124 (N_7124,N_3158,N_3152);
nor U7125 (N_7125,N_4557,N_4060);
or U7126 (N_7126,N_2600,N_3077);
and U7127 (N_7127,N_4489,N_2955);
nor U7128 (N_7128,N_3975,N_3555);
nand U7129 (N_7129,N_3755,N_4368);
nand U7130 (N_7130,N_4193,N_2557);
and U7131 (N_7131,N_3313,N_2690);
xor U7132 (N_7132,N_4312,N_3196);
nor U7133 (N_7133,N_4581,N_4664);
nand U7134 (N_7134,N_3459,N_2752);
and U7135 (N_7135,N_3181,N_4461);
or U7136 (N_7136,N_4396,N_4635);
nand U7137 (N_7137,N_3042,N_4222);
nor U7138 (N_7138,N_4080,N_4023);
xor U7139 (N_7139,N_4690,N_2908);
and U7140 (N_7140,N_2720,N_4020);
xnor U7141 (N_7141,N_4138,N_4806);
and U7142 (N_7142,N_4228,N_3210);
nor U7143 (N_7143,N_3635,N_3706);
or U7144 (N_7144,N_4212,N_3423);
nand U7145 (N_7145,N_3607,N_2643);
nand U7146 (N_7146,N_2682,N_3049);
xor U7147 (N_7147,N_3294,N_4182);
and U7148 (N_7148,N_2939,N_4190);
nor U7149 (N_7149,N_3820,N_3026);
or U7150 (N_7150,N_2943,N_4184);
nor U7151 (N_7151,N_4690,N_3791);
or U7152 (N_7152,N_4799,N_4656);
nor U7153 (N_7153,N_4134,N_3955);
xnor U7154 (N_7154,N_3858,N_3583);
nor U7155 (N_7155,N_4687,N_2710);
or U7156 (N_7156,N_3924,N_3983);
and U7157 (N_7157,N_3373,N_3140);
or U7158 (N_7158,N_2734,N_4473);
xor U7159 (N_7159,N_4044,N_4454);
xor U7160 (N_7160,N_3766,N_3476);
nor U7161 (N_7161,N_4665,N_3975);
xor U7162 (N_7162,N_3621,N_3256);
nand U7163 (N_7163,N_3522,N_2856);
xnor U7164 (N_7164,N_3216,N_4042);
nor U7165 (N_7165,N_3745,N_3926);
and U7166 (N_7166,N_3351,N_4897);
nor U7167 (N_7167,N_3539,N_4500);
or U7168 (N_7168,N_4418,N_4291);
or U7169 (N_7169,N_3115,N_3451);
nand U7170 (N_7170,N_3841,N_4646);
nand U7171 (N_7171,N_3416,N_3639);
nor U7172 (N_7172,N_2802,N_4328);
nor U7173 (N_7173,N_3524,N_4035);
nand U7174 (N_7174,N_2935,N_3006);
or U7175 (N_7175,N_2843,N_3745);
and U7176 (N_7176,N_3883,N_3310);
nor U7177 (N_7177,N_4284,N_3903);
xor U7178 (N_7178,N_3732,N_4488);
nor U7179 (N_7179,N_2711,N_3079);
nand U7180 (N_7180,N_2848,N_4034);
or U7181 (N_7181,N_3412,N_4174);
xor U7182 (N_7182,N_3836,N_3468);
or U7183 (N_7183,N_4915,N_4250);
or U7184 (N_7184,N_3911,N_4311);
or U7185 (N_7185,N_4954,N_2644);
or U7186 (N_7186,N_3433,N_2553);
or U7187 (N_7187,N_4509,N_3947);
nor U7188 (N_7188,N_4960,N_2678);
xor U7189 (N_7189,N_3758,N_4117);
xor U7190 (N_7190,N_2673,N_2529);
xnor U7191 (N_7191,N_2894,N_3798);
and U7192 (N_7192,N_4382,N_4626);
nand U7193 (N_7193,N_3602,N_4063);
nor U7194 (N_7194,N_3967,N_3997);
and U7195 (N_7195,N_4721,N_3700);
nand U7196 (N_7196,N_4987,N_4340);
nor U7197 (N_7197,N_3984,N_3955);
nand U7198 (N_7198,N_3140,N_3286);
or U7199 (N_7199,N_3900,N_4360);
xnor U7200 (N_7200,N_2726,N_4180);
xor U7201 (N_7201,N_4150,N_3214);
or U7202 (N_7202,N_4038,N_3988);
xor U7203 (N_7203,N_3169,N_2695);
nor U7204 (N_7204,N_3583,N_3518);
nand U7205 (N_7205,N_4827,N_3729);
xor U7206 (N_7206,N_4650,N_2762);
nand U7207 (N_7207,N_3481,N_4296);
and U7208 (N_7208,N_3928,N_3406);
and U7209 (N_7209,N_3201,N_4770);
nor U7210 (N_7210,N_3616,N_4628);
nand U7211 (N_7211,N_3426,N_4055);
and U7212 (N_7212,N_4076,N_3715);
nor U7213 (N_7213,N_3946,N_3157);
or U7214 (N_7214,N_3931,N_4714);
xor U7215 (N_7215,N_3076,N_3314);
and U7216 (N_7216,N_3133,N_3359);
xor U7217 (N_7217,N_3436,N_3241);
or U7218 (N_7218,N_4987,N_2707);
or U7219 (N_7219,N_3410,N_4464);
and U7220 (N_7220,N_4534,N_3569);
and U7221 (N_7221,N_4896,N_3581);
and U7222 (N_7222,N_4316,N_3556);
nand U7223 (N_7223,N_4054,N_4473);
or U7224 (N_7224,N_3536,N_2646);
xnor U7225 (N_7225,N_4949,N_2986);
or U7226 (N_7226,N_4447,N_4368);
nand U7227 (N_7227,N_3041,N_2840);
nand U7228 (N_7228,N_3807,N_3750);
xor U7229 (N_7229,N_3510,N_2780);
or U7230 (N_7230,N_4575,N_3441);
or U7231 (N_7231,N_3554,N_3455);
or U7232 (N_7232,N_4952,N_3490);
xnor U7233 (N_7233,N_2717,N_3323);
and U7234 (N_7234,N_4931,N_2831);
and U7235 (N_7235,N_2705,N_3459);
nor U7236 (N_7236,N_3858,N_4863);
and U7237 (N_7237,N_4936,N_3183);
xor U7238 (N_7238,N_3602,N_4502);
or U7239 (N_7239,N_2630,N_2877);
or U7240 (N_7240,N_3277,N_2969);
xor U7241 (N_7241,N_4907,N_3494);
and U7242 (N_7242,N_2707,N_4112);
and U7243 (N_7243,N_4916,N_4060);
or U7244 (N_7244,N_2503,N_4630);
and U7245 (N_7245,N_2606,N_3551);
xor U7246 (N_7246,N_3164,N_4299);
xnor U7247 (N_7247,N_4974,N_2518);
or U7248 (N_7248,N_3789,N_2794);
nor U7249 (N_7249,N_4168,N_3010);
and U7250 (N_7250,N_4116,N_3716);
xnor U7251 (N_7251,N_2990,N_4998);
or U7252 (N_7252,N_3812,N_3337);
nand U7253 (N_7253,N_4390,N_3459);
or U7254 (N_7254,N_2562,N_3986);
and U7255 (N_7255,N_3527,N_4130);
xor U7256 (N_7256,N_3103,N_4046);
and U7257 (N_7257,N_2721,N_3458);
nor U7258 (N_7258,N_4753,N_4290);
nor U7259 (N_7259,N_4177,N_4170);
xor U7260 (N_7260,N_3277,N_3743);
nor U7261 (N_7261,N_3963,N_4139);
nor U7262 (N_7262,N_2989,N_4274);
nor U7263 (N_7263,N_3448,N_2740);
xnor U7264 (N_7264,N_2591,N_3176);
and U7265 (N_7265,N_3647,N_3711);
nand U7266 (N_7266,N_3947,N_2832);
xor U7267 (N_7267,N_4327,N_2578);
nand U7268 (N_7268,N_2606,N_4426);
or U7269 (N_7269,N_4150,N_3200);
xor U7270 (N_7270,N_4014,N_4947);
and U7271 (N_7271,N_4510,N_4533);
nor U7272 (N_7272,N_2620,N_2989);
nand U7273 (N_7273,N_3908,N_2645);
nor U7274 (N_7274,N_3892,N_4111);
nor U7275 (N_7275,N_2605,N_3452);
or U7276 (N_7276,N_3470,N_4026);
or U7277 (N_7277,N_2576,N_3578);
and U7278 (N_7278,N_3886,N_4034);
xnor U7279 (N_7279,N_4395,N_4036);
and U7280 (N_7280,N_3250,N_4633);
or U7281 (N_7281,N_4596,N_4254);
xnor U7282 (N_7282,N_4678,N_2642);
xnor U7283 (N_7283,N_4741,N_3898);
and U7284 (N_7284,N_2790,N_3793);
nor U7285 (N_7285,N_2820,N_3350);
nand U7286 (N_7286,N_2864,N_4427);
nand U7287 (N_7287,N_4433,N_4686);
xor U7288 (N_7288,N_2568,N_3003);
xor U7289 (N_7289,N_2877,N_3817);
nand U7290 (N_7290,N_3244,N_2856);
and U7291 (N_7291,N_4597,N_4493);
nand U7292 (N_7292,N_3664,N_3431);
nor U7293 (N_7293,N_3522,N_3711);
or U7294 (N_7294,N_3555,N_2882);
xnor U7295 (N_7295,N_3501,N_3143);
nand U7296 (N_7296,N_4251,N_3029);
nand U7297 (N_7297,N_3066,N_4958);
nor U7298 (N_7298,N_4505,N_4142);
or U7299 (N_7299,N_4131,N_4113);
and U7300 (N_7300,N_3757,N_4141);
xnor U7301 (N_7301,N_4000,N_2809);
and U7302 (N_7302,N_4964,N_2744);
nor U7303 (N_7303,N_2939,N_2504);
and U7304 (N_7304,N_4841,N_2697);
nor U7305 (N_7305,N_4547,N_2706);
or U7306 (N_7306,N_4990,N_3491);
and U7307 (N_7307,N_3765,N_3808);
or U7308 (N_7308,N_3185,N_3004);
xor U7309 (N_7309,N_3497,N_4163);
and U7310 (N_7310,N_3697,N_4537);
xor U7311 (N_7311,N_2980,N_4809);
or U7312 (N_7312,N_3130,N_4986);
nor U7313 (N_7313,N_4813,N_3076);
nand U7314 (N_7314,N_4206,N_4821);
xor U7315 (N_7315,N_2558,N_3807);
and U7316 (N_7316,N_4009,N_4106);
nand U7317 (N_7317,N_4301,N_3124);
nor U7318 (N_7318,N_3257,N_3261);
xnor U7319 (N_7319,N_4588,N_2992);
and U7320 (N_7320,N_2718,N_4246);
nand U7321 (N_7321,N_3523,N_2506);
or U7322 (N_7322,N_2692,N_3037);
and U7323 (N_7323,N_3573,N_3246);
and U7324 (N_7324,N_3573,N_3623);
and U7325 (N_7325,N_4601,N_2975);
xnor U7326 (N_7326,N_3342,N_3416);
nor U7327 (N_7327,N_3610,N_4316);
nor U7328 (N_7328,N_2869,N_3072);
nand U7329 (N_7329,N_3371,N_3290);
xor U7330 (N_7330,N_2822,N_3803);
nand U7331 (N_7331,N_3534,N_4561);
xor U7332 (N_7332,N_3624,N_2645);
nand U7333 (N_7333,N_4024,N_4610);
xnor U7334 (N_7334,N_2876,N_4054);
xor U7335 (N_7335,N_3108,N_2788);
xnor U7336 (N_7336,N_3359,N_3499);
nand U7337 (N_7337,N_4715,N_3152);
xor U7338 (N_7338,N_4057,N_2552);
and U7339 (N_7339,N_2774,N_2708);
and U7340 (N_7340,N_3928,N_2817);
nand U7341 (N_7341,N_4457,N_4073);
nor U7342 (N_7342,N_4251,N_3896);
and U7343 (N_7343,N_3587,N_2666);
or U7344 (N_7344,N_4279,N_4568);
nand U7345 (N_7345,N_4055,N_2714);
nand U7346 (N_7346,N_4300,N_2576);
or U7347 (N_7347,N_4303,N_3538);
and U7348 (N_7348,N_4358,N_3671);
nand U7349 (N_7349,N_3152,N_4709);
and U7350 (N_7350,N_4150,N_2926);
nand U7351 (N_7351,N_4584,N_3683);
and U7352 (N_7352,N_2609,N_3849);
nor U7353 (N_7353,N_3260,N_2622);
xor U7354 (N_7354,N_4360,N_2528);
nand U7355 (N_7355,N_3599,N_4365);
and U7356 (N_7356,N_4129,N_3961);
and U7357 (N_7357,N_3199,N_4436);
nand U7358 (N_7358,N_4120,N_4059);
and U7359 (N_7359,N_2962,N_3627);
or U7360 (N_7360,N_4972,N_4580);
and U7361 (N_7361,N_3615,N_3852);
and U7362 (N_7362,N_3252,N_4388);
or U7363 (N_7363,N_4746,N_4638);
nand U7364 (N_7364,N_4506,N_4864);
nand U7365 (N_7365,N_2982,N_3321);
xor U7366 (N_7366,N_2586,N_4880);
xor U7367 (N_7367,N_3725,N_3236);
or U7368 (N_7368,N_4507,N_3832);
or U7369 (N_7369,N_3136,N_4454);
nor U7370 (N_7370,N_4252,N_2978);
and U7371 (N_7371,N_3569,N_3475);
xor U7372 (N_7372,N_2801,N_3745);
nor U7373 (N_7373,N_4610,N_4472);
nor U7374 (N_7374,N_3109,N_2524);
nor U7375 (N_7375,N_3771,N_4900);
nand U7376 (N_7376,N_3257,N_2993);
nor U7377 (N_7377,N_2752,N_3222);
or U7378 (N_7378,N_3681,N_3558);
or U7379 (N_7379,N_3340,N_3462);
or U7380 (N_7380,N_4136,N_3047);
and U7381 (N_7381,N_4830,N_4720);
xnor U7382 (N_7382,N_3873,N_4534);
and U7383 (N_7383,N_2951,N_3606);
nor U7384 (N_7384,N_2853,N_3499);
and U7385 (N_7385,N_2706,N_4998);
or U7386 (N_7386,N_3031,N_2784);
and U7387 (N_7387,N_3162,N_4086);
nor U7388 (N_7388,N_4899,N_4985);
nand U7389 (N_7389,N_4134,N_4192);
nor U7390 (N_7390,N_3309,N_3230);
or U7391 (N_7391,N_4596,N_4066);
nand U7392 (N_7392,N_4619,N_2936);
or U7393 (N_7393,N_3873,N_3978);
and U7394 (N_7394,N_3126,N_3534);
xor U7395 (N_7395,N_3741,N_3791);
nor U7396 (N_7396,N_3373,N_3808);
and U7397 (N_7397,N_4660,N_3653);
nand U7398 (N_7398,N_3630,N_3123);
xnor U7399 (N_7399,N_3328,N_4737);
and U7400 (N_7400,N_3669,N_3531);
nand U7401 (N_7401,N_4966,N_2569);
and U7402 (N_7402,N_4417,N_4665);
or U7403 (N_7403,N_4552,N_4252);
nand U7404 (N_7404,N_3719,N_2635);
and U7405 (N_7405,N_4352,N_4024);
or U7406 (N_7406,N_2776,N_3201);
nor U7407 (N_7407,N_2887,N_3896);
and U7408 (N_7408,N_4763,N_4025);
or U7409 (N_7409,N_3928,N_2630);
nor U7410 (N_7410,N_3404,N_4182);
nor U7411 (N_7411,N_2956,N_4254);
xor U7412 (N_7412,N_3145,N_4221);
nor U7413 (N_7413,N_4995,N_4480);
or U7414 (N_7414,N_4009,N_4006);
xnor U7415 (N_7415,N_4357,N_4805);
nor U7416 (N_7416,N_4139,N_3388);
nand U7417 (N_7417,N_3855,N_3731);
xnor U7418 (N_7418,N_4789,N_4393);
or U7419 (N_7419,N_4169,N_3131);
xor U7420 (N_7420,N_4364,N_3790);
xor U7421 (N_7421,N_3997,N_4783);
xor U7422 (N_7422,N_3168,N_4325);
xnor U7423 (N_7423,N_4488,N_2653);
or U7424 (N_7424,N_4343,N_2699);
xor U7425 (N_7425,N_3828,N_4495);
xor U7426 (N_7426,N_2701,N_3496);
xor U7427 (N_7427,N_4518,N_4272);
and U7428 (N_7428,N_3034,N_3137);
and U7429 (N_7429,N_3983,N_4376);
and U7430 (N_7430,N_3695,N_3322);
nand U7431 (N_7431,N_4831,N_2544);
or U7432 (N_7432,N_3589,N_2543);
and U7433 (N_7433,N_2875,N_4536);
xor U7434 (N_7434,N_3316,N_3729);
nor U7435 (N_7435,N_4143,N_4804);
or U7436 (N_7436,N_3983,N_3798);
nor U7437 (N_7437,N_4631,N_4741);
xnor U7438 (N_7438,N_3329,N_4827);
nand U7439 (N_7439,N_3392,N_3079);
xnor U7440 (N_7440,N_3128,N_4049);
xor U7441 (N_7441,N_2547,N_4618);
nor U7442 (N_7442,N_3665,N_3266);
or U7443 (N_7443,N_2663,N_4741);
nand U7444 (N_7444,N_4778,N_4587);
xnor U7445 (N_7445,N_4745,N_2977);
and U7446 (N_7446,N_3071,N_4057);
or U7447 (N_7447,N_3578,N_4767);
nor U7448 (N_7448,N_3425,N_2808);
nand U7449 (N_7449,N_3010,N_2820);
nand U7450 (N_7450,N_4699,N_3608);
or U7451 (N_7451,N_4803,N_3491);
nor U7452 (N_7452,N_4490,N_3034);
nor U7453 (N_7453,N_2782,N_2712);
or U7454 (N_7454,N_3676,N_3419);
nand U7455 (N_7455,N_4295,N_4740);
nand U7456 (N_7456,N_2652,N_3848);
and U7457 (N_7457,N_3212,N_3580);
nor U7458 (N_7458,N_4275,N_4737);
xor U7459 (N_7459,N_4598,N_4812);
nand U7460 (N_7460,N_4281,N_3264);
and U7461 (N_7461,N_3740,N_3215);
nor U7462 (N_7462,N_3449,N_3100);
and U7463 (N_7463,N_4092,N_4677);
or U7464 (N_7464,N_4495,N_4864);
nand U7465 (N_7465,N_4552,N_4366);
and U7466 (N_7466,N_3562,N_3956);
or U7467 (N_7467,N_4740,N_4434);
and U7468 (N_7468,N_2737,N_3954);
and U7469 (N_7469,N_4519,N_2882);
and U7470 (N_7470,N_4450,N_4728);
nor U7471 (N_7471,N_4351,N_3425);
and U7472 (N_7472,N_4103,N_4024);
or U7473 (N_7473,N_3546,N_4222);
nand U7474 (N_7474,N_3166,N_3586);
nor U7475 (N_7475,N_3236,N_3563);
and U7476 (N_7476,N_2928,N_4190);
xor U7477 (N_7477,N_4320,N_4072);
nor U7478 (N_7478,N_3793,N_2669);
xor U7479 (N_7479,N_4657,N_2628);
xor U7480 (N_7480,N_3480,N_2907);
or U7481 (N_7481,N_2822,N_3132);
and U7482 (N_7482,N_4858,N_2598);
and U7483 (N_7483,N_3577,N_3088);
nand U7484 (N_7484,N_2779,N_2934);
and U7485 (N_7485,N_4572,N_3296);
xnor U7486 (N_7486,N_4690,N_4932);
and U7487 (N_7487,N_4510,N_4993);
or U7488 (N_7488,N_3154,N_4430);
and U7489 (N_7489,N_4294,N_4711);
and U7490 (N_7490,N_3799,N_4343);
nor U7491 (N_7491,N_2698,N_4100);
or U7492 (N_7492,N_4086,N_4747);
nand U7493 (N_7493,N_3481,N_4521);
xnor U7494 (N_7494,N_4215,N_4125);
or U7495 (N_7495,N_3685,N_3139);
nor U7496 (N_7496,N_4169,N_3925);
or U7497 (N_7497,N_3169,N_4604);
xnor U7498 (N_7498,N_4696,N_2548);
nor U7499 (N_7499,N_4580,N_2865);
nor U7500 (N_7500,N_7201,N_5103);
nand U7501 (N_7501,N_6099,N_6459);
xor U7502 (N_7502,N_5212,N_5666);
nor U7503 (N_7503,N_5803,N_7106);
and U7504 (N_7504,N_7044,N_6771);
xnor U7505 (N_7505,N_5407,N_5262);
xnor U7506 (N_7506,N_6644,N_6097);
or U7507 (N_7507,N_5137,N_6108);
or U7508 (N_7508,N_5129,N_5758);
and U7509 (N_7509,N_6996,N_5729);
nand U7510 (N_7510,N_7089,N_7261);
nor U7511 (N_7511,N_6123,N_5419);
nor U7512 (N_7512,N_6820,N_5352);
and U7513 (N_7513,N_6679,N_7097);
xnor U7514 (N_7514,N_5717,N_6483);
or U7515 (N_7515,N_5934,N_6785);
nor U7516 (N_7516,N_6737,N_6125);
nand U7517 (N_7517,N_6580,N_6310);
and U7518 (N_7518,N_6609,N_5404);
nor U7519 (N_7519,N_7477,N_6723);
nand U7520 (N_7520,N_6654,N_6727);
and U7521 (N_7521,N_5799,N_7391);
or U7522 (N_7522,N_5764,N_6308);
nor U7523 (N_7523,N_7026,N_5241);
nand U7524 (N_7524,N_5821,N_7077);
or U7525 (N_7525,N_6700,N_7240);
nand U7526 (N_7526,N_5181,N_6544);
xnor U7527 (N_7527,N_7205,N_5588);
or U7528 (N_7528,N_7098,N_5708);
nand U7529 (N_7529,N_6074,N_5230);
and U7530 (N_7530,N_6047,N_5070);
or U7531 (N_7531,N_5011,N_7046);
nor U7532 (N_7532,N_5528,N_5947);
nor U7533 (N_7533,N_6332,N_5557);
and U7534 (N_7534,N_7042,N_6427);
or U7535 (N_7535,N_6300,N_5013);
or U7536 (N_7536,N_7185,N_6627);
or U7537 (N_7537,N_6681,N_5487);
and U7538 (N_7538,N_5967,N_5919);
or U7539 (N_7539,N_5582,N_7305);
nor U7540 (N_7540,N_7085,N_7349);
nor U7541 (N_7541,N_6794,N_5603);
nand U7542 (N_7542,N_6695,N_6792);
nand U7543 (N_7543,N_5434,N_5672);
or U7544 (N_7544,N_6212,N_6960);
xor U7545 (N_7545,N_7276,N_6676);
nor U7546 (N_7546,N_6063,N_7417);
nand U7547 (N_7547,N_6592,N_5598);
or U7548 (N_7548,N_6736,N_5705);
or U7549 (N_7549,N_6796,N_6340);
xor U7550 (N_7550,N_6640,N_6827);
nor U7551 (N_7551,N_5001,N_5278);
nand U7552 (N_7552,N_6545,N_5246);
xnor U7553 (N_7553,N_6263,N_5161);
and U7554 (N_7554,N_6940,N_5136);
and U7555 (N_7555,N_6957,N_5222);
nor U7556 (N_7556,N_5523,N_6755);
nor U7557 (N_7557,N_5816,N_6614);
or U7558 (N_7558,N_7292,N_7296);
or U7559 (N_7559,N_6174,N_7306);
nand U7560 (N_7560,N_5219,N_7142);
nand U7561 (N_7561,N_6774,N_7108);
nand U7562 (N_7562,N_6721,N_7325);
xnor U7563 (N_7563,N_6604,N_5951);
nand U7564 (N_7564,N_6902,N_6510);
and U7565 (N_7565,N_7423,N_5558);
or U7566 (N_7566,N_6479,N_6012);
nor U7567 (N_7567,N_6216,N_7063);
or U7568 (N_7568,N_5301,N_7490);
and U7569 (N_7569,N_6987,N_6296);
nand U7570 (N_7570,N_5379,N_6042);
nand U7571 (N_7571,N_5865,N_6766);
nand U7572 (N_7572,N_6178,N_6487);
nor U7573 (N_7573,N_6250,N_5007);
nand U7574 (N_7574,N_6936,N_5418);
and U7575 (N_7575,N_6791,N_5955);
or U7576 (N_7576,N_7177,N_5574);
and U7577 (N_7577,N_5913,N_6611);
or U7578 (N_7578,N_5794,N_5331);
or U7579 (N_7579,N_7485,N_6550);
nor U7580 (N_7580,N_6722,N_5525);
nand U7581 (N_7581,N_7336,N_5220);
nand U7582 (N_7582,N_7304,N_7147);
and U7583 (N_7583,N_6847,N_5748);
nand U7584 (N_7584,N_6666,N_6145);
and U7585 (N_7585,N_6441,N_6704);
or U7586 (N_7586,N_5151,N_6066);
or U7587 (N_7587,N_6151,N_7343);
nor U7588 (N_7588,N_5361,N_7429);
or U7589 (N_7589,N_6931,N_5494);
nand U7590 (N_7590,N_5527,N_6589);
or U7591 (N_7591,N_7321,N_5704);
xor U7592 (N_7592,N_5045,N_6092);
nand U7593 (N_7593,N_6008,N_6734);
and U7594 (N_7594,N_6065,N_5185);
nor U7595 (N_7595,N_6593,N_6435);
and U7596 (N_7596,N_5180,N_5746);
nor U7597 (N_7597,N_5747,N_7441);
or U7598 (N_7598,N_7288,N_6900);
and U7599 (N_7599,N_5012,N_7311);
xnor U7600 (N_7600,N_6881,N_6196);
and U7601 (N_7601,N_5818,N_6061);
xor U7602 (N_7602,N_5787,N_6130);
or U7603 (N_7603,N_6651,N_6619);
nand U7604 (N_7604,N_5398,N_5421);
xnor U7605 (N_7605,N_6261,N_7341);
nand U7606 (N_7606,N_5992,N_7189);
and U7607 (N_7607,N_6730,N_5851);
xor U7608 (N_7608,N_6307,N_5099);
nand U7609 (N_7609,N_6970,N_5192);
and U7610 (N_7610,N_6757,N_5941);
xnor U7611 (N_7611,N_5830,N_6244);
xnor U7612 (N_7612,N_6428,N_6558);
xnor U7613 (N_7613,N_6673,N_6852);
or U7614 (N_7614,N_6623,N_5634);
and U7615 (N_7615,N_7266,N_5432);
or U7616 (N_7616,N_5139,N_5786);
and U7617 (N_7617,N_6274,N_5079);
nor U7618 (N_7618,N_6253,N_7235);
or U7619 (N_7619,N_6457,N_6362);
and U7620 (N_7620,N_5148,N_7277);
or U7621 (N_7621,N_6056,N_5459);
nor U7622 (N_7622,N_5046,N_5107);
and U7623 (N_7623,N_5997,N_5422);
xor U7624 (N_7624,N_7209,N_6058);
or U7625 (N_7625,N_7264,N_7482);
nand U7626 (N_7626,N_5238,N_7013);
or U7627 (N_7627,N_6348,N_5145);
or U7628 (N_7628,N_6742,N_5049);
xor U7629 (N_7629,N_6893,N_6976);
and U7630 (N_7630,N_5840,N_5882);
xnor U7631 (N_7631,N_5338,N_5990);
xor U7632 (N_7632,N_7076,N_5092);
and U7633 (N_7633,N_6333,N_6193);
nor U7634 (N_7634,N_5020,N_6343);
nor U7635 (N_7635,N_6284,N_5184);
or U7636 (N_7636,N_5686,N_7181);
nand U7637 (N_7637,N_5682,N_5549);
or U7638 (N_7638,N_7080,N_6490);
nor U7639 (N_7639,N_7048,N_5206);
nand U7640 (N_7640,N_5548,N_6385);
and U7641 (N_7641,N_6769,N_5085);
xnor U7642 (N_7642,N_6842,N_6799);
and U7643 (N_7643,N_5039,N_6366);
nand U7644 (N_7644,N_5059,N_5820);
and U7645 (N_7645,N_7130,N_6773);
or U7646 (N_7646,N_7213,N_6001);
xor U7647 (N_7647,N_5502,N_5568);
or U7648 (N_7648,N_7449,N_6447);
and U7649 (N_7649,N_5730,N_5838);
xnor U7650 (N_7650,N_7475,N_5199);
xnor U7651 (N_7651,N_5295,N_5975);
nand U7652 (N_7652,N_6551,N_5797);
xnor U7653 (N_7653,N_6153,N_6071);
xnor U7654 (N_7654,N_5369,N_5844);
xor U7655 (N_7655,N_6152,N_7432);
nand U7656 (N_7656,N_6918,N_5625);
nand U7657 (N_7657,N_5687,N_6320);
or U7658 (N_7658,N_5669,N_5442);
or U7659 (N_7659,N_5304,N_7144);
xor U7660 (N_7660,N_7195,N_5940);
and U7661 (N_7661,N_6353,N_5963);
and U7662 (N_7662,N_6677,N_6210);
nor U7663 (N_7663,N_6562,N_6613);
nor U7664 (N_7664,N_5647,N_7274);
nand U7665 (N_7665,N_5397,N_5097);
nand U7666 (N_7666,N_7050,N_6475);
xor U7667 (N_7667,N_6607,N_6057);
and U7668 (N_7668,N_7236,N_7134);
nand U7669 (N_7669,N_5347,N_6655);
xnor U7670 (N_7670,N_5058,N_5389);
or U7671 (N_7671,N_5544,N_6081);
xor U7672 (N_7672,N_5133,N_5954);
xnor U7673 (N_7673,N_6669,N_5760);
nor U7674 (N_7674,N_7180,N_7334);
and U7675 (N_7675,N_7251,N_7453);
nand U7676 (N_7676,N_6121,N_5392);
and U7677 (N_7677,N_5564,N_5035);
or U7678 (N_7678,N_6361,N_5655);
and U7679 (N_7679,N_7102,N_7227);
or U7680 (N_7680,N_6197,N_6854);
xor U7681 (N_7681,N_6392,N_5567);
nand U7682 (N_7682,N_6582,N_6078);
xnor U7683 (N_7683,N_5885,N_6059);
and U7684 (N_7684,N_7281,N_6237);
nand U7685 (N_7685,N_6405,N_5073);
xnor U7686 (N_7686,N_6207,N_6528);
nand U7687 (N_7687,N_6860,N_6387);
nand U7688 (N_7688,N_6663,N_5646);
or U7689 (N_7689,N_5834,N_7173);
nor U7690 (N_7690,N_5929,N_5636);
and U7691 (N_7691,N_6961,N_5839);
and U7692 (N_7692,N_5066,N_5120);
nand U7693 (N_7693,N_7022,N_5871);
and U7694 (N_7694,N_6840,N_5330);
nor U7695 (N_7695,N_6922,N_7123);
and U7696 (N_7696,N_5341,N_6950);
nor U7697 (N_7697,N_5648,N_7265);
nor U7698 (N_7698,N_5062,N_5375);
nor U7699 (N_7699,N_6468,N_6920);
nand U7700 (N_7700,N_5431,N_5956);
nor U7701 (N_7701,N_6632,N_7388);
and U7702 (N_7702,N_7379,N_5436);
nand U7703 (N_7703,N_6530,N_7069);
or U7704 (N_7704,N_7182,N_5460);
nor U7705 (N_7705,N_6132,N_5287);
or U7706 (N_7706,N_7335,N_6648);
nor U7707 (N_7707,N_5660,N_6466);
xnor U7708 (N_7708,N_7090,N_6705);
nor U7709 (N_7709,N_5978,N_5470);
xnor U7710 (N_7710,N_7163,N_7405);
or U7711 (N_7711,N_5365,N_6981);
xnor U7712 (N_7712,N_5521,N_6511);
xnor U7713 (N_7713,N_5089,N_5401);
nand U7714 (N_7714,N_7132,N_6371);
or U7715 (N_7715,N_5350,N_5877);
and U7716 (N_7716,N_6618,N_7499);
or U7717 (N_7717,N_6233,N_6815);
and U7718 (N_7718,N_6688,N_5325);
or U7719 (N_7719,N_5736,N_7148);
nand U7720 (N_7720,N_7114,N_6911);
and U7721 (N_7721,N_5363,N_6497);
nor U7722 (N_7722,N_5609,N_5115);
and U7723 (N_7723,N_6650,N_5987);
xnor U7724 (N_7724,N_5353,N_6040);
or U7725 (N_7725,N_7422,N_7184);
nor U7726 (N_7726,N_7060,N_6697);
nor U7727 (N_7727,N_5541,N_6195);
and U7728 (N_7728,N_5626,N_6819);
nor U7729 (N_7729,N_6298,N_5328);
nor U7730 (N_7730,N_5154,N_6455);
nor U7731 (N_7731,N_7316,N_6994);
and U7732 (N_7732,N_6539,N_5600);
nand U7733 (N_7733,N_6703,N_6763);
nor U7734 (N_7734,N_6407,N_6044);
nand U7735 (N_7735,N_5677,N_6281);
nor U7736 (N_7736,N_5750,N_5004);
nor U7737 (N_7737,N_6738,N_7027);
and U7738 (N_7738,N_7263,N_5033);
xnor U7739 (N_7739,N_5909,N_6275);
or U7740 (N_7740,N_7474,N_5996);
or U7741 (N_7741,N_7468,N_5171);
nand U7742 (N_7742,N_6805,N_5593);
nor U7743 (N_7743,N_6485,N_6778);
nand U7744 (N_7744,N_7062,N_7197);
or U7745 (N_7745,N_5825,N_5195);
nor U7746 (N_7746,N_5141,N_6595);
and U7747 (N_7747,N_5356,N_6579);
nor U7748 (N_7748,N_7283,N_5500);
nor U7749 (N_7749,N_5320,N_6780);
or U7750 (N_7750,N_6553,N_7394);
or U7751 (N_7751,N_5713,N_7176);
or U7752 (N_7752,N_7211,N_7471);
xor U7753 (N_7753,N_7293,N_5991);
and U7754 (N_7754,N_5780,N_6315);
xor U7755 (N_7755,N_5306,N_6027);
nand U7756 (N_7756,N_7437,N_5209);
nor U7757 (N_7757,N_5025,N_6873);
or U7758 (N_7758,N_7245,N_6083);
nor U7759 (N_7759,N_5125,N_7234);
or U7760 (N_7760,N_6127,N_5800);
nor U7761 (N_7761,N_5441,N_6921);
and U7762 (N_7762,N_6807,N_7220);
xnor U7763 (N_7763,N_7014,N_7055);
and U7764 (N_7764,N_6895,N_6601);
and U7765 (N_7765,N_6830,N_6594);
and U7766 (N_7766,N_7366,N_6100);
and U7767 (N_7767,N_5057,N_5709);
and U7768 (N_7768,N_5453,N_7435);
nand U7769 (N_7769,N_7011,N_6329);
nand U7770 (N_7770,N_5444,N_7465);
nand U7771 (N_7771,N_7492,N_5901);
nor U7772 (N_7772,N_5715,N_6825);
nor U7773 (N_7773,N_6832,N_6512);
or U7774 (N_7774,N_6519,N_7020);
and U7775 (N_7775,N_6710,N_6255);
and U7776 (N_7776,N_5198,N_5552);
nor U7777 (N_7777,N_7150,N_6509);
xnor U7778 (N_7778,N_5783,N_7312);
and U7779 (N_7779,N_6844,N_7346);
or U7780 (N_7780,N_7156,N_6942);
nand U7781 (N_7781,N_5152,N_5305);
nor U7782 (N_7782,N_6891,N_5386);
nand U7783 (N_7783,N_5086,N_5428);
xor U7784 (N_7784,N_5205,N_6414);
and U7785 (N_7785,N_6449,N_6713);
and U7786 (N_7786,N_5383,N_5740);
nor U7787 (N_7787,N_5989,N_7408);
xor U7788 (N_7788,N_6653,N_6469);
xnor U7789 (N_7789,N_5359,N_7337);
nor U7790 (N_7790,N_6659,N_5250);
and U7791 (N_7791,N_6880,N_5894);
and U7792 (N_7792,N_7479,N_7302);
or U7793 (N_7793,N_6735,N_5981);
xor U7794 (N_7794,N_6876,N_5875);
or U7795 (N_7795,N_5316,N_7496);
or U7796 (N_7796,N_7332,N_6326);
xor U7797 (N_7797,N_6213,N_7291);
and U7798 (N_7798,N_5081,N_5255);
xor U7799 (N_7799,N_7088,N_6913);
nand U7800 (N_7800,N_5000,N_6200);
xnor U7801 (N_7801,N_5679,N_7255);
nand U7802 (N_7802,N_6184,N_6146);
and U7803 (N_7803,N_6919,N_6616);
nand U7804 (N_7804,N_6941,N_5067);
xnor U7805 (N_7805,N_7112,N_6947);
nand U7806 (N_7806,N_7351,N_5024);
nor U7807 (N_7807,N_5455,N_6055);
nor U7808 (N_7808,N_6465,N_6354);
or U7809 (N_7809,N_6016,N_6529);
xnor U7810 (N_7810,N_7420,N_6583);
xor U7811 (N_7811,N_5656,N_6818);
and U7812 (N_7812,N_6328,N_7052);
nor U7813 (N_7813,N_5360,N_5368);
and U7814 (N_7814,N_5961,N_5477);
xnor U7815 (N_7815,N_5326,N_5569);
nand U7816 (N_7816,N_5918,N_6024);
xor U7817 (N_7817,N_5591,N_6954);
and U7818 (N_7818,N_5869,N_5906);
or U7819 (N_7819,N_5972,N_5256);
or U7820 (N_7820,N_6576,N_7393);
nand U7821 (N_7821,N_7442,N_7212);
nand U7822 (N_7822,N_6495,N_7401);
xor U7823 (N_7823,N_6339,N_5400);
or U7824 (N_7824,N_6090,N_5769);
or U7825 (N_7825,N_5566,N_5619);
xor U7826 (N_7826,N_6002,N_6462);
or U7827 (N_7827,N_7072,N_6882);
and U7828 (N_7828,N_6101,N_7171);
or U7829 (N_7829,N_5638,N_5364);
nand U7830 (N_7830,N_6128,N_6686);
nand U7831 (N_7831,N_5688,N_6064);
xor U7832 (N_7832,N_6559,N_7071);
or U7833 (N_7833,N_5560,N_6242);
nand U7834 (N_7834,N_6452,N_5731);
xor U7835 (N_7835,N_6404,N_5578);
or U7836 (N_7836,N_6772,N_5795);
nand U7837 (N_7837,N_7010,N_5102);
xor U7838 (N_7838,N_5118,N_5068);
xnor U7839 (N_7839,N_6739,N_5908);
and U7840 (N_7840,N_7323,N_5433);
nand U7841 (N_7841,N_5023,N_6269);
or U7842 (N_7842,N_7233,N_5244);
xnor U7843 (N_7843,N_7258,N_6522);
or U7844 (N_7844,N_5737,N_7051);
nand U7845 (N_7845,N_7015,N_7404);
or U7846 (N_7846,N_6980,N_6965);
or U7847 (N_7847,N_5604,N_6998);
nor U7848 (N_7848,N_6678,N_7356);
and U7849 (N_7849,N_5545,N_6481);
nor U7850 (N_7850,N_5164,N_7095);
nor U7851 (N_7851,N_6273,N_7398);
nor U7852 (N_7852,N_5165,N_7457);
xor U7853 (N_7853,N_5738,N_5707);
nand U7854 (N_7854,N_5060,N_5734);
and U7855 (N_7855,N_5468,N_6630);
and U7856 (N_7856,N_5083,N_6859);
and U7857 (N_7857,N_6206,N_6718);
and U7858 (N_7858,N_6227,N_6508);
nand U7859 (N_7859,N_6926,N_6603);
nor U7860 (N_7860,N_5970,N_5505);
nand U7861 (N_7861,N_5718,N_6394);
nand U7862 (N_7862,N_6496,N_6674);
or U7863 (N_7863,N_5105,N_5607);
nor U7864 (N_7864,N_6637,N_7267);
or U7865 (N_7865,N_5644,N_6163);
or U7866 (N_7866,N_5358,N_5514);
and U7867 (N_7867,N_5334,N_6527);
or U7868 (N_7868,N_6743,N_5637);
xnor U7869 (N_7869,N_6500,N_6471);
or U7870 (N_7870,N_7428,N_6868);
and U7871 (N_7871,N_6937,N_6685);
nor U7872 (N_7872,N_6748,N_5510);
nor U7873 (N_7873,N_7023,N_5823);
and U7874 (N_7874,N_7152,N_6573);
xnor U7875 (N_7875,N_7074,N_6089);
xor U7876 (N_7876,N_5778,N_5503);
nand U7877 (N_7877,N_6857,N_5131);
nor U7878 (N_7878,N_5518,N_6235);
nand U7879 (N_7879,N_5631,N_5275);
and U7880 (N_7880,N_5156,N_7295);
nand U7881 (N_7881,N_6246,N_7116);
or U7882 (N_7882,N_6075,N_5022);
nand U7883 (N_7883,N_6955,N_5471);
and U7884 (N_7884,N_6491,N_7355);
nand U7885 (N_7885,N_5651,N_6124);
nor U7886 (N_7886,N_6378,N_5583);
nand U7887 (N_7887,N_6817,N_7068);
nor U7888 (N_7888,N_6399,N_6964);
nand U7889 (N_7889,N_6069,N_5168);
and U7890 (N_7890,N_7057,N_5610);
and U7891 (N_7891,N_6276,N_7438);
or U7892 (N_7892,N_5050,N_6989);
and U7893 (N_7893,N_5504,N_6978);
xnor U7894 (N_7894,N_5917,N_6549);
nor U7895 (N_7895,N_5466,N_5472);
nand U7896 (N_7896,N_6232,N_5010);
and U7897 (N_7897,N_6265,N_6953);
or U7898 (N_7898,N_6105,N_6203);
and U7899 (N_7899,N_5700,N_6706);
nor U7900 (N_7900,N_6547,N_5124);
or U7901 (N_7901,N_6716,N_6758);
xor U7902 (N_7902,N_6289,N_7115);
xnor U7903 (N_7903,N_5339,N_6806);
xor U7904 (N_7904,N_6999,N_5891);
and U7905 (N_7905,N_5411,N_7330);
nor U7906 (N_7906,N_7183,N_5114);
or U7907 (N_7907,N_6131,N_6183);
or U7908 (N_7908,N_6661,N_7118);
and U7909 (N_7909,N_5333,N_6241);
or U7910 (N_7910,N_5935,N_6162);
nand U7911 (N_7911,N_7472,N_5971);
and U7912 (N_7912,N_6386,N_7228);
xor U7913 (N_7913,N_6897,N_6513);
nor U7914 (N_7914,N_6341,N_6260);
nor U7915 (N_7915,N_7459,N_6973);
nand U7916 (N_7916,N_7392,N_6812);
xnor U7917 (N_7917,N_5930,N_5678);
xor U7918 (N_7918,N_6336,N_5053);
and U7919 (N_7919,N_6988,N_7287);
and U7920 (N_7920,N_5807,N_6556);
and U7921 (N_7921,N_5848,N_6762);
nand U7922 (N_7922,N_6541,N_7386);
or U7923 (N_7923,N_5692,N_7226);
nor U7924 (N_7924,N_6238,N_6109);
and U7925 (N_7925,N_7455,N_5135);
nand U7926 (N_7926,N_5367,N_6903);
and U7927 (N_7927,N_5123,N_5710);
nand U7928 (N_7928,N_6413,N_6605);
xor U7929 (N_7929,N_6759,N_5489);
nor U7930 (N_7930,N_7488,N_5966);
nor U7931 (N_7931,N_5868,N_6804);
xor U7932 (N_7932,N_6137,N_5041);
or U7933 (N_7933,N_6194,N_7053);
xnor U7934 (N_7934,N_6231,N_5897);
and U7935 (N_7935,N_5061,N_5064);
nand U7936 (N_7936,N_7324,N_6294);
nand U7937 (N_7937,N_5695,N_7091);
or U7938 (N_7938,N_6768,N_6888);
and U7939 (N_7939,N_5801,N_5052);
and U7940 (N_7940,N_5481,N_5349);
xnor U7941 (N_7941,N_6085,N_7446);
nor U7942 (N_7942,N_6221,N_7411);
xnor U7943 (N_7943,N_5071,N_7344);
nand U7944 (N_7944,N_7041,N_5814);
xor U7945 (N_7945,N_7476,N_5577);
or U7946 (N_7946,N_5841,N_5292);
xnor U7947 (N_7947,N_6641,N_6568);
and U7948 (N_7948,N_5486,N_5575);
and U7949 (N_7949,N_7206,N_6201);
or U7950 (N_7950,N_6323,N_5296);
nor U7951 (N_7951,N_5706,N_6956);
or U7952 (N_7952,N_7252,N_6094);
xnor U7953 (N_7953,N_6262,N_6358);
xnor U7954 (N_7954,N_5146,N_5265);
nor U7955 (N_7955,N_6486,N_6014);
xnor U7956 (N_7956,N_5533,N_6438);
or U7957 (N_7957,N_6161,N_5374);
nand U7958 (N_7958,N_5149,N_5988);
nor U7959 (N_7959,N_6802,N_6835);
nor U7960 (N_7960,N_5535,N_5158);
and U7961 (N_7961,N_5615,N_6301);
and U7962 (N_7962,N_6403,N_6561);
or U7963 (N_7963,N_6138,N_5924);
and U7964 (N_7964,N_6581,N_5539);
nand U7965 (N_7965,N_7329,N_5017);
nand U7966 (N_7966,N_5828,N_6297);
and U7967 (N_7967,N_6598,N_5307);
and U7968 (N_7968,N_6098,N_6456);
or U7969 (N_7969,N_5405,N_6220);
and U7970 (N_7970,N_6177,N_6389);
or U7971 (N_7971,N_5040,N_6744);
xor U7972 (N_7972,N_5259,N_7430);
xor U7973 (N_7973,N_6377,N_7162);
nand U7974 (N_7974,N_6949,N_7169);
or U7975 (N_7975,N_7421,N_5283);
nor U7976 (N_7976,N_6464,N_7038);
nand U7977 (N_7977,N_7259,N_5670);
xor U7978 (N_7978,N_7113,N_6420);
nor U7979 (N_7979,N_6570,N_6434);
and U7980 (N_7980,N_6687,N_5658);
nor U7981 (N_7981,N_6437,N_6072);
and U7982 (N_7982,N_5775,N_5298);
or U7983 (N_7983,N_5624,N_5649);
nor U7984 (N_7984,N_7003,N_6367);
and U7985 (N_7985,N_6173,N_7406);
and U7986 (N_7986,N_6877,N_5417);
xor U7987 (N_7987,N_5112,N_5620);
or U7988 (N_7988,N_7122,N_6375);
nand U7989 (N_7989,N_7390,N_5571);
and U7990 (N_7990,N_6597,N_6446);
nand U7991 (N_7991,N_5597,N_5993);
xnor U7992 (N_7992,N_7443,N_6181);
or U7993 (N_7993,N_7047,N_5888);
xor U7994 (N_7994,N_6102,N_6645);
nand U7995 (N_7995,N_7460,N_7061);
and U7996 (N_7996,N_5529,N_5811);
and U7997 (N_7997,N_5138,N_5870);
or U7998 (N_7998,N_7275,N_6110);
nand U7999 (N_7999,N_7229,N_5332);
nor U8000 (N_8000,N_6565,N_7307);
xnor U8001 (N_8001,N_6566,N_6525);
and U8002 (N_8002,N_6370,N_6425);
and U8003 (N_8003,N_5754,N_7214);
or U8004 (N_8004,N_7222,N_6277);
and U8005 (N_8005,N_5110,N_7188);
and U8006 (N_8006,N_5284,N_5663);
xor U8007 (N_8007,N_6652,N_7400);
or U8008 (N_8008,N_5380,N_7489);
and U8009 (N_8009,N_5898,N_7269);
nand U8010 (N_8010,N_5479,N_6176);
or U8011 (N_8011,N_5813,N_5080);
nor U8012 (N_8012,N_5446,N_7225);
xnor U8013 (N_8013,N_5237,N_5534);
nor U8014 (N_8014,N_5030,N_7143);
and U8015 (N_8015,N_5735,N_6192);
or U8016 (N_8016,N_6187,N_6571);
xor U8017 (N_8017,N_6963,N_5457);
xnor U8018 (N_8018,N_5458,N_6866);
and U8019 (N_8019,N_7049,N_6388);
and U8020 (N_8020,N_7375,N_6788);
or U8021 (N_8021,N_6741,N_5394);
nand U8022 (N_8022,N_5408,N_6314);
nand U8023 (N_8023,N_6731,N_5104);
or U8024 (N_8024,N_6728,N_6076);
and U8025 (N_8025,N_5815,N_6114);
nand U8026 (N_8026,N_5055,N_6808);
nand U8027 (N_8027,N_6005,N_5895);
and U8028 (N_8028,N_7216,N_7359);
nor U8029 (N_8029,N_7110,N_6144);
and U8030 (N_8030,N_6638,N_7194);
and U8031 (N_8031,N_6560,N_6312);
xnor U8032 (N_8032,N_5182,N_5042);
nor U8033 (N_8033,N_5665,N_6790);
xnor U8034 (N_8034,N_5785,N_5480);
nand U8035 (N_8035,N_6331,N_6346);
or U8036 (N_8036,N_6383,N_5200);
or U8037 (N_8037,N_5088,N_6930);
nand U8038 (N_8038,N_5822,N_5618);
and U8039 (N_8039,N_5999,N_5308);
or U8040 (N_8040,N_5054,N_5570);
and U8041 (N_8041,N_5712,N_6856);
nor U8042 (N_8042,N_5832,N_5240);
nor U8043 (N_8043,N_5765,N_6251);
or U8044 (N_8044,N_5303,N_5281);
and U8045 (N_8045,N_7456,N_6974);
or U8046 (N_8046,N_7362,N_5409);
nand U8047 (N_8047,N_5986,N_6885);
nor U8048 (N_8048,N_5804,N_7272);
nand U8049 (N_8049,N_6675,N_6875);
or U8050 (N_8050,N_5627,N_6683);
nand U8051 (N_8051,N_7187,N_5142);
xor U8052 (N_8052,N_5346,N_6453);
nor U8053 (N_8053,N_7407,N_7320);
or U8054 (N_8054,N_6908,N_7029);
xnor U8055 (N_8055,N_7299,N_5810);
nor U8056 (N_8056,N_5854,N_5725);
or U8057 (N_8057,N_6429,N_6038);
xnor U8058 (N_8058,N_5202,N_7270);
nor U8059 (N_8059,N_5561,N_6430);
or U8060 (N_8060,N_5743,N_5274);
xor U8061 (N_8061,N_6691,N_6168);
xor U8062 (N_8062,N_6306,N_5351);
xnor U8063 (N_8063,N_5236,N_5884);
and U8064 (N_8064,N_6169,N_7444);
xnor U8065 (N_8065,N_6523,N_5953);
or U8066 (N_8066,N_5002,N_5973);
or U8067 (N_8067,N_6170,N_7202);
nor U8068 (N_8068,N_6282,N_6628);
nand U8069 (N_8069,N_5449,N_6849);
nor U8070 (N_8070,N_6190,N_5196);
and U8071 (N_8071,N_7434,N_5464);
nand U8072 (N_8072,N_7093,N_7371);
nand U8073 (N_8073,N_7354,N_6382);
and U8074 (N_8074,N_6499,N_6458);
and U8075 (N_8075,N_6803,N_5921);
nand U8076 (N_8076,N_5792,N_6629);
xor U8077 (N_8077,N_6033,N_5980);
and U8078 (N_8078,N_7018,N_6770);
nor U8079 (N_8079,N_5983,N_6118);
nor U8080 (N_8080,N_6436,N_7294);
xnor U8081 (N_8081,N_5447,N_7413);
xnor U8082 (N_8082,N_6816,N_6858);
xor U8083 (N_8083,N_7157,N_7369);
and U8084 (N_8084,N_6958,N_6256);
nor U8085 (N_8085,N_7105,N_6801);
xor U8086 (N_8086,N_6480,N_5269);
xor U8087 (N_8087,N_6322,N_6694);
or U8088 (N_8088,N_6962,N_7254);
nand U8089 (N_8089,N_6711,N_7491);
xnor U8090 (N_8090,N_7248,N_5866);
nor U8091 (N_8091,N_5177,N_5323);
xnor U8092 (N_8092,N_6381,N_6208);
xor U8093 (N_8093,N_5362,N_6658);
nor U8094 (N_8094,N_7317,N_6062);
xor U8095 (N_8095,N_7483,N_7378);
nand U8096 (N_8096,N_5858,N_6423);
nor U8097 (N_8097,N_7452,N_7200);
and U8098 (N_8098,N_7120,N_5019);
nand U8099 (N_8099,N_5957,N_6945);
xor U8100 (N_8100,N_5874,N_6935);
and U8101 (N_8101,N_6997,N_5217);
xor U8102 (N_8102,N_6342,N_5886);
xnor U8103 (N_8103,N_5159,N_5109);
nor U8104 (N_8104,N_6898,N_5632);
nand U8105 (N_8105,N_5853,N_6712);
nor U8106 (N_8106,N_5289,N_5872);
or U8107 (N_8107,N_5044,N_5291);
or U8108 (N_8108,N_5623,N_7387);
and U8109 (N_8109,N_5772,N_5257);
or U8110 (N_8110,N_5420,N_7131);
or U8111 (N_8111,N_6234,N_6984);
nor U8112 (N_8112,N_6051,N_5629);
and U8113 (N_8113,N_5005,N_5793);
and U8114 (N_8114,N_6717,N_6543);
nor U8115 (N_8115,N_5856,N_5208);
and U8116 (N_8116,N_5694,N_6117);
xnor U8117 (N_8117,N_6372,N_5267);
nand U8118 (N_8118,N_7040,N_7243);
xnor U8119 (N_8119,N_6909,N_6927);
nand U8120 (N_8120,N_6800,N_5861);
or U8121 (N_8121,N_6148,N_6247);
nor U8122 (N_8122,N_5440,N_6548);
nor U8123 (N_8123,N_6225,N_6878);
xor U8124 (N_8124,N_6087,N_6321);
xnor U8125 (N_8125,N_6134,N_5532);
xor U8126 (N_8126,N_6018,N_5370);
nor U8127 (N_8127,N_6907,N_6043);
and U8128 (N_8128,N_5399,N_5995);
or U8129 (N_8129,N_5524,N_6280);
or U8130 (N_8130,N_5319,N_6944);
nor U8131 (N_8131,N_6222,N_5722);
nor U8132 (N_8132,N_6702,N_5312);
nor U8133 (N_8133,N_5314,N_7347);
or U8134 (N_8134,N_6243,N_7462);
or U8135 (N_8135,N_5507,N_6209);
and U8136 (N_8136,N_5642,N_5662);
or U8137 (N_8137,N_6442,N_5667);
nand U8138 (N_8138,N_6380,N_6271);
and U8139 (N_8139,N_5675,N_5761);
and U8140 (N_8140,N_5488,N_5454);
nand U8141 (N_8141,N_5430,N_6337);
nand U8142 (N_8142,N_6082,N_5482);
nor U8143 (N_8143,N_6356,N_6503);
and U8144 (N_8144,N_5936,N_5258);
nand U8145 (N_8145,N_7230,N_7019);
and U8146 (N_8146,N_6670,N_6848);
nor U8147 (N_8147,N_5766,N_5095);
or U8148 (N_8148,N_5461,N_7215);
nand U8149 (N_8149,N_6096,N_6506);
and U8150 (N_8150,N_5122,N_5563);
xnor U8151 (N_8151,N_7463,N_6412);
nand U8152 (N_8152,N_5438,N_6606);
nor U8153 (N_8153,N_6460,N_6657);
and U8154 (N_8154,N_6959,N_5197);
nor U8155 (N_8155,N_5857,N_6521);
and U8156 (N_8156,N_7239,N_6990);
and U8157 (N_8157,N_7124,N_6439);
xnor U8158 (N_8158,N_7383,N_6303);
nand U8159 (N_8159,N_6635,N_6030);
and U8160 (N_8160,N_7094,N_5286);
or U8161 (N_8161,N_7340,N_6224);
nand U8162 (N_8162,N_6890,N_5210);
or U8163 (N_8163,N_5923,N_7286);
and U8164 (N_8164,N_5538,N_7361);
nand U8165 (N_8165,N_5952,N_5231);
nor U8166 (N_8166,N_6448,N_5849);
nand U8167 (N_8167,N_6482,N_7253);
nor U8168 (N_8168,N_5031,N_6175);
and U8169 (N_8169,N_6865,N_6517);
nor U8170 (N_8170,N_6313,N_6290);
nor U8171 (N_8171,N_5594,N_7313);
xor U8172 (N_8172,N_5998,N_5659);
xor U8173 (N_8173,N_5491,N_6398);
xor U8174 (N_8174,N_5213,N_7161);
nor U8175 (N_8175,N_6636,N_5587);
and U8176 (N_8176,N_5391,N_5806);
nand U8177 (N_8177,N_7058,N_5467);
and U8178 (N_8178,N_6732,N_6472);
and U8179 (N_8179,N_7374,N_5911);
nand U8180 (N_8180,N_5193,N_5390);
nor U8181 (N_8181,N_5904,N_6349);
nand U8182 (N_8182,N_6985,N_6833);
nor U8183 (N_8183,N_6843,N_7466);
nor U8184 (N_8184,N_5452,N_5203);
nand U8185 (N_8185,N_5628,N_5429);
xor U8186 (N_8186,N_6749,N_6838);
xnor U8187 (N_8187,N_7199,N_7121);
nor U8188 (N_8188,N_6664,N_6376);
nand U8189 (N_8189,N_6218,N_5224);
xnor U8190 (N_8190,N_5008,N_7043);
and U8191 (N_8191,N_5643,N_5382);
or U8192 (N_8192,N_6113,N_5580);
nand U8193 (N_8193,N_7409,N_7416);
xor U8194 (N_8194,N_7001,N_6248);
xor U8195 (N_8195,N_7005,N_5768);
and U8196 (N_8196,N_5311,N_6440);
xnor U8197 (N_8197,N_7099,N_5721);
and U8198 (N_8198,N_6054,N_5513);
and U8199 (N_8199,N_6133,N_6784);
xnor U8200 (N_8200,N_5728,N_6408);
nor U8201 (N_8201,N_6526,N_5753);
and U8202 (N_8202,N_7168,N_5711);
and U8203 (N_8203,N_6564,N_5423);
or U8204 (N_8204,N_5096,N_6968);
nor U8205 (N_8205,N_7450,N_5641);
and U8206 (N_8206,N_5762,N_7190);
nor U8207 (N_8207,N_7223,N_7458);
or U8208 (N_8208,N_5106,N_6596);
nand U8209 (N_8209,N_7360,N_5693);
or U8210 (N_8210,N_6286,N_7327);
nor U8211 (N_8211,N_6896,N_5029);
or U8212 (N_8212,N_6690,N_6951);
and U8213 (N_8213,N_6726,N_6318);
and U8214 (N_8214,N_5490,N_5342);
and U8215 (N_8215,N_6330,N_7352);
or U8216 (N_8216,N_5279,N_7493);
and U8217 (N_8217,N_7191,N_5661);
or U8218 (N_8218,N_6837,N_6364);
nand U8219 (N_8219,N_6390,N_7480);
and U8220 (N_8220,N_5959,N_6714);
nand U8221 (N_8221,N_5896,N_7364);
xor U8222 (N_8222,N_7487,N_6139);
nor U8223 (N_8223,N_7192,N_6292);
and U8224 (N_8224,N_5416,N_6760);
nand U8225 (N_8225,N_6202,N_5119);
xnor U8226 (N_8226,N_7384,N_5779);
xor U8227 (N_8227,N_5697,N_7141);
nand U8228 (N_8228,N_5579,N_5819);
nand U8229 (N_8229,N_6924,N_6514);
nand U8230 (N_8230,N_5774,N_5690);
nand U8231 (N_8231,N_6967,N_7024);
nand U8232 (N_8232,N_6786,N_6285);
xor U8233 (N_8233,N_5985,N_5859);
nor U8234 (N_8234,N_7363,N_6540);
xor U8235 (N_8235,N_6359,N_7415);
or U8236 (N_8236,N_6259,N_6905);
nand U8237 (N_8237,N_7280,N_5469);
and U8238 (N_8238,N_5691,N_5976);
and U8239 (N_8239,N_5300,N_5565);
and U8240 (N_8240,N_6116,N_6050);
xnor U8241 (N_8241,N_6906,N_7418);
or U8242 (N_8242,N_5584,N_5613);
nor U8243 (N_8243,N_5611,N_6295);
nand U8244 (N_8244,N_6013,N_5167);
nand U8245 (N_8245,N_7498,N_5297);
nor U8246 (N_8246,N_5724,N_7339);
xor U8247 (N_8247,N_6590,N_6140);
and U8248 (N_8248,N_5633,N_6156);
nor U8249 (N_8249,N_5384,N_5939);
xor U8250 (N_8250,N_5727,N_5355);
nand U8251 (N_8251,N_5069,N_6324);
nand U8252 (N_8252,N_6524,N_7059);
and U8253 (N_8253,N_6186,N_6928);
and U8254 (N_8254,N_5437,N_5701);
nand U8255 (N_8255,N_6258,N_7308);
nand U8256 (N_8256,N_6095,N_5645);
nor U8257 (N_8257,N_5962,N_5302);
xor U8258 (N_8258,N_6810,N_5555);
nor U8259 (N_8259,N_5048,N_7037);
and U8260 (N_8260,N_6239,N_5551);
nand U8261 (N_8261,N_6916,N_5497);
xnor U8262 (N_8262,N_7160,N_6662);
nor U8263 (N_8263,N_6272,N_5026);
nor U8264 (N_8264,N_6397,N_6557);
nand U8265 (N_8265,N_6115,N_7389);
and U8266 (N_8266,N_6478,N_5476);
xor U8267 (N_8267,N_6534,N_7310);
and U8268 (N_8268,N_5852,N_7469);
xnor U8269 (N_8269,N_5671,N_5047);
or U8270 (N_8270,N_5251,N_7345);
xnor U8271 (N_8271,N_5403,N_5522);
or U8272 (N_8272,N_7309,N_6003);
nor U8273 (N_8273,N_6991,N_7410);
and U8274 (N_8274,N_6620,N_6536);
nor U8275 (N_8275,N_5261,N_6518);
or U8276 (N_8276,N_5128,N_7007);
and U8277 (N_8277,N_6135,N_5247);
nor U8278 (N_8278,N_7414,N_5932);
or U8279 (N_8279,N_5945,N_6871);
nor U8280 (N_8280,N_6391,N_7232);
nor U8281 (N_8281,N_5664,N_7380);
nand U8282 (N_8282,N_5835,N_7137);
nand U8283 (N_8283,N_5556,N_6185);
nand U8284 (N_8284,N_6172,N_6041);
nor U8285 (N_8285,N_6424,N_6889);
nor U8286 (N_8286,N_6080,N_5234);
nand U8287 (N_8287,N_5435,N_6923);
and U8288 (N_8288,N_5268,N_6841);
or U8289 (N_8289,N_7224,N_6418);
or U8290 (N_8290,N_6166,N_6829);
nand U8291 (N_8291,N_7377,N_5140);
nand U8292 (N_8292,N_5475,N_5335);
nor U8293 (N_8293,N_5689,N_5276);
nand U8294 (N_8294,N_5887,N_6572);
nor U8295 (N_8295,N_6776,N_6761);
xnor U8296 (N_8296,N_5372,N_5902);
xnor U8297 (N_8297,N_6473,N_5867);
xnor U8298 (N_8298,N_5742,N_7031);
and U8299 (N_8299,N_5183,N_5021);
nand U8300 (N_8300,N_7056,N_5091);
or U8301 (N_8301,N_5817,N_6680);
nand U8302 (N_8302,N_6198,N_6591);
xnor U8303 (N_8303,N_6091,N_7328);
nor U8304 (N_8304,N_6019,N_5445);
nand U8305 (N_8305,N_6334,N_5554);
and U8306 (N_8306,N_6360,N_6846);
nand U8307 (N_8307,N_5243,N_6709);
xnor U8308 (N_8308,N_5227,N_5680);
or U8309 (N_8309,N_6395,N_7145);
and U8310 (N_8310,N_6751,N_7082);
and U8311 (N_8311,N_6288,N_7045);
and U8312 (N_8312,N_7250,N_7136);
nand U8313 (N_8313,N_5673,N_6787);
and U8314 (N_8314,N_5425,N_5674);
xor U8315 (N_8315,N_5218,N_7025);
and U8316 (N_8316,N_7244,N_5880);
nor U8317 (N_8317,N_6781,N_6402);
or U8318 (N_8318,N_5337,N_5340);
or U8319 (N_8319,N_7279,N_5617);
and U8320 (N_8320,N_7238,N_7125);
nand U8321 (N_8321,N_5831,N_6671);
and U8322 (N_8322,N_5547,N_6304);
xnor U8323 (N_8323,N_7382,N_5038);
nand U8324 (N_8324,N_5927,N_6396);
nand U8325 (N_8325,N_6291,N_5396);
or U8326 (N_8326,N_5890,N_5946);
and U8327 (N_8327,N_6914,N_6179);
nand U8328 (N_8328,N_6068,N_5493);
nor U8329 (N_8329,N_6915,N_6707);
xor U8330 (N_8330,N_5899,N_6910);
xor U8331 (N_8331,N_5414,N_5016);
nor U8332 (N_8332,N_7273,N_5280);
xnor U8333 (N_8333,N_7032,N_5925);
and U8334 (N_8334,N_6498,N_6350);
or U8335 (N_8335,N_6729,N_7314);
xnor U8336 (N_8336,N_5833,N_7427);
nand U8337 (N_8337,N_6575,N_6347);
nor U8338 (N_8338,N_6104,N_7070);
xnor U8339 (N_8339,N_6979,N_6266);
xor U8340 (N_8340,N_6432,N_5499);
nand U8341 (N_8341,N_7436,N_5696);
xor U8342 (N_8342,N_5948,N_7111);
nand U8343 (N_8343,N_5395,N_5260);
xnor U8344 (N_8344,N_5915,N_6938);
nor U8345 (N_8345,N_6982,N_5117);
or U8346 (N_8346,N_7372,N_5366);
xnor U8347 (N_8347,N_5075,N_5492);
xor U8348 (N_8348,N_5702,N_6489);
and U8349 (N_8349,N_7473,N_7155);
nand U8350 (N_8350,N_5526,N_5776);
and U8351 (N_8351,N_5796,N_6143);
nand U8352 (N_8352,N_5937,N_5090);
and U8353 (N_8353,N_5170,N_5511);
or U8354 (N_8354,N_6665,N_6649);
nor U8355 (N_8355,N_6445,N_6507);
and U8356 (N_8356,N_7175,N_5344);
xnor U8357 (N_8357,N_6765,N_6443);
or U8358 (N_8358,N_5150,N_5829);
or U8359 (N_8359,N_5272,N_6492);
nand U8360 (N_8360,N_5842,N_5512);
nor U8361 (N_8361,N_5484,N_6715);
xor U8362 (N_8362,N_5881,N_5608);
or U8363 (N_8363,N_5676,N_5153);
nand U8364 (N_8364,N_5540,N_6775);
or U8365 (N_8365,N_5169,N_5354);
nand U8366 (N_8366,N_5893,N_6720);
nand U8367 (N_8367,N_5699,N_5456);
xnor U8368 (N_8368,N_5406,N_7174);
xnor U8369 (N_8369,N_7412,N_5322);
nand U8370 (N_8370,N_5232,N_7333);
and U8371 (N_8371,N_7289,N_5006);
nand U8372 (N_8372,N_6867,N_5744);
xnor U8373 (N_8373,N_6421,N_5763);
nand U8374 (N_8374,N_6698,N_5739);
nand U8375 (N_8375,N_6783,N_7439);
and U8376 (N_8376,N_7318,N_7301);
nor U8377 (N_8377,N_5530,N_6567);
nand U8378 (N_8378,N_5373,N_5944);
nand U8379 (N_8379,N_5519,N_6164);
and U8380 (N_8380,N_6205,N_6745);
nand U8381 (N_8381,N_6626,N_5933);
or U8382 (N_8382,N_5448,N_5984);
or U8383 (N_8383,N_6643,N_6103);
and U8384 (N_8384,N_5716,N_5860);
xor U8385 (N_8385,N_5850,N_6352);
or U8386 (N_8386,N_5393,N_6992);
nor U8387 (N_8387,N_5752,N_5108);
and U8388 (N_8388,N_6035,N_7448);
nand U8389 (N_8389,N_7064,N_6719);
and U8390 (N_8390,N_5843,N_6634);
nor U8391 (N_8391,N_7006,N_6625);
and U8392 (N_8392,N_6814,N_6037);
or U8393 (N_8393,N_5263,N_5501);
and U8394 (N_8394,N_5266,N_5111);
or U8395 (N_8395,N_6204,N_6129);
nor U8396 (N_8396,N_5223,N_6136);
or U8397 (N_8397,N_6855,N_5264);
nor U8398 (N_8398,N_5155,N_7117);
and U8399 (N_8399,N_5982,N_6532);
and U8400 (N_8400,N_7376,N_6624);
xnor U8401 (N_8401,N_5950,N_6226);
or U8402 (N_8402,N_5595,N_7033);
or U8403 (N_8403,N_5789,N_6569);
xnor U8404 (N_8404,N_5271,N_5698);
nor U8405 (N_8405,N_5463,N_5703);
and U8406 (N_8406,N_5376,N_6824);
nand U8407 (N_8407,N_6850,N_5515);
or U8408 (N_8408,N_6049,N_6777);
nor U8409 (N_8409,N_5270,N_5309);
nand U8410 (N_8410,N_6191,N_6077);
nor U8411 (N_8411,N_6007,N_5321);
nor U8412 (N_8412,N_5254,N_5683);
xnor U8413 (N_8413,N_5187,N_7139);
nand U8414 (N_8414,N_5015,N_5965);
nand U8415 (N_8415,N_7079,N_5134);
or U8416 (N_8416,N_6126,N_6584);
nor U8417 (N_8417,N_6939,N_6107);
nand U8418 (N_8418,N_7140,N_6283);
or U8419 (N_8419,N_5537,N_6159);
nand U8420 (N_8420,N_6839,N_6901);
or U8421 (N_8421,N_5027,N_5883);
or U8422 (N_8422,N_6267,N_6211);
nor U8423 (N_8423,N_6317,N_5317);
and U8424 (N_8424,N_6585,N_6693);
xor U8425 (N_8425,N_6070,N_6045);
nand U8426 (N_8426,N_7067,N_6599);
and U8427 (N_8427,N_7034,N_6836);
nor U8428 (N_8428,N_6393,N_6554);
and U8429 (N_8429,N_7154,N_5979);
or U8430 (N_8430,N_5229,N_5032);
nor U8431 (N_8431,N_7358,N_5756);
nor U8432 (N_8432,N_5862,N_6245);
or U8433 (N_8433,N_5076,N_5864);
or U8434 (N_8434,N_7285,N_5616);
nor U8435 (N_8435,N_7073,N_7119);
or U8436 (N_8436,N_6149,N_6165);
nor U8437 (N_8437,N_6764,N_5282);
nor U8438 (N_8438,N_6067,N_7447);
nand U8439 (N_8439,N_6171,N_7164);
nor U8440 (N_8440,N_6983,N_5586);
xor U8441 (N_8441,N_7084,N_5100);
nor U8442 (N_8442,N_5905,N_5876);
nor U8443 (N_8443,N_7247,N_5116);
and U8444 (N_8444,N_5777,N_6029);
or U8445 (N_8445,N_6684,N_6384);
or U8446 (N_8446,N_6182,N_5836);
nor U8447 (N_8447,N_6588,N_7204);
xor U8448 (N_8448,N_5974,N_7107);
nor U8449 (N_8449,N_6752,N_6409);
or U8450 (N_8450,N_6355,N_5313);
or U8451 (N_8451,N_5249,N_7196);
and U8452 (N_8452,N_5074,N_7101);
xnor U8453 (N_8453,N_7365,N_6932);
nor U8454 (N_8454,N_5808,N_7178);
nor U8455 (N_8455,N_6120,N_5847);
nor U8456 (N_8456,N_6552,N_5043);
nand U8457 (N_8457,N_6444,N_5837);
nor U8458 (N_8458,N_7081,N_7036);
nor U8459 (N_8459,N_6270,N_5508);
xnor U8460 (N_8460,N_7065,N_6293);
nand U8461 (N_8461,N_5573,N_6365);
nand U8462 (N_8462,N_6060,N_7242);
xnor U8463 (N_8463,N_5443,N_5606);
and U8464 (N_8464,N_5410,N_6416);
or U8465 (N_8465,N_7300,N_5147);
nor U8466 (N_8466,N_6111,N_5784);
or U8467 (N_8467,N_5473,N_6555);
nor U8468 (N_8468,N_6943,N_7440);
or U8469 (N_8469,N_5639,N_5173);
xor U8470 (N_8470,N_6422,N_5413);
xor U8471 (N_8471,N_6887,N_7425);
and U8472 (N_8472,N_7271,N_5179);
nand U8473 (N_8473,N_5242,N_5907);
or U8474 (N_8474,N_6899,N_5176);
or U8475 (N_8475,N_6009,N_6756);
or U8476 (N_8476,N_6287,N_6006);
nor U8477 (N_8477,N_5190,N_7451);
or U8478 (N_8478,N_5900,N_7326);
nor U8479 (N_8479,N_5654,N_7338);
and U8480 (N_8480,N_6410,N_5130);
xnor U8481 (N_8481,N_5969,N_5290);
or U8482 (N_8482,N_6879,N_6533);
xor U8483 (N_8483,N_7179,N_5226);
xor U8484 (N_8484,N_6401,N_7017);
or U8485 (N_8485,N_6531,N_5132);
nand U8486 (N_8486,N_5653,N_6869);
or U8487 (N_8487,N_6725,N_7484);
or U8488 (N_8488,N_6488,N_5077);
nor U8489 (N_8489,N_7424,N_5174);
nor U8490 (N_8490,N_6079,N_5812);
nand U8491 (N_8491,N_6039,N_5798);
or U8492 (N_8492,N_5113,N_6966);
xnor U8493 (N_8493,N_6157,N_6608);
and U8494 (N_8494,N_6022,N_5163);
xnor U8495 (N_8495,N_7028,N_6053);
xnor U8496 (N_8496,N_5590,N_6011);
nor U8497 (N_8497,N_5233,N_6577);
or U8498 (N_8498,N_6821,N_7478);
or U8499 (N_8499,N_5723,N_7186);
or U8500 (N_8500,N_7092,N_7083);
and U8501 (N_8501,N_5402,N_7153);
or U8502 (N_8502,N_5928,N_5788);
xor U8503 (N_8503,N_5720,N_6369);
and U8504 (N_8504,N_6021,N_5635);
xnor U8505 (N_8505,N_5098,N_5093);
and U8506 (N_8506,N_7221,N_7127);
or U8507 (N_8507,N_6325,N_5439);
or U8508 (N_8508,N_5640,N_5612);
xor U8509 (N_8509,N_6746,N_5749);
and U8510 (N_8510,N_5157,N_5191);
and U8511 (N_8511,N_7241,N_5621);
xor U8512 (N_8512,N_5790,N_6279);
nand U8513 (N_8513,N_5087,N_7086);
or U8514 (N_8514,N_6870,N_6642);
nor U8515 (N_8515,N_5630,N_5770);
xor U8516 (N_8516,N_5585,N_5496);
or U8517 (N_8517,N_6311,N_5977);
or U8518 (N_8518,N_5755,N_5914);
xnor U8519 (N_8519,N_6793,N_5826);
xor U8520 (N_8520,N_5681,N_6160);
or U8521 (N_8521,N_5542,N_7397);
xor U8522 (N_8522,N_5426,N_7315);
xnor U8523 (N_8523,N_5188,N_7193);
nand U8524 (N_8524,N_6587,N_5520);
xor U8525 (N_8525,N_7207,N_6689);
xnor U8526 (N_8526,N_5028,N_6917);
and U8527 (N_8527,N_6451,N_5543);
or U8528 (N_8528,N_7350,N_7035);
and U8529 (N_8529,N_5878,N_5451);
nand U8530 (N_8530,N_7016,N_7495);
xor U8531 (N_8531,N_6463,N_5931);
xnor U8532 (N_8532,N_5485,N_6733);
nand U8533 (N_8533,N_5288,N_7012);
nor U8534 (N_8534,N_7135,N_5596);
nand U8535 (N_8535,N_6946,N_7431);
or U8536 (N_8536,N_6701,N_6419);
or U8537 (N_8537,N_7385,N_7260);
and U8538 (N_8538,N_5166,N_6305);
or U8539 (N_8539,N_5388,N_5357);
and U8540 (N_8540,N_5964,N_6150);
xor U8541 (N_8541,N_6215,N_5378);
and U8542 (N_8542,N_6344,N_6750);
nor U8543 (N_8543,N_5294,N_6933);
or U8544 (N_8544,N_7039,N_7172);
nand U8545 (N_8545,N_5387,N_5845);
nand U8546 (N_8546,N_6667,N_5873);
or U8547 (N_8547,N_7419,N_6023);
nand U8548 (N_8548,N_5498,N_7373);
or U8549 (N_8549,N_6327,N_6264);
or U8550 (N_8550,N_5175,N_6345);
nor U8551 (N_8551,N_6505,N_6894);
nand U8552 (N_8552,N_7268,N_6032);
xnor U8553 (N_8553,N_6025,N_5879);
xnor U8554 (N_8554,N_6335,N_5767);
nor U8555 (N_8555,N_6199,N_6219);
and U8556 (N_8556,N_7357,N_5741);
or U8557 (N_8557,N_7297,N_6546);
xor U8558 (N_8558,N_7303,N_6740);
nand U8559 (N_8559,N_7368,N_7481);
nor U8560 (N_8560,N_6502,N_6000);
or U8561 (N_8561,N_5474,N_6026);
or U8562 (N_8562,N_5942,N_6823);
nand U8563 (N_8563,N_6086,N_5903);
nor U8564 (N_8564,N_5343,N_7217);
or U8565 (N_8565,N_5034,N_6031);
nor U8566 (N_8566,N_5143,N_5299);
nor U8567 (N_8567,N_6612,N_5009);
and U8568 (N_8568,N_6217,N_6046);
and U8569 (N_8569,N_5381,N_7008);
nand U8570 (N_8570,N_6782,N_6986);
or U8571 (N_8571,N_6797,N_5782);
nand U8572 (N_8572,N_7284,N_5221);
nand U8573 (N_8573,N_5824,N_6600);
nor U8574 (N_8574,N_5949,N_5248);
or U8575 (N_8575,N_6892,N_5652);
xor U8576 (N_8576,N_7159,N_6574);
and U8577 (N_8577,N_6048,N_6724);
xnor U8578 (N_8578,N_7246,N_5745);
nor U8579 (N_8579,N_6229,N_5204);
or U8580 (N_8580,N_6853,N_6036);
and U8581 (N_8581,N_5912,N_6017);
nand U8582 (N_8582,N_6338,N_5450);
nor U8583 (N_8583,N_5277,N_7231);
or U8584 (N_8584,N_5214,N_7461);
nand U8585 (N_8585,N_6863,N_5315);
nand U8586 (N_8586,N_6975,N_5225);
nor U8587 (N_8587,N_7170,N_5327);
nand U8588 (N_8588,N_5684,N_7403);
nand U8589 (N_8589,N_5072,N_7096);
xor U8590 (N_8590,N_6316,N_6813);
nor U8591 (N_8591,N_7151,N_6610);
xnor U8592 (N_8592,N_7218,N_6052);
nand U8593 (N_8593,N_5318,N_6309);
nand U8594 (N_8594,N_5773,N_5802);
or U8595 (N_8595,N_6374,N_6972);
nand U8596 (N_8596,N_7087,N_6180);
nor U8597 (N_8597,N_5516,N_5791);
or U8598 (N_8598,N_7138,N_6020);
nand U8599 (N_8599,N_5827,N_7370);
and U8600 (N_8600,N_6668,N_5336);
xnor U8601 (N_8601,N_6257,N_7256);
xnor U8602 (N_8602,N_6537,N_7104);
xor U8603 (N_8603,N_5889,N_5014);
nand U8604 (N_8604,N_5324,N_5051);
xnor U8605 (N_8605,N_5759,N_5685);
nor U8606 (N_8606,N_6084,N_5245);
and U8607 (N_8607,N_6252,N_7467);
nand U8608 (N_8608,N_6621,N_6106);
or U8609 (N_8609,N_5509,N_7426);
xnor U8610 (N_8610,N_6494,N_7078);
and U8611 (N_8611,N_6299,N_6692);
nor U8612 (N_8612,N_5178,N_5172);
nand U8613 (N_8613,N_5385,N_6779);
nor U8614 (N_8614,N_6158,N_6516);
xor U8615 (N_8615,N_5235,N_6798);
and U8616 (N_8616,N_7381,N_5056);
and U8617 (N_8617,N_6167,N_6477);
or U8618 (N_8618,N_5726,N_7149);
or U8619 (N_8619,N_5506,N_5121);
or U8620 (N_8620,N_6426,N_5968);
or U8621 (N_8621,N_5994,N_5036);
and U8622 (N_8622,N_7319,N_5216);
and U8623 (N_8623,N_7000,N_5194);
and U8624 (N_8624,N_5348,N_5650);
and U8625 (N_8625,N_5189,N_5733);
or U8626 (N_8626,N_5253,N_7009);
or U8627 (N_8627,N_6155,N_6474);
or U8628 (N_8628,N_5063,N_7396);
and U8629 (N_8629,N_6929,N_6538);
and U8630 (N_8630,N_6154,N_5424);
nor U8631 (N_8631,N_6406,N_5546);
nand U8632 (N_8632,N_6230,N_6602);
xor U8633 (N_8633,N_5082,N_7203);
nor U8634 (N_8634,N_6433,N_5732);
nor U8635 (N_8635,N_6699,N_5614);
nand U8636 (N_8636,N_7342,N_6119);
nand U8637 (N_8637,N_5562,N_6993);
nor U8638 (N_8638,N_6223,N_6834);
nor U8639 (N_8639,N_5605,N_5714);
or U8640 (N_8640,N_5938,N_7219);
and U8641 (N_8641,N_7322,N_6249);
nor U8642 (N_8642,N_5273,N_6969);
xor U8643 (N_8643,N_6925,N_7198);
nor U8644 (N_8644,N_7158,N_7290);
xor U8645 (N_8645,N_7353,N_6351);
nor U8646 (N_8646,N_6368,N_6948);
nand U8647 (N_8647,N_6515,N_7109);
nand U8648 (N_8648,N_7257,N_6268);
xnor U8649 (N_8649,N_7399,N_5201);
nor U8650 (N_8650,N_6015,N_7054);
nor U8651 (N_8651,N_7278,N_6363);
nor U8652 (N_8652,N_7133,N_7146);
nand U8653 (N_8653,N_7262,N_7470);
or U8654 (N_8654,N_5846,N_6415);
nor U8655 (N_8655,N_6952,N_5037);
nor U8656 (N_8656,N_6883,N_7066);
nor U8657 (N_8657,N_6753,N_7237);
nor U8658 (N_8658,N_6476,N_5855);
or U8659 (N_8659,N_5916,N_7100);
or U8660 (N_8660,N_5228,N_5581);
or U8661 (N_8661,N_6656,N_6493);
nor U8662 (N_8662,N_5252,N_6028);
and U8663 (N_8663,N_5805,N_5757);
or U8664 (N_8664,N_6886,N_6672);
xor U8665 (N_8665,N_6622,N_7210);
and U8666 (N_8666,N_6484,N_6417);
and U8667 (N_8667,N_6789,N_6971);
and U8668 (N_8668,N_7348,N_6617);
nor U8669 (N_8669,N_6795,N_7395);
nor U8670 (N_8670,N_5126,N_5719);
or U8671 (N_8671,N_6501,N_5207);
nand U8672 (N_8672,N_6122,N_6826);
nor U8673 (N_8673,N_6811,N_5483);
nor U8674 (N_8674,N_7494,N_6142);
or U8675 (N_8675,N_5589,N_7331);
xor U8676 (N_8676,N_5602,N_6431);
and U8677 (N_8677,N_7166,N_6278);
nor U8678 (N_8678,N_5601,N_7464);
nor U8679 (N_8679,N_5160,N_6977);
xnor U8680 (N_8680,N_5553,N_6563);
and U8681 (N_8681,N_6754,N_5239);
xor U8682 (N_8682,N_7002,N_6851);
nand U8683 (N_8683,N_6400,N_5465);
and U8684 (N_8684,N_6254,N_6214);
or U8685 (N_8685,N_5657,N_5478);
nor U8686 (N_8686,N_6586,N_7249);
nor U8687 (N_8687,N_6112,N_5495);
or U8688 (N_8688,N_5576,N_5186);
xor U8689 (N_8689,N_6578,N_7129);
nor U8690 (N_8690,N_7167,N_6088);
xor U8691 (N_8691,N_6828,N_6708);
nor U8692 (N_8692,N_6520,N_5781);
nor U8693 (N_8693,N_6682,N_5550);
nand U8694 (N_8694,N_6147,N_7298);
nor U8695 (N_8695,N_5078,N_7030);
and U8696 (N_8696,N_5572,N_5094);
nor U8697 (N_8697,N_6747,N_6454);
xnor U8698 (N_8698,N_6872,N_6934);
or U8699 (N_8699,N_5412,N_7367);
and U8700 (N_8700,N_6822,N_5329);
nor U8701 (N_8701,N_5809,N_6357);
xor U8702 (N_8702,N_6141,N_5622);
xnor U8703 (N_8703,N_7128,N_7282);
nand U8704 (N_8704,N_5958,N_6845);
xor U8705 (N_8705,N_6411,N_6373);
or U8706 (N_8706,N_6647,N_5920);
and U8707 (N_8707,N_5599,N_5377);
nor U8708 (N_8708,N_5892,N_7075);
nand U8709 (N_8709,N_6004,N_6639);
and U8710 (N_8710,N_7402,N_6093);
nand U8711 (N_8711,N_6240,N_5960);
xnor U8712 (N_8712,N_6809,N_5668);
or U8713 (N_8713,N_7126,N_5943);
and U8714 (N_8714,N_5415,N_7004);
xnor U8715 (N_8715,N_7445,N_7486);
or U8716 (N_8716,N_5751,N_7103);
nand U8717 (N_8717,N_6831,N_5084);
xor U8718 (N_8718,N_6861,N_7021);
xnor U8719 (N_8719,N_6633,N_7208);
nand U8720 (N_8720,N_6884,N_5018);
or U8721 (N_8721,N_5559,N_6504);
nand U8722 (N_8722,N_6646,N_6696);
or U8723 (N_8723,N_5215,N_5531);
or U8724 (N_8724,N_6073,N_6535);
or U8725 (N_8725,N_6010,N_6995);
nand U8726 (N_8726,N_5162,N_6862);
xnor U8727 (N_8727,N_5285,N_5427);
nand U8728 (N_8728,N_6904,N_7433);
xnor U8729 (N_8729,N_5310,N_6302);
or U8730 (N_8730,N_5592,N_6874);
nand U8731 (N_8731,N_6631,N_7454);
and U8732 (N_8732,N_5926,N_5922);
nor U8733 (N_8733,N_5065,N_6034);
xor U8734 (N_8734,N_6461,N_5910);
nand U8735 (N_8735,N_6767,N_6542);
nand U8736 (N_8736,N_6188,N_5211);
xnor U8737 (N_8737,N_6379,N_5863);
or U8738 (N_8738,N_6912,N_6236);
xnor U8739 (N_8739,N_5127,N_7165);
xor U8740 (N_8740,N_5462,N_6615);
nor U8741 (N_8741,N_6319,N_6189);
or U8742 (N_8742,N_6470,N_6660);
or U8743 (N_8743,N_5003,N_5144);
or U8744 (N_8744,N_6864,N_6228);
and U8745 (N_8745,N_5101,N_6467);
nand U8746 (N_8746,N_5536,N_5771);
nor U8747 (N_8747,N_5517,N_6450);
or U8748 (N_8748,N_7497,N_5345);
xor U8749 (N_8749,N_5371,N_5293);
nor U8750 (N_8750,N_6583,N_5037);
xnor U8751 (N_8751,N_6765,N_5252);
and U8752 (N_8752,N_5411,N_5842);
or U8753 (N_8753,N_5447,N_6060);
xnor U8754 (N_8754,N_5422,N_7095);
or U8755 (N_8755,N_5246,N_5014);
xnor U8756 (N_8756,N_6812,N_7213);
xnor U8757 (N_8757,N_5327,N_7262);
and U8758 (N_8758,N_5807,N_7098);
nand U8759 (N_8759,N_5330,N_6540);
nor U8760 (N_8760,N_5143,N_6357);
xnor U8761 (N_8761,N_5499,N_5483);
or U8762 (N_8762,N_6487,N_6245);
and U8763 (N_8763,N_5442,N_5512);
nand U8764 (N_8764,N_5865,N_5419);
or U8765 (N_8765,N_5834,N_5077);
and U8766 (N_8766,N_7483,N_5627);
xor U8767 (N_8767,N_6613,N_5608);
or U8768 (N_8768,N_5916,N_6241);
and U8769 (N_8769,N_6506,N_5110);
nor U8770 (N_8770,N_7469,N_6669);
xor U8771 (N_8771,N_7470,N_6662);
or U8772 (N_8772,N_5891,N_7289);
nand U8773 (N_8773,N_6682,N_7354);
nor U8774 (N_8774,N_6120,N_5267);
nor U8775 (N_8775,N_6204,N_6352);
xnor U8776 (N_8776,N_6872,N_6689);
xnor U8777 (N_8777,N_7366,N_6826);
or U8778 (N_8778,N_6823,N_6121);
nand U8779 (N_8779,N_6269,N_5647);
nand U8780 (N_8780,N_6320,N_7484);
nor U8781 (N_8781,N_5325,N_6166);
xor U8782 (N_8782,N_5347,N_6615);
nand U8783 (N_8783,N_6789,N_6423);
xnor U8784 (N_8784,N_5038,N_5386);
or U8785 (N_8785,N_5792,N_7388);
or U8786 (N_8786,N_5589,N_6556);
and U8787 (N_8787,N_5288,N_5716);
and U8788 (N_8788,N_7104,N_5377);
nand U8789 (N_8789,N_5567,N_6700);
and U8790 (N_8790,N_7399,N_7195);
or U8791 (N_8791,N_6786,N_6755);
and U8792 (N_8792,N_5473,N_5730);
or U8793 (N_8793,N_5788,N_5596);
and U8794 (N_8794,N_6977,N_5028);
nor U8795 (N_8795,N_7491,N_5016);
nor U8796 (N_8796,N_5375,N_7222);
nor U8797 (N_8797,N_6727,N_5854);
or U8798 (N_8798,N_5307,N_5394);
xor U8799 (N_8799,N_6297,N_5800);
or U8800 (N_8800,N_6616,N_6285);
nor U8801 (N_8801,N_7314,N_5802);
nand U8802 (N_8802,N_6577,N_5816);
nand U8803 (N_8803,N_7487,N_6038);
xor U8804 (N_8804,N_6998,N_5206);
xor U8805 (N_8805,N_6395,N_7359);
or U8806 (N_8806,N_5776,N_6372);
or U8807 (N_8807,N_6292,N_5678);
or U8808 (N_8808,N_6094,N_5754);
or U8809 (N_8809,N_5535,N_6850);
and U8810 (N_8810,N_5387,N_5105);
nor U8811 (N_8811,N_6829,N_5566);
nand U8812 (N_8812,N_6470,N_7467);
xor U8813 (N_8813,N_5337,N_6150);
xor U8814 (N_8814,N_6918,N_6874);
xnor U8815 (N_8815,N_5761,N_7326);
or U8816 (N_8816,N_5352,N_7396);
nor U8817 (N_8817,N_5152,N_5686);
xor U8818 (N_8818,N_5098,N_6363);
nand U8819 (N_8819,N_6384,N_6171);
and U8820 (N_8820,N_5321,N_5514);
nor U8821 (N_8821,N_6417,N_5935);
nor U8822 (N_8822,N_7148,N_6153);
nand U8823 (N_8823,N_7311,N_7482);
nor U8824 (N_8824,N_6008,N_6491);
xor U8825 (N_8825,N_6158,N_7387);
or U8826 (N_8826,N_7439,N_6660);
and U8827 (N_8827,N_7077,N_5696);
xnor U8828 (N_8828,N_6401,N_6095);
and U8829 (N_8829,N_5472,N_5482);
nor U8830 (N_8830,N_6944,N_5270);
xnor U8831 (N_8831,N_7222,N_6749);
nor U8832 (N_8832,N_7055,N_5834);
or U8833 (N_8833,N_7092,N_6229);
and U8834 (N_8834,N_6068,N_6978);
or U8835 (N_8835,N_6735,N_6550);
nor U8836 (N_8836,N_5215,N_6867);
xor U8837 (N_8837,N_6430,N_6937);
xnor U8838 (N_8838,N_7366,N_6171);
and U8839 (N_8839,N_6253,N_6989);
and U8840 (N_8840,N_6734,N_6589);
nor U8841 (N_8841,N_5488,N_5290);
nand U8842 (N_8842,N_5363,N_7493);
xor U8843 (N_8843,N_6662,N_7299);
nor U8844 (N_8844,N_6487,N_6589);
or U8845 (N_8845,N_5138,N_5007);
nand U8846 (N_8846,N_7445,N_5214);
xor U8847 (N_8847,N_6320,N_7141);
or U8848 (N_8848,N_6782,N_6200);
xor U8849 (N_8849,N_5744,N_6053);
nand U8850 (N_8850,N_7349,N_5999);
nand U8851 (N_8851,N_7407,N_7152);
or U8852 (N_8852,N_7467,N_5351);
xor U8853 (N_8853,N_6549,N_6387);
nor U8854 (N_8854,N_5629,N_6494);
nor U8855 (N_8855,N_6954,N_6168);
nor U8856 (N_8856,N_6110,N_5417);
nand U8857 (N_8857,N_7077,N_6932);
nand U8858 (N_8858,N_7266,N_7069);
or U8859 (N_8859,N_6146,N_5333);
xnor U8860 (N_8860,N_7126,N_6969);
xor U8861 (N_8861,N_5260,N_7498);
or U8862 (N_8862,N_5617,N_5769);
and U8863 (N_8863,N_6989,N_6567);
xnor U8864 (N_8864,N_5227,N_7275);
nand U8865 (N_8865,N_5147,N_5393);
nand U8866 (N_8866,N_7326,N_5095);
and U8867 (N_8867,N_6993,N_5059);
or U8868 (N_8868,N_6643,N_5629);
xnor U8869 (N_8869,N_5590,N_6390);
or U8870 (N_8870,N_7417,N_6182);
nand U8871 (N_8871,N_6576,N_5898);
nor U8872 (N_8872,N_6690,N_5639);
nand U8873 (N_8873,N_6732,N_5090);
xnor U8874 (N_8874,N_5822,N_6578);
or U8875 (N_8875,N_6898,N_5354);
nor U8876 (N_8876,N_5633,N_6944);
and U8877 (N_8877,N_5354,N_5098);
or U8878 (N_8878,N_5197,N_5154);
and U8879 (N_8879,N_6380,N_5818);
or U8880 (N_8880,N_5242,N_6296);
nand U8881 (N_8881,N_5133,N_5615);
or U8882 (N_8882,N_7382,N_5320);
nor U8883 (N_8883,N_5770,N_5358);
nand U8884 (N_8884,N_6307,N_6218);
nor U8885 (N_8885,N_6062,N_6131);
nand U8886 (N_8886,N_5324,N_6392);
xnor U8887 (N_8887,N_6882,N_6203);
nand U8888 (N_8888,N_5336,N_7162);
xnor U8889 (N_8889,N_7010,N_7138);
nand U8890 (N_8890,N_7362,N_5784);
and U8891 (N_8891,N_6518,N_5473);
and U8892 (N_8892,N_6980,N_5594);
nand U8893 (N_8893,N_5679,N_6731);
nand U8894 (N_8894,N_5158,N_6629);
nand U8895 (N_8895,N_7257,N_5554);
and U8896 (N_8896,N_6398,N_5240);
or U8897 (N_8897,N_5715,N_6464);
or U8898 (N_8898,N_5708,N_6441);
nor U8899 (N_8899,N_6252,N_6008);
and U8900 (N_8900,N_6721,N_6055);
or U8901 (N_8901,N_7345,N_6066);
nor U8902 (N_8902,N_6621,N_5833);
nand U8903 (N_8903,N_7401,N_6293);
and U8904 (N_8904,N_6013,N_5386);
nor U8905 (N_8905,N_6791,N_7062);
xnor U8906 (N_8906,N_6841,N_6453);
nand U8907 (N_8907,N_7418,N_7343);
and U8908 (N_8908,N_7250,N_6842);
nand U8909 (N_8909,N_7095,N_5877);
nor U8910 (N_8910,N_5188,N_6337);
or U8911 (N_8911,N_7384,N_5922);
or U8912 (N_8912,N_6533,N_5920);
xor U8913 (N_8913,N_6092,N_5324);
xnor U8914 (N_8914,N_7450,N_6323);
or U8915 (N_8915,N_6958,N_5781);
xnor U8916 (N_8916,N_5384,N_6786);
nor U8917 (N_8917,N_6189,N_6328);
xor U8918 (N_8918,N_5567,N_6883);
xor U8919 (N_8919,N_5541,N_5662);
and U8920 (N_8920,N_6356,N_7242);
or U8921 (N_8921,N_5636,N_7026);
or U8922 (N_8922,N_5523,N_6988);
and U8923 (N_8923,N_5223,N_5416);
xor U8924 (N_8924,N_6135,N_5222);
nor U8925 (N_8925,N_7144,N_6480);
xnor U8926 (N_8926,N_5985,N_7337);
or U8927 (N_8927,N_7202,N_7076);
and U8928 (N_8928,N_6738,N_6439);
and U8929 (N_8929,N_7202,N_5584);
nand U8930 (N_8930,N_6691,N_6563);
xor U8931 (N_8931,N_6227,N_6228);
xor U8932 (N_8932,N_7282,N_5552);
or U8933 (N_8933,N_5783,N_6531);
nor U8934 (N_8934,N_5403,N_5731);
and U8935 (N_8935,N_5824,N_6925);
and U8936 (N_8936,N_5985,N_5387);
xor U8937 (N_8937,N_7205,N_6857);
xor U8938 (N_8938,N_6619,N_5308);
or U8939 (N_8939,N_5060,N_5316);
xnor U8940 (N_8940,N_5814,N_6918);
and U8941 (N_8941,N_7330,N_5387);
and U8942 (N_8942,N_5876,N_5223);
or U8943 (N_8943,N_5347,N_7172);
nor U8944 (N_8944,N_6449,N_6914);
xnor U8945 (N_8945,N_7070,N_5748);
nor U8946 (N_8946,N_6239,N_7467);
xnor U8947 (N_8947,N_5129,N_5557);
nor U8948 (N_8948,N_5967,N_6004);
and U8949 (N_8949,N_7142,N_7182);
nand U8950 (N_8950,N_5969,N_7367);
nor U8951 (N_8951,N_6876,N_7336);
xor U8952 (N_8952,N_6181,N_7368);
xnor U8953 (N_8953,N_5767,N_5921);
nor U8954 (N_8954,N_5045,N_5947);
nand U8955 (N_8955,N_6596,N_6489);
or U8956 (N_8956,N_7087,N_7262);
xnor U8957 (N_8957,N_5391,N_5449);
nand U8958 (N_8958,N_5534,N_5329);
nor U8959 (N_8959,N_5100,N_5044);
xor U8960 (N_8960,N_5720,N_5565);
or U8961 (N_8961,N_5441,N_6888);
xnor U8962 (N_8962,N_5540,N_5308);
nor U8963 (N_8963,N_5614,N_6723);
and U8964 (N_8964,N_7092,N_6090);
or U8965 (N_8965,N_6021,N_6215);
xnor U8966 (N_8966,N_7480,N_6950);
and U8967 (N_8967,N_5463,N_6956);
and U8968 (N_8968,N_7179,N_5536);
or U8969 (N_8969,N_6854,N_7476);
or U8970 (N_8970,N_6221,N_5651);
nand U8971 (N_8971,N_7351,N_6236);
nor U8972 (N_8972,N_5348,N_6563);
nor U8973 (N_8973,N_6297,N_5640);
or U8974 (N_8974,N_5969,N_6040);
or U8975 (N_8975,N_6628,N_5766);
nand U8976 (N_8976,N_7202,N_7242);
or U8977 (N_8977,N_5052,N_5916);
or U8978 (N_8978,N_5745,N_5592);
nor U8979 (N_8979,N_5146,N_6584);
nand U8980 (N_8980,N_5073,N_6930);
or U8981 (N_8981,N_6699,N_5290);
nand U8982 (N_8982,N_6526,N_7487);
and U8983 (N_8983,N_6880,N_7459);
xnor U8984 (N_8984,N_6980,N_6109);
nor U8985 (N_8985,N_5361,N_7449);
nand U8986 (N_8986,N_5726,N_6570);
and U8987 (N_8987,N_6526,N_5957);
and U8988 (N_8988,N_5092,N_7190);
or U8989 (N_8989,N_5073,N_5891);
nand U8990 (N_8990,N_6973,N_6021);
nand U8991 (N_8991,N_6312,N_6883);
and U8992 (N_8992,N_5627,N_6787);
nand U8993 (N_8993,N_5779,N_5140);
or U8994 (N_8994,N_6313,N_6139);
and U8995 (N_8995,N_5851,N_5338);
nand U8996 (N_8996,N_5468,N_6850);
and U8997 (N_8997,N_5705,N_6909);
nor U8998 (N_8998,N_6025,N_7318);
or U8999 (N_8999,N_6279,N_6625);
xor U9000 (N_9000,N_5165,N_5377);
and U9001 (N_9001,N_6581,N_6143);
nor U9002 (N_9002,N_5093,N_6510);
and U9003 (N_9003,N_5577,N_7128);
nand U9004 (N_9004,N_6481,N_5274);
and U9005 (N_9005,N_5774,N_6519);
xor U9006 (N_9006,N_5726,N_6143);
xor U9007 (N_9007,N_5264,N_6608);
or U9008 (N_9008,N_5967,N_7236);
xor U9009 (N_9009,N_5568,N_5520);
xor U9010 (N_9010,N_6504,N_5319);
and U9011 (N_9011,N_6388,N_5134);
nand U9012 (N_9012,N_6087,N_6956);
xor U9013 (N_9013,N_6192,N_5983);
xnor U9014 (N_9014,N_5455,N_7377);
and U9015 (N_9015,N_5480,N_6440);
or U9016 (N_9016,N_6356,N_5964);
or U9017 (N_9017,N_5429,N_7475);
nand U9018 (N_9018,N_5103,N_5484);
and U9019 (N_9019,N_5048,N_5715);
xnor U9020 (N_9020,N_6263,N_7118);
or U9021 (N_9021,N_5410,N_6913);
nand U9022 (N_9022,N_6374,N_6711);
xnor U9023 (N_9023,N_5480,N_5372);
and U9024 (N_9024,N_6694,N_6348);
nor U9025 (N_9025,N_7111,N_7075);
or U9026 (N_9026,N_7173,N_7053);
nand U9027 (N_9027,N_6958,N_5996);
xor U9028 (N_9028,N_6596,N_5511);
and U9029 (N_9029,N_6416,N_6298);
nand U9030 (N_9030,N_5950,N_6042);
or U9031 (N_9031,N_5700,N_7181);
xor U9032 (N_9032,N_5816,N_5436);
nor U9033 (N_9033,N_6420,N_7424);
and U9034 (N_9034,N_7439,N_5185);
xor U9035 (N_9035,N_5449,N_5606);
nor U9036 (N_9036,N_7054,N_6560);
nand U9037 (N_9037,N_6860,N_5118);
or U9038 (N_9038,N_5377,N_5839);
nand U9039 (N_9039,N_7476,N_7206);
xor U9040 (N_9040,N_5436,N_5712);
nor U9041 (N_9041,N_5115,N_6583);
xnor U9042 (N_9042,N_7085,N_7003);
xnor U9043 (N_9043,N_5856,N_7241);
or U9044 (N_9044,N_6127,N_6848);
xnor U9045 (N_9045,N_5506,N_5416);
nor U9046 (N_9046,N_6864,N_5856);
and U9047 (N_9047,N_6335,N_5489);
or U9048 (N_9048,N_5393,N_5453);
and U9049 (N_9049,N_7196,N_6609);
or U9050 (N_9050,N_6640,N_7079);
xor U9051 (N_9051,N_5970,N_7152);
and U9052 (N_9052,N_5876,N_7204);
and U9053 (N_9053,N_6286,N_6648);
nor U9054 (N_9054,N_5501,N_6050);
nand U9055 (N_9055,N_5701,N_5625);
or U9056 (N_9056,N_5161,N_5737);
and U9057 (N_9057,N_7309,N_5587);
and U9058 (N_9058,N_5720,N_6247);
nor U9059 (N_9059,N_6632,N_6660);
xnor U9060 (N_9060,N_6044,N_5920);
or U9061 (N_9061,N_6435,N_6594);
nor U9062 (N_9062,N_7389,N_6802);
or U9063 (N_9063,N_6247,N_7494);
nor U9064 (N_9064,N_5168,N_6650);
and U9065 (N_9065,N_7044,N_5603);
nand U9066 (N_9066,N_5902,N_5549);
nand U9067 (N_9067,N_5772,N_6599);
xnor U9068 (N_9068,N_6993,N_6450);
nor U9069 (N_9069,N_5889,N_7339);
nand U9070 (N_9070,N_6330,N_5050);
nor U9071 (N_9071,N_7254,N_5702);
xnor U9072 (N_9072,N_7356,N_7201);
nor U9073 (N_9073,N_7068,N_7001);
nor U9074 (N_9074,N_6225,N_6123);
nor U9075 (N_9075,N_6571,N_7165);
and U9076 (N_9076,N_6790,N_6795);
and U9077 (N_9077,N_5627,N_6550);
nor U9078 (N_9078,N_6950,N_5854);
nor U9079 (N_9079,N_7057,N_5640);
and U9080 (N_9080,N_6070,N_5229);
or U9081 (N_9081,N_5801,N_5208);
xnor U9082 (N_9082,N_7348,N_7355);
nor U9083 (N_9083,N_5472,N_6641);
and U9084 (N_9084,N_5836,N_5790);
nor U9085 (N_9085,N_6044,N_5467);
nor U9086 (N_9086,N_5741,N_5745);
nand U9087 (N_9087,N_5321,N_5750);
xnor U9088 (N_9088,N_5404,N_7435);
or U9089 (N_9089,N_5004,N_7042);
and U9090 (N_9090,N_5884,N_6709);
xnor U9091 (N_9091,N_5568,N_6094);
and U9092 (N_9092,N_7262,N_5089);
nand U9093 (N_9093,N_6461,N_6582);
and U9094 (N_9094,N_5381,N_6667);
and U9095 (N_9095,N_6684,N_5372);
nor U9096 (N_9096,N_6197,N_6749);
xnor U9097 (N_9097,N_5022,N_6932);
nor U9098 (N_9098,N_6220,N_5977);
nand U9099 (N_9099,N_6107,N_6916);
or U9100 (N_9100,N_6708,N_5871);
nand U9101 (N_9101,N_6626,N_5433);
xnor U9102 (N_9102,N_5825,N_5539);
xor U9103 (N_9103,N_5558,N_6403);
nand U9104 (N_9104,N_5797,N_7246);
xnor U9105 (N_9105,N_7428,N_7429);
and U9106 (N_9106,N_5851,N_6712);
and U9107 (N_9107,N_7020,N_5757);
or U9108 (N_9108,N_6248,N_6729);
nand U9109 (N_9109,N_6785,N_5373);
nor U9110 (N_9110,N_6809,N_6519);
and U9111 (N_9111,N_6342,N_5133);
and U9112 (N_9112,N_5836,N_5515);
and U9113 (N_9113,N_6427,N_6597);
nand U9114 (N_9114,N_6219,N_6254);
xnor U9115 (N_9115,N_6616,N_6775);
or U9116 (N_9116,N_7070,N_7084);
and U9117 (N_9117,N_7186,N_5828);
or U9118 (N_9118,N_5061,N_6210);
nand U9119 (N_9119,N_7282,N_5675);
and U9120 (N_9120,N_5433,N_6537);
nor U9121 (N_9121,N_5629,N_5668);
xnor U9122 (N_9122,N_5659,N_5147);
or U9123 (N_9123,N_6153,N_6049);
and U9124 (N_9124,N_6242,N_6983);
nand U9125 (N_9125,N_6651,N_7441);
nor U9126 (N_9126,N_5960,N_5539);
or U9127 (N_9127,N_6753,N_5461);
nand U9128 (N_9128,N_5630,N_6123);
nor U9129 (N_9129,N_5492,N_7326);
or U9130 (N_9130,N_5502,N_6129);
nand U9131 (N_9131,N_5989,N_5839);
or U9132 (N_9132,N_6054,N_6889);
xnor U9133 (N_9133,N_6089,N_7297);
xor U9134 (N_9134,N_5669,N_5701);
nor U9135 (N_9135,N_7115,N_7407);
xor U9136 (N_9136,N_5799,N_6091);
and U9137 (N_9137,N_6194,N_6439);
and U9138 (N_9138,N_6505,N_7060);
nand U9139 (N_9139,N_5362,N_7184);
or U9140 (N_9140,N_6595,N_6559);
and U9141 (N_9141,N_7051,N_5770);
xor U9142 (N_9142,N_6451,N_5377);
nand U9143 (N_9143,N_7487,N_6660);
nor U9144 (N_9144,N_6994,N_7164);
nor U9145 (N_9145,N_6702,N_5163);
and U9146 (N_9146,N_6510,N_5366);
xnor U9147 (N_9147,N_7295,N_5104);
and U9148 (N_9148,N_5564,N_6984);
xnor U9149 (N_9149,N_6858,N_5462);
nor U9150 (N_9150,N_5891,N_6243);
nand U9151 (N_9151,N_7479,N_6556);
nor U9152 (N_9152,N_5212,N_5183);
xnor U9153 (N_9153,N_7039,N_5005);
nand U9154 (N_9154,N_5901,N_7371);
and U9155 (N_9155,N_6856,N_5075);
nor U9156 (N_9156,N_5156,N_6626);
nor U9157 (N_9157,N_5518,N_6047);
and U9158 (N_9158,N_5199,N_6068);
or U9159 (N_9159,N_7069,N_6700);
nor U9160 (N_9160,N_5146,N_6156);
xnor U9161 (N_9161,N_6592,N_5916);
nor U9162 (N_9162,N_6652,N_5709);
xnor U9163 (N_9163,N_6100,N_7106);
nor U9164 (N_9164,N_6505,N_7141);
and U9165 (N_9165,N_5088,N_6922);
nor U9166 (N_9166,N_6426,N_7216);
nand U9167 (N_9167,N_6164,N_6770);
or U9168 (N_9168,N_6992,N_7266);
nor U9169 (N_9169,N_7252,N_6962);
nor U9170 (N_9170,N_6898,N_6686);
or U9171 (N_9171,N_6670,N_6154);
nand U9172 (N_9172,N_6843,N_6321);
or U9173 (N_9173,N_5953,N_7357);
or U9174 (N_9174,N_5433,N_7235);
nand U9175 (N_9175,N_5277,N_5895);
and U9176 (N_9176,N_5497,N_5216);
nand U9177 (N_9177,N_6542,N_6481);
or U9178 (N_9178,N_5357,N_7336);
nor U9179 (N_9179,N_5749,N_6090);
nand U9180 (N_9180,N_7373,N_5261);
or U9181 (N_9181,N_6684,N_5787);
and U9182 (N_9182,N_6414,N_6227);
or U9183 (N_9183,N_6705,N_5059);
and U9184 (N_9184,N_5442,N_7095);
nor U9185 (N_9185,N_7017,N_5155);
nand U9186 (N_9186,N_6366,N_6554);
nor U9187 (N_9187,N_7139,N_5430);
and U9188 (N_9188,N_7227,N_7172);
and U9189 (N_9189,N_5285,N_5642);
nand U9190 (N_9190,N_5994,N_5073);
xnor U9191 (N_9191,N_6787,N_6992);
or U9192 (N_9192,N_5820,N_5396);
and U9193 (N_9193,N_5497,N_5372);
nand U9194 (N_9194,N_5581,N_7417);
nor U9195 (N_9195,N_5077,N_5995);
or U9196 (N_9196,N_7169,N_5023);
nor U9197 (N_9197,N_5325,N_7179);
nand U9198 (N_9198,N_5341,N_7054);
or U9199 (N_9199,N_5985,N_5307);
nor U9200 (N_9200,N_6395,N_6440);
or U9201 (N_9201,N_5087,N_5432);
or U9202 (N_9202,N_6766,N_7158);
nand U9203 (N_9203,N_7472,N_5432);
nor U9204 (N_9204,N_7314,N_6658);
xor U9205 (N_9205,N_7128,N_7054);
xor U9206 (N_9206,N_5176,N_6384);
nor U9207 (N_9207,N_6622,N_5327);
or U9208 (N_9208,N_6704,N_6859);
or U9209 (N_9209,N_7289,N_7276);
xnor U9210 (N_9210,N_7428,N_5950);
xnor U9211 (N_9211,N_6003,N_6060);
xor U9212 (N_9212,N_6375,N_5055);
and U9213 (N_9213,N_5740,N_5508);
nand U9214 (N_9214,N_6843,N_5741);
and U9215 (N_9215,N_5647,N_6841);
or U9216 (N_9216,N_5647,N_5589);
nand U9217 (N_9217,N_6043,N_7307);
and U9218 (N_9218,N_6816,N_6705);
and U9219 (N_9219,N_5821,N_5091);
nand U9220 (N_9220,N_6858,N_6376);
nor U9221 (N_9221,N_6885,N_6943);
or U9222 (N_9222,N_5644,N_6304);
nand U9223 (N_9223,N_5085,N_5707);
nand U9224 (N_9224,N_6713,N_5348);
and U9225 (N_9225,N_5968,N_5482);
nand U9226 (N_9226,N_6346,N_6520);
nand U9227 (N_9227,N_6468,N_6032);
nand U9228 (N_9228,N_5748,N_5859);
or U9229 (N_9229,N_7152,N_7119);
nand U9230 (N_9230,N_6122,N_5570);
or U9231 (N_9231,N_6598,N_5093);
and U9232 (N_9232,N_6671,N_5961);
or U9233 (N_9233,N_6461,N_7002);
nor U9234 (N_9234,N_5460,N_7229);
xor U9235 (N_9235,N_6403,N_6816);
and U9236 (N_9236,N_5395,N_6781);
nor U9237 (N_9237,N_6875,N_5614);
or U9238 (N_9238,N_5912,N_6597);
nor U9239 (N_9239,N_6409,N_7262);
or U9240 (N_9240,N_6916,N_5825);
and U9241 (N_9241,N_6723,N_6170);
and U9242 (N_9242,N_5964,N_6166);
and U9243 (N_9243,N_6834,N_7187);
nand U9244 (N_9244,N_6236,N_5130);
or U9245 (N_9245,N_7353,N_6992);
nand U9246 (N_9246,N_5159,N_5640);
and U9247 (N_9247,N_6099,N_5476);
nand U9248 (N_9248,N_5010,N_5016);
and U9249 (N_9249,N_5370,N_5977);
and U9250 (N_9250,N_6775,N_5830);
nand U9251 (N_9251,N_5627,N_5019);
or U9252 (N_9252,N_5939,N_5623);
nand U9253 (N_9253,N_6713,N_5769);
and U9254 (N_9254,N_6641,N_5899);
and U9255 (N_9255,N_5321,N_5220);
nand U9256 (N_9256,N_5875,N_5184);
and U9257 (N_9257,N_6556,N_7163);
xor U9258 (N_9258,N_5462,N_6969);
nor U9259 (N_9259,N_7209,N_5511);
or U9260 (N_9260,N_6360,N_6830);
nand U9261 (N_9261,N_5010,N_6397);
nor U9262 (N_9262,N_5252,N_7252);
nor U9263 (N_9263,N_7400,N_6539);
nor U9264 (N_9264,N_6242,N_5500);
nand U9265 (N_9265,N_6623,N_7147);
or U9266 (N_9266,N_5285,N_7404);
nand U9267 (N_9267,N_5170,N_5222);
or U9268 (N_9268,N_6291,N_6223);
nand U9269 (N_9269,N_5325,N_5323);
xor U9270 (N_9270,N_6285,N_7129);
and U9271 (N_9271,N_6063,N_5156);
nor U9272 (N_9272,N_7044,N_6341);
nand U9273 (N_9273,N_6459,N_5502);
or U9274 (N_9274,N_7266,N_6022);
nor U9275 (N_9275,N_7248,N_5692);
nand U9276 (N_9276,N_7279,N_6520);
or U9277 (N_9277,N_6518,N_6776);
and U9278 (N_9278,N_5777,N_5562);
nand U9279 (N_9279,N_6809,N_6172);
xor U9280 (N_9280,N_7194,N_6187);
and U9281 (N_9281,N_7378,N_6955);
nand U9282 (N_9282,N_6634,N_7211);
nor U9283 (N_9283,N_5894,N_5309);
and U9284 (N_9284,N_6202,N_5508);
or U9285 (N_9285,N_7099,N_6620);
and U9286 (N_9286,N_6307,N_7432);
nand U9287 (N_9287,N_5654,N_5116);
and U9288 (N_9288,N_5749,N_5999);
and U9289 (N_9289,N_6774,N_7026);
or U9290 (N_9290,N_5190,N_6609);
nor U9291 (N_9291,N_7245,N_5793);
nand U9292 (N_9292,N_6817,N_6115);
and U9293 (N_9293,N_5085,N_5773);
nand U9294 (N_9294,N_6150,N_6099);
nand U9295 (N_9295,N_7179,N_5510);
nand U9296 (N_9296,N_6862,N_5944);
xor U9297 (N_9297,N_6540,N_6135);
and U9298 (N_9298,N_5494,N_5448);
nor U9299 (N_9299,N_5562,N_7048);
and U9300 (N_9300,N_6960,N_5195);
xor U9301 (N_9301,N_7202,N_7491);
nand U9302 (N_9302,N_6962,N_5172);
and U9303 (N_9303,N_5367,N_5201);
nor U9304 (N_9304,N_5918,N_6228);
nand U9305 (N_9305,N_7489,N_6285);
nor U9306 (N_9306,N_5858,N_5663);
nor U9307 (N_9307,N_5215,N_7374);
or U9308 (N_9308,N_5682,N_6336);
nor U9309 (N_9309,N_5552,N_6478);
or U9310 (N_9310,N_5940,N_6269);
or U9311 (N_9311,N_7088,N_7136);
and U9312 (N_9312,N_5114,N_6648);
xor U9313 (N_9313,N_5060,N_7107);
and U9314 (N_9314,N_5079,N_6908);
nor U9315 (N_9315,N_6735,N_5581);
xor U9316 (N_9316,N_5568,N_6254);
or U9317 (N_9317,N_5182,N_6881);
nand U9318 (N_9318,N_6234,N_6683);
nor U9319 (N_9319,N_5667,N_6701);
nor U9320 (N_9320,N_7114,N_6299);
and U9321 (N_9321,N_5223,N_5279);
xnor U9322 (N_9322,N_5855,N_5972);
or U9323 (N_9323,N_7118,N_7435);
nand U9324 (N_9324,N_5144,N_7010);
xnor U9325 (N_9325,N_7109,N_5303);
nand U9326 (N_9326,N_6383,N_7079);
xor U9327 (N_9327,N_6620,N_7264);
xnor U9328 (N_9328,N_5263,N_5057);
nand U9329 (N_9329,N_6628,N_6358);
nand U9330 (N_9330,N_7259,N_5988);
and U9331 (N_9331,N_5994,N_7192);
nor U9332 (N_9332,N_6650,N_6415);
nor U9333 (N_9333,N_6464,N_6377);
and U9334 (N_9334,N_5432,N_6230);
xnor U9335 (N_9335,N_7258,N_6047);
nand U9336 (N_9336,N_6626,N_7087);
nor U9337 (N_9337,N_6443,N_5766);
and U9338 (N_9338,N_6657,N_5025);
nand U9339 (N_9339,N_7327,N_5672);
and U9340 (N_9340,N_5557,N_5152);
nor U9341 (N_9341,N_7212,N_5856);
and U9342 (N_9342,N_5744,N_7230);
nand U9343 (N_9343,N_5412,N_6340);
and U9344 (N_9344,N_5976,N_6410);
nor U9345 (N_9345,N_5341,N_6382);
nor U9346 (N_9346,N_6442,N_5907);
or U9347 (N_9347,N_6869,N_6984);
and U9348 (N_9348,N_7170,N_6900);
or U9349 (N_9349,N_5203,N_7368);
or U9350 (N_9350,N_6954,N_5851);
xnor U9351 (N_9351,N_7466,N_7080);
nor U9352 (N_9352,N_5622,N_7061);
nor U9353 (N_9353,N_5596,N_6115);
nand U9354 (N_9354,N_7354,N_6250);
xor U9355 (N_9355,N_6509,N_6663);
or U9356 (N_9356,N_6524,N_6668);
and U9357 (N_9357,N_5424,N_5559);
and U9358 (N_9358,N_7078,N_7262);
nand U9359 (N_9359,N_5280,N_7266);
and U9360 (N_9360,N_5749,N_5312);
nor U9361 (N_9361,N_5371,N_5707);
or U9362 (N_9362,N_5448,N_5903);
nor U9363 (N_9363,N_7187,N_6575);
nand U9364 (N_9364,N_5705,N_7012);
xnor U9365 (N_9365,N_5933,N_7057);
xor U9366 (N_9366,N_5731,N_6157);
or U9367 (N_9367,N_5884,N_6959);
and U9368 (N_9368,N_6149,N_5219);
and U9369 (N_9369,N_6117,N_5779);
and U9370 (N_9370,N_6658,N_6816);
nand U9371 (N_9371,N_6320,N_7248);
xor U9372 (N_9372,N_7417,N_6148);
nor U9373 (N_9373,N_6321,N_6448);
and U9374 (N_9374,N_5548,N_6913);
nand U9375 (N_9375,N_5677,N_5724);
and U9376 (N_9376,N_7293,N_6968);
xnor U9377 (N_9377,N_5264,N_6503);
and U9378 (N_9378,N_5428,N_5764);
and U9379 (N_9379,N_6070,N_7070);
and U9380 (N_9380,N_6679,N_6304);
xnor U9381 (N_9381,N_6961,N_5716);
xor U9382 (N_9382,N_6326,N_7423);
xnor U9383 (N_9383,N_5857,N_5852);
nor U9384 (N_9384,N_7104,N_7243);
or U9385 (N_9385,N_7017,N_7452);
or U9386 (N_9386,N_5861,N_6222);
and U9387 (N_9387,N_7401,N_5235);
nand U9388 (N_9388,N_7257,N_7206);
nand U9389 (N_9389,N_7140,N_6623);
nor U9390 (N_9390,N_6798,N_6069);
nand U9391 (N_9391,N_5901,N_5511);
or U9392 (N_9392,N_5591,N_5905);
nand U9393 (N_9393,N_6957,N_6034);
or U9394 (N_9394,N_6787,N_7314);
or U9395 (N_9395,N_5526,N_6397);
nor U9396 (N_9396,N_6968,N_6031);
nor U9397 (N_9397,N_5622,N_6358);
and U9398 (N_9398,N_5454,N_6291);
and U9399 (N_9399,N_7060,N_6867);
or U9400 (N_9400,N_6443,N_7233);
xnor U9401 (N_9401,N_5273,N_6463);
and U9402 (N_9402,N_6408,N_5766);
xor U9403 (N_9403,N_7399,N_5235);
or U9404 (N_9404,N_6805,N_7038);
nor U9405 (N_9405,N_7292,N_6697);
and U9406 (N_9406,N_7180,N_5655);
xor U9407 (N_9407,N_6795,N_6417);
or U9408 (N_9408,N_5727,N_6111);
nand U9409 (N_9409,N_5485,N_7441);
or U9410 (N_9410,N_7004,N_6201);
xor U9411 (N_9411,N_6869,N_5838);
xor U9412 (N_9412,N_5480,N_6741);
nand U9413 (N_9413,N_5134,N_6055);
and U9414 (N_9414,N_7435,N_5115);
xnor U9415 (N_9415,N_7214,N_7097);
and U9416 (N_9416,N_7351,N_6633);
or U9417 (N_9417,N_7356,N_6830);
or U9418 (N_9418,N_6141,N_5540);
and U9419 (N_9419,N_5137,N_6643);
nand U9420 (N_9420,N_6680,N_6965);
nand U9421 (N_9421,N_5067,N_6960);
and U9422 (N_9422,N_5871,N_7036);
or U9423 (N_9423,N_5257,N_6328);
or U9424 (N_9424,N_5057,N_6987);
or U9425 (N_9425,N_5854,N_6384);
and U9426 (N_9426,N_5270,N_7391);
nand U9427 (N_9427,N_5934,N_5436);
or U9428 (N_9428,N_6404,N_6435);
xor U9429 (N_9429,N_5901,N_6749);
nand U9430 (N_9430,N_5125,N_5939);
or U9431 (N_9431,N_5817,N_7119);
xor U9432 (N_9432,N_6932,N_6971);
xor U9433 (N_9433,N_6216,N_7399);
or U9434 (N_9434,N_7292,N_6346);
nor U9435 (N_9435,N_6285,N_5388);
nor U9436 (N_9436,N_5121,N_6261);
nand U9437 (N_9437,N_5334,N_6601);
xor U9438 (N_9438,N_7292,N_6140);
and U9439 (N_9439,N_5075,N_5467);
and U9440 (N_9440,N_5932,N_7439);
nand U9441 (N_9441,N_5240,N_7060);
and U9442 (N_9442,N_6151,N_5382);
xnor U9443 (N_9443,N_5407,N_7236);
nor U9444 (N_9444,N_5531,N_6049);
nand U9445 (N_9445,N_6088,N_6721);
and U9446 (N_9446,N_5707,N_7268);
xnor U9447 (N_9447,N_6099,N_5204);
nor U9448 (N_9448,N_5420,N_6196);
nand U9449 (N_9449,N_5840,N_6618);
xor U9450 (N_9450,N_5778,N_5506);
xor U9451 (N_9451,N_6120,N_5572);
and U9452 (N_9452,N_5773,N_5025);
and U9453 (N_9453,N_7105,N_5074);
xnor U9454 (N_9454,N_5638,N_7357);
xor U9455 (N_9455,N_6600,N_6006);
and U9456 (N_9456,N_5238,N_6867);
xnor U9457 (N_9457,N_6137,N_6247);
nand U9458 (N_9458,N_5375,N_5379);
and U9459 (N_9459,N_6021,N_5976);
and U9460 (N_9460,N_5368,N_5042);
nand U9461 (N_9461,N_6352,N_6525);
and U9462 (N_9462,N_5614,N_5641);
nand U9463 (N_9463,N_7046,N_6486);
nand U9464 (N_9464,N_6038,N_6254);
and U9465 (N_9465,N_5483,N_5306);
nand U9466 (N_9466,N_5761,N_5493);
nand U9467 (N_9467,N_5671,N_5283);
and U9468 (N_9468,N_6550,N_6325);
nor U9469 (N_9469,N_5625,N_5165);
nand U9470 (N_9470,N_5991,N_6875);
and U9471 (N_9471,N_5342,N_6373);
xnor U9472 (N_9472,N_6919,N_5358);
or U9473 (N_9473,N_5824,N_6930);
and U9474 (N_9474,N_7004,N_7136);
xnor U9475 (N_9475,N_6209,N_6679);
or U9476 (N_9476,N_6831,N_6725);
and U9477 (N_9477,N_6075,N_5102);
and U9478 (N_9478,N_6479,N_5495);
xor U9479 (N_9479,N_5500,N_7129);
nand U9480 (N_9480,N_7461,N_6286);
or U9481 (N_9481,N_5156,N_5253);
nor U9482 (N_9482,N_5103,N_6317);
or U9483 (N_9483,N_7417,N_6277);
nor U9484 (N_9484,N_7438,N_6968);
and U9485 (N_9485,N_7415,N_5948);
xnor U9486 (N_9486,N_5097,N_6109);
or U9487 (N_9487,N_6212,N_6766);
or U9488 (N_9488,N_5915,N_6209);
nor U9489 (N_9489,N_6989,N_6730);
nor U9490 (N_9490,N_6595,N_6215);
or U9491 (N_9491,N_5884,N_7039);
nor U9492 (N_9492,N_7050,N_7212);
and U9493 (N_9493,N_5487,N_5533);
or U9494 (N_9494,N_5591,N_7380);
nor U9495 (N_9495,N_5577,N_7452);
nor U9496 (N_9496,N_7080,N_5489);
xnor U9497 (N_9497,N_7361,N_6022);
xnor U9498 (N_9498,N_5726,N_6118);
nand U9499 (N_9499,N_5816,N_6448);
or U9500 (N_9500,N_5643,N_6605);
nand U9501 (N_9501,N_6986,N_5472);
and U9502 (N_9502,N_7063,N_7213);
xnor U9503 (N_9503,N_7149,N_7010);
or U9504 (N_9504,N_6105,N_5477);
or U9505 (N_9505,N_5717,N_5651);
and U9506 (N_9506,N_6374,N_5044);
xnor U9507 (N_9507,N_7405,N_6000);
or U9508 (N_9508,N_7168,N_6737);
nor U9509 (N_9509,N_5417,N_7233);
nor U9510 (N_9510,N_6775,N_5071);
and U9511 (N_9511,N_6459,N_6794);
xor U9512 (N_9512,N_5640,N_5487);
xnor U9513 (N_9513,N_7055,N_5833);
and U9514 (N_9514,N_6439,N_7242);
nor U9515 (N_9515,N_6175,N_6664);
or U9516 (N_9516,N_6520,N_6415);
nand U9517 (N_9517,N_6243,N_5494);
xnor U9518 (N_9518,N_6839,N_7013);
or U9519 (N_9519,N_6130,N_6472);
nor U9520 (N_9520,N_7088,N_6371);
or U9521 (N_9521,N_6774,N_6260);
xnor U9522 (N_9522,N_6323,N_5399);
xnor U9523 (N_9523,N_7237,N_5549);
nor U9524 (N_9524,N_7359,N_5694);
and U9525 (N_9525,N_6909,N_6505);
xor U9526 (N_9526,N_7324,N_5342);
or U9527 (N_9527,N_6288,N_6916);
and U9528 (N_9528,N_6760,N_6461);
xnor U9529 (N_9529,N_6844,N_6980);
xnor U9530 (N_9530,N_6067,N_5948);
nand U9531 (N_9531,N_6089,N_6917);
or U9532 (N_9532,N_6533,N_6778);
nor U9533 (N_9533,N_5772,N_5295);
xnor U9534 (N_9534,N_6693,N_5689);
or U9535 (N_9535,N_6031,N_6159);
nand U9536 (N_9536,N_5990,N_7079);
or U9537 (N_9537,N_7315,N_5506);
nand U9538 (N_9538,N_7073,N_5884);
nand U9539 (N_9539,N_6926,N_5254);
nand U9540 (N_9540,N_6670,N_7394);
xnor U9541 (N_9541,N_7336,N_6728);
or U9542 (N_9542,N_5104,N_5914);
or U9543 (N_9543,N_5962,N_6942);
nor U9544 (N_9544,N_7322,N_6460);
nand U9545 (N_9545,N_5304,N_6480);
xor U9546 (N_9546,N_7178,N_5140);
or U9547 (N_9547,N_6922,N_7399);
or U9548 (N_9548,N_6466,N_5579);
or U9549 (N_9549,N_6019,N_6920);
nand U9550 (N_9550,N_6289,N_6015);
nor U9551 (N_9551,N_6926,N_5968);
and U9552 (N_9552,N_6788,N_5480);
xor U9553 (N_9553,N_6008,N_6633);
xor U9554 (N_9554,N_6278,N_5805);
nand U9555 (N_9555,N_7423,N_6614);
xnor U9556 (N_9556,N_6541,N_5805);
nand U9557 (N_9557,N_7338,N_5987);
or U9558 (N_9558,N_6108,N_6876);
or U9559 (N_9559,N_5403,N_5280);
nor U9560 (N_9560,N_6997,N_5666);
and U9561 (N_9561,N_5195,N_5656);
nand U9562 (N_9562,N_5295,N_6590);
xor U9563 (N_9563,N_5451,N_6701);
nor U9564 (N_9564,N_5328,N_6293);
or U9565 (N_9565,N_6514,N_5950);
or U9566 (N_9566,N_7467,N_5092);
nor U9567 (N_9567,N_6694,N_6182);
nand U9568 (N_9568,N_5852,N_7273);
and U9569 (N_9569,N_5151,N_5167);
nand U9570 (N_9570,N_6298,N_5205);
xor U9571 (N_9571,N_5130,N_7475);
or U9572 (N_9572,N_6339,N_5423);
nor U9573 (N_9573,N_5981,N_7446);
and U9574 (N_9574,N_7055,N_6195);
nor U9575 (N_9575,N_6528,N_7305);
nor U9576 (N_9576,N_5663,N_6376);
or U9577 (N_9577,N_5376,N_6689);
and U9578 (N_9578,N_5011,N_6049);
nor U9579 (N_9579,N_5370,N_6390);
nand U9580 (N_9580,N_7413,N_7481);
and U9581 (N_9581,N_6180,N_6019);
or U9582 (N_9582,N_7475,N_5071);
and U9583 (N_9583,N_7357,N_5843);
and U9584 (N_9584,N_7479,N_6885);
xor U9585 (N_9585,N_5590,N_6383);
xor U9586 (N_9586,N_5730,N_6608);
nor U9587 (N_9587,N_5689,N_6594);
nor U9588 (N_9588,N_5176,N_7309);
nor U9589 (N_9589,N_6402,N_5884);
nor U9590 (N_9590,N_5873,N_5769);
or U9591 (N_9591,N_5881,N_5297);
xor U9592 (N_9592,N_5940,N_6970);
and U9593 (N_9593,N_6709,N_7267);
nand U9594 (N_9594,N_6516,N_6246);
and U9595 (N_9595,N_5556,N_5726);
or U9596 (N_9596,N_7262,N_6960);
nand U9597 (N_9597,N_7151,N_7032);
nand U9598 (N_9598,N_5705,N_6562);
and U9599 (N_9599,N_5272,N_5872);
nor U9600 (N_9600,N_6524,N_5361);
nand U9601 (N_9601,N_6277,N_7213);
xor U9602 (N_9602,N_5670,N_7483);
or U9603 (N_9603,N_7247,N_6433);
or U9604 (N_9604,N_5268,N_6636);
nand U9605 (N_9605,N_5648,N_5201);
xor U9606 (N_9606,N_6147,N_6510);
or U9607 (N_9607,N_5737,N_6044);
xor U9608 (N_9608,N_7240,N_7126);
or U9609 (N_9609,N_5296,N_7159);
nor U9610 (N_9610,N_7496,N_7381);
and U9611 (N_9611,N_5199,N_6115);
nand U9612 (N_9612,N_5092,N_5223);
or U9613 (N_9613,N_7063,N_5568);
nor U9614 (N_9614,N_5887,N_5300);
xor U9615 (N_9615,N_6228,N_5730);
and U9616 (N_9616,N_6109,N_5127);
nor U9617 (N_9617,N_7477,N_5551);
or U9618 (N_9618,N_6811,N_6826);
nor U9619 (N_9619,N_7233,N_6321);
xor U9620 (N_9620,N_6552,N_7061);
or U9621 (N_9621,N_6722,N_5918);
and U9622 (N_9622,N_5584,N_5469);
and U9623 (N_9623,N_5445,N_6984);
and U9624 (N_9624,N_7054,N_5021);
xnor U9625 (N_9625,N_5635,N_5956);
or U9626 (N_9626,N_5149,N_5394);
or U9627 (N_9627,N_6306,N_6959);
xnor U9628 (N_9628,N_7461,N_5324);
nor U9629 (N_9629,N_7009,N_6001);
nor U9630 (N_9630,N_7091,N_6044);
nand U9631 (N_9631,N_5735,N_6574);
or U9632 (N_9632,N_5167,N_5795);
xnor U9633 (N_9633,N_6926,N_7294);
and U9634 (N_9634,N_6007,N_5273);
and U9635 (N_9635,N_6372,N_5964);
xor U9636 (N_9636,N_7465,N_6423);
nor U9637 (N_9637,N_6739,N_5865);
or U9638 (N_9638,N_5432,N_7414);
nand U9639 (N_9639,N_6464,N_6926);
and U9640 (N_9640,N_6347,N_6950);
or U9641 (N_9641,N_6415,N_5334);
xnor U9642 (N_9642,N_5021,N_5412);
and U9643 (N_9643,N_5830,N_7256);
or U9644 (N_9644,N_6218,N_6174);
xnor U9645 (N_9645,N_6742,N_6534);
nand U9646 (N_9646,N_6085,N_5451);
and U9647 (N_9647,N_6525,N_6446);
or U9648 (N_9648,N_6751,N_6357);
and U9649 (N_9649,N_5081,N_5391);
xor U9650 (N_9650,N_5718,N_5280);
and U9651 (N_9651,N_5725,N_5218);
xor U9652 (N_9652,N_6513,N_7357);
xnor U9653 (N_9653,N_6081,N_6619);
nor U9654 (N_9654,N_7420,N_5479);
and U9655 (N_9655,N_6546,N_7157);
or U9656 (N_9656,N_7434,N_7308);
nand U9657 (N_9657,N_5471,N_7421);
xor U9658 (N_9658,N_5713,N_6364);
nand U9659 (N_9659,N_6703,N_7277);
nand U9660 (N_9660,N_5546,N_5336);
xor U9661 (N_9661,N_6845,N_6998);
or U9662 (N_9662,N_5315,N_6099);
nand U9663 (N_9663,N_5743,N_7173);
nor U9664 (N_9664,N_7081,N_7180);
nor U9665 (N_9665,N_6294,N_6369);
and U9666 (N_9666,N_6422,N_7438);
or U9667 (N_9667,N_6948,N_6181);
nor U9668 (N_9668,N_7195,N_7177);
nand U9669 (N_9669,N_7179,N_6504);
nand U9670 (N_9670,N_5434,N_7218);
xnor U9671 (N_9671,N_7426,N_7351);
or U9672 (N_9672,N_5037,N_6312);
and U9673 (N_9673,N_6465,N_5831);
nor U9674 (N_9674,N_5829,N_6698);
and U9675 (N_9675,N_5874,N_5680);
and U9676 (N_9676,N_6621,N_7414);
and U9677 (N_9677,N_5590,N_6204);
nor U9678 (N_9678,N_5694,N_6059);
xnor U9679 (N_9679,N_5932,N_7087);
or U9680 (N_9680,N_6150,N_5083);
and U9681 (N_9681,N_6430,N_5650);
xor U9682 (N_9682,N_7386,N_6432);
nand U9683 (N_9683,N_7349,N_5306);
nand U9684 (N_9684,N_7121,N_6387);
xnor U9685 (N_9685,N_5284,N_7159);
or U9686 (N_9686,N_5457,N_6379);
or U9687 (N_9687,N_5638,N_6559);
and U9688 (N_9688,N_6720,N_7196);
or U9689 (N_9689,N_5748,N_6664);
nor U9690 (N_9690,N_5724,N_6397);
and U9691 (N_9691,N_6364,N_5602);
nand U9692 (N_9692,N_6333,N_7144);
or U9693 (N_9693,N_5181,N_5483);
nand U9694 (N_9694,N_6699,N_5319);
nor U9695 (N_9695,N_6204,N_6752);
nor U9696 (N_9696,N_5498,N_7487);
or U9697 (N_9697,N_5285,N_5517);
or U9698 (N_9698,N_5540,N_6652);
and U9699 (N_9699,N_6976,N_7202);
and U9700 (N_9700,N_5778,N_6435);
or U9701 (N_9701,N_6020,N_6328);
nor U9702 (N_9702,N_6615,N_6360);
nand U9703 (N_9703,N_6617,N_6118);
nor U9704 (N_9704,N_6071,N_6316);
nor U9705 (N_9705,N_5904,N_6836);
and U9706 (N_9706,N_7472,N_6655);
nand U9707 (N_9707,N_6650,N_6812);
nor U9708 (N_9708,N_6140,N_5095);
nor U9709 (N_9709,N_7314,N_6372);
and U9710 (N_9710,N_5087,N_6153);
nor U9711 (N_9711,N_7077,N_6488);
and U9712 (N_9712,N_6699,N_6375);
xor U9713 (N_9713,N_6065,N_5050);
and U9714 (N_9714,N_5481,N_5560);
or U9715 (N_9715,N_7077,N_6274);
nor U9716 (N_9716,N_6716,N_5043);
and U9717 (N_9717,N_7008,N_5445);
nand U9718 (N_9718,N_6989,N_7240);
nor U9719 (N_9719,N_5116,N_7487);
or U9720 (N_9720,N_5812,N_6461);
nor U9721 (N_9721,N_5506,N_6173);
and U9722 (N_9722,N_5241,N_7319);
and U9723 (N_9723,N_6113,N_7082);
xnor U9724 (N_9724,N_5012,N_5315);
nor U9725 (N_9725,N_5168,N_5726);
and U9726 (N_9726,N_5363,N_5190);
and U9727 (N_9727,N_5596,N_6538);
nand U9728 (N_9728,N_5327,N_6343);
and U9729 (N_9729,N_5228,N_5986);
and U9730 (N_9730,N_7073,N_7152);
nor U9731 (N_9731,N_6903,N_7487);
or U9732 (N_9732,N_7388,N_7267);
or U9733 (N_9733,N_5373,N_7271);
xor U9734 (N_9734,N_7084,N_6118);
nand U9735 (N_9735,N_5093,N_7288);
nand U9736 (N_9736,N_5753,N_6736);
xor U9737 (N_9737,N_7302,N_6331);
xnor U9738 (N_9738,N_6120,N_7411);
and U9739 (N_9739,N_6662,N_7453);
xnor U9740 (N_9740,N_5004,N_5184);
nor U9741 (N_9741,N_6539,N_6900);
xnor U9742 (N_9742,N_7035,N_6156);
nor U9743 (N_9743,N_6577,N_7451);
nor U9744 (N_9744,N_6118,N_7237);
xor U9745 (N_9745,N_7347,N_6505);
nor U9746 (N_9746,N_5052,N_6787);
xor U9747 (N_9747,N_6393,N_5963);
nand U9748 (N_9748,N_7467,N_5710);
and U9749 (N_9749,N_7427,N_7464);
xor U9750 (N_9750,N_6991,N_5190);
nand U9751 (N_9751,N_7476,N_6375);
and U9752 (N_9752,N_7206,N_6599);
and U9753 (N_9753,N_7402,N_6992);
xor U9754 (N_9754,N_6839,N_6821);
xor U9755 (N_9755,N_6825,N_5906);
xnor U9756 (N_9756,N_7125,N_6923);
xnor U9757 (N_9757,N_5836,N_5163);
nor U9758 (N_9758,N_5574,N_5989);
nand U9759 (N_9759,N_6717,N_6696);
xnor U9760 (N_9760,N_6757,N_6093);
or U9761 (N_9761,N_6446,N_6628);
nor U9762 (N_9762,N_5165,N_5792);
xnor U9763 (N_9763,N_6391,N_7060);
and U9764 (N_9764,N_5151,N_5866);
nand U9765 (N_9765,N_5620,N_7326);
nor U9766 (N_9766,N_5469,N_6823);
xor U9767 (N_9767,N_5627,N_5961);
or U9768 (N_9768,N_6106,N_6226);
nor U9769 (N_9769,N_7335,N_7461);
xnor U9770 (N_9770,N_6725,N_6796);
and U9771 (N_9771,N_6580,N_6196);
nor U9772 (N_9772,N_6214,N_5838);
or U9773 (N_9773,N_5754,N_5019);
nor U9774 (N_9774,N_6473,N_5380);
and U9775 (N_9775,N_6630,N_5377);
and U9776 (N_9776,N_5468,N_5935);
nand U9777 (N_9777,N_7418,N_5358);
nor U9778 (N_9778,N_6780,N_6965);
and U9779 (N_9779,N_7223,N_5123);
xnor U9780 (N_9780,N_7301,N_5062);
nand U9781 (N_9781,N_7091,N_5264);
nor U9782 (N_9782,N_5445,N_7449);
nand U9783 (N_9783,N_7158,N_5751);
or U9784 (N_9784,N_5494,N_7451);
or U9785 (N_9785,N_5944,N_5515);
nand U9786 (N_9786,N_6121,N_7409);
nand U9787 (N_9787,N_5203,N_5132);
xnor U9788 (N_9788,N_5084,N_6415);
nand U9789 (N_9789,N_7148,N_5701);
or U9790 (N_9790,N_5091,N_5362);
nand U9791 (N_9791,N_6566,N_5464);
or U9792 (N_9792,N_7038,N_6595);
nand U9793 (N_9793,N_5248,N_5806);
nand U9794 (N_9794,N_6733,N_7238);
nand U9795 (N_9795,N_5507,N_7167);
xnor U9796 (N_9796,N_5812,N_6447);
nand U9797 (N_9797,N_5481,N_5313);
nor U9798 (N_9798,N_7384,N_7449);
and U9799 (N_9799,N_7468,N_7156);
nand U9800 (N_9800,N_5179,N_6468);
nand U9801 (N_9801,N_5738,N_5876);
xor U9802 (N_9802,N_7069,N_5789);
and U9803 (N_9803,N_7127,N_6168);
nor U9804 (N_9804,N_7433,N_6684);
xor U9805 (N_9805,N_7406,N_6396);
or U9806 (N_9806,N_6084,N_5171);
or U9807 (N_9807,N_6735,N_5405);
or U9808 (N_9808,N_7340,N_6968);
nand U9809 (N_9809,N_7360,N_6431);
nor U9810 (N_9810,N_7251,N_7370);
nor U9811 (N_9811,N_5990,N_5932);
nor U9812 (N_9812,N_5405,N_6932);
and U9813 (N_9813,N_5638,N_5894);
and U9814 (N_9814,N_7030,N_5631);
and U9815 (N_9815,N_6041,N_7462);
nand U9816 (N_9816,N_6903,N_5988);
nand U9817 (N_9817,N_6042,N_6603);
nor U9818 (N_9818,N_6934,N_6351);
xor U9819 (N_9819,N_6620,N_5355);
xnor U9820 (N_9820,N_7266,N_7453);
xor U9821 (N_9821,N_6325,N_5482);
or U9822 (N_9822,N_5092,N_7030);
xnor U9823 (N_9823,N_6713,N_6310);
nand U9824 (N_9824,N_6973,N_6574);
nand U9825 (N_9825,N_6296,N_5128);
xnor U9826 (N_9826,N_6652,N_6879);
and U9827 (N_9827,N_7079,N_6238);
nor U9828 (N_9828,N_6015,N_5951);
nand U9829 (N_9829,N_6985,N_5974);
and U9830 (N_9830,N_5127,N_6749);
and U9831 (N_9831,N_6473,N_7195);
nor U9832 (N_9832,N_5718,N_7169);
and U9833 (N_9833,N_6073,N_6378);
or U9834 (N_9834,N_6337,N_5208);
and U9835 (N_9835,N_5347,N_7157);
and U9836 (N_9836,N_7492,N_6512);
nand U9837 (N_9837,N_6126,N_6134);
nor U9838 (N_9838,N_5262,N_7472);
nor U9839 (N_9839,N_7423,N_5725);
or U9840 (N_9840,N_6191,N_5046);
nand U9841 (N_9841,N_7351,N_6747);
nand U9842 (N_9842,N_6325,N_5552);
and U9843 (N_9843,N_5419,N_5853);
or U9844 (N_9844,N_6504,N_5465);
nor U9845 (N_9845,N_5519,N_6870);
and U9846 (N_9846,N_5315,N_6841);
and U9847 (N_9847,N_6086,N_7205);
xor U9848 (N_9848,N_7075,N_6345);
xor U9849 (N_9849,N_5312,N_6985);
xor U9850 (N_9850,N_5760,N_6759);
or U9851 (N_9851,N_6077,N_6792);
nand U9852 (N_9852,N_6991,N_5087);
xnor U9853 (N_9853,N_5243,N_6214);
and U9854 (N_9854,N_5675,N_5182);
or U9855 (N_9855,N_5002,N_5109);
nor U9856 (N_9856,N_5338,N_7114);
xor U9857 (N_9857,N_5203,N_6384);
xnor U9858 (N_9858,N_6688,N_6876);
xnor U9859 (N_9859,N_6828,N_5343);
and U9860 (N_9860,N_6447,N_5789);
or U9861 (N_9861,N_6253,N_5327);
and U9862 (N_9862,N_5108,N_7226);
nand U9863 (N_9863,N_6385,N_7014);
xor U9864 (N_9864,N_6666,N_6542);
or U9865 (N_9865,N_5974,N_6102);
nand U9866 (N_9866,N_5446,N_6894);
nor U9867 (N_9867,N_5264,N_5163);
and U9868 (N_9868,N_5942,N_5672);
nor U9869 (N_9869,N_5824,N_5632);
nand U9870 (N_9870,N_6910,N_6182);
nor U9871 (N_9871,N_6985,N_6083);
nand U9872 (N_9872,N_7089,N_5454);
or U9873 (N_9873,N_6242,N_5888);
nor U9874 (N_9874,N_5318,N_6947);
and U9875 (N_9875,N_5498,N_7386);
and U9876 (N_9876,N_5513,N_5879);
nand U9877 (N_9877,N_5272,N_7143);
xnor U9878 (N_9878,N_6104,N_5522);
nor U9879 (N_9879,N_6873,N_7279);
nand U9880 (N_9880,N_5548,N_5868);
or U9881 (N_9881,N_6812,N_6199);
or U9882 (N_9882,N_6814,N_5336);
and U9883 (N_9883,N_5703,N_6972);
nand U9884 (N_9884,N_6724,N_7000);
and U9885 (N_9885,N_5592,N_6937);
nand U9886 (N_9886,N_6738,N_6136);
and U9887 (N_9887,N_6176,N_7024);
xnor U9888 (N_9888,N_5568,N_6421);
and U9889 (N_9889,N_7449,N_6728);
or U9890 (N_9890,N_6598,N_5966);
nor U9891 (N_9891,N_6972,N_6598);
nor U9892 (N_9892,N_5074,N_6003);
nand U9893 (N_9893,N_6503,N_5351);
nor U9894 (N_9894,N_7033,N_5000);
or U9895 (N_9895,N_7258,N_6268);
and U9896 (N_9896,N_6273,N_5058);
or U9897 (N_9897,N_5202,N_5571);
nor U9898 (N_9898,N_7207,N_5257);
nor U9899 (N_9899,N_5283,N_6596);
and U9900 (N_9900,N_7496,N_5943);
xor U9901 (N_9901,N_6277,N_6205);
and U9902 (N_9902,N_5116,N_7441);
or U9903 (N_9903,N_7479,N_7427);
nor U9904 (N_9904,N_6266,N_7230);
and U9905 (N_9905,N_7033,N_6956);
nor U9906 (N_9906,N_5392,N_6591);
or U9907 (N_9907,N_5714,N_7418);
xor U9908 (N_9908,N_5378,N_5498);
xor U9909 (N_9909,N_6892,N_5752);
xor U9910 (N_9910,N_6713,N_7491);
xor U9911 (N_9911,N_5296,N_6683);
nand U9912 (N_9912,N_5610,N_5223);
or U9913 (N_9913,N_6924,N_6543);
nand U9914 (N_9914,N_5663,N_6248);
or U9915 (N_9915,N_7108,N_6664);
and U9916 (N_9916,N_6647,N_6973);
nor U9917 (N_9917,N_6405,N_5794);
nand U9918 (N_9918,N_5401,N_6274);
xor U9919 (N_9919,N_6391,N_5986);
nor U9920 (N_9920,N_6151,N_6524);
xor U9921 (N_9921,N_5517,N_6175);
and U9922 (N_9922,N_7339,N_5738);
and U9923 (N_9923,N_6599,N_7265);
or U9924 (N_9924,N_5388,N_7460);
nor U9925 (N_9925,N_6293,N_7381);
or U9926 (N_9926,N_7137,N_6897);
xor U9927 (N_9927,N_5915,N_6341);
nand U9928 (N_9928,N_5509,N_5903);
or U9929 (N_9929,N_6976,N_7020);
and U9930 (N_9930,N_5322,N_5911);
or U9931 (N_9931,N_6302,N_7299);
xor U9932 (N_9932,N_5696,N_6577);
and U9933 (N_9933,N_5464,N_6072);
xor U9934 (N_9934,N_7254,N_6380);
nor U9935 (N_9935,N_5434,N_6108);
and U9936 (N_9936,N_5990,N_5862);
xnor U9937 (N_9937,N_6730,N_7423);
nand U9938 (N_9938,N_6045,N_5406);
nor U9939 (N_9939,N_6858,N_7037);
nand U9940 (N_9940,N_5992,N_6824);
xnor U9941 (N_9941,N_6675,N_6362);
and U9942 (N_9942,N_7232,N_5939);
and U9943 (N_9943,N_6438,N_6058);
nor U9944 (N_9944,N_7270,N_5333);
nor U9945 (N_9945,N_7353,N_5098);
and U9946 (N_9946,N_5621,N_6916);
nand U9947 (N_9947,N_6387,N_5807);
and U9948 (N_9948,N_7316,N_6744);
nand U9949 (N_9949,N_7401,N_5392);
nand U9950 (N_9950,N_5593,N_6119);
nor U9951 (N_9951,N_5087,N_5405);
and U9952 (N_9952,N_6551,N_6371);
and U9953 (N_9953,N_6990,N_6877);
or U9954 (N_9954,N_5214,N_6206);
nor U9955 (N_9955,N_6805,N_7253);
nand U9956 (N_9956,N_6374,N_5978);
nand U9957 (N_9957,N_7100,N_5695);
nor U9958 (N_9958,N_5892,N_6916);
nand U9959 (N_9959,N_6814,N_5422);
or U9960 (N_9960,N_7418,N_5395);
nand U9961 (N_9961,N_6654,N_5634);
xor U9962 (N_9962,N_6292,N_6092);
and U9963 (N_9963,N_5900,N_7396);
nand U9964 (N_9964,N_5978,N_6473);
or U9965 (N_9965,N_6516,N_6012);
and U9966 (N_9966,N_6798,N_7243);
or U9967 (N_9967,N_6377,N_7285);
or U9968 (N_9968,N_7048,N_6039);
or U9969 (N_9969,N_5211,N_7203);
xor U9970 (N_9970,N_6147,N_6470);
or U9971 (N_9971,N_6318,N_6123);
nor U9972 (N_9972,N_5509,N_6589);
or U9973 (N_9973,N_6799,N_5841);
or U9974 (N_9974,N_5661,N_5635);
and U9975 (N_9975,N_6376,N_6968);
nand U9976 (N_9976,N_5689,N_5666);
nor U9977 (N_9977,N_5565,N_6934);
nand U9978 (N_9978,N_6362,N_6552);
or U9979 (N_9979,N_7175,N_6295);
nand U9980 (N_9980,N_7429,N_5079);
nand U9981 (N_9981,N_7281,N_5660);
xor U9982 (N_9982,N_5625,N_7200);
nor U9983 (N_9983,N_7411,N_7090);
and U9984 (N_9984,N_7405,N_5472);
and U9985 (N_9985,N_6594,N_7193);
and U9986 (N_9986,N_5462,N_6514);
xor U9987 (N_9987,N_6563,N_6618);
xnor U9988 (N_9988,N_5497,N_5042);
and U9989 (N_9989,N_7044,N_6289);
and U9990 (N_9990,N_5629,N_7063);
nand U9991 (N_9991,N_6764,N_6412);
nor U9992 (N_9992,N_5018,N_6745);
xor U9993 (N_9993,N_6648,N_6833);
and U9994 (N_9994,N_5409,N_6917);
and U9995 (N_9995,N_5317,N_5730);
xnor U9996 (N_9996,N_5393,N_6458);
and U9997 (N_9997,N_5790,N_7272);
and U9998 (N_9998,N_6471,N_5700);
nand U9999 (N_9999,N_5123,N_5148);
nand U10000 (N_10000,N_8763,N_9265);
xor U10001 (N_10001,N_8820,N_8313);
and U10002 (N_10002,N_8621,N_9121);
and U10003 (N_10003,N_8261,N_7533);
or U10004 (N_10004,N_8776,N_8493);
and U10005 (N_10005,N_8685,N_8837);
and U10006 (N_10006,N_9344,N_7678);
xnor U10007 (N_10007,N_9490,N_8538);
or U10008 (N_10008,N_9492,N_9623);
or U10009 (N_10009,N_8600,N_7827);
xor U10010 (N_10010,N_9014,N_9363);
or U10011 (N_10011,N_7980,N_8233);
and U10012 (N_10012,N_8753,N_9205);
nand U10013 (N_10013,N_9092,N_8570);
nand U10014 (N_10014,N_9432,N_9782);
and U10015 (N_10015,N_9139,N_8551);
and U10016 (N_10016,N_9062,N_8043);
xnor U10017 (N_10017,N_9952,N_9064);
nor U10018 (N_10018,N_9898,N_8698);
nand U10019 (N_10019,N_9099,N_8929);
xor U10020 (N_10020,N_9727,N_9241);
or U10021 (N_10021,N_8396,N_9210);
and U10022 (N_10022,N_7527,N_9115);
nand U10023 (N_10023,N_7724,N_9017);
nand U10024 (N_10024,N_9221,N_9454);
nand U10025 (N_10025,N_7515,N_9076);
xor U10026 (N_10026,N_7816,N_8176);
nand U10027 (N_10027,N_9060,N_9132);
nor U10028 (N_10028,N_7855,N_7665);
xnor U10029 (N_10029,N_7556,N_7657);
and U10030 (N_10030,N_7634,N_9571);
xnor U10031 (N_10031,N_9788,N_9588);
nor U10032 (N_10032,N_7680,N_8772);
nand U10033 (N_10033,N_8849,N_8499);
or U10034 (N_10034,N_7535,N_8650);
nor U10035 (N_10035,N_8979,N_9854);
and U10036 (N_10036,N_9528,N_8535);
nand U10037 (N_10037,N_9359,N_9860);
and U10038 (N_10038,N_7615,N_9762);
nor U10039 (N_10039,N_9504,N_8879);
xnor U10040 (N_10040,N_8153,N_9067);
xor U10041 (N_10041,N_8874,N_7581);
xor U10042 (N_10042,N_9270,N_9969);
nor U10043 (N_10043,N_8523,N_9581);
nor U10044 (N_10044,N_7631,N_7741);
and U10045 (N_10045,N_9821,N_8182);
and U10046 (N_10046,N_8920,N_8652);
and U10047 (N_10047,N_9760,N_8312);
and U10048 (N_10048,N_8397,N_9983);
xor U10049 (N_10049,N_8302,N_7561);
nand U10050 (N_10050,N_9390,N_9547);
nor U10051 (N_10051,N_8567,N_8150);
nand U10052 (N_10052,N_8568,N_7997);
and U10053 (N_10053,N_9050,N_8077);
nor U10054 (N_10054,N_7887,N_9382);
and U10055 (N_10055,N_7956,N_8280);
nor U10056 (N_10056,N_8664,N_8234);
nor U10057 (N_10057,N_7659,N_9033);
nand U10058 (N_10058,N_8923,N_7675);
xnor U10059 (N_10059,N_7745,N_8980);
and U10060 (N_10060,N_9240,N_9140);
nor U10061 (N_10061,N_9219,N_9849);
nor U10062 (N_10062,N_9365,N_8156);
xor U10063 (N_10063,N_9745,N_7846);
nor U10064 (N_10064,N_7786,N_9930);
or U10065 (N_10065,N_7583,N_9790);
or U10066 (N_10066,N_7722,N_9312);
nor U10067 (N_10067,N_9595,N_9187);
and U10068 (N_10068,N_7594,N_8735);
or U10069 (N_10069,N_8269,N_9423);
nand U10070 (N_10070,N_9027,N_8033);
or U10071 (N_10071,N_8936,N_8554);
and U10072 (N_10072,N_9560,N_8368);
and U10073 (N_10073,N_9124,N_7946);
or U10074 (N_10074,N_9502,N_9280);
xor U10075 (N_10075,N_9512,N_8612);
or U10076 (N_10076,N_9942,N_9810);
nand U10077 (N_10077,N_8505,N_7670);
nand U10078 (N_10078,N_7560,N_7972);
or U10079 (N_10079,N_9051,N_8005);
nor U10080 (N_10080,N_8022,N_7942);
and U10081 (N_10081,N_7682,N_9933);
or U10082 (N_10082,N_8818,N_8447);
or U10083 (N_10083,N_9328,N_8046);
or U10084 (N_10084,N_9081,N_8216);
nor U10085 (N_10085,N_8205,N_9193);
or U10086 (N_10086,N_8995,N_9425);
and U10087 (N_10087,N_8266,N_9799);
xnor U10088 (N_10088,N_9052,N_7730);
xor U10089 (N_10089,N_8669,N_8301);
nor U10090 (N_10090,N_7517,N_8560);
xnor U10091 (N_10091,N_8789,N_8648);
or U10092 (N_10092,N_9204,N_9072);
xor U10093 (N_10093,N_8133,N_8056);
or U10094 (N_10094,N_8031,N_8985);
nand U10095 (N_10095,N_8157,N_9475);
nor U10096 (N_10096,N_9003,N_9738);
nor U10097 (N_10097,N_8802,N_9447);
nor U10098 (N_10098,N_9726,N_9729);
nand U10099 (N_10099,N_9215,N_7669);
or U10100 (N_10100,N_8581,N_7822);
nand U10101 (N_10101,N_8214,N_7812);
and U10102 (N_10102,N_9255,N_8722);
or U10103 (N_10103,N_7829,N_9961);
nand U10104 (N_10104,N_7947,N_8681);
nor U10105 (N_10105,N_9886,N_9178);
nand U10106 (N_10106,N_8132,N_8574);
or U10107 (N_10107,N_8419,N_8773);
nand U10108 (N_10108,N_8898,N_8781);
nor U10109 (N_10109,N_9833,N_7712);
nor U10110 (N_10110,N_8503,N_9181);
or U10111 (N_10111,N_8335,N_9922);
xnor U10112 (N_10112,N_8298,N_9574);
nand U10113 (N_10113,N_8712,N_8543);
or U10114 (N_10114,N_7937,N_8836);
or U10115 (N_10115,N_9201,N_7723);
nor U10116 (N_10116,N_8519,N_8974);
and U10117 (N_10117,N_7610,N_9755);
and U10118 (N_10118,N_9628,N_9674);
or U10119 (N_10119,N_7731,N_8321);
nand U10120 (N_10120,N_9895,N_8194);
nor U10121 (N_10121,N_8555,N_8012);
nand U10122 (N_10122,N_8891,N_9348);
and U10123 (N_10123,N_8666,N_9303);
nand U10124 (N_10124,N_7969,N_8798);
nor U10125 (N_10125,N_8809,N_9836);
or U10126 (N_10126,N_8792,N_7949);
nand U10127 (N_10127,N_8921,N_7586);
or U10128 (N_10128,N_7679,N_9576);
nor U10129 (N_10129,N_9398,N_9989);
nand U10130 (N_10130,N_7746,N_8162);
or U10131 (N_10131,N_7565,N_8528);
xor U10132 (N_10132,N_8453,N_9352);
nand U10133 (N_10133,N_7952,N_8747);
nand U10134 (N_10134,N_8464,N_9339);
and U10135 (N_10135,N_8177,N_7709);
or U10136 (N_10136,N_8721,N_9144);
and U10137 (N_10137,N_8801,N_9236);
and U10138 (N_10138,N_8160,N_8074);
nand U10139 (N_10139,N_9406,N_8673);
nand U10140 (N_10140,N_8127,N_9226);
and U10141 (N_10141,N_7697,N_7606);
or U10142 (N_10142,N_9884,N_9386);
and U10143 (N_10143,N_9596,N_8358);
and U10144 (N_10144,N_8830,N_9822);
nand U10145 (N_10145,N_8889,N_9349);
or U10146 (N_10146,N_9346,N_9702);
or U10147 (N_10147,N_7871,N_9223);
and U10148 (N_10148,N_7771,N_9307);
nand U10149 (N_10149,N_8649,N_7874);
nor U10150 (N_10150,N_9414,N_7803);
or U10151 (N_10151,N_9951,N_9258);
or U10152 (N_10152,N_8846,N_7708);
xor U10153 (N_10153,N_8126,N_7693);
or U10154 (N_10154,N_9217,N_8223);
or U10155 (N_10155,N_8040,N_8691);
or U10156 (N_10156,N_9921,N_9582);
nor U10157 (N_10157,N_9880,N_9503);
nor U10158 (N_10158,N_8224,N_8314);
xor U10159 (N_10159,N_8512,N_7611);
and U10160 (N_10160,N_7845,N_9722);
or U10161 (N_10161,N_8190,N_9834);
and U10162 (N_10162,N_9636,N_8151);
nor U10163 (N_10163,N_7639,N_7655);
nand U10164 (N_10164,N_8333,N_8938);
nor U10165 (N_10165,N_7976,N_7948);
nor U10166 (N_10166,N_9474,N_8690);
nand U10167 (N_10167,N_8785,N_8963);
nor U10168 (N_10168,N_9608,N_9681);
nor U10169 (N_10169,N_9486,N_8263);
or U10170 (N_10170,N_9924,N_7849);
nand U10171 (N_10171,N_7826,N_8348);
xnor U10172 (N_10172,N_8508,N_8706);
and U10173 (N_10173,N_7961,N_9794);
nor U10174 (N_10174,N_9230,N_7960);
xnor U10175 (N_10175,N_8981,N_9616);
xor U10176 (N_10176,N_9527,N_8482);
xor U10177 (N_10177,N_8588,N_9604);
nor U10178 (N_10178,N_8622,N_8563);
or U10179 (N_10179,N_7766,N_7760);
nor U10180 (N_10180,N_8867,N_8851);
xnor U10181 (N_10181,N_9610,N_8810);
and U10182 (N_10182,N_7792,N_7643);
or U10183 (N_10183,N_9536,N_9514);
xor U10184 (N_10184,N_9387,N_8848);
nand U10185 (N_10185,N_9764,N_9036);
and U10186 (N_10186,N_7881,N_7676);
nor U10187 (N_10187,N_8948,N_9519);
or U10188 (N_10188,N_8273,N_8219);
xor U10189 (N_10189,N_8096,N_8517);
or U10190 (N_10190,N_8500,N_9974);
nand U10191 (N_10191,N_9698,N_8367);
and U10192 (N_10192,N_8978,N_8684);
nor U10193 (N_10193,N_9809,N_9332);
or U10194 (N_10194,N_9059,N_9781);
xor U10195 (N_10195,N_8495,N_8520);
and U10196 (N_10196,N_9626,N_7981);
and U10197 (N_10197,N_9295,N_8217);
nor U10198 (N_10198,N_8199,N_8770);
nor U10199 (N_10199,N_8530,N_8803);
nand U10200 (N_10200,N_9257,N_8148);
and U10201 (N_10201,N_9057,N_9195);
nand U10202 (N_10202,N_9479,N_8433);
and U10203 (N_10203,N_8972,N_9366);
xor U10204 (N_10204,N_8470,N_9102);
and U10205 (N_10205,N_9997,N_8839);
nor U10206 (N_10206,N_9859,N_9850);
nor U10207 (N_10207,N_7711,N_9553);
xnor U10208 (N_10208,N_9721,N_8865);
xor U10209 (N_10209,N_9373,N_8346);
and U10210 (N_10210,N_8427,N_7988);
nand U10211 (N_10211,N_7662,N_9773);
xor U10212 (N_10212,N_9237,N_8062);
and U10213 (N_10213,N_8525,N_9499);
nand U10214 (N_10214,N_7649,N_7970);
and U10215 (N_10215,N_9744,N_9966);
and U10216 (N_10216,N_8221,N_8870);
xor U10217 (N_10217,N_8052,N_9111);
xor U10218 (N_10218,N_9523,N_9956);
nor U10219 (N_10219,N_9965,N_9125);
and U10220 (N_10220,N_8276,N_9761);
or U10221 (N_10221,N_8483,N_8643);
and U10222 (N_10222,N_9070,N_7735);
and U10223 (N_10223,N_9182,N_8039);
or U10224 (N_10224,N_9866,N_9973);
xnor U10225 (N_10225,N_7895,N_9899);
and U10226 (N_10226,N_8458,N_7577);
nor U10227 (N_10227,N_9007,N_9090);
and U10228 (N_10228,N_8328,N_8204);
nor U10229 (N_10229,N_7526,N_8001);
nor U10230 (N_10230,N_9500,N_8063);
xnor U10231 (N_10231,N_7602,N_8539);
nor U10232 (N_10232,N_8169,N_9540);
nor U10233 (N_10233,N_7836,N_9273);
xor U10234 (N_10234,N_9700,N_9709);
nand U10235 (N_10235,N_7914,N_7633);
or U10236 (N_10236,N_9220,N_9167);
nand U10237 (N_10237,N_9460,N_7592);
and U10238 (N_10238,N_8415,N_9559);
xor U10239 (N_10239,N_8641,N_7739);
nand U10240 (N_10240,N_8275,N_9483);
xnor U10241 (N_10241,N_9106,N_7617);
nand U10242 (N_10242,N_8585,N_9618);
nor U10243 (N_10243,N_8872,N_8060);
and U10244 (N_10244,N_9287,N_8890);
nor U10245 (N_10245,N_8754,N_9671);
nor U10246 (N_10246,N_7523,N_8324);
or U10247 (N_10247,N_8278,N_9994);
nand U10248 (N_10248,N_7572,N_9877);
xor U10249 (N_10249,N_8767,N_8198);
xnor U10250 (N_10250,N_9345,N_8013);
and U10251 (N_10251,N_9658,N_7777);
nor U10252 (N_10252,N_8845,N_8000);
xor U10253 (N_10253,N_8394,N_8454);
nand U10254 (N_10254,N_9645,N_7768);
nor U10255 (N_10255,N_9413,N_9879);
xnor U10256 (N_10256,N_8674,N_8137);
or U10257 (N_10257,N_9455,N_7753);
or U10258 (N_10258,N_8120,N_8431);
xnor U10259 (N_10259,N_9998,N_8203);
xnor U10260 (N_10260,N_9024,N_7886);
nor U10261 (N_10261,N_8507,N_8953);
nand U10262 (N_10262,N_9048,N_9823);
xnor U10263 (N_10263,N_8697,N_9196);
nor U10264 (N_10264,N_7548,N_9557);
nor U10265 (N_10265,N_8784,N_8315);
and U10266 (N_10266,N_9861,N_9131);
or U10267 (N_10267,N_9278,N_9640);
and U10268 (N_10268,N_8759,N_7719);
xnor U10269 (N_10269,N_9575,N_7628);
or U10270 (N_10270,N_9279,N_8533);
or U10271 (N_10271,N_9775,N_8518);
nand U10272 (N_10272,N_8240,N_8758);
or U10273 (N_10273,N_8576,N_8626);
and U10274 (N_10274,N_8951,N_9362);
nand U10275 (N_10275,N_8918,N_9228);
or U10276 (N_10276,N_9937,N_8277);
or U10277 (N_10277,N_7504,N_9152);
nor U10278 (N_10278,N_8756,N_8462);
and U10279 (N_10279,N_8195,N_8465);
or U10280 (N_10280,N_8192,N_8049);
nor U10281 (N_10281,N_9372,N_8187);
nor U10282 (N_10282,N_8322,N_8343);
and U10283 (N_10283,N_8893,N_9683);
and U10284 (N_10284,N_9157,N_8937);
nor U10285 (N_10285,N_9569,N_8687);
nor U10286 (N_10286,N_9056,N_9171);
and U10287 (N_10287,N_8511,N_8596);
nand U10288 (N_10288,N_8619,N_9495);
and U10289 (N_10289,N_9094,N_7685);
and U10290 (N_10290,N_8252,N_7637);
nor U10291 (N_10291,N_7806,N_8943);
and U10292 (N_10292,N_9692,N_8279);
xnor U10293 (N_10293,N_9355,N_8091);
nor U10294 (N_10294,N_7957,N_9396);
or U10295 (N_10295,N_9199,N_9511);
nor U10296 (N_10296,N_7817,N_8099);
xor U10297 (N_10297,N_7557,N_7522);
nor U10298 (N_10298,N_9768,N_9785);
nand U10299 (N_10299,N_9804,N_8124);
or U10300 (N_10300,N_8375,N_9754);
nor U10301 (N_10301,N_8434,N_9939);
nor U10302 (N_10302,N_8496,N_7654);
nor U10303 (N_10303,N_7773,N_7530);
or U10304 (N_10304,N_8268,N_9958);
or U10305 (N_10305,N_9103,N_8579);
nand U10306 (N_10306,N_8877,N_9246);
or U10307 (N_10307,N_9548,N_9192);
nand U10308 (N_10308,N_7564,N_8966);
or U10309 (N_10309,N_7793,N_7933);
or U10310 (N_10310,N_7707,N_7541);
xnor U10311 (N_10311,N_9837,N_9710);
or U10312 (N_10312,N_9964,N_8924);
xor U10313 (N_10313,N_8603,N_8961);
or U10314 (N_10314,N_7732,N_9112);
nor U10315 (N_10315,N_9530,N_8633);
or U10316 (N_10316,N_8249,N_8693);
nand U10317 (N_10317,N_9686,N_9868);
xnor U10318 (N_10318,N_8862,N_7779);
xnor U10319 (N_10319,N_9224,N_7906);
nor U10320 (N_10320,N_8718,N_7733);
and U10321 (N_10321,N_9133,N_9395);
xnor U10322 (N_10322,N_8125,N_8983);
nor U10323 (N_10323,N_8702,N_8954);
or U10324 (N_10324,N_9637,N_9286);
nor U10325 (N_10325,N_8391,N_9408);
nor U10326 (N_10326,N_8976,N_9107);
nor U10327 (N_10327,N_9206,N_8286);
and U10328 (N_10328,N_9542,N_9429);
xor U10329 (N_10329,N_9233,N_7700);
nor U10330 (N_10330,N_9872,N_7798);
nor U10331 (N_10331,N_8474,N_8880);
or U10332 (N_10332,N_7668,N_7959);
nor U10333 (N_10333,N_8984,N_8740);
or U10334 (N_10334,N_7683,N_9855);
and U10335 (N_10335,N_7562,N_9962);
nor U10336 (N_10336,N_7772,N_9767);
or U10337 (N_10337,N_8208,N_7532);
nand U10338 (N_10338,N_8410,N_9579);
or U10339 (N_10339,N_8061,N_8259);
nor U10340 (N_10340,N_8294,N_9337);
and U10341 (N_10341,N_8429,N_8683);
nand U10342 (N_10342,N_9119,N_9218);
xnor U10343 (N_10343,N_7630,N_8293);
nand U10344 (N_10344,N_7944,N_8804);
nor U10345 (N_10345,N_8509,N_9302);
xnor U10346 (N_10346,N_8360,N_8181);
nand U10347 (N_10347,N_7831,N_7998);
and U10348 (N_10348,N_8311,N_7783);
xnor U10349 (N_10349,N_8786,N_9129);
xnor U10350 (N_10350,N_9802,N_9725);
or U10351 (N_10351,N_8009,N_9720);
nand U10352 (N_10352,N_7842,N_9696);
or U10353 (N_10353,N_9585,N_8371);
and U10354 (N_10354,N_8308,N_9970);
and U10355 (N_10355,N_9805,N_9538);
or U10356 (N_10356,N_7785,N_9870);
nand U10357 (N_10357,N_8537,N_7646);
xor U10358 (N_10358,N_8841,N_8264);
xor U10359 (N_10359,N_9083,N_9156);
and U10360 (N_10360,N_9838,N_9465);
and U10361 (N_10361,N_9315,N_9290);
xor U10362 (N_10362,N_8138,N_8689);
nand U10363 (N_10363,N_7703,N_9308);
nand U10364 (N_10364,N_9065,N_9874);
nand U10365 (N_10365,N_8292,N_9501);
nor U10366 (N_10366,N_8032,N_7977);
nor U10367 (N_10367,N_8631,N_9082);
xnor U10368 (N_10368,N_8919,N_8935);
nand U10369 (N_10369,N_8143,N_8004);
xor U10370 (N_10370,N_9096,N_8858);
xnor U10371 (N_10371,N_9740,N_9126);
or U10372 (N_10372,N_9282,N_7814);
and U10373 (N_10373,N_8144,N_9545);
xnor U10374 (N_10374,N_8670,N_8154);
or U10375 (N_10375,N_8905,N_8010);
nand U10376 (N_10376,N_9748,N_7767);
nand U10377 (N_10377,N_8593,N_7689);
nor U10378 (N_10378,N_7726,N_7923);
xor U10379 (N_10379,N_8957,N_8986);
xor U10380 (N_10380,N_8656,N_7913);
nor U10381 (N_10381,N_9587,N_9418);
xnor U10382 (N_10382,N_9409,N_8017);
and U10383 (N_10383,N_7716,N_8220);
or U10384 (N_10384,N_7559,N_7549);
and U10385 (N_10385,N_9778,N_9202);
nor U10386 (N_10386,N_7811,N_8244);
and U10387 (N_10387,N_7922,N_8088);
nand U10388 (N_10388,N_8828,N_9049);
and U10389 (N_10389,N_8882,N_8296);
nor U10390 (N_10390,N_9960,N_8534);
nand U10391 (N_10391,N_8078,N_7607);
xnor U10392 (N_10392,N_8466,N_9467);
or U10393 (N_10393,N_9622,N_9586);
xnor U10394 (N_10394,N_9943,N_7930);
and U10395 (N_10395,N_9814,N_8553);
nand U10396 (N_10396,N_9992,N_9589);
nand U10397 (N_10397,N_9967,N_8896);
nor U10398 (N_10398,N_8305,N_9630);
nor U10399 (N_10399,N_7908,N_7671);
and U10400 (N_10400,N_9166,N_9304);
and U10401 (N_10401,N_7996,N_9824);
nor U10402 (N_10402,N_8339,N_8541);
nand U10403 (N_10403,N_7815,N_8742);
nand U10404 (N_10404,N_8559,N_9292);
and U10405 (N_10405,N_7694,N_8881);
nand U10406 (N_10406,N_9032,N_9285);
nor U10407 (N_10407,N_9815,N_9599);
nand U10408 (N_10408,N_8734,N_8737);
xor U10409 (N_10409,N_8284,N_7544);
nand U10410 (N_10410,N_9949,N_8393);
or U10411 (N_10411,N_9252,N_9333);
or U10412 (N_10412,N_9819,N_8939);
or U10413 (N_10413,N_9926,N_8100);
or U10414 (N_10414,N_8575,N_9058);
nand U10415 (N_10415,N_9914,N_7832);
xnor U10416 (N_10416,N_7984,N_9276);
xor U10417 (N_10417,N_8178,N_7904);
xnor U10418 (N_10418,N_8340,N_9468);
and U10419 (N_10419,N_8744,N_9708);
nand U10420 (N_10420,N_9020,N_9335);
nand U10421 (N_10421,N_7851,N_9300);
or U10422 (N_10422,N_8232,N_8445);
or U10423 (N_10423,N_7626,N_8444);
or U10424 (N_10424,N_7859,N_7931);
nor U10425 (N_10425,N_9361,N_7938);
nor U10426 (N_10426,N_8136,N_8123);
and U10427 (N_10427,N_7663,N_8826);
or U10428 (N_10428,N_8486,N_9912);
or U10429 (N_10429,N_7576,N_7860);
xor U10430 (N_10430,N_8775,N_8788);
nor U10431 (N_10431,N_9040,N_8726);
or U10432 (N_10432,N_8569,N_8583);
nor U10433 (N_10433,N_8404,N_9869);
nand U10434 (N_10434,N_9143,N_9045);
and U10435 (N_10435,N_9077,N_8374);
nor U10436 (N_10436,N_9981,N_9200);
or U10437 (N_10437,N_7775,N_7691);
and U10438 (N_10438,N_7713,N_9897);
nor U10439 (N_10439,N_7876,N_9505);
xnor U10440 (N_10440,N_8873,N_9243);
xor U10441 (N_10441,N_9054,N_9347);
or U10442 (N_10442,N_8871,N_9289);
and U10443 (N_10443,N_9403,N_8527);
nor U10444 (N_10444,N_9158,N_8956);
nor U10445 (N_10445,N_9325,N_9263);
and U10446 (N_10446,N_8186,N_8868);
or U10447 (N_10447,N_8614,N_9110);
nand U10448 (N_10448,N_9247,N_7995);
or U10449 (N_10449,N_9660,N_8632);
or U10450 (N_10450,N_9421,N_8813);
or U10451 (N_10451,N_9741,N_7762);
and U10452 (N_10452,N_8502,N_8065);
or U10453 (N_10453,N_7717,N_9118);
xor U10454 (N_10454,N_9602,N_9625);
or U10455 (N_10455,N_8455,N_8736);
or U10456 (N_10456,N_8058,N_7748);
nor U10457 (N_10457,N_8959,N_8594);
nand U10458 (N_10458,N_9953,N_8987);
and U10459 (N_10459,N_9491,N_8129);
or U10460 (N_10460,N_9004,N_8330);
or U10461 (N_10461,N_8488,N_8657);
nand U10462 (N_10462,N_9774,N_7585);
nand U10463 (N_10463,N_7640,N_9480);
and U10464 (N_10464,N_9902,N_8790);
nor U10465 (N_10465,N_8437,N_8420);
xor U10466 (N_10466,N_7941,N_9911);
and U10467 (N_10467,N_9259,N_9177);
nand U10468 (N_10468,N_8679,N_7764);
nor U10469 (N_10469,N_7840,N_8051);
nand U10470 (N_10470,N_8634,N_9842);
or U10471 (N_10471,N_8732,N_9841);
or U10472 (N_10472,N_7936,N_8226);
nor U10473 (N_10473,N_8498,N_8636);
xnor U10474 (N_10474,N_8101,N_9010);
and U10475 (N_10475,N_9305,N_8625);
or U10476 (N_10476,N_7858,N_8930);
nor U10477 (N_10477,N_8942,N_8070);
nor U10478 (N_10478,N_9168,N_8696);
or U10479 (N_10479,N_9524,N_7701);
nand U10480 (N_10480,N_9030,N_8762);
or U10481 (N_10481,N_9063,N_8605);
xnor U10482 (N_10482,N_8272,N_8536);
nor U10483 (N_10483,N_7967,N_9648);
nor U10484 (N_10484,N_8069,N_8036);
nor U10485 (N_10485,N_7833,N_7677);
nor U10486 (N_10486,N_8714,N_7774);
nand U10487 (N_10487,N_9714,N_8895);
nand U10488 (N_10488,N_8202,N_9456);
and U10489 (N_10489,N_9670,N_8200);
nor U10490 (N_10490,N_8095,N_8316);
nand U10491 (N_10491,N_9901,N_8900);
and U10492 (N_10492,N_8651,N_9776);
xor U10493 (N_10493,N_8338,N_8440);
xor U10494 (N_10494,N_8089,N_7943);
nor U10495 (N_10495,N_8728,N_9319);
and U10496 (N_10496,N_9294,N_8377);
xnor U10497 (N_10497,N_8422,N_9717);
nand U10498 (N_10498,N_8183,N_8675);
xor U10499 (N_10499,N_8430,N_8692);
nand U10500 (N_10500,N_9183,N_9935);
xor U10501 (N_10501,N_7605,N_8059);
or U10502 (N_10502,N_9370,N_8540);
and U10503 (N_10503,N_7964,N_8155);
or U10504 (N_10504,N_8323,N_8586);
nand U10505 (N_10505,N_9448,N_7695);
or U10506 (N_10506,N_9894,N_8635);
and U10507 (N_10507,N_9232,N_7536);
xnor U10508 (N_10508,N_8122,N_7958);
xnor U10509 (N_10509,N_8327,N_9412);
or U10510 (N_10510,N_8840,N_9369);
or U10511 (N_10511,N_9878,N_9411);
nand U10512 (N_10512,N_8805,N_7656);
nand U10513 (N_10513,N_8045,N_8428);
xor U10514 (N_10514,N_7704,N_8011);
or U10515 (N_10515,N_9662,N_8794);
and U10516 (N_10516,N_7818,N_7761);
xnor U10517 (N_10517,N_7917,N_8452);
and U10518 (N_10518,N_7608,N_8640);
xor U10519 (N_10519,N_7892,N_9123);
and U10520 (N_10520,N_9546,N_9175);
and U10521 (N_10521,N_9401,N_9567);
nand U10522 (N_10522,N_8085,N_7935);
or U10523 (N_10523,N_8128,N_8071);
or U10524 (N_10524,N_9055,N_7516);
nor U10525 (N_10525,N_8236,N_8970);
or U10526 (N_10526,N_9564,N_8513);
or U10527 (N_10527,N_9179,N_7890);
nor U10528 (N_10528,N_9254,N_8908);
or U10529 (N_10529,N_8090,N_7974);
nand U10530 (N_10530,N_8925,N_9507);
xor U10531 (N_10531,N_9797,N_7505);
nor U10532 (N_10532,N_7919,N_8285);
and U10533 (N_10533,N_7720,N_9825);
and U10534 (N_10534,N_8875,N_8587);
or U10535 (N_10535,N_9578,N_8412);
nand U10536 (N_10536,N_8899,N_8564);
and U10537 (N_10537,N_8663,N_8325);
and U10538 (N_10538,N_8345,N_7993);
xnor U10539 (N_10539,N_8532,N_9013);
nor U10540 (N_10540,N_9851,N_9174);
and U10541 (N_10541,N_8876,N_8075);
or U10542 (N_10542,N_8102,N_7924);
or U10543 (N_10543,N_9991,N_9863);
and U10544 (N_10544,N_8149,N_9358);
or U10545 (N_10545,N_7983,N_8299);
nand U10546 (N_10546,N_9871,N_9881);
xnor U10547 (N_10547,N_8073,N_8647);
nor U10548 (N_10548,N_8146,N_7912);
nor U10549 (N_10549,N_9194,N_7721);
and U10550 (N_10550,N_9617,N_7578);
or U10551 (N_10551,N_9169,N_8379);
and U10552 (N_10552,N_7807,N_9719);
nor U10553 (N_10553,N_7511,N_9407);
nand U10554 (N_10554,N_8709,N_8812);
and U10555 (N_10555,N_9478,N_8719);
xor U10556 (N_10556,N_9813,N_7620);
nor U10557 (N_10557,N_9451,N_9556);
xnor U10558 (N_10558,N_8725,N_9526);
xnor U10559 (N_10559,N_8573,N_9685);
nand U10560 (N_10560,N_9306,N_9443);
and U10561 (N_10561,N_8418,N_7910);
and U10562 (N_10562,N_9917,N_9397);
nor U10563 (N_10563,N_8355,N_7804);
and U10564 (N_10564,N_9136,N_7901);
nor U10565 (N_10565,N_9812,N_9803);
or U10566 (N_10566,N_8475,N_8050);
nand U10567 (N_10567,N_8222,N_8850);
nor U10568 (N_10568,N_7614,N_9261);
or U10569 (N_10569,N_8897,N_8246);
and U10570 (N_10570,N_8741,N_8592);
xnor U10571 (N_10571,N_8115,N_9605);
or U10572 (N_10572,N_8406,N_7673);
or U10573 (N_10573,N_9439,N_9453);
xnor U10574 (N_10574,N_8460,N_7879);
nand U10575 (N_10575,N_8238,N_7765);
xnor U10576 (N_10576,N_8861,N_9379);
nor U10577 (N_10577,N_8081,N_9155);
nand U10578 (N_10578,N_7755,N_9262);
or U10579 (N_10579,N_8707,N_7575);
or U10580 (N_10580,N_8912,N_7600);
and U10581 (N_10581,N_8212,N_8584);
xnor U10582 (N_10582,N_8515,N_9985);
nor U10583 (N_10583,N_9577,N_8254);
xor U10584 (N_10584,N_8598,N_9795);
or U10585 (N_10585,N_8667,N_8931);
and U10586 (N_10586,N_9378,N_7644);
or U10587 (N_10587,N_9022,N_9404);
nand U10588 (N_10588,N_9242,N_8996);
nand U10589 (N_10589,N_8903,N_7973);
nor U10590 (N_10590,N_8602,N_8711);
and U10591 (N_10591,N_8514,N_8274);
or U10592 (N_10592,N_8552,N_9384);
xnor U10593 (N_10593,N_9915,N_7763);
nand U10594 (N_10594,N_9149,N_7945);
nand U10595 (N_10595,N_9002,N_9274);
nor U10596 (N_10596,N_7555,N_7553);
or U10597 (N_10597,N_8265,N_9634);
nand U10598 (N_10598,N_7570,N_9853);
and U10599 (N_10599,N_8724,N_8550);
and U10600 (N_10600,N_8832,N_8910);
and U10601 (N_10601,N_9712,N_8381);
nor U10602 (N_10602,N_9646,N_9963);
or U10603 (N_10603,N_9376,N_9919);
xnor U10604 (N_10604,N_8353,N_8386);
xor U10605 (N_10605,N_7542,N_9089);
or U10606 (N_10606,N_9927,N_9713);
nand U10607 (N_10607,N_8962,N_7869);
or U10608 (N_10608,N_9517,N_8119);
or U10609 (N_10609,N_7591,N_9458);
nand U10610 (N_10610,N_7690,N_7878);
xnor U10611 (N_10611,N_8161,N_7514);
xor U10612 (N_10612,N_7508,N_8947);
or U10613 (N_10613,N_9100,N_9627);
and U10614 (N_10614,N_9513,N_8811);
nand U10615 (N_10615,N_9529,N_8441);
xnor U10616 (N_10616,N_9946,N_9612);
nor U10617 (N_10617,N_9104,N_8782);
and U10618 (N_10618,N_8489,N_9955);
nor U10619 (N_10619,N_8516,N_9108);
nor U10620 (N_10620,N_8578,N_9808);
xnor U10621 (N_10621,N_9137,N_8041);
and U10622 (N_10622,N_9561,N_9765);
nand U10623 (N_10623,N_7622,N_7987);
xor U10624 (N_10624,N_7698,N_9669);
nand U10625 (N_10625,N_9750,N_9449);
xnor U10626 (N_10626,N_8411,N_8914);
or U10627 (N_10627,N_9298,N_8565);
nor U10628 (N_10628,N_9235,N_9520);
and U10629 (N_10629,N_8363,N_8915);
or U10630 (N_10630,N_9791,N_8822);
nor U10631 (N_10631,N_8218,N_9704);
nand U10632 (N_10632,N_9271,N_9105);
nand U10633 (N_10633,N_9975,N_8185);
nor U10634 (N_10634,N_8791,N_8907);
or U10635 (N_10635,N_8864,N_9856);
and U10636 (N_10636,N_9078,N_9857);
or U10637 (N_10637,N_8751,N_7790);
or U10638 (N_10638,N_8179,N_8270);
or U10639 (N_10639,N_7621,N_8020);
xor U10640 (N_10640,N_9817,N_9555);
nor U10641 (N_10641,N_9093,N_8019);
xnor U10642 (N_10642,N_7603,N_9896);
nor U10643 (N_10643,N_7580,N_9839);
and U10644 (N_10644,N_8531,N_9891);
nand U10645 (N_10645,N_9843,N_8023);
and U10646 (N_10646,N_8407,N_8400);
nand U10647 (N_10647,N_9984,N_9145);
or U10648 (N_10648,N_9549,N_8171);
and U10649 (N_10649,N_7747,N_9929);
nand U10650 (N_10650,N_9716,N_9473);
or U10651 (N_10651,N_9260,N_8795);
or U10652 (N_10652,N_8816,N_7820);
xnor U10653 (N_10653,N_9356,N_9959);
and U10654 (N_10654,N_9668,N_9086);
or U10655 (N_10655,N_8589,N_9807);
xnor U10656 (N_10656,N_9170,N_8960);
nand U10657 (N_10657,N_8958,N_9916);
nand U10658 (N_10658,N_7734,N_7579);
xnor U10659 (N_10659,N_8357,N_7797);
xor U10660 (N_10660,N_8524,N_8723);
nand U10661 (N_10661,N_9715,N_8457);
or U10662 (N_10662,N_7838,N_9619);
nand U10663 (N_10663,N_7926,N_7563);
xnor U10664 (N_10664,N_8739,N_8170);
nor U10665 (N_10665,N_9739,N_9753);
nor U10666 (N_10666,N_9436,N_8885);
and U10667 (N_10667,N_7558,N_8716);
or U10668 (N_10668,N_8624,N_9497);
xnor U10669 (N_10669,N_8613,N_8941);
or U10670 (N_10670,N_7791,N_8620);
and U10671 (N_10671,N_7645,N_7501);
xnor U10672 (N_10672,N_9583,N_8799);
nor U10673 (N_10673,N_9665,N_9430);
and U10674 (N_10674,N_9239,N_7925);
and U10675 (N_10675,N_7540,N_8764);
and U10676 (N_10676,N_9084,N_7571);
or U10677 (N_10677,N_8174,N_8118);
nand U10678 (N_10678,N_9887,N_9173);
or U10679 (N_10679,N_9999,N_7687);
nand U10680 (N_10680,N_8104,N_9554);
nand U10681 (N_10681,N_9786,N_8291);
nand U10682 (N_10682,N_8267,N_9350);
nand U10683 (N_10683,N_9338,N_9353);
nand U10684 (N_10684,N_9734,N_9482);
nor U10685 (N_10685,N_7568,N_7990);
or U10686 (N_10686,N_8351,N_8504);
nor U10687 (N_10687,N_9165,N_7883);
xor U10688 (N_10688,N_8968,N_9977);
or U10689 (N_10689,N_7978,N_9611);
nand U10690 (N_10690,N_9873,N_7975);
and U10691 (N_10691,N_7582,N_9128);
nor U10692 (N_10692,N_9591,N_9888);
and U10693 (N_10693,N_9766,N_9367);
nor U10694 (N_10694,N_9222,N_9180);
nand U10695 (N_10695,N_8206,N_7900);
and U10696 (N_10696,N_9694,N_8892);
nor U10697 (N_10697,N_8599,N_7781);
and U10698 (N_10698,N_9566,N_9109);
nand U10699 (N_10699,N_8364,N_8034);
or U10700 (N_10700,N_9769,N_8660);
and U10701 (N_10701,N_9161,N_8201);
and U10702 (N_10702,N_7864,N_8468);
and U10703 (N_10703,N_8977,N_8435);
nand U10704 (N_10704,N_9890,N_8998);
and U10705 (N_10705,N_8855,N_9299);
or U10706 (N_10706,N_8147,N_9489);
and U10707 (N_10707,N_8366,N_7819);
xnor U10708 (N_10708,N_9392,N_8833);
xor U10709 (N_10709,N_8901,N_8637);
nand U10710 (N_10710,N_7823,N_8478);
xor U10711 (N_10711,N_9831,N_8713);
or U10712 (N_10712,N_7648,N_8952);
or U10713 (N_10713,N_9091,N_8306);
or U10714 (N_10714,N_8117,N_8743);
nand U10715 (N_10715,N_7598,N_8843);
nor U10716 (N_10716,N_8601,N_9368);
nand U10717 (N_10717,N_9213,N_8401);
nor U10718 (N_10718,N_9798,N_8571);
and U10719 (N_10719,N_7629,N_9296);
nand U10720 (N_10720,N_8193,N_7954);
and U10721 (N_10721,N_8997,N_8035);
and U10722 (N_10722,N_8695,N_8755);
or U10723 (N_10723,N_8629,N_8940);
xor U10724 (N_10724,N_9954,N_7905);
xnor U10725 (N_10725,N_8164,N_8165);
nand U10726 (N_10726,N_7503,N_7710);
xnor U10727 (N_10727,N_9042,N_8082);
nor U10728 (N_10728,N_8271,N_7623);
and U10729 (N_10729,N_8370,N_9488);
nand U10730 (N_10730,N_8704,N_8990);
nor U10731 (N_10731,N_8337,N_7599);
nor U10732 (N_10732,N_8392,N_8037);
xor U10733 (N_10733,N_8448,N_8319);
nor U10734 (N_10734,N_8446,N_8159);
nand U10735 (N_10735,N_9153,N_8310);
nor U10736 (N_10736,N_9730,N_8395);
or U10737 (N_10737,N_9190,N_9987);
nor U10738 (N_10738,N_8745,N_9940);
or U10739 (N_10739,N_7813,N_9250);
nor U10740 (N_10740,N_8175,N_9464);
or U10741 (N_10741,N_9659,N_8655);
nor U10742 (N_10742,N_8038,N_9724);
and U10743 (N_10743,N_8591,N_8015);
nor U10744 (N_10744,N_9531,N_8439);
nor U10745 (N_10745,N_9597,N_8191);
nand U10746 (N_10746,N_8645,N_7911);
xor U10747 (N_10747,N_9584,N_9508);
xnor U10748 (N_10748,N_7543,N_9445);
xnor U10749 (N_10749,N_8965,N_9317);
nand U10750 (N_10750,N_8072,N_9663);
xnor U10751 (N_10751,N_9046,N_9789);
xor U10752 (N_10752,N_9044,N_9657);
nand U10753 (N_10753,N_8545,N_9148);
or U10754 (N_10754,N_9707,N_9928);
nor U10755 (N_10755,N_9426,N_8424);
or U10756 (N_10756,N_8354,N_7660);
and U10757 (N_10757,N_8860,N_7661);
xnor U10758 (N_10758,N_9909,N_9718);
nor U10759 (N_10759,N_8021,N_9268);
nand U10760 (N_10760,N_9703,N_9080);
xnor U10761 (N_10761,N_8479,N_8548);
nor U10762 (N_10762,N_9322,N_8079);
or U10763 (N_10763,N_9840,N_9023);
or U10764 (N_10764,N_9457,N_9327);
xnor U10765 (N_10765,N_9518,N_7778);
xor U10766 (N_10766,N_8853,N_9818);
or U10767 (N_10767,N_9532,N_9649);
nand U10768 (N_10768,N_8245,N_8800);
xnor U10769 (N_10769,N_9986,N_8442);
and U10770 (N_10770,N_9422,N_7986);
nand U10771 (N_10771,N_8066,N_8607);
nand U10772 (N_10772,N_7744,N_9164);
xnor U10773 (N_10773,N_9521,N_7940);
and U10774 (N_10774,N_9639,N_9198);
xor U10775 (N_10775,N_7889,N_8329);
nand U10776 (N_10776,N_9208,N_9689);
nor U10777 (N_10777,N_7567,N_9419);
and U10778 (N_10778,N_7547,N_8026);
xnor U10779 (N_10779,N_8662,N_9087);
and U10780 (N_10780,N_8255,N_7590);
xnor U10781 (N_10781,N_9227,N_7759);
xnor U10782 (N_10782,N_8934,N_8093);
or U10783 (N_10783,N_7861,N_7953);
nand U10784 (N_10784,N_8720,N_8057);
and U10785 (N_10785,N_9141,N_7554);
and U10786 (N_10786,N_8113,N_8611);
nor U10787 (N_10787,N_7934,N_7872);
nor U10788 (N_10788,N_9780,N_8779);
nor U10789 (N_10789,N_9679,N_7740);
or U10790 (N_10790,N_7604,N_9053);
xor U10791 (N_10791,N_8213,N_9827);
and U10792 (N_10792,N_8387,N_8210);
nor U10793 (N_10793,N_9021,N_9238);
nor U10794 (N_10794,N_9918,N_9134);
nand U10795 (N_10795,N_9435,N_8821);
nor U10796 (N_10796,N_9472,N_8971);
or U10797 (N_10797,N_9459,N_8361);
xnor U10798 (N_10798,N_8054,N_8449);
nand U10799 (N_10799,N_7539,N_9652);
xnor U10800 (N_10800,N_8003,N_9424);
or U10801 (N_10801,N_9142,N_9621);
or U10802 (N_10802,N_9968,N_8916);
xor U10803 (N_10803,N_9427,N_7593);
or U10804 (N_10804,N_8869,N_9098);
nand U10805 (N_10805,N_9672,N_7776);
nand U10806 (N_10806,N_9310,N_7574);
or U10807 (N_10807,N_7985,N_8944);
nor U10808 (N_10808,N_8922,N_9651);
and U10809 (N_10809,N_7758,N_9678);
xor U10810 (N_10810,N_9079,N_9151);
and U10811 (N_10811,N_9537,N_9095);
xor U10812 (N_10812,N_8256,N_7989);
xnor U10813 (N_10813,N_7821,N_9947);
nor U10814 (N_10814,N_8703,N_9214);
or U10815 (N_10815,N_9341,N_7750);
or U10816 (N_10816,N_7500,N_8638);
or U10817 (N_10817,N_8109,N_7616);
nand U10818 (N_10818,N_8863,N_8617);
nand U10819 (N_10819,N_8933,N_8825);
nor U10820 (N_10820,N_9197,N_8443);
nor U10821 (N_10821,N_8909,N_9736);
or U10822 (N_10822,N_8973,N_9437);
and U10823 (N_10823,N_7787,N_9229);
and U10824 (N_10824,N_8894,N_9284);
xnor U10825 (N_10825,N_8257,N_9399);
and U10826 (N_10826,N_9620,N_9590);
or U10827 (N_10827,N_9675,N_9493);
nand U10828 (N_10828,N_8064,N_7519);
and U10829 (N_10829,N_7625,N_9688);
and U10830 (N_10830,N_7856,N_7962);
nor U10831 (N_10831,N_8130,N_9127);
or U10832 (N_10832,N_9309,N_9978);
xor U10833 (N_10833,N_9920,N_7714);
or U10834 (N_10834,N_8653,N_8682);
or U10835 (N_10835,N_9749,N_7715);
xor U10836 (N_10836,N_8362,N_8700);
nor U10837 (N_10837,N_9673,N_8608);
nand U10838 (N_10838,N_9638,N_8492);
xnor U10839 (N_10839,N_8911,N_8006);
or U10840 (N_10840,N_7866,N_9757);
nand U10841 (N_10841,N_8086,N_8783);
nor U10842 (N_10842,N_7898,N_7524);
xor U10843 (N_10843,N_7552,N_9931);
or U10844 (N_10844,N_9009,N_9948);
xor U10845 (N_10845,N_9075,N_8932);
xnor U10846 (N_10846,N_8857,N_7612);
nor U10847 (N_10847,N_9330,N_8477);
xor U10848 (N_10848,N_8260,N_9442);
and U10849 (N_10849,N_9598,N_7854);
and U10850 (N_10850,N_7770,N_8526);
and U10851 (N_10851,N_8926,N_9534);
xor U10852 (N_10852,N_9029,N_7518);
nor U10853 (N_10853,N_9275,N_9043);
xor U10854 (N_10854,N_9535,N_7950);
xnor U10855 (N_10855,N_9551,N_7613);
nand U10856 (N_10856,N_9865,N_8024);
and U10857 (N_10857,N_7636,N_9037);
xnor U10858 (N_10858,N_9122,N_7857);
or U10859 (N_10859,N_8884,N_7796);
nand U10860 (N_10860,N_7870,N_8529);
and U10861 (N_10861,N_8107,N_9162);
or U10862 (N_10862,N_9905,N_9297);
nand U10863 (N_10863,N_9188,N_8556);
xor U10864 (N_10864,N_7538,N_7966);
nor U10865 (N_10865,N_9469,N_8184);
or U10866 (N_10866,N_9320,N_8806);
xnor U10867 (N_10867,N_8028,N_8797);
xor U10868 (N_10868,N_9624,N_8152);
or U10869 (N_10869,N_9291,N_8577);
and U10870 (N_10870,N_9941,N_9541);
xor U10871 (N_10871,N_9471,N_9130);
nand U10872 (N_10872,N_8262,N_9883);
xnor U10873 (N_10873,N_9699,N_7550);
nor U10874 (N_10874,N_8807,N_8173);
xor U10875 (N_10875,N_9976,N_9701);
and U10876 (N_10876,N_7529,N_8604);
nand U10877 (N_10877,N_8999,N_7546);
nor U10878 (N_10878,N_8388,N_7844);
xnor U10879 (N_10879,N_8627,N_8644);
xor U10880 (N_10880,N_8414,N_9900);
xor U10881 (N_10881,N_9594,N_9147);
and U10882 (N_10882,N_7706,N_7853);
or U10883 (N_10883,N_7520,N_8859);
nor U10884 (N_10884,N_9892,N_9381);
and U10885 (N_10885,N_9828,N_7834);
nand U10886 (N_10886,N_8417,N_7868);
nand U10887 (N_10887,N_9006,N_9374);
and U10888 (N_10888,N_8134,N_9770);
xor U10889 (N_10889,N_9420,N_9431);
nand U10890 (N_10890,N_8838,N_7652);
nand U10891 (N_10891,N_9485,N_9209);
nand U10892 (N_10892,N_8309,N_9743);
nor U10893 (N_10893,N_7907,N_9272);
nor U10894 (N_10894,N_9015,N_7569);
nor U10895 (N_10895,N_9038,N_8510);
nand U10896 (N_10896,N_9867,N_8092);
or U10897 (N_10897,N_8002,N_8141);
and U10898 (N_10898,N_9733,N_8053);
nand U10899 (N_10899,N_9677,N_7929);
nand U10900 (N_10900,N_8852,N_8317);
and U10901 (N_10901,N_7799,N_9073);
xnor U10902 (N_10902,N_7696,N_8111);
nor U10903 (N_10903,N_8904,N_8044);
xnor U10904 (N_10904,N_7751,N_8087);
nor U10905 (N_10905,N_8835,N_9820);
xor U10906 (N_10906,N_8522,N_7754);
and U10907 (N_10907,N_8334,N_9568);
nor U10908 (N_10908,N_7800,N_8659);
or U10909 (N_10909,N_8562,N_8350);
or U10910 (N_10910,N_9031,N_8746);
nor U10911 (N_10911,N_8572,N_8352);
xnor U10912 (N_10912,N_9606,N_9433);
or U10913 (N_10913,N_9697,N_8777);
or U10914 (N_10914,N_8331,N_9380);
nor U10915 (N_10915,N_8661,N_9120);
nor U10916 (N_10916,N_8398,N_9163);
xnor U10917 (N_10917,N_9498,N_9787);
nand U10918 (N_10918,N_9644,N_8402);
nor U10919 (N_10919,N_8768,N_8139);
and U10920 (N_10920,N_9515,N_8250);
and U10921 (N_10921,N_7835,N_7647);
nor U10922 (N_10922,N_9572,N_9441);
xor U10923 (N_10923,N_7736,N_8288);
xor U10924 (N_10924,N_8975,N_7674);
xor U10925 (N_10925,N_8131,N_7828);
and U10926 (N_10926,N_9680,N_8796);
nor U10927 (N_10927,N_8646,N_7551);
and U10928 (N_10928,N_8172,N_8927);
nor U10929 (N_10929,N_8484,N_9071);
or U10930 (N_10930,N_7916,N_8686);
nand U10931 (N_10931,N_7688,N_9329);
and U10932 (N_10932,N_7743,N_9643);
nor U10933 (N_10933,N_7880,N_8106);
nor U10934 (N_10934,N_7601,N_9088);
nand U10935 (N_10935,N_7897,N_7865);
xor U10936 (N_10936,N_8769,N_9923);
xor U10937 (N_10937,N_8103,N_8727);
nor U10938 (N_10938,N_9615,N_8542);
nor U10939 (N_10939,N_7903,N_7839);
xnor U10940 (N_10940,N_7939,N_8609);
nor U10941 (N_10941,N_8752,N_8780);
or U10942 (N_10942,N_8694,N_8142);
and U10943 (N_10943,N_8778,N_9793);
and U10944 (N_10944,N_9806,N_8671);
or U10945 (N_10945,N_7534,N_9383);
nor U10946 (N_10946,N_8623,N_9288);
and U10947 (N_10947,N_8558,N_7862);
xor U10948 (N_10948,N_9661,N_9847);
nor U10949 (N_10949,N_8042,N_9533);
nand U10950 (N_10950,N_7902,N_7588);
nand U10951 (N_10951,N_9385,N_9035);
or U10952 (N_10952,N_7802,N_9248);
or U10953 (N_10953,N_9462,N_9028);
nand U10954 (N_10954,N_9377,N_9340);
nand U10955 (N_10955,N_8228,N_8561);
xor U10956 (N_10956,N_9728,N_7684);
or U10957 (N_10957,N_7531,N_7882);
or U10958 (N_10958,N_7837,N_8094);
or U10959 (N_10959,N_8341,N_7597);
xor U10960 (N_10960,N_9846,N_9391);
xnor U10961 (N_10961,N_9466,N_8823);
or U10962 (N_10962,N_7788,N_8461);
or U10963 (N_10963,N_8678,N_9746);
or U10964 (N_10964,N_8708,N_8808);
nor U10965 (N_10965,N_9751,N_9522);
nand U10966 (N_10966,N_8618,N_8557);
nand U10967 (N_10967,N_7737,N_9629);
or U10968 (N_10968,N_8580,N_8993);
nand U10969 (N_10969,N_9394,N_8405);
and U10970 (N_10970,N_8365,N_9101);
xor U10971 (N_10971,N_7632,N_8231);
nand U10972 (N_10972,N_9191,N_8856);
and U10973 (N_10973,N_9440,N_9826);
or U10974 (N_10974,N_8385,N_9331);
nand U10975 (N_10975,N_7587,N_8994);
xor U10976 (N_10976,N_7843,N_8076);
xor U10977 (N_10977,N_8701,N_9906);
and U10978 (N_10978,N_9470,N_7506);
nor U10979 (N_10979,N_9313,N_8450);
and U10980 (N_10980,N_8582,N_9784);
nand U10981 (N_10981,N_9324,N_8318);
nand U10982 (N_10982,N_8167,N_9667);
nand U10983 (N_10983,N_9047,N_9552);
xnor U10984 (N_10984,N_9256,N_9184);
xnor U10985 (N_10985,N_9811,N_8369);
and U10986 (N_10986,N_9647,N_9026);
nor U10987 (N_10987,N_9687,N_7894);
and U10988 (N_10988,N_9543,N_9012);
xnor U10989 (N_10989,N_8408,N_9580);
or U10990 (N_10990,N_8389,N_8688);
or U10991 (N_10991,N_8665,N_8463);
xor U10992 (N_10992,N_9225,N_8967);
xor U10993 (N_10993,N_8295,N_9903);
nand U10994 (N_10994,N_7850,N_9019);
or U10995 (N_10995,N_8121,N_8467);
and U10996 (N_10996,N_9150,N_8438);
nor U10997 (N_10997,N_8372,N_8084);
nor U10998 (N_10998,N_8342,N_8116);
xnor U10999 (N_10999,N_9207,N_7729);
or U11000 (N_11000,N_8243,N_7738);
nand U11001 (N_11001,N_9160,N_9097);
or U11002 (N_11002,N_8988,N_8765);
nor U11003 (N_11003,N_9938,N_8456);
nor U11004 (N_11004,N_8731,N_8886);
and U11005 (N_11005,N_9463,N_8158);
and U11006 (N_11006,N_9000,N_8227);
nor U11007 (N_11007,N_9450,N_8491);
nor U11008 (N_11008,N_8831,N_9438);
and U11009 (N_11009,N_9510,N_7769);
nor U11010 (N_11010,N_7545,N_8878);
nand U11011 (N_11011,N_9654,N_8715);
nor U11012 (N_11012,N_7885,N_8787);
nand U11013 (N_11013,N_9360,N_8991);
nor U11014 (N_11014,N_9573,N_9848);
nor U11015 (N_11015,N_7681,N_9357);
xor U11016 (N_11016,N_9034,N_7847);
nor U11017 (N_11017,N_9783,N_9434);
and U11018 (N_11018,N_9539,N_8403);
nor U11019 (N_11019,N_9417,N_8472);
xnor U11020 (N_11020,N_8668,N_8610);
and U11021 (N_11021,N_8114,N_8844);
nor U11022 (N_11022,N_8029,N_9779);
nand U11023 (N_11023,N_8373,N_9506);
and U11024 (N_11024,N_8320,N_9154);
xnor U11025 (N_11025,N_8730,N_8229);
xor U11026 (N_11026,N_8251,N_7528);
and U11027 (N_11027,N_9653,N_7651);
or U11028 (N_11028,N_8654,N_8188);
nor U11029 (N_11029,N_8383,N_9172);
nand U11030 (N_11030,N_7502,N_8761);
or U11031 (N_11031,N_9613,N_9316);
and U11032 (N_11032,N_7932,N_8738);
nor U11033 (N_11033,N_7979,N_8888);
nor U11034 (N_11034,N_8819,N_9655);
nand U11035 (N_11035,N_8964,N_7658);
and U11036 (N_11036,N_8055,N_9844);
xnor U11037 (N_11037,N_8196,N_8766);
and U11038 (N_11038,N_8382,N_9607);
and U11039 (N_11039,N_8239,N_8390);
nand U11040 (N_11040,N_9945,N_8025);
nor U11041 (N_11041,N_9641,N_8950);
nor U11042 (N_11042,N_7877,N_9972);
and U11043 (N_11043,N_8854,N_8423);
and U11044 (N_11044,N_8699,N_8717);
or U11045 (N_11045,N_9005,N_7825);
xnor U11046 (N_11046,N_8949,N_9635);
and U11047 (N_11047,N_8282,N_9016);
nor U11048 (N_11048,N_8297,N_8628);
and U11049 (N_11049,N_7808,N_8928);
or U11050 (N_11050,N_9862,N_8774);
and U11051 (N_11051,N_8887,N_9601);
nand U11052 (N_11052,N_8140,N_8108);
nand U11053 (N_11053,N_8955,N_9908);
and U11054 (N_11054,N_8237,N_8359);
nor U11055 (N_11055,N_7510,N_9907);
nand U11056 (N_11056,N_9041,N_7650);
and U11057 (N_11057,N_8098,N_9114);
nor U11058 (N_11058,N_7782,N_9614);
xnor U11059 (N_11059,N_9801,N_9293);
nor U11060 (N_11060,N_9875,N_9957);
nand U11061 (N_11061,N_8241,N_9609);
and U11062 (N_11062,N_9711,N_7909);
and U11063 (N_11063,N_9266,N_7584);
and U11064 (N_11064,N_9666,N_9550);
and U11065 (N_11065,N_7664,N_7809);
and U11066 (N_11066,N_7638,N_7915);
nand U11067 (N_11067,N_9146,N_9354);
and U11068 (N_11068,N_7928,N_8566);
nand U11069 (N_11069,N_9001,N_8501);
and U11070 (N_11070,N_9910,N_9477);
nor U11071 (N_11071,N_7692,N_8672);
xor U11072 (N_11072,N_8110,N_9737);
nor U11073 (N_11073,N_8189,N_9845);
nand U11074 (N_11074,N_8546,N_8068);
or U11075 (N_11075,N_8356,N_7968);
nor U11076 (N_11076,N_9138,N_8290);
nand U11077 (N_11077,N_8658,N_8135);
and U11078 (N_11078,N_7635,N_8235);
or U11079 (N_11079,N_9684,N_7752);
xor U11080 (N_11080,N_8521,N_7521);
and U11081 (N_11081,N_7852,N_8326);
nand U11082 (N_11082,N_9267,N_7875);
nand U11083 (N_11083,N_7795,N_7686);
nand U11084 (N_11084,N_9664,N_7992);
or U11085 (N_11085,N_9759,N_7728);
or U11086 (N_11086,N_9444,N_9777);
and U11087 (N_11087,N_9415,N_7873);
nand U11088 (N_11088,N_9203,N_9446);
or U11089 (N_11089,N_9245,N_9732);
xnor U11090 (N_11090,N_9388,N_9944);
xnor U11091 (N_11091,N_7756,N_9496);
xor U11092 (N_11092,N_9069,N_8814);
or U11093 (N_11093,N_8416,N_9185);
nor U11094 (N_11094,N_8547,N_7884);
nor U11095 (N_11095,N_9889,N_8485);
nor U11096 (N_11096,N_8494,N_9835);
nor U11097 (N_11097,N_9830,N_8982);
xnor U11098 (N_11098,N_8180,N_9690);
or U11099 (N_11099,N_9936,N_9068);
nor U11100 (N_11100,N_9253,N_9693);
or U11101 (N_11101,N_9993,N_7965);
xnor U11102 (N_11102,N_9742,N_8027);
and U11103 (N_11103,N_9375,N_8230);
or U11104 (N_11104,N_8459,N_9558);
xor U11105 (N_11105,N_9025,N_8705);
xor U11106 (N_11106,N_7867,N_7955);
nor U11107 (N_11107,N_9428,N_8606);
xor U11108 (N_11108,N_7641,N_8750);
nor U11109 (N_11109,N_9800,N_9314);
nor U11110 (N_11110,N_9832,N_9979);
and U11111 (N_11111,N_8842,N_9189);
or U11112 (N_11112,N_9885,N_9212);
nor U11113 (N_11113,N_9735,N_7667);
xor U11114 (N_11114,N_9277,N_9563);
nor U11115 (N_11115,N_9321,N_8757);
or U11116 (N_11116,N_7672,N_7619);
and U11117 (N_11117,N_9342,N_7920);
nor U11118 (N_11118,N_8680,N_8487);
and U11119 (N_11119,N_7537,N_9336);
or U11120 (N_11120,N_9950,N_8112);
nand U11121 (N_11121,N_8347,N_8815);
and U11122 (N_11122,N_7699,N_7653);
or U11123 (N_11123,N_7824,N_9393);
nand U11124 (N_11124,N_9525,N_9676);
nor U11125 (N_11125,N_8506,N_8677);
xnor U11126 (N_11126,N_9251,N_8030);
xnor U11127 (N_11127,N_8480,N_7963);
nand U11128 (N_11128,N_7566,N_8902);
and U11129 (N_11129,N_9593,N_8376);
xor U11130 (N_11130,N_8197,N_8425);
xor U11131 (N_11131,N_9758,N_8749);
xnor U11132 (N_11132,N_9705,N_9980);
or U11133 (N_11133,N_9600,N_9632);
nand U11134 (N_11134,N_9706,N_7589);
nor U11135 (N_11135,N_8595,N_8166);
and U11136 (N_11136,N_8303,N_8018);
nor U11137 (N_11137,N_9509,N_7971);
nor U11138 (N_11138,N_8105,N_9516);
nand U11139 (N_11139,N_9400,N_9633);
xor U11140 (N_11140,N_9481,N_9264);
or U11141 (N_11141,N_9756,N_9476);
xor U11142 (N_11142,N_8642,N_8597);
nor U11143 (N_11143,N_7725,N_8917);
or U11144 (N_11144,N_7780,N_9932);
or U11145 (N_11145,N_7991,N_7951);
nor U11146 (N_11146,N_8432,N_8413);
and U11147 (N_11147,N_8332,N_9249);
nor U11148 (N_11148,N_8906,N_8258);
xor U11149 (N_11149,N_9864,N_7888);
and U11150 (N_11150,N_9410,N_8913);
nor U11151 (N_11151,N_8426,N_9996);
nand U11152 (N_11152,N_8289,N_8616);
and U11153 (N_11153,N_8209,N_9792);
nand U11154 (N_11154,N_9631,N_7848);
and U11155 (N_11155,N_9592,N_8163);
or U11156 (N_11156,N_8378,N_7830);
nor U11157 (N_11157,N_9747,N_9039);
nor U11158 (N_11158,N_9343,N_7727);
nand U11159 (N_11159,N_8883,N_7642);
xnor U11160 (N_11160,N_7784,N_8946);
nand U11161 (N_11161,N_8047,N_8590);
nand U11162 (N_11162,N_9995,N_9283);
or U11163 (N_11163,N_8242,N_9650);
nor U11164 (N_11164,N_9018,N_9269);
and U11165 (N_11165,N_7921,N_8615);
nor U11166 (N_11166,N_8771,N_9893);
xnor U11167 (N_11167,N_7618,N_8436);
nor U11168 (N_11168,N_8945,N_7742);
nor U11169 (N_11169,N_8215,N_9117);
nor U11170 (N_11170,N_8349,N_8989);
or U11171 (N_11171,N_8497,N_7512);
and U11172 (N_11172,N_7805,N_9752);
and U11173 (N_11173,N_7789,N_9988);
nor U11174 (N_11174,N_9934,N_7757);
and U11175 (N_11175,N_9405,N_9402);
xor U11176 (N_11176,N_8336,N_7595);
and U11177 (N_11177,N_9389,N_9176);
nand U11178 (N_11178,N_8793,N_9461);
nand U11179 (N_11179,N_8014,N_8168);
or U11180 (N_11180,N_9008,N_9816);
xnor U11181 (N_11181,N_8639,N_8549);
or U11182 (N_11182,N_9135,N_8409);
and U11183 (N_11183,N_9695,N_7794);
and U11184 (N_11184,N_7899,N_8829);
nor U11185 (N_11185,N_7982,N_9723);
or U11186 (N_11186,N_7702,N_8817);
or U11187 (N_11187,N_8283,N_9982);
xor U11188 (N_11188,N_8225,N_7627);
nand U11189 (N_11189,N_8007,N_8287);
or U11190 (N_11190,N_9913,N_8676);
and U11191 (N_11191,N_9326,N_9318);
nand U11192 (N_11192,N_8344,N_7749);
nand U11193 (N_11193,N_8384,N_9771);
or U11194 (N_11194,N_8247,N_7841);
and U11195 (N_11195,N_8248,N_7999);
nand U11196 (N_11196,N_9494,N_8834);
xnor U11197 (N_11197,N_8421,N_7801);
and U11198 (N_11198,N_9691,N_8207);
nand U11199 (N_11199,N_8481,N_8469);
or U11200 (N_11200,N_9334,N_9971);
nor U11201 (N_11201,N_9544,N_8083);
and U11202 (N_11202,N_9925,N_7994);
nor U11203 (N_11203,N_8544,N_8097);
nor U11204 (N_11204,N_8630,N_8490);
nand U11205 (N_11205,N_8476,N_8827);
nor U11206 (N_11206,N_8471,N_8281);
nand U11207 (N_11207,N_9113,N_8866);
nor U11208 (N_11208,N_8211,N_9570);
nand U11209 (N_11209,N_9085,N_7718);
or U11210 (N_11210,N_7513,N_9452);
nor U11211 (N_11211,N_8307,N_8733);
or U11212 (N_11212,N_9642,N_9159);
nor U11213 (N_11213,N_7705,N_9311);
xor U11214 (N_11214,N_7863,N_8451);
nor U11215 (N_11215,N_7624,N_7927);
or U11216 (N_11216,N_8473,N_8080);
nand U11217 (N_11217,N_9061,N_8729);
nor U11218 (N_11218,N_9858,N_9074);
xor U11219 (N_11219,N_7609,N_8145);
nor U11220 (N_11220,N_9731,N_9603);
xnor U11221 (N_11221,N_7507,N_8710);
xor U11222 (N_11222,N_7891,N_7596);
nand U11223 (N_11223,N_8067,N_8760);
and U11224 (N_11224,N_7525,N_9772);
and U11225 (N_11225,N_8304,N_9876);
nor U11226 (N_11226,N_9301,N_9990);
nor U11227 (N_11227,N_9066,N_9656);
xnor U11228 (N_11228,N_8992,N_9351);
nor U11229 (N_11229,N_9281,N_9904);
or U11230 (N_11230,N_9852,N_9211);
nand U11231 (N_11231,N_9116,N_9763);
or U11232 (N_11232,N_9487,N_9416);
nand U11233 (N_11233,N_8048,N_9562);
and U11234 (N_11234,N_8380,N_9484);
nand U11235 (N_11235,N_7573,N_9244);
nor U11236 (N_11236,N_8300,N_9323);
nor U11237 (N_11237,N_9682,N_9231);
or U11238 (N_11238,N_7896,N_9011);
or U11239 (N_11239,N_7893,N_7666);
or U11240 (N_11240,N_8969,N_9186);
nor U11241 (N_11241,N_9882,N_8847);
and U11242 (N_11242,N_9796,N_8824);
or U11243 (N_11243,N_8748,N_9234);
nor U11244 (N_11244,N_8008,N_7810);
and U11245 (N_11245,N_8399,N_9565);
and U11246 (N_11246,N_9829,N_9364);
nor U11247 (N_11247,N_7918,N_9216);
nor U11248 (N_11248,N_8016,N_9371);
nor U11249 (N_11249,N_7509,N_8253);
nor U11250 (N_11250,N_7614,N_9018);
nand U11251 (N_11251,N_9747,N_8099);
nor U11252 (N_11252,N_8168,N_8489);
xnor U11253 (N_11253,N_9335,N_8949);
xor U11254 (N_11254,N_8444,N_8939);
and U11255 (N_11255,N_9174,N_9971);
and U11256 (N_11256,N_8148,N_8765);
or U11257 (N_11257,N_7785,N_7766);
xnor U11258 (N_11258,N_8872,N_8242);
nor U11259 (N_11259,N_9420,N_8070);
or U11260 (N_11260,N_9791,N_9611);
nand U11261 (N_11261,N_9582,N_7959);
nand U11262 (N_11262,N_9781,N_8300);
nand U11263 (N_11263,N_9691,N_9024);
nor U11264 (N_11264,N_7781,N_9841);
nand U11265 (N_11265,N_9559,N_8014);
nor U11266 (N_11266,N_7718,N_9860);
nor U11267 (N_11267,N_8637,N_8066);
xor U11268 (N_11268,N_8283,N_9964);
or U11269 (N_11269,N_8133,N_9813);
and U11270 (N_11270,N_9875,N_9650);
xor U11271 (N_11271,N_8078,N_9256);
nand U11272 (N_11272,N_9461,N_7746);
and U11273 (N_11273,N_7713,N_9879);
or U11274 (N_11274,N_8118,N_9461);
xnor U11275 (N_11275,N_8685,N_7995);
nand U11276 (N_11276,N_7800,N_9197);
or U11277 (N_11277,N_7694,N_8967);
or U11278 (N_11278,N_9503,N_8967);
nor U11279 (N_11279,N_8566,N_8374);
or U11280 (N_11280,N_7978,N_7692);
nand U11281 (N_11281,N_9996,N_9786);
nand U11282 (N_11282,N_8990,N_8646);
or U11283 (N_11283,N_9008,N_8299);
nor U11284 (N_11284,N_7689,N_9717);
xnor U11285 (N_11285,N_9114,N_9386);
and U11286 (N_11286,N_8216,N_8111);
or U11287 (N_11287,N_9040,N_7531);
nand U11288 (N_11288,N_8446,N_8527);
xnor U11289 (N_11289,N_8463,N_9237);
or U11290 (N_11290,N_8502,N_7893);
or U11291 (N_11291,N_7540,N_9921);
nor U11292 (N_11292,N_8682,N_8022);
and U11293 (N_11293,N_7816,N_7552);
xnor U11294 (N_11294,N_9937,N_7985);
nor U11295 (N_11295,N_7930,N_8572);
xnor U11296 (N_11296,N_7668,N_9866);
nor U11297 (N_11297,N_7798,N_8487);
nand U11298 (N_11298,N_7913,N_9660);
and U11299 (N_11299,N_9835,N_9959);
nor U11300 (N_11300,N_8618,N_9864);
or U11301 (N_11301,N_9810,N_8221);
nand U11302 (N_11302,N_8221,N_8904);
nand U11303 (N_11303,N_7984,N_8092);
nand U11304 (N_11304,N_7560,N_9022);
and U11305 (N_11305,N_8902,N_8291);
nand U11306 (N_11306,N_9200,N_8460);
nand U11307 (N_11307,N_8698,N_9049);
xnor U11308 (N_11308,N_8236,N_8032);
and U11309 (N_11309,N_9187,N_7731);
nand U11310 (N_11310,N_9206,N_7769);
xor U11311 (N_11311,N_7970,N_8100);
nor U11312 (N_11312,N_7898,N_9305);
or U11313 (N_11313,N_8961,N_9535);
xnor U11314 (N_11314,N_9722,N_8464);
and U11315 (N_11315,N_7532,N_8249);
nor U11316 (N_11316,N_9908,N_7569);
xor U11317 (N_11317,N_7856,N_7664);
nor U11318 (N_11318,N_9455,N_8745);
or U11319 (N_11319,N_9195,N_9712);
nand U11320 (N_11320,N_8746,N_9646);
or U11321 (N_11321,N_8284,N_9415);
and U11322 (N_11322,N_9866,N_8975);
or U11323 (N_11323,N_8622,N_8340);
nor U11324 (N_11324,N_7941,N_8345);
nand U11325 (N_11325,N_8866,N_9679);
nand U11326 (N_11326,N_7873,N_9027);
xnor U11327 (N_11327,N_9225,N_9996);
and U11328 (N_11328,N_8072,N_8471);
and U11329 (N_11329,N_9168,N_9632);
nor U11330 (N_11330,N_7664,N_8027);
xnor U11331 (N_11331,N_9646,N_7793);
nor U11332 (N_11332,N_8692,N_8781);
or U11333 (N_11333,N_9814,N_7801);
or U11334 (N_11334,N_9089,N_9643);
nand U11335 (N_11335,N_9840,N_9245);
nand U11336 (N_11336,N_8840,N_7758);
nor U11337 (N_11337,N_9788,N_9227);
or U11338 (N_11338,N_9317,N_8547);
xor U11339 (N_11339,N_9499,N_9995);
xor U11340 (N_11340,N_9841,N_7778);
and U11341 (N_11341,N_9272,N_9680);
or U11342 (N_11342,N_9789,N_7607);
and U11343 (N_11343,N_7553,N_9850);
nor U11344 (N_11344,N_8125,N_9389);
nand U11345 (N_11345,N_8562,N_7855);
and U11346 (N_11346,N_8052,N_9686);
and U11347 (N_11347,N_9740,N_8117);
xnor U11348 (N_11348,N_8962,N_8968);
nand U11349 (N_11349,N_7565,N_9965);
xor U11350 (N_11350,N_7938,N_9998);
or U11351 (N_11351,N_7839,N_8344);
nor U11352 (N_11352,N_8522,N_9950);
nand U11353 (N_11353,N_9554,N_7941);
xnor U11354 (N_11354,N_9822,N_9043);
or U11355 (N_11355,N_9965,N_9247);
xor U11356 (N_11356,N_8133,N_7854);
nand U11357 (N_11357,N_7931,N_7845);
or U11358 (N_11358,N_9525,N_9008);
nor U11359 (N_11359,N_8897,N_7623);
and U11360 (N_11360,N_9191,N_9608);
and U11361 (N_11361,N_8164,N_8500);
xnor U11362 (N_11362,N_9849,N_8757);
or U11363 (N_11363,N_9127,N_7736);
nor U11364 (N_11364,N_9741,N_9972);
xnor U11365 (N_11365,N_8770,N_7735);
nand U11366 (N_11366,N_7794,N_8139);
and U11367 (N_11367,N_9554,N_9297);
nand U11368 (N_11368,N_7814,N_8706);
xor U11369 (N_11369,N_8902,N_8766);
nand U11370 (N_11370,N_9015,N_8393);
nand U11371 (N_11371,N_9228,N_9810);
and U11372 (N_11372,N_9019,N_9380);
xor U11373 (N_11373,N_9489,N_7809);
or U11374 (N_11374,N_7800,N_8082);
nand U11375 (N_11375,N_9994,N_8637);
or U11376 (N_11376,N_8032,N_9635);
or U11377 (N_11377,N_8293,N_7963);
nand U11378 (N_11378,N_7930,N_8145);
xnor U11379 (N_11379,N_9299,N_9396);
or U11380 (N_11380,N_8818,N_9269);
xor U11381 (N_11381,N_9082,N_7707);
or U11382 (N_11382,N_9053,N_8064);
nor U11383 (N_11383,N_7856,N_8076);
or U11384 (N_11384,N_8493,N_7836);
and U11385 (N_11385,N_7690,N_9922);
nor U11386 (N_11386,N_8927,N_9110);
xnor U11387 (N_11387,N_7908,N_8438);
nand U11388 (N_11388,N_7779,N_9109);
nand U11389 (N_11389,N_8087,N_7770);
or U11390 (N_11390,N_8029,N_9080);
or U11391 (N_11391,N_9514,N_9577);
nand U11392 (N_11392,N_9926,N_8777);
and U11393 (N_11393,N_8444,N_8566);
or U11394 (N_11394,N_9831,N_7881);
and U11395 (N_11395,N_7636,N_8222);
and U11396 (N_11396,N_8144,N_8633);
xor U11397 (N_11397,N_8429,N_9763);
nand U11398 (N_11398,N_8080,N_9957);
nand U11399 (N_11399,N_8854,N_9960);
and U11400 (N_11400,N_8298,N_7746);
nand U11401 (N_11401,N_8923,N_7559);
nor U11402 (N_11402,N_8149,N_9442);
or U11403 (N_11403,N_7582,N_9104);
xnor U11404 (N_11404,N_8119,N_8366);
or U11405 (N_11405,N_9039,N_7988);
or U11406 (N_11406,N_8247,N_7586);
or U11407 (N_11407,N_9649,N_7620);
or U11408 (N_11408,N_9496,N_7612);
xor U11409 (N_11409,N_9132,N_9861);
nor U11410 (N_11410,N_8538,N_8995);
and U11411 (N_11411,N_8257,N_9169);
nand U11412 (N_11412,N_8602,N_7514);
xnor U11413 (N_11413,N_8360,N_8554);
nor U11414 (N_11414,N_9772,N_9545);
xor U11415 (N_11415,N_9471,N_8033);
or U11416 (N_11416,N_9161,N_7726);
nor U11417 (N_11417,N_8834,N_8998);
nand U11418 (N_11418,N_7609,N_8370);
xnor U11419 (N_11419,N_9664,N_9571);
and U11420 (N_11420,N_8011,N_7879);
and U11421 (N_11421,N_9768,N_7600);
nand U11422 (N_11422,N_8945,N_9112);
and U11423 (N_11423,N_7511,N_8277);
nor U11424 (N_11424,N_9017,N_7896);
nor U11425 (N_11425,N_7714,N_9530);
nor U11426 (N_11426,N_7685,N_8427);
or U11427 (N_11427,N_9816,N_8618);
nand U11428 (N_11428,N_8557,N_7775);
xor U11429 (N_11429,N_8068,N_8694);
nor U11430 (N_11430,N_8046,N_7654);
nand U11431 (N_11431,N_9233,N_9745);
nand U11432 (N_11432,N_9516,N_7672);
xor U11433 (N_11433,N_8618,N_8770);
or U11434 (N_11434,N_9874,N_8359);
xor U11435 (N_11435,N_8944,N_9129);
or U11436 (N_11436,N_8187,N_9692);
nor U11437 (N_11437,N_7707,N_8599);
nor U11438 (N_11438,N_7753,N_9990);
nand U11439 (N_11439,N_9249,N_7771);
xor U11440 (N_11440,N_9141,N_8795);
xor U11441 (N_11441,N_9578,N_7602);
or U11442 (N_11442,N_8844,N_9711);
or U11443 (N_11443,N_9811,N_8271);
or U11444 (N_11444,N_9591,N_9057);
xnor U11445 (N_11445,N_9640,N_8160);
and U11446 (N_11446,N_9067,N_8695);
xnor U11447 (N_11447,N_9073,N_9179);
and U11448 (N_11448,N_9946,N_9953);
xor U11449 (N_11449,N_9488,N_8102);
or U11450 (N_11450,N_9680,N_9312);
or U11451 (N_11451,N_8497,N_8708);
nand U11452 (N_11452,N_7721,N_8448);
nand U11453 (N_11453,N_9662,N_7603);
or U11454 (N_11454,N_8297,N_9430);
nor U11455 (N_11455,N_8199,N_9204);
xor U11456 (N_11456,N_9296,N_9857);
xor U11457 (N_11457,N_7654,N_9560);
nand U11458 (N_11458,N_9429,N_8844);
nand U11459 (N_11459,N_8451,N_8839);
nand U11460 (N_11460,N_8693,N_8176);
nand U11461 (N_11461,N_8323,N_8332);
xor U11462 (N_11462,N_9738,N_9329);
and U11463 (N_11463,N_9971,N_9120);
xnor U11464 (N_11464,N_9586,N_8421);
and U11465 (N_11465,N_8207,N_7992);
and U11466 (N_11466,N_8246,N_7700);
and U11467 (N_11467,N_7616,N_9283);
nor U11468 (N_11468,N_9634,N_8095);
or U11469 (N_11469,N_9883,N_8986);
and U11470 (N_11470,N_8335,N_8241);
nor U11471 (N_11471,N_9939,N_9424);
xnor U11472 (N_11472,N_8196,N_9289);
nor U11473 (N_11473,N_9360,N_9974);
xnor U11474 (N_11474,N_8406,N_7562);
nor U11475 (N_11475,N_8319,N_8814);
nand U11476 (N_11476,N_9058,N_8999);
and U11477 (N_11477,N_8155,N_9374);
and U11478 (N_11478,N_8369,N_9794);
xnor U11479 (N_11479,N_9856,N_8536);
nor U11480 (N_11480,N_9257,N_8383);
nor U11481 (N_11481,N_7928,N_9033);
nor U11482 (N_11482,N_8134,N_7620);
and U11483 (N_11483,N_9152,N_7620);
or U11484 (N_11484,N_8662,N_8918);
nor U11485 (N_11485,N_8431,N_8696);
nor U11486 (N_11486,N_7519,N_9498);
nor U11487 (N_11487,N_8191,N_9978);
xnor U11488 (N_11488,N_9393,N_9929);
xor U11489 (N_11489,N_8148,N_8936);
xor U11490 (N_11490,N_9756,N_7774);
or U11491 (N_11491,N_7653,N_7802);
nor U11492 (N_11492,N_9345,N_7733);
or U11493 (N_11493,N_9594,N_8636);
or U11494 (N_11494,N_9670,N_8895);
or U11495 (N_11495,N_8140,N_9783);
and U11496 (N_11496,N_8868,N_8402);
or U11497 (N_11497,N_8822,N_9348);
nor U11498 (N_11498,N_7805,N_7551);
xnor U11499 (N_11499,N_7622,N_9057);
or U11500 (N_11500,N_7997,N_7763);
or U11501 (N_11501,N_8342,N_8190);
xor U11502 (N_11502,N_8266,N_8655);
nor U11503 (N_11503,N_8009,N_9150);
or U11504 (N_11504,N_9517,N_8561);
xor U11505 (N_11505,N_9235,N_9709);
and U11506 (N_11506,N_8464,N_8462);
xor U11507 (N_11507,N_9963,N_8282);
and U11508 (N_11508,N_7521,N_8736);
and U11509 (N_11509,N_7738,N_7979);
nand U11510 (N_11510,N_7932,N_7827);
or U11511 (N_11511,N_8286,N_8087);
nand U11512 (N_11512,N_8279,N_9945);
nor U11513 (N_11513,N_8881,N_8735);
or U11514 (N_11514,N_8013,N_9018);
xnor U11515 (N_11515,N_9831,N_8492);
and U11516 (N_11516,N_9259,N_9719);
or U11517 (N_11517,N_8659,N_9834);
and U11518 (N_11518,N_7752,N_8377);
and U11519 (N_11519,N_8058,N_9050);
or U11520 (N_11520,N_9816,N_9279);
and U11521 (N_11521,N_9441,N_8376);
xnor U11522 (N_11522,N_9353,N_9712);
nand U11523 (N_11523,N_8607,N_9857);
nand U11524 (N_11524,N_9794,N_7954);
or U11525 (N_11525,N_8500,N_8374);
or U11526 (N_11526,N_9837,N_8703);
nand U11527 (N_11527,N_9300,N_7526);
or U11528 (N_11528,N_9049,N_7740);
or U11529 (N_11529,N_9992,N_7834);
nor U11530 (N_11530,N_9642,N_9387);
or U11531 (N_11531,N_9848,N_9291);
nand U11532 (N_11532,N_9182,N_8832);
and U11533 (N_11533,N_9110,N_9146);
and U11534 (N_11534,N_8405,N_7760);
and U11535 (N_11535,N_9583,N_8367);
and U11536 (N_11536,N_9634,N_8830);
xnor U11537 (N_11537,N_7904,N_8001);
xnor U11538 (N_11538,N_9473,N_9131);
nand U11539 (N_11539,N_9579,N_7548);
xor U11540 (N_11540,N_9925,N_8549);
or U11541 (N_11541,N_9265,N_7638);
nor U11542 (N_11542,N_7919,N_7669);
and U11543 (N_11543,N_9265,N_7762);
xnor U11544 (N_11544,N_9959,N_8427);
xnor U11545 (N_11545,N_8900,N_9049);
nand U11546 (N_11546,N_9284,N_9415);
and U11547 (N_11547,N_8947,N_7843);
or U11548 (N_11548,N_7909,N_9775);
or U11549 (N_11549,N_9705,N_7585);
nand U11550 (N_11550,N_8259,N_9240);
or U11551 (N_11551,N_8865,N_8433);
or U11552 (N_11552,N_9639,N_9894);
nor U11553 (N_11553,N_7673,N_8066);
nand U11554 (N_11554,N_9314,N_8733);
xor U11555 (N_11555,N_9463,N_7772);
nor U11556 (N_11556,N_8464,N_9405);
nor U11557 (N_11557,N_9224,N_8548);
nand U11558 (N_11558,N_7831,N_8604);
nand U11559 (N_11559,N_9753,N_7517);
xor U11560 (N_11560,N_9787,N_8439);
or U11561 (N_11561,N_7582,N_9035);
nand U11562 (N_11562,N_7800,N_8593);
nand U11563 (N_11563,N_8642,N_8928);
nor U11564 (N_11564,N_8400,N_8405);
nand U11565 (N_11565,N_9958,N_7575);
nand U11566 (N_11566,N_9858,N_8249);
and U11567 (N_11567,N_9992,N_9526);
nand U11568 (N_11568,N_7733,N_7790);
nand U11569 (N_11569,N_9549,N_8589);
nand U11570 (N_11570,N_9067,N_8575);
nand U11571 (N_11571,N_8570,N_7655);
nor U11572 (N_11572,N_8168,N_8142);
nor U11573 (N_11573,N_8066,N_7975);
nor U11574 (N_11574,N_8870,N_7781);
nor U11575 (N_11575,N_8844,N_7704);
nor U11576 (N_11576,N_8672,N_8469);
and U11577 (N_11577,N_9329,N_8768);
or U11578 (N_11578,N_8174,N_9335);
xor U11579 (N_11579,N_9371,N_9909);
xnor U11580 (N_11580,N_9784,N_7856);
and U11581 (N_11581,N_8582,N_7774);
and U11582 (N_11582,N_8362,N_7505);
or U11583 (N_11583,N_9572,N_8208);
or U11584 (N_11584,N_9546,N_8480);
or U11585 (N_11585,N_7802,N_8100);
or U11586 (N_11586,N_9592,N_9353);
nand U11587 (N_11587,N_7625,N_9259);
xnor U11588 (N_11588,N_8534,N_7558);
xnor U11589 (N_11589,N_8264,N_8400);
or U11590 (N_11590,N_8617,N_8394);
or U11591 (N_11591,N_7650,N_9879);
nand U11592 (N_11592,N_9274,N_9244);
xnor U11593 (N_11593,N_9952,N_9780);
nor U11594 (N_11594,N_8342,N_8058);
and U11595 (N_11595,N_9943,N_8288);
or U11596 (N_11596,N_7966,N_9693);
and U11597 (N_11597,N_9610,N_7943);
or U11598 (N_11598,N_8126,N_9982);
or U11599 (N_11599,N_7858,N_7802);
nand U11600 (N_11600,N_7965,N_7887);
or U11601 (N_11601,N_9484,N_9235);
nor U11602 (N_11602,N_9801,N_7752);
or U11603 (N_11603,N_8113,N_8199);
or U11604 (N_11604,N_9754,N_7778);
nor U11605 (N_11605,N_8235,N_8275);
nor U11606 (N_11606,N_9468,N_7823);
nor U11607 (N_11607,N_9431,N_9469);
nor U11608 (N_11608,N_8685,N_8586);
nor U11609 (N_11609,N_7868,N_9579);
xnor U11610 (N_11610,N_8651,N_9967);
nand U11611 (N_11611,N_8047,N_7970);
and U11612 (N_11612,N_9203,N_8753);
and U11613 (N_11613,N_9256,N_9835);
nor U11614 (N_11614,N_7572,N_9411);
xor U11615 (N_11615,N_9514,N_8301);
xnor U11616 (N_11616,N_8320,N_9787);
xor U11617 (N_11617,N_7500,N_9415);
xor U11618 (N_11618,N_8047,N_8668);
xnor U11619 (N_11619,N_9652,N_9038);
or U11620 (N_11620,N_8398,N_9789);
nor U11621 (N_11621,N_8601,N_8090);
xor U11622 (N_11622,N_9939,N_8594);
and U11623 (N_11623,N_7543,N_9502);
and U11624 (N_11624,N_7718,N_7545);
or U11625 (N_11625,N_8231,N_9215);
nor U11626 (N_11626,N_8187,N_8032);
nand U11627 (N_11627,N_8694,N_9704);
xor U11628 (N_11628,N_9917,N_7649);
and U11629 (N_11629,N_8154,N_9757);
or U11630 (N_11630,N_8206,N_8474);
and U11631 (N_11631,N_7829,N_8910);
nand U11632 (N_11632,N_7963,N_9266);
or U11633 (N_11633,N_8786,N_7500);
and U11634 (N_11634,N_8327,N_7767);
or U11635 (N_11635,N_9963,N_9593);
and U11636 (N_11636,N_8254,N_7649);
nand U11637 (N_11637,N_8853,N_7674);
and U11638 (N_11638,N_8563,N_9965);
and U11639 (N_11639,N_8845,N_8292);
and U11640 (N_11640,N_9083,N_9562);
nand U11641 (N_11641,N_9190,N_7883);
and U11642 (N_11642,N_9327,N_8596);
xor U11643 (N_11643,N_8165,N_9965);
and U11644 (N_11644,N_8759,N_7953);
and U11645 (N_11645,N_7596,N_8460);
xor U11646 (N_11646,N_8560,N_8129);
or U11647 (N_11647,N_8814,N_7501);
nand U11648 (N_11648,N_7811,N_8321);
xor U11649 (N_11649,N_8367,N_8187);
or U11650 (N_11650,N_8049,N_8521);
and U11651 (N_11651,N_9834,N_8074);
xnor U11652 (N_11652,N_7503,N_7954);
xor U11653 (N_11653,N_8753,N_8670);
nor U11654 (N_11654,N_8695,N_8499);
or U11655 (N_11655,N_8537,N_8669);
or U11656 (N_11656,N_9307,N_9781);
nand U11657 (N_11657,N_9532,N_9603);
xnor U11658 (N_11658,N_8891,N_9261);
or U11659 (N_11659,N_7861,N_7936);
or U11660 (N_11660,N_8864,N_8527);
or U11661 (N_11661,N_8671,N_9011);
and U11662 (N_11662,N_9595,N_9740);
or U11663 (N_11663,N_8169,N_7685);
and U11664 (N_11664,N_7784,N_7546);
and U11665 (N_11665,N_7861,N_8949);
xor U11666 (N_11666,N_9078,N_7749);
nand U11667 (N_11667,N_9090,N_7956);
xor U11668 (N_11668,N_7523,N_8823);
or U11669 (N_11669,N_8517,N_9915);
nor U11670 (N_11670,N_9510,N_7502);
nor U11671 (N_11671,N_7724,N_9863);
nand U11672 (N_11672,N_9027,N_7509);
nor U11673 (N_11673,N_7931,N_9889);
xnor U11674 (N_11674,N_8323,N_9069);
and U11675 (N_11675,N_8753,N_8308);
nor U11676 (N_11676,N_7907,N_7652);
nor U11677 (N_11677,N_8018,N_8823);
nand U11678 (N_11678,N_9104,N_8563);
or U11679 (N_11679,N_8681,N_7706);
and U11680 (N_11680,N_9002,N_8409);
or U11681 (N_11681,N_8361,N_7900);
or U11682 (N_11682,N_8254,N_8732);
nand U11683 (N_11683,N_8310,N_8691);
nand U11684 (N_11684,N_8857,N_9350);
xor U11685 (N_11685,N_8883,N_8253);
nand U11686 (N_11686,N_9846,N_7611);
nand U11687 (N_11687,N_9190,N_8858);
nand U11688 (N_11688,N_7851,N_8289);
nor U11689 (N_11689,N_9136,N_9725);
nor U11690 (N_11690,N_8926,N_9900);
nor U11691 (N_11691,N_8478,N_7875);
or U11692 (N_11692,N_8887,N_9168);
xnor U11693 (N_11693,N_7542,N_7937);
and U11694 (N_11694,N_7629,N_8026);
xnor U11695 (N_11695,N_8872,N_8735);
or U11696 (N_11696,N_9031,N_8050);
xor U11697 (N_11697,N_9343,N_7959);
nand U11698 (N_11698,N_7530,N_9117);
or U11699 (N_11699,N_8913,N_9636);
nor U11700 (N_11700,N_8927,N_9070);
xnor U11701 (N_11701,N_8883,N_7907);
xnor U11702 (N_11702,N_9191,N_8527);
xnor U11703 (N_11703,N_8878,N_8996);
xor U11704 (N_11704,N_8703,N_7953);
nor U11705 (N_11705,N_9362,N_9796);
and U11706 (N_11706,N_9045,N_7964);
or U11707 (N_11707,N_8573,N_8476);
nand U11708 (N_11708,N_7755,N_9295);
and U11709 (N_11709,N_9818,N_7512);
nor U11710 (N_11710,N_7621,N_7705);
or U11711 (N_11711,N_9002,N_9658);
xor U11712 (N_11712,N_7788,N_7916);
or U11713 (N_11713,N_9156,N_8365);
and U11714 (N_11714,N_9809,N_8418);
xnor U11715 (N_11715,N_9752,N_7527);
xnor U11716 (N_11716,N_9262,N_8733);
nor U11717 (N_11717,N_8003,N_9269);
nand U11718 (N_11718,N_9286,N_8577);
and U11719 (N_11719,N_7547,N_8527);
nand U11720 (N_11720,N_8349,N_9635);
or U11721 (N_11721,N_9503,N_9931);
or U11722 (N_11722,N_7783,N_9880);
and U11723 (N_11723,N_8731,N_8459);
xnor U11724 (N_11724,N_8012,N_8908);
nor U11725 (N_11725,N_7861,N_7781);
nor U11726 (N_11726,N_9123,N_9973);
or U11727 (N_11727,N_7993,N_7758);
and U11728 (N_11728,N_7947,N_8214);
nor U11729 (N_11729,N_8593,N_7559);
and U11730 (N_11730,N_9947,N_7767);
nor U11731 (N_11731,N_9247,N_9465);
nand U11732 (N_11732,N_8918,N_9441);
xnor U11733 (N_11733,N_7584,N_7827);
or U11734 (N_11734,N_8104,N_9835);
nand U11735 (N_11735,N_8659,N_9686);
nor U11736 (N_11736,N_8096,N_7618);
xor U11737 (N_11737,N_8558,N_8895);
nand U11738 (N_11738,N_8783,N_7787);
nand U11739 (N_11739,N_9213,N_7938);
nand U11740 (N_11740,N_8163,N_7964);
and U11741 (N_11741,N_9338,N_8576);
xor U11742 (N_11742,N_9168,N_9531);
nor U11743 (N_11743,N_9487,N_7691);
or U11744 (N_11744,N_9574,N_8114);
nor U11745 (N_11745,N_9035,N_9642);
xnor U11746 (N_11746,N_7780,N_8746);
nand U11747 (N_11747,N_9659,N_8195);
nand U11748 (N_11748,N_8647,N_8291);
and U11749 (N_11749,N_9673,N_9475);
or U11750 (N_11750,N_7863,N_7836);
or U11751 (N_11751,N_7862,N_8700);
nand U11752 (N_11752,N_9950,N_8479);
and U11753 (N_11753,N_8412,N_8984);
nand U11754 (N_11754,N_8322,N_9874);
xor U11755 (N_11755,N_8159,N_7942);
nor U11756 (N_11756,N_8902,N_8892);
and U11757 (N_11757,N_9728,N_9747);
nand U11758 (N_11758,N_7685,N_7818);
or U11759 (N_11759,N_8743,N_8314);
nor U11760 (N_11760,N_9751,N_7641);
or U11761 (N_11761,N_9794,N_8830);
nand U11762 (N_11762,N_9631,N_9374);
xnor U11763 (N_11763,N_8021,N_8967);
xor U11764 (N_11764,N_7931,N_8017);
and U11765 (N_11765,N_8892,N_8710);
xnor U11766 (N_11766,N_8288,N_7904);
and U11767 (N_11767,N_8932,N_9391);
nand U11768 (N_11768,N_7816,N_8165);
nand U11769 (N_11769,N_8302,N_8766);
and U11770 (N_11770,N_7944,N_7513);
nor U11771 (N_11771,N_9578,N_9434);
nand U11772 (N_11772,N_9849,N_7562);
or U11773 (N_11773,N_7567,N_9939);
and U11774 (N_11774,N_9022,N_8423);
nor U11775 (N_11775,N_9623,N_9654);
nand U11776 (N_11776,N_9836,N_8107);
or U11777 (N_11777,N_8714,N_9778);
xor U11778 (N_11778,N_8704,N_9046);
or U11779 (N_11779,N_9454,N_7974);
and U11780 (N_11780,N_9984,N_7699);
or U11781 (N_11781,N_9746,N_9959);
nor U11782 (N_11782,N_9866,N_8438);
and U11783 (N_11783,N_8753,N_7542);
xor U11784 (N_11784,N_9157,N_8461);
and U11785 (N_11785,N_7886,N_8745);
or U11786 (N_11786,N_7567,N_8080);
nand U11787 (N_11787,N_9793,N_9415);
nor U11788 (N_11788,N_8677,N_8170);
xnor U11789 (N_11789,N_8379,N_9992);
nor U11790 (N_11790,N_7505,N_7968);
nand U11791 (N_11791,N_9135,N_7826);
nand U11792 (N_11792,N_9330,N_9649);
nand U11793 (N_11793,N_8262,N_9448);
nor U11794 (N_11794,N_9898,N_8079);
xnor U11795 (N_11795,N_9823,N_8270);
or U11796 (N_11796,N_8344,N_9509);
nand U11797 (N_11797,N_9892,N_9878);
and U11798 (N_11798,N_8546,N_7738);
nor U11799 (N_11799,N_9042,N_9810);
nor U11800 (N_11800,N_8274,N_8947);
xor U11801 (N_11801,N_8621,N_9654);
xnor U11802 (N_11802,N_8748,N_8836);
xnor U11803 (N_11803,N_7625,N_9386);
and U11804 (N_11804,N_9535,N_9427);
nor U11805 (N_11805,N_9618,N_7886);
nor U11806 (N_11806,N_7627,N_8786);
and U11807 (N_11807,N_9352,N_9516);
or U11808 (N_11808,N_9520,N_8411);
xor U11809 (N_11809,N_7875,N_9093);
nand U11810 (N_11810,N_9742,N_9938);
xnor U11811 (N_11811,N_9374,N_9250);
nand U11812 (N_11812,N_8953,N_9137);
nor U11813 (N_11813,N_9635,N_8171);
xor U11814 (N_11814,N_7908,N_9218);
or U11815 (N_11815,N_9223,N_7704);
nand U11816 (N_11816,N_9568,N_9024);
nand U11817 (N_11817,N_9865,N_9790);
xnor U11818 (N_11818,N_9453,N_8888);
nor U11819 (N_11819,N_9343,N_8355);
and U11820 (N_11820,N_8304,N_9917);
nand U11821 (N_11821,N_9714,N_8840);
nor U11822 (N_11822,N_7577,N_8360);
xnor U11823 (N_11823,N_8321,N_9850);
nand U11824 (N_11824,N_8821,N_8812);
nor U11825 (N_11825,N_7745,N_7930);
nand U11826 (N_11826,N_9844,N_9359);
and U11827 (N_11827,N_8600,N_8867);
or U11828 (N_11828,N_9758,N_8340);
nor U11829 (N_11829,N_8962,N_9459);
or U11830 (N_11830,N_8777,N_7590);
nand U11831 (N_11831,N_8809,N_7817);
nor U11832 (N_11832,N_9155,N_8680);
and U11833 (N_11833,N_8880,N_9192);
and U11834 (N_11834,N_9406,N_9408);
and U11835 (N_11835,N_8668,N_8547);
or U11836 (N_11836,N_7648,N_8488);
and U11837 (N_11837,N_7644,N_8452);
and U11838 (N_11838,N_9369,N_8797);
or U11839 (N_11839,N_8131,N_9989);
and U11840 (N_11840,N_8372,N_9282);
nand U11841 (N_11841,N_8113,N_8502);
nor U11842 (N_11842,N_7938,N_9615);
nand U11843 (N_11843,N_7768,N_8436);
and U11844 (N_11844,N_7964,N_9862);
nand U11845 (N_11845,N_9448,N_8878);
nand U11846 (N_11846,N_9117,N_7604);
and U11847 (N_11847,N_9261,N_8122);
or U11848 (N_11848,N_8840,N_7690);
and U11849 (N_11849,N_8786,N_9551);
xnor U11850 (N_11850,N_7943,N_9286);
or U11851 (N_11851,N_7864,N_8000);
nand U11852 (N_11852,N_8172,N_7504);
or U11853 (N_11853,N_9874,N_8885);
or U11854 (N_11854,N_7861,N_9032);
xor U11855 (N_11855,N_7773,N_9715);
nand U11856 (N_11856,N_7544,N_7666);
xor U11857 (N_11857,N_7986,N_7732);
xnor U11858 (N_11858,N_9968,N_9272);
nor U11859 (N_11859,N_8196,N_7768);
and U11860 (N_11860,N_9258,N_7649);
nor U11861 (N_11861,N_8203,N_8103);
nand U11862 (N_11862,N_8555,N_7914);
and U11863 (N_11863,N_8742,N_7958);
and U11864 (N_11864,N_9906,N_9505);
nor U11865 (N_11865,N_8037,N_8992);
or U11866 (N_11866,N_9451,N_8238);
nand U11867 (N_11867,N_8215,N_8594);
and U11868 (N_11868,N_8969,N_9065);
and U11869 (N_11869,N_7832,N_8180);
xnor U11870 (N_11870,N_9667,N_9221);
xnor U11871 (N_11871,N_9924,N_9717);
and U11872 (N_11872,N_7731,N_8982);
or U11873 (N_11873,N_9737,N_8075);
nor U11874 (N_11874,N_7997,N_8617);
nand U11875 (N_11875,N_8344,N_9131);
and U11876 (N_11876,N_9618,N_7803);
nor U11877 (N_11877,N_9177,N_9241);
xor U11878 (N_11878,N_7828,N_9108);
nand U11879 (N_11879,N_8658,N_8302);
nand U11880 (N_11880,N_9751,N_9626);
or U11881 (N_11881,N_9016,N_7584);
and U11882 (N_11882,N_7991,N_8075);
nor U11883 (N_11883,N_8831,N_7704);
and U11884 (N_11884,N_9352,N_7564);
or U11885 (N_11885,N_7882,N_9248);
and U11886 (N_11886,N_9098,N_8433);
and U11887 (N_11887,N_8634,N_8769);
or U11888 (N_11888,N_8922,N_8668);
xnor U11889 (N_11889,N_8177,N_7944);
nand U11890 (N_11890,N_9919,N_8935);
or U11891 (N_11891,N_9150,N_9605);
xor U11892 (N_11892,N_8228,N_7998);
nor U11893 (N_11893,N_8079,N_8784);
xor U11894 (N_11894,N_8630,N_7851);
nand U11895 (N_11895,N_7624,N_7640);
and U11896 (N_11896,N_9500,N_8896);
or U11897 (N_11897,N_9244,N_8947);
nand U11898 (N_11898,N_8076,N_7520);
or U11899 (N_11899,N_8025,N_9514);
xnor U11900 (N_11900,N_7637,N_8747);
xnor U11901 (N_11901,N_8944,N_9663);
or U11902 (N_11902,N_9536,N_8426);
and U11903 (N_11903,N_7694,N_8987);
and U11904 (N_11904,N_8972,N_8049);
and U11905 (N_11905,N_7660,N_9984);
nor U11906 (N_11906,N_7740,N_8729);
nand U11907 (N_11907,N_9545,N_7911);
nand U11908 (N_11908,N_7551,N_8066);
and U11909 (N_11909,N_8635,N_8748);
and U11910 (N_11910,N_7533,N_9621);
or U11911 (N_11911,N_7590,N_8712);
nor U11912 (N_11912,N_9464,N_9194);
and U11913 (N_11913,N_9480,N_9248);
xor U11914 (N_11914,N_7770,N_8100);
nand U11915 (N_11915,N_7744,N_8452);
nor U11916 (N_11916,N_8814,N_8535);
nand U11917 (N_11917,N_8956,N_8127);
nand U11918 (N_11918,N_7661,N_8451);
nand U11919 (N_11919,N_9975,N_9295);
and U11920 (N_11920,N_7878,N_8275);
nor U11921 (N_11921,N_7808,N_8288);
or U11922 (N_11922,N_9976,N_7853);
xnor U11923 (N_11923,N_8443,N_9424);
xnor U11924 (N_11924,N_9602,N_7938);
nand U11925 (N_11925,N_8209,N_9621);
nor U11926 (N_11926,N_9748,N_8689);
or U11927 (N_11927,N_9457,N_9687);
or U11928 (N_11928,N_8934,N_7597);
and U11929 (N_11929,N_7885,N_8732);
and U11930 (N_11930,N_9564,N_9249);
xnor U11931 (N_11931,N_7526,N_7548);
xnor U11932 (N_11932,N_8389,N_8090);
xor U11933 (N_11933,N_9759,N_8305);
nand U11934 (N_11934,N_8301,N_8306);
or U11935 (N_11935,N_8423,N_7635);
nand U11936 (N_11936,N_8432,N_7563);
or U11937 (N_11937,N_7628,N_9310);
and U11938 (N_11938,N_8081,N_7591);
or U11939 (N_11939,N_9863,N_9105);
nand U11940 (N_11940,N_9323,N_9450);
or U11941 (N_11941,N_9994,N_8781);
and U11942 (N_11942,N_8926,N_9687);
or U11943 (N_11943,N_9081,N_9838);
nand U11944 (N_11944,N_8760,N_9389);
and U11945 (N_11945,N_8618,N_9615);
nand U11946 (N_11946,N_8114,N_8675);
nand U11947 (N_11947,N_8141,N_9882);
nor U11948 (N_11948,N_8120,N_8720);
nor U11949 (N_11949,N_7825,N_7682);
nand U11950 (N_11950,N_9796,N_9193);
or U11951 (N_11951,N_9558,N_9340);
nor U11952 (N_11952,N_8443,N_8913);
or U11953 (N_11953,N_9595,N_8158);
or U11954 (N_11954,N_9570,N_8036);
nor U11955 (N_11955,N_8894,N_9996);
nand U11956 (N_11956,N_9114,N_7909);
or U11957 (N_11957,N_7630,N_9455);
nand U11958 (N_11958,N_9383,N_8270);
or U11959 (N_11959,N_9142,N_9528);
nor U11960 (N_11960,N_7814,N_9169);
nor U11961 (N_11961,N_7639,N_8618);
xor U11962 (N_11962,N_7970,N_9856);
nand U11963 (N_11963,N_9388,N_7994);
nor U11964 (N_11964,N_8646,N_9587);
xnor U11965 (N_11965,N_8299,N_7976);
xor U11966 (N_11966,N_9286,N_8179);
nor U11967 (N_11967,N_8037,N_9117);
or U11968 (N_11968,N_8990,N_9936);
or U11969 (N_11969,N_9488,N_8756);
nor U11970 (N_11970,N_9549,N_9882);
nor U11971 (N_11971,N_8091,N_9604);
and U11972 (N_11972,N_9484,N_7821);
nand U11973 (N_11973,N_8397,N_9035);
or U11974 (N_11974,N_7919,N_7521);
nand U11975 (N_11975,N_7873,N_9880);
or U11976 (N_11976,N_8883,N_8401);
xnor U11977 (N_11977,N_9023,N_8472);
or U11978 (N_11978,N_9231,N_7598);
xnor U11979 (N_11979,N_9045,N_9165);
nor U11980 (N_11980,N_7681,N_9811);
xnor U11981 (N_11981,N_9759,N_9127);
xor U11982 (N_11982,N_8802,N_8979);
nand U11983 (N_11983,N_8969,N_7889);
xor U11984 (N_11984,N_8526,N_8350);
and U11985 (N_11985,N_7659,N_9877);
nor U11986 (N_11986,N_8740,N_9579);
or U11987 (N_11987,N_9936,N_9093);
or U11988 (N_11988,N_9331,N_9702);
nand U11989 (N_11989,N_8984,N_7828);
and U11990 (N_11990,N_7735,N_8681);
nand U11991 (N_11991,N_7511,N_9241);
xnor U11992 (N_11992,N_7766,N_8095);
nor U11993 (N_11993,N_9444,N_9380);
nand U11994 (N_11994,N_8815,N_9624);
or U11995 (N_11995,N_9878,N_7995);
nor U11996 (N_11996,N_7799,N_7789);
and U11997 (N_11997,N_9755,N_9067);
or U11998 (N_11998,N_9851,N_8858);
nand U11999 (N_11999,N_9160,N_8228);
nor U12000 (N_12000,N_9133,N_8187);
nor U12001 (N_12001,N_9149,N_8922);
or U12002 (N_12002,N_9453,N_8261);
nor U12003 (N_12003,N_9194,N_8687);
or U12004 (N_12004,N_9492,N_8118);
and U12005 (N_12005,N_9511,N_9286);
or U12006 (N_12006,N_8305,N_7876);
xnor U12007 (N_12007,N_8727,N_9431);
nor U12008 (N_12008,N_9656,N_8853);
and U12009 (N_12009,N_9385,N_9715);
xor U12010 (N_12010,N_7514,N_9881);
nor U12011 (N_12011,N_9927,N_8606);
nor U12012 (N_12012,N_9019,N_8577);
nor U12013 (N_12013,N_8479,N_8585);
and U12014 (N_12014,N_9988,N_7580);
nand U12015 (N_12015,N_8466,N_9570);
and U12016 (N_12016,N_9364,N_7627);
and U12017 (N_12017,N_8970,N_9667);
nand U12018 (N_12018,N_7591,N_7717);
and U12019 (N_12019,N_8214,N_9270);
nand U12020 (N_12020,N_9792,N_8210);
nor U12021 (N_12021,N_9212,N_7727);
xor U12022 (N_12022,N_9761,N_7530);
or U12023 (N_12023,N_7734,N_8957);
nand U12024 (N_12024,N_8365,N_9864);
xnor U12025 (N_12025,N_9792,N_9023);
and U12026 (N_12026,N_7599,N_9527);
or U12027 (N_12027,N_7810,N_9589);
nand U12028 (N_12028,N_9531,N_8135);
or U12029 (N_12029,N_8341,N_9355);
and U12030 (N_12030,N_8317,N_9876);
nor U12031 (N_12031,N_8484,N_7578);
and U12032 (N_12032,N_7857,N_9344);
nor U12033 (N_12033,N_8457,N_7528);
or U12034 (N_12034,N_9108,N_8979);
or U12035 (N_12035,N_8169,N_8473);
and U12036 (N_12036,N_7969,N_7583);
nor U12037 (N_12037,N_8270,N_8838);
nand U12038 (N_12038,N_7676,N_8103);
xnor U12039 (N_12039,N_7761,N_9692);
and U12040 (N_12040,N_7786,N_9626);
nand U12041 (N_12041,N_9116,N_9571);
and U12042 (N_12042,N_8856,N_9805);
or U12043 (N_12043,N_9458,N_8101);
nand U12044 (N_12044,N_9640,N_7659);
nor U12045 (N_12045,N_9103,N_8843);
and U12046 (N_12046,N_9952,N_9696);
and U12047 (N_12047,N_8438,N_9017);
nand U12048 (N_12048,N_8122,N_9050);
nor U12049 (N_12049,N_7502,N_8177);
nand U12050 (N_12050,N_9072,N_8002);
and U12051 (N_12051,N_7587,N_8510);
nand U12052 (N_12052,N_8565,N_7731);
xnor U12053 (N_12053,N_9367,N_7990);
nand U12054 (N_12054,N_8644,N_8887);
or U12055 (N_12055,N_9190,N_9878);
xnor U12056 (N_12056,N_8473,N_7722);
and U12057 (N_12057,N_8670,N_8289);
nor U12058 (N_12058,N_9684,N_8520);
nand U12059 (N_12059,N_9797,N_7682);
xnor U12060 (N_12060,N_7743,N_7639);
nand U12061 (N_12061,N_9154,N_8467);
or U12062 (N_12062,N_9042,N_7686);
or U12063 (N_12063,N_8733,N_9900);
and U12064 (N_12064,N_9748,N_9364);
nor U12065 (N_12065,N_7933,N_7735);
nor U12066 (N_12066,N_8266,N_9745);
and U12067 (N_12067,N_9314,N_7760);
nor U12068 (N_12068,N_9885,N_9228);
and U12069 (N_12069,N_8177,N_8217);
nor U12070 (N_12070,N_8796,N_7532);
and U12071 (N_12071,N_9162,N_9793);
nor U12072 (N_12072,N_9875,N_9259);
and U12073 (N_12073,N_8754,N_9143);
xnor U12074 (N_12074,N_7516,N_8498);
nor U12075 (N_12075,N_9610,N_9020);
nand U12076 (N_12076,N_7816,N_9400);
nand U12077 (N_12077,N_8305,N_9571);
or U12078 (N_12078,N_8988,N_8693);
nor U12079 (N_12079,N_9724,N_9281);
xnor U12080 (N_12080,N_7863,N_9829);
xnor U12081 (N_12081,N_9959,N_7711);
and U12082 (N_12082,N_7890,N_9858);
nor U12083 (N_12083,N_8653,N_9194);
nand U12084 (N_12084,N_9289,N_9095);
nand U12085 (N_12085,N_7878,N_8677);
nand U12086 (N_12086,N_8331,N_7591);
nor U12087 (N_12087,N_9100,N_8226);
and U12088 (N_12088,N_7524,N_9222);
and U12089 (N_12089,N_8397,N_9351);
nand U12090 (N_12090,N_9424,N_9258);
nor U12091 (N_12091,N_8840,N_9580);
and U12092 (N_12092,N_9079,N_7514);
or U12093 (N_12093,N_7829,N_9239);
xor U12094 (N_12094,N_8306,N_8429);
nand U12095 (N_12095,N_7723,N_9955);
nor U12096 (N_12096,N_9030,N_7755);
xor U12097 (N_12097,N_9271,N_7576);
xor U12098 (N_12098,N_8655,N_9847);
or U12099 (N_12099,N_8876,N_9973);
nand U12100 (N_12100,N_8684,N_8775);
nor U12101 (N_12101,N_9654,N_9747);
or U12102 (N_12102,N_8798,N_9988);
xnor U12103 (N_12103,N_9138,N_7972);
xnor U12104 (N_12104,N_7772,N_9679);
nand U12105 (N_12105,N_9192,N_7980);
nand U12106 (N_12106,N_8689,N_8760);
and U12107 (N_12107,N_7523,N_9894);
xor U12108 (N_12108,N_9055,N_8918);
or U12109 (N_12109,N_9341,N_8635);
nor U12110 (N_12110,N_8074,N_9911);
nor U12111 (N_12111,N_7573,N_9181);
nand U12112 (N_12112,N_8294,N_9612);
nand U12113 (N_12113,N_9156,N_8590);
xnor U12114 (N_12114,N_8822,N_7975);
xor U12115 (N_12115,N_9643,N_9382);
or U12116 (N_12116,N_8472,N_9707);
or U12117 (N_12117,N_9366,N_8067);
nand U12118 (N_12118,N_7717,N_9126);
or U12119 (N_12119,N_8525,N_9391);
and U12120 (N_12120,N_9907,N_9069);
xnor U12121 (N_12121,N_8139,N_7729);
nor U12122 (N_12122,N_9441,N_7789);
nor U12123 (N_12123,N_9947,N_9100);
nand U12124 (N_12124,N_8370,N_9906);
or U12125 (N_12125,N_8117,N_8493);
and U12126 (N_12126,N_9909,N_8099);
nand U12127 (N_12127,N_9401,N_8338);
and U12128 (N_12128,N_8604,N_9082);
or U12129 (N_12129,N_9318,N_9881);
nor U12130 (N_12130,N_8143,N_8991);
nand U12131 (N_12131,N_8208,N_8069);
xor U12132 (N_12132,N_8135,N_7746);
xor U12133 (N_12133,N_9709,N_8450);
nand U12134 (N_12134,N_7690,N_7580);
xor U12135 (N_12135,N_8845,N_9419);
and U12136 (N_12136,N_8238,N_8857);
nand U12137 (N_12137,N_9629,N_7573);
or U12138 (N_12138,N_7585,N_9691);
or U12139 (N_12139,N_9149,N_8792);
and U12140 (N_12140,N_8026,N_8547);
nand U12141 (N_12141,N_9786,N_8259);
and U12142 (N_12142,N_8142,N_7649);
nand U12143 (N_12143,N_7515,N_7911);
nand U12144 (N_12144,N_7637,N_8079);
or U12145 (N_12145,N_8986,N_8177);
nor U12146 (N_12146,N_8063,N_9516);
or U12147 (N_12147,N_7779,N_7620);
and U12148 (N_12148,N_7930,N_8156);
xor U12149 (N_12149,N_8648,N_7986);
nor U12150 (N_12150,N_7540,N_7806);
and U12151 (N_12151,N_8892,N_7752);
nor U12152 (N_12152,N_9485,N_8554);
and U12153 (N_12153,N_9479,N_8981);
nand U12154 (N_12154,N_8003,N_9939);
nor U12155 (N_12155,N_8854,N_9213);
nor U12156 (N_12156,N_7823,N_8568);
nand U12157 (N_12157,N_8261,N_8537);
nand U12158 (N_12158,N_9829,N_8433);
nor U12159 (N_12159,N_9093,N_9227);
xor U12160 (N_12160,N_8379,N_9821);
xor U12161 (N_12161,N_8899,N_9920);
nand U12162 (N_12162,N_7715,N_9410);
or U12163 (N_12163,N_9086,N_9081);
or U12164 (N_12164,N_9852,N_8288);
and U12165 (N_12165,N_8623,N_9881);
nor U12166 (N_12166,N_8010,N_9251);
nor U12167 (N_12167,N_7777,N_8632);
nor U12168 (N_12168,N_8817,N_8664);
nor U12169 (N_12169,N_8076,N_8581);
or U12170 (N_12170,N_9351,N_8021);
xnor U12171 (N_12171,N_8434,N_8083);
xnor U12172 (N_12172,N_9144,N_9247);
nand U12173 (N_12173,N_9847,N_9037);
or U12174 (N_12174,N_7832,N_7888);
or U12175 (N_12175,N_8000,N_7597);
xnor U12176 (N_12176,N_7704,N_8840);
nor U12177 (N_12177,N_9399,N_8475);
and U12178 (N_12178,N_9114,N_8006);
nand U12179 (N_12179,N_9540,N_8997);
or U12180 (N_12180,N_9541,N_9517);
and U12181 (N_12181,N_9555,N_9883);
nor U12182 (N_12182,N_9011,N_9533);
xnor U12183 (N_12183,N_7984,N_8999);
xnor U12184 (N_12184,N_7991,N_9491);
and U12185 (N_12185,N_8587,N_9429);
or U12186 (N_12186,N_8894,N_7645);
nor U12187 (N_12187,N_8880,N_8069);
nor U12188 (N_12188,N_8136,N_8014);
and U12189 (N_12189,N_9206,N_9189);
and U12190 (N_12190,N_8241,N_9337);
or U12191 (N_12191,N_9277,N_7796);
nor U12192 (N_12192,N_9351,N_7617);
nand U12193 (N_12193,N_9606,N_7651);
nor U12194 (N_12194,N_8653,N_7716);
nand U12195 (N_12195,N_9025,N_7720);
nor U12196 (N_12196,N_7676,N_7924);
and U12197 (N_12197,N_9626,N_9969);
and U12198 (N_12198,N_9639,N_8719);
nor U12199 (N_12199,N_8500,N_9658);
nor U12200 (N_12200,N_8654,N_8299);
nor U12201 (N_12201,N_7861,N_9578);
xnor U12202 (N_12202,N_9949,N_9454);
nor U12203 (N_12203,N_8020,N_8443);
or U12204 (N_12204,N_7532,N_8658);
and U12205 (N_12205,N_9343,N_8236);
and U12206 (N_12206,N_8558,N_8419);
or U12207 (N_12207,N_7899,N_8586);
and U12208 (N_12208,N_9268,N_7727);
nor U12209 (N_12209,N_7714,N_8636);
or U12210 (N_12210,N_9399,N_8500);
nand U12211 (N_12211,N_8547,N_8591);
xnor U12212 (N_12212,N_9886,N_8497);
and U12213 (N_12213,N_9073,N_8595);
nor U12214 (N_12214,N_8300,N_8376);
xnor U12215 (N_12215,N_8767,N_8182);
or U12216 (N_12216,N_9019,N_7592);
nor U12217 (N_12217,N_9469,N_8827);
xnor U12218 (N_12218,N_7867,N_8288);
nand U12219 (N_12219,N_8615,N_7509);
nor U12220 (N_12220,N_9573,N_8070);
nand U12221 (N_12221,N_8759,N_9244);
xnor U12222 (N_12222,N_8199,N_8909);
nor U12223 (N_12223,N_8183,N_9439);
xnor U12224 (N_12224,N_7769,N_8365);
and U12225 (N_12225,N_8724,N_8336);
or U12226 (N_12226,N_8720,N_9958);
or U12227 (N_12227,N_9082,N_9171);
nand U12228 (N_12228,N_9267,N_7527);
or U12229 (N_12229,N_8643,N_9337);
or U12230 (N_12230,N_9021,N_8849);
xor U12231 (N_12231,N_8976,N_9401);
or U12232 (N_12232,N_8459,N_9541);
nand U12233 (N_12233,N_8882,N_9706);
or U12234 (N_12234,N_8039,N_7991);
nor U12235 (N_12235,N_8079,N_7658);
or U12236 (N_12236,N_9702,N_9973);
xor U12237 (N_12237,N_9095,N_9049);
nand U12238 (N_12238,N_8719,N_8730);
nand U12239 (N_12239,N_9036,N_8578);
nor U12240 (N_12240,N_9411,N_8126);
nand U12241 (N_12241,N_8872,N_8609);
and U12242 (N_12242,N_7855,N_8267);
xor U12243 (N_12243,N_7813,N_8445);
nand U12244 (N_12244,N_8605,N_8246);
and U12245 (N_12245,N_8899,N_9179);
nor U12246 (N_12246,N_7681,N_7966);
nand U12247 (N_12247,N_7796,N_7726);
and U12248 (N_12248,N_8130,N_8973);
and U12249 (N_12249,N_9995,N_8716);
or U12250 (N_12250,N_9589,N_9437);
or U12251 (N_12251,N_8944,N_7619);
and U12252 (N_12252,N_8398,N_9521);
or U12253 (N_12253,N_8904,N_9047);
nor U12254 (N_12254,N_8573,N_9514);
nor U12255 (N_12255,N_8145,N_7776);
xnor U12256 (N_12256,N_9892,N_8323);
nand U12257 (N_12257,N_8595,N_8209);
xnor U12258 (N_12258,N_8279,N_9963);
nor U12259 (N_12259,N_9979,N_9287);
or U12260 (N_12260,N_9418,N_7627);
nor U12261 (N_12261,N_7748,N_8204);
nand U12262 (N_12262,N_9270,N_8366);
nor U12263 (N_12263,N_7720,N_9914);
and U12264 (N_12264,N_8545,N_9704);
xnor U12265 (N_12265,N_8367,N_9080);
xor U12266 (N_12266,N_9247,N_9127);
nor U12267 (N_12267,N_7556,N_9105);
nor U12268 (N_12268,N_9654,N_8545);
nand U12269 (N_12269,N_9580,N_7815);
and U12270 (N_12270,N_9722,N_9835);
nand U12271 (N_12271,N_7865,N_9473);
and U12272 (N_12272,N_9072,N_7582);
nand U12273 (N_12273,N_9501,N_9565);
and U12274 (N_12274,N_8072,N_9027);
xnor U12275 (N_12275,N_9145,N_8181);
and U12276 (N_12276,N_8148,N_8069);
nor U12277 (N_12277,N_9350,N_7652);
xor U12278 (N_12278,N_8569,N_9315);
xnor U12279 (N_12279,N_8088,N_7932);
nand U12280 (N_12280,N_9108,N_8749);
nor U12281 (N_12281,N_9774,N_7926);
xor U12282 (N_12282,N_8187,N_9603);
nor U12283 (N_12283,N_9121,N_8888);
xor U12284 (N_12284,N_8307,N_8831);
nand U12285 (N_12285,N_8409,N_9257);
nand U12286 (N_12286,N_8622,N_9232);
nand U12287 (N_12287,N_9742,N_7652);
and U12288 (N_12288,N_9619,N_8990);
and U12289 (N_12289,N_8781,N_9351);
and U12290 (N_12290,N_9036,N_8615);
or U12291 (N_12291,N_8149,N_9134);
nor U12292 (N_12292,N_9367,N_7659);
xnor U12293 (N_12293,N_9991,N_8410);
xnor U12294 (N_12294,N_8307,N_8504);
or U12295 (N_12295,N_9818,N_8728);
xor U12296 (N_12296,N_9029,N_9266);
nor U12297 (N_12297,N_7719,N_9370);
and U12298 (N_12298,N_9105,N_9237);
xnor U12299 (N_12299,N_9551,N_9518);
nor U12300 (N_12300,N_9894,N_9859);
nor U12301 (N_12301,N_7608,N_9712);
or U12302 (N_12302,N_8841,N_7918);
xnor U12303 (N_12303,N_7887,N_8688);
nand U12304 (N_12304,N_9138,N_8188);
nor U12305 (N_12305,N_7912,N_9823);
nand U12306 (N_12306,N_9502,N_8557);
or U12307 (N_12307,N_8116,N_9108);
or U12308 (N_12308,N_8110,N_7645);
nor U12309 (N_12309,N_8561,N_9146);
nor U12310 (N_12310,N_9608,N_8187);
and U12311 (N_12311,N_7624,N_7632);
xor U12312 (N_12312,N_9643,N_7521);
and U12313 (N_12313,N_8999,N_9266);
nand U12314 (N_12314,N_9748,N_9243);
nand U12315 (N_12315,N_7843,N_9172);
nor U12316 (N_12316,N_9360,N_8225);
nor U12317 (N_12317,N_9756,N_7556);
nor U12318 (N_12318,N_8893,N_8030);
and U12319 (N_12319,N_7949,N_8388);
nor U12320 (N_12320,N_7692,N_9354);
or U12321 (N_12321,N_7886,N_8846);
nor U12322 (N_12322,N_8102,N_8644);
xnor U12323 (N_12323,N_8458,N_7514);
or U12324 (N_12324,N_8413,N_7563);
and U12325 (N_12325,N_8172,N_8334);
xor U12326 (N_12326,N_8370,N_8693);
xor U12327 (N_12327,N_8976,N_8864);
xor U12328 (N_12328,N_7967,N_8431);
xor U12329 (N_12329,N_9130,N_9421);
nand U12330 (N_12330,N_8316,N_8309);
and U12331 (N_12331,N_8514,N_9072);
and U12332 (N_12332,N_9828,N_7929);
and U12333 (N_12333,N_8961,N_9048);
nor U12334 (N_12334,N_8878,N_8934);
nand U12335 (N_12335,N_8303,N_9474);
xor U12336 (N_12336,N_7828,N_7993);
xnor U12337 (N_12337,N_8416,N_9143);
and U12338 (N_12338,N_9728,N_9229);
nand U12339 (N_12339,N_8847,N_7884);
or U12340 (N_12340,N_7611,N_9087);
xnor U12341 (N_12341,N_8767,N_9519);
nor U12342 (N_12342,N_7906,N_9067);
or U12343 (N_12343,N_9194,N_8954);
or U12344 (N_12344,N_9025,N_7639);
nor U12345 (N_12345,N_9914,N_9946);
or U12346 (N_12346,N_7837,N_8927);
xnor U12347 (N_12347,N_8852,N_7914);
nor U12348 (N_12348,N_9043,N_8771);
xor U12349 (N_12349,N_9317,N_9009);
and U12350 (N_12350,N_9768,N_8272);
nor U12351 (N_12351,N_8537,N_8532);
nor U12352 (N_12352,N_8931,N_7955);
or U12353 (N_12353,N_8411,N_8730);
or U12354 (N_12354,N_7895,N_8609);
xor U12355 (N_12355,N_7503,N_8974);
xor U12356 (N_12356,N_7767,N_9498);
and U12357 (N_12357,N_8408,N_7916);
nand U12358 (N_12358,N_8638,N_8601);
xor U12359 (N_12359,N_9185,N_8995);
or U12360 (N_12360,N_8773,N_9022);
or U12361 (N_12361,N_9687,N_9810);
and U12362 (N_12362,N_8279,N_9316);
nor U12363 (N_12363,N_9793,N_8970);
nor U12364 (N_12364,N_8214,N_7512);
or U12365 (N_12365,N_7938,N_7841);
nand U12366 (N_12366,N_8989,N_9086);
xnor U12367 (N_12367,N_8189,N_8805);
and U12368 (N_12368,N_8362,N_9693);
and U12369 (N_12369,N_8611,N_7860);
nand U12370 (N_12370,N_7974,N_8535);
or U12371 (N_12371,N_9867,N_8943);
xnor U12372 (N_12372,N_9682,N_8907);
xor U12373 (N_12373,N_9811,N_9889);
xnor U12374 (N_12374,N_9581,N_8382);
xor U12375 (N_12375,N_7548,N_7707);
nand U12376 (N_12376,N_9288,N_8657);
nand U12377 (N_12377,N_9734,N_8586);
xnor U12378 (N_12378,N_9361,N_9352);
and U12379 (N_12379,N_8498,N_8466);
nor U12380 (N_12380,N_8740,N_9054);
xnor U12381 (N_12381,N_7838,N_8536);
xor U12382 (N_12382,N_7832,N_8034);
or U12383 (N_12383,N_9972,N_9784);
and U12384 (N_12384,N_9348,N_9580);
and U12385 (N_12385,N_8899,N_8713);
or U12386 (N_12386,N_7958,N_7756);
or U12387 (N_12387,N_8525,N_9589);
nor U12388 (N_12388,N_8160,N_7656);
and U12389 (N_12389,N_9614,N_8769);
or U12390 (N_12390,N_9644,N_8867);
nand U12391 (N_12391,N_8878,N_8401);
nor U12392 (N_12392,N_8916,N_8409);
or U12393 (N_12393,N_7630,N_9508);
and U12394 (N_12394,N_7961,N_8603);
or U12395 (N_12395,N_8431,N_8773);
nor U12396 (N_12396,N_9209,N_8106);
nor U12397 (N_12397,N_8196,N_8234);
and U12398 (N_12398,N_9243,N_9608);
nor U12399 (N_12399,N_8132,N_8787);
and U12400 (N_12400,N_8202,N_9784);
and U12401 (N_12401,N_8930,N_7674);
or U12402 (N_12402,N_7949,N_9723);
nand U12403 (N_12403,N_8928,N_8998);
xor U12404 (N_12404,N_7764,N_9096);
or U12405 (N_12405,N_7718,N_9978);
xor U12406 (N_12406,N_7776,N_8428);
nor U12407 (N_12407,N_8829,N_8700);
or U12408 (N_12408,N_8504,N_7903);
xor U12409 (N_12409,N_7573,N_8961);
nor U12410 (N_12410,N_9041,N_8833);
or U12411 (N_12411,N_7968,N_9887);
and U12412 (N_12412,N_7545,N_9836);
and U12413 (N_12413,N_9356,N_7562);
or U12414 (N_12414,N_8816,N_8125);
and U12415 (N_12415,N_7976,N_9445);
nor U12416 (N_12416,N_8118,N_9187);
and U12417 (N_12417,N_9360,N_7998);
nor U12418 (N_12418,N_7722,N_7913);
or U12419 (N_12419,N_8971,N_7546);
nand U12420 (N_12420,N_7791,N_9607);
nor U12421 (N_12421,N_9286,N_9631);
and U12422 (N_12422,N_8805,N_9505);
xor U12423 (N_12423,N_9233,N_8149);
and U12424 (N_12424,N_9427,N_9937);
nand U12425 (N_12425,N_9568,N_8782);
nand U12426 (N_12426,N_8774,N_8986);
nand U12427 (N_12427,N_7848,N_8573);
nand U12428 (N_12428,N_8346,N_8830);
xor U12429 (N_12429,N_7670,N_9505);
nor U12430 (N_12430,N_9574,N_9339);
and U12431 (N_12431,N_8162,N_9076);
nor U12432 (N_12432,N_8638,N_9367);
xor U12433 (N_12433,N_7642,N_8063);
and U12434 (N_12434,N_7591,N_8495);
nand U12435 (N_12435,N_9529,N_8636);
nor U12436 (N_12436,N_8603,N_8259);
xor U12437 (N_12437,N_9825,N_9983);
or U12438 (N_12438,N_8233,N_8446);
xor U12439 (N_12439,N_9942,N_7893);
xnor U12440 (N_12440,N_8907,N_8614);
nor U12441 (N_12441,N_7982,N_9604);
xnor U12442 (N_12442,N_7827,N_7943);
nor U12443 (N_12443,N_8980,N_8352);
or U12444 (N_12444,N_9164,N_9385);
xnor U12445 (N_12445,N_8699,N_9641);
and U12446 (N_12446,N_8336,N_8445);
nor U12447 (N_12447,N_9528,N_9515);
nand U12448 (N_12448,N_9914,N_9169);
nor U12449 (N_12449,N_9530,N_8766);
nand U12450 (N_12450,N_8248,N_9005);
nand U12451 (N_12451,N_8732,N_8507);
or U12452 (N_12452,N_9439,N_9978);
or U12453 (N_12453,N_9477,N_8291);
or U12454 (N_12454,N_7980,N_9023);
or U12455 (N_12455,N_9771,N_9673);
nor U12456 (N_12456,N_8427,N_8597);
or U12457 (N_12457,N_8032,N_9817);
or U12458 (N_12458,N_8149,N_8625);
xor U12459 (N_12459,N_9595,N_7821);
or U12460 (N_12460,N_9544,N_8329);
nand U12461 (N_12461,N_9875,N_8285);
nor U12462 (N_12462,N_7869,N_9012);
nand U12463 (N_12463,N_7527,N_8100);
or U12464 (N_12464,N_8605,N_8914);
nor U12465 (N_12465,N_9673,N_9885);
xor U12466 (N_12466,N_9631,N_7974);
or U12467 (N_12467,N_8030,N_8739);
nor U12468 (N_12468,N_8163,N_9939);
nand U12469 (N_12469,N_9310,N_9213);
or U12470 (N_12470,N_7674,N_8981);
nand U12471 (N_12471,N_8819,N_7507);
nand U12472 (N_12472,N_8459,N_7509);
xor U12473 (N_12473,N_8180,N_9058);
and U12474 (N_12474,N_8068,N_8299);
xor U12475 (N_12475,N_9205,N_9597);
nand U12476 (N_12476,N_7565,N_8842);
nand U12477 (N_12477,N_8502,N_8693);
xor U12478 (N_12478,N_9094,N_8538);
or U12479 (N_12479,N_8099,N_8218);
and U12480 (N_12480,N_9803,N_7893);
xor U12481 (N_12481,N_7630,N_9968);
nor U12482 (N_12482,N_9518,N_9221);
nor U12483 (N_12483,N_9938,N_8018);
or U12484 (N_12484,N_7568,N_8353);
nor U12485 (N_12485,N_7782,N_7697);
or U12486 (N_12486,N_8526,N_9466);
nand U12487 (N_12487,N_8869,N_8112);
or U12488 (N_12488,N_8333,N_8872);
or U12489 (N_12489,N_9763,N_8737);
nand U12490 (N_12490,N_9071,N_9286);
and U12491 (N_12491,N_9062,N_8383);
and U12492 (N_12492,N_9793,N_8117);
nand U12493 (N_12493,N_8883,N_7845);
and U12494 (N_12494,N_9595,N_8042);
or U12495 (N_12495,N_9817,N_9647);
nand U12496 (N_12496,N_8634,N_8730);
nand U12497 (N_12497,N_8481,N_7751);
or U12498 (N_12498,N_8165,N_9872);
and U12499 (N_12499,N_8284,N_9200);
and U12500 (N_12500,N_11520,N_12351);
nand U12501 (N_12501,N_10880,N_10411);
and U12502 (N_12502,N_10009,N_11730);
or U12503 (N_12503,N_11772,N_11685);
or U12504 (N_12504,N_10339,N_12352);
and U12505 (N_12505,N_11139,N_10913);
nor U12506 (N_12506,N_10324,N_11953);
and U12507 (N_12507,N_11480,N_11185);
or U12508 (N_12508,N_10772,N_11711);
nor U12509 (N_12509,N_10056,N_10771);
and U12510 (N_12510,N_10791,N_10370);
nand U12511 (N_12511,N_11177,N_12224);
and U12512 (N_12512,N_12250,N_12493);
and U12513 (N_12513,N_12385,N_11717);
xor U12514 (N_12514,N_11737,N_10741);
nor U12515 (N_12515,N_12217,N_12077);
and U12516 (N_12516,N_10679,N_11962);
nor U12517 (N_12517,N_10724,N_11227);
nor U12518 (N_12518,N_12497,N_10361);
and U12519 (N_12519,N_12173,N_10357);
nor U12520 (N_12520,N_11947,N_12128);
or U12521 (N_12521,N_11254,N_11651);
xor U12522 (N_12522,N_10836,N_12009);
nor U12523 (N_12523,N_11178,N_11092);
nand U12524 (N_12524,N_10181,N_12482);
xor U12525 (N_12525,N_10206,N_10519);
or U12526 (N_12526,N_10802,N_11538);
xnor U12527 (N_12527,N_10360,N_11558);
xnor U12528 (N_12528,N_11066,N_11061);
xnor U12529 (N_12529,N_11755,N_11171);
xnor U12530 (N_12530,N_12285,N_10337);
xor U12531 (N_12531,N_10329,N_10254);
xor U12532 (N_12532,N_11463,N_11720);
xnor U12533 (N_12533,N_11549,N_11854);
or U12534 (N_12534,N_11359,N_10248);
or U12535 (N_12535,N_10010,N_11332);
or U12536 (N_12536,N_10905,N_11161);
and U12537 (N_12537,N_12345,N_11202);
nor U12538 (N_12538,N_11942,N_10582);
and U12539 (N_12539,N_10420,N_10968);
or U12540 (N_12540,N_10143,N_10467);
xor U12541 (N_12541,N_11676,N_11602);
nand U12542 (N_12542,N_11133,N_11277);
or U12543 (N_12543,N_10767,N_10302);
nand U12544 (N_12544,N_11808,N_10222);
nand U12545 (N_12545,N_12498,N_10655);
and U12546 (N_12546,N_10027,N_10053);
nand U12547 (N_12547,N_10850,N_10389);
xor U12548 (N_12548,N_10901,N_11909);
nor U12549 (N_12549,N_12304,N_10640);
or U12550 (N_12550,N_11247,N_11539);
and U12551 (N_12551,N_10769,N_10536);
nor U12552 (N_12552,N_10753,N_11762);
and U12553 (N_12553,N_12241,N_11391);
xor U12554 (N_12554,N_12338,N_12181);
and U12555 (N_12555,N_11355,N_11191);
nor U12556 (N_12556,N_12000,N_11877);
nor U12557 (N_12557,N_10658,N_11036);
and U12558 (N_12558,N_10689,N_12073);
and U12559 (N_12559,N_11484,N_11243);
nor U12560 (N_12560,N_10390,N_11504);
nand U12561 (N_12561,N_10030,N_10817);
nor U12562 (N_12562,N_11938,N_10933);
xnor U12563 (N_12563,N_12177,N_12264);
and U12564 (N_12564,N_10867,N_10780);
nand U12565 (N_12565,N_12136,N_10726);
nand U12566 (N_12566,N_10505,N_12303);
or U12567 (N_12567,N_12278,N_10977);
and U12568 (N_12568,N_10957,N_12336);
and U12569 (N_12569,N_11124,N_11940);
or U12570 (N_12570,N_10683,N_10935);
xor U12571 (N_12571,N_10888,N_10177);
or U12572 (N_12572,N_11271,N_12066);
nor U12573 (N_12573,N_10629,N_11159);
or U12574 (N_12574,N_10362,N_12216);
and U12575 (N_12575,N_11014,N_11879);
nor U12576 (N_12576,N_11205,N_11352);
nand U12577 (N_12577,N_12448,N_10576);
xor U12578 (N_12578,N_10623,N_11491);
and U12579 (N_12579,N_10703,N_11663);
nor U12580 (N_12580,N_10785,N_11279);
or U12581 (N_12581,N_11715,N_10507);
xnor U12582 (N_12582,N_10837,N_10891);
or U12583 (N_12583,N_10033,N_12170);
xor U12584 (N_12584,N_10534,N_11103);
and U12585 (N_12585,N_12317,N_10923);
nand U12586 (N_12586,N_10155,N_10454);
or U12587 (N_12587,N_11871,N_11620);
and U12588 (N_12588,N_11401,N_11180);
nand U12589 (N_12589,N_10607,N_11326);
nor U12590 (N_12590,N_10555,N_12373);
nand U12591 (N_12591,N_10131,N_10456);
nor U12592 (N_12592,N_11437,N_12394);
or U12593 (N_12593,N_10103,N_10075);
and U12594 (N_12594,N_11059,N_11422);
or U12595 (N_12595,N_11550,N_10947);
or U12596 (N_12596,N_11988,N_11402);
nand U12597 (N_12597,N_12244,N_12310);
or U12598 (N_12598,N_10224,N_11725);
nor U12599 (N_12599,N_11980,N_10427);
nand U12600 (N_12600,N_11246,N_10061);
or U12601 (N_12601,N_11276,N_10062);
xor U12602 (N_12602,N_10770,N_12123);
nor U12603 (N_12603,N_11691,N_10100);
and U12604 (N_12604,N_10425,N_11547);
xnor U12605 (N_12605,N_11971,N_10488);
nand U12606 (N_12606,N_12455,N_10765);
nand U12607 (N_12607,N_11374,N_11848);
xor U12608 (N_12608,N_10015,N_11849);
nor U12609 (N_12609,N_11423,N_10101);
and U12610 (N_12610,N_10147,N_12006);
xnor U12611 (N_12611,N_10333,N_10599);
or U12612 (N_12612,N_10966,N_10719);
nand U12613 (N_12613,N_10069,N_11232);
nor U12614 (N_12614,N_10717,N_11987);
nor U12615 (N_12615,N_10188,N_11412);
nand U12616 (N_12616,N_11206,N_11233);
nor U12617 (N_12617,N_11065,N_10478);
nand U12618 (N_12618,N_10554,N_10512);
nor U12619 (N_12619,N_10669,N_10274);
xnor U12620 (N_12620,N_10032,N_10443);
and U12621 (N_12621,N_10471,N_11572);
nand U12622 (N_12622,N_10906,N_11687);
and U12623 (N_12623,N_11740,N_10190);
nand U12624 (N_12624,N_10676,N_12486);
nand U12625 (N_12625,N_11381,N_11021);
nand U12626 (N_12626,N_11496,N_11797);
or U12627 (N_12627,N_10170,N_10296);
or U12628 (N_12628,N_11783,N_12419);
nor U12629 (N_12629,N_10474,N_12207);
or U12630 (N_12630,N_12214,N_10077);
and U12631 (N_12631,N_10725,N_11302);
nor U12632 (N_12632,N_11071,N_11111);
nor U12633 (N_12633,N_10870,N_12021);
and U12634 (N_12634,N_11472,N_10498);
xor U12635 (N_12635,N_11880,N_10135);
nand U12636 (N_12636,N_10315,N_10593);
nand U12637 (N_12637,N_12218,N_12042);
nor U12638 (N_12638,N_10985,N_11989);
or U12639 (N_12639,N_11904,N_10440);
nor U12640 (N_12640,N_10996,N_11869);
xnor U12641 (N_12641,N_12478,N_10145);
or U12642 (N_12642,N_11767,N_11050);
and U12643 (N_12643,N_10876,N_12197);
nor U12644 (N_12644,N_11827,N_12434);
or U12645 (N_12645,N_10070,N_12456);
nand U12646 (N_12646,N_11333,N_11300);
nor U12647 (N_12647,N_12089,N_10861);
and U12648 (N_12648,N_10183,N_11739);
and U12649 (N_12649,N_12382,N_12225);
and U12650 (N_12650,N_11918,N_10338);
nand U12651 (N_12651,N_11228,N_10732);
or U12652 (N_12652,N_10429,N_11366);
or U12653 (N_12653,N_11765,N_10908);
or U12654 (N_12654,N_10482,N_11757);
or U12655 (N_12655,N_11444,N_12034);
or U12656 (N_12656,N_10815,N_10270);
xnor U12657 (N_12657,N_11492,N_11107);
and U12658 (N_12658,N_12029,N_10355);
or U12659 (N_12659,N_11590,N_11314);
nand U12660 (N_12660,N_12143,N_10079);
xor U12661 (N_12661,N_11217,N_11046);
nand U12662 (N_12662,N_10028,N_10094);
nand U12663 (N_12663,N_12255,N_11514);
xnor U12664 (N_12664,N_10714,N_11670);
nor U12665 (N_12665,N_12316,N_11821);
nor U12666 (N_12666,N_10843,N_10723);
nor U12667 (N_12667,N_11612,N_11210);
nand U12668 (N_12668,N_11501,N_10890);
nand U12669 (N_12669,N_10763,N_11749);
xor U12670 (N_12670,N_10783,N_12182);
nand U12671 (N_12671,N_12124,N_12023);
nand U12672 (N_12672,N_11203,N_12201);
and U12673 (N_12673,N_11331,N_10937);
and U12674 (N_12674,N_11703,N_11097);
xnor U12675 (N_12675,N_11712,N_10489);
nand U12676 (N_12676,N_11468,N_10911);
and U12677 (N_12677,N_12044,N_10757);
and U12678 (N_12678,N_11011,N_11702);
xor U12679 (N_12679,N_12413,N_11681);
or U12680 (N_12680,N_11127,N_12298);
or U12681 (N_12681,N_10014,N_11536);
or U12682 (N_12682,N_12240,N_11546);
or U12683 (N_12683,N_10039,N_11897);
nor U12684 (N_12684,N_11796,N_12393);
nand U12685 (N_12685,N_11321,N_11335);
or U12686 (N_12686,N_10684,N_10118);
nand U12687 (N_12687,N_11045,N_10195);
nor U12688 (N_12688,N_10899,N_12375);
xor U12689 (N_12689,N_11769,N_12194);
or U12690 (N_12690,N_11995,N_10169);
nand U12691 (N_12691,N_12347,N_10350);
nand U12692 (N_12692,N_11922,N_12049);
or U12693 (N_12693,N_12301,N_11308);
nand U12694 (N_12694,N_11642,N_12152);
nor U12695 (N_12695,N_10262,N_10213);
nand U12696 (N_12696,N_11174,N_11950);
or U12697 (N_12697,N_10813,N_10748);
and U12698 (N_12698,N_11519,N_10305);
nand U12699 (N_12699,N_11616,N_11750);
or U12700 (N_12700,N_11035,N_11598);
and U12701 (N_12701,N_11009,N_12221);
or U12702 (N_12702,N_11242,N_12184);
or U12703 (N_12703,N_10711,N_12071);
and U12704 (N_12704,N_12453,N_10191);
or U12705 (N_12705,N_11378,N_11441);
nand U12706 (N_12706,N_11664,N_10267);
nor U12707 (N_12707,N_11701,N_10619);
or U12708 (N_12708,N_11179,N_11680);
nor U12709 (N_12709,N_11407,N_10250);
nand U12710 (N_12710,N_10886,N_12109);
xnor U12711 (N_12711,N_10106,N_12357);
nand U12712 (N_12712,N_11710,N_10497);
xor U12713 (N_12713,N_10826,N_10904);
nand U12714 (N_12714,N_12280,N_11760);
or U12715 (N_12715,N_10496,N_10462);
nand U12716 (N_12716,N_10940,N_11489);
and U12717 (N_12717,N_10006,N_10000);
or U12718 (N_12718,N_10561,N_11853);
and U12719 (N_12719,N_12212,N_10522);
xor U12720 (N_12720,N_10225,N_10406);
xnor U12721 (N_12721,N_10102,N_11636);
nor U12722 (N_12722,N_11917,N_11033);
or U12723 (N_12723,N_10217,N_11025);
nand U12724 (N_12724,N_11650,N_12459);
xnor U12725 (N_12725,N_10089,N_10893);
nand U12726 (N_12726,N_10961,N_11905);
and U12727 (N_12727,N_11292,N_10375);
nand U12728 (N_12728,N_12169,N_12239);
and U12729 (N_12729,N_11047,N_11813);
nand U12730 (N_12730,N_11340,N_10639);
nand U12731 (N_12731,N_11460,N_11955);
nand U12732 (N_12732,N_10245,N_11728);
nand U12733 (N_12733,N_11199,N_12268);
and U12734 (N_12734,N_10112,N_11928);
nand U12735 (N_12735,N_12174,N_11012);
or U12736 (N_12736,N_11447,N_10946);
xnor U12737 (N_12737,N_10625,N_10604);
nor U12738 (N_12738,N_10986,N_12472);
nor U12739 (N_12739,N_10351,N_11529);
nor U12740 (N_12740,N_12294,N_10749);
and U12741 (N_12741,N_11263,N_11259);
or U12742 (N_12742,N_12064,N_10883);
or U12743 (N_12743,N_11068,N_12245);
and U12744 (N_12744,N_10043,N_11056);
or U12745 (N_12745,N_11418,N_10007);
nand U12746 (N_12746,N_10394,N_10571);
nor U12747 (N_12747,N_10445,N_10068);
nor U12748 (N_12748,N_10203,N_11048);
nor U12749 (N_12749,N_11992,N_11709);
or U12750 (N_12750,N_10588,N_10052);
nor U12751 (N_12751,N_11163,N_10279);
xor U12752 (N_12752,N_11777,N_10927);
or U12753 (N_12753,N_10150,N_11957);
nor U12754 (N_12754,N_11822,N_11260);
and U12755 (N_12755,N_10346,N_12401);
and U12756 (N_12756,N_10779,N_10918);
nor U12757 (N_12757,N_11951,N_11522);
and U12758 (N_12758,N_11115,N_11360);
and U12759 (N_12759,N_11138,N_11884);
nand U12760 (N_12760,N_11991,N_11336);
xnor U12761 (N_12761,N_11090,N_10437);
and U12762 (N_12762,N_10857,N_11688);
nor U12763 (N_12763,N_10175,N_12376);
xnor U12764 (N_12764,N_10278,N_10326);
xnor U12765 (N_12765,N_10202,N_10016);
or U12766 (N_12766,N_12463,N_11224);
and U12767 (N_12767,N_11113,N_10408);
and U12768 (N_12768,N_10781,N_11920);
xor U12769 (N_12769,N_11110,N_11555);
or U12770 (N_12770,N_10840,N_10520);
xnor U12771 (N_12771,N_10049,N_12289);
nor U12772 (N_12772,N_11038,N_11086);
and U12773 (N_12773,N_12113,N_11387);
xnor U12774 (N_12774,N_11858,N_11840);
nand U12775 (N_12775,N_11996,N_11278);
xnor U12776 (N_12776,N_10999,N_11888);
xor U12777 (N_12777,N_11781,N_11515);
or U12778 (N_12778,N_12074,N_11791);
and U12779 (N_12779,N_11317,N_11846);
nand U12780 (N_12780,N_11774,N_10677);
or U12781 (N_12781,N_11235,N_10592);
nand U12782 (N_12782,N_11830,N_12112);
xor U12783 (N_12783,N_10548,N_11325);
xor U12784 (N_12784,N_11288,N_11633);
and U12785 (N_12785,N_12187,N_11924);
xor U12786 (N_12786,N_12386,N_10651);
and U12787 (N_12787,N_10113,N_11250);
nand U12788 (N_12788,N_10167,N_10613);
nor U12789 (N_12789,N_11010,N_10879);
nor U12790 (N_12790,N_10776,N_10307);
nand U12791 (N_12791,N_10388,N_10570);
xor U12792 (N_12792,N_10690,N_12390);
xnor U12793 (N_12793,N_11528,N_12360);
nand U12794 (N_12794,N_10382,N_11426);
or U12795 (N_12795,N_11104,N_12223);
xnor U12796 (N_12796,N_12062,N_10092);
xnor U12797 (N_12797,N_11882,N_12037);
nor U12798 (N_12798,N_10345,N_11764);
nand U12799 (N_12799,N_10896,N_11756);
xnor U12800 (N_12800,N_10553,N_10415);
nor U12801 (N_12801,N_10981,N_10795);
nor U12802 (N_12802,N_10805,N_10281);
and U12803 (N_12803,N_11132,N_11208);
nor U12804 (N_12804,N_11109,N_10759);
xor U12805 (N_12805,N_11446,N_10494);
and U12806 (N_12806,N_11576,N_11872);
or U12807 (N_12807,N_11493,N_11386);
nor U12808 (N_12808,N_11147,N_11022);
nor U12809 (N_12809,N_10695,N_12059);
and U12810 (N_12810,N_11075,N_11763);
nand U12811 (N_12811,N_11274,N_11617);
or U12812 (N_12812,N_10319,N_11399);
nor U12813 (N_12813,N_10585,N_10137);
xnor U12814 (N_12814,N_12231,N_12363);
xor U12815 (N_12815,N_12243,N_10929);
xor U12816 (N_12816,N_10897,N_11442);
or U12817 (N_12817,N_11170,N_12052);
and U12818 (N_12818,N_11815,N_10855);
nand U12819 (N_12819,N_10313,N_10814);
xnor U12820 (N_12820,N_10473,N_10451);
nor U12821 (N_12821,N_10434,N_11149);
nand U12822 (N_12822,N_10410,N_11084);
nor U12823 (N_12823,N_12148,N_10697);
xnor U12824 (N_12824,N_12334,N_11679);
xor U12825 (N_12825,N_11741,N_12101);
xor U12826 (N_12826,N_10589,N_10654);
or U12827 (N_12827,N_12114,N_11385);
xnor U12828 (N_12828,N_10269,N_10441);
or U12829 (N_12829,N_11272,N_10648);
nor U12830 (N_12830,N_11860,N_11482);
or U12831 (N_12831,N_10902,N_10164);
xor U12832 (N_12832,N_10852,N_10894);
or U12833 (N_12833,N_10866,N_12251);
nor U12834 (N_12834,N_12020,N_10675);
or U12835 (N_12835,N_11868,N_11560);
and U12836 (N_12836,N_12175,N_10212);
nor U12837 (N_12837,N_11912,N_12305);
or U12838 (N_12838,N_11622,N_10393);
or U12839 (N_12839,N_10887,N_11850);
or U12840 (N_12840,N_11742,N_11162);
or U12841 (N_12841,N_11098,N_11672);
nand U12842 (N_12842,N_11934,N_10127);
nand U12843 (N_12843,N_11220,N_10875);
nand U12844 (N_12844,N_11478,N_12265);
nand U12845 (N_12845,N_11586,N_10931);
or U12846 (N_12846,N_12164,N_11275);
nand U12847 (N_12847,N_10997,N_12208);
or U12848 (N_12848,N_10403,N_12185);
and U12849 (N_12849,N_10688,N_12499);
nor U12850 (N_12850,N_10258,N_11674);
and U12851 (N_12851,N_12428,N_10829);
nand U12852 (N_12852,N_11420,N_10341);
nand U12853 (N_12853,N_11972,N_10128);
nor U12854 (N_12854,N_10354,N_10737);
xor U12855 (N_12855,N_10559,N_10895);
and U12856 (N_12856,N_10988,N_11062);
and U12857 (N_12857,N_10332,N_10466);
or U12858 (N_12858,N_12365,N_11117);
xnor U12859 (N_12859,N_10823,N_10287);
xor U12860 (N_12860,N_12254,N_12322);
and U12861 (N_12861,N_12438,N_10708);
xor U12862 (N_12862,N_10597,N_10325);
nor U12863 (N_12863,N_12171,N_12327);
or U12864 (N_12864,N_12132,N_12421);
xnor U12865 (N_12865,N_11017,N_11878);
nand U12866 (N_12866,N_11212,N_10458);
nor U12867 (N_12867,N_12086,N_10513);
nor U12868 (N_12868,N_11531,N_10461);
nand U12869 (N_12869,N_11583,N_11265);
nand U12870 (N_12870,N_10130,N_10421);
or U12871 (N_12871,N_11559,N_10139);
nor U12872 (N_12872,N_11876,N_12468);
or U12873 (N_12873,N_11291,N_10707);
and U12874 (N_12874,N_11665,N_10398);
nand U12875 (N_12875,N_11207,N_11627);
or U12876 (N_12876,N_10808,N_12417);
or U12877 (N_12877,N_10058,N_10706);
xor U12878 (N_12878,N_10146,N_12331);
or U12879 (N_12879,N_10086,N_10331);
xnor U12880 (N_12880,N_12195,N_12209);
nand U12881 (N_12881,N_11875,N_10407);
nand U12882 (N_12882,N_11319,N_11338);
nor U12883 (N_12883,N_11584,N_11443);
xor U12884 (N_12884,N_11776,N_11006);
or U12885 (N_12885,N_10686,N_10673);
or U12886 (N_12886,N_12444,N_12247);
and U12887 (N_12887,N_10636,N_12105);
nor U12888 (N_12888,N_10249,N_11900);
nand U12889 (N_12889,N_11055,N_10965);
xor U12890 (N_12890,N_10359,N_10209);
or U12891 (N_12891,N_11524,N_11719);
or U12892 (N_12892,N_11511,N_10263);
nand U12893 (N_12893,N_11505,N_11044);
xnor U12894 (N_12894,N_11637,N_11383);
and U12895 (N_12895,N_10704,N_11350);
nor U12896 (N_12896,N_10608,N_12356);
and U12897 (N_12897,N_11095,N_11356);
and U12898 (N_12898,N_10500,N_10903);
nor U12899 (N_12899,N_11836,N_11731);
or U12900 (N_12900,N_10612,N_10044);
and U12901 (N_12901,N_11395,N_11790);
or U12902 (N_12902,N_10793,N_11394);
nor U12903 (N_12903,N_12033,N_10252);
or U12904 (N_12904,N_10975,N_11348);
or U12905 (N_12905,N_12041,N_10868);
nand U12906 (N_12906,N_11419,N_10530);
and U12907 (N_12907,N_11997,N_11994);
nor U12908 (N_12908,N_10702,N_11736);
and U12909 (N_12909,N_10801,N_10297);
or U12910 (N_12910,N_11248,N_12423);
and U12911 (N_12911,N_10934,N_12362);
nand U12912 (N_12912,N_11082,N_11824);
and U12913 (N_12913,N_10566,N_11693);
nand U12914 (N_12914,N_10944,N_11581);
and U12915 (N_12915,N_10125,N_11771);
or U12916 (N_12916,N_11015,N_10994);
nor U12917 (N_12917,N_10084,N_11379);
and U12918 (N_12918,N_11659,N_11600);
nand U12919 (N_12919,N_10615,N_12013);
or U12920 (N_12920,N_11431,N_11838);
xnor U12921 (N_12921,N_11434,N_12203);
or U12922 (N_12922,N_11502,N_10849);
nand U12923 (N_12923,N_11122,N_10760);
nor U12924 (N_12924,N_10951,N_10255);
xor U12925 (N_12925,N_11969,N_12081);
and U12926 (N_12926,N_12258,N_11847);
nor U12927 (N_12927,N_11436,N_10956);
xor U12928 (N_12928,N_10091,N_10960);
nand U12929 (N_12929,N_10465,N_11594);
and U12930 (N_12930,N_12312,N_11655);
xor U12931 (N_12931,N_10081,N_10120);
and U12932 (N_12932,N_11453,N_10384);
xor U12933 (N_12933,N_10787,N_12172);
or U12934 (N_12934,N_10614,N_11251);
or U12935 (N_12935,N_10020,N_12107);
nor U12936 (N_12936,N_10515,N_10609);
or U12937 (N_12937,N_11329,N_12252);
nor U12938 (N_12938,N_10539,N_10898);
xnor U12939 (N_12939,N_11892,N_10179);
or U12940 (N_12940,N_12155,N_11887);
and U12941 (N_12941,N_11935,N_10162);
and U12942 (N_12942,N_11456,N_12068);
nand U12943 (N_12943,N_10369,N_10036);
xnor U12944 (N_12944,N_11753,N_10066);
xor U12945 (N_12945,N_10533,N_11222);
xnor U12946 (N_12946,N_10037,N_11438);
or U12947 (N_12947,N_11105,N_12139);
or U12948 (N_12948,N_11722,N_10716);
or U12949 (N_12949,N_12485,N_11956);
or U12950 (N_12950,N_11816,N_11005);
and U12951 (N_12951,N_10914,N_11101);
and U12952 (N_12952,N_11462,N_11985);
or U12953 (N_12953,N_12093,N_11981);
and U12954 (N_12954,N_11999,N_11964);
or U12955 (N_12955,N_10303,N_11389);
or U12956 (N_12956,N_10563,N_11164);
or U12957 (N_12957,N_11414,N_10864);
nor U12958 (N_12958,N_10631,N_11613);
or U12959 (N_12959,N_11428,N_11196);
nor U12960 (N_12960,N_12420,N_11049);
nor U12961 (N_12961,N_11069,N_11927);
xnor U12962 (N_12962,N_10735,N_11020);
nand U12963 (N_12963,N_10080,N_10976);
nor U12964 (N_12964,N_11324,N_11610);
xnor U12965 (N_12965,N_10739,N_12308);
xnor U12966 (N_12966,N_12379,N_11952);
xnor U12967 (N_12967,N_11193,N_10881);
xnor U12968 (N_12968,N_10945,N_10057);
and U12969 (N_12969,N_11024,N_12002);
nor U12970 (N_12970,N_11269,N_12057);
nand U12971 (N_12971,N_10733,N_10211);
nand U12972 (N_12972,N_11628,N_10157);
xnor U12973 (N_12973,N_12321,N_10626);
xor U12974 (N_12974,N_10132,N_11939);
nor U12975 (N_12975,N_11509,N_11320);
xnor U12976 (N_12976,N_11435,N_11239);
or U12977 (N_12977,N_11735,N_10405);
or U12978 (N_12978,N_12481,N_10122);
xnor U12979 (N_12979,N_12069,N_10827);
nand U12980 (N_12980,N_10344,N_10353);
xnor U12981 (N_12981,N_10644,N_11353);
and U12982 (N_12982,N_11266,N_10096);
and U12983 (N_12983,N_10356,N_11141);
nor U12984 (N_12984,N_11345,N_11945);
xor U12985 (N_12985,N_11782,N_12306);
xor U12986 (N_12986,N_10266,N_10982);
nor U12987 (N_12987,N_11675,N_11304);
nand U12988 (N_12988,N_10051,N_10792);
nand U12989 (N_12989,N_10308,N_10798);
nand U12990 (N_12990,N_11770,N_11330);
xor U12991 (N_12991,N_11237,N_11649);
or U12992 (N_12992,N_10283,N_10199);
or U12993 (N_12993,N_10348,N_10192);
or U12994 (N_12994,N_11318,N_11218);
nand U12995 (N_12995,N_11123,N_11365);
and U12996 (N_12996,N_11388,N_11019);
nand U12997 (N_12997,N_11802,N_11784);
and U12998 (N_12998,N_11571,N_10844);
or U12999 (N_12999,N_10277,N_10368);
nand U13000 (N_13000,N_10055,N_12426);
nor U13001 (N_13001,N_11487,N_12070);
and U13002 (N_13002,N_11295,N_11864);
or U13003 (N_13003,N_12380,N_11798);
or U13004 (N_13004,N_12409,N_11601);
nor U13005 (N_13005,N_10453,N_12028);
xor U13006 (N_13006,N_10071,N_12416);
nor U13007 (N_13007,N_11188,N_11192);
xnor U13008 (N_13008,N_12084,N_10314);
xor U13009 (N_13009,N_10076,N_11214);
xor U13010 (N_13010,N_10484,N_11297);
nand U13011 (N_13011,N_11226,N_10973);
or U13012 (N_13012,N_11832,N_10450);
and U13013 (N_13013,N_10859,N_11656);
and U13014 (N_13014,N_12364,N_12083);
nor U13015 (N_13015,N_11469,N_12159);
xor U13016 (N_13016,N_11057,N_11803);
nor U13017 (N_13017,N_10204,N_10025);
or U13018 (N_13018,N_10509,N_12001);
and U13019 (N_13019,N_11591,N_10618);
xnor U13020 (N_13020,N_10021,N_10751);
xor U13021 (N_13021,N_10387,N_11729);
nor U13022 (N_13022,N_12490,N_11384);
or U13023 (N_13023,N_10380,N_11789);
xnor U13024 (N_13024,N_10715,N_12094);
nor U13025 (N_13025,N_10309,N_11721);
nor U13026 (N_13026,N_11053,N_10138);
nand U13027 (N_13027,N_11458,N_10635);
and U13028 (N_13028,N_10114,N_11157);
or U13029 (N_13029,N_11527,N_12460);
and U13030 (N_13030,N_12349,N_10178);
and U13031 (N_13031,N_11289,N_12025);
or U13032 (N_13032,N_11373,N_12205);
nand U13033 (N_13033,N_11758,N_10232);
nor U13034 (N_13034,N_10449,N_12215);
xor U13035 (N_13035,N_11400,N_11673);
xor U13036 (N_13036,N_12313,N_10117);
nor U13037 (N_13037,N_11608,N_11173);
nor U13038 (N_13038,N_12344,N_11216);
xor U13039 (N_13039,N_10201,N_12477);
and U13040 (N_13040,N_10334,N_10105);
and U13041 (N_13041,N_10523,N_11483);
or U13042 (N_13042,N_10573,N_12135);
nand U13043 (N_13043,N_10758,N_11376);
xor U13044 (N_13044,N_11016,N_11751);
nand U13045 (N_13045,N_11966,N_11042);
or U13046 (N_13046,N_11844,N_11778);
and U13047 (N_13047,N_11933,N_12496);
xor U13048 (N_13048,N_10300,N_11404);
xor U13049 (N_13049,N_10532,N_10754);
or U13050 (N_13050,N_12178,N_10430);
nor U13051 (N_13051,N_11894,N_11833);
nand U13052 (N_13052,N_10470,N_11857);
nand U13053 (N_13053,N_11327,N_12063);
nor U13054 (N_13054,N_10642,N_11167);
and U13055 (N_13055,N_11371,N_11919);
and U13056 (N_13056,N_11085,N_10622);
or U13057 (N_13057,N_11100,N_11074);
nand U13058 (N_13058,N_10271,N_11614);
and U13059 (N_13059,N_12075,N_10562);
and U13060 (N_13060,N_10745,N_10712);
xnor U13061 (N_13061,N_10241,N_10264);
or U13062 (N_13062,N_12092,N_10853);
nor U13063 (N_13063,N_10371,N_11172);
nand U13064 (N_13064,N_11677,N_10820);
or U13065 (N_13065,N_10115,N_11883);
xnor U13066 (N_13066,N_11958,N_11114);
nand U13067 (N_13067,N_10005,N_11564);
nand U13068 (N_13068,N_10939,N_10819);
and U13069 (N_13069,N_10803,N_11644);
xnor U13070 (N_13070,N_10119,N_10882);
or U13071 (N_13071,N_10672,N_11346);
nor U13072 (N_13072,N_11099,N_12297);
nand U13073 (N_13073,N_11593,N_12154);
and U13074 (N_13074,N_11580,N_11975);
or U13075 (N_13075,N_10537,N_10108);
xnor U13076 (N_13076,N_12326,N_10775);
nand U13077 (N_13077,N_10546,N_12279);
nor U13078 (N_13078,N_10696,N_12192);
and U13079 (N_13079,N_12036,N_12213);
or U13080 (N_13080,N_11241,N_11030);
xnor U13081 (N_13081,N_10008,N_10156);
or U13082 (N_13082,N_12353,N_10477);
nand U13083 (N_13083,N_12149,N_11323);
or U13084 (N_13084,N_12035,N_10662);
nor U13085 (N_13085,N_12102,N_10652);
nand U13086 (N_13086,N_10510,N_11152);
or U13087 (N_13087,N_10987,N_12127);
xnor U13088 (N_13088,N_12072,N_11370);
xnor U13089 (N_13089,N_10166,N_11595);
xor U13090 (N_13090,N_12090,N_10954);
and U13091 (N_13091,N_12492,N_10871);
nor U13092 (N_13092,N_12466,N_11358);
xor U13093 (N_13093,N_10479,N_10653);
or U13094 (N_13094,N_10231,N_10928);
or U13095 (N_13095,N_11984,N_11624);
and U13096 (N_13096,N_10123,N_10383);
nor U13097 (N_13097,N_10667,N_12377);
xnor U13098 (N_13098,N_11965,N_10740);
and U13099 (N_13099,N_10874,N_10832);
nor U13100 (N_13100,N_10692,N_11603);
nand U13101 (N_13101,N_10402,N_10833);
and U13102 (N_13102,N_10374,N_10804);
nand U13103 (N_13103,N_10784,N_11852);
or U13104 (N_13104,N_12300,N_11240);
or U13105 (N_13105,N_10744,N_10565);
xor U13106 (N_13106,N_11819,N_10932);
or U13107 (N_13107,N_12473,N_10289);
nor U13108 (N_13108,N_11229,N_12436);
nor U13109 (N_13109,N_12381,N_11804);
and U13110 (N_13110,N_11565,N_10634);
or U13111 (N_13111,N_12058,N_10807);
and U13112 (N_13112,N_10503,N_11837);
nand U13113 (N_13113,N_12323,N_11856);
xor U13114 (N_13114,N_12435,N_12372);
and U13115 (N_13115,N_11578,N_11165);
xnor U13116 (N_13116,N_12383,N_11316);
xor U13117 (N_13117,N_12050,N_10646);
or U13118 (N_13118,N_11060,N_10316);
nand U13119 (N_13119,N_12189,N_10290);
and U13120 (N_13120,N_12480,N_12055);
and U13121 (N_13121,N_10885,N_10835);
nand U13122 (N_13122,N_10574,N_11129);
nor U13123 (N_13123,N_11817,N_10799);
and U13124 (N_13124,N_10547,N_12311);
nor U13125 (N_13125,N_11267,N_11579);
xor U13126 (N_13126,N_11160,N_11530);
and U13127 (N_13127,N_10149,N_10605);
nor U13128 (N_13128,N_12030,N_12230);
xor U13129 (N_13129,N_12080,N_10306);
xor U13130 (N_13130,N_10261,N_10378);
nor U13131 (N_13131,N_10794,N_10073);
nor U13132 (N_13132,N_11700,N_11621);
nand U13133 (N_13133,N_11311,N_11041);
nand U13134 (N_13134,N_10409,N_10611);
nand U13135 (N_13135,N_12119,N_10432);
nor U13136 (N_13136,N_11296,N_11126);
xnor U13137 (N_13137,N_10417,N_12088);
xnor U13138 (N_13138,N_10218,N_11648);
and U13139 (N_13139,N_11724,N_10168);
nor U13140 (N_13140,N_11119,N_10969);
nor U13141 (N_13141,N_10072,N_11851);
nand U13142 (N_13142,N_11548,N_10436);
and U13143 (N_13143,N_11990,N_10038);
or U13144 (N_13144,N_11696,N_11153);
xnor U13145 (N_13145,N_10060,N_10990);
and U13146 (N_13146,N_12065,N_12199);
or U13147 (N_13147,N_11541,N_11766);
and U13148 (N_13148,N_10971,N_12236);
or U13149 (N_13149,N_10910,N_11903);
and U13150 (N_13150,N_12186,N_10433);
xnor U13151 (N_13151,N_11396,N_12431);
xnor U13152 (N_13152,N_12176,N_10811);
nand U13153 (N_13153,N_11977,N_10363);
and U13154 (N_13154,N_12325,N_11282);
nor U13155 (N_13155,N_10974,N_12467);
nand U13156 (N_13156,N_10491,N_10366);
nand U13157 (N_13157,N_10093,N_11245);
or U13158 (N_13158,N_11341,N_10627);
xor U13159 (N_13159,N_11439,N_12017);
nand U13160 (N_13160,N_10180,N_11054);
nand U13161 (N_13161,N_10260,N_11343);
or U13162 (N_13162,N_10685,N_10148);
or U13163 (N_13163,N_11716,N_11512);
nor U13164 (N_13164,N_10590,N_11754);
nor U13165 (N_13165,N_11003,N_11108);
xor U13166 (N_13166,N_10797,N_12146);
xnor U13167 (N_13167,N_12424,N_10736);
or U13168 (N_13168,N_10431,N_10884);
nand U13169 (N_13169,N_10647,N_10670);
nor U13170 (N_13170,N_11175,N_12442);
xor U13171 (N_13171,N_10050,N_10328);
and U13172 (N_13172,N_11051,N_10054);
nor U13173 (N_13173,N_11574,N_10244);
nor U13174 (N_13174,N_11499,N_10728);
nor U13175 (N_13175,N_12163,N_11186);
xor U13176 (N_13176,N_12281,N_11517);
nor U13177 (N_13177,N_10518,N_12452);
or U13178 (N_13178,N_11886,N_10970);
nand U13179 (N_13179,N_12087,N_11623);
xnor U13180 (N_13180,N_10630,N_11398);
nor U13181 (N_13181,N_10734,N_11982);
or U13182 (N_13182,N_10294,N_11592);
nor U13183 (N_13183,N_10578,N_11845);
xnor U13184 (N_13184,N_12219,N_12359);
and U13185 (N_13185,N_11902,N_11625);
or U13186 (N_13186,N_11142,N_12166);
xnor U13187 (N_13187,N_10134,N_12246);
nand U13188 (N_13188,N_10938,N_10789);
and U13189 (N_13189,N_11262,N_12193);
or U13190 (N_13190,N_11198,N_10525);
nor U13191 (N_13191,N_10097,N_10778);
nor U13192 (N_13192,N_12402,N_10011);
xnor U13193 (N_13193,N_10786,N_11923);
nor U13194 (N_13194,N_10452,N_10034);
and U13195 (N_13195,N_10577,N_11201);
or U13196 (N_13196,N_10774,N_12440);
nand U13197 (N_13197,N_10317,N_10216);
and U13198 (N_13198,N_11500,N_12309);
nor U13199 (N_13199,N_11561,N_11761);
and U13200 (N_13200,N_12091,N_10506);
and U13201 (N_13201,N_11079,N_10579);
xnor U13202 (N_13202,N_10463,N_11307);
xnor U13203 (N_13203,N_11023,N_10839);
nor U13204 (N_13204,N_10773,N_10730);
nor U13205 (N_13205,N_10142,N_10718);
xnor U13206 (N_13206,N_10173,N_11773);
nand U13207 (N_13207,N_11925,N_11136);
and U13208 (N_13208,N_10412,N_12054);
xnor U13209 (N_13209,N_10621,N_10273);
and U13210 (N_13210,N_11885,N_11273);
xnor U13211 (N_13211,N_10680,N_10495);
or U13212 (N_13212,N_12040,N_10660);
nor U13213 (N_13213,N_10024,N_10788);
or U13214 (N_13214,N_11793,N_11861);
nor U13215 (N_13215,N_11645,N_11197);
nor U13216 (N_13216,N_12097,N_10983);
nor U13217 (N_13217,N_11448,N_10182);
xnor U13218 (N_13218,N_11089,N_10018);
nand U13219 (N_13219,N_12446,N_11088);
xnor U13220 (N_13220,N_10502,N_12126);
nand U13221 (N_13221,N_12461,N_10721);
and U13222 (N_13222,N_10645,N_10659);
and U13223 (N_13223,N_11380,N_11344);
and U13224 (N_13224,N_10208,N_12008);
nand U13225 (N_13225,N_10842,N_11695);
nor U13226 (N_13226,N_12232,N_10099);
nand U13227 (N_13227,N_12259,N_11258);
or U13228 (N_13228,N_11169,N_11823);
nor U13229 (N_13229,N_11299,N_10460);
nand U13230 (N_13230,N_10246,N_11072);
xor U13231 (N_13231,N_11270,N_11211);
nand U13232 (N_13232,N_11029,N_10504);
or U13233 (N_13233,N_10386,N_10090);
nand U13234 (N_13234,N_11639,N_10153);
nand U13235 (N_13235,N_10838,N_10019);
xor U13236 (N_13236,N_10226,N_11759);
or U13237 (N_13237,N_10700,N_12198);
or U13238 (N_13238,N_10816,N_12016);
and U13239 (N_13239,N_10280,N_11707);
nor U13240 (N_13240,N_11087,N_11094);
or U13241 (N_13241,N_12151,N_10858);
nor U13242 (N_13242,N_10863,N_12378);
or U13243 (N_13243,N_12295,N_11305);
and U13244 (N_13244,N_11284,N_11873);
and U13245 (N_13245,N_11286,N_11252);
nor U13246 (N_13246,N_11310,N_11037);
xnor U13247 (N_13247,N_10755,N_11234);
xor U13248 (N_13248,N_11775,N_11473);
xnor U13249 (N_13249,N_12369,N_10581);
or U13250 (N_13250,N_12014,N_11657);
and U13251 (N_13251,N_10575,N_11334);
nand U13252 (N_13252,N_11026,N_12122);
and U13253 (N_13253,N_12333,N_12387);
or U13254 (N_13254,N_11190,N_10845);
xor U13255 (N_13255,N_11494,N_10637);
or U13256 (N_13256,N_10243,N_12427);
or U13257 (N_13257,N_11826,N_10233);
xnor U13258 (N_13258,N_11632,N_11134);
nand U13259 (N_13259,N_11256,N_11863);
nor U13260 (N_13260,N_10439,N_10230);
nand U13261 (N_13261,N_11184,N_11589);
nand U13262 (N_13262,N_10320,N_10268);
or U13263 (N_13263,N_11290,N_10722);
and U13264 (N_13264,N_10796,N_11450);
nand U13265 (N_13265,N_10508,N_12341);
and U13266 (N_13266,N_11889,N_10606);
xor U13267 (N_13267,N_12445,N_11121);
and U13268 (N_13268,N_10327,N_11131);
or U13269 (N_13269,N_12188,N_11526);
and U13270 (N_13270,N_12263,N_12328);
or U13271 (N_13271,N_11906,N_11605);
nor U13272 (N_13272,N_11429,N_10012);
nand U13273 (N_13273,N_11930,N_11293);
nand U13274 (N_13274,N_11787,N_10064);
nor U13275 (N_13275,N_12320,N_10521);
nand U13276 (N_13276,N_11459,N_11706);
and U13277 (N_13277,N_11552,N_11425);
nand U13278 (N_13278,N_10395,N_11692);
and U13279 (N_13279,N_10160,N_10917);
and U13280 (N_13280,N_11630,N_12211);
xnor U13281 (N_13281,N_10159,N_11921);
or U13282 (N_13282,N_11911,N_12429);
and U13283 (N_13283,N_10661,N_11916);
nor U13284 (N_13284,N_11570,N_11485);
nor U13285 (N_13285,N_12011,N_12430);
nand U13286 (N_13286,N_11806,N_10185);
nand U13287 (N_13287,N_12227,N_11168);
nor U13288 (N_13288,N_10993,N_12479);
nor U13289 (N_13289,N_12010,N_11467);
nand U13290 (N_13290,N_12183,N_10941);
nor U13291 (N_13291,N_12141,N_10595);
or U13292 (N_13292,N_10198,N_11954);
or U13293 (N_13293,N_12238,N_11535);
nor U13294 (N_13294,N_12339,N_11411);
nand U13295 (N_13295,N_11970,N_10942);
or U13296 (N_13296,N_10569,N_10638);
and U13297 (N_13297,N_12293,N_10687);
xnor U13298 (N_13298,N_11794,N_10551);
and U13299 (N_13299,N_10550,N_12019);
xnor U13300 (N_13300,N_10953,N_11080);
xnor U13301 (N_13301,N_11654,N_12096);
nor U13302 (N_13302,N_11585,N_10220);
xnor U13303 (N_13303,N_10682,N_11145);
or U13304 (N_13304,N_11640,N_10860);
and U13305 (N_13305,N_11834,N_10979);
nor U13306 (N_13306,N_10746,N_10256);
nand U13307 (N_13307,N_12076,N_11405);
xnor U13308 (N_13308,N_11150,N_10442);
and U13309 (N_13309,N_11200,N_12161);
xor U13310 (N_13310,N_12039,N_10215);
or U13311 (N_13311,N_10729,N_12007);
and U13312 (N_13312,N_10152,N_11810);
and U13313 (N_13313,N_11281,N_11181);
nand U13314 (N_13314,N_10397,N_12418);
nand U13315 (N_13315,N_10632,N_10336);
xnor U13316 (N_13316,N_12190,N_10641);
or U13317 (N_13317,N_10616,N_10624);
xnor U13318 (N_13318,N_12274,N_12454);
nor U13319 (N_13319,N_11039,N_12425);
or U13320 (N_13320,N_11008,N_11077);
nor U13321 (N_13321,N_10967,N_11818);
nand U13322 (N_13322,N_11238,N_12450);
xor U13323 (N_13323,N_11587,N_11667);
or U13324 (N_13324,N_11936,N_10543);
nor U13325 (N_13325,N_10110,N_10889);
nor U13326 (N_13326,N_12324,N_10856);
or U13327 (N_13327,N_11983,N_11596);
nor U13328 (N_13328,N_12012,N_11466);
or U13329 (N_13329,N_10731,N_10426);
nand U13330 (N_13330,N_11698,N_11481);
and U13331 (N_13331,N_11867,N_10285);
nor U13332 (N_13332,N_12342,N_11507);
nand U13333 (N_13333,N_10584,N_10189);
nand U13334 (N_13334,N_12433,N_10681);
xor U13335 (N_13335,N_10276,N_12015);
nand U13336 (N_13336,N_11669,N_11554);
xor U13337 (N_13337,N_10541,N_11941);
or U13338 (N_13338,N_11814,N_12206);
nor U13339 (N_13339,N_11926,N_11372);
xor U13340 (N_13340,N_11949,N_11083);
and U13341 (N_13341,N_10121,N_12368);
nand U13342 (N_13342,N_10742,N_11727);
or U13343 (N_13343,N_10259,N_10750);
nand U13344 (N_13344,N_10924,N_11874);
nor U13345 (N_13345,N_11475,N_10766);
nand U13346 (N_13346,N_11828,N_11257);
or U13347 (N_13347,N_10984,N_11413);
and U13348 (N_13348,N_11315,N_12156);
nor U13349 (N_13349,N_11031,N_12226);
and U13350 (N_13350,N_11686,N_10825);
xnor U13351 (N_13351,N_10691,N_12296);
or U13352 (N_13352,N_10877,N_12022);
xor U13353 (N_13353,N_11959,N_10221);
xor U13354 (N_13354,N_10492,N_11968);
nand U13355 (N_13355,N_10995,N_11364);
and U13356 (N_13356,N_10416,N_12350);
nor U13357 (N_13357,N_12374,N_12400);
or U13358 (N_13358,N_11452,N_11375);
and U13359 (N_13359,N_12314,N_12489);
nand U13360 (N_13360,N_11351,N_11120);
xnor U13361 (N_13361,N_11018,N_11743);
nand U13362 (N_13362,N_10372,N_10764);
and U13363 (N_13363,N_11301,N_11568);
nor U13364 (N_13364,N_11313,N_11430);
nor U13365 (N_13365,N_10223,N_10187);
nor U13366 (N_13366,N_11835,N_12266);
xor U13367 (N_13367,N_12291,N_10602);
and U13368 (N_13368,N_12051,N_10438);
xor U13369 (N_13369,N_11545,N_10295);
xor U13370 (N_13370,N_12389,N_11910);
nor U13371 (N_13371,N_10572,N_12043);
nor U13372 (N_13372,N_10311,N_11143);
and U13373 (N_13373,N_12125,N_10557);
or U13374 (N_13374,N_11619,N_11932);
nor U13375 (N_13375,N_10365,N_10257);
nor U13376 (N_13376,N_12284,N_10936);
nand U13377 (N_13377,N_12235,N_12204);
nor U13378 (N_13378,N_11244,N_12140);
or U13379 (N_13379,N_11597,N_12407);
nand U13380 (N_13380,N_12053,N_11312);
xnor U13381 (N_13381,N_11733,N_10617);
nor U13382 (N_13382,N_12157,N_11309);
xnor U13383 (N_13383,N_10435,N_12120);
nand U13384 (N_13384,N_12103,N_11540);
nor U13385 (N_13385,N_11785,N_11194);
nor U13386 (N_13386,N_10531,N_11455);
or U13387 (N_13387,N_10926,N_11799);
nor U13388 (N_13388,N_11154,N_11678);
xor U13389 (N_13389,N_11615,N_11779);
xnor U13390 (N_13390,N_11839,N_10738);
nand U13391 (N_13391,N_11490,N_10048);
nand U13392 (N_13392,N_12270,N_11829);
xor U13393 (N_13393,N_10210,N_12410);
xor U13394 (N_13394,N_12354,N_12361);
nor U13395 (N_13395,N_11342,N_10529);
or U13396 (N_13396,N_12412,N_11476);
and U13397 (N_13397,N_12346,N_10693);
xor U13398 (N_13398,N_11899,N_10872);
nand U13399 (N_13399,N_11895,N_11408);
or U13400 (N_13400,N_10992,N_10247);
and U13401 (N_13401,N_12038,N_10964);
nor U13402 (N_13402,N_12242,N_12138);
or U13403 (N_13403,N_11537,N_11638);
and U13404 (N_13404,N_12249,N_11704);
and U13405 (N_13405,N_12443,N_10564);
nand U13406 (N_13406,N_10475,N_11495);
nor U13407 (N_13407,N_11007,N_11189);
nand U13408 (N_13408,N_11513,N_11268);
and U13409 (N_13409,N_12487,N_10921);
or U13410 (N_13410,N_10067,N_10163);
or U13411 (N_13411,N_12116,N_10472);
xor U13412 (N_13412,N_12398,N_10948);
nor U13413 (N_13413,N_11236,N_10228);
xnor U13414 (N_13414,N_10330,N_11708);
xnor U13415 (N_13415,N_12302,N_10487);
and U13416 (N_13416,N_10958,N_12100);
or U13417 (N_13417,N_11034,N_10251);
xnor U13418 (N_13418,N_10912,N_11397);
nor U13419 (N_13419,N_10869,N_11215);
nor U13420 (N_13420,N_11699,N_11713);
or U13421 (N_13421,N_11410,N_10490);
nand U13422 (N_13422,N_10457,N_12129);
xor U13423 (N_13423,N_10705,N_12168);
nor U13424 (N_13424,N_10065,N_10665);
xor U13425 (N_13425,N_10962,N_11457);
nor U13426 (N_13426,N_12332,N_12343);
or U13427 (N_13427,N_12098,N_10818);
or U13428 (N_13428,N_10768,N_12290);
nand U13429 (N_13429,N_10126,N_10193);
and U13430 (N_13430,N_11841,N_10323);
and U13431 (N_13431,N_11349,N_10486);
or U13432 (N_13432,N_10567,N_11582);
nor U13433 (N_13433,N_10831,N_12018);
nand U13434 (N_13434,N_12260,N_12256);
xnor U13435 (N_13435,N_10526,N_12078);
nand U13436 (N_13436,N_11786,N_10253);
xnor U13437 (N_13437,N_10583,N_10628);
nor U13438 (N_13438,N_12047,N_11454);
nor U13439 (N_13439,N_12005,N_12391);
xor U13440 (N_13440,N_11811,N_10580);
nand U13441 (N_13441,N_10668,N_11403);
xnor U13442 (N_13442,N_12488,N_11805);
or U13443 (N_13443,N_10419,N_11306);
and U13444 (N_13444,N_11421,N_11788);
nand U13445 (N_13445,N_11427,N_10650);
nor U13446 (N_13446,N_12282,N_10424);
nand U13447 (N_13447,N_11209,N_11744);
xnor U13448 (N_13448,N_11652,N_11231);
nand U13449 (N_13449,N_10828,N_10423);
and U13450 (N_13450,N_10978,N_10980);
nand U13451 (N_13451,N_10291,N_10501);
and U13452 (N_13452,N_10900,N_12276);
nand U13453 (N_13453,N_11562,N_11634);
xnor U13454 (N_13454,N_10286,N_10560);
or U13455 (N_13455,N_11183,N_12269);
xor U13456 (N_13456,N_12469,N_10483);
nor U13457 (N_13457,N_11508,N_10082);
or U13458 (N_13458,N_10596,N_10916);
nand U13459 (N_13459,N_11204,N_10046);
xnor U13460 (N_13460,N_12257,N_10591);
nor U13461 (N_13461,N_10528,N_10558);
nor U13462 (N_13462,N_12133,N_11433);
and U13463 (N_13463,N_12275,N_10777);
xor U13464 (N_13464,N_10045,N_10556);
xor U13465 (N_13465,N_11093,N_12355);
nor U13466 (N_13466,N_10540,N_12283);
nor U13467 (N_13467,N_10373,N_10448);
xnor U13468 (N_13468,N_11451,N_10663);
xor U13469 (N_13469,N_11362,N_10310);
or U13470 (N_13470,N_10414,N_12476);
and U13471 (N_13471,N_11865,N_11151);
and U13472 (N_13472,N_10878,N_10743);
xor U13473 (N_13473,N_12406,N_10227);
or U13474 (N_13474,N_10598,N_12117);
nand U13475 (N_13475,N_10184,N_12210);
and U13476 (N_13476,N_10455,N_11606);
nor U13477 (N_13477,N_11557,N_12106);
nor U13478 (N_13478,N_11058,N_11569);
and U13479 (N_13479,N_10922,N_10643);
xnor U13480 (N_13480,N_12384,N_11261);
nor U13481 (N_13481,N_11747,N_11668);
or U13482 (N_13482,N_11577,N_10404);
xor U13483 (N_13483,N_11800,N_12370);
nor U13484 (N_13484,N_12441,N_10377);
or U13485 (N_13485,N_10088,N_12121);
nand U13486 (N_13486,N_10041,N_10376);
or U13487 (N_13487,N_12196,N_10322);
nand U13488 (N_13488,N_12272,N_10229);
or U13489 (N_13489,N_11553,N_10950);
xor U13490 (N_13490,N_11498,N_11322);
xnor U13491 (N_13491,N_10299,N_10418);
and U13492 (N_13492,N_10292,N_11219);
xnor U13493 (N_13493,N_11461,N_11812);
and U13494 (N_13494,N_11609,N_11525);
nor U13495 (N_13495,N_11734,N_11156);
and U13496 (N_13496,N_11807,N_11367);
xnor U13497 (N_13497,N_12191,N_10161);
nor U13498 (N_13498,N_11146,N_11859);
nand U13499 (N_13499,N_11298,N_11963);
and U13500 (N_13500,N_11660,N_12267);
or U13501 (N_13501,N_10610,N_10275);
and U13502 (N_13502,N_11102,N_11944);
nor U13503 (N_13503,N_12495,N_10136);
nor U13504 (N_13504,N_12367,N_12167);
nand U13505 (N_13505,N_10129,N_12414);
xor U13506 (N_13506,N_12180,N_10026);
xor U13507 (N_13507,N_10095,N_11449);
nor U13508 (N_13508,N_12358,N_11611);
nor U13509 (N_13509,N_10017,N_10234);
xnor U13510 (N_13510,N_12079,N_11510);
or U13511 (N_13511,N_12060,N_11563);
xnor U13512 (N_13512,N_11866,N_10727);
or U13513 (N_13513,N_10549,N_11723);
xnor U13514 (N_13514,N_11690,N_12229);
and U13515 (N_13515,N_10480,N_10542);
nor U13516 (N_13516,N_11973,N_11532);
nor U13517 (N_13517,N_11907,N_10282);
nand U13518 (N_13518,N_10538,N_10001);
or U13519 (N_13519,N_10476,N_11140);
xor U13520 (N_13520,N_12474,N_11416);
and U13521 (N_13521,N_10809,N_11144);
or U13522 (N_13522,N_10237,N_10925);
xnor U13523 (N_13523,N_11825,N_11067);
nor U13524 (N_13524,N_10151,N_11106);
nand U13525 (N_13525,N_12248,N_11195);
or U13526 (N_13526,N_12288,N_12024);
nor U13527 (N_13527,N_10527,N_12439);
xnor U13528 (N_13528,N_11937,N_11542);
nand U13529 (N_13529,N_11694,N_11842);
nor U13530 (N_13530,N_10002,N_11726);
nand U13531 (N_13531,N_10240,N_11626);
xnor U13532 (N_13532,N_12415,N_11409);
and U13533 (N_13533,N_10709,N_10422);
nand U13534 (N_13534,N_11363,N_12432);
nor U13535 (N_13535,N_10154,N_12292);
xor U13536 (N_13536,N_11870,N_11470);
nor U13537 (N_13537,N_11629,N_10919);
or U13538 (N_13538,N_11801,N_10821);
nor U13539 (N_13539,N_12319,N_12108);
xnor U13540 (N_13540,N_12458,N_11979);
xnor U13541 (N_13541,N_10186,N_10568);
and U13542 (N_13542,N_10846,N_11795);
and U13543 (N_13543,N_11948,N_10761);
or U13544 (N_13544,N_11148,N_11417);
or U13545 (N_13545,N_11368,N_12158);
xor U13546 (N_13546,N_11855,N_11732);
nor U13547 (N_13547,N_10236,N_11653);
or U13548 (N_13548,N_12449,N_12451);
nand U13549 (N_13549,N_11831,N_11890);
and U13550 (N_13550,N_10074,N_10031);
nor U13551 (N_13551,N_12335,N_12340);
xor U13552 (N_13552,N_11187,N_12318);
nor U13553 (N_13553,N_11369,N_11908);
xnor U13554 (N_13554,N_10340,N_10633);
and U13555 (N_13555,N_12027,N_10694);
or U13556 (N_13556,N_10873,N_12237);
and U13557 (N_13557,N_10035,N_12233);
and U13558 (N_13558,N_11646,N_12153);
or U13559 (N_13559,N_11551,N_12299);
nor U13560 (N_13560,N_12160,N_10392);
xnor U13561 (N_13561,N_11961,N_11929);
nand U13562 (N_13562,N_11477,N_11683);
nor U13563 (N_13563,N_10955,N_10288);
and U13564 (N_13564,N_12115,N_11662);
nor U13565 (N_13565,N_10907,N_10447);
xnor U13566 (N_13566,N_11497,N_11682);
xor U13567 (N_13567,N_12271,N_10587);
or U13568 (N_13568,N_10165,N_12220);
nor U13569 (N_13569,N_10358,N_10892);
and U13570 (N_13570,N_11960,N_11738);
nand U13571 (N_13571,N_12404,N_11898);
nor U13572 (N_13572,N_10381,N_10342);
nand U13573 (N_13573,N_10401,N_11943);
nand U13574 (N_13574,N_10293,N_10400);
xnor U13575 (N_13575,N_10915,N_11474);
and U13576 (N_13576,N_11544,N_10600);
and U13577 (N_13577,N_11125,N_12437);
nand U13578 (N_13578,N_11745,N_10219);
nor U13579 (N_13579,N_10197,N_10022);
or U13580 (N_13580,N_10171,N_11993);
nor U13581 (N_13581,N_10747,N_12475);
xor U13582 (N_13582,N_10552,N_12277);
and U13583 (N_13583,N_11752,N_10516);
xor U13584 (N_13584,N_10699,N_11641);
and U13585 (N_13585,N_10848,N_12315);
or U13586 (N_13586,N_12287,N_11643);
and U13587 (N_13587,N_10144,N_11432);
or U13588 (N_13588,N_12330,N_12004);
nand U13589 (N_13589,N_12470,N_10318);
xnor U13590 (N_13590,N_12273,N_12253);
or U13591 (N_13591,N_12056,N_11354);
nand U13592 (N_13592,N_11974,N_10133);
or U13593 (N_13593,N_10304,N_11027);
xor U13594 (N_13594,N_12422,N_11780);
xnor U13595 (N_13595,N_11440,N_10963);
nor U13596 (N_13596,N_10762,N_11213);
xor U13597 (N_13597,N_11128,N_12003);
nand U13598 (N_13598,N_11506,N_11915);
or U13599 (N_13599,N_10972,N_11521);
xnor U13600 (N_13600,N_10834,N_11091);
nor U13601 (N_13601,N_10824,N_10013);
xor U13602 (N_13602,N_12399,N_12329);
nor U13603 (N_13603,N_11986,N_10349);
nor U13604 (N_13604,N_10800,N_12162);
nor U13605 (N_13605,N_11503,N_10446);
xor U13606 (N_13606,N_10029,N_10399);
nand U13607 (N_13607,N_10023,N_11998);
nand U13608 (N_13608,N_12234,N_11287);
and U13609 (N_13609,N_10172,N_12131);
xnor U13610 (N_13610,N_12031,N_10511);
nand U13611 (N_13611,N_11768,N_11862);
nand U13612 (N_13612,N_10499,N_12408);
nor U13613 (N_13613,N_11294,N_11534);
nand U13614 (N_13614,N_10493,N_11689);
nand U13615 (N_13615,N_11303,N_12061);
and U13616 (N_13616,N_10959,N_12134);
or U13617 (N_13617,N_11573,N_12085);
nand U13618 (N_13618,N_11946,N_10124);
nand U13619 (N_13619,N_12286,N_10098);
nor U13620 (N_13620,N_10174,N_10756);
or U13621 (N_13621,N_12366,N_11471);
xnor U13622 (N_13622,N_10004,N_10459);
or U13623 (N_13623,N_12307,N_11896);
xor U13624 (N_13624,N_12395,N_11533);
nor U13625 (N_13625,N_10321,N_11881);
and U13626 (N_13626,N_11967,N_12484);
and U13627 (N_13627,N_11415,N_10367);
xnor U13628 (N_13628,N_11635,N_11820);
xnor U13629 (N_13629,N_11073,N_11249);
and U13630 (N_13630,N_11118,N_10176);
and U13631 (N_13631,N_10854,N_10656);
or U13632 (N_13632,N_12405,N_11043);
and U13633 (N_13633,N_11264,N_11028);
or U13634 (N_13634,N_11255,N_12494);
xor U13635 (N_13635,N_12032,N_12396);
xnor U13636 (N_13636,N_10720,N_11543);
nor U13637 (N_13637,N_11070,N_11479);
nor U13638 (N_13638,N_10469,N_11337);
nor U13639 (N_13639,N_12337,N_12026);
nor U13640 (N_13640,N_11064,N_10207);
nor U13641 (N_13641,N_11913,N_10865);
nor U13642 (N_13642,N_10214,N_12165);
xnor U13643 (N_13643,N_10671,N_10943);
nand U13644 (N_13644,N_12045,N_11424);
or U13645 (N_13645,N_10920,N_10042);
or U13646 (N_13646,N_10909,N_10930);
xor U13647 (N_13647,N_11382,N_11280);
nand U13648 (N_13648,N_11078,N_11697);
or U13649 (N_13649,N_11032,N_12099);
nor U13650 (N_13650,N_10514,N_11155);
and U13651 (N_13651,N_11464,N_11390);
xor U13652 (N_13652,N_10085,N_10312);
and U13653 (N_13653,N_10428,N_10468);
nand U13654 (N_13654,N_12348,N_10379);
or U13655 (N_13655,N_11004,N_10352);
nor U13656 (N_13656,N_10701,N_10586);
xnor U13657 (N_13657,N_11283,N_11176);
nor U13658 (N_13658,N_11843,N_10678);
nand U13659 (N_13659,N_11000,N_11901);
or U13660 (N_13660,N_10524,N_11230);
nand U13661 (N_13661,N_11040,N_10485);
nor U13662 (N_13662,N_10790,N_12228);
nand U13663 (N_13663,N_10991,N_10385);
or U13664 (N_13664,N_10949,N_10989);
and U13665 (N_13665,N_10649,N_11705);
and U13666 (N_13666,N_12462,N_10620);
nor U13667 (N_13667,N_10594,N_11518);
xor U13668 (N_13668,N_11978,N_10841);
xor U13669 (N_13669,N_12403,N_12447);
or U13670 (N_13670,N_11339,N_11406);
xnor U13671 (N_13671,N_11357,N_10003);
xor U13672 (N_13672,N_11002,N_10464);
nand U13673 (N_13673,N_11347,N_12147);
xor U13674 (N_13674,N_11631,N_10812);
nor U13675 (N_13675,N_11166,N_10298);
xnor U13676 (N_13676,N_10391,N_10830);
nand U13677 (N_13677,N_12222,N_10657);
and U13678 (N_13678,N_10284,N_10109);
xor U13679 (N_13679,N_12464,N_10698);
nor U13680 (N_13680,N_11445,N_11566);
or U13681 (N_13681,N_10601,N_12095);
xnor U13682 (N_13682,N_10545,N_12411);
and U13683 (N_13683,N_11130,N_12262);
xor U13684 (N_13684,N_11746,N_12110);
nor U13685 (N_13685,N_10535,N_11523);
and U13686 (N_13686,N_10200,N_10603);
nand U13687 (N_13687,N_10364,N_10272);
or U13688 (N_13688,N_10413,N_10347);
nor U13689 (N_13689,N_11575,N_10713);
xnor U13690 (N_13690,N_12371,N_10301);
and U13691 (N_13691,N_10196,N_12471);
or U13692 (N_13692,N_12118,N_10481);
xnor U13693 (N_13693,N_11465,N_11253);
nand U13694 (N_13694,N_12150,N_10444);
nand U13695 (N_13695,N_10998,N_10059);
nand U13696 (N_13696,N_10343,N_10140);
nand U13697 (N_13697,N_11931,N_12145);
and U13698 (N_13698,N_10782,N_10822);
or U13699 (N_13699,N_11599,N_12137);
xor U13700 (N_13700,N_11588,N_10087);
nor U13701 (N_13701,N_12144,N_11604);
and U13702 (N_13702,N_11116,N_12202);
nor U13703 (N_13703,N_11392,N_11714);
nor U13704 (N_13704,N_10040,N_11658);
nor U13705 (N_13705,N_10235,N_11112);
nor U13706 (N_13706,N_10083,N_10810);
nor U13707 (N_13707,N_10666,N_11618);
nor U13708 (N_13708,N_11182,N_10107);
nor U13709 (N_13709,N_10111,N_11684);
and U13710 (N_13710,N_11661,N_10710);
or U13711 (N_13711,N_11221,N_11076);
nor U13712 (N_13712,N_12392,N_10544);
nor U13713 (N_13713,N_11488,N_10238);
nand U13714 (N_13714,N_10847,N_10806);
and U13715 (N_13715,N_12261,N_11893);
xor U13716 (N_13716,N_10116,N_10752);
nor U13717 (N_13717,N_10078,N_11647);
and U13718 (N_13718,N_11001,N_11081);
xor U13719 (N_13719,N_10063,N_10396);
nor U13720 (N_13720,N_12111,N_11666);
or U13721 (N_13721,N_12046,N_12142);
or U13722 (N_13722,N_11748,N_11567);
nor U13723 (N_13723,N_12491,N_11393);
nand U13724 (N_13724,N_11914,N_10664);
nand U13725 (N_13725,N_11285,N_10239);
nand U13726 (N_13726,N_11013,N_11809);
xor U13727 (N_13727,N_12200,N_11225);
or U13728 (N_13728,N_12465,N_10862);
and U13729 (N_13729,N_11137,N_12483);
or U13730 (N_13730,N_11976,N_11516);
nand U13731 (N_13731,N_11361,N_11891);
nor U13732 (N_13732,N_10141,N_10517);
nor U13733 (N_13733,N_11486,N_11792);
nor U13734 (N_13734,N_10047,N_11063);
xor U13735 (N_13735,N_11377,N_11607);
nand U13736 (N_13736,N_11671,N_12388);
nand U13737 (N_13737,N_10952,N_12397);
nand U13738 (N_13738,N_11223,N_12457);
or U13739 (N_13739,N_10104,N_10205);
or U13740 (N_13740,N_11718,N_11328);
xnor U13741 (N_13741,N_11052,N_10194);
and U13742 (N_13742,N_12104,N_12082);
xnor U13743 (N_13743,N_12067,N_10158);
and U13744 (N_13744,N_11096,N_10674);
or U13745 (N_13745,N_11556,N_10335);
nand U13746 (N_13746,N_10851,N_11158);
nand U13747 (N_13747,N_12179,N_10242);
nand U13748 (N_13748,N_10265,N_11135);
nor U13749 (N_13749,N_12130,N_12048);
xor U13750 (N_13750,N_11618,N_11664);
nand U13751 (N_13751,N_11737,N_12306);
and U13752 (N_13752,N_10257,N_12341);
xor U13753 (N_13753,N_10789,N_11856);
and U13754 (N_13754,N_12036,N_11741);
nand U13755 (N_13755,N_12161,N_10355);
xnor U13756 (N_13756,N_12239,N_11149);
and U13757 (N_13757,N_11563,N_10573);
or U13758 (N_13758,N_11150,N_10288);
nor U13759 (N_13759,N_11120,N_11517);
or U13760 (N_13760,N_11486,N_10710);
and U13761 (N_13761,N_10910,N_11970);
or U13762 (N_13762,N_10098,N_10996);
and U13763 (N_13763,N_10159,N_11611);
nand U13764 (N_13764,N_11005,N_11333);
nand U13765 (N_13765,N_10105,N_10009);
or U13766 (N_13766,N_11248,N_10542);
xnor U13767 (N_13767,N_10659,N_12090);
or U13768 (N_13768,N_10639,N_10500);
xnor U13769 (N_13769,N_11909,N_10905);
nand U13770 (N_13770,N_12328,N_12095);
and U13771 (N_13771,N_10122,N_10142);
and U13772 (N_13772,N_12224,N_12306);
xor U13773 (N_13773,N_11233,N_11523);
nand U13774 (N_13774,N_10634,N_10477);
xor U13775 (N_13775,N_10567,N_10872);
and U13776 (N_13776,N_10691,N_11110);
or U13777 (N_13777,N_11913,N_11521);
nor U13778 (N_13778,N_10281,N_10616);
or U13779 (N_13779,N_12237,N_11414);
and U13780 (N_13780,N_12387,N_10251);
nor U13781 (N_13781,N_11574,N_12381);
nand U13782 (N_13782,N_12362,N_11268);
or U13783 (N_13783,N_11274,N_11171);
or U13784 (N_13784,N_12463,N_11918);
and U13785 (N_13785,N_10690,N_11324);
and U13786 (N_13786,N_10263,N_11001);
or U13787 (N_13787,N_11538,N_10695);
or U13788 (N_13788,N_10623,N_10496);
or U13789 (N_13789,N_10798,N_12444);
xnor U13790 (N_13790,N_10977,N_10030);
nor U13791 (N_13791,N_10573,N_10628);
nor U13792 (N_13792,N_10868,N_12100);
nor U13793 (N_13793,N_11934,N_11175);
xor U13794 (N_13794,N_10566,N_11732);
and U13795 (N_13795,N_11692,N_10069);
xor U13796 (N_13796,N_12051,N_10951);
nand U13797 (N_13797,N_12107,N_10377);
or U13798 (N_13798,N_11989,N_11894);
nor U13799 (N_13799,N_10063,N_11429);
or U13800 (N_13800,N_12328,N_11773);
and U13801 (N_13801,N_11096,N_12325);
and U13802 (N_13802,N_10487,N_10952);
or U13803 (N_13803,N_10490,N_10967);
nor U13804 (N_13804,N_10996,N_12452);
xnor U13805 (N_13805,N_11406,N_10041);
xnor U13806 (N_13806,N_12004,N_12169);
or U13807 (N_13807,N_11995,N_10938);
and U13808 (N_13808,N_10783,N_12342);
or U13809 (N_13809,N_10464,N_11368);
nand U13810 (N_13810,N_11558,N_10234);
nor U13811 (N_13811,N_10720,N_11200);
or U13812 (N_13812,N_11862,N_11014);
and U13813 (N_13813,N_11483,N_11907);
nor U13814 (N_13814,N_10530,N_10422);
nor U13815 (N_13815,N_12148,N_11008);
nand U13816 (N_13816,N_10454,N_12325);
nor U13817 (N_13817,N_10315,N_11295);
nor U13818 (N_13818,N_10574,N_12448);
or U13819 (N_13819,N_12124,N_10643);
xor U13820 (N_13820,N_12151,N_11441);
or U13821 (N_13821,N_11181,N_10092);
nor U13822 (N_13822,N_12106,N_10976);
and U13823 (N_13823,N_10258,N_11165);
or U13824 (N_13824,N_11392,N_10974);
or U13825 (N_13825,N_12309,N_12198);
xnor U13826 (N_13826,N_10851,N_10342);
or U13827 (N_13827,N_11309,N_11379);
or U13828 (N_13828,N_10519,N_10065);
xnor U13829 (N_13829,N_11060,N_10373);
and U13830 (N_13830,N_12125,N_10140);
xor U13831 (N_13831,N_12153,N_11106);
nor U13832 (N_13832,N_10052,N_10253);
nor U13833 (N_13833,N_11183,N_10412);
or U13834 (N_13834,N_11121,N_10701);
and U13835 (N_13835,N_11673,N_10095);
or U13836 (N_13836,N_11136,N_11338);
nor U13837 (N_13837,N_10886,N_11925);
and U13838 (N_13838,N_11401,N_10183);
nand U13839 (N_13839,N_11478,N_11929);
nor U13840 (N_13840,N_10384,N_12137);
nor U13841 (N_13841,N_12101,N_12139);
nor U13842 (N_13842,N_10807,N_10609);
xnor U13843 (N_13843,N_10181,N_10620);
nand U13844 (N_13844,N_11638,N_11506);
nor U13845 (N_13845,N_11716,N_10180);
nor U13846 (N_13846,N_10856,N_12057);
xnor U13847 (N_13847,N_12059,N_11067);
xor U13848 (N_13848,N_10129,N_12411);
and U13849 (N_13849,N_10239,N_11589);
nand U13850 (N_13850,N_10846,N_12309);
xnor U13851 (N_13851,N_10284,N_10817);
nor U13852 (N_13852,N_12416,N_12094);
nor U13853 (N_13853,N_11873,N_12153);
and U13854 (N_13854,N_10001,N_10443);
nor U13855 (N_13855,N_11258,N_10313);
and U13856 (N_13856,N_12399,N_12304);
or U13857 (N_13857,N_11245,N_11817);
and U13858 (N_13858,N_10716,N_11214);
or U13859 (N_13859,N_10250,N_10524);
nand U13860 (N_13860,N_10921,N_11503);
and U13861 (N_13861,N_10142,N_11123);
xor U13862 (N_13862,N_10647,N_12265);
nor U13863 (N_13863,N_10354,N_11005);
and U13864 (N_13864,N_12296,N_10584);
xnor U13865 (N_13865,N_11000,N_11736);
and U13866 (N_13866,N_12238,N_10532);
or U13867 (N_13867,N_11944,N_10203);
or U13868 (N_13868,N_11235,N_11018);
nand U13869 (N_13869,N_10322,N_11347);
nand U13870 (N_13870,N_10736,N_11144);
and U13871 (N_13871,N_10395,N_10193);
xor U13872 (N_13872,N_11504,N_10583);
xnor U13873 (N_13873,N_11505,N_11226);
xnor U13874 (N_13874,N_11181,N_11839);
or U13875 (N_13875,N_10513,N_11240);
and U13876 (N_13876,N_10215,N_10515);
and U13877 (N_13877,N_10106,N_12449);
xnor U13878 (N_13878,N_10610,N_11254);
xnor U13879 (N_13879,N_12322,N_12037);
nor U13880 (N_13880,N_12240,N_11451);
xnor U13881 (N_13881,N_12427,N_12199);
or U13882 (N_13882,N_11857,N_10446);
nor U13883 (N_13883,N_10593,N_11479);
nor U13884 (N_13884,N_10966,N_10855);
and U13885 (N_13885,N_10216,N_10314);
xnor U13886 (N_13886,N_12118,N_10792);
xnor U13887 (N_13887,N_10809,N_11740);
nand U13888 (N_13888,N_11377,N_11208);
nor U13889 (N_13889,N_11815,N_10826);
nand U13890 (N_13890,N_11982,N_10337);
xnor U13891 (N_13891,N_10402,N_12355);
xnor U13892 (N_13892,N_11234,N_10076);
xnor U13893 (N_13893,N_10281,N_11247);
nor U13894 (N_13894,N_11320,N_12437);
or U13895 (N_13895,N_11795,N_10772);
nor U13896 (N_13896,N_10585,N_11671);
or U13897 (N_13897,N_10564,N_12174);
or U13898 (N_13898,N_12412,N_10471);
xnor U13899 (N_13899,N_10835,N_10536);
or U13900 (N_13900,N_10517,N_12211);
and U13901 (N_13901,N_10416,N_11933);
or U13902 (N_13902,N_12445,N_11167);
nand U13903 (N_13903,N_12279,N_11500);
nor U13904 (N_13904,N_10030,N_11281);
xnor U13905 (N_13905,N_10793,N_11095);
xnor U13906 (N_13906,N_10205,N_12341);
nor U13907 (N_13907,N_11911,N_12498);
xnor U13908 (N_13908,N_12270,N_10141);
and U13909 (N_13909,N_11324,N_12408);
nor U13910 (N_13910,N_10583,N_11484);
nor U13911 (N_13911,N_10671,N_10732);
and U13912 (N_13912,N_10890,N_10755);
and U13913 (N_13913,N_10842,N_11252);
or U13914 (N_13914,N_11011,N_10961);
xor U13915 (N_13915,N_11189,N_11855);
or U13916 (N_13916,N_11068,N_11336);
or U13917 (N_13917,N_10288,N_12163);
xor U13918 (N_13918,N_11316,N_12414);
and U13919 (N_13919,N_10503,N_10343);
or U13920 (N_13920,N_11902,N_10379);
nand U13921 (N_13921,N_11222,N_12308);
or U13922 (N_13922,N_11566,N_10150);
and U13923 (N_13923,N_10753,N_10401);
or U13924 (N_13924,N_12459,N_10625);
and U13925 (N_13925,N_10700,N_11830);
nand U13926 (N_13926,N_12455,N_12320);
xnor U13927 (N_13927,N_11021,N_11188);
nor U13928 (N_13928,N_11539,N_10307);
and U13929 (N_13929,N_12276,N_10035);
nand U13930 (N_13930,N_11777,N_10365);
nand U13931 (N_13931,N_12493,N_10888);
xnor U13932 (N_13932,N_10706,N_11208);
nand U13933 (N_13933,N_10044,N_11112);
and U13934 (N_13934,N_11222,N_11395);
or U13935 (N_13935,N_12045,N_10192);
nor U13936 (N_13936,N_12382,N_10843);
and U13937 (N_13937,N_12145,N_12248);
or U13938 (N_13938,N_10300,N_10266);
xor U13939 (N_13939,N_12216,N_10649);
and U13940 (N_13940,N_11940,N_11888);
nor U13941 (N_13941,N_10640,N_10371);
nand U13942 (N_13942,N_11988,N_10044);
nor U13943 (N_13943,N_10785,N_11940);
xor U13944 (N_13944,N_11965,N_10259);
nand U13945 (N_13945,N_11990,N_10969);
xnor U13946 (N_13946,N_11771,N_12369);
nand U13947 (N_13947,N_12258,N_11734);
nor U13948 (N_13948,N_11692,N_11815);
and U13949 (N_13949,N_11972,N_11166);
nand U13950 (N_13950,N_10909,N_10305);
nand U13951 (N_13951,N_10364,N_10619);
nand U13952 (N_13952,N_11222,N_12195);
nand U13953 (N_13953,N_12012,N_12319);
or U13954 (N_13954,N_11799,N_10026);
xor U13955 (N_13955,N_10342,N_10789);
or U13956 (N_13956,N_11391,N_10450);
or U13957 (N_13957,N_11435,N_10316);
xor U13958 (N_13958,N_10196,N_10144);
or U13959 (N_13959,N_10547,N_11269);
and U13960 (N_13960,N_10128,N_11304);
or U13961 (N_13961,N_12080,N_10149);
or U13962 (N_13962,N_11281,N_10059);
or U13963 (N_13963,N_11812,N_12184);
or U13964 (N_13964,N_10401,N_10250);
and U13965 (N_13965,N_12382,N_11246);
nand U13966 (N_13966,N_10422,N_10168);
and U13967 (N_13967,N_11636,N_12226);
nor U13968 (N_13968,N_10756,N_10105);
and U13969 (N_13969,N_10163,N_11573);
and U13970 (N_13970,N_11465,N_11286);
xnor U13971 (N_13971,N_10580,N_11368);
xnor U13972 (N_13972,N_10911,N_10481);
or U13973 (N_13973,N_11355,N_10519);
xnor U13974 (N_13974,N_11925,N_12432);
nand U13975 (N_13975,N_11713,N_12456);
or U13976 (N_13976,N_11450,N_11237);
or U13977 (N_13977,N_11317,N_12245);
nand U13978 (N_13978,N_10583,N_10367);
and U13979 (N_13979,N_11540,N_10539);
xnor U13980 (N_13980,N_12242,N_10922);
nand U13981 (N_13981,N_11876,N_12268);
or U13982 (N_13982,N_11515,N_10307);
or U13983 (N_13983,N_10699,N_10114);
or U13984 (N_13984,N_12145,N_12211);
and U13985 (N_13985,N_12232,N_10708);
nand U13986 (N_13986,N_12039,N_12338);
nand U13987 (N_13987,N_11449,N_12065);
xnor U13988 (N_13988,N_11707,N_10352);
and U13989 (N_13989,N_10002,N_11472);
nand U13990 (N_13990,N_10499,N_12212);
xor U13991 (N_13991,N_12114,N_10604);
nor U13992 (N_13992,N_10217,N_10535);
xor U13993 (N_13993,N_12014,N_11088);
nand U13994 (N_13994,N_11448,N_10996);
nor U13995 (N_13995,N_11543,N_11733);
and U13996 (N_13996,N_11398,N_11361);
nand U13997 (N_13997,N_10928,N_11245);
nor U13998 (N_13998,N_12376,N_11573);
and U13999 (N_13999,N_11477,N_10827);
nor U14000 (N_14000,N_10788,N_11865);
and U14001 (N_14001,N_11427,N_11785);
and U14002 (N_14002,N_10654,N_10997);
nand U14003 (N_14003,N_11882,N_11761);
xnor U14004 (N_14004,N_11776,N_12312);
xor U14005 (N_14005,N_11393,N_11614);
or U14006 (N_14006,N_11525,N_12265);
nor U14007 (N_14007,N_11812,N_11624);
and U14008 (N_14008,N_12490,N_12475);
and U14009 (N_14009,N_10652,N_11119);
nor U14010 (N_14010,N_11760,N_10003);
xor U14011 (N_14011,N_12300,N_10095);
nand U14012 (N_14012,N_11405,N_11199);
xor U14013 (N_14013,N_10631,N_12005);
nor U14014 (N_14014,N_10147,N_11846);
nand U14015 (N_14015,N_12197,N_11265);
nand U14016 (N_14016,N_10461,N_11351);
nor U14017 (N_14017,N_11591,N_10553);
nand U14018 (N_14018,N_10113,N_10746);
or U14019 (N_14019,N_11866,N_11002);
xnor U14020 (N_14020,N_10854,N_11124);
nor U14021 (N_14021,N_11397,N_10136);
xor U14022 (N_14022,N_11451,N_11640);
nand U14023 (N_14023,N_12186,N_11525);
nand U14024 (N_14024,N_10883,N_10763);
or U14025 (N_14025,N_10317,N_11814);
or U14026 (N_14026,N_11687,N_12308);
or U14027 (N_14027,N_11064,N_10089);
xnor U14028 (N_14028,N_10995,N_10877);
and U14029 (N_14029,N_10075,N_10562);
or U14030 (N_14030,N_10207,N_10909);
nand U14031 (N_14031,N_11027,N_11263);
nand U14032 (N_14032,N_10981,N_10518);
and U14033 (N_14033,N_12067,N_12274);
nor U14034 (N_14034,N_12062,N_11604);
nand U14035 (N_14035,N_10590,N_12413);
nor U14036 (N_14036,N_10776,N_11398);
xnor U14037 (N_14037,N_11203,N_11356);
xnor U14038 (N_14038,N_11888,N_10045);
nor U14039 (N_14039,N_12076,N_12436);
nor U14040 (N_14040,N_11917,N_10562);
nand U14041 (N_14041,N_11605,N_11249);
and U14042 (N_14042,N_11198,N_12361);
nand U14043 (N_14043,N_12170,N_11560);
xor U14044 (N_14044,N_12277,N_10819);
nand U14045 (N_14045,N_10438,N_12250);
nor U14046 (N_14046,N_10857,N_10635);
nor U14047 (N_14047,N_10670,N_10512);
nor U14048 (N_14048,N_11904,N_11154);
xnor U14049 (N_14049,N_10393,N_11488);
xor U14050 (N_14050,N_12216,N_11977);
xnor U14051 (N_14051,N_11594,N_11148);
and U14052 (N_14052,N_11309,N_11033);
and U14053 (N_14053,N_11046,N_10179);
nand U14054 (N_14054,N_12470,N_10734);
nand U14055 (N_14055,N_11249,N_10498);
xor U14056 (N_14056,N_10164,N_10340);
xnor U14057 (N_14057,N_10247,N_11266);
and U14058 (N_14058,N_11093,N_12490);
nand U14059 (N_14059,N_10647,N_11787);
nor U14060 (N_14060,N_12131,N_11031);
nor U14061 (N_14061,N_11223,N_10640);
nand U14062 (N_14062,N_10605,N_12311);
xor U14063 (N_14063,N_11901,N_11698);
nand U14064 (N_14064,N_10172,N_11585);
or U14065 (N_14065,N_10950,N_11837);
xor U14066 (N_14066,N_11974,N_12377);
nand U14067 (N_14067,N_10385,N_12352);
and U14068 (N_14068,N_10127,N_11040);
nand U14069 (N_14069,N_10332,N_10744);
nor U14070 (N_14070,N_10340,N_11967);
nor U14071 (N_14071,N_11827,N_11574);
xnor U14072 (N_14072,N_10339,N_11966);
nand U14073 (N_14073,N_12143,N_10129);
nor U14074 (N_14074,N_10957,N_10703);
nand U14075 (N_14075,N_10739,N_12139);
nor U14076 (N_14076,N_11893,N_10879);
nand U14077 (N_14077,N_10640,N_12365);
and U14078 (N_14078,N_12211,N_11923);
or U14079 (N_14079,N_11211,N_11406);
xnor U14080 (N_14080,N_11243,N_12426);
xor U14081 (N_14081,N_11400,N_10379);
nand U14082 (N_14082,N_10935,N_12232);
xor U14083 (N_14083,N_11919,N_11804);
nor U14084 (N_14084,N_10698,N_12112);
xnor U14085 (N_14085,N_10296,N_10352);
nand U14086 (N_14086,N_12417,N_12241);
and U14087 (N_14087,N_11531,N_11527);
xnor U14088 (N_14088,N_10994,N_11629);
xor U14089 (N_14089,N_10367,N_10165);
or U14090 (N_14090,N_10573,N_12478);
nor U14091 (N_14091,N_12202,N_12321);
xor U14092 (N_14092,N_12179,N_11847);
nand U14093 (N_14093,N_11562,N_10569);
nor U14094 (N_14094,N_11076,N_11540);
xnor U14095 (N_14095,N_10999,N_11308);
nor U14096 (N_14096,N_10044,N_11573);
or U14097 (N_14097,N_11085,N_11467);
or U14098 (N_14098,N_12143,N_11210);
nand U14099 (N_14099,N_12126,N_10956);
nand U14100 (N_14100,N_11778,N_10406);
and U14101 (N_14101,N_12467,N_10703);
nand U14102 (N_14102,N_12357,N_12288);
nand U14103 (N_14103,N_11100,N_10568);
nand U14104 (N_14104,N_10625,N_11191);
xor U14105 (N_14105,N_10072,N_10491);
xnor U14106 (N_14106,N_11964,N_10050);
nor U14107 (N_14107,N_11451,N_11128);
xnor U14108 (N_14108,N_12141,N_11908);
nor U14109 (N_14109,N_11241,N_12247);
nand U14110 (N_14110,N_11885,N_11994);
xor U14111 (N_14111,N_12318,N_12139);
nand U14112 (N_14112,N_10282,N_10828);
nor U14113 (N_14113,N_11884,N_10342);
nand U14114 (N_14114,N_12338,N_10643);
nand U14115 (N_14115,N_12262,N_10552);
xnor U14116 (N_14116,N_11813,N_10163);
nor U14117 (N_14117,N_11898,N_12405);
and U14118 (N_14118,N_11051,N_12013);
or U14119 (N_14119,N_10135,N_10148);
nand U14120 (N_14120,N_10657,N_12429);
nor U14121 (N_14121,N_10060,N_11576);
and U14122 (N_14122,N_11240,N_11167);
or U14123 (N_14123,N_12013,N_10472);
nand U14124 (N_14124,N_10329,N_11220);
nor U14125 (N_14125,N_10762,N_10896);
or U14126 (N_14126,N_11313,N_11153);
nor U14127 (N_14127,N_10477,N_12401);
xor U14128 (N_14128,N_11265,N_12424);
nor U14129 (N_14129,N_10551,N_12169);
and U14130 (N_14130,N_10536,N_10200);
or U14131 (N_14131,N_10956,N_12386);
nor U14132 (N_14132,N_12450,N_11939);
nor U14133 (N_14133,N_11464,N_10947);
xnor U14134 (N_14134,N_11421,N_10009);
xor U14135 (N_14135,N_12301,N_12228);
nand U14136 (N_14136,N_10227,N_11858);
nand U14137 (N_14137,N_10989,N_12337);
xnor U14138 (N_14138,N_11335,N_11225);
xor U14139 (N_14139,N_10107,N_11570);
and U14140 (N_14140,N_11906,N_10965);
xnor U14141 (N_14141,N_11172,N_10086);
nor U14142 (N_14142,N_10901,N_10629);
and U14143 (N_14143,N_11863,N_11804);
xnor U14144 (N_14144,N_12087,N_11359);
or U14145 (N_14145,N_10555,N_11328);
or U14146 (N_14146,N_11999,N_12465);
nand U14147 (N_14147,N_12427,N_11568);
nor U14148 (N_14148,N_11601,N_11884);
xnor U14149 (N_14149,N_10203,N_10184);
nand U14150 (N_14150,N_11382,N_12059);
and U14151 (N_14151,N_12240,N_10993);
and U14152 (N_14152,N_11230,N_11254);
xor U14153 (N_14153,N_11751,N_11003);
and U14154 (N_14154,N_11208,N_11712);
nor U14155 (N_14155,N_11053,N_12289);
or U14156 (N_14156,N_12180,N_11243);
or U14157 (N_14157,N_10991,N_11303);
or U14158 (N_14158,N_10833,N_12155);
nor U14159 (N_14159,N_12038,N_12473);
or U14160 (N_14160,N_11223,N_11980);
nor U14161 (N_14161,N_10771,N_12447);
xnor U14162 (N_14162,N_11518,N_10818);
and U14163 (N_14163,N_10773,N_12487);
nor U14164 (N_14164,N_10552,N_12104);
nor U14165 (N_14165,N_11360,N_11793);
xnor U14166 (N_14166,N_10309,N_11266);
and U14167 (N_14167,N_11927,N_10187);
and U14168 (N_14168,N_10429,N_12374);
nor U14169 (N_14169,N_10436,N_11781);
nor U14170 (N_14170,N_10786,N_11984);
nand U14171 (N_14171,N_11345,N_11999);
and U14172 (N_14172,N_11201,N_10418);
nor U14173 (N_14173,N_11591,N_10674);
xnor U14174 (N_14174,N_10804,N_11781);
nor U14175 (N_14175,N_10369,N_11764);
nand U14176 (N_14176,N_11517,N_10860);
and U14177 (N_14177,N_12128,N_11925);
or U14178 (N_14178,N_10945,N_11438);
xor U14179 (N_14179,N_12043,N_12298);
nand U14180 (N_14180,N_11346,N_11171);
nor U14181 (N_14181,N_12373,N_10023);
and U14182 (N_14182,N_12332,N_12483);
xor U14183 (N_14183,N_11955,N_11424);
and U14184 (N_14184,N_12046,N_11866);
or U14185 (N_14185,N_12114,N_11695);
and U14186 (N_14186,N_11555,N_10957);
xor U14187 (N_14187,N_11827,N_11704);
or U14188 (N_14188,N_11024,N_10631);
and U14189 (N_14189,N_11937,N_12322);
and U14190 (N_14190,N_11398,N_11219);
and U14191 (N_14191,N_12265,N_10096);
nor U14192 (N_14192,N_10523,N_10953);
nand U14193 (N_14193,N_11746,N_11566);
xor U14194 (N_14194,N_10658,N_11041);
or U14195 (N_14195,N_11983,N_11694);
or U14196 (N_14196,N_11657,N_11266);
nor U14197 (N_14197,N_11490,N_11904);
nand U14198 (N_14198,N_10754,N_12448);
nand U14199 (N_14199,N_11257,N_10519);
or U14200 (N_14200,N_12137,N_11573);
and U14201 (N_14201,N_10613,N_10763);
nand U14202 (N_14202,N_12453,N_10500);
or U14203 (N_14203,N_11577,N_10804);
or U14204 (N_14204,N_10514,N_12333);
nor U14205 (N_14205,N_11579,N_12306);
nor U14206 (N_14206,N_10002,N_10985);
nand U14207 (N_14207,N_10457,N_12152);
or U14208 (N_14208,N_10407,N_10428);
or U14209 (N_14209,N_11526,N_12110);
nand U14210 (N_14210,N_12438,N_12330);
and U14211 (N_14211,N_11037,N_10223);
nor U14212 (N_14212,N_10373,N_11821);
or U14213 (N_14213,N_10361,N_10664);
xor U14214 (N_14214,N_10296,N_11857);
nor U14215 (N_14215,N_12492,N_10530);
xor U14216 (N_14216,N_11210,N_11729);
or U14217 (N_14217,N_11442,N_10610);
and U14218 (N_14218,N_10739,N_11803);
xnor U14219 (N_14219,N_11900,N_11460);
or U14220 (N_14220,N_10385,N_11722);
or U14221 (N_14221,N_10685,N_11519);
xor U14222 (N_14222,N_10932,N_11163);
nor U14223 (N_14223,N_12055,N_10142);
xor U14224 (N_14224,N_10170,N_12065);
or U14225 (N_14225,N_11238,N_10629);
or U14226 (N_14226,N_10446,N_12287);
or U14227 (N_14227,N_12427,N_10789);
or U14228 (N_14228,N_10409,N_11023);
nor U14229 (N_14229,N_11914,N_10862);
or U14230 (N_14230,N_12130,N_11739);
nand U14231 (N_14231,N_11062,N_11268);
or U14232 (N_14232,N_10898,N_10239);
nor U14233 (N_14233,N_10016,N_11936);
and U14234 (N_14234,N_12146,N_11398);
xor U14235 (N_14235,N_10611,N_12331);
or U14236 (N_14236,N_11514,N_11759);
or U14237 (N_14237,N_10423,N_12132);
xor U14238 (N_14238,N_12416,N_11633);
or U14239 (N_14239,N_11185,N_10986);
nor U14240 (N_14240,N_12084,N_10152);
or U14241 (N_14241,N_12373,N_11334);
nor U14242 (N_14242,N_11189,N_11645);
xor U14243 (N_14243,N_10722,N_12034);
or U14244 (N_14244,N_12179,N_12127);
nor U14245 (N_14245,N_11806,N_11373);
nor U14246 (N_14246,N_11865,N_10084);
and U14247 (N_14247,N_10149,N_10264);
nand U14248 (N_14248,N_12262,N_12097);
or U14249 (N_14249,N_12275,N_12001);
or U14250 (N_14250,N_12463,N_11775);
xor U14251 (N_14251,N_12290,N_10903);
nor U14252 (N_14252,N_11543,N_11497);
or U14253 (N_14253,N_11045,N_11518);
and U14254 (N_14254,N_12034,N_10692);
xnor U14255 (N_14255,N_12089,N_10925);
nor U14256 (N_14256,N_10170,N_12330);
and U14257 (N_14257,N_10779,N_10687);
nor U14258 (N_14258,N_12298,N_11008);
xor U14259 (N_14259,N_10848,N_11190);
nand U14260 (N_14260,N_10864,N_11379);
or U14261 (N_14261,N_11775,N_11810);
or U14262 (N_14262,N_10183,N_10141);
xor U14263 (N_14263,N_10922,N_10426);
or U14264 (N_14264,N_11153,N_11929);
and U14265 (N_14265,N_11313,N_10244);
nand U14266 (N_14266,N_12256,N_10552);
nor U14267 (N_14267,N_11269,N_10593);
xnor U14268 (N_14268,N_10819,N_10535);
nand U14269 (N_14269,N_11353,N_10863);
nor U14270 (N_14270,N_10109,N_10982);
and U14271 (N_14271,N_12430,N_10150);
nor U14272 (N_14272,N_11491,N_11681);
and U14273 (N_14273,N_11284,N_10431);
nand U14274 (N_14274,N_11350,N_10460);
nand U14275 (N_14275,N_10845,N_12438);
nor U14276 (N_14276,N_10161,N_10000);
or U14277 (N_14277,N_11098,N_10853);
xor U14278 (N_14278,N_10575,N_12323);
and U14279 (N_14279,N_10355,N_10563);
xnor U14280 (N_14280,N_10898,N_12457);
nor U14281 (N_14281,N_10631,N_10829);
nand U14282 (N_14282,N_11409,N_11638);
nand U14283 (N_14283,N_11288,N_11860);
xor U14284 (N_14284,N_10177,N_11352);
xor U14285 (N_14285,N_10592,N_11994);
nor U14286 (N_14286,N_10603,N_12102);
xor U14287 (N_14287,N_10446,N_10736);
xor U14288 (N_14288,N_10635,N_10273);
nand U14289 (N_14289,N_12217,N_11398);
and U14290 (N_14290,N_11279,N_10495);
or U14291 (N_14291,N_11448,N_11604);
or U14292 (N_14292,N_10820,N_11628);
or U14293 (N_14293,N_11136,N_10992);
or U14294 (N_14294,N_11687,N_10955);
or U14295 (N_14295,N_10224,N_11405);
or U14296 (N_14296,N_11751,N_10306);
and U14297 (N_14297,N_10542,N_11389);
and U14298 (N_14298,N_11515,N_11808);
and U14299 (N_14299,N_10859,N_11337);
nand U14300 (N_14300,N_12015,N_12371);
or U14301 (N_14301,N_10971,N_11203);
nand U14302 (N_14302,N_10515,N_10038);
nand U14303 (N_14303,N_10666,N_10919);
nand U14304 (N_14304,N_11454,N_11653);
xnor U14305 (N_14305,N_10898,N_11969);
and U14306 (N_14306,N_12240,N_10867);
and U14307 (N_14307,N_10369,N_11928);
nand U14308 (N_14308,N_11650,N_11522);
and U14309 (N_14309,N_10678,N_10739);
nand U14310 (N_14310,N_11346,N_11299);
xor U14311 (N_14311,N_10656,N_10086);
xor U14312 (N_14312,N_10885,N_11684);
nor U14313 (N_14313,N_10994,N_11155);
nand U14314 (N_14314,N_12021,N_12334);
xnor U14315 (N_14315,N_10156,N_10605);
or U14316 (N_14316,N_11572,N_11769);
or U14317 (N_14317,N_10768,N_11965);
or U14318 (N_14318,N_11003,N_10450);
or U14319 (N_14319,N_11218,N_12490);
and U14320 (N_14320,N_11628,N_12060);
and U14321 (N_14321,N_10638,N_11646);
or U14322 (N_14322,N_12271,N_10111);
nor U14323 (N_14323,N_12153,N_12163);
xnor U14324 (N_14324,N_11273,N_11772);
nor U14325 (N_14325,N_12042,N_12417);
xor U14326 (N_14326,N_11561,N_12245);
or U14327 (N_14327,N_10864,N_12232);
nor U14328 (N_14328,N_12127,N_11785);
nor U14329 (N_14329,N_11903,N_11332);
xor U14330 (N_14330,N_12177,N_11304);
nand U14331 (N_14331,N_10860,N_10266);
nand U14332 (N_14332,N_10804,N_11630);
and U14333 (N_14333,N_11488,N_10149);
nand U14334 (N_14334,N_12143,N_11507);
nand U14335 (N_14335,N_10855,N_10874);
nand U14336 (N_14336,N_11903,N_10529);
nor U14337 (N_14337,N_10130,N_10860);
and U14338 (N_14338,N_12442,N_12263);
nand U14339 (N_14339,N_11003,N_10002);
or U14340 (N_14340,N_11961,N_11439);
nand U14341 (N_14341,N_11054,N_11964);
xor U14342 (N_14342,N_11854,N_10991);
nor U14343 (N_14343,N_10270,N_10123);
or U14344 (N_14344,N_10552,N_11119);
nor U14345 (N_14345,N_12153,N_11621);
or U14346 (N_14346,N_10221,N_11336);
or U14347 (N_14347,N_10911,N_12027);
nand U14348 (N_14348,N_10491,N_11348);
or U14349 (N_14349,N_12186,N_12300);
nand U14350 (N_14350,N_12102,N_10001);
and U14351 (N_14351,N_10901,N_11743);
and U14352 (N_14352,N_10436,N_11845);
xor U14353 (N_14353,N_10983,N_11283);
nor U14354 (N_14354,N_11345,N_11272);
and U14355 (N_14355,N_11634,N_10633);
or U14356 (N_14356,N_12144,N_10374);
nand U14357 (N_14357,N_11251,N_10262);
nand U14358 (N_14358,N_12482,N_10892);
or U14359 (N_14359,N_11001,N_10144);
and U14360 (N_14360,N_10111,N_10425);
nor U14361 (N_14361,N_10277,N_12163);
xor U14362 (N_14362,N_10487,N_11038);
nor U14363 (N_14363,N_11863,N_11357);
nor U14364 (N_14364,N_10751,N_10231);
nor U14365 (N_14365,N_10458,N_11099);
xor U14366 (N_14366,N_12104,N_12397);
nand U14367 (N_14367,N_12123,N_10316);
nor U14368 (N_14368,N_10020,N_11535);
xor U14369 (N_14369,N_12042,N_11657);
xnor U14370 (N_14370,N_11724,N_11795);
and U14371 (N_14371,N_12138,N_11073);
xnor U14372 (N_14372,N_10521,N_10358);
nor U14373 (N_14373,N_10692,N_11635);
nor U14374 (N_14374,N_10117,N_11077);
xor U14375 (N_14375,N_12471,N_11733);
and U14376 (N_14376,N_11655,N_11046);
and U14377 (N_14377,N_11345,N_11757);
xor U14378 (N_14378,N_10814,N_12225);
nand U14379 (N_14379,N_12206,N_11122);
xnor U14380 (N_14380,N_11203,N_11132);
or U14381 (N_14381,N_10835,N_12428);
and U14382 (N_14382,N_10377,N_10464);
and U14383 (N_14383,N_10013,N_11406);
xor U14384 (N_14384,N_12105,N_12486);
nor U14385 (N_14385,N_11977,N_10895);
and U14386 (N_14386,N_10306,N_11859);
nor U14387 (N_14387,N_11673,N_11667);
nor U14388 (N_14388,N_10852,N_10413);
or U14389 (N_14389,N_10453,N_11681);
nor U14390 (N_14390,N_11555,N_10410);
nand U14391 (N_14391,N_10580,N_10227);
xor U14392 (N_14392,N_12068,N_12001);
nand U14393 (N_14393,N_11417,N_12194);
and U14394 (N_14394,N_12116,N_12492);
xor U14395 (N_14395,N_10505,N_11063);
xor U14396 (N_14396,N_12109,N_10641);
nand U14397 (N_14397,N_11838,N_10530);
or U14398 (N_14398,N_11803,N_10844);
nand U14399 (N_14399,N_11321,N_12324);
or U14400 (N_14400,N_11526,N_10935);
and U14401 (N_14401,N_10808,N_11621);
nand U14402 (N_14402,N_10192,N_10360);
xor U14403 (N_14403,N_10133,N_10351);
nor U14404 (N_14404,N_10441,N_10786);
and U14405 (N_14405,N_12236,N_11502);
xor U14406 (N_14406,N_11812,N_11430);
nor U14407 (N_14407,N_10774,N_10371);
nor U14408 (N_14408,N_11789,N_11886);
or U14409 (N_14409,N_11295,N_11471);
nand U14410 (N_14410,N_10046,N_11736);
and U14411 (N_14411,N_10813,N_12471);
nand U14412 (N_14412,N_12131,N_10797);
xor U14413 (N_14413,N_11204,N_12213);
nand U14414 (N_14414,N_10831,N_10245);
nor U14415 (N_14415,N_12133,N_11949);
nor U14416 (N_14416,N_11256,N_10461);
nand U14417 (N_14417,N_10003,N_11834);
nor U14418 (N_14418,N_10932,N_10874);
xnor U14419 (N_14419,N_10782,N_10074);
or U14420 (N_14420,N_12159,N_11187);
nor U14421 (N_14421,N_10099,N_12413);
or U14422 (N_14422,N_11350,N_12466);
and U14423 (N_14423,N_10457,N_11710);
xor U14424 (N_14424,N_11482,N_11903);
nor U14425 (N_14425,N_11297,N_10489);
xnor U14426 (N_14426,N_11816,N_11710);
or U14427 (N_14427,N_10761,N_11722);
and U14428 (N_14428,N_10227,N_12378);
nor U14429 (N_14429,N_10200,N_11561);
and U14430 (N_14430,N_10757,N_11732);
or U14431 (N_14431,N_11012,N_10398);
xnor U14432 (N_14432,N_11026,N_11908);
nor U14433 (N_14433,N_11418,N_10714);
nand U14434 (N_14434,N_10212,N_12150);
or U14435 (N_14435,N_12215,N_10558);
nand U14436 (N_14436,N_10625,N_12022);
xnor U14437 (N_14437,N_11331,N_10234);
nand U14438 (N_14438,N_12308,N_10934);
nand U14439 (N_14439,N_11477,N_10097);
nand U14440 (N_14440,N_11761,N_11892);
or U14441 (N_14441,N_10437,N_12060);
or U14442 (N_14442,N_12036,N_10694);
nand U14443 (N_14443,N_12453,N_12270);
nor U14444 (N_14444,N_10298,N_10270);
and U14445 (N_14445,N_10717,N_10828);
nand U14446 (N_14446,N_12225,N_11141);
nand U14447 (N_14447,N_11775,N_10459);
nor U14448 (N_14448,N_11627,N_11864);
and U14449 (N_14449,N_12414,N_12465);
nor U14450 (N_14450,N_10898,N_10130);
and U14451 (N_14451,N_11543,N_11241);
nor U14452 (N_14452,N_12383,N_10803);
or U14453 (N_14453,N_11540,N_11459);
xnor U14454 (N_14454,N_11878,N_11464);
and U14455 (N_14455,N_11263,N_11209);
and U14456 (N_14456,N_11857,N_10481);
nand U14457 (N_14457,N_10946,N_10173);
nor U14458 (N_14458,N_11082,N_10527);
nand U14459 (N_14459,N_10207,N_10619);
nand U14460 (N_14460,N_10634,N_10648);
or U14461 (N_14461,N_11420,N_11999);
and U14462 (N_14462,N_12062,N_11950);
and U14463 (N_14463,N_10260,N_10637);
nand U14464 (N_14464,N_12225,N_10533);
nor U14465 (N_14465,N_11603,N_11059);
nand U14466 (N_14466,N_11227,N_11286);
nor U14467 (N_14467,N_10237,N_11810);
or U14468 (N_14468,N_11619,N_11060);
xor U14469 (N_14469,N_11582,N_10959);
nand U14470 (N_14470,N_11112,N_11991);
and U14471 (N_14471,N_11288,N_12014);
and U14472 (N_14472,N_11070,N_12191);
nand U14473 (N_14473,N_11818,N_11202);
nand U14474 (N_14474,N_11837,N_11682);
xor U14475 (N_14475,N_10903,N_12453);
and U14476 (N_14476,N_10971,N_12241);
or U14477 (N_14477,N_11494,N_10737);
or U14478 (N_14478,N_10343,N_11823);
or U14479 (N_14479,N_12217,N_11448);
or U14480 (N_14480,N_12012,N_10194);
xor U14481 (N_14481,N_12080,N_10372);
and U14482 (N_14482,N_10758,N_12346);
or U14483 (N_14483,N_11323,N_12173);
nand U14484 (N_14484,N_10542,N_12281);
nor U14485 (N_14485,N_12384,N_11202);
and U14486 (N_14486,N_10975,N_10020);
or U14487 (N_14487,N_11185,N_11170);
nor U14488 (N_14488,N_10027,N_11600);
and U14489 (N_14489,N_10155,N_11409);
nand U14490 (N_14490,N_10978,N_11821);
or U14491 (N_14491,N_12098,N_11691);
nor U14492 (N_14492,N_11086,N_11290);
nand U14493 (N_14493,N_10886,N_10975);
nor U14494 (N_14494,N_11630,N_11940);
nor U14495 (N_14495,N_10769,N_11214);
xnor U14496 (N_14496,N_10601,N_11664);
xnor U14497 (N_14497,N_12058,N_11950);
nand U14498 (N_14498,N_11436,N_10165);
xor U14499 (N_14499,N_10684,N_10179);
xor U14500 (N_14500,N_12326,N_10500);
and U14501 (N_14501,N_12424,N_12182);
xor U14502 (N_14502,N_11162,N_10752);
and U14503 (N_14503,N_11654,N_12363);
xnor U14504 (N_14504,N_12322,N_10683);
nor U14505 (N_14505,N_12085,N_10121);
nor U14506 (N_14506,N_11998,N_12048);
nand U14507 (N_14507,N_10574,N_11479);
nor U14508 (N_14508,N_11020,N_12348);
or U14509 (N_14509,N_10819,N_11781);
nor U14510 (N_14510,N_11005,N_10670);
nand U14511 (N_14511,N_11099,N_10187);
or U14512 (N_14512,N_10538,N_11444);
nand U14513 (N_14513,N_12041,N_10613);
and U14514 (N_14514,N_10779,N_12301);
nand U14515 (N_14515,N_11254,N_12060);
nand U14516 (N_14516,N_11301,N_11934);
or U14517 (N_14517,N_10469,N_11487);
and U14518 (N_14518,N_10903,N_11854);
or U14519 (N_14519,N_10862,N_11861);
nor U14520 (N_14520,N_10044,N_11807);
and U14521 (N_14521,N_11982,N_11229);
xor U14522 (N_14522,N_10084,N_10426);
nor U14523 (N_14523,N_10906,N_11034);
nand U14524 (N_14524,N_12022,N_10375);
nor U14525 (N_14525,N_11975,N_10989);
nor U14526 (N_14526,N_10672,N_11359);
or U14527 (N_14527,N_10570,N_12478);
nor U14528 (N_14528,N_11771,N_12402);
or U14529 (N_14529,N_10528,N_10339);
nand U14530 (N_14530,N_11795,N_10262);
and U14531 (N_14531,N_10354,N_10106);
and U14532 (N_14532,N_10137,N_11676);
xnor U14533 (N_14533,N_11973,N_11335);
or U14534 (N_14534,N_10643,N_12450);
and U14535 (N_14535,N_11084,N_11015);
and U14536 (N_14536,N_11713,N_11718);
and U14537 (N_14537,N_10276,N_11930);
xnor U14538 (N_14538,N_10733,N_11309);
and U14539 (N_14539,N_10037,N_11201);
and U14540 (N_14540,N_10404,N_11368);
and U14541 (N_14541,N_10486,N_10703);
nor U14542 (N_14542,N_10709,N_12387);
or U14543 (N_14543,N_10798,N_10736);
xor U14544 (N_14544,N_11533,N_11285);
or U14545 (N_14545,N_11363,N_10623);
xnor U14546 (N_14546,N_11792,N_10368);
nand U14547 (N_14547,N_10548,N_10709);
nand U14548 (N_14548,N_12180,N_10909);
nand U14549 (N_14549,N_11195,N_12458);
and U14550 (N_14550,N_12262,N_10846);
or U14551 (N_14551,N_10207,N_10988);
or U14552 (N_14552,N_11810,N_10656);
or U14553 (N_14553,N_10862,N_10632);
and U14554 (N_14554,N_10449,N_11772);
xnor U14555 (N_14555,N_12014,N_10862);
xnor U14556 (N_14556,N_10312,N_11250);
and U14557 (N_14557,N_12303,N_10172);
and U14558 (N_14558,N_10143,N_11845);
xor U14559 (N_14559,N_10046,N_11730);
nand U14560 (N_14560,N_10917,N_11873);
nand U14561 (N_14561,N_11224,N_12137);
xnor U14562 (N_14562,N_11395,N_11682);
nand U14563 (N_14563,N_12311,N_10975);
xor U14564 (N_14564,N_11748,N_10443);
xor U14565 (N_14565,N_12129,N_10781);
xor U14566 (N_14566,N_10731,N_10678);
nand U14567 (N_14567,N_11427,N_11524);
or U14568 (N_14568,N_10365,N_11704);
nor U14569 (N_14569,N_11411,N_11141);
xnor U14570 (N_14570,N_10832,N_12032);
nand U14571 (N_14571,N_10047,N_12196);
or U14572 (N_14572,N_11857,N_11642);
and U14573 (N_14573,N_11384,N_11788);
or U14574 (N_14574,N_12484,N_12080);
and U14575 (N_14575,N_10948,N_10646);
nand U14576 (N_14576,N_10972,N_10603);
and U14577 (N_14577,N_11199,N_11502);
nor U14578 (N_14578,N_10851,N_10493);
xnor U14579 (N_14579,N_11803,N_12451);
xnor U14580 (N_14580,N_10864,N_12331);
or U14581 (N_14581,N_12040,N_12490);
and U14582 (N_14582,N_10521,N_10284);
xnor U14583 (N_14583,N_11720,N_10209);
nand U14584 (N_14584,N_10559,N_12465);
xor U14585 (N_14585,N_11916,N_10146);
xnor U14586 (N_14586,N_11941,N_11038);
xnor U14587 (N_14587,N_11732,N_12144);
nand U14588 (N_14588,N_11699,N_12050);
xor U14589 (N_14589,N_11548,N_11232);
nor U14590 (N_14590,N_12428,N_12325);
nand U14591 (N_14591,N_11027,N_10167);
nor U14592 (N_14592,N_11472,N_10373);
xor U14593 (N_14593,N_12412,N_10967);
nor U14594 (N_14594,N_11329,N_11391);
nand U14595 (N_14595,N_11246,N_12051);
nand U14596 (N_14596,N_10813,N_10317);
nand U14597 (N_14597,N_11400,N_10123);
or U14598 (N_14598,N_12495,N_12393);
xnor U14599 (N_14599,N_10017,N_12342);
nor U14600 (N_14600,N_10482,N_11902);
xor U14601 (N_14601,N_12157,N_11803);
or U14602 (N_14602,N_11123,N_11812);
or U14603 (N_14603,N_10963,N_11547);
xor U14604 (N_14604,N_11734,N_11545);
or U14605 (N_14605,N_12016,N_12021);
and U14606 (N_14606,N_12121,N_12419);
and U14607 (N_14607,N_10199,N_12081);
xnor U14608 (N_14608,N_10826,N_11562);
and U14609 (N_14609,N_12013,N_10502);
nor U14610 (N_14610,N_11491,N_11288);
and U14611 (N_14611,N_10246,N_12236);
and U14612 (N_14612,N_11647,N_11851);
nor U14613 (N_14613,N_10329,N_12470);
nor U14614 (N_14614,N_12256,N_11724);
or U14615 (N_14615,N_10789,N_10008);
or U14616 (N_14616,N_11198,N_11570);
xor U14617 (N_14617,N_11650,N_11335);
or U14618 (N_14618,N_11729,N_11544);
or U14619 (N_14619,N_10816,N_11343);
nor U14620 (N_14620,N_10429,N_11785);
xor U14621 (N_14621,N_12496,N_10721);
xor U14622 (N_14622,N_11108,N_12450);
xnor U14623 (N_14623,N_11052,N_10282);
nor U14624 (N_14624,N_10192,N_12458);
nand U14625 (N_14625,N_11131,N_10417);
or U14626 (N_14626,N_10844,N_12322);
xor U14627 (N_14627,N_11471,N_10246);
and U14628 (N_14628,N_10935,N_11269);
xnor U14629 (N_14629,N_11659,N_11431);
or U14630 (N_14630,N_12288,N_11340);
and U14631 (N_14631,N_11473,N_12243);
or U14632 (N_14632,N_12477,N_10720);
nor U14633 (N_14633,N_11173,N_11099);
nand U14634 (N_14634,N_11437,N_10558);
or U14635 (N_14635,N_11918,N_10332);
nand U14636 (N_14636,N_11727,N_11421);
xnor U14637 (N_14637,N_10812,N_10481);
or U14638 (N_14638,N_11032,N_11509);
and U14639 (N_14639,N_11287,N_11751);
and U14640 (N_14640,N_10393,N_11958);
nand U14641 (N_14641,N_11266,N_12251);
and U14642 (N_14642,N_10948,N_10339);
xnor U14643 (N_14643,N_10875,N_10296);
nor U14644 (N_14644,N_11443,N_10124);
or U14645 (N_14645,N_11893,N_11302);
and U14646 (N_14646,N_10956,N_11991);
nand U14647 (N_14647,N_11189,N_11469);
nor U14648 (N_14648,N_12250,N_11543);
and U14649 (N_14649,N_11659,N_11364);
xnor U14650 (N_14650,N_11658,N_12111);
or U14651 (N_14651,N_10372,N_11855);
or U14652 (N_14652,N_10368,N_10039);
xnor U14653 (N_14653,N_10265,N_11023);
and U14654 (N_14654,N_11472,N_12301);
and U14655 (N_14655,N_12398,N_10721);
xnor U14656 (N_14656,N_10591,N_11385);
and U14657 (N_14657,N_12445,N_12452);
or U14658 (N_14658,N_11258,N_12367);
xnor U14659 (N_14659,N_11443,N_11986);
nor U14660 (N_14660,N_11381,N_11967);
nor U14661 (N_14661,N_10609,N_11344);
nand U14662 (N_14662,N_11500,N_10182);
or U14663 (N_14663,N_11997,N_11161);
nor U14664 (N_14664,N_11947,N_10208);
or U14665 (N_14665,N_10588,N_10222);
nand U14666 (N_14666,N_12449,N_12037);
and U14667 (N_14667,N_10815,N_11719);
nand U14668 (N_14668,N_11486,N_11151);
nor U14669 (N_14669,N_10431,N_12406);
nor U14670 (N_14670,N_10251,N_10777);
or U14671 (N_14671,N_10257,N_12494);
nand U14672 (N_14672,N_11631,N_11417);
or U14673 (N_14673,N_12270,N_12121);
or U14674 (N_14674,N_12414,N_10310);
nand U14675 (N_14675,N_12208,N_11871);
and U14676 (N_14676,N_11644,N_11101);
nand U14677 (N_14677,N_10405,N_12001);
nand U14678 (N_14678,N_10823,N_11389);
or U14679 (N_14679,N_11474,N_12296);
and U14680 (N_14680,N_10288,N_11394);
xnor U14681 (N_14681,N_11442,N_10191);
and U14682 (N_14682,N_10312,N_10041);
or U14683 (N_14683,N_11865,N_10414);
or U14684 (N_14684,N_10890,N_11274);
and U14685 (N_14685,N_10230,N_11389);
xor U14686 (N_14686,N_11291,N_10783);
xor U14687 (N_14687,N_12100,N_10194);
nand U14688 (N_14688,N_10900,N_11220);
and U14689 (N_14689,N_10274,N_10212);
xnor U14690 (N_14690,N_10742,N_11920);
nor U14691 (N_14691,N_11529,N_12494);
nand U14692 (N_14692,N_10415,N_10203);
xor U14693 (N_14693,N_11777,N_10933);
nand U14694 (N_14694,N_10288,N_10665);
or U14695 (N_14695,N_11031,N_10792);
or U14696 (N_14696,N_12335,N_12007);
xnor U14697 (N_14697,N_10603,N_10635);
nor U14698 (N_14698,N_11760,N_10081);
nand U14699 (N_14699,N_10645,N_12037);
and U14700 (N_14700,N_11019,N_11044);
xnor U14701 (N_14701,N_10500,N_12071);
nor U14702 (N_14702,N_12113,N_10413);
and U14703 (N_14703,N_11122,N_12437);
nor U14704 (N_14704,N_12435,N_11918);
nor U14705 (N_14705,N_12109,N_10154);
and U14706 (N_14706,N_11487,N_12432);
xor U14707 (N_14707,N_11376,N_10025);
or U14708 (N_14708,N_10193,N_10246);
and U14709 (N_14709,N_12257,N_10280);
or U14710 (N_14710,N_10621,N_12467);
or U14711 (N_14711,N_11861,N_12048);
or U14712 (N_14712,N_10389,N_10872);
or U14713 (N_14713,N_11625,N_12306);
xnor U14714 (N_14714,N_11848,N_10303);
and U14715 (N_14715,N_10155,N_11456);
nand U14716 (N_14716,N_10010,N_10761);
nor U14717 (N_14717,N_12054,N_11038);
xnor U14718 (N_14718,N_10027,N_10504);
nand U14719 (N_14719,N_12203,N_11667);
nand U14720 (N_14720,N_12258,N_10479);
nor U14721 (N_14721,N_10074,N_10834);
nand U14722 (N_14722,N_12039,N_11594);
xor U14723 (N_14723,N_12267,N_10235);
nor U14724 (N_14724,N_12250,N_10876);
or U14725 (N_14725,N_10076,N_11634);
nor U14726 (N_14726,N_10319,N_11270);
or U14727 (N_14727,N_11323,N_10029);
nor U14728 (N_14728,N_10247,N_11840);
or U14729 (N_14729,N_12429,N_11408);
nor U14730 (N_14730,N_10156,N_11191);
and U14731 (N_14731,N_11554,N_11012);
nor U14732 (N_14732,N_10357,N_12301);
nor U14733 (N_14733,N_12493,N_12272);
nand U14734 (N_14734,N_10082,N_12487);
and U14735 (N_14735,N_11044,N_10089);
xor U14736 (N_14736,N_12165,N_11738);
nand U14737 (N_14737,N_11659,N_10199);
or U14738 (N_14738,N_10454,N_11369);
and U14739 (N_14739,N_11062,N_11235);
xor U14740 (N_14740,N_10958,N_11077);
nand U14741 (N_14741,N_10175,N_11909);
or U14742 (N_14742,N_12033,N_12046);
nand U14743 (N_14743,N_11930,N_10229);
nand U14744 (N_14744,N_11925,N_10451);
or U14745 (N_14745,N_11235,N_12149);
and U14746 (N_14746,N_10063,N_10666);
or U14747 (N_14747,N_11578,N_11749);
and U14748 (N_14748,N_11670,N_12369);
nor U14749 (N_14749,N_11135,N_11594);
nor U14750 (N_14750,N_12252,N_11433);
xnor U14751 (N_14751,N_11227,N_12467);
and U14752 (N_14752,N_11687,N_10623);
nand U14753 (N_14753,N_11306,N_10263);
nand U14754 (N_14754,N_12484,N_10384);
and U14755 (N_14755,N_10512,N_10277);
xnor U14756 (N_14756,N_11602,N_10220);
or U14757 (N_14757,N_12091,N_11457);
or U14758 (N_14758,N_12366,N_10469);
or U14759 (N_14759,N_10576,N_10354);
xnor U14760 (N_14760,N_11102,N_11932);
xor U14761 (N_14761,N_11370,N_12043);
and U14762 (N_14762,N_10188,N_11063);
xnor U14763 (N_14763,N_11490,N_10698);
xor U14764 (N_14764,N_12155,N_10031);
or U14765 (N_14765,N_10542,N_12025);
and U14766 (N_14766,N_11432,N_10705);
or U14767 (N_14767,N_11419,N_10091);
and U14768 (N_14768,N_12258,N_10849);
xor U14769 (N_14769,N_10554,N_10608);
or U14770 (N_14770,N_10114,N_12322);
nor U14771 (N_14771,N_10935,N_10710);
nor U14772 (N_14772,N_11927,N_10161);
xnor U14773 (N_14773,N_11790,N_11291);
nor U14774 (N_14774,N_11288,N_10008);
xor U14775 (N_14775,N_12462,N_11321);
xor U14776 (N_14776,N_12303,N_11453);
and U14777 (N_14777,N_11377,N_11330);
nor U14778 (N_14778,N_10600,N_11684);
nand U14779 (N_14779,N_12376,N_10970);
and U14780 (N_14780,N_11022,N_12123);
and U14781 (N_14781,N_10633,N_10003);
or U14782 (N_14782,N_10839,N_11275);
or U14783 (N_14783,N_12438,N_12221);
nor U14784 (N_14784,N_10501,N_11978);
and U14785 (N_14785,N_10513,N_12421);
nor U14786 (N_14786,N_11374,N_10979);
nand U14787 (N_14787,N_12246,N_10382);
nor U14788 (N_14788,N_10916,N_11515);
nand U14789 (N_14789,N_10186,N_11075);
or U14790 (N_14790,N_12350,N_10407);
or U14791 (N_14791,N_10951,N_11553);
xor U14792 (N_14792,N_10057,N_12079);
nor U14793 (N_14793,N_12440,N_10717);
nor U14794 (N_14794,N_12153,N_10410);
nand U14795 (N_14795,N_10150,N_10987);
nor U14796 (N_14796,N_10394,N_11035);
or U14797 (N_14797,N_11673,N_11194);
nand U14798 (N_14798,N_10092,N_12311);
xnor U14799 (N_14799,N_11100,N_11231);
and U14800 (N_14800,N_11717,N_10318);
nor U14801 (N_14801,N_10106,N_11375);
nand U14802 (N_14802,N_11579,N_11553);
and U14803 (N_14803,N_11468,N_11690);
nand U14804 (N_14804,N_11541,N_10177);
nor U14805 (N_14805,N_10417,N_10530);
or U14806 (N_14806,N_12463,N_11029);
nor U14807 (N_14807,N_11116,N_10392);
nor U14808 (N_14808,N_10187,N_12133);
nor U14809 (N_14809,N_10922,N_11287);
nand U14810 (N_14810,N_11374,N_11876);
nor U14811 (N_14811,N_12272,N_12028);
and U14812 (N_14812,N_11199,N_12277);
nand U14813 (N_14813,N_10761,N_11959);
or U14814 (N_14814,N_10599,N_10624);
or U14815 (N_14815,N_11185,N_10808);
nand U14816 (N_14816,N_12439,N_12158);
and U14817 (N_14817,N_10814,N_11674);
nand U14818 (N_14818,N_11206,N_11218);
xor U14819 (N_14819,N_11814,N_11113);
nor U14820 (N_14820,N_11924,N_11857);
xnor U14821 (N_14821,N_10088,N_11645);
or U14822 (N_14822,N_10640,N_11363);
or U14823 (N_14823,N_11861,N_10481);
xnor U14824 (N_14824,N_12375,N_10369);
xor U14825 (N_14825,N_11197,N_11640);
xor U14826 (N_14826,N_12279,N_12068);
and U14827 (N_14827,N_11929,N_10064);
nor U14828 (N_14828,N_10595,N_12051);
xnor U14829 (N_14829,N_12208,N_10245);
and U14830 (N_14830,N_10283,N_10754);
xnor U14831 (N_14831,N_10169,N_10621);
xor U14832 (N_14832,N_11767,N_11420);
nand U14833 (N_14833,N_10903,N_11148);
nand U14834 (N_14834,N_12017,N_12376);
nand U14835 (N_14835,N_11723,N_11200);
nor U14836 (N_14836,N_10435,N_11791);
nor U14837 (N_14837,N_11712,N_12147);
and U14838 (N_14838,N_11799,N_11079);
nor U14839 (N_14839,N_11446,N_10393);
nand U14840 (N_14840,N_10319,N_11854);
nor U14841 (N_14841,N_12347,N_11274);
and U14842 (N_14842,N_10052,N_11566);
or U14843 (N_14843,N_11254,N_10467);
nand U14844 (N_14844,N_10470,N_10308);
nor U14845 (N_14845,N_11420,N_11938);
xnor U14846 (N_14846,N_11976,N_10263);
nor U14847 (N_14847,N_10706,N_11809);
nand U14848 (N_14848,N_10550,N_10637);
or U14849 (N_14849,N_11803,N_11708);
nor U14850 (N_14850,N_12384,N_10750);
or U14851 (N_14851,N_11913,N_10598);
and U14852 (N_14852,N_10921,N_10953);
nor U14853 (N_14853,N_10697,N_10310);
xor U14854 (N_14854,N_11299,N_10548);
and U14855 (N_14855,N_10205,N_10191);
xor U14856 (N_14856,N_11509,N_11941);
nand U14857 (N_14857,N_11775,N_11210);
xor U14858 (N_14858,N_10307,N_11876);
nor U14859 (N_14859,N_11177,N_11094);
and U14860 (N_14860,N_10822,N_10498);
nor U14861 (N_14861,N_11727,N_10589);
nor U14862 (N_14862,N_10162,N_10114);
nand U14863 (N_14863,N_10732,N_10858);
nand U14864 (N_14864,N_10042,N_11645);
nand U14865 (N_14865,N_12160,N_11226);
nor U14866 (N_14866,N_10421,N_11405);
xnor U14867 (N_14867,N_10920,N_12191);
nor U14868 (N_14868,N_11481,N_11491);
or U14869 (N_14869,N_10188,N_11838);
nand U14870 (N_14870,N_11424,N_11909);
nand U14871 (N_14871,N_12487,N_12155);
or U14872 (N_14872,N_10722,N_11961);
and U14873 (N_14873,N_10370,N_10289);
xor U14874 (N_14874,N_12089,N_11835);
or U14875 (N_14875,N_10748,N_12397);
and U14876 (N_14876,N_10597,N_11879);
nand U14877 (N_14877,N_11316,N_10813);
nor U14878 (N_14878,N_12030,N_10695);
nand U14879 (N_14879,N_11021,N_10812);
and U14880 (N_14880,N_10082,N_11517);
or U14881 (N_14881,N_12071,N_10455);
or U14882 (N_14882,N_12016,N_11925);
or U14883 (N_14883,N_10280,N_10563);
xor U14884 (N_14884,N_11257,N_12269);
and U14885 (N_14885,N_11018,N_11691);
xor U14886 (N_14886,N_10339,N_12312);
xnor U14887 (N_14887,N_10311,N_11268);
nand U14888 (N_14888,N_10551,N_11064);
or U14889 (N_14889,N_10628,N_10513);
or U14890 (N_14890,N_12058,N_10043);
xnor U14891 (N_14891,N_12302,N_12101);
xor U14892 (N_14892,N_11277,N_11976);
nand U14893 (N_14893,N_11821,N_11864);
xor U14894 (N_14894,N_11772,N_10120);
and U14895 (N_14895,N_11966,N_11056);
or U14896 (N_14896,N_11825,N_11427);
xor U14897 (N_14897,N_10219,N_12317);
nand U14898 (N_14898,N_10634,N_10254);
or U14899 (N_14899,N_11616,N_11658);
and U14900 (N_14900,N_10936,N_11646);
nand U14901 (N_14901,N_10853,N_11724);
nand U14902 (N_14902,N_11328,N_10989);
nand U14903 (N_14903,N_11993,N_12033);
and U14904 (N_14904,N_11405,N_11742);
nor U14905 (N_14905,N_12080,N_10506);
and U14906 (N_14906,N_11070,N_11418);
and U14907 (N_14907,N_12378,N_11146);
nor U14908 (N_14908,N_10173,N_10054);
nor U14909 (N_14909,N_11590,N_12496);
xor U14910 (N_14910,N_11854,N_10561);
nand U14911 (N_14911,N_12357,N_12000);
nor U14912 (N_14912,N_12176,N_12347);
nand U14913 (N_14913,N_11341,N_11619);
nand U14914 (N_14914,N_11963,N_11966);
and U14915 (N_14915,N_11945,N_11517);
or U14916 (N_14916,N_10985,N_11703);
or U14917 (N_14917,N_11578,N_11025);
nand U14918 (N_14918,N_10583,N_12172);
nor U14919 (N_14919,N_12389,N_12128);
and U14920 (N_14920,N_12496,N_12202);
or U14921 (N_14921,N_11423,N_10401);
nor U14922 (N_14922,N_11118,N_10675);
nor U14923 (N_14923,N_10243,N_11963);
and U14924 (N_14924,N_11484,N_10538);
nand U14925 (N_14925,N_11146,N_11610);
or U14926 (N_14926,N_10545,N_12470);
or U14927 (N_14927,N_10379,N_12453);
or U14928 (N_14928,N_10611,N_12182);
nand U14929 (N_14929,N_12070,N_11643);
xor U14930 (N_14930,N_11746,N_12035);
nand U14931 (N_14931,N_11857,N_10494);
xor U14932 (N_14932,N_12332,N_10198);
nor U14933 (N_14933,N_10728,N_12251);
nand U14934 (N_14934,N_12164,N_10558);
xnor U14935 (N_14935,N_12419,N_12249);
nand U14936 (N_14936,N_10559,N_10169);
and U14937 (N_14937,N_11448,N_10426);
nor U14938 (N_14938,N_11285,N_10113);
xnor U14939 (N_14939,N_10014,N_11299);
xor U14940 (N_14940,N_11821,N_12415);
or U14941 (N_14941,N_12215,N_10916);
nand U14942 (N_14942,N_11682,N_11899);
xor U14943 (N_14943,N_10022,N_11663);
xor U14944 (N_14944,N_12033,N_12018);
nor U14945 (N_14945,N_10417,N_11277);
xor U14946 (N_14946,N_10452,N_10493);
nor U14947 (N_14947,N_10140,N_11047);
and U14948 (N_14948,N_11189,N_10876);
nand U14949 (N_14949,N_10144,N_12372);
xnor U14950 (N_14950,N_10609,N_10814);
and U14951 (N_14951,N_11487,N_11019);
and U14952 (N_14952,N_12226,N_11116);
nor U14953 (N_14953,N_11061,N_10017);
or U14954 (N_14954,N_11477,N_10269);
or U14955 (N_14955,N_11207,N_12471);
nand U14956 (N_14956,N_10154,N_12294);
nand U14957 (N_14957,N_11068,N_10993);
or U14958 (N_14958,N_11752,N_11946);
xnor U14959 (N_14959,N_11883,N_11205);
or U14960 (N_14960,N_11802,N_11734);
or U14961 (N_14961,N_11200,N_10007);
or U14962 (N_14962,N_11756,N_11912);
and U14963 (N_14963,N_11989,N_10597);
xor U14964 (N_14964,N_11214,N_10610);
nand U14965 (N_14965,N_10959,N_12384);
nand U14966 (N_14966,N_12457,N_11641);
xnor U14967 (N_14967,N_11966,N_10578);
nand U14968 (N_14968,N_10679,N_10878);
xor U14969 (N_14969,N_11806,N_10975);
or U14970 (N_14970,N_12213,N_11532);
nand U14971 (N_14971,N_10072,N_10596);
nand U14972 (N_14972,N_11707,N_10869);
and U14973 (N_14973,N_11926,N_11427);
and U14974 (N_14974,N_11732,N_11001);
or U14975 (N_14975,N_11278,N_11048);
and U14976 (N_14976,N_12262,N_12417);
xor U14977 (N_14977,N_11330,N_10098);
nor U14978 (N_14978,N_11518,N_11146);
nand U14979 (N_14979,N_12109,N_10365);
or U14980 (N_14980,N_11181,N_11675);
nand U14981 (N_14981,N_12020,N_12363);
nor U14982 (N_14982,N_11781,N_10384);
nor U14983 (N_14983,N_12047,N_10786);
nand U14984 (N_14984,N_11363,N_10891);
or U14985 (N_14985,N_10701,N_11730);
xnor U14986 (N_14986,N_12065,N_10184);
and U14987 (N_14987,N_12157,N_11517);
nor U14988 (N_14988,N_10326,N_11991);
and U14989 (N_14989,N_10343,N_11280);
nor U14990 (N_14990,N_10222,N_11546);
or U14991 (N_14991,N_10900,N_11773);
nor U14992 (N_14992,N_10841,N_11897);
nor U14993 (N_14993,N_11750,N_12092);
or U14994 (N_14994,N_10534,N_11705);
xnor U14995 (N_14995,N_10828,N_12363);
xor U14996 (N_14996,N_10314,N_10520);
nand U14997 (N_14997,N_10418,N_10801);
xor U14998 (N_14998,N_12328,N_11612);
xnor U14999 (N_14999,N_10881,N_11225);
or U15000 (N_15000,N_13016,N_13308);
nor U15001 (N_15001,N_14555,N_12826);
nor U15002 (N_15002,N_14452,N_13196);
nand U15003 (N_15003,N_12715,N_14250);
xnor U15004 (N_15004,N_14462,N_14771);
nand U15005 (N_15005,N_12643,N_13784);
nor U15006 (N_15006,N_12530,N_12984);
nand U15007 (N_15007,N_13568,N_14357);
nand U15008 (N_15008,N_13488,N_13075);
xnor U15009 (N_15009,N_14308,N_13053);
or U15010 (N_15010,N_14664,N_13124);
nor U15011 (N_15011,N_14483,N_13634);
and U15012 (N_15012,N_14439,N_14090);
nand U15013 (N_15013,N_12939,N_12982);
nand U15014 (N_15014,N_13723,N_12674);
nand U15015 (N_15015,N_13062,N_13870);
and U15016 (N_15016,N_13325,N_14054);
nor U15017 (N_15017,N_13306,N_12535);
xnor U15018 (N_15018,N_12523,N_13435);
or U15019 (N_15019,N_12808,N_14823);
nand U15020 (N_15020,N_13892,N_14454);
nand U15021 (N_15021,N_14861,N_13839);
or U15022 (N_15022,N_14020,N_13057);
and U15023 (N_15023,N_13254,N_14038);
or U15024 (N_15024,N_13300,N_13363);
nand U15025 (N_15025,N_14348,N_13327);
nand U15026 (N_15026,N_12917,N_12508);
or U15027 (N_15027,N_13763,N_14925);
and U15028 (N_15028,N_13921,N_12698);
and U15029 (N_15029,N_14947,N_14616);
or U15030 (N_15030,N_13394,N_14293);
nand U15031 (N_15031,N_13460,N_13206);
xnor U15032 (N_15032,N_13333,N_13790);
and U15033 (N_15033,N_13910,N_14184);
nand U15034 (N_15034,N_13466,N_14652);
and U15035 (N_15035,N_13964,N_14882);
xor U15036 (N_15036,N_12832,N_13923);
nor U15037 (N_15037,N_13750,N_13098);
and U15038 (N_15038,N_12851,N_14165);
xor U15039 (N_15039,N_14353,N_13848);
or U15040 (N_15040,N_14239,N_14690);
and U15041 (N_15041,N_13485,N_14696);
or U15042 (N_15042,N_12944,N_13503);
nor U15043 (N_15043,N_12782,N_14494);
nand U15044 (N_15044,N_14758,N_12668);
nand U15045 (N_15045,N_13258,N_13480);
xor U15046 (N_15046,N_13153,N_13822);
xnor U15047 (N_15047,N_13904,N_14106);
nand U15048 (N_15048,N_14301,N_13428);
nor U15049 (N_15049,N_13102,N_13849);
or U15050 (N_15050,N_14116,N_13146);
xnor U15051 (N_15051,N_14952,N_14496);
or U15052 (N_15052,N_14962,N_13886);
or U15053 (N_15053,N_13513,N_13352);
nand U15054 (N_15054,N_12701,N_12956);
xnor U15055 (N_15055,N_12614,N_14344);
nor U15056 (N_15056,N_13190,N_14892);
and U15057 (N_15057,N_14501,N_12713);
and U15058 (N_15058,N_13317,N_13626);
xnor U15059 (N_15059,N_13105,N_13445);
or U15060 (N_15060,N_14248,N_13699);
xor U15061 (N_15061,N_12626,N_13698);
nor U15062 (N_15062,N_14334,N_13693);
or U15063 (N_15063,N_14727,N_13748);
xor U15064 (N_15064,N_13156,N_13932);
and U15065 (N_15065,N_14506,N_14644);
nand U15066 (N_15066,N_13252,N_13358);
nand U15067 (N_15067,N_14586,N_14889);
or U15068 (N_15068,N_12800,N_13453);
nand U15069 (N_15069,N_14241,N_13611);
nor U15070 (N_15070,N_13228,N_13584);
and U15071 (N_15071,N_13419,N_12551);
nand U15072 (N_15072,N_12850,N_13040);
xor U15073 (N_15073,N_14631,N_12986);
and U15074 (N_15074,N_14738,N_13391);
nor U15075 (N_15075,N_13337,N_12803);
and U15076 (N_15076,N_14992,N_13167);
nor U15077 (N_15077,N_13007,N_14317);
or U15078 (N_15078,N_13783,N_13773);
xnor U15079 (N_15079,N_14863,N_13341);
or U15080 (N_15080,N_13999,N_13437);
xor U15081 (N_15081,N_13881,N_13967);
nand U15082 (N_15082,N_14589,N_13244);
xor U15083 (N_15083,N_13052,N_12930);
or U15084 (N_15084,N_14729,N_13395);
nand U15085 (N_15085,N_14431,N_14540);
and U15086 (N_15086,N_14814,N_14078);
and U15087 (N_15087,N_13301,N_14599);
nor U15088 (N_15088,N_13820,N_12899);
nand U15089 (N_15089,N_13665,N_14595);
or U15090 (N_15090,N_14796,N_13262);
nand U15091 (N_15091,N_14660,N_12766);
or U15092 (N_15092,N_14836,N_13446);
nand U15093 (N_15093,N_14529,N_13674);
nor U15094 (N_15094,N_14959,N_13774);
or U15095 (N_15095,N_13170,N_12750);
and U15096 (N_15096,N_13613,N_14743);
nand U15097 (N_15097,N_13782,N_14413);
nand U15098 (N_15098,N_13478,N_14989);
nand U15099 (N_15099,N_13652,N_14950);
nand U15100 (N_15100,N_12838,N_14022);
xor U15101 (N_15101,N_13424,N_14192);
or U15102 (N_15102,N_13943,N_14811);
or U15103 (N_15103,N_14695,N_14759);
nor U15104 (N_15104,N_13928,N_12743);
and U15105 (N_15105,N_13083,N_13987);
or U15106 (N_15106,N_13577,N_12682);
xnor U15107 (N_15107,N_12860,N_13314);
nand U15108 (N_15108,N_12973,N_14709);
or U15109 (N_15109,N_14786,N_13548);
or U15110 (N_15110,N_13771,N_13149);
xor U15111 (N_15111,N_12672,N_14866);
xnor U15112 (N_15112,N_12932,N_13058);
nor U15113 (N_15113,N_14582,N_14522);
xnor U15114 (N_15114,N_12964,N_13609);
or U15115 (N_15115,N_14670,N_14173);
and U15116 (N_15116,N_14922,N_14915);
nand U15117 (N_15117,N_14155,N_12854);
or U15118 (N_15118,N_14570,N_13209);
or U15119 (N_15119,N_12656,N_14156);
nand U15120 (N_15120,N_13302,N_12799);
nand U15121 (N_15121,N_14645,N_13544);
nand U15122 (N_15122,N_14363,N_13799);
or U15123 (N_15123,N_14810,N_12874);
and U15124 (N_15124,N_12895,N_12764);
or U15125 (N_15125,N_14006,N_14651);
nand U15126 (N_15126,N_14369,N_14126);
or U15127 (N_15127,N_13659,N_14457);
or U15128 (N_15128,N_12796,N_14879);
xor U15129 (N_15129,N_12681,N_13742);
xor U15130 (N_15130,N_14531,N_14321);
or U15131 (N_15131,N_13617,N_13565);
xor U15132 (N_15132,N_14665,N_14404);
and U15133 (N_15133,N_12848,N_14532);
xor U15134 (N_15134,N_12654,N_12852);
or U15135 (N_15135,N_14217,N_14027);
nand U15136 (N_15136,N_14557,N_13861);
xnor U15137 (N_15137,N_14444,N_13767);
or U15138 (N_15138,N_14869,N_13347);
nor U15139 (N_15139,N_12640,N_14639);
xor U15140 (N_15140,N_14753,N_14568);
nand U15141 (N_15141,N_14517,N_14115);
or U15142 (N_15142,N_13487,N_14658);
nor U15143 (N_15143,N_13408,N_14957);
and U15144 (N_15144,N_13991,N_12566);
nand U15145 (N_15145,N_14847,N_13778);
xor U15146 (N_15146,N_14953,N_14898);
nor U15147 (N_15147,N_13425,N_12507);
or U15148 (N_15148,N_13013,N_14492);
and U15149 (N_15149,N_14990,N_14030);
nor U15150 (N_15150,N_14841,N_13184);
nor U15151 (N_15151,N_14234,N_14040);
xnor U15152 (N_15152,N_14306,N_13801);
or U15153 (N_15153,N_12897,N_13458);
and U15154 (N_15154,N_14421,N_12509);
and U15155 (N_15155,N_13482,N_14168);
nor U15156 (N_15156,N_13322,N_13712);
nor U15157 (N_15157,N_12876,N_14045);
nand U15158 (N_15158,N_12671,N_13403);
nor U15159 (N_15159,N_13789,N_12663);
nand U15160 (N_15160,N_13139,N_14839);
and U15161 (N_15161,N_14222,N_12928);
nor U15162 (N_15162,N_12568,N_13281);
nor U15163 (N_15163,N_12555,N_12631);
or U15164 (N_15164,N_14605,N_13941);
xnor U15165 (N_15165,N_13265,N_14859);
or U15166 (N_15166,N_13351,N_12721);
nor U15167 (N_15167,N_14577,N_13433);
xor U15168 (N_15168,N_13837,N_14319);
nand U15169 (N_15169,N_13655,N_12922);
or U15170 (N_15170,N_13705,N_14946);
and U15171 (N_15171,N_14337,N_13387);
and U15172 (N_15172,N_13441,N_12923);
nand U15173 (N_15173,N_14851,N_12697);
or U15174 (N_15174,N_14713,N_12572);
xor U15175 (N_15175,N_14060,N_13236);
nor U15176 (N_15176,N_12584,N_14827);
nand U15177 (N_15177,N_14587,N_13727);
or U15178 (N_15178,N_14097,N_13498);
or U15179 (N_15179,N_13444,N_14507);
xnor U15180 (N_15180,N_12898,N_13025);
and U15181 (N_15181,N_13818,N_14114);
xor U15182 (N_15182,N_14987,N_12521);
xnor U15183 (N_15183,N_13541,N_14411);
and U15184 (N_15184,N_14292,N_13050);
nand U15185 (N_15185,N_12995,N_14888);
and U15186 (N_15186,N_14967,N_12905);
nand U15187 (N_15187,N_13077,N_13169);
nand U15188 (N_15188,N_12841,N_12567);
nand U15189 (N_15189,N_12807,N_14926);
xor U15190 (N_15190,N_14893,N_13519);
xnor U15191 (N_15191,N_13587,N_13555);
or U15192 (N_15192,N_13942,N_13234);
and U15193 (N_15193,N_14955,N_13936);
or U15194 (N_15194,N_13724,N_13869);
nor U15195 (N_15195,N_12615,N_13827);
or U15196 (N_15196,N_14381,N_14681);
and U15197 (N_15197,N_14277,N_13131);
nand U15198 (N_15198,N_14976,N_14464);
or U15199 (N_15199,N_14152,N_12763);
nand U15200 (N_15200,N_14780,N_13618);
or U15201 (N_15201,N_13760,N_13147);
xnor U15202 (N_15202,N_13866,N_12975);
nor U15203 (N_15203,N_14091,N_13142);
or U15204 (N_15204,N_14552,N_14453);
or U15205 (N_15205,N_13957,N_13495);
nand U15206 (N_15206,N_12795,N_13035);
xnor U15207 (N_15207,N_12954,N_13830);
and U15208 (N_15208,N_14933,N_13512);
nor U15209 (N_15209,N_13218,N_13751);
and U15210 (N_15210,N_13261,N_14218);
nand U15211 (N_15211,N_14736,N_13323);
and U15212 (N_15212,N_13321,N_13372);
xnor U15213 (N_15213,N_13385,N_12506);
and U15214 (N_15214,N_12546,N_13030);
nor U15215 (N_15215,N_12692,N_13183);
and U15216 (N_15216,N_13907,N_12934);
nand U15217 (N_15217,N_12694,N_12936);
and U15218 (N_15218,N_13112,N_12933);
xor U15219 (N_15219,N_14145,N_14612);
or U15220 (N_15220,N_14716,N_14829);
nand U15221 (N_15221,N_14133,N_13654);
xnor U15222 (N_15222,N_14161,N_13217);
and U15223 (N_15223,N_13477,N_13536);
xor U15224 (N_15224,N_14674,N_14186);
xnor U15225 (N_15225,N_13974,N_13993);
xor U15226 (N_15226,N_14554,N_14895);
and U15227 (N_15227,N_13235,N_14305);
nor U15228 (N_15228,N_13481,N_13803);
xnor U15229 (N_15229,N_14415,N_13733);
nor U15230 (N_15230,N_14262,N_14638);
or U15231 (N_15231,N_14806,N_14164);
xnor U15232 (N_15232,N_13073,N_13992);
or U15233 (N_15233,N_13243,N_13821);
nand U15234 (N_15234,N_14273,N_14376);
or U15235 (N_15235,N_12557,N_13679);
and U15236 (N_15236,N_12779,N_14767);
or U15237 (N_15237,N_14868,N_14580);
or U15238 (N_15238,N_13645,N_13895);
and U15239 (N_15239,N_14949,N_13687);
nand U15240 (N_15240,N_13707,N_13451);
and U15241 (N_15241,N_14936,N_13880);
nor U15242 (N_15242,N_14757,N_12574);
xnor U15243 (N_15243,N_12849,N_14258);
xor U15244 (N_15244,N_13396,N_14979);
xor U15245 (N_15245,N_13474,N_13336);
nor U15246 (N_15246,N_14977,N_14052);
and U15247 (N_15247,N_12617,N_14023);
or U15248 (N_15248,N_14768,N_13549);
nor U15249 (N_15249,N_14528,N_13177);
nand U15250 (N_15250,N_14158,N_14538);
and U15251 (N_15251,N_13873,N_14190);
nor U15252 (N_15252,N_14443,N_14562);
nand U15253 (N_15253,N_13179,N_14880);
and U15254 (N_15254,N_13292,N_14831);
nor U15255 (N_15255,N_12739,N_13684);
xnor U15256 (N_15256,N_12998,N_14590);
and U15257 (N_15257,N_14844,N_14551);
nor U15258 (N_15258,N_13889,N_14733);
xnor U15259 (N_15259,N_13214,N_14336);
nor U15260 (N_15260,N_14072,N_14378);
xnor U15261 (N_15261,N_13635,N_12983);
and U15262 (N_15262,N_12591,N_13402);
nand U15263 (N_15263,N_14702,N_12911);
nand U15264 (N_15264,N_12503,N_14712);
and U15265 (N_15265,N_14360,N_12729);
or U15266 (N_15266,N_14260,N_14726);
xnor U15267 (N_15267,N_13975,N_14320);
and U15268 (N_15268,N_13702,N_13329);
and U15269 (N_15269,N_14084,N_13127);
nand U15270 (N_15270,N_14899,N_12888);
nor U15271 (N_15271,N_14025,N_14988);
nand U15272 (N_15272,N_13026,N_14153);
or U15273 (N_15273,N_12554,N_12828);
or U15274 (N_15274,N_13996,N_14750);
nor U15275 (N_15275,N_12968,N_14487);
or U15276 (N_15276,N_14731,N_13295);
or U15277 (N_15277,N_14636,N_13809);
xnor U15278 (N_15278,N_12789,N_13864);
nand U15279 (N_15279,N_14510,N_13109);
nand U15280 (N_15280,N_12802,N_14104);
nand U15281 (N_15281,N_13423,N_13906);
nor U15282 (N_15282,N_14986,N_13182);
nor U15283 (N_15283,N_13560,N_12606);
nand U15284 (N_15284,N_14666,N_14400);
and U15285 (N_15285,N_13832,N_14255);
or U15286 (N_15286,N_13643,N_12505);
xor U15287 (N_15287,N_14896,N_14734);
and U15288 (N_15288,N_13042,N_12561);
and U15289 (N_15289,N_14930,N_13031);
or U15290 (N_15290,N_14323,N_14704);
and U15291 (N_15291,N_12532,N_13715);
and U15292 (N_15292,N_13787,N_13111);
xnor U15293 (N_15293,N_13990,N_14219);
xor U15294 (N_15294,N_12902,N_12938);
xor U15295 (N_15295,N_14520,N_14601);
or U15296 (N_15296,N_12823,N_13067);
xor U15297 (N_15297,N_14256,N_13484);
and U15298 (N_15298,N_14914,N_12903);
nor U15299 (N_15299,N_14203,N_13074);
xnor U15300 (N_15300,N_13540,N_12861);
nor U15301 (N_15301,N_12929,N_14070);
or U15302 (N_15302,N_13346,N_13373);
or U15303 (N_15303,N_14455,N_12913);
and U15304 (N_15304,N_13867,N_13877);
or U15305 (N_15305,N_14212,N_12773);
and U15306 (N_15306,N_13316,N_13890);
or U15307 (N_15307,N_12599,N_14923);
and U15308 (N_15308,N_12650,N_14667);
or U15309 (N_15309,N_13045,N_13623);
and U15310 (N_15310,N_12625,N_14762);
nand U15311 (N_15311,N_13836,N_14581);
or U15312 (N_15312,N_14909,N_14263);
and U15313 (N_15313,N_14139,N_13299);
and U15314 (N_15314,N_13667,N_12699);
nand U15315 (N_15315,N_12621,N_14650);
and U15316 (N_15316,N_14172,N_14504);
nand U15317 (N_15317,N_13104,N_13759);
or U15318 (N_15318,N_13905,N_13411);
and U15319 (N_15319,N_13753,N_13651);
and U15320 (N_15320,N_14178,N_14794);
nand U15321 (N_15321,N_12686,N_14063);
or U15322 (N_15322,N_12833,N_13229);
nor U15323 (N_15323,N_13014,N_12517);
nor U15324 (N_15324,N_14721,N_13469);
or U15325 (N_15325,N_12748,N_13048);
xor U15326 (N_15326,N_13514,N_14275);
nand U15327 (N_15327,N_12562,N_14067);
nor U15328 (N_15328,N_13187,N_13279);
xnor U15329 (N_15329,N_14686,N_14633);
xor U15330 (N_15330,N_14610,N_14399);
and U15331 (N_15331,N_12690,N_14420);
nor U15332 (N_15332,N_14085,N_13653);
or U15333 (N_15333,N_14683,N_12673);
nand U15334 (N_15334,N_13714,N_13858);
and U15335 (N_15335,N_14548,N_13219);
and U15336 (N_15336,N_14295,N_13995);
or U15337 (N_15337,N_13011,N_14701);
nand U15338 (N_15338,N_13128,N_12735);
and U15339 (N_15339,N_14322,N_14718);
nor U15340 (N_15340,N_14565,N_13537);
xnor U15341 (N_15341,N_14858,N_12585);
nor U15342 (N_15342,N_14053,N_13489);
and U15343 (N_15343,N_14931,N_12787);
and U15344 (N_15344,N_12527,N_12855);
xor U15345 (N_15345,N_14698,N_14774);
nor U15346 (N_15346,N_12520,N_13289);
xor U15347 (N_15347,N_12988,N_13949);
xnor U15348 (N_15348,N_13193,N_14625);
or U15349 (N_15349,N_13972,N_12525);
and U15350 (N_15350,N_14668,N_12609);
xor U15351 (N_15351,N_13464,N_14237);
and U15352 (N_15352,N_13271,N_14901);
and U15353 (N_15353,N_14635,N_13959);
or U15354 (N_15354,N_13133,N_13616);
nand U15355 (N_15355,N_14876,N_13911);
nand U15356 (N_15356,N_14900,N_14437);
or U15357 (N_15357,N_12996,N_12538);
xnor U15358 (N_15358,N_14845,N_13150);
xnor U15359 (N_15359,N_12845,N_14533);
nor U15360 (N_15360,N_14170,N_13092);
nand U15361 (N_15361,N_12647,N_13130);
and U15362 (N_15362,N_13981,N_14553);
or U15363 (N_15363,N_13951,N_13834);
and U15364 (N_15364,N_13572,N_13853);
xnor U15365 (N_15365,N_14547,N_14384);
and U15366 (N_15366,N_14333,N_13612);
or U15367 (N_15367,N_13671,N_13304);
or U15368 (N_15368,N_13971,N_13041);
xnor U15369 (N_15369,N_14885,N_13202);
nor U15370 (N_15370,N_14101,N_12737);
xor U15371 (N_15371,N_13494,N_14943);
or U15372 (N_15372,N_12644,N_14179);
nor U15373 (N_15373,N_12827,N_14166);
or U15374 (N_15374,N_12926,N_14782);
xor U15375 (N_15375,N_12866,N_13937);
nor U15376 (N_15376,N_13815,N_13159);
xnor U15377 (N_15377,N_13510,N_13249);
xnor U15378 (N_15378,N_14613,N_14406);
nand U15379 (N_15379,N_14846,N_14993);
and U15380 (N_15380,N_12871,N_14672);
nand U15381 (N_15381,N_12502,N_13794);
xor U15382 (N_15382,N_14951,N_14387);
nand U15383 (N_15383,N_14112,N_14770);
or U15384 (N_15384,N_14999,N_14430);
and U15385 (N_15385,N_14500,N_14883);
nand U15386 (N_15386,N_13644,N_13273);
nor U15387 (N_15387,N_14611,N_13418);
nor U15388 (N_15388,N_14629,N_13005);
or U15389 (N_15389,N_14373,N_13500);
nand U15390 (N_15390,N_13700,N_13093);
xnor U15391 (N_15391,N_14778,N_13162);
xor U15392 (N_15392,N_13224,N_13377);
or U15393 (N_15393,N_13800,N_13546);
and U15394 (N_15394,N_12967,N_13843);
and U15395 (N_15395,N_14432,N_13539);
and U15396 (N_15396,N_13239,N_13132);
xnor U15397 (N_15397,N_14677,N_13294);
nor U15398 (N_15398,N_12708,N_13189);
nor U15399 (N_15399,N_14223,N_14254);
xor U15400 (N_15400,N_14862,N_13476);
and U15401 (N_15401,N_12613,N_14603);
or U15402 (N_15402,N_14800,N_13155);
xnor U15403 (N_15403,N_13472,N_14825);
xnor U15404 (N_15404,N_14566,N_14146);
and U15405 (N_15405,N_14226,N_12889);
xnor U15406 (N_15406,N_13796,N_13602);
nor U15407 (N_15407,N_13625,N_12925);
and U15408 (N_15408,N_13554,N_13020);
and U15409 (N_15409,N_14312,N_12948);
xnor U15410 (N_15410,N_14539,N_14544);
xnor U15411 (N_15411,N_12705,N_13983);
nand U15412 (N_15412,N_14130,N_12859);
xor U15413 (N_15413,N_12839,N_14534);
xor U15414 (N_15414,N_14798,N_12540);
and U15415 (N_15415,N_12950,N_13661);
and U15416 (N_15416,N_14332,N_13569);
or U15417 (N_15417,N_14428,N_14535);
or U15418 (N_15418,N_13378,N_12586);
xnor U15419 (N_15419,N_12772,N_13909);
or U15420 (N_15420,N_12563,N_14474);
nand U15421 (N_15421,N_13736,N_14064);
nor U15422 (N_15422,N_13831,N_14151);
or U15423 (N_15423,N_14215,N_12738);
and U15424 (N_15424,N_14075,N_14004);
or U15425 (N_15425,N_13594,N_12665);
and U15426 (N_15426,N_14077,N_12759);
or U15427 (N_15427,N_12723,N_12843);
xnor U15428 (N_15428,N_14089,N_14408);
xnor U15429 (N_15429,N_13735,N_14129);
xor U15430 (N_15430,N_13208,N_14189);
and U15431 (N_15431,N_12588,N_14604);
xor U15432 (N_15432,N_12989,N_12653);
nand U15433 (N_15433,N_13097,N_14291);
nand U15434 (N_15434,N_14177,N_14824);
or U15435 (N_15435,N_14790,N_13499);
and U15436 (N_15436,N_14124,N_14837);
and U15437 (N_15437,N_13647,N_14479);
nand U15438 (N_15438,N_13920,N_12891);
nor U15439 (N_15439,N_14382,N_13312);
or U15440 (N_15440,N_14183,N_13175);
nand U15441 (N_15441,N_12951,N_13533);
nor U15442 (N_15442,N_14325,N_13966);
nor U15443 (N_15443,N_13749,N_13608);
xor U15444 (N_15444,N_13191,N_13897);
nor U15445 (N_15445,N_14154,N_13251);
xnor U15446 (N_15446,N_13164,N_14200);
xnor U15447 (N_15447,N_13017,N_13380);
nor U15448 (N_15448,N_12731,N_13681);
nand U15449 (N_15449,N_12769,N_12662);
and U15450 (N_15450,N_12688,N_13267);
xnor U15451 (N_15451,N_12725,N_13772);
or U15452 (N_15452,N_12678,N_12620);
nand U15453 (N_15453,N_14475,N_13666);
or U15454 (N_15454,N_13465,N_12652);
and U15455 (N_15455,N_14187,N_13204);
nand U15456 (N_15456,N_13934,N_13947);
or U15457 (N_15457,N_13597,N_13579);
nand U15458 (N_15458,N_14358,N_13037);
and U15459 (N_15459,N_12675,N_13056);
and U15460 (N_15460,N_12556,N_13326);
and U15461 (N_15461,N_14017,N_13331);
and U15462 (N_15462,N_13640,N_13989);
xnor U15463 (N_15463,N_13770,N_14073);
nand U15464 (N_15464,N_13406,N_13070);
xor U15465 (N_15465,N_13738,N_13961);
or U15466 (N_15466,N_14434,N_13365);
nor U15467 (N_15467,N_13280,N_13237);
or U15468 (N_15468,N_13180,N_12840);
nor U15469 (N_15469,N_12858,N_13390);
and U15470 (N_15470,N_13574,N_14281);
nand U15471 (N_15471,N_12639,N_12870);
or U15472 (N_15472,N_13792,N_13582);
nand U15473 (N_15473,N_13604,N_12857);
and U15474 (N_15474,N_14495,N_14985);
xor U15475 (N_15475,N_13125,N_13592);
xor U15476 (N_15476,N_13194,N_14471);
and U15477 (N_15477,N_14802,N_14752);
nor U15478 (N_15478,N_14875,N_14285);
nor U15479 (N_15479,N_14484,N_14316);
xor U15480 (N_15480,N_13675,N_12767);
nand U15481 (N_15481,N_14894,N_13690);
xor U15482 (N_15482,N_12791,N_12777);
nor U15483 (N_15483,N_14385,N_13581);
or U15484 (N_15484,N_13256,N_13950);
or U15485 (N_15485,N_14359,N_12537);
nor U15486 (N_15486,N_12970,N_14427);
nor U15487 (N_15487,N_13161,N_14745);
nand U15488 (N_15488,N_14036,N_13059);
nor U15489 (N_15489,N_14511,N_14365);
nor U15490 (N_15490,N_14232,N_14488);
xnor U15491 (N_15491,N_13362,N_13288);
or U15492 (N_15492,N_13449,N_13006);
xnor U15493 (N_15493,N_14937,N_14403);
or U15494 (N_15494,N_13158,N_14671);
and U15495 (N_15495,N_13361,N_13859);
xor U15496 (N_15496,N_13072,N_12515);
or U15497 (N_15497,N_14034,N_14903);
nand U15498 (N_15498,N_12985,N_13455);
nand U15499 (N_15499,N_14131,N_13743);
and U15500 (N_15500,N_14433,N_12768);
nor U15501 (N_15501,N_14654,N_13978);
nand U15502 (N_15502,N_12638,N_12862);
nand U15503 (N_15503,N_13368,N_14366);
or U15504 (N_15504,N_13285,N_12992);
nand U15505 (N_15505,N_13412,N_12830);
xnor U15506 (N_15506,N_14723,N_14110);
nand U15507 (N_15507,N_14461,N_12797);
or U15508 (N_15508,N_14247,N_14185);
or U15509 (N_15509,N_14368,N_14784);
nor U15510 (N_15510,N_12733,N_13917);
xor U15511 (N_15511,N_12894,N_12762);
xnor U15512 (N_15512,N_13526,N_14730);
xor U15513 (N_15513,N_13151,N_13883);
nor U15514 (N_15514,N_13078,N_13908);
nor U15515 (N_15515,N_14527,N_14537);
and U15516 (N_15516,N_13780,N_13211);
xor U15517 (N_15517,N_12648,N_12593);
nor U15518 (N_15518,N_13071,N_13296);
and U15519 (N_15519,N_13230,N_14118);
nor U15520 (N_15520,N_14523,N_14361);
xor U15521 (N_15521,N_14148,N_14593);
and U15522 (N_15522,N_13855,N_13094);
or U15523 (N_15523,N_14928,N_12522);
xnor U15524 (N_15524,N_12825,N_12607);
nor U15525 (N_15525,N_13844,N_13009);
or U15526 (N_15526,N_13049,N_13222);
nor U15527 (N_15527,N_13434,N_14700);
or U15528 (N_15528,N_13828,N_14220);
nand U15529 (N_15529,N_14065,N_14264);
nand U15530 (N_15530,N_14035,N_12837);
and U15531 (N_15531,N_13430,N_14505);
and U15532 (N_15532,N_13266,N_13108);
or U15533 (N_15533,N_12863,N_14349);
or U15534 (N_15534,N_14422,N_14840);
nand U15535 (N_15535,N_13117,N_13970);
and U15536 (N_15536,N_13003,N_12543);
xor U15537 (N_15537,N_14490,N_13741);
xor U15538 (N_15538,N_12518,N_13367);
and U15539 (N_15539,N_13432,N_13835);
nor U15540 (N_15540,N_12619,N_12884);
nor U15541 (N_15541,N_13232,N_14195);
or U15542 (N_15542,N_13134,N_13694);
nand U15543 (N_15543,N_12576,N_14578);
nand U15544 (N_15544,N_12910,N_12702);
or U15545 (N_15545,N_13779,N_14596);
nand U15546 (N_15546,N_14509,N_14579);
and U15547 (N_15547,N_13573,N_13532);
nand U15548 (N_15548,N_13710,N_13000);
nand U15549 (N_15549,N_14111,N_13940);
nor U15550 (N_15550,N_14597,N_13802);
nor U15551 (N_15551,N_13518,N_14873);
or U15552 (N_15552,N_14140,N_13065);
and U15553 (N_15553,N_13722,N_13717);
nand U15554 (N_15554,N_13021,N_12582);
or U15555 (N_15555,N_14379,N_13023);
xor U15556 (N_15556,N_14047,N_13080);
nor U15557 (N_15557,N_13825,N_14508);
and U15558 (N_15558,N_13588,N_13649);
nor U15559 (N_15559,N_13213,N_13099);
or U15560 (N_15560,N_13930,N_13393);
xor U15561 (N_15561,N_14764,N_13530);
xor U15562 (N_15562,N_13882,N_12501);
nor U15563 (N_15563,N_14600,N_13938);
and U15564 (N_15564,N_12778,N_14856);
and U15565 (N_15565,N_14588,N_13274);
or U15566 (N_15566,N_14904,N_13871);
or U15567 (N_15567,N_13726,N_12958);
and U15568 (N_15568,N_13315,N_13334);
xnor U15569 (N_15569,N_13948,N_14685);
xor U15570 (N_15570,N_14477,N_13845);
nor U15571 (N_15571,N_14491,N_12842);
and U15572 (N_15572,N_13247,N_13463);
xor U15573 (N_15573,N_13253,N_12991);
and U15574 (N_15574,N_13123,N_13388);
xnor U15575 (N_15575,N_14128,N_13721);
or U15576 (N_15576,N_14449,N_14797);
or U15577 (N_15577,N_14707,N_13320);
nor U15578 (N_15578,N_13840,N_14249);
and U15579 (N_15579,N_13107,N_12512);
nand U15580 (N_15580,N_12977,N_14472);
nand U15581 (N_15581,N_14917,N_14678);
nand U15582 (N_15582,N_13242,N_14706);
xor U15583 (N_15583,N_14619,N_14748);
xor U15584 (N_15584,N_13885,N_14015);
xnor U15585 (N_15585,N_14965,N_12962);
or U15586 (N_15586,N_12879,N_13564);
or U15587 (N_15587,N_14739,N_12770);
and U15588 (N_15588,N_14805,N_13330);
and U15589 (N_15589,N_12504,N_13701);
nand U15590 (N_15590,N_12868,N_14087);
or U15591 (N_15591,N_13517,N_14961);
nor U15592 (N_15592,N_13324,N_14290);
or U15593 (N_15593,N_14278,N_14628);
nor U15594 (N_15594,N_14968,N_14299);
xnor U15595 (N_15595,N_13355,N_13525);
and U15596 (N_15596,N_12784,N_13879);
nand U15597 (N_15597,N_12811,N_13775);
nor U15598 (N_15598,N_14419,N_13740);
xnor U15599 (N_15599,N_13205,N_14545);
nor U15600 (N_15600,N_14994,N_14692);
nand U15601 (N_15601,N_14637,N_13442);
xor U15602 (N_15602,N_14725,N_14041);
or U15603 (N_15603,N_14804,N_12560);
and U15604 (N_15604,N_14057,N_13379);
xor U15605 (N_15605,N_14594,N_13814);
or U15606 (N_15606,N_12655,N_13963);
nor U15607 (N_15607,N_12670,N_12990);
nor U15608 (N_15608,N_13764,N_14550);
nor U15609 (N_15609,N_13737,N_14812);
nor U15610 (N_15610,N_14855,N_14235);
or U15611 (N_15611,N_13297,N_14913);
or U15612 (N_15612,N_14502,N_13583);
nor U15613 (N_15613,N_14852,N_14018);
and U15614 (N_15614,N_12624,N_14513);
nand U15615 (N_15615,N_14575,N_14149);
xor U15616 (N_15616,N_14591,N_12896);
or U15617 (N_15617,N_13282,N_14298);
or U15618 (N_15618,N_13163,N_13901);
nand U15619 (N_15619,N_14283,N_14370);
nand U15620 (N_15620,N_14956,N_14940);
or U15621 (N_15621,N_12920,N_14279);
nor U15622 (N_15622,N_13309,N_14417);
nor U15623 (N_15623,N_13457,N_14367);
nand U15624 (N_15624,N_13414,N_12603);
nor U15625 (N_15625,N_13122,N_13891);
nand U15626 (N_15626,N_14626,N_13269);
nand U15627 (N_15627,N_14530,N_13508);
or U15628 (N_15628,N_14769,N_14171);
or U15629 (N_15629,N_13758,N_14372);
nor U15630 (N_15630,N_13087,N_14964);
xnor U15631 (N_15631,N_14280,N_12793);
nor U15632 (N_15632,N_12676,N_14801);
xnor U15633 (N_15633,N_13468,N_14567);
xnor U15634 (N_15634,N_14728,N_14000);
or U15635 (N_15635,N_12596,N_13216);
nor U15636 (N_15636,N_12916,N_12853);
nor U15637 (N_15637,N_13144,N_12552);
xnor U15638 (N_15638,N_13676,N_13290);
nor U15639 (N_15639,N_13374,N_13918);
and U15640 (N_15640,N_14679,N_13570);
xor U15641 (N_15641,N_14657,N_14043);
xnor U15642 (N_15642,N_12633,N_13605);
nor U15643 (N_15643,N_13043,N_12707);
or U15644 (N_15644,N_14448,N_14772);
nor U15645 (N_15645,N_14356,N_14150);
or U15646 (N_15646,N_13392,N_14300);
nand U15647 (N_15647,N_14469,N_13250);
xor U15648 (N_15648,N_13257,N_12700);
nand U15649 (N_15649,N_14098,N_13283);
or U15650 (N_15650,N_14374,N_14355);
nand U15651 (N_15651,N_14242,N_12940);
nor U15652 (N_15652,N_12516,N_13847);
xnor U15653 (N_15653,N_12752,N_14082);
nor U15654 (N_15654,N_14857,N_12687);
and U15655 (N_15655,N_14559,N_14737);
xnor U15656 (N_15656,N_13019,N_12628);
nand U15657 (N_15657,N_14345,N_13893);
or U15658 (N_15658,N_14058,N_14818);
or U15659 (N_15659,N_13032,N_13231);
and U15660 (N_15660,N_13955,N_13593);
or U15661 (N_15661,N_13614,N_13709);
nand U15662 (N_15662,N_13811,N_13033);
xnor U15663 (N_15663,N_13793,N_14196);
nor U15664 (N_15664,N_13984,N_13319);
and U15665 (N_15665,N_12798,N_14315);
nand U15666 (N_15666,N_13004,N_13015);
and U15667 (N_15667,N_14583,N_13805);
nor U15668 (N_15668,N_13766,N_13353);
nand U15669 (N_15669,N_13143,N_12528);
and U15670 (N_15670,N_14607,N_14445);
nor U15671 (N_15671,N_14364,N_12878);
xnor U15672 (N_15672,N_12602,N_13542);
or U15673 (N_15673,N_13638,N_12935);
xor U15674 (N_15674,N_13381,N_14287);
nand U15675 (N_15675,N_14618,N_14792);
or U15676 (N_15676,N_12915,N_14687);
xnor U15677 (N_15677,N_14029,N_14975);
or U15678 (N_15678,N_12819,N_13591);
and U15679 (N_15679,N_13090,N_14438);
nand U15680 (N_15680,N_13900,N_13027);
or U15681 (N_15681,N_14643,N_14887);
and U15682 (N_15682,N_14105,N_13945);
and U15683 (N_15683,N_14079,N_13360);
and U15684 (N_15684,N_12817,N_13806);
xnor U15685 (N_15685,N_13185,N_13571);
xnor U15686 (N_15686,N_12893,N_13912);
or U15687 (N_15687,N_14585,N_12571);
nor U15688 (N_15688,N_13754,N_13884);
or U15689 (N_15689,N_14939,N_14966);
xor U15690 (N_15690,N_12544,N_13563);
nand U15691 (N_15691,N_14257,N_14971);
xnor U15692 (N_15692,N_14673,N_13047);
and U15693 (N_15693,N_13670,N_12931);
nor U15694 (N_15694,N_12924,N_14435);
nand U15695 (N_15695,N_12820,N_12953);
xnor U15696 (N_15696,N_12809,N_14617);
nor U15697 (N_15697,N_14815,N_14092);
nor U15698 (N_15698,N_14525,N_12881);
or U15699 (N_15699,N_14542,N_13819);
nor U15700 (N_15700,N_12728,N_12918);
xor U15701 (N_15701,N_14194,N_13875);
or U15702 (N_15702,N_13550,N_14623);
nor U15703 (N_15703,N_13473,N_12869);
nor U15704 (N_15704,N_12912,N_14874);
nor U15705 (N_15705,N_14388,N_14108);
and U15706 (N_15706,N_14927,N_13725);
nand U15707 (N_15707,N_14560,N_12720);
or U15708 (N_15708,N_14902,N_13538);
xor U15709 (N_15709,N_14013,N_13559);
nand U15710 (N_15710,N_14756,N_14689);
or U15711 (N_15711,N_12627,N_14655);
nand U15712 (N_15712,N_13739,N_14125);
nor U15713 (N_15713,N_13238,N_14307);
xor U15714 (N_15714,N_14396,N_12844);
xor U15715 (N_15715,N_13448,N_13195);
and U15716 (N_15716,N_12775,N_14783);
nor U15717 (N_15717,N_12616,N_13259);
xnor U15718 (N_15718,N_14423,N_13791);
and U15719 (N_15719,N_12683,N_12717);
xnor U15720 (N_15720,N_14715,N_13462);
nand U15721 (N_15721,N_14835,N_14390);
nand U15722 (N_15722,N_13416,N_12691);
and U15723 (N_15723,N_13447,N_14002);
and U15724 (N_15724,N_13404,N_14302);
or U15725 (N_15725,N_14615,N_13348);
and U15726 (N_15726,N_14207,N_13100);
or U15727 (N_15727,N_13553,N_13913);
nand U15728 (N_15728,N_13038,N_12904);
nand U15729 (N_15729,N_13939,N_13287);
xnor U15730 (N_15730,N_13340,N_12914);
or U15731 (N_15731,N_13095,N_14205);
nand U15732 (N_15732,N_14069,N_13575);
nand U15733 (N_15733,N_13657,N_13356);
or U15734 (N_15734,N_14157,N_13470);
and U15735 (N_15735,N_12669,N_13688);
nand U15736 (N_15736,N_12623,N_12821);
or U15737 (N_15737,N_14122,N_14251);
and U15738 (N_15738,N_14793,N_13096);
and U15739 (N_15739,N_12947,N_13350);
and U15740 (N_15740,N_14897,N_14478);
and U15741 (N_15741,N_14884,N_12711);
and U15742 (N_15742,N_13807,N_14828);
or U15743 (N_15743,N_13769,N_13931);
and U15744 (N_15744,N_14918,N_14867);
xor U15745 (N_15745,N_14331,N_14259);
or U15746 (N_15746,N_12810,N_13422);
or U15747 (N_15747,N_14608,N_13926);
xnor U15748 (N_15748,N_12730,N_13902);
nor U15749 (N_15749,N_14048,N_13504);
xnor U15750 (N_15750,N_12754,N_14329);
nand U15751 (N_15751,N_13804,N_12533);
nand U15752 (N_15752,N_13629,N_14473);
nand U15753 (N_15753,N_13543,N_13887);
nand U15754 (N_15754,N_14910,N_14908);
nand U15755 (N_15755,N_14995,N_13255);
nor U15756 (N_15756,N_14008,N_14467);
and U15757 (N_15757,N_12771,N_13417);
or U15758 (N_15758,N_12834,N_14121);
or U15759 (N_15759,N_14697,N_14641);
and U15760 (N_15760,N_14714,N_13246);
xnor U15761 (N_15761,N_13141,N_13106);
and U15762 (N_15762,N_13944,N_12836);
and U15763 (N_15763,N_14480,N_14182);
nand U15764 (N_15764,N_13878,N_14676);
or U15765 (N_15765,N_12511,N_12867);
xor U15766 (N_15766,N_12997,N_12781);
nor U15767 (N_15767,N_12760,N_14777);
or U15768 (N_15768,N_13731,N_14088);
nor U15769 (N_15769,N_14978,N_14191);
and U15770 (N_15770,N_14574,N_14005);
nand U15771 (N_15771,N_14788,N_13245);
xor U15772 (N_15772,N_12589,N_13576);
or U15773 (N_15773,N_13706,N_12722);
or U15774 (N_15774,N_14180,N_14826);
nand U15775 (N_15775,N_12677,N_14132);
nand U15776 (N_15776,N_13952,N_14208);
or U15777 (N_15777,N_14606,N_14942);
and U15778 (N_15778,N_14193,N_13746);
nand U15779 (N_15779,N_13833,N_13303);
nor U15780 (N_15780,N_13729,N_12804);
nand U15781 (N_15781,N_14310,N_13286);
or U15782 (N_15782,N_14021,N_13716);
or U15783 (N_15783,N_14109,N_14414);
nand U15784 (N_15784,N_12877,N_14934);
and U15785 (N_15785,N_12726,N_14911);
nand U15786 (N_15786,N_13695,N_13085);
and U15787 (N_15787,N_14742,N_13034);
nand U15788 (N_15788,N_13421,N_13600);
and U15789 (N_15789,N_14708,N_14338);
nor U15790 (N_15790,N_14526,N_14266);
nor U15791 (N_15791,N_12666,N_13173);
nand U15792 (N_15792,N_12661,N_12553);
and U15793 (N_15793,N_14138,N_14819);
xnor U15794 (N_15794,N_13927,N_14833);
or U15795 (N_15795,N_14094,N_12646);
and U15796 (N_15796,N_13744,N_14272);
and U15797 (N_15797,N_14252,N_13311);
nand U15798 (N_15798,N_14497,N_13637);
nor U15799 (N_15799,N_12847,N_13960);
nand U15800 (N_15800,N_13354,N_14515);
and U15801 (N_15801,N_14974,N_14973);
or U15802 (N_15802,N_13603,N_14760);
or U15803 (N_15803,N_14236,N_13452);
xor U15804 (N_15804,N_13976,N_13619);
or U15805 (N_15805,N_13145,N_13491);
xor U15806 (N_15806,N_13401,N_13270);
nand U15807 (N_15807,N_12664,N_14199);
nand U15808 (N_15808,N_13113,N_13172);
xnor U15809 (N_15809,N_12636,N_14997);
nand U15810 (N_15810,N_12806,N_14627);
or U15811 (N_15811,N_13761,N_13607);
or U15812 (N_15812,N_14352,N_12635);
or U15813 (N_15813,N_12801,N_14465);
or U15814 (N_15814,N_13483,N_13310);
or U15815 (N_15815,N_14808,N_12927);
nand U15816 (N_15816,N_13552,N_13860);
nor U15817 (N_15817,N_13233,N_13456);
and U15818 (N_15818,N_12608,N_13284);
nand U15819 (N_15819,N_14051,N_13384);
and U15820 (N_15820,N_13628,N_14773);
xor U15821 (N_15821,N_14398,N_14944);
or U15822 (N_15822,N_14984,N_12630);
nand U15823 (N_15823,N_12818,N_13343);
nand U15824 (N_15824,N_14854,N_13567);
and U15825 (N_15825,N_14059,N_13136);
xnor U15826 (N_15826,N_13055,N_13622);
and U15827 (N_15827,N_14225,N_12513);
and U15828 (N_15828,N_14921,N_12575);
or U15829 (N_15829,N_13086,N_12907);
nand U15830 (N_15830,N_13630,N_14563);
and U15831 (N_15831,N_13589,N_12960);
or U15832 (N_15832,N_13066,N_14347);
nand U15833 (N_15833,N_13954,N_13979);
nor U15834 (N_15834,N_14046,N_14080);
or U15835 (N_15835,N_12987,N_12993);
xnor U15836 (N_15836,N_14891,N_14489);
nand U15837 (N_15837,N_14684,N_13454);
and U15838 (N_15838,N_14144,N_14503);
and U15839 (N_15839,N_14521,N_14747);
nand U15840 (N_15840,N_14703,N_13490);
nand U15841 (N_15841,N_14834,N_14447);
or U15842 (N_15842,N_14693,N_14919);
and U15843 (N_15843,N_13919,N_13140);
and U15844 (N_15844,N_13121,N_12959);
nand U15845 (N_15845,N_13192,N_14912);
nand U15846 (N_15846,N_14881,N_14799);
nand U15847 (N_15847,N_14485,N_12564);
nor U15848 (N_15848,N_14807,N_13207);
xnor U15849 (N_15849,N_13063,N_13029);
and U15850 (N_15850,N_13426,N_13051);
nor U15851 (N_15851,N_14458,N_14204);
nor U15852 (N_15852,N_13001,N_12632);
xnor U15853 (N_15853,N_14838,N_13677);
and U15854 (N_15854,N_13060,N_14963);
xnor U15855 (N_15855,N_14647,N_12583);
xor U15856 (N_15856,N_12689,N_12578);
or U15857 (N_15857,N_12887,N_14201);
or U15858 (N_15858,N_12696,N_12882);
and U15859 (N_15859,N_13339,N_13492);
nand U15860 (N_15860,N_12590,N_14749);
xnor U15861 (N_15861,N_12892,N_14311);
and U15862 (N_15862,N_13101,N_14282);
nor U15863 (N_15863,N_13765,N_12937);
nor U15864 (N_15864,N_14877,N_14803);
nand U15865 (N_15865,N_13376,N_14412);
nand U15866 (N_15866,N_12703,N_13198);
and U15867 (N_15867,N_13786,N_14099);
nand U15868 (N_15868,N_14549,N_13439);
nor U15869 (N_15869,N_13116,N_14498);
or U15870 (N_15870,N_13946,N_14663);
nand U15871 (N_15871,N_12812,N_14231);
and U15872 (N_15872,N_12706,N_14391);
and U15873 (N_15873,N_12649,N_12900);
xnor U15874 (N_15874,N_13977,N_13668);
or U15875 (N_15875,N_12549,N_14066);
nor U15876 (N_15876,N_12742,N_14330);
or U15877 (N_15877,N_13226,N_12736);
and U15878 (N_15878,N_13012,N_13157);
and U15879 (N_15879,N_14229,N_14340);
and U15880 (N_15880,N_14791,N_14470);
xor U15881 (N_15881,N_13221,N_13496);
and U15882 (N_15882,N_14042,N_14143);
and U15883 (N_15883,N_13357,N_13689);
or U15884 (N_15884,N_14809,N_13785);
and U15885 (N_15885,N_13872,N_12718);
nor U15886 (N_15886,N_14561,N_14395);
and U15887 (N_15887,N_14028,N_14646);
or U15888 (N_15888,N_14343,N_13010);
xnor U15889 (N_15889,N_13631,N_14720);
or U15890 (N_15890,N_14107,N_13383);
nor U15891 (N_15891,N_12955,N_14304);
nor U15892 (N_15892,N_13718,N_13443);
or U15893 (N_15893,N_14853,N_14014);
nand U15894 (N_15894,N_14929,N_12941);
or U15895 (N_15895,N_13648,N_14482);
nand U15896 (N_15896,N_13138,N_13018);
nand U15897 (N_15897,N_12657,N_13263);
xor U15898 (N_15898,N_14214,N_12745);
nor U15899 (N_15899,N_13227,N_13728);
and U15900 (N_15900,N_14776,N_12942);
xor U15901 (N_15901,N_14440,N_13210);
nand U15902 (N_15902,N_14056,N_13186);
or U15903 (N_15903,N_14744,N_14870);
or U15904 (N_15904,N_13865,N_13399);
or U15905 (N_15905,N_13225,N_12783);
nor U15906 (N_15906,N_12755,N_14787);
or U15907 (N_15907,N_13197,N_14246);
xnor U15908 (N_15908,N_14970,N_14055);
nor U15909 (N_15909,N_14062,N_12716);
or U15910 (N_15910,N_14339,N_13762);
or U15911 (N_15911,N_14163,N_13755);
xor U15912 (N_15912,N_14640,N_14860);
nor U15913 (N_15913,N_13962,N_13561);
or U15914 (N_15914,N_14303,N_14717);
xnor U15915 (N_15915,N_13084,N_12856);
or U15916 (N_15916,N_13069,N_14680);
nand U15917 (N_15917,N_14820,N_13929);
xnor U15918 (N_15918,N_14392,N_14103);
nand U15919 (N_15919,N_12545,N_13956);
nand U15920 (N_15920,N_14705,N_14209);
or U15921 (N_15921,N_14982,N_14050);
nor U15922 (N_15922,N_13531,N_12679);
nand U15923 (N_15923,N_13181,N_13590);
nand U15924 (N_15924,N_14735,N_13682);
xnor U15925 (N_15925,N_14649,N_14159);
nor U15926 (N_15926,N_13896,N_12651);
xor U15927 (N_15927,N_13459,N_14416);
nor U15928 (N_15928,N_13344,N_12751);
nand U15929 (N_15929,N_14197,N_12824);
nand U15930 (N_15930,N_13509,N_13022);
nand U15931 (N_15931,N_14864,N_13562);
and U15932 (N_15932,N_13397,N_14377);
nand U15933 (N_15933,N_14418,N_13044);
nor U15934 (N_15934,N_14409,N_13115);
and U15935 (N_15935,N_12595,N_13342);
xnor U15936 (N_15936,N_13826,N_14160);
xor U15937 (N_15937,N_14424,N_13615);
xor U15938 (N_15938,N_14935,N_13461);
and U15939 (N_15939,N_12519,N_13816);
xor U15940 (N_15940,N_14456,N_12680);
nand U15941 (N_15941,N_12999,N_13998);
xor U15942 (N_15942,N_12756,N_14019);
and U15943 (N_15943,N_12890,N_13152);
xor U15944 (N_15944,N_13520,N_14878);
and U15945 (N_15945,N_13620,N_12813);
nor U15946 (N_15946,N_12909,N_13166);
nor U15947 (N_15947,N_14710,N_13660);
xnor U15948 (N_15948,N_12712,N_14958);
and U15949 (N_15949,N_14761,N_12659);
xor U15950 (N_15950,N_13305,N_14102);
xor U15951 (N_15951,N_13757,N_14216);
nor U15952 (N_15952,N_12883,N_13633);
and U15953 (N_15953,N_14722,N_13313);
or U15954 (N_15954,N_14632,N_13965);
nand U15955 (N_15955,N_14314,N_12921);
or U15956 (N_15956,N_14240,N_14294);
and U15957 (N_15957,N_14682,N_14068);
nor U15958 (N_15958,N_13720,N_14789);
nand U15959 (N_15959,N_12865,N_13359);
nand U15960 (N_15960,N_14346,N_14659);
or U15961 (N_15961,N_13110,N_14499);
and U15962 (N_15962,N_14031,N_13413);
nor U15963 (N_15963,N_13366,N_13685);
and U15964 (N_15964,N_12611,N_14972);
xor U15965 (N_15965,N_13126,N_13810);
xnor U15966 (N_15966,N_14945,N_14516);
or U15967 (N_15967,N_13165,N_14468);
or U15968 (N_15968,N_12757,N_12548);
nor U15969 (N_15969,N_14371,N_14120);
and U15970 (N_15970,N_13201,N_14543);
nand U15971 (N_15971,N_13662,N_13168);
nand U15972 (N_15972,N_14230,N_12873);
or U15973 (N_15973,N_12550,N_12780);
nor U15974 (N_15974,N_13663,N_13747);
xor U15975 (N_15975,N_14719,N_13969);
xnor U15976 (N_15976,N_14998,N_12776);
nand U15977 (N_15977,N_12542,N_12637);
or U15978 (N_15978,N_13137,N_12886);
nand U15979 (N_15979,N_14136,N_14905);
or U15980 (N_15980,N_13854,N_13524);
nand U15981 (N_15981,N_12514,N_14244);
xor U15982 (N_15982,N_12753,N_13415);
and U15983 (N_15983,N_14074,N_13824);
or U15984 (N_15984,N_14402,N_14576);
nor U15985 (N_15985,N_14147,N_12864);
nand U15986 (N_15986,N_14751,N_14119);
nor U15987 (N_15987,N_13409,N_13856);
xor U15988 (N_15988,N_13371,N_13708);
or U15989 (N_15989,N_14890,N_13986);
or U15990 (N_15990,N_12580,N_13547);
xor U15991 (N_15991,N_13692,N_14653);
and U15992 (N_15992,N_12618,N_13338);
or U15993 (N_15993,N_14007,N_14318);
and U15994 (N_15994,N_13089,N_13407);
or U15995 (N_15995,N_12610,N_13627);
or U15996 (N_15996,N_13120,N_13876);
nor U15997 (N_15997,N_12790,N_14268);
nand U15998 (N_15998,N_14466,N_14991);
or U15999 (N_15999,N_14167,N_13440);
nand U16000 (N_16000,N_12765,N_14375);
nor U16001 (N_16001,N_12634,N_13980);
nand U16002 (N_16002,N_14463,N_14871);
or U16003 (N_16003,N_14061,N_13915);
and U16004 (N_16004,N_12524,N_13585);
nand U16005 (N_16005,N_14446,N_13656);
xor U16006 (N_16006,N_13400,N_14224);
and U16007 (N_16007,N_12641,N_13046);
xor U16008 (N_16008,N_13535,N_12979);
nand U16009 (N_16009,N_13697,N_13982);
and U16010 (N_16010,N_12594,N_12536);
nand U16011 (N_16011,N_14746,N_12714);
nor U16012 (N_16012,N_14198,N_14011);
and U16013 (N_16013,N_14724,N_14850);
nand U16014 (N_16014,N_14174,N_13506);
and U16015 (N_16015,N_13586,N_13088);
and U16016 (N_16016,N_13119,N_14083);
nor U16017 (N_16017,N_13420,N_14426);
and U16018 (N_16018,N_13212,N_14872);
or U16019 (N_16019,N_13318,N_13632);
and U16020 (N_16020,N_13566,N_13405);
nor U16021 (N_16021,N_12612,N_12957);
nor U16022 (N_16022,N_12746,N_14569);
or U16023 (N_16023,N_13054,N_13933);
and U16024 (N_16024,N_14924,N_14383);
xor U16025 (N_16025,N_12829,N_14785);
and U16026 (N_16026,N_14476,N_13678);
nand U16027 (N_16027,N_14514,N_13850);
nor U16028 (N_16028,N_12710,N_12604);
and U16029 (N_16029,N_13664,N_13272);
xnor U16030 (N_16030,N_12758,N_12816);
nor U16031 (N_16031,N_13862,N_14622);
xnor U16032 (N_16032,N_14442,N_13711);
nor U16033 (N_16033,N_14181,N_13505);
or U16034 (N_16034,N_13475,N_13382);
xnor U16035 (N_16035,N_13730,N_14288);
nand U16036 (N_16036,N_12547,N_13752);
xnor U16037 (N_16037,N_13596,N_13008);
or U16038 (N_16038,N_14960,N_14609);
and U16039 (N_16039,N_13795,N_13813);
and U16040 (N_16040,N_14327,N_14313);
nor U16041 (N_16041,N_13278,N_13064);
and U16042 (N_16042,N_14481,N_13268);
or U16043 (N_16043,N_12526,N_12539);
xnor U16044 (N_16044,N_12685,N_14032);
xor U16045 (N_16045,N_14309,N_14518);
or U16046 (N_16046,N_13486,N_13502);
and U16047 (N_16047,N_13264,N_12500);
nand U16048 (N_16048,N_14648,N_14228);
and U16049 (N_16049,N_13680,N_14694);
nand U16050 (N_16050,N_13841,N_14983);
or U16051 (N_16051,N_14271,N_14699);
xor U16052 (N_16052,N_14213,N_12774);
nor U16053 (N_16053,N_14350,N_14137);
xnor U16054 (N_16054,N_13364,N_14162);
or U16055 (N_16055,N_14634,N_14661);
nor U16056 (N_16056,N_12978,N_14779);
or U16057 (N_16057,N_12966,N_14270);
nor U16058 (N_16058,N_13788,N_14081);
nand U16059 (N_16059,N_14100,N_13851);
xor U16060 (N_16060,N_14393,N_14326);
xor U16061 (N_16061,N_13160,N_12994);
and U16062 (N_16062,N_13973,N_13997);
or U16063 (N_16063,N_13894,N_13497);
and U16064 (N_16064,N_13703,N_12815);
nand U16065 (N_16065,N_13823,N_12788);
xnor U16066 (N_16066,N_12642,N_12693);
or U16067 (N_16067,N_14781,N_13515);
nor U16068 (N_16068,N_13683,N_13812);
nand U16069 (N_16069,N_14571,N_13028);
nor U16070 (N_16070,N_13868,N_13178);
or U16071 (N_16071,N_13410,N_13276);
or U16072 (N_16072,N_13200,N_13345);
or U16073 (N_16073,N_12658,N_14401);
or U16074 (N_16074,N_12740,N_13493);
nor U16075 (N_16075,N_13291,N_14436);
xnor U16076 (N_16076,N_13335,N_14341);
and U16077 (N_16077,N_13240,N_13610);
nor U16078 (N_16078,N_12972,N_14765);
nor U16079 (N_16079,N_13429,N_14584);
and U16080 (N_16080,N_13528,N_14886);
nand U16081 (N_16081,N_14546,N_14397);
and U16082 (N_16082,N_13673,N_12822);
nand U16083 (N_16083,N_14113,N_14556);
xnor U16084 (N_16084,N_12885,N_13386);
and U16085 (N_16085,N_14711,N_13798);
or U16086 (N_16086,N_14842,N_13068);
xnor U16087 (N_16087,N_12529,N_14261);
nor U16088 (N_16088,N_13039,N_13438);
nand U16089 (N_16089,N_14335,N_14740);
or U16090 (N_16090,N_13389,N_14407);
xnor U16091 (N_16091,N_13545,N_14688);
and U16092 (N_16092,N_13369,N_14766);
nor U16093 (N_16093,N_12510,N_13328);
or U16094 (N_16094,N_14211,N_13241);
or U16095 (N_16095,N_13450,N_12831);
or U16096 (N_16096,N_13557,N_14822);
nand U16097 (N_16097,N_14351,N_13129);
xnor U16098 (N_16098,N_14001,N_14741);
or U16099 (N_16099,N_13061,N_13199);
and U16100 (N_16100,N_12981,N_12573);
or U16101 (N_16101,N_14037,N_14675);
nor U16102 (N_16102,N_13148,N_13277);
or U16103 (N_16103,N_13985,N_13781);
or U16104 (N_16104,N_14405,N_13777);
nor U16105 (N_16105,N_12814,N_13081);
or U16106 (N_16106,N_14265,N_13829);
or U16107 (N_16107,N_13076,N_12541);
and U16108 (N_16108,N_14134,N_14938);
nand U16109 (N_16109,N_13135,N_13650);
nand U16110 (N_16110,N_13534,N_13036);
and U16111 (N_16111,N_14524,N_14169);
or U16112 (N_16112,N_12565,N_14536);
xor U16113 (N_16113,N_12946,N_13696);
nand U16114 (N_16114,N_14076,N_12597);
nand U16115 (N_16115,N_12734,N_14754);
nand U16116 (N_16116,N_14630,N_13899);
nand U16117 (N_16117,N_14175,N_12741);
or U16118 (N_16118,N_14202,N_14486);
or U16119 (N_16119,N_14849,N_12976);
nand U16120 (N_16120,N_13578,N_14460);
xor U16121 (N_16121,N_12581,N_14621);
nor U16122 (N_16122,N_13669,N_13734);
and U16123 (N_16123,N_14512,N_14907);
or U16124 (N_16124,N_12971,N_14848);
xnor U16125 (N_16125,N_14920,N_13863);
nand U16126 (N_16126,N_14243,N_14286);
and U16127 (N_16127,N_12600,N_14071);
and U16128 (N_16128,N_14135,N_13838);
nand U16129 (N_16129,N_12974,N_13558);
or U16130 (N_16130,N_14564,N_13293);
or U16131 (N_16131,N_12598,N_14558);
and U16132 (N_16132,N_12747,N_13431);
xor U16133 (N_16133,N_14324,N_12695);
or U16134 (N_16134,N_13888,N_13914);
nand U16135 (N_16135,N_13846,N_14253);
xnor U16136 (N_16136,N_13598,N_14832);
or U16137 (N_16137,N_14328,N_12587);
nand U16138 (N_16138,N_14233,N_12835);
and U16139 (N_16139,N_14127,N_13903);
and U16140 (N_16140,N_12660,N_13174);
xnor U16141 (N_16141,N_13223,N_14289);
nand U16142 (N_16142,N_13658,N_14429);
nor U16143 (N_16143,N_14010,N_13691);
nand U16144 (N_16144,N_14614,N_14830);
or U16145 (N_16145,N_12744,N_13176);
nor U16146 (N_16146,N_14297,N_14954);
and U16147 (N_16147,N_13507,N_14227);
and U16148 (N_16148,N_12605,N_12684);
nor U16149 (N_16149,N_14123,N_13275);
or U16150 (N_16150,N_12579,N_13471);
or U16151 (N_16151,N_13248,N_14843);
nor U16152 (N_16152,N_13898,N_13079);
nor U16153 (N_16153,N_12908,N_14024);
nor U16154 (N_16154,N_12732,N_14093);
and U16155 (N_16155,N_13808,N_12719);
nand U16156 (N_16156,N_14394,N_13307);
xnor U16157 (N_16157,N_14141,N_13501);
nor U16158 (N_16158,N_12846,N_13522);
and U16159 (N_16159,N_14763,N_12558);
nand U16160 (N_16160,N_14816,N_13215);
and U16161 (N_16161,N_13260,N_13595);
xor U16162 (N_16162,N_14493,N_13953);
or U16163 (N_16163,N_12724,N_12901);
and U16164 (N_16164,N_12980,N_13922);
and U16165 (N_16165,N_13516,N_13704);
nor U16166 (N_16166,N_14642,N_13621);
nor U16167 (N_16167,N_13599,N_14296);
nor U16168 (N_16168,N_13857,N_13601);
xnor U16169 (N_16169,N_14865,N_13398);
or U16170 (N_16170,N_13935,N_13852);
nand U16171 (N_16171,N_14624,N_12943);
or U16172 (N_16172,N_13580,N_13114);
and U16173 (N_16173,N_13479,N_13842);
nor U16174 (N_16174,N_14044,N_14996);
nand U16175 (N_16175,N_14026,N_12963);
xnor U16176 (N_16176,N_14598,N_14980);
xor U16177 (N_16177,N_14441,N_14267);
nand U16178 (N_16178,N_14095,N_14206);
and U16179 (N_16179,N_14691,N_12965);
nor U16180 (N_16180,N_14342,N_13203);
nor U16181 (N_16181,N_13375,N_13817);
nor U16182 (N_16182,N_14380,N_12952);
xor U16183 (N_16183,N_13958,N_14142);
nor U16184 (N_16184,N_12792,N_12601);
and U16185 (N_16185,N_13370,N_13171);
nand U16186 (N_16186,N_12761,N_13511);
nand U16187 (N_16187,N_14732,N_12805);
nand U16188 (N_16188,N_13103,N_12749);
xnor U16189 (N_16189,N_14541,N_14795);
or U16190 (N_16190,N_14817,N_12629);
or U16191 (N_16191,N_14117,N_13606);
xor U16192 (N_16192,N_14941,N_14906);
and U16193 (N_16193,N_13002,N_13188);
xnor U16194 (N_16194,N_12880,N_13091);
nor U16195 (N_16195,N_13642,N_12949);
nor U16196 (N_16196,N_14755,N_13924);
and U16197 (N_16197,N_14602,N_13523);
nand U16198 (N_16198,N_13436,N_13732);
nand U16199 (N_16199,N_12622,N_12704);
nand U16200 (N_16200,N_14176,N_13024);
xor U16201 (N_16201,N_13556,N_13082);
nand U16202 (N_16202,N_13427,N_12570);
xor U16203 (N_16203,N_14269,N_12667);
nand U16204 (N_16204,N_14362,N_12945);
or U16205 (N_16205,N_14813,N_14238);
nand U16206 (N_16206,N_13994,N_14620);
nand U16207 (N_16207,N_13988,N_13672);
nand U16208 (N_16208,N_13154,N_14049);
and U16209 (N_16209,N_12645,N_14969);
and U16210 (N_16210,N_12969,N_14033);
nand U16211 (N_16211,N_14669,N_14096);
xnor U16212 (N_16212,N_13118,N_14245);
and U16213 (N_16213,N_14188,N_14451);
nand U16214 (N_16214,N_12577,N_14450);
and U16215 (N_16215,N_13298,N_14003);
nor U16216 (N_16216,N_14039,N_13529);
and U16217 (N_16217,N_14948,N_13925);
xor U16218 (N_16218,N_14459,N_14210);
nand U16219 (N_16219,N_13527,N_14572);
nor U16220 (N_16220,N_14276,N_14012);
xnor U16221 (N_16221,N_14389,N_13797);
nor U16222 (N_16222,N_13646,N_12872);
or U16223 (N_16223,N_12592,N_14932);
or U16224 (N_16224,N_14016,N_14410);
and U16225 (N_16225,N_14354,N_12961);
or U16226 (N_16226,N_13467,N_13624);
and U16227 (N_16227,N_14775,N_14386);
and U16228 (N_16228,N_14573,N_13776);
nor U16229 (N_16229,N_13521,N_12906);
and U16230 (N_16230,N_14086,N_13713);
or U16231 (N_16231,N_12559,N_13968);
nor U16232 (N_16232,N_14981,N_13332);
and U16233 (N_16233,N_12709,N_14662);
nand U16234 (N_16234,N_13686,N_12786);
or U16235 (N_16235,N_14221,N_14519);
and U16236 (N_16236,N_13916,N_13768);
nand U16237 (N_16237,N_14274,N_12727);
nand U16238 (N_16238,N_13719,N_12794);
nand U16239 (N_16239,N_12785,N_12875);
and U16240 (N_16240,N_13636,N_12569);
nand U16241 (N_16241,N_13639,N_13745);
and U16242 (N_16242,N_13874,N_12534);
or U16243 (N_16243,N_13349,N_14284);
or U16244 (N_16244,N_12531,N_13220);
nand U16245 (N_16245,N_13756,N_14009);
xnor U16246 (N_16246,N_14916,N_14821);
nor U16247 (N_16247,N_14592,N_14656);
nor U16248 (N_16248,N_13551,N_14425);
nand U16249 (N_16249,N_12919,N_13641);
xor U16250 (N_16250,N_14863,N_14852);
xnor U16251 (N_16251,N_14912,N_13892);
nand U16252 (N_16252,N_13589,N_14456);
and U16253 (N_16253,N_14289,N_14473);
nand U16254 (N_16254,N_13158,N_14258);
nor U16255 (N_16255,N_13552,N_14309);
xor U16256 (N_16256,N_12936,N_13309);
and U16257 (N_16257,N_13664,N_13997);
or U16258 (N_16258,N_12702,N_12916);
and U16259 (N_16259,N_14636,N_12700);
and U16260 (N_16260,N_14917,N_14623);
nand U16261 (N_16261,N_13762,N_13045);
nor U16262 (N_16262,N_14022,N_12772);
xor U16263 (N_16263,N_12622,N_14567);
or U16264 (N_16264,N_12727,N_12856);
or U16265 (N_16265,N_12812,N_13140);
nor U16266 (N_16266,N_12894,N_12732);
and U16267 (N_16267,N_13972,N_12892);
xor U16268 (N_16268,N_12963,N_13662);
xnor U16269 (N_16269,N_13362,N_14318);
and U16270 (N_16270,N_12594,N_13080);
xnor U16271 (N_16271,N_13626,N_13766);
xor U16272 (N_16272,N_14799,N_13464);
nor U16273 (N_16273,N_14125,N_14313);
or U16274 (N_16274,N_14310,N_13196);
nor U16275 (N_16275,N_14304,N_12607);
and U16276 (N_16276,N_12573,N_14310);
or U16277 (N_16277,N_14943,N_14500);
and U16278 (N_16278,N_14310,N_13647);
nand U16279 (N_16279,N_13548,N_14113);
xor U16280 (N_16280,N_12621,N_13273);
and U16281 (N_16281,N_13173,N_13374);
nor U16282 (N_16282,N_14952,N_14797);
xor U16283 (N_16283,N_14683,N_12832);
xor U16284 (N_16284,N_14683,N_13059);
or U16285 (N_16285,N_13785,N_13478);
and U16286 (N_16286,N_13247,N_14517);
and U16287 (N_16287,N_14576,N_13732);
and U16288 (N_16288,N_13630,N_13555);
nand U16289 (N_16289,N_14527,N_12591);
and U16290 (N_16290,N_14187,N_14043);
xor U16291 (N_16291,N_14776,N_14866);
xnor U16292 (N_16292,N_14609,N_14768);
xnor U16293 (N_16293,N_13639,N_13481);
nor U16294 (N_16294,N_14335,N_13942);
or U16295 (N_16295,N_13388,N_13763);
nand U16296 (N_16296,N_14474,N_14054);
and U16297 (N_16297,N_13718,N_14814);
nor U16298 (N_16298,N_14560,N_14266);
or U16299 (N_16299,N_13026,N_14846);
nand U16300 (N_16300,N_13384,N_13082);
nor U16301 (N_16301,N_13766,N_14347);
nand U16302 (N_16302,N_14935,N_14017);
nor U16303 (N_16303,N_12653,N_12690);
nor U16304 (N_16304,N_14978,N_13773);
xnor U16305 (N_16305,N_12805,N_14148);
xor U16306 (N_16306,N_12892,N_12650);
xnor U16307 (N_16307,N_14751,N_14334);
xor U16308 (N_16308,N_13160,N_14775);
or U16309 (N_16309,N_14127,N_14935);
nor U16310 (N_16310,N_14881,N_14430);
or U16311 (N_16311,N_12862,N_14591);
nand U16312 (N_16312,N_14364,N_13446);
nor U16313 (N_16313,N_13989,N_13361);
nor U16314 (N_16314,N_13227,N_14627);
and U16315 (N_16315,N_13628,N_14273);
or U16316 (N_16316,N_14855,N_14254);
or U16317 (N_16317,N_14519,N_13726);
nor U16318 (N_16318,N_14189,N_13475);
xor U16319 (N_16319,N_12872,N_12741);
xor U16320 (N_16320,N_14309,N_13894);
or U16321 (N_16321,N_13495,N_14253);
or U16322 (N_16322,N_13170,N_14803);
or U16323 (N_16323,N_14804,N_14394);
or U16324 (N_16324,N_14111,N_12860);
or U16325 (N_16325,N_13928,N_12524);
nor U16326 (N_16326,N_14811,N_12970);
or U16327 (N_16327,N_14255,N_13010);
xnor U16328 (N_16328,N_13185,N_12644);
xor U16329 (N_16329,N_13780,N_14791);
and U16330 (N_16330,N_14757,N_13092);
xnor U16331 (N_16331,N_13170,N_13430);
nor U16332 (N_16332,N_12534,N_13701);
or U16333 (N_16333,N_14018,N_14897);
and U16334 (N_16334,N_12641,N_13465);
xor U16335 (N_16335,N_14189,N_12653);
and U16336 (N_16336,N_13097,N_14958);
and U16337 (N_16337,N_13455,N_13663);
or U16338 (N_16338,N_13058,N_12937);
or U16339 (N_16339,N_12696,N_13255);
or U16340 (N_16340,N_13424,N_14557);
nor U16341 (N_16341,N_13881,N_12717);
nand U16342 (N_16342,N_12637,N_13069);
nand U16343 (N_16343,N_13770,N_12677);
nor U16344 (N_16344,N_13118,N_12883);
xor U16345 (N_16345,N_12906,N_13569);
or U16346 (N_16346,N_13625,N_14034);
xor U16347 (N_16347,N_13830,N_12659);
nor U16348 (N_16348,N_12947,N_14595);
and U16349 (N_16349,N_14602,N_13565);
nand U16350 (N_16350,N_14983,N_14172);
and U16351 (N_16351,N_14675,N_14875);
nor U16352 (N_16352,N_14487,N_13119);
nand U16353 (N_16353,N_13595,N_13145);
xnor U16354 (N_16354,N_14472,N_12612);
nand U16355 (N_16355,N_14543,N_12715);
xnor U16356 (N_16356,N_14736,N_14892);
or U16357 (N_16357,N_13737,N_14274);
and U16358 (N_16358,N_13044,N_14976);
and U16359 (N_16359,N_12755,N_13449);
xnor U16360 (N_16360,N_13931,N_14060);
xnor U16361 (N_16361,N_14956,N_12765);
and U16362 (N_16362,N_13122,N_14652);
xor U16363 (N_16363,N_12679,N_13845);
and U16364 (N_16364,N_14843,N_12571);
nand U16365 (N_16365,N_12739,N_14035);
or U16366 (N_16366,N_13407,N_14247);
xor U16367 (N_16367,N_14688,N_13987);
nor U16368 (N_16368,N_14428,N_14029);
or U16369 (N_16369,N_12601,N_13671);
nand U16370 (N_16370,N_13472,N_14045);
and U16371 (N_16371,N_14116,N_14367);
xnor U16372 (N_16372,N_14031,N_14422);
and U16373 (N_16373,N_13772,N_14914);
or U16374 (N_16374,N_13654,N_12624);
nand U16375 (N_16375,N_12933,N_14242);
and U16376 (N_16376,N_13931,N_14488);
xor U16377 (N_16377,N_14913,N_14891);
xor U16378 (N_16378,N_14562,N_12669);
nand U16379 (N_16379,N_12655,N_13519);
nand U16380 (N_16380,N_14512,N_13833);
and U16381 (N_16381,N_13550,N_12547);
nand U16382 (N_16382,N_12839,N_13574);
xor U16383 (N_16383,N_12821,N_12881);
and U16384 (N_16384,N_12564,N_14145);
nand U16385 (N_16385,N_13262,N_13278);
nand U16386 (N_16386,N_12909,N_13261);
xnor U16387 (N_16387,N_14119,N_12902);
and U16388 (N_16388,N_13821,N_14024);
or U16389 (N_16389,N_13694,N_12724);
nor U16390 (N_16390,N_13852,N_13942);
nor U16391 (N_16391,N_12722,N_13816);
or U16392 (N_16392,N_12516,N_13875);
and U16393 (N_16393,N_14460,N_12922);
or U16394 (N_16394,N_14979,N_14495);
xor U16395 (N_16395,N_14401,N_14986);
or U16396 (N_16396,N_14175,N_12781);
nand U16397 (N_16397,N_14464,N_14605);
xor U16398 (N_16398,N_13495,N_14907);
nand U16399 (N_16399,N_12597,N_14164);
xor U16400 (N_16400,N_12629,N_12898);
xor U16401 (N_16401,N_14088,N_13673);
and U16402 (N_16402,N_12566,N_14494);
or U16403 (N_16403,N_12895,N_14169);
nand U16404 (N_16404,N_13295,N_13443);
and U16405 (N_16405,N_14171,N_14563);
nor U16406 (N_16406,N_12928,N_14294);
nand U16407 (N_16407,N_13615,N_12971);
xnor U16408 (N_16408,N_13478,N_13719);
nand U16409 (N_16409,N_13933,N_13333);
nor U16410 (N_16410,N_14991,N_13027);
nor U16411 (N_16411,N_13916,N_14612);
nor U16412 (N_16412,N_14185,N_14560);
nor U16413 (N_16413,N_13797,N_14171);
xnor U16414 (N_16414,N_13090,N_13105);
nand U16415 (N_16415,N_13549,N_13184);
xnor U16416 (N_16416,N_14381,N_14948);
nand U16417 (N_16417,N_13674,N_14713);
nand U16418 (N_16418,N_14185,N_14491);
and U16419 (N_16419,N_13829,N_13428);
nor U16420 (N_16420,N_14584,N_13740);
nand U16421 (N_16421,N_13204,N_13282);
or U16422 (N_16422,N_12831,N_14984);
nor U16423 (N_16423,N_12571,N_13545);
xor U16424 (N_16424,N_12771,N_14052);
or U16425 (N_16425,N_12988,N_12631);
and U16426 (N_16426,N_14282,N_13742);
or U16427 (N_16427,N_14974,N_14039);
nand U16428 (N_16428,N_14345,N_14361);
xor U16429 (N_16429,N_13466,N_12601);
nor U16430 (N_16430,N_13911,N_13217);
and U16431 (N_16431,N_14910,N_14307);
nand U16432 (N_16432,N_13603,N_14263);
or U16433 (N_16433,N_14072,N_13166);
nor U16434 (N_16434,N_13515,N_13987);
and U16435 (N_16435,N_14308,N_14482);
and U16436 (N_16436,N_14830,N_14691);
nor U16437 (N_16437,N_13470,N_12582);
nand U16438 (N_16438,N_14913,N_14601);
and U16439 (N_16439,N_12874,N_12762);
and U16440 (N_16440,N_14807,N_12891);
nand U16441 (N_16441,N_13020,N_13273);
xnor U16442 (N_16442,N_14167,N_14183);
nor U16443 (N_16443,N_14942,N_13912);
nand U16444 (N_16444,N_14543,N_13822);
nor U16445 (N_16445,N_13859,N_12885);
xor U16446 (N_16446,N_14794,N_13800);
and U16447 (N_16447,N_13901,N_14581);
nand U16448 (N_16448,N_13950,N_13633);
and U16449 (N_16449,N_14413,N_14201);
nor U16450 (N_16450,N_14427,N_14760);
and U16451 (N_16451,N_14241,N_13303);
and U16452 (N_16452,N_13286,N_14328);
and U16453 (N_16453,N_14285,N_14932);
xnor U16454 (N_16454,N_13016,N_12809);
nor U16455 (N_16455,N_13458,N_13225);
and U16456 (N_16456,N_12979,N_13129);
xor U16457 (N_16457,N_14959,N_12995);
xor U16458 (N_16458,N_13645,N_14743);
nand U16459 (N_16459,N_14948,N_13693);
nand U16460 (N_16460,N_13342,N_13212);
or U16461 (N_16461,N_13525,N_14697);
xnor U16462 (N_16462,N_12663,N_13209);
or U16463 (N_16463,N_12766,N_13819);
and U16464 (N_16464,N_13205,N_13127);
nand U16465 (N_16465,N_13971,N_13638);
xnor U16466 (N_16466,N_14221,N_13638);
xor U16467 (N_16467,N_12799,N_13657);
or U16468 (N_16468,N_13120,N_12503);
nor U16469 (N_16469,N_14592,N_13324);
or U16470 (N_16470,N_14897,N_13035);
nand U16471 (N_16471,N_14788,N_13444);
nand U16472 (N_16472,N_13855,N_13642);
nand U16473 (N_16473,N_14805,N_14107);
nor U16474 (N_16474,N_13643,N_13012);
and U16475 (N_16475,N_14832,N_13647);
nor U16476 (N_16476,N_14434,N_12779);
nor U16477 (N_16477,N_12782,N_13956);
or U16478 (N_16478,N_14514,N_13752);
nor U16479 (N_16479,N_12707,N_12760);
xnor U16480 (N_16480,N_12525,N_14706);
nor U16481 (N_16481,N_13818,N_13959);
nor U16482 (N_16482,N_13886,N_14279);
xnor U16483 (N_16483,N_13297,N_13770);
nor U16484 (N_16484,N_14552,N_14539);
xnor U16485 (N_16485,N_13633,N_13427);
or U16486 (N_16486,N_13536,N_12597);
nand U16487 (N_16487,N_12926,N_13050);
nand U16488 (N_16488,N_13543,N_14068);
xnor U16489 (N_16489,N_13164,N_13989);
and U16490 (N_16490,N_14447,N_14665);
or U16491 (N_16491,N_13168,N_12741);
and U16492 (N_16492,N_14743,N_13506);
or U16493 (N_16493,N_13083,N_12727);
or U16494 (N_16494,N_12979,N_13750);
nor U16495 (N_16495,N_14707,N_12884);
or U16496 (N_16496,N_13452,N_14305);
and U16497 (N_16497,N_14437,N_14847);
and U16498 (N_16498,N_14279,N_14582);
or U16499 (N_16499,N_12866,N_14139);
or U16500 (N_16500,N_14763,N_13049);
and U16501 (N_16501,N_13222,N_13597);
and U16502 (N_16502,N_13746,N_12628);
and U16503 (N_16503,N_12622,N_14000);
xor U16504 (N_16504,N_14844,N_14149);
nand U16505 (N_16505,N_13365,N_13880);
xnor U16506 (N_16506,N_13206,N_14103);
and U16507 (N_16507,N_13338,N_13208);
nand U16508 (N_16508,N_14870,N_12863);
or U16509 (N_16509,N_14865,N_14599);
or U16510 (N_16510,N_14408,N_13175);
nor U16511 (N_16511,N_12758,N_14803);
nor U16512 (N_16512,N_13910,N_13904);
or U16513 (N_16513,N_14799,N_13728);
or U16514 (N_16514,N_13500,N_14942);
nor U16515 (N_16515,N_14904,N_12707);
or U16516 (N_16516,N_14915,N_13881);
xnor U16517 (N_16517,N_14795,N_14867);
and U16518 (N_16518,N_13628,N_13605);
and U16519 (N_16519,N_13833,N_12987);
or U16520 (N_16520,N_12606,N_12560);
or U16521 (N_16521,N_14097,N_14939);
nor U16522 (N_16522,N_13127,N_13352);
nor U16523 (N_16523,N_14338,N_13375);
nand U16524 (N_16524,N_13792,N_12954);
xnor U16525 (N_16525,N_13635,N_13893);
nor U16526 (N_16526,N_14438,N_14587);
nand U16527 (N_16527,N_14486,N_12953);
or U16528 (N_16528,N_13625,N_13283);
nand U16529 (N_16529,N_13500,N_14191);
nand U16530 (N_16530,N_13243,N_13902);
or U16531 (N_16531,N_13810,N_12988);
or U16532 (N_16532,N_13020,N_13763);
or U16533 (N_16533,N_14555,N_14308);
and U16534 (N_16534,N_12571,N_13009);
xnor U16535 (N_16535,N_12668,N_14716);
and U16536 (N_16536,N_14804,N_14726);
or U16537 (N_16537,N_13809,N_14965);
nor U16538 (N_16538,N_14402,N_12928);
xnor U16539 (N_16539,N_12600,N_12993);
nand U16540 (N_16540,N_13846,N_12624);
nor U16541 (N_16541,N_12979,N_12960);
nand U16542 (N_16542,N_12706,N_12724);
and U16543 (N_16543,N_12967,N_14837);
nor U16544 (N_16544,N_14233,N_13129);
and U16545 (N_16545,N_12924,N_12510);
nand U16546 (N_16546,N_14739,N_14852);
nand U16547 (N_16547,N_13309,N_14351);
and U16548 (N_16548,N_14271,N_14464);
or U16549 (N_16549,N_14365,N_14210);
or U16550 (N_16550,N_13334,N_12883);
xor U16551 (N_16551,N_12901,N_14283);
nor U16552 (N_16552,N_13123,N_12609);
or U16553 (N_16553,N_12685,N_13928);
or U16554 (N_16554,N_14024,N_14263);
nand U16555 (N_16555,N_14133,N_13313);
nand U16556 (N_16556,N_14516,N_14597);
nand U16557 (N_16557,N_13685,N_14686);
nor U16558 (N_16558,N_13456,N_14265);
xor U16559 (N_16559,N_12533,N_14010);
xor U16560 (N_16560,N_13632,N_13518);
and U16561 (N_16561,N_12649,N_12663);
and U16562 (N_16562,N_13412,N_14580);
nand U16563 (N_16563,N_14146,N_14746);
or U16564 (N_16564,N_12531,N_14097);
xnor U16565 (N_16565,N_14330,N_14805);
xnor U16566 (N_16566,N_12527,N_12517);
nand U16567 (N_16567,N_12818,N_13763);
and U16568 (N_16568,N_12556,N_14038);
nand U16569 (N_16569,N_14134,N_12941);
and U16570 (N_16570,N_12720,N_13137);
and U16571 (N_16571,N_14270,N_14600);
nor U16572 (N_16572,N_13580,N_12698);
or U16573 (N_16573,N_13240,N_14395);
xnor U16574 (N_16574,N_14397,N_12758);
and U16575 (N_16575,N_12570,N_12792);
nand U16576 (N_16576,N_14106,N_13661);
nand U16577 (N_16577,N_12545,N_13337);
or U16578 (N_16578,N_14450,N_12554);
and U16579 (N_16579,N_13520,N_13164);
nand U16580 (N_16580,N_14491,N_13888);
nor U16581 (N_16581,N_12730,N_12818);
xor U16582 (N_16582,N_13253,N_12628);
nand U16583 (N_16583,N_12646,N_13298);
xnor U16584 (N_16584,N_12512,N_13499);
xor U16585 (N_16585,N_13000,N_14853);
nand U16586 (N_16586,N_13792,N_13972);
nor U16587 (N_16587,N_13295,N_13544);
nand U16588 (N_16588,N_12619,N_12773);
and U16589 (N_16589,N_14170,N_14634);
or U16590 (N_16590,N_14827,N_13307);
nand U16591 (N_16591,N_12533,N_13923);
nor U16592 (N_16592,N_13825,N_12521);
xor U16593 (N_16593,N_13071,N_14699);
xor U16594 (N_16594,N_13237,N_13505);
nand U16595 (N_16595,N_13533,N_13309);
and U16596 (N_16596,N_12864,N_14946);
or U16597 (N_16597,N_14146,N_13897);
or U16598 (N_16598,N_14030,N_12659);
or U16599 (N_16599,N_14756,N_13279);
xor U16600 (N_16600,N_12546,N_12621);
and U16601 (N_16601,N_14590,N_12597);
and U16602 (N_16602,N_13859,N_13536);
and U16603 (N_16603,N_13024,N_14731);
nor U16604 (N_16604,N_14614,N_13012);
nand U16605 (N_16605,N_14792,N_14287);
xor U16606 (N_16606,N_14112,N_14253);
and U16607 (N_16607,N_13361,N_13462);
xnor U16608 (N_16608,N_12762,N_14916);
and U16609 (N_16609,N_14522,N_13230);
or U16610 (N_16610,N_13601,N_12665);
nand U16611 (N_16611,N_12561,N_13393);
and U16612 (N_16612,N_14291,N_14209);
or U16613 (N_16613,N_14534,N_14676);
xor U16614 (N_16614,N_12637,N_14107);
or U16615 (N_16615,N_14503,N_13199);
or U16616 (N_16616,N_14756,N_12937);
or U16617 (N_16617,N_14279,N_14435);
nor U16618 (N_16618,N_14635,N_12744);
nand U16619 (N_16619,N_12505,N_12503);
and U16620 (N_16620,N_12769,N_13450);
nand U16621 (N_16621,N_14462,N_13674);
nand U16622 (N_16622,N_13289,N_13332);
and U16623 (N_16623,N_13949,N_12753);
or U16624 (N_16624,N_12849,N_14295);
and U16625 (N_16625,N_14884,N_13044);
nand U16626 (N_16626,N_13384,N_14793);
nor U16627 (N_16627,N_13080,N_14846);
nand U16628 (N_16628,N_14013,N_12673);
xnor U16629 (N_16629,N_13025,N_14242);
nor U16630 (N_16630,N_14183,N_14401);
xor U16631 (N_16631,N_14577,N_14594);
nor U16632 (N_16632,N_13307,N_12614);
and U16633 (N_16633,N_14505,N_12888);
and U16634 (N_16634,N_12650,N_14350);
and U16635 (N_16635,N_14232,N_14472);
and U16636 (N_16636,N_12786,N_14652);
or U16637 (N_16637,N_14055,N_13307);
nand U16638 (N_16638,N_14389,N_13381);
and U16639 (N_16639,N_12895,N_13456);
or U16640 (N_16640,N_12509,N_13489);
or U16641 (N_16641,N_12636,N_12799);
xnor U16642 (N_16642,N_14915,N_14142);
xnor U16643 (N_16643,N_12912,N_13982);
nor U16644 (N_16644,N_14165,N_14764);
nand U16645 (N_16645,N_12699,N_13940);
xor U16646 (N_16646,N_13992,N_14198);
or U16647 (N_16647,N_13010,N_13260);
and U16648 (N_16648,N_13986,N_13300);
or U16649 (N_16649,N_13688,N_14767);
nand U16650 (N_16650,N_14188,N_14323);
xor U16651 (N_16651,N_13421,N_14082);
nand U16652 (N_16652,N_14612,N_13882);
nand U16653 (N_16653,N_13303,N_13943);
or U16654 (N_16654,N_12900,N_14759);
nor U16655 (N_16655,N_12914,N_14644);
and U16656 (N_16656,N_14009,N_14151);
nor U16657 (N_16657,N_13803,N_13869);
xnor U16658 (N_16658,N_13792,N_13822);
or U16659 (N_16659,N_13466,N_14026);
xnor U16660 (N_16660,N_13308,N_12584);
or U16661 (N_16661,N_14723,N_13125);
or U16662 (N_16662,N_12790,N_12969);
nand U16663 (N_16663,N_12789,N_12656);
xor U16664 (N_16664,N_14170,N_14520);
and U16665 (N_16665,N_14955,N_13482);
and U16666 (N_16666,N_14691,N_14106);
or U16667 (N_16667,N_14026,N_13949);
nor U16668 (N_16668,N_12931,N_13402);
or U16669 (N_16669,N_13249,N_14589);
and U16670 (N_16670,N_14274,N_14490);
nand U16671 (N_16671,N_14114,N_14807);
and U16672 (N_16672,N_13043,N_13969);
nor U16673 (N_16673,N_13901,N_13664);
nand U16674 (N_16674,N_13398,N_13182);
or U16675 (N_16675,N_13848,N_12838);
nand U16676 (N_16676,N_13714,N_13530);
nor U16677 (N_16677,N_14694,N_12659);
nor U16678 (N_16678,N_12688,N_13137);
or U16679 (N_16679,N_12700,N_14974);
xnor U16680 (N_16680,N_12814,N_13576);
or U16681 (N_16681,N_12796,N_13004);
and U16682 (N_16682,N_14846,N_14198);
nand U16683 (N_16683,N_13053,N_12916);
nor U16684 (N_16684,N_13992,N_14426);
or U16685 (N_16685,N_12504,N_13131);
nand U16686 (N_16686,N_14300,N_12864);
and U16687 (N_16687,N_14227,N_12650);
nor U16688 (N_16688,N_13087,N_14566);
xnor U16689 (N_16689,N_14491,N_12611);
xor U16690 (N_16690,N_13825,N_13786);
or U16691 (N_16691,N_13130,N_13186);
xnor U16692 (N_16692,N_14367,N_13101);
nand U16693 (N_16693,N_14056,N_12913);
nor U16694 (N_16694,N_13662,N_12925);
and U16695 (N_16695,N_13921,N_14438);
nor U16696 (N_16696,N_14258,N_13656);
and U16697 (N_16697,N_13332,N_14988);
or U16698 (N_16698,N_14894,N_13129);
and U16699 (N_16699,N_14252,N_14294);
and U16700 (N_16700,N_13589,N_13424);
nor U16701 (N_16701,N_13938,N_13176);
or U16702 (N_16702,N_13298,N_12954);
nor U16703 (N_16703,N_14622,N_13631);
and U16704 (N_16704,N_13064,N_13451);
nand U16705 (N_16705,N_13290,N_14083);
and U16706 (N_16706,N_14910,N_14435);
nand U16707 (N_16707,N_13897,N_14778);
nand U16708 (N_16708,N_12690,N_13405);
nand U16709 (N_16709,N_12756,N_13248);
nand U16710 (N_16710,N_13629,N_14543);
nand U16711 (N_16711,N_14209,N_13914);
xnor U16712 (N_16712,N_13256,N_14402);
and U16713 (N_16713,N_12940,N_13897);
or U16714 (N_16714,N_13627,N_13619);
nor U16715 (N_16715,N_14558,N_13195);
xnor U16716 (N_16716,N_13913,N_13269);
nor U16717 (N_16717,N_13436,N_13304);
xnor U16718 (N_16718,N_14278,N_14050);
nand U16719 (N_16719,N_13211,N_13673);
and U16720 (N_16720,N_14341,N_12673);
xnor U16721 (N_16721,N_12986,N_14032);
or U16722 (N_16722,N_13807,N_13119);
nand U16723 (N_16723,N_14416,N_14510);
and U16724 (N_16724,N_14570,N_14894);
or U16725 (N_16725,N_13236,N_12781);
nor U16726 (N_16726,N_14603,N_12748);
xor U16727 (N_16727,N_14624,N_14265);
nor U16728 (N_16728,N_13613,N_13178);
or U16729 (N_16729,N_12611,N_14038);
nor U16730 (N_16730,N_13237,N_12929);
nand U16731 (N_16731,N_13761,N_14507);
nor U16732 (N_16732,N_12879,N_12505);
nor U16733 (N_16733,N_14156,N_12824);
nand U16734 (N_16734,N_12736,N_12787);
or U16735 (N_16735,N_13203,N_13579);
or U16736 (N_16736,N_13601,N_14765);
nor U16737 (N_16737,N_12910,N_13532);
nand U16738 (N_16738,N_13994,N_14215);
and U16739 (N_16739,N_14385,N_14875);
nand U16740 (N_16740,N_12885,N_14128);
xor U16741 (N_16741,N_13352,N_13514);
nand U16742 (N_16742,N_13949,N_14579);
nor U16743 (N_16743,N_13176,N_14050);
and U16744 (N_16744,N_13200,N_13911);
nand U16745 (N_16745,N_14443,N_12759);
nand U16746 (N_16746,N_14705,N_12790);
nor U16747 (N_16747,N_13851,N_12566);
nor U16748 (N_16748,N_14047,N_12692);
or U16749 (N_16749,N_13306,N_13273);
and U16750 (N_16750,N_13533,N_13911);
xnor U16751 (N_16751,N_14048,N_14747);
nor U16752 (N_16752,N_12918,N_13165);
nand U16753 (N_16753,N_12772,N_13889);
and U16754 (N_16754,N_14419,N_14601);
nor U16755 (N_16755,N_13522,N_12973);
or U16756 (N_16756,N_13462,N_13623);
or U16757 (N_16757,N_13029,N_13931);
nand U16758 (N_16758,N_14414,N_14475);
or U16759 (N_16759,N_14584,N_12792);
nand U16760 (N_16760,N_13910,N_12752);
and U16761 (N_16761,N_13279,N_13689);
and U16762 (N_16762,N_14214,N_14628);
nand U16763 (N_16763,N_13219,N_13860);
xor U16764 (N_16764,N_14085,N_12873);
nor U16765 (N_16765,N_14988,N_13280);
nand U16766 (N_16766,N_13490,N_13678);
xnor U16767 (N_16767,N_14710,N_12810);
nor U16768 (N_16768,N_13666,N_14036);
or U16769 (N_16769,N_14279,N_14237);
nor U16770 (N_16770,N_13311,N_14793);
or U16771 (N_16771,N_13234,N_12652);
nand U16772 (N_16772,N_14176,N_14128);
and U16773 (N_16773,N_14213,N_14519);
nand U16774 (N_16774,N_13065,N_14431);
nor U16775 (N_16775,N_14452,N_13093);
and U16776 (N_16776,N_13467,N_13928);
nor U16777 (N_16777,N_14558,N_13016);
xnor U16778 (N_16778,N_14195,N_14319);
and U16779 (N_16779,N_12943,N_12502);
nand U16780 (N_16780,N_12941,N_12618);
and U16781 (N_16781,N_12915,N_12966);
and U16782 (N_16782,N_13278,N_12566);
xnor U16783 (N_16783,N_14132,N_14599);
nand U16784 (N_16784,N_12894,N_13231);
xnor U16785 (N_16785,N_12763,N_13296);
xor U16786 (N_16786,N_12942,N_13519);
nand U16787 (N_16787,N_14172,N_14042);
xor U16788 (N_16788,N_12604,N_12594);
nand U16789 (N_16789,N_13965,N_14645);
xnor U16790 (N_16790,N_14081,N_14836);
or U16791 (N_16791,N_13275,N_13016);
or U16792 (N_16792,N_13438,N_13959);
nor U16793 (N_16793,N_13062,N_14725);
xnor U16794 (N_16794,N_13348,N_14607);
nand U16795 (N_16795,N_13227,N_14240);
nor U16796 (N_16796,N_12949,N_12620);
nor U16797 (N_16797,N_14035,N_12870);
or U16798 (N_16798,N_13429,N_13114);
nor U16799 (N_16799,N_14240,N_13904);
or U16800 (N_16800,N_13305,N_13569);
nand U16801 (N_16801,N_14532,N_12509);
nand U16802 (N_16802,N_12515,N_14935);
nand U16803 (N_16803,N_13623,N_13265);
nand U16804 (N_16804,N_13008,N_13814);
and U16805 (N_16805,N_13947,N_13007);
nand U16806 (N_16806,N_12622,N_14659);
or U16807 (N_16807,N_12627,N_13664);
nor U16808 (N_16808,N_14041,N_14607);
nand U16809 (N_16809,N_12520,N_12630);
xor U16810 (N_16810,N_14535,N_14170);
and U16811 (N_16811,N_14210,N_14705);
nor U16812 (N_16812,N_14375,N_13573);
nand U16813 (N_16813,N_13866,N_14475);
or U16814 (N_16814,N_13154,N_13302);
nor U16815 (N_16815,N_13678,N_14440);
nor U16816 (N_16816,N_14136,N_12906);
or U16817 (N_16817,N_14765,N_13349);
and U16818 (N_16818,N_14065,N_14306);
and U16819 (N_16819,N_13656,N_12768);
nor U16820 (N_16820,N_14774,N_14000);
or U16821 (N_16821,N_14547,N_13410);
and U16822 (N_16822,N_13775,N_13999);
nand U16823 (N_16823,N_14869,N_13695);
nor U16824 (N_16824,N_14996,N_14610);
and U16825 (N_16825,N_14972,N_13157);
or U16826 (N_16826,N_13363,N_12717);
or U16827 (N_16827,N_14493,N_12985);
and U16828 (N_16828,N_13463,N_14042);
nor U16829 (N_16829,N_13639,N_14279);
nand U16830 (N_16830,N_13991,N_13870);
or U16831 (N_16831,N_13951,N_12683);
or U16832 (N_16832,N_12591,N_12592);
xnor U16833 (N_16833,N_14676,N_13393);
nor U16834 (N_16834,N_13986,N_12501);
or U16835 (N_16835,N_14870,N_12647);
xnor U16836 (N_16836,N_13755,N_13818);
xnor U16837 (N_16837,N_14540,N_13108);
and U16838 (N_16838,N_13350,N_14677);
or U16839 (N_16839,N_14517,N_13046);
and U16840 (N_16840,N_13931,N_14567);
or U16841 (N_16841,N_14637,N_14354);
and U16842 (N_16842,N_14199,N_14268);
and U16843 (N_16843,N_14328,N_14014);
nand U16844 (N_16844,N_12663,N_12559);
xor U16845 (N_16845,N_14564,N_14686);
nor U16846 (N_16846,N_14041,N_13728);
nor U16847 (N_16847,N_12882,N_14121);
nand U16848 (N_16848,N_14988,N_13049);
xnor U16849 (N_16849,N_14568,N_13699);
or U16850 (N_16850,N_13634,N_13052);
nor U16851 (N_16851,N_13386,N_13902);
nand U16852 (N_16852,N_14821,N_13996);
nand U16853 (N_16853,N_12780,N_12611);
nor U16854 (N_16854,N_13594,N_14000);
nor U16855 (N_16855,N_12790,N_14052);
nor U16856 (N_16856,N_13917,N_14818);
or U16857 (N_16857,N_14815,N_12554);
nand U16858 (N_16858,N_14152,N_13996);
and U16859 (N_16859,N_14898,N_13152);
and U16860 (N_16860,N_14703,N_14939);
nor U16861 (N_16861,N_13870,N_14835);
or U16862 (N_16862,N_14694,N_13082);
and U16863 (N_16863,N_14478,N_12841);
or U16864 (N_16864,N_12864,N_12775);
and U16865 (N_16865,N_13704,N_13261);
nor U16866 (N_16866,N_14823,N_14485);
nand U16867 (N_16867,N_12817,N_13305);
and U16868 (N_16868,N_12966,N_13978);
xnor U16869 (N_16869,N_13144,N_12548);
or U16870 (N_16870,N_14278,N_13276);
and U16871 (N_16871,N_13529,N_13678);
or U16872 (N_16872,N_14545,N_12772);
and U16873 (N_16873,N_13507,N_14253);
xor U16874 (N_16874,N_12807,N_14397);
or U16875 (N_16875,N_13928,N_13775);
or U16876 (N_16876,N_14216,N_14419);
nor U16877 (N_16877,N_12824,N_14099);
and U16878 (N_16878,N_14545,N_14498);
and U16879 (N_16879,N_12803,N_13145);
nor U16880 (N_16880,N_14932,N_13971);
nor U16881 (N_16881,N_14466,N_13698);
xor U16882 (N_16882,N_12623,N_12917);
nor U16883 (N_16883,N_12610,N_13630);
and U16884 (N_16884,N_12806,N_14016);
nor U16885 (N_16885,N_13663,N_13807);
nand U16886 (N_16886,N_13573,N_13856);
nor U16887 (N_16887,N_14919,N_13650);
nor U16888 (N_16888,N_14099,N_13053);
xnor U16889 (N_16889,N_13077,N_13643);
xnor U16890 (N_16890,N_12770,N_13803);
nor U16891 (N_16891,N_12944,N_13854);
or U16892 (N_16892,N_12765,N_14941);
nand U16893 (N_16893,N_13160,N_13843);
nand U16894 (N_16894,N_14418,N_13417);
nand U16895 (N_16895,N_14311,N_13600);
xnor U16896 (N_16896,N_14386,N_13204);
and U16897 (N_16897,N_13602,N_14040);
and U16898 (N_16898,N_12912,N_13919);
and U16899 (N_16899,N_14108,N_14500);
and U16900 (N_16900,N_13623,N_14331);
or U16901 (N_16901,N_13903,N_14299);
or U16902 (N_16902,N_12663,N_12874);
or U16903 (N_16903,N_12611,N_14443);
nor U16904 (N_16904,N_14181,N_12848);
and U16905 (N_16905,N_13657,N_13740);
and U16906 (N_16906,N_12786,N_14146);
xnor U16907 (N_16907,N_14547,N_13117);
nand U16908 (N_16908,N_13199,N_12798);
nand U16909 (N_16909,N_14259,N_14557);
or U16910 (N_16910,N_13619,N_14246);
and U16911 (N_16911,N_13815,N_13002);
xor U16912 (N_16912,N_14243,N_14830);
nand U16913 (N_16913,N_14813,N_12696);
and U16914 (N_16914,N_13690,N_12869);
and U16915 (N_16915,N_13887,N_14434);
nor U16916 (N_16916,N_13289,N_13853);
xor U16917 (N_16917,N_14948,N_14897);
xnor U16918 (N_16918,N_14071,N_14261);
nor U16919 (N_16919,N_14562,N_12939);
or U16920 (N_16920,N_14611,N_14873);
and U16921 (N_16921,N_13632,N_14312);
nand U16922 (N_16922,N_14342,N_13134);
and U16923 (N_16923,N_13421,N_14436);
nor U16924 (N_16924,N_12524,N_13377);
xor U16925 (N_16925,N_12653,N_14839);
and U16926 (N_16926,N_14314,N_14552);
nor U16927 (N_16927,N_13016,N_14397);
and U16928 (N_16928,N_13397,N_14757);
nand U16929 (N_16929,N_13012,N_13709);
nor U16930 (N_16930,N_13301,N_14927);
nand U16931 (N_16931,N_13603,N_14558);
nand U16932 (N_16932,N_14334,N_13476);
nor U16933 (N_16933,N_13142,N_14324);
nand U16934 (N_16934,N_12784,N_12651);
or U16935 (N_16935,N_14736,N_12571);
nor U16936 (N_16936,N_14746,N_13679);
and U16937 (N_16937,N_14381,N_12938);
and U16938 (N_16938,N_14200,N_12862);
xor U16939 (N_16939,N_13428,N_13814);
nor U16940 (N_16940,N_13724,N_13065);
or U16941 (N_16941,N_13438,N_14611);
nor U16942 (N_16942,N_13588,N_13215);
or U16943 (N_16943,N_13447,N_12829);
nor U16944 (N_16944,N_12606,N_14648);
nor U16945 (N_16945,N_12853,N_13316);
and U16946 (N_16946,N_13808,N_14929);
or U16947 (N_16947,N_13169,N_13032);
nand U16948 (N_16948,N_13398,N_12746);
xnor U16949 (N_16949,N_13285,N_13422);
and U16950 (N_16950,N_13796,N_14653);
or U16951 (N_16951,N_13296,N_14753);
or U16952 (N_16952,N_12531,N_14535);
nor U16953 (N_16953,N_14115,N_12626);
xnor U16954 (N_16954,N_13795,N_14595);
xor U16955 (N_16955,N_14730,N_13087);
nand U16956 (N_16956,N_12616,N_14147);
nor U16957 (N_16957,N_12744,N_13568);
nand U16958 (N_16958,N_14479,N_13363);
or U16959 (N_16959,N_14523,N_14595);
nand U16960 (N_16960,N_14909,N_13019);
and U16961 (N_16961,N_14420,N_13033);
or U16962 (N_16962,N_13039,N_14477);
xor U16963 (N_16963,N_13203,N_13605);
or U16964 (N_16964,N_14646,N_13797);
nand U16965 (N_16965,N_13944,N_13598);
nor U16966 (N_16966,N_13101,N_12761);
nor U16967 (N_16967,N_14371,N_12719);
nor U16968 (N_16968,N_13295,N_14830);
nand U16969 (N_16969,N_13799,N_14431);
xor U16970 (N_16970,N_13078,N_13776);
nor U16971 (N_16971,N_13650,N_14932);
and U16972 (N_16972,N_14707,N_13937);
or U16973 (N_16973,N_12826,N_13280);
xor U16974 (N_16974,N_14842,N_13408);
and U16975 (N_16975,N_14732,N_12740);
or U16976 (N_16976,N_14590,N_14844);
nand U16977 (N_16977,N_13090,N_14429);
and U16978 (N_16978,N_14253,N_13246);
nor U16979 (N_16979,N_13533,N_13679);
and U16980 (N_16980,N_12582,N_14557);
and U16981 (N_16981,N_12768,N_14826);
nand U16982 (N_16982,N_12501,N_12571);
or U16983 (N_16983,N_14100,N_13581);
nand U16984 (N_16984,N_14161,N_13864);
and U16985 (N_16985,N_12768,N_12991);
xor U16986 (N_16986,N_12994,N_14132);
nand U16987 (N_16987,N_14128,N_14973);
nor U16988 (N_16988,N_14027,N_13724);
or U16989 (N_16989,N_13245,N_13106);
nand U16990 (N_16990,N_12889,N_13595);
and U16991 (N_16991,N_13955,N_13081);
xnor U16992 (N_16992,N_14772,N_13557);
nand U16993 (N_16993,N_14295,N_13833);
xor U16994 (N_16994,N_13889,N_12538);
nor U16995 (N_16995,N_13404,N_13906);
and U16996 (N_16996,N_14691,N_14873);
or U16997 (N_16997,N_14017,N_13535);
xor U16998 (N_16998,N_12973,N_12623);
xnor U16999 (N_16999,N_14427,N_13892);
nand U17000 (N_17000,N_14744,N_13397);
xnor U17001 (N_17001,N_14978,N_13338);
nand U17002 (N_17002,N_14119,N_14395);
nand U17003 (N_17003,N_14044,N_13228);
nor U17004 (N_17004,N_13364,N_14392);
or U17005 (N_17005,N_13115,N_13802);
or U17006 (N_17006,N_13719,N_14565);
nor U17007 (N_17007,N_13879,N_13309);
xnor U17008 (N_17008,N_13312,N_13672);
and U17009 (N_17009,N_13396,N_14947);
nor U17010 (N_17010,N_13122,N_13045);
and U17011 (N_17011,N_14386,N_13778);
xnor U17012 (N_17012,N_12551,N_13777);
xnor U17013 (N_17013,N_14783,N_13182);
and U17014 (N_17014,N_14153,N_13564);
and U17015 (N_17015,N_13783,N_13928);
nand U17016 (N_17016,N_12712,N_12533);
nor U17017 (N_17017,N_13468,N_13260);
xor U17018 (N_17018,N_14203,N_13266);
and U17019 (N_17019,N_13723,N_14595);
or U17020 (N_17020,N_14556,N_13740);
and U17021 (N_17021,N_13849,N_14421);
and U17022 (N_17022,N_12815,N_14662);
nor U17023 (N_17023,N_13944,N_14605);
nor U17024 (N_17024,N_12969,N_12981);
or U17025 (N_17025,N_12610,N_13721);
or U17026 (N_17026,N_13949,N_12894);
and U17027 (N_17027,N_13841,N_14585);
nor U17028 (N_17028,N_12555,N_13634);
xnor U17029 (N_17029,N_13901,N_13927);
nand U17030 (N_17030,N_13135,N_12696);
and U17031 (N_17031,N_13269,N_12798);
xnor U17032 (N_17032,N_14022,N_13029);
and U17033 (N_17033,N_13010,N_12572);
and U17034 (N_17034,N_14700,N_13925);
and U17035 (N_17035,N_13775,N_13652);
nand U17036 (N_17036,N_13418,N_14751);
nand U17037 (N_17037,N_14525,N_14058);
and U17038 (N_17038,N_12742,N_14507);
or U17039 (N_17039,N_14193,N_14324);
and U17040 (N_17040,N_13113,N_14698);
nor U17041 (N_17041,N_13676,N_14384);
nand U17042 (N_17042,N_12654,N_12887);
or U17043 (N_17043,N_13128,N_13276);
xor U17044 (N_17044,N_13089,N_12769);
nand U17045 (N_17045,N_13221,N_13860);
xnor U17046 (N_17046,N_14311,N_13407);
nand U17047 (N_17047,N_14240,N_14501);
nand U17048 (N_17048,N_13001,N_14231);
xor U17049 (N_17049,N_13704,N_12551);
nand U17050 (N_17050,N_14725,N_14583);
and U17051 (N_17051,N_13141,N_13084);
nand U17052 (N_17052,N_13775,N_13398);
nand U17053 (N_17053,N_12517,N_13681);
nor U17054 (N_17054,N_12533,N_12577);
or U17055 (N_17055,N_14917,N_12601);
nand U17056 (N_17056,N_14764,N_13672);
or U17057 (N_17057,N_14881,N_12658);
or U17058 (N_17058,N_13674,N_14833);
or U17059 (N_17059,N_14045,N_13057);
and U17060 (N_17060,N_14846,N_14327);
or U17061 (N_17061,N_13325,N_14963);
nor U17062 (N_17062,N_12818,N_14504);
xor U17063 (N_17063,N_12702,N_12715);
and U17064 (N_17064,N_14264,N_14281);
xor U17065 (N_17065,N_13481,N_14501);
nor U17066 (N_17066,N_13071,N_13195);
xor U17067 (N_17067,N_14630,N_13292);
and U17068 (N_17068,N_14618,N_14764);
or U17069 (N_17069,N_12976,N_14484);
nor U17070 (N_17070,N_13250,N_12934);
nor U17071 (N_17071,N_13559,N_14055);
xor U17072 (N_17072,N_14507,N_14799);
xnor U17073 (N_17073,N_14351,N_13737);
nand U17074 (N_17074,N_13636,N_14618);
xnor U17075 (N_17075,N_14252,N_13892);
nand U17076 (N_17076,N_14730,N_14117);
and U17077 (N_17077,N_13271,N_13863);
nor U17078 (N_17078,N_12566,N_14785);
and U17079 (N_17079,N_14447,N_14019);
nor U17080 (N_17080,N_12680,N_13550);
and U17081 (N_17081,N_13270,N_14000);
xnor U17082 (N_17082,N_13634,N_14711);
nand U17083 (N_17083,N_12740,N_14977);
and U17084 (N_17084,N_13991,N_14375);
nor U17085 (N_17085,N_13217,N_14096);
and U17086 (N_17086,N_13519,N_13426);
xnor U17087 (N_17087,N_14424,N_13627);
nor U17088 (N_17088,N_14168,N_14731);
nor U17089 (N_17089,N_12580,N_13000);
nor U17090 (N_17090,N_14209,N_13641);
and U17091 (N_17091,N_14771,N_14589);
xnor U17092 (N_17092,N_13127,N_12598);
nor U17093 (N_17093,N_14407,N_14181);
xnor U17094 (N_17094,N_14510,N_12975);
nand U17095 (N_17095,N_13241,N_14186);
xnor U17096 (N_17096,N_12784,N_13508);
xnor U17097 (N_17097,N_14565,N_12591);
xor U17098 (N_17098,N_13626,N_14250);
nand U17099 (N_17099,N_14923,N_14609);
nor U17100 (N_17100,N_13513,N_14439);
nand U17101 (N_17101,N_14487,N_14300);
nor U17102 (N_17102,N_14972,N_13904);
nor U17103 (N_17103,N_12865,N_14058);
xor U17104 (N_17104,N_14654,N_14608);
or U17105 (N_17105,N_13981,N_14747);
and U17106 (N_17106,N_14185,N_13063);
xnor U17107 (N_17107,N_14177,N_14086);
and U17108 (N_17108,N_13235,N_13096);
or U17109 (N_17109,N_14222,N_14817);
and U17110 (N_17110,N_14389,N_13932);
or U17111 (N_17111,N_13696,N_12595);
or U17112 (N_17112,N_12765,N_12685);
and U17113 (N_17113,N_13535,N_12779);
or U17114 (N_17114,N_14073,N_13471);
and U17115 (N_17115,N_13684,N_14103);
nor U17116 (N_17116,N_13134,N_13653);
xor U17117 (N_17117,N_12627,N_13312);
nor U17118 (N_17118,N_13257,N_13719);
or U17119 (N_17119,N_14357,N_12944);
nor U17120 (N_17120,N_12880,N_12812);
nand U17121 (N_17121,N_13178,N_12707);
or U17122 (N_17122,N_12858,N_13065);
nor U17123 (N_17123,N_12891,N_12553);
nand U17124 (N_17124,N_13852,N_12561);
xnor U17125 (N_17125,N_14316,N_14085);
nand U17126 (N_17126,N_14181,N_14530);
nor U17127 (N_17127,N_12608,N_14096);
nor U17128 (N_17128,N_12980,N_13612);
or U17129 (N_17129,N_14440,N_13727);
or U17130 (N_17130,N_13546,N_13625);
xnor U17131 (N_17131,N_12912,N_12707);
and U17132 (N_17132,N_13731,N_12878);
or U17133 (N_17133,N_13438,N_12871);
or U17134 (N_17134,N_14961,N_14499);
nor U17135 (N_17135,N_13383,N_14473);
and U17136 (N_17136,N_13070,N_12532);
and U17137 (N_17137,N_14325,N_13875);
nor U17138 (N_17138,N_13021,N_13848);
xnor U17139 (N_17139,N_14178,N_13831);
nor U17140 (N_17140,N_14423,N_13629);
xnor U17141 (N_17141,N_12802,N_14339);
nand U17142 (N_17142,N_12892,N_12949);
or U17143 (N_17143,N_13151,N_14779);
xnor U17144 (N_17144,N_13427,N_13515);
nand U17145 (N_17145,N_13222,N_13689);
nor U17146 (N_17146,N_13677,N_14027);
nor U17147 (N_17147,N_13257,N_13114);
nand U17148 (N_17148,N_14061,N_13964);
or U17149 (N_17149,N_14367,N_13346);
nand U17150 (N_17150,N_13094,N_12620);
or U17151 (N_17151,N_12531,N_14658);
nor U17152 (N_17152,N_12926,N_14399);
xnor U17153 (N_17153,N_13182,N_14946);
nand U17154 (N_17154,N_14516,N_12648);
nand U17155 (N_17155,N_13560,N_12884);
or U17156 (N_17156,N_13511,N_13676);
nand U17157 (N_17157,N_12579,N_14065);
nand U17158 (N_17158,N_12564,N_13744);
nor U17159 (N_17159,N_13142,N_13044);
nand U17160 (N_17160,N_12636,N_13073);
xor U17161 (N_17161,N_14787,N_12943);
and U17162 (N_17162,N_13726,N_13124);
or U17163 (N_17163,N_13358,N_14318);
or U17164 (N_17164,N_14659,N_13339);
xnor U17165 (N_17165,N_14321,N_14268);
xnor U17166 (N_17166,N_13895,N_13828);
nand U17167 (N_17167,N_13793,N_14801);
nor U17168 (N_17168,N_13116,N_14031);
nor U17169 (N_17169,N_14773,N_13768);
nor U17170 (N_17170,N_12627,N_14822);
nor U17171 (N_17171,N_13027,N_13194);
nand U17172 (N_17172,N_14057,N_13236);
and U17173 (N_17173,N_13565,N_13194);
xor U17174 (N_17174,N_14298,N_13658);
and U17175 (N_17175,N_13835,N_12520);
nor U17176 (N_17176,N_14575,N_12533);
and U17177 (N_17177,N_13602,N_14921);
xnor U17178 (N_17178,N_13144,N_12860);
nand U17179 (N_17179,N_14014,N_13397);
and U17180 (N_17180,N_14942,N_12582);
and U17181 (N_17181,N_12862,N_14420);
or U17182 (N_17182,N_14482,N_14237);
nor U17183 (N_17183,N_13018,N_14254);
nor U17184 (N_17184,N_13587,N_14382);
xnor U17185 (N_17185,N_13890,N_12745);
nand U17186 (N_17186,N_13940,N_13308);
nand U17187 (N_17187,N_14641,N_13790);
nor U17188 (N_17188,N_14097,N_13302);
xor U17189 (N_17189,N_13903,N_14380);
and U17190 (N_17190,N_14979,N_13281);
and U17191 (N_17191,N_13153,N_12568);
xor U17192 (N_17192,N_13496,N_12618);
xnor U17193 (N_17193,N_13716,N_14315);
nand U17194 (N_17194,N_13835,N_14000);
nor U17195 (N_17195,N_12518,N_14391);
nand U17196 (N_17196,N_13019,N_14817);
nand U17197 (N_17197,N_14529,N_14270);
xnor U17198 (N_17198,N_13588,N_13926);
nor U17199 (N_17199,N_14573,N_12717);
xnor U17200 (N_17200,N_13006,N_14126);
and U17201 (N_17201,N_12696,N_12598);
and U17202 (N_17202,N_13238,N_14732);
nand U17203 (N_17203,N_14236,N_12620);
nand U17204 (N_17204,N_13761,N_13677);
nor U17205 (N_17205,N_13268,N_13197);
nand U17206 (N_17206,N_13360,N_13713);
xnor U17207 (N_17207,N_14188,N_12570);
nand U17208 (N_17208,N_13666,N_13530);
or U17209 (N_17209,N_14412,N_13456);
or U17210 (N_17210,N_12662,N_14126);
xnor U17211 (N_17211,N_13104,N_12890);
nand U17212 (N_17212,N_12946,N_14475);
nor U17213 (N_17213,N_13360,N_14403);
xnor U17214 (N_17214,N_12876,N_13024);
and U17215 (N_17215,N_13758,N_13075);
nor U17216 (N_17216,N_13722,N_12508);
nand U17217 (N_17217,N_13675,N_13412);
nor U17218 (N_17218,N_12738,N_12646);
nand U17219 (N_17219,N_14227,N_13406);
nor U17220 (N_17220,N_13193,N_13257);
and U17221 (N_17221,N_14344,N_14528);
and U17222 (N_17222,N_14163,N_13083);
and U17223 (N_17223,N_13719,N_14439);
nand U17224 (N_17224,N_12779,N_12517);
xnor U17225 (N_17225,N_13020,N_13456);
or U17226 (N_17226,N_13631,N_12594);
and U17227 (N_17227,N_13414,N_13809);
xor U17228 (N_17228,N_14413,N_13067);
xor U17229 (N_17229,N_12898,N_13314);
and U17230 (N_17230,N_14244,N_14996);
xnor U17231 (N_17231,N_14307,N_12732);
xor U17232 (N_17232,N_12536,N_13599);
and U17233 (N_17233,N_14122,N_13824);
nor U17234 (N_17234,N_12769,N_13720);
xor U17235 (N_17235,N_13041,N_12716);
nor U17236 (N_17236,N_14320,N_12982);
nand U17237 (N_17237,N_12596,N_14340);
xor U17238 (N_17238,N_14708,N_14577);
and U17239 (N_17239,N_14580,N_13709);
and U17240 (N_17240,N_12657,N_13969);
or U17241 (N_17241,N_13024,N_14355);
xor U17242 (N_17242,N_14213,N_14318);
nor U17243 (N_17243,N_14093,N_13726);
or U17244 (N_17244,N_14415,N_13574);
and U17245 (N_17245,N_14049,N_13101);
xor U17246 (N_17246,N_13694,N_14983);
and U17247 (N_17247,N_14243,N_14522);
nand U17248 (N_17248,N_13789,N_14666);
nand U17249 (N_17249,N_13838,N_13042);
xnor U17250 (N_17250,N_14950,N_13202);
xnor U17251 (N_17251,N_14339,N_14021);
and U17252 (N_17252,N_13985,N_14052);
or U17253 (N_17253,N_12744,N_12609);
nand U17254 (N_17254,N_12839,N_13057);
nand U17255 (N_17255,N_13684,N_13601);
and U17256 (N_17256,N_14833,N_13001);
nor U17257 (N_17257,N_13707,N_13708);
and U17258 (N_17258,N_14374,N_14603);
nand U17259 (N_17259,N_13868,N_13180);
nand U17260 (N_17260,N_13594,N_13380);
nand U17261 (N_17261,N_12539,N_14183);
nand U17262 (N_17262,N_14097,N_13355);
nor U17263 (N_17263,N_14485,N_13503);
nor U17264 (N_17264,N_12978,N_12726);
and U17265 (N_17265,N_14001,N_13039);
or U17266 (N_17266,N_12901,N_13715);
nand U17267 (N_17267,N_13020,N_13341);
or U17268 (N_17268,N_13872,N_12702);
and U17269 (N_17269,N_12776,N_14160);
and U17270 (N_17270,N_12579,N_13633);
nor U17271 (N_17271,N_14294,N_12979);
nand U17272 (N_17272,N_13477,N_13468);
nor U17273 (N_17273,N_14447,N_14129);
and U17274 (N_17274,N_12980,N_13247);
nand U17275 (N_17275,N_14612,N_13783);
xnor U17276 (N_17276,N_12926,N_13302);
nand U17277 (N_17277,N_13547,N_13942);
xnor U17278 (N_17278,N_13702,N_12956);
xor U17279 (N_17279,N_14616,N_14771);
nand U17280 (N_17280,N_13564,N_14919);
nand U17281 (N_17281,N_14740,N_14273);
nor U17282 (N_17282,N_13820,N_14949);
and U17283 (N_17283,N_13220,N_13768);
xnor U17284 (N_17284,N_13797,N_13087);
and U17285 (N_17285,N_13645,N_14976);
nor U17286 (N_17286,N_12820,N_14860);
xnor U17287 (N_17287,N_12537,N_12959);
nor U17288 (N_17288,N_12956,N_13211);
nand U17289 (N_17289,N_14295,N_12841);
nand U17290 (N_17290,N_14366,N_14033);
nand U17291 (N_17291,N_13768,N_13536);
or U17292 (N_17292,N_13058,N_12557);
xor U17293 (N_17293,N_13358,N_13404);
xnor U17294 (N_17294,N_12930,N_13575);
nand U17295 (N_17295,N_13271,N_14483);
nand U17296 (N_17296,N_13736,N_14262);
and U17297 (N_17297,N_13186,N_13385);
xor U17298 (N_17298,N_12821,N_13391);
or U17299 (N_17299,N_13121,N_12968);
xor U17300 (N_17300,N_13153,N_13033);
xnor U17301 (N_17301,N_14572,N_13182);
nor U17302 (N_17302,N_13598,N_12518);
nand U17303 (N_17303,N_14796,N_13094);
nand U17304 (N_17304,N_14913,N_13995);
or U17305 (N_17305,N_13797,N_13736);
and U17306 (N_17306,N_14260,N_13285);
or U17307 (N_17307,N_14567,N_12795);
nand U17308 (N_17308,N_13960,N_12636);
nor U17309 (N_17309,N_13093,N_14781);
or U17310 (N_17310,N_13998,N_13816);
nor U17311 (N_17311,N_12643,N_13497);
and U17312 (N_17312,N_14176,N_13745);
or U17313 (N_17313,N_14379,N_12759);
nor U17314 (N_17314,N_14019,N_14218);
xor U17315 (N_17315,N_13699,N_13721);
or U17316 (N_17316,N_14326,N_12629);
nor U17317 (N_17317,N_14441,N_14459);
and U17318 (N_17318,N_13006,N_13090);
xor U17319 (N_17319,N_14259,N_14097);
nand U17320 (N_17320,N_12713,N_14652);
nand U17321 (N_17321,N_14707,N_14980);
nand U17322 (N_17322,N_13852,N_12510);
or U17323 (N_17323,N_14778,N_12878);
nand U17324 (N_17324,N_13197,N_14253);
nor U17325 (N_17325,N_12929,N_14779);
and U17326 (N_17326,N_14083,N_13642);
and U17327 (N_17327,N_13369,N_12855);
nor U17328 (N_17328,N_12575,N_13166);
nor U17329 (N_17329,N_14309,N_14461);
or U17330 (N_17330,N_12829,N_14478);
xor U17331 (N_17331,N_14245,N_14242);
or U17332 (N_17332,N_13675,N_14088);
nand U17333 (N_17333,N_12943,N_13136);
nor U17334 (N_17334,N_13415,N_13229);
nand U17335 (N_17335,N_14168,N_14555);
and U17336 (N_17336,N_14518,N_14625);
xor U17337 (N_17337,N_13807,N_14983);
xnor U17338 (N_17338,N_14781,N_12931);
xor U17339 (N_17339,N_13343,N_14879);
or U17340 (N_17340,N_13361,N_13749);
xor U17341 (N_17341,N_13764,N_12684);
or U17342 (N_17342,N_13736,N_13555);
nand U17343 (N_17343,N_13819,N_13241);
or U17344 (N_17344,N_13518,N_13213);
nor U17345 (N_17345,N_14497,N_14139);
xor U17346 (N_17346,N_13478,N_13175);
nor U17347 (N_17347,N_14167,N_12733);
or U17348 (N_17348,N_12677,N_14796);
nand U17349 (N_17349,N_14982,N_14051);
nand U17350 (N_17350,N_13583,N_14006);
nand U17351 (N_17351,N_12859,N_13760);
nor U17352 (N_17352,N_14396,N_14127);
xor U17353 (N_17353,N_12877,N_14254);
nand U17354 (N_17354,N_14085,N_14240);
nand U17355 (N_17355,N_13237,N_13666);
xor U17356 (N_17356,N_13905,N_12987);
nand U17357 (N_17357,N_13628,N_13787);
and U17358 (N_17358,N_14415,N_14220);
nand U17359 (N_17359,N_14607,N_13086);
nor U17360 (N_17360,N_13844,N_12700);
and U17361 (N_17361,N_14097,N_14953);
nor U17362 (N_17362,N_13772,N_13955);
nor U17363 (N_17363,N_12683,N_13727);
or U17364 (N_17364,N_12674,N_14101);
nor U17365 (N_17365,N_12562,N_14604);
nand U17366 (N_17366,N_13812,N_12765);
nor U17367 (N_17367,N_13611,N_12548);
and U17368 (N_17368,N_14354,N_13530);
or U17369 (N_17369,N_14415,N_13940);
xor U17370 (N_17370,N_13401,N_13884);
and U17371 (N_17371,N_14984,N_13838);
nand U17372 (N_17372,N_13982,N_12651);
xnor U17373 (N_17373,N_12539,N_13475);
nand U17374 (N_17374,N_13635,N_13980);
and U17375 (N_17375,N_14941,N_14237);
nor U17376 (N_17376,N_13387,N_14857);
or U17377 (N_17377,N_14970,N_12501);
nor U17378 (N_17378,N_14203,N_12677);
nand U17379 (N_17379,N_12933,N_13825);
and U17380 (N_17380,N_14269,N_14079);
xnor U17381 (N_17381,N_13589,N_14933);
nor U17382 (N_17382,N_13935,N_12617);
nor U17383 (N_17383,N_14999,N_13027);
and U17384 (N_17384,N_13395,N_12506);
and U17385 (N_17385,N_14547,N_14260);
nor U17386 (N_17386,N_12865,N_13020);
nor U17387 (N_17387,N_12727,N_13631);
or U17388 (N_17388,N_14703,N_14627);
and U17389 (N_17389,N_12982,N_14331);
and U17390 (N_17390,N_13145,N_13238);
or U17391 (N_17391,N_14235,N_14795);
and U17392 (N_17392,N_14945,N_12579);
and U17393 (N_17393,N_14123,N_13109);
nand U17394 (N_17394,N_14018,N_14660);
xor U17395 (N_17395,N_13396,N_12537);
xnor U17396 (N_17396,N_14321,N_14353);
nand U17397 (N_17397,N_13847,N_14734);
nor U17398 (N_17398,N_14719,N_12595);
nor U17399 (N_17399,N_13996,N_13842);
or U17400 (N_17400,N_13633,N_13875);
xnor U17401 (N_17401,N_14935,N_14020);
or U17402 (N_17402,N_13629,N_12625);
nor U17403 (N_17403,N_14378,N_13693);
nor U17404 (N_17404,N_12866,N_14099);
nand U17405 (N_17405,N_13695,N_14671);
and U17406 (N_17406,N_13626,N_13455);
or U17407 (N_17407,N_13820,N_14639);
nand U17408 (N_17408,N_14611,N_12691);
xnor U17409 (N_17409,N_13264,N_13372);
nor U17410 (N_17410,N_12867,N_13909);
nor U17411 (N_17411,N_12863,N_14473);
nand U17412 (N_17412,N_13000,N_13239);
nand U17413 (N_17413,N_13155,N_14566);
xor U17414 (N_17414,N_12971,N_12803);
nor U17415 (N_17415,N_14678,N_12816);
or U17416 (N_17416,N_14610,N_12953);
xnor U17417 (N_17417,N_13205,N_12959);
and U17418 (N_17418,N_13184,N_12870);
and U17419 (N_17419,N_13805,N_14768);
and U17420 (N_17420,N_12953,N_14322);
xor U17421 (N_17421,N_12955,N_13408);
or U17422 (N_17422,N_12938,N_13987);
or U17423 (N_17423,N_14725,N_13156);
xnor U17424 (N_17424,N_12744,N_13126);
nor U17425 (N_17425,N_14320,N_12912);
nor U17426 (N_17426,N_13136,N_13788);
or U17427 (N_17427,N_13331,N_13680);
xnor U17428 (N_17428,N_13760,N_12609);
nand U17429 (N_17429,N_14025,N_13340);
xor U17430 (N_17430,N_12539,N_14553);
xor U17431 (N_17431,N_14015,N_13611);
nor U17432 (N_17432,N_12682,N_14123);
nor U17433 (N_17433,N_14344,N_13726);
xnor U17434 (N_17434,N_13806,N_12503);
xor U17435 (N_17435,N_14599,N_14169);
nor U17436 (N_17436,N_13703,N_12935);
nor U17437 (N_17437,N_14174,N_14841);
xnor U17438 (N_17438,N_14782,N_14098);
nor U17439 (N_17439,N_12696,N_13550);
or U17440 (N_17440,N_14647,N_14854);
nor U17441 (N_17441,N_14384,N_12771);
and U17442 (N_17442,N_12959,N_14340);
nor U17443 (N_17443,N_12695,N_13071);
nand U17444 (N_17444,N_12505,N_12968);
nor U17445 (N_17445,N_14730,N_14651);
and U17446 (N_17446,N_14678,N_13381);
and U17447 (N_17447,N_14746,N_14256);
xnor U17448 (N_17448,N_14167,N_13546);
and U17449 (N_17449,N_13500,N_14734);
xor U17450 (N_17450,N_14417,N_14068);
xor U17451 (N_17451,N_13101,N_14121);
nor U17452 (N_17452,N_14101,N_14585);
xor U17453 (N_17453,N_12809,N_12848);
or U17454 (N_17454,N_13166,N_13722);
xor U17455 (N_17455,N_12653,N_12875);
xnor U17456 (N_17456,N_14961,N_14401);
and U17457 (N_17457,N_12548,N_13568);
nand U17458 (N_17458,N_14412,N_12698);
nand U17459 (N_17459,N_13380,N_14091);
or U17460 (N_17460,N_12616,N_13972);
xor U17461 (N_17461,N_13017,N_14347);
or U17462 (N_17462,N_13867,N_14069);
xnor U17463 (N_17463,N_13858,N_13785);
and U17464 (N_17464,N_13269,N_13336);
nor U17465 (N_17465,N_14215,N_14524);
xnor U17466 (N_17466,N_14997,N_13931);
or U17467 (N_17467,N_13729,N_14295);
and U17468 (N_17468,N_13427,N_13913);
xnor U17469 (N_17469,N_14924,N_13867);
nand U17470 (N_17470,N_14894,N_14719);
or U17471 (N_17471,N_13527,N_13080);
nand U17472 (N_17472,N_14339,N_14722);
nand U17473 (N_17473,N_13859,N_13721);
nand U17474 (N_17474,N_12825,N_13452);
xor U17475 (N_17475,N_12571,N_14053);
xnor U17476 (N_17476,N_14634,N_12797);
or U17477 (N_17477,N_13177,N_14458);
nor U17478 (N_17478,N_12510,N_13095);
xor U17479 (N_17479,N_13443,N_14520);
nand U17480 (N_17480,N_13388,N_14646);
or U17481 (N_17481,N_14920,N_13223);
and U17482 (N_17482,N_13547,N_14743);
or U17483 (N_17483,N_13205,N_13922);
and U17484 (N_17484,N_13999,N_14335);
xnor U17485 (N_17485,N_13472,N_13246);
or U17486 (N_17486,N_13600,N_12865);
or U17487 (N_17487,N_13088,N_14095);
nand U17488 (N_17488,N_12698,N_14509);
nor U17489 (N_17489,N_12766,N_14513);
xnor U17490 (N_17490,N_14407,N_14857);
and U17491 (N_17491,N_12502,N_12893);
nand U17492 (N_17492,N_13076,N_14381);
xor U17493 (N_17493,N_13589,N_12892);
nand U17494 (N_17494,N_14624,N_12643);
xnor U17495 (N_17495,N_13801,N_14103);
and U17496 (N_17496,N_14712,N_12862);
and U17497 (N_17497,N_13399,N_13861);
and U17498 (N_17498,N_12758,N_13821);
xnor U17499 (N_17499,N_13257,N_14157);
and U17500 (N_17500,N_15711,N_16882);
nand U17501 (N_17501,N_15006,N_17443);
or U17502 (N_17502,N_17003,N_16721);
or U17503 (N_17503,N_15094,N_17041);
nor U17504 (N_17504,N_16264,N_17284);
nor U17505 (N_17505,N_17249,N_15222);
and U17506 (N_17506,N_17319,N_16683);
nor U17507 (N_17507,N_17416,N_15944);
and U17508 (N_17508,N_17239,N_17316);
nor U17509 (N_17509,N_15990,N_17179);
nand U17510 (N_17510,N_15244,N_15730);
nand U17511 (N_17511,N_17260,N_17430);
xor U17512 (N_17512,N_16612,N_16821);
or U17513 (N_17513,N_17195,N_16674);
and U17514 (N_17514,N_15699,N_16074);
and U17515 (N_17515,N_16896,N_15855);
nor U17516 (N_17516,N_15241,N_15032);
nand U17517 (N_17517,N_15100,N_15782);
or U17518 (N_17518,N_15559,N_17445);
xnor U17519 (N_17519,N_16258,N_15258);
or U17520 (N_17520,N_16504,N_15727);
xor U17521 (N_17521,N_15012,N_17196);
and U17522 (N_17522,N_16594,N_17476);
and U17523 (N_17523,N_15413,N_16075);
xor U17524 (N_17524,N_16667,N_16278);
or U17525 (N_17525,N_16414,N_17061);
nor U17526 (N_17526,N_15824,N_15147);
or U17527 (N_17527,N_15407,N_17202);
or U17528 (N_17528,N_15203,N_17494);
nor U17529 (N_17529,N_15941,N_16960);
and U17530 (N_17530,N_16863,N_16608);
nor U17531 (N_17531,N_16233,N_15485);
nand U17532 (N_17532,N_16870,N_16575);
nor U17533 (N_17533,N_15090,N_15969);
or U17534 (N_17534,N_15024,N_17111);
nor U17535 (N_17535,N_16828,N_17221);
nand U17536 (N_17536,N_17299,N_15743);
nand U17537 (N_17537,N_15405,N_15349);
xor U17538 (N_17538,N_16627,N_17408);
xor U17539 (N_17539,N_17368,N_16623);
nand U17540 (N_17540,N_17357,N_16364);
xnor U17541 (N_17541,N_16423,N_16565);
nor U17542 (N_17542,N_17164,N_16046);
nor U17543 (N_17543,N_15048,N_16617);
xnor U17544 (N_17544,N_15393,N_16665);
or U17545 (N_17545,N_16010,N_16970);
nor U17546 (N_17546,N_16854,N_16611);
nor U17547 (N_17547,N_17081,N_16006);
xor U17548 (N_17548,N_16374,N_16697);
xor U17549 (N_17549,N_15380,N_15851);
or U17550 (N_17550,N_16957,N_16492);
or U17551 (N_17551,N_16985,N_17049);
xor U17552 (N_17552,N_16950,N_16929);
or U17553 (N_17553,N_16535,N_16057);
nand U17554 (N_17554,N_15123,N_15338);
and U17555 (N_17555,N_17488,N_16124);
xnor U17556 (N_17556,N_17439,N_15301);
xnor U17557 (N_17557,N_16591,N_15604);
and U17558 (N_17558,N_16754,N_15206);
nand U17559 (N_17559,N_17293,N_17112);
nor U17560 (N_17560,N_15544,N_16867);
or U17561 (N_17561,N_17171,N_16537);
xor U17562 (N_17562,N_15273,N_16467);
or U17563 (N_17563,N_15976,N_16241);
and U17564 (N_17564,N_15850,N_17103);
or U17565 (N_17565,N_16853,N_15908);
xor U17566 (N_17566,N_16779,N_15849);
nor U17567 (N_17567,N_17248,N_15439);
nand U17568 (N_17568,N_16732,N_15932);
or U17569 (N_17569,N_17339,N_16763);
xor U17570 (N_17570,N_15326,N_15109);
nor U17571 (N_17571,N_16631,N_15419);
xor U17572 (N_17572,N_16085,N_15539);
xnor U17573 (N_17573,N_15896,N_17089);
nor U17574 (N_17574,N_16687,N_15418);
nor U17575 (N_17575,N_15140,N_16522);
xor U17576 (N_17576,N_17331,N_17454);
and U17577 (N_17577,N_16357,N_15592);
nand U17578 (N_17578,N_16941,N_17148);
or U17579 (N_17579,N_15160,N_16373);
nor U17580 (N_17580,N_16688,N_17124);
xnor U17581 (N_17581,N_16826,N_17129);
xor U17582 (N_17582,N_16160,N_15839);
and U17583 (N_17583,N_15830,N_16829);
nand U17584 (N_17584,N_16865,N_17270);
nand U17585 (N_17585,N_16254,N_16165);
and U17586 (N_17586,N_15083,N_15387);
nor U17587 (N_17587,N_17345,N_16028);
nand U17588 (N_17588,N_15848,N_17291);
nor U17589 (N_17589,N_16061,N_15398);
nor U17590 (N_17590,N_17477,N_17093);
nand U17591 (N_17591,N_15101,N_17166);
or U17592 (N_17592,N_16093,N_16992);
xor U17593 (N_17593,N_16285,N_15652);
nor U17594 (N_17594,N_15069,N_16243);
nor U17595 (N_17595,N_17037,N_16933);
and U17596 (N_17596,N_15589,N_16881);
nand U17597 (N_17597,N_16066,N_17203);
nor U17598 (N_17598,N_15721,N_16224);
and U17599 (N_17599,N_16604,N_16544);
and U17600 (N_17600,N_17432,N_15605);
nor U17601 (N_17601,N_15564,N_17114);
and U17602 (N_17602,N_16184,N_15579);
nor U17603 (N_17603,N_17255,N_15498);
nor U17604 (N_17604,N_17096,N_17243);
or U17605 (N_17605,N_15474,N_15791);
nand U17606 (N_17606,N_17022,N_16990);
or U17607 (N_17607,N_16847,N_17176);
xnor U17608 (N_17608,N_15845,N_17306);
or U17609 (N_17609,N_17446,N_15557);
and U17610 (N_17610,N_17383,N_15171);
or U17611 (N_17611,N_15622,N_16446);
or U17612 (N_17612,N_16197,N_16448);
and U17613 (N_17613,N_16416,N_16549);
nor U17614 (N_17614,N_15285,N_15663);
and U17615 (N_17615,N_17286,N_15490);
or U17616 (N_17616,N_15831,N_16155);
and U17617 (N_17617,N_15449,N_16482);
xnor U17618 (N_17618,N_17363,N_16660);
and U17619 (N_17619,N_15630,N_15166);
xor U17620 (N_17620,N_15187,N_15263);
or U17621 (N_17621,N_15547,N_16669);
xor U17622 (N_17622,N_15017,N_16104);
nand U17623 (N_17623,N_15129,N_16478);
nor U17624 (N_17624,N_17138,N_16410);
nand U17625 (N_17625,N_16917,N_16681);
xor U17626 (N_17626,N_15808,N_17263);
and U17627 (N_17627,N_17497,N_17487);
xor U17628 (N_17628,N_16495,N_16808);
nand U17629 (N_17629,N_15164,N_16127);
xnor U17630 (N_17630,N_16561,N_16043);
and U17631 (N_17631,N_16056,N_16550);
or U17632 (N_17632,N_16835,N_16791);
nor U17633 (N_17633,N_16520,N_15108);
xor U17634 (N_17634,N_17119,N_16106);
nor U17635 (N_17635,N_16614,N_17174);
or U17636 (N_17636,N_16015,N_16920);
or U17637 (N_17637,N_16477,N_16441);
nor U17638 (N_17638,N_15395,N_16206);
nand U17639 (N_17639,N_16111,N_15335);
xor U17640 (N_17640,N_17123,N_16768);
and U17641 (N_17641,N_15517,N_16217);
and U17642 (N_17642,N_16137,N_16432);
nor U17643 (N_17643,N_16359,N_17144);
or U17644 (N_17644,N_15359,N_16459);
nor U17645 (N_17645,N_15327,N_16802);
and U17646 (N_17646,N_17264,N_16112);
and U17647 (N_17647,N_16142,N_16260);
or U17648 (N_17648,N_17104,N_15909);
or U17649 (N_17649,N_17281,N_15228);
and U17650 (N_17650,N_15370,N_17370);
or U17651 (N_17651,N_15722,N_15814);
nor U17652 (N_17652,N_16943,N_15163);
nor U17653 (N_17653,N_15766,N_16782);
nand U17654 (N_17654,N_17462,N_17475);
and U17655 (N_17655,N_16783,N_17317);
nor U17656 (N_17656,N_16038,N_16023);
and U17657 (N_17657,N_16274,N_17464);
xor U17658 (N_17658,N_15642,N_15607);
xor U17659 (N_17659,N_16437,N_17163);
nand U17660 (N_17660,N_15177,N_17389);
nand U17661 (N_17661,N_15501,N_16343);
nand U17662 (N_17662,N_17038,N_15535);
nand U17663 (N_17663,N_17063,N_15023);
nor U17664 (N_17664,N_17091,N_15575);
or U17665 (N_17665,N_15971,N_15060);
and U17666 (N_17666,N_15865,N_16116);
nand U17667 (N_17667,N_15613,N_15266);
nor U17668 (N_17668,N_16319,N_16794);
and U17669 (N_17669,N_17455,N_16816);
and U17670 (N_17670,N_16238,N_16346);
nand U17671 (N_17671,N_15219,N_17180);
or U17672 (N_17672,N_16766,N_16480);
and U17673 (N_17673,N_15999,N_16348);
nand U17674 (N_17674,N_17391,N_15392);
and U17675 (N_17675,N_15960,N_15581);
xnor U17676 (N_17676,N_17242,N_16566);
and U17677 (N_17677,N_16257,N_17159);
xnor U17678 (N_17678,N_16713,N_17109);
or U17679 (N_17679,N_15625,N_16354);
or U17680 (N_17680,N_17360,N_16649);
or U17681 (N_17681,N_16693,N_16898);
and U17682 (N_17682,N_16607,N_15578);
or U17683 (N_17683,N_17080,N_17398);
or U17684 (N_17684,N_16152,N_16251);
nor U17685 (N_17685,N_15681,N_17405);
xor U17686 (N_17686,N_16685,N_16020);
nand U17687 (N_17687,N_17214,N_16235);
or U17688 (N_17688,N_15074,N_15977);
and U17689 (N_17689,N_15441,N_16965);
or U17690 (N_17690,N_16261,N_16626);
xor U17691 (N_17691,N_15443,N_16715);
xnor U17692 (N_17692,N_15486,N_16954);
nor U17693 (N_17693,N_17338,N_16281);
xnor U17694 (N_17694,N_15084,N_15704);
and U17695 (N_17695,N_16939,N_17418);
xor U17696 (N_17696,N_16171,N_17285);
or U17697 (N_17697,N_16486,N_15788);
or U17698 (N_17698,N_16641,N_17267);
or U17699 (N_17699,N_15841,N_16600);
nand U17700 (N_17700,N_17006,N_15323);
xor U17701 (N_17701,N_16318,N_16032);
or U17702 (N_17702,N_16145,N_17305);
xor U17703 (N_17703,N_16122,N_16174);
nand U17704 (N_17704,N_15626,N_16398);
nand U17705 (N_17705,N_15106,N_15803);
xor U17706 (N_17706,N_15789,N_15343);
and U17707 (N_17707,N_15513,N_15353);
xnor U17708 (N_17708,N_15384,N_15801);
and U17709 (N_17709,N_16275,N_15321);
and U17710 (N_17710,N_15471,N_15299);
xor U17711 (N_17711,N_16878,N_16556);
or U17712 (N_17712,N_15616,N_15958);
nor U17713 (N_17713,N_16638,N_17051);
and U17714 (N_17714,N_17002,N_16977);
nand U17715 (N_17715,N_17327,N_15341);
and U17716 (N_17716,N_15448,N_15889);
xor U17717 (N_17717,N_16519,N_15793);
and U17718 (N_17718,N_16008,N_16119);
and U17719 (N_17719,N_17431,N_15333);
nand U17720 (N_17720,N_16923,N_15256);
or U17721 (N_17721,N_15033,N_16762);
nand U17722 (N_17722,N_17482,N_15097);
and U17723 (N_17723,N_15252,N_15388);
nand U17724 (N_17724,N_16725,N_17131);
or U17725 (N_17725,N_17412,N_17486);
or U17726 (N_17726,N_15606,N_15758);
and U17727 (N_17727,N_16317,N_15938);
nor U17728 (N_17728,N_16864,N_15041);
nand U17729 (N_17729,N_15105,N_17272);
or U17730 (N_17730,N_16512,N_16956);
or U17731 (N_17731,N_15061,N_15895);
or U17732 (N_17732,N_17329,N_17034);
or U17733 (N_17733,N_15132,N_15249);
and U17734 (N_17734,N_15408,N_15885);
or U17735 (N_17735,N_15042,N_17499);
nand U17736 (N_17736,N_16942,N_16190);
nand U17737 (N_17737,N_17340,N_17492);
nor U17738 (N_17738,N_16005,N_16105);
xor U17739 (N_17739,N_16505,N_16324);
xor U17740 (N_17740,N_16962,N_17085);
xor U17741 (N_17741,N_16312,N_15718);
or U17742 (N_17742,N_15942,N_16026);
nor U17743 (N_17743,N_16201,N_15157);
nor U17744 (N_17744,N_15601,N_16579);
nor U17745 (N_17745,N_16525,N_17266);
nor U17746 (N_17746,N_15165,N_17358);
or U17747 (N_17747,N_16288,N_15858);
nor U17748 (N_17748,N_15227,N_16961);
nor U17749 (N_17749,N_16514,N_15638);
or U17750 (N_17750,N_17436,N_16680);
and U17751 (N_17751,N_16383,N_16788);
nor U17752 (N_17752,N_16823,N_15598);
nor U17753 (N_17753,N_15970,N_15734);
or U17754 (N_17754,N_16048,N_17355);
and U17755 (N_17755,N_16314,N_16449);
xor U17756 (N_17756,N_15747,N_17297);
nand U17757 (N_17757,N_15153,N_15319);
nor U17758 (N_17758,N_17254,N_15135);
and U17759 (N_17759,N_16371,N_17438);
or U17760 (N_17760,N_17273,N_17382);
or U17761 (N_17761,N_15530,N_17146);
xor U17762 (N_17762,N_17035,N_16889);
and U17763 (N_17763,N_16179,N_15586);
nand U17764 (N_17764,N_16738,N_16971);
xor U17765 (N_17765,N_15450,N_15641);
nand U17766 (N_17766,N_16000,N_15792);
nand U17767 (N_17767,N_17082,N_15700);
xnor U17768 (N_17768,N_15212,N_17478);
xor U17769 (N_17769,N_15685,N_16306);
nor U17770 (N_17770,N_17328,N_16709);
and U17771 (N_17771,N_17133,N_15200);
or U17772 (N_17772,N_16904,N_15494);
xnor U17773 (N_17773,N_17184,N_16734);
nand U17774 (N_17774,N_15468,N_15840);
and U17775 (N_17775,N_17298,N_15279);
nor U17776 (N_17776,N_15152,N_17156);
nor U17777 (N_17777,N_16866,N_15373);
and U17778 (N_17778,N_15125,N_15647);
nor U17779 (N_17779,N_17224,N_17162);
nor U17780 (N_17780,N_16948,N_16490);
nand U17781 (N_17781,N_15378,N_15102);
nand U17782 (N_17782,N_15962,N_16379);
or U17783 (N_17783,N_17077,N_16799);
xnor U17784 (N_17784,N_16913,N_17287);
nand U17785 (N_17785,N_15811,N_16474);
or U17786 (N_17786,N_15778,N_15190);
xor U17787 (N_17787,N_16220,N_15692);
xor U17788 (N_17788,N_15198,N_17359);
nor U17789 (N_17789,N_16417,N_15205);
nand U17790 (N_17790,N_17021,N_15141);
and U17791 (N_17791,N_16237,N_16265);
xor U17792 (N_17792,N_17350,N_16894);
nand U17793 (N_17793,N_16701,N_15176);
nor U17794 (N_17794,N_16389,N_17092);
nor U17795 (N_17795,N_17252,N_16402);
or U17796 (N_17796,N_15864,N_15917);
and U17797 (N_17797,N_16129,N_17090);
and U17798 (N_17798,N_17033,N_16749);
nor U17799 (N_17799,N_15317,N_16924);
or U17800 (N_17800,N_17247,N_15644);
or U17801 (N_17801,N_16330,N_17110);
and U17802 (N_17802,N_15079,N_15281);
xor U17803 (N_17803,N_16516,N_15804);
or U17804 (N_17804,N_16936,N_16506);
nor U17805 (N_17805,N_17017,N_16745);
xnor U17806 (N_17806,N_17458,N_17495);
and U17807 (N_17807,N_15093,N_15320);
or U17808 (N_17808,N_16590,N_16425);
nand U17809 (N_17809,N_15051,N_17466);
nor U17810 (N_17810,N_17228,N_16031);
nand U17811 (N_17811,N_16729,N_16926);
nor U17812 (N_17812,N_16905,N_15666);
nand U17813 (N_17813,N_17216,N_16349);
xnor U17814 (N_17814,N_17150,N_17351);
or U17815 (N_17815,N_15553,N_17422);
and U17816 (N_17816,N_15213,N_17256);
or U17817 (N_17817,N_16805,N_17045);
nand U17818 (N_17818,N_15843,N_16931);
nor U17819 (N_17819,N_15207,N_16430);
or U17820 (N_17820,N_15270,N_16757);
nor U17821 (N_17821,N_16072,N_15362);
or U17822 (N_17822,N_15142,N_15826);
nor U17823 (N_17823,N_16148,N_17240);
nor U17824 (N_17824,N_15974,N_16356);
or U17825 (N_17825,N_15175,N_15812);
nor U17826 (N_17826,N_16753,N_15701);
xor U17827 (N_17827,N_16045,N_16433);
xnor U17828 (N_17828,N_15275,N_15055);
nor U17829 (N_17829,N_15661,N_16121);
and U17830 (N_17830,N_16321,N_16044);
nand U17831 (N_17831,N_15107,N_16750);
or U17832 (N_17832,N_16986,N_16648);
and U17833 (N_17833,N_15324,N_16355);
nor U17834 (N_17834,N_16170,N_17457);
and U17835 (N_17835,N_15593,N_16880);
and U17836 (N_17836,N_15375,N_17313);
xnor U17837 (N_17837,N_15195,N_15807);
or U17838 (N_17838,N_16294,N_17075);
xnor U17839 (N_17839,N_15943,N_15532);
xor U17840 (N_17840,N_15117,N_16593);
xnor U17841 (N_17841,N_17460,N_17258);
xnor U17842 (N_17842,N_15907,N_16645);
xnor U17843 (N_17843,N_16922,N_15777);
xnor U17844 (N_17844,N_15478,N_15994);
or U17845 (N_17845,N_15355,N_17121);
nand U17846 (N_17846,N_16135,N_16707);
xnor U17847 (N_17847,N_16178,N_16021);
xor U17848 (N_17848,N_17292,N_15649);
nor U17849 (N_17849,N_15716,N_16067);
xnor U17850 (N_17850,N_17087,N_17116);
nand U17851 (N_17851,N_16029,N_16091);
and U17852 (N_17852,N_15550,N_17213);
and U17853 (N_17853,N_16655,N_15627);
nand U17854 (N_17854,N_16299,N_16921);
or U17855 (N_17855,N_15732,N_15487);
or U17856 (N_17856,N_15143,N_15512);
nand U17857 (N_17857,N_16457,N_17411);
and U17858 (N_17858,N_17068,N_15679);
and U17859 (N_17859,N_15364,N_15950);
nor U17860 (N_17860,N_15914,N_16778);
or U17861 (N_17861,N_15134,N_17118);
and U17862 (N_17862,N_15576,N_16256);
and U17863 (N_17863,N_15755,N_16606);
or U17864 (N_17864,N_16222,N_15447);
nand U17865 (N_17865,N_15984,N_16369);
nand U17866 (N_17866,N_17052,N_15991);
nor U17867 (N_17867,N_15306,N_17283);
or U17868 (N_17868,N_16559,N_15297);
nand U17869 (N_17869,N_17467,N_15172);
nor U17870 (N_17870,N_16110,N_15080);
nor U17871 (N_17871,N_15703,N_15401);
nand U17872 (N_17872,N_15431,N_15688);
or U17873 (N_17873,N_17199,N_17449);
xor U17874 (N_17874,N_17296,N_16156);
or U17875 (N_17875,N_15128,N_15352);
and U17876 (N_17876,N_15585,N_17354);
nand U17877 (N_17877,N_15762,N_16017);
and U17878 (N_17878,N_15796,N_15274);
and U17879 (N_17879,N_15870,N_16862);
nand U17880 (N_17880,N_15633,N_17208);
nor U17881 (N_17881,N_16071,N_17294);
or U17882 (N_17882,N_15561,N_15185);
nand U17883 (N_17883,N_16511,N_15590);
nor U17884 (N_17884,N_16166,N_16973);
xor U17885 (N_17885,N_16194,N_15706);
and U17886 (N_17886,N_15693,N_17440);
or U17887 (N_17887,N_16313,N_15571);
nor U17888 (N_17888,N_17126,N_16158);
xnor U17889 (N_17889,N_15288,N_15295);
nor U17890 (N_17890,N_17369,N_17388);
xnor U17891 (N_17891,N_15037,N_15538);
nand U17892 (N_17892,N_17059,N_15987);
or U17893 (N_17893,N_16436,N_16149);
xor U17894 (N_17894,N_15020,N_16557);
or U17895 (N_17895,N_15566,N_15837);
or U17896 (N_17896,N_15247,N_16405);
nor U17897 (N_17897,N_16475,N_16891);
nand U17898 (N_17898,N_15953,N_16874);
and U17899 (N_17899,N_16613,N_16438);
or U17900 (N_17900,N_17001,N_15307);
nand U17901 (N_17901,N_16994,N_16297);
or U17902 (N_17902,N_15669,N_15610);
nand U17903 (N_17903,N_15660,N_15502);
or U17904 (N_17904,N_15124,N_16700);
or U17905 (N_17905,N_16050,N_16375);
and U17906 (N_17906,N_15199,N_16822);
xor U17907 (N_17907,N_15952,N_17130);
nor U17908 (N_17908,N_16684,N_16376);
or U17909 (N_17909,N_15947,N_16770);
xnor U17910 (N_17910,N_15923,N_16654);
or U17911 (N_17911,N_15329,N_15754);
or U17912 (N_17912,N_16214,N_17374);
nand U17913 (N_17913,N_16789,N_15149);
xor U17914 (N_17914,N_16837,N_15912);
or U17915 (N_17915,N_15897,N_15096);
nand U17916 (N_17916,N_17117,N_15126);
nand U17917 (N_17917,N_15815,N_16207);
nor U17918 (N_17918,N_15186,N_17218);
or U17919 (N_17919,N_15903,N_15525);
and U17920 (N_17920,N_16532,N_15071);
or U17921 (N_17921,N_15052,N_16706);
xnor U17922 (N_17922,N_16102,N_15304);
xor U17923 (N_17923,N_15381,N_16997);
nor U17924 (N_17924,N_15058,N_16139);
and U17925 (N_17925,N_16065,N_15066);
and U17926 (N_17926,N_16501,N_16548);
and U17927 (N_17927,N_15597,N_15505);
and U17928 (N_17928,N_16596,N_16897);
and U17929 (N_17929,N_15340,N_16203);
or U17930 (N_17930,N_16813,N_16925);
or U17931 (N_17931,N_16711,N_17188);
nand U17932 (N_17932,N_16640,N_15549);
or U17933 (N_17933,N_15847,N_15150);
nor U17934 (N_17934,N_15739,N_15600);
nand U17935 (N_17935,N_15519,N_16581);
nand U17936 (N_17936,N_16338,N_17365);
or U17937 (N_17937,N_15565,N_15371);
and U17938 (N_17938,N_16598,N_17421);
or U17939 (N_17939,N_15940,N_16928);
or U17940 (N_17940,N_15531,N_16618);
xnor U17941 (N_17941,N_15933,N_16714);
nand U17942 (N_17942,N_16434,N_16195);
nor U17943 (N_17943,N_16670,N_16814);
nor U17944 (N_17944,N_15455,N_15735);
xnor U17945 (N_17945,N_15728,N_15534);
and U17946 (N_17946,N_15440,N_15982);
nand U17947 (N_17947,N_15181,N_17404);
xor U17948 (N_17948,N_17465,N_16455);
xor U17949 (N_17949,N_17145,N_17183);
xnor U17950 (N_17950,N_15078,N_16529);
or U17951 (N_17951,N_17450,N_16803);
nand U17952 (N_17952,N_15194,N_15560);
nor U17953 (N_17953,N_16047,N_17399);
nand U17954 (N_17954,N_15516,N_16993);
or U17955 (N_17955,N_16984,N_16817);
and U17956 (N_17956,N_16421,N_17217);
and U17957 (N_17957,N_17044,N_16487);
or U17958 (N_17958,N_15878,N_15621);
and U17959 (N_17959,N_16678,N_15072);
nor U17960 (N_17960,N_17489,N_16695);
nand U17961 (N_17961,N_16850,N_15753);
xnor U17962 (N_17962,N_16058,N_16528);
or U17963 (N_17963,N_15001,N_15312);
nand U17964 (N_17964,N_16760,N_15346);
and U17965 (N_17965,N_15523,N_16088);
and U17966 (N_17966,N_15363,N_16797);
nand U17967 (N_17967,N_15827,N_16196);
or U17968 (N_17968,N_15188,N_15000);
and U17969 (N_17969,N_15609,N_16401);
xor U17970 (N_17970,N_15664,N_16539);
and U17971 (N_17971,N_17004,N_16756);
and U17972 (N_17972,N_17342,N_16588);
or U17973 (N_17973,N_16886,N_17324);
or U17974 (N_17974,N_15904,N_16301);
and U17975 (N_17975,N_17414,N_16983);
and U17976 (N_17976,N_16025,N_17197);
nor U17977 (N_17977,N_15082,N_17057);
nand U17978 (N_17978,N_16530,N_16328);
xor U17979 (N_17979,N_15334,N_15076);
nand U17980 (N_17980,N_16176,N_15667);
nor U17981 (N_17981,N_16839,N_15540);
or U17982 (N_17982,N_16245,N_16646);
or U17983 (N_17983,N_16764,N_16743);
and U17984 (N_17984,N_17390,N_16834);
nor U17985 (N_17985,N_15764,N_17447);
xor U17986 (N_17986,N_17105,N_15546);
or U17987 (N_17987,N_15253,N_15310);
and U17988 (N_17988,N_16465,N_16408);
nor U17989 (N_17989,N_15283,N_15665);
and U17990 (N_17990,N_16053,N_15262);
nor U17991 (N_17991,N_15828,N_15239);
nand U17992 (N_17992,N_16533,N_15202);
or U17993 (N_17993,N_15174,N_15913);
and U17994 (N_17994,N_15745,N_15013);
or U17995 (N_17995,N_16615,N_15838);
nor U17996 (N_17996,N_16974,N_15951);
and U17997 (N_17997,N_15491,N_16114);
and U17998 (N_17998,N_15302,N_17452);
and U17999 (N_17999,N_17381,N_15336);
xnor U18000 (N_18000,N_15910,N_16976);
nand U18001 (N_18001,N_16335,N_16639);
nor U18002 (N_18002,N_15608,N_16271);
or U18003 (N_18003,N_15457,N_15030);
and U18004 (N_18004,N_15127,N_15813);
nand U18005 (N_18005,N_16087,N_15308);
nand U18006 (N_18006,N_16751,N_15508);
nand U18007 (N_18007,N_16167,N_17178);
nand U18008 (N_18008,N_15278,N_17149);
and U18009 (N_18009,N_15620,N_15386);
and U18010 (N_18010,N_15488,N_16471);
nor U18011 (N_18011,N_15853,N_17311);
or U18012 (N_18012,N_16409,N_16382);
xor U18013 (N_18013,N_15316,N_17172);
or U18014 (N_18014,N_15678,N_17282);
or U18015 (N_18015,N_16951,N_17187);
and U18016 (N_18016,N_15467,N_16543);
or U18017 (N_18017,N_16848,N_15573);
and U18018 (N_18018,N_16812,N_16981);
or U18019 (N_18019,N_15780,N_16443);
xor U18020 (N_18020,N_16347,N_16716);
nor U18021 (N_18021,N_16629,N_16541);
xor U18022 (N_18022,N_15231,N_17018);
nor U18023 (N_18023,N_15835,N_15115);
nor U18024 (N_18024,N_17198,N_16427);
nand U18025 (N_18025,N_15783,N_16286);
xor U18026 (N_18026,N_17301,N_15551);
xor U18027 (N_18027,N_17334,N_17401);
nand U18028 (N_18028,N_15927,N_16571);
xnor U18029 (N_18029,N_17441,N_16442);
and U18030 (N_18030,N_16002,N_15103);
xnor U18031 (N_18031,N_17277,N_17168);
xor U18032 (N_18032,N_16554,N_17097);
or U18033 (N_18033,N_16164,N_16724);
or U18034 (N_18034,N_16555,N_15682);
nor U18035 (N_18035,N_16741,N_16054);
and U18036 (N_18036,N_17410,N_17205);
nand U18037 (N_18037,N_16439,N_15861);
and U18038 (N_18038,N_16836,N_15817);
xor U18039 (N_18039,N_16240,N_15255);
nor U18040 (N_18040,N_17241,N_15291);
xnor U18041 (N_18041,N_15372,N_16500);
nand U18042 (N_18042,N_16051,N_15110);
nor U18043 (N_18043,N_16466,N_16070);
xnor U18044 (N_18044,N_16209,N_15463);
nor U18045 (N_18045,N_16049,N_15475);
nor U18046 (N_18046,N_15612,N_16063);
nor U18047 (N_18047,N_16811,N_15717);
and U18048 (N_18048,N_15872,N_16394);
and U18049 (N_18049,N_17335,N_15330);
or U18050 (N_18050,N_15043,N_16022);
or U18051 (N_18051,N_17276,N_15672);
or U18052 (N_18052,N_15242,N_16413);
xnor U18053 (N_18053,N_16429,N_17028);
nor U18054 (N_18054,N_16128,N_15369);
or U18055 (N_18055,N_15028,N_15092);
and U18056 (N_18056,N_15645,N_15854);
nand U18057 (N_18057,N_15116,N_15047);
nand U18058 (N_18058,N_16801,N_17009);
xnor U18059 (N_18059,N_16100,N_15918);
nand U18060 (N_18060,N_16605,N_17269);
xnor U18061 (N_18061,N_17362,N_17229);
nand U18062 (N_18062,N_16852,N_16192);
or U18063 (N_18063,N_17419,N_17177);
nand U18064 (N_18064,N_15640,N_15158);
nor U18065 (N_18065,N_16573,N_15624);
and U18066 (N_18066,N_15365,N_15760);
nand U18067 (N_18067,N_16079,N_16996);
or U18068 (N_18068,N_15635,N_17023);
xnor U18069 (N_18069,N_16226,N_16918);
and U18070 (N_18070,N_16147,N_15035);
or U18071 (N_18071,N_15825,N_15429);
or U18072 (N_18072,N_15623,N_17207);
and U18073 (N_18073,N_15738,N_15121);
xnor U18074 (N_18074,N_15629,N_16247);
and U18075 (N_18075,N_15472,N_17013);
nand U18076 (N_18076,N_16968,N_15122);
and U18077 (N_18077,N_15930,N_17008);
and U18078 (N_18078,N_16123,N_16177);
nor U18079 (N_18079,N_17300,N_16907);
or U18080 (N_18080,N_15257,N_16873);
or U18081 (N_18081,N_15964,N_15900);
xnor U18082 (N_18082,N_15710,N_16987);
or U18083 (N_18083,N_16830,N_15995);
or U18084 (N_18084,N_15420,N_16576);
and U18085 (N_18085,N_16503,N_17341);
xnor U18086 (N_18086,N_17053,N_15877);
or U18087 (N_18087,N_15003,N_17005);
nand U18088 (N_18088,N_16513,N_17086);
nand U18089 (N_18089,N_16902,N_15053);
nor U18090 (N_18090,N_15415,N_16585);
nand U18091 (N_18091,N_16352,N_17403);
nor U18092 (N_18092,N_15892,N_15325);
nor U18093 (N_18093,N_15752,N_16208);
xor U18094 (N_18094,N_15775,N_15170);
nand U18095 (N_18095,N_15965,N_16246);
nor U18096 (N_18096,N_16932,N_16689);
nor U18097 (N_18097,N_15018,N_15887);
and U18098 (N_18098,N_16771,N_16719);
xnor U18099 (N_18099,N_17106,N_16908);
nor U18100 (N_18100,N_15397,N_16899);
or U18101 (N_18101,N_16189,N_15954);
nor U18102 (N_18102,N_15021,N_16334);
nor U18103 (N_18103,N_15684,N_15138);
nor U18104 (N_18104,N_15554,N_16563);
or U18105 (N_18105,N_15216,N_15810);
xnor U18106 (N_18106,N_15756,N_16508);
nand U18107 (N_18107,N_16269,N_16315);
nor U18108 (N_18108,N_15087,N_16577);
xnor U18109 (N_18109,N_16509,N_16125);
and U18110 (N_18110,N_15411,N_15968);
and U18111 (N_18111,N_16643,N_16033);
or U18112 (N_18112,N_15002,N_15691);
and U18113 (N_18113,N_16173,N_15054);
and U18114 (N_18114,N_16153,N_15799);
xor U18115 (N_18115,N_15869,N_17194);
nor U18116 (N_18116,N_15805,N_16731);
and U18117 (N_18117,N_16710,N_15599);
nor U18118 (N_18118,N_17158,N_17429);
or U18119 (N_18119,N_15785,N_16252);
nor U18120 (N_18120,N_16569,N_15476);
or U18121 (N_18121,N_15757,N_16526);
and U18122 (N_18122,N_16963,N_17043);
or U18123 (N_18123,N_15461,N_16476);
nand U18124 (N_18124,N_16491,N_15347);
and U18125 (N_18125,N_17115,N_17046);
nor U18126 (N_18126,N_16041,N_15026);
or U18127 (N_18127,N_15211,N_16211);
or U18128 (N_18128,N_15875,N_15770);
xnor U18129 (N_18129,N_16634,N_15705);
or U18130 (N_18130,N_15636,N_16212);
xor U18131 (N_18131,N_16527,N_16773);
and U18132 (N_18132,N_16858,N_16747);
nor U18133 (N_18133,N_17326,N_16042);
or U18134 (N_18134,N_16964,N_17417);
nand U18135 (N_18135,N_17226,N_15267);
or U18136 (N_18136,N_15670,N_15015);
or U18137 (N_18137,N_16291,N_16151);
xor U18138 (N_18138,N_15311,N_15524);
and U18139 (N_18139,N_16239,N_16856);
or U18140 (N_18140,N_15484,N_15577);
and U18141 (N_18141,N_16726,N_16378);
nor U18142 (N_18142,N_16775,N_16326);
xnor U18143 (N_18143,N_16632,N_17020);
and U18144 (N_18144,N_17396,N_16746);
nand U18145 (N_18145,N_15860,N_16946);
nand U18146 (N_18146,N_16117,N_15973);
nor U18147 (N_18147,N_15526,N_15277);
nand U18148 (N_18148,N_16888,N_17120);
xor U18149 (N_18149,N_16131,N_15574);
and U18150 (N_18150,N_17386,N_15740);
and U18151 (N_18151,N_16625,N_16483);
or U18152 (N_18152,N_15077,N_15111);
or U18153 (N_18153,N_16325,N_15820);
xor U18154 (N_18154,N_15394,N_16454);
and U18155 (N_18155,N_17275,N_15034);
and U18156 (N_18156,N_17375,N_16293);
nor U18157 (N_18157,N_16785,N_16277);
nand U18158 (N_18158,N_16146,N_17420);
nor U18159 (N_18159,N_15208,N_16582);
nor U18160 (N_18160,N_15201,N_16162);
nor U18161 (N_18161,N_16861,N_17409);
or U18162 (N_18162,N_15309,N_15541);
or U18163 (N_18163,N_15983,N_16855);
and U18164 (N_18164,N_15781,N_16672);
and U18165 (N_18165,N_17303,N_15883);
and U18166 (N_18166,N_15751,N_16630);
or U18167 (N_18167,N_16287,N_15955);
or U18168 (N_18168,N_17125,N_15480);
and U18169 (N_18169,N_16958,N_17237);
or U18170 (N_18170,N_16134,N_16081);
nor U18171 (N_18171,N_17246,N_16340);
or U18172 (N_18172,N_17181,N_16360);
and U18173 (N_18173,N_17434,N_16407);
and U18174 (N_18174,N_15477,N_15133);
nor U18175 (N_18175,N_15059,N_16161);
xor U18176 (N_18176,N_16650,N_15161);
or U18177 (N_18177,N_15428,N_15243);
xnor U18178 (N_18178,N_16887,N_15421);
nor U18179 (N_18179,N_16193,N_17485);
nand U18180 (N_18180,N_16795,N_17236);
nand U18181 (N_18181,N_15919,N_16759);
or U18182 (N_18182,N_17084,N_15619);
nand U18183 (N_18183,N_17472,N_16884);
nor U18184 (N_18184,N_16831,N_15773);
nand U18185 (N_18185,N_16266,N_17425);
and U18186 (N_18186,N_16909,N_15331);
and U18187 (N_18187,N_16228,N_16883);
nor U18188 (N_18188,N_17384,N_15424);
nand U18189 (N_18189,N_16083,N_15859);
nand U18190 (N_18190,N_15271,N_15979);
nand U18191 (N_18191,N_16198,N_15648);
xor U18192 (N_18192,N_17192,N_15655);
nand U18193 (N_18193,N_15432,N_15067);
nor U18194 (N_18194,N_15410,N_15857);
and U18195 (N_18195,N_15235,N_16096);
nor U18196 (N_18196,N_15009,N_15404);
or U18197 (N_18197,N_16037,N_15496);
xor U18198 (N_18198,N_15357,N_15719);
and U18199 (N_18199,N_15354,N_16744);
nand U18200 (N_18200,N_16113,N_15091);
nand U18201 (N_18201,N_15050,N_15434);
nand U18202 (N_18202,N_16635,N_16221);
or U18203 (N_18203,N_15768,N_16272);
nand U18204 (N_18204,N_17175,N_15436);
nand U18205 (N_18205,N_16479,N_15011);
or U18206 (N_18206,N_15967,N_16404);
nor U18207 (N_18207,N_16076,N_16035);
xor U18208 (N_18208,N_15708,N_15136);
nand U18209 (N_18209,N_15795,N_15438);
nand U18210 (N_18210,N_16666,N_17395);
xnor U18211 (N_18211,N_16959,N_15567);
or U18212 (N_18212,N_15423,N_17474);
xor U18213 (N_18213,N_15926,N_16901);
or U18214 (N_18214,N_15587,N_16493);
or U18215 (N_18215,N_15146,N_15131);
or U18216 (N_18216,N_16333,N_16636);
xor U18217 (N_18217,N_17190,N_15215);
nand U18218 (N_18218,N_15412,N_15668);
nor U18219 (N_18219,N_16912,N_15650);
nand U18220 (N_18220,N_17227,N_15383);
nand U18221 (N_18221,N_16236,N_15765);
and U18222 (N_18222,N_15068,N_17094);
nand U18223 (N_18223,N_16944,N_16084);
xnor U18224 (N_18224,N_15657,N_16388);
nor U18225 (N_18225,N_16098,N_15975);
and U18226 (N_18226,N_17137,N_15698);
xnor U18227 (N_18227,N_16521,N_16767);
xor U18228 (N_18228,N_17377,N_17325);
and U18229 (N_18229,N_15493,N_15173);
or U18230 (N_18230,N_16982,N_15873);
nor U18231 (N_18231,N_17308,N_15806);
and U18232 (N_18232,N_17219,N_16447);
nand U18233 (N_18233,N_16007,N_15075);
nand U18234 (N_18234,N_16219,N_16735);
nor U18235 (N_18235,N_16601,N_16080);
nor U18236 (N_18236,N_15736,N_15823);
nor U18237 (N_18237,N_17261,N_17244);
or U18238 (N_18238,N_16099,N_16720);
and U18239 (N_18239,N_15862,N_15866);
and U18240 (N_18240,N_15025,N_16518);
nand U18241 (N_18241,N_17200,N_15948);
nand U18242 (N_18242,N_17071,N_16769);
or U18243 (N_18243,N_17372,N_16733);
xnor U18244 (N_18244,N_16403,N_16304);
xor U18245 (N_18245,N_16280,N_16798);
xnor U18246 (N_18246,N_15709,N_16001);
nor U18247 (N_18247,N_16586,N_15966);
or U18248 (N_18248,N_17047,N_16819);
xor U18249 (N_18249,N_15602,N_16686);
xor U18250 (N_18250,N_15240,N_15533);
nor U18251 (N_18251,N_17036,N_15902);
nand U18252 (N_18252,N_16181,N_15293);
xor U18253 (N_18253,N_16399,N_16820);
nand U18254 (N_18254,N_15269,N_15921);
nor U18255 (N_18255,N_16547,N_15435);
and U18256 (N_18256,N_15742,N_15632);
nor U18257 (N_18257,N_16270,N_15332);
nand U18258 (N_18258,N_17107,N_15639);
or U18259 (N_18259,N_17127,N_15374);
nand U18260 (N_18260,N_15809,N_16302);
and U18261 (N_18261,N_15871,N_15993);
xor U18262 (N_18262,N_15726,N_15856);
or U18263 (N_18263,N_15929,N_15759);
or U18264 (N_18264,N_16464,N_15771);
nor U18265 (N_18265,N_16742,N_16242);
xnor U18266 (N_18266,N_15528,N_16273);
xor U18267 (N_18267,N_16337,N_15680);
nor U18268 (N_18268,N_16777,N_15963);
nand U18269 (N_18269,N_16412,N_17442);
or U18270 (N_18270,N_16004,N_16642);
nor U18271 (N_18271,N_17173,N_16717);
xnor U18272 (N_18272,N_16497,N_15939);
xor U18273 (N_18273,N_16914,N_15615);
or U18274 (N_18274,N_16851,N_16510);
and U18275 (N_18275,N_15007,N_15382);
xnor U18276 (N_18276,N_17238,N_15039);
or U18277 (N_18277,N_16101,N_17069);
nand U18278 (N_18278,N_15715,N_17152);
xor U18279 (N_18279,N_16089,N_17361);
xor U18280 (N_18280,N_16584,N_16790);
xor U18281 (N_18281,N_15104,N_15744);
or U18282 (N_18282,N_15934,N_16838);
and U18283 (N_18283,N_17031,N_17012);
nand U18284 (N_18284,N_17170,N_15981);
and U18285 (N_18285,N_16900,N_16524);
or U18286 (N_18286,N_16892,N_15769);
nor U18287 (N_18287,N_16481,N_17295);
or U18288 (N_18288,N_15469,N_15818);
nor U18289 (N_18289,N_15250,N_15694);
or U18290 (N_18290,N_16120,N_15834);
nor U18291 (N_18291,N_16183,N_15822);
or U18292 (N_18292,N_15403,N_16570);
or U18293 (N_18293,N_17223,N_15073);
and U18294 (N_18294,N_16496,N_17448);
or U18295 (N_18295,N_16540,N_16656);
or U18296 (N_18296,N_17193,N_16191);
or U18297 (N_18297,N_15784,N_15406);
and U18298 (N_18298,N_16456,N_15891);
nand U18299 (N_18299,N_15842,N_16204);
nand U18300 (N_18300,N_15130,N_15989);
nand U18301 (N_18301,N_15588,N_16804);
or U18302 (N_18302,N_15998,N_17397);
or U18303 (N_18303,N_15481,N_16560);
or U18304 (N_18304,N_16353,N_17070);
nand U18305 (N_18305,N_16927,N_16276);
nand U18306 (N_18306,N_16345,N_15065);
or U18307 (N_18307,N_17233,N_16978);
and U18308 (N_18308,N_16327,N_16824);
nor U18309 (N_18309,N_17378,N_15580);
nand U18310 (N_18310,N_17011,N_16910);
and U18311 (N_18311,N_16546,N_16662);
or U18312 (N_18312,N_16248,N_16657);
or U18313 (N_18313,N_15460,N_17076);
nand U18314 (N_18314,N_15746,N_17289);
and U18315 (N_18315,N_15687,N_15453);
or U18316 (N_18316,N_16872,N_16937);
or U18317 (N_18317,N_16292,N_16633);
nand U18318 (N_18318,N_15881,N_16622);
xnor U18319 (N_18319,N_17102,N_15303);
and U18320 (N_18320,N_16890,N_17483);
nand U18321 (N_18321,N_16755,N_16300);
xnor U18322 (N_18322,N_16308,N_15562);
nor U18323 (N_18323,N_16268,N_15064);
or U18324 (N_18324,N_15482,N_16133);
nor U18325 (N_18325,N_16138,N_16199);
nor U18326 (N_18326,N_17333,N_15686);
and U18327 (N_18327,N_15189,N_16841);
nor U18328 (N_18328,N_16915,N_16132);
nor U18329 (N_18329,N_16077,N_17435);
or U18330 (N_18330,N_16336,N_15399);
xor U18331 (N_18331,N_15422,N_15289);
xor U18332 (N_18332,N_15376,N_16027);
nand U18333 (N_18333,N_15010,N_16718);
and U18334 (N_18334,N_17014,N_15425);
or U18335 (N_18335,N_17322,N_15696);
and U18336 (N_18336,N_17470,N_16661);
nor U18337 (N_18337,N_16776,N_16107);
xor U18338 (N_18338,N_17330,N_15005);
or U18339 (N_18339,N_16784,N_16796);
nor U18340 (N_18340,N_16969,N_16316);
nor U18341 (N_18341,N_15099,N_16339);
or U18342 (N_18342,N_17424,N_15920);
nand U18343 (N_18343,N_16673,N_16322);
and U18344 (N_18344,N_16295,N_16692);
and U18345 (N_18345,N_15572,N_17185);
xor U18346 (N_18346,N_16163,N_15167);
nand U18347 (N_18347,N_17128,N_16704);
or U18348 (N_18348,N_17095,N_15402);
nor U18349 (N_18349,N_15287,N_15816);
xnor U18350 (N_18350,N_15391,N_16073);
nand U18351 (N_18351,N_16411,N_15433);
nand U18352 (N_18352,N_15906,N_17461);
nand U18353 (N_18353,N_16350,N_16450);
and U18354 (N_18354,N_15154,N_16832);
xnor U18355 (N_18355,N_16460,N_15725);
nand U18356 (N_18356,N_15924,N_16972);
and U18357 (N_18357,N_16840,N_15582);
and U18358 (N_18358,N_15209,N_15344);
nor U18359 (N_18359,N_16279,N_16682);
xor U18360 (N_18360,N_15563,N_16458);
or U18361 (N_18361,N_17032,N_17139);
xnor U18362 (N_18362,N_15925,N_16342);
nor U18363 (N_18363,N_15144,N_16934);
nor U18364 (N_18364,N_15254,N_16833);
and U18365 (N_18365,N_16418,N_15886);
nand U18366 (N_18366,N_15675,N_15458);
and U18367 (N_18367,N_16130,N_16472);
nand U18368 (N_18368,N_15114,N_15348);
or U18369 (N_18369,N_17407,N_17367);
xnor U18370 (N_18370,N_16668,N_16938);
or U18371 (N_18371,N_16064,N_16078);
nor U18372 (N_18372,N_15282,N_15569);
nor U18373 (N_18373,N_15527,N_16420);
nor U18374 (N_18374,N_16580,N_17468);
xnor U18375 (N_18375,N_16534,N_17490);
nor U18376 (N_18376,N_16392,N_15786);
nor U18377 (N_18377,N_17079,N_16469);
and U18378 (N_18378,N_17025,N_15637);
nor U18379 (N_18379,N_15454,N_16967);
xnor U18380 (N_18380,N_16876,N_17167);
and U18381 (N_18381,N_16599,N_17473);
nand U18382 (N_18382,N_16761,N_15345);
xnor U18383 (N_18383,N_15452,N_16461);
or U18384 (N_18384,N_16574,N_17157);
and U18385 (N_18385,N_17320,N_16216);
or U18386 (N_18386,N_17235,N_15916);
xnor U18387 (N_18387,N_16305,N_16703);
xor U18388 (N_18388,N_17058,N_15537);
and U18389 (N_18389,N_15492,N_16232);
or U18390 (N_18390,N_15868,N_16052);
xor U18391 (N_18391,N_16568,N_16444);
nor U18392 (N_18392,N_15296,N_15430);
xnor U18393 (N_18393,N_15507,N_16014);
and U18394 (N_18394,N_17321,N_16488);
xnor U18395 (N_18395,N_16810,N_17039);
and U18396 (N_18396,N_17212,N_16966);
xor U18397 (N_18397,N_16141,N_17364);
nand U18398 (N_18398,N_15713,N_17463);
nand U18399 (N_18399,N_15656,N_15479);
or U18400 (N_18400,N_16542,N_15707);
and U18401 (N_18401,N_15197,N_16426);
and U18402 (N_18402,N_17232,N_15497);
xor U18403 (N_18403,N_15674,N_16202);
nand U18404 (N_18404,N_15223,N_16024);
xor U18405 (N_18405,N_16664,N_15019);
xnor U18406 (N_18406,N_16370,N_15888);
and U18407 (N_18407,N_16628,N_17346);
xnor U18408 (N_18408,N_15846,N_15714);
nor U18409 (N_18409,N_16230,N_15276);
xnor U18410 (N_18410,N_16871,N_16616);
or U18411 (N_18411,N_15978,N_16895);
nand U18412 (N_18412,N_16842,N_15673);
nand U18413 (N_18413,N_17332,N_17204);
nand U18414 (N_18414,N_16911,N_16188);
and U18415 (N_18415,N_15339,N_15145);
or U18416 (N_18416,N_17376,N_16143);
and U18417 (N_18417,N_17498,N_15720);
nor U18418 (N_18418,N_16545,N_17310);
xnor U18419 (N_18419,N_16991,N_16126);
or U18420 (N_18420,N_15044,N_15451);
or U18421 (N_18421,N_16103,N_16229);
xnor U18422 (N_18422,N_16587,N_15631);
xnor U18423 (N_18423,N_17010,N_15852);
nor U18424 (N_18424,N_15238,N_17385);
nor U18425 (N_18425,N_15204,N_15268);
nor U18426 (N_18426,N_17402,N_15596);
nand U18427 (N_18427,N_15518,N_16473);
xor U18428 (N_18428,N_17113,N_17366);
nand U18429 (N_18429,N_15570,N_15225);
or U18430 (N_18430,N_17257,N_15368);
or U18431 (N_18431,N_17373,N_15794);
nor U18432 (N_18432,N_15396,N_15658);
xnor U18433 (N_18433,N_16361,N_15915);
and U18434 (N_18434,N_15045,N_16538);
and U18435 (N_18435,N_15509,N_15118);
nor U18436 (N_18436,N_15400,N_15290);
xor U18437 (N_18437,N_16652,N_16857);
nand U18438 (N_18438,N_15536,N_15483);
and U18439 (N_18439,N_16980,N_16552);
or U18440 (N_18440,N_16323,N_17108);
nor U18441 (N_18441,N_17182,N_17083);
xnor U18442 (N_18442,N_16154,N_15821);
nand U18443 (N_18443,N_16415,N_16722);
and U18444 (N_18444,N_16393,N_15556);
and U18445 (N_18445,N_17141,N_15683);
or U18446 (N_18446,N_17406,N_16030);
nor U18447 (N_18447,N_16752,N_15500);
and U18448 (N_18448,N_16780,N_16723);
nor U18449 (N_18449,N_17302,N_17393);
nor U18450 (N_18450,N_15095,N_15248);
or U18451 (N_18451,N_17211,N_16517);
xnor U18452 (N_18452,N_16422,N_16036);
or U18453 (N_18453,N_15221,N_15465);
or U18454 (N_18454,N_15520,N_15056);
or U18455 (N_18455,N_15120,N_15779);
nor U18456 (N_18456,N_15763,N_15729);
and U18457 (N_18457,N_15733,N_17201);
and U18458 (N_18458,N_16424,N_15322);
or U18459 (N_18459,N_15081,N_15555);
nor U18460 (N_18460,N_17100,N_16311);
and U18461 (N_18461,N_15617,N_17491);
nor U18462 (N_18462,N_15584,N_16108);
and U18463 (N_18463,N_16597,N_15611);
xor U18464 (N_18464,N_16435,N_16453);
xor U18465 (N_18465,N_17066,N_16589);
xor U18466 (N_18466,N_15591,N_17394);
nand U18467 (N_18467,N_17245,N_15183);
and U18468 (N_18468,N_15437,N_16069);
xnor U18469 (N_18469,N_16223,N_16055);
and U18470 (N_18470,N_15552,N_16885);
nor U18471 (N_18471,N_15456,N_17169);
nor U18472 (N_18472,N_15358,N_16610);
xnor U18473 (N_18473,N_17099,N_16384);
and U18474 (N_18474,N_16115,N_15305);
nand U18475 (N_18475,N_16440,N_15089);
xnor U18476 (N_18476,N_17048,N_15218);
nand U18477 (N_18477,N_15265,N_16094);
or U18478 (N_18478,N_15776,N_15884);
or U18479 (N_18479,N_15379,N_16893);
xor U18480 (N_18480,N_15761,N_16331);
nand U18481 (N_18481,N_15772,N_16515);
nor U18482 (N_18482,N_15594,N_16564);
xor U18483 (N_18483,N_16807,N_16567);
xor U18484 (N_18484,N_17337,N_16647);
nor U18485 (N_18485,N_17134,N_15390);
and U18486 (N_18486,N_16309,N_15874);
nand U18487 (N_18487,N_16827,N_15690);
nand U18488 (N_18488,N_15992,N_16708);
nand U18489 (N_18489,N_15997,N_17348);
and U18490 (N_18490,N_17209,N_15911);
or U18491 (N_18491,N_15342,N_17186);
xor U18492 (N_18492,N_15543,N_15473);
and U18493 (N_18493,N_16419,N_17215);
nand U18494 (N_18494,N_16298,N_15931);
xnor U18495 (N_18495,N_17060,N_16507);
nand U18496 (N_18496,N_15314,N_16169);
nor U18497 (N_18497,N_16180,N_16395);
xnor U18498 (N_18498,N_15651,N_15836);
xnor U18499 (N_18499,N_16367,N_15260);
and U18500 (N_18500,N_16621,N_16385);
xnor U18501 (N_18501,N_16787,N_16748);
nor U18502 (N_18502,N_17280,N_15361);
or U18503 (N_18503,N_16234,N_16060);
and U18504 (N_18504,N_17349,N_15178);
xor U18505 (N_18505,N_17307,N_15844);
xnor U18506 (N_18506,N_15832,N_16727);
or U18507 (N_18507,N_16879,N_15671);
and U18508 (N_18508,N_15945,N_16663);
or U18509 (N_18509,N_16947,N_15800);
xnor U18510 (N_18510,N_17225,N_15272);
and U18511 (N_18511,N_17042,N_15184);
and U18512 (N_18512,N_17387,N_17352);
or U18513 (N_18513,N_16772,N_15180);
nor U18514 (N_18514,N_15168,N_17323);
and U18515 (N_18515,N_16906,N_15360);
and U18516 (N_18516,N_16536,N_17078);
xnor U18517 (N_18517,N_15935,N_15499);
xnor U18518 (N_18518,N_15802,N_17161);
and U18519 (N_18519,N_15503,N_16019);
or U18520 (N_18520,N_15444,N_17456);
xor U18521 (N_18521,N_17027,N_15972);
nand U18522 (N_18522,N_15957,N_15750);
and U18523 (N_18523,N_16818,N_17210);
and U18524 (N_18524,N_17067,N_17484);
nand U18525 (N_18525,N_16086,N_16225);
xnor U18526 (N_18526,N_15038,N_15898);
and U18527 (N_18527,N_17356,N_16068);
nor U18528 (N_18528,N_17259,N_15098);
or U18529 (N_18529,N_15049,N_15232);
xor U18530 (N_18530,N_16284,N_15366);
xor U18531 (N_18531,N_17459,N_16231);
nor U18532 (N_18532,N_16603,N_15169);
and U18533 (N_18533,N_15731,N_17493);
nor U18534 (N_18534,N_15790,N_17428);
xor U18535 (N_18535,N_15767,N_17073);
nor U18536 (N_18536,N_15712,N_16062);
nand U18537 (N_18537,N_17000,N_16303);
nand U18538 (N_18538,N_15016,N_15464);
nand U18539 (N_18539,N_15220,N_16218);
xor U18540 (N_18540,N_17288,N_17469);
or U18541 (N_18541,N_16690,N_17392);
or U18542 (N_18542,N_16307,N_16011);
xnor U18543 (N_18543,N_15980,N_16849);
xor U18544 (N_18544,N_16737,N_16489);
and U18545 (N_18545,N_16310,N_17050);
and U18546 (N_18546,N_16016,N_16676);
and U18547 (N_18547,N_16999,N_15749);
and U18548 (N_18548,N_17132,N_15879);
and U18549 (N_18549,N_15959,N_17347);
xnor U18550 (N_18550,N_16825,N_16945);
nand U18551 (N_18551,N_16843,N_16815);
and U18552 (N_18552,N_16877,N_17007);
nor U18553 (N_18553,N_15985,N_17437);
and U18554 (N_18554,N_17318,N_17234);
nor U18555 (N_18555,N_16736,N_16875);
and U18556 (N_18556,N_16013,N_16092);
or U18557 (N_18557,N_16462,N_16792);
nand U18558 (N_18558,N_15937,N_17413);
nand U18559 (N_18559,N_15192,N_16988);
xor U18560 (N_18560,N_16494,N_16320);
nor U18561 (N_18561,N_17142,N_15119);
and U18562 (N_18562,N_16558,N_15446);
nand U18563 (N_18563,N_15653,N_16498);
and U18564 (N_18564,N_15787,N_16644);
nand U18565 (N_18565,N_15417,N_16809);
nand U18566 (N_18566,N_16362,N_16157);
or U18567 (N_18567,N_15063,N_17143);
or U18568 (N_18568,N_15148,N_16739);
nand U18569 (N_18569,N_17344,N_16463);
nor U18570 (N_18570,N_16406,N_16358);
nor U18571 (N_18571,N_15737,N_15351);
nor U18572 (N_18572,N_17253,N_17423);
or U18573 (N_18573,N_16696,N_16012);
nand U18574 (N_18574,N_16903,N_16351);
or U18575 (N_18575,N_16651,N_16609);
xnor U18576 (N_18576,N_16989,N_17015);
and U18577 (N_18577,N_17206,N_16186);
nor U18578 (N_18578,N_16975,N_17290);
and U18579 (N_18579,N_15489,N_15085);
or U18580 (N_18580,N_15416,N_16675);
and U18581 (N_18581,N_16387,N_15882);
xnor U18582 (N_18582,N_16953,N_15442);
or U18583 (N_18583,N_17380,N_16259);
or U18584 (N_18584,N_15230,N_15797);
nand U18585 (N_18585,N_16619,N_15748);
or U18586 (N_18586,N_15377,N_15086);
nand U18587 (N_18587,N_15004,N_16583);
or U18588 (N_18588,N_16368,N_16363);
nor U18589 (N_18589,N_17230,N_17479);
and U18590 (N_18590,N_15798,N_16391);
nand U18591 (N_18591,N_16200,N_17088);
xor U18592 (N_18592,N_16806,N_16845);
or U18593 (N_18593,N_17165,N_16624);
and U18594 (N_18594,N_15880,N_15294);
nor U18595 (N_18595,N_16740,N_15466);
xnor U18596 (N_18596,N_15229,N_16390);
nand U18597 (N_18597,N_17314,N_15462);
and U18598 (N_18598,N_15300,N_16916);
and U18599 (N_18599,N_15236,N_16227);
xor U18600 (N_18600,N_17315,N_15356);
nand U18601 (N_18601,N_16620,N_16332);
nand U18602 (N_18602,N_16059,N_16677);
nor U18603 (N_18603,N_17135,N_15529);
or U18604 (N_18604,N_17271,N_16283);
or U18605 (N_18605,N_15337,N_15155);
xor U18606 (N_18606,N_15233,N_16572);
or U18607 (N_18607,N_17016,N_17055);
and U18608 (N_18608,N_15689,N_15261);
nand U18609 (N_18609,N_15677,N_15515);
or U18610 (N_18610,N_15315,N_17278);
or U18611 (N_18611,N_16728,N_16168);
nand U18612 (N_18612,N_17026,N_17072);
nand U18613 (N_18613,N_16868,N_16263);
nor U18614 (N_18614,N_16296,N_16702);
nand U18615 (N_18615,N_16470,N_15774);
nor U18616 (N_18616,N_17444,N_16955);
or U18617 (N_18617,N_17155,N_15070);
nand U18618 (N_18618,N_17160,N_15014);
nand U18619 (N_18619,N_16377,N_16919);
nor U18620 (N_18620,N_16499,N_17054);
xnor U18621 (N_18621,N_15628,N_15318);
xor U18622 (N_18622,N_15259,N_17019);
xor U18623 (N_18623,N_17400,N_16213);
nand U18624 (N_18624,N_15036,N_15506);
or U18625 (N_18625,N_15504,N_16445);
or U18626 (N_18626,N_17415,N_15196);
xnor U18627 (N_18627,N_17279,N_17262);
nor U18628 (N_18628,N_15583,N_17353);
and U18629 (N_18629,N_15643,N_15905);
and U18630 (N_18630,N_15426,N_16658);
or U18631 (N_18631,N_15162,N_15234);
xnor U18632 (N_18632,N_15409,N_16859);
nor U18633 (N_18633,N_15890,N_15040);
and U18634 (N_18634,N_17122,N_17426);
or U18635 (N_18635,N_17098,N_17056);
or U18636 (N_18636,N_16262,N_16380);
xor U18637 (N_18637,N_15867,N_15137);
and U18638 (N_18638,N_15899,N_15470);
nor U18639 (N_18639,N_15956,N_16431);
or U18640 (N_18640,N_16979,N_16118);
nor U18641 (N_18641,N_17274,N_15251);
and U18642 (N_18642,N_15246,N_17496);
xnor U18643 (N_18643,N_15193,N_16018);
xnor U18644 (N_18644,N_15113,N_15286);
nor U18645 (N_18645,N_15210,N_15522);
xnor U18646 (N_18646,N_15697,N_17453);
nor U18647 (N_18647,N_16578,N_16341);
nand U18648 (N_18648,N_17136,N_15495);
xor U18649 (N_18649,N_16860,N_15057);
and U18650 (N_18650,N_15676,N_15224);
nand U18651 (N_18651,N_15961,N_16144);
nand U18652 (N_18652,N_15946,N_15245);
and U18653 (N_18653,N_15654,N_16290);
nor U18654 (N_18654,N_16551,N_16372);
or U18655 (N_18655,N_17189,N_16502);
nand U18656 (N_18656,N_16694,N_15901);
xnor U18657 (N_18657,N_15723,N_15514);
nand U18658 (N_18658,N_16282,N_16595);
nand U18659 (N_18659,N_15313,N_15695);
nor U18660 (N_18660,N_15008,N_16562);
or U18661 (N_18661,N_16995,N_16691);
xor U18662 (N_18662,N_16090,N_17062);
nor U18663 (N_18663,N_17074,N_16267);
or U18664 (N_18664,N_15741,N_17064);
nor U18665 (N_18665,N_15662,N_15298);
and U18666 (N_18666,N_15988,N_16255);
and U18667 (N_18667,N_16249,N_16428);
nand U18668 (N_18668,N_16949,N_17371);
or U18669 (N_18669,N_15350,N_15031);
or U18670 (N_18670,N_17379,N_16187);
xor U18671 (N_18671,N_17231,N_16531);
or U18672 (N_18672,N_16774,N_16039);
or U18673 (N_18673,N_15996,N_16712);
or U18674 (N_18674,N_17153,N_15088);
nor U18675 (N_18675,N_15922,N_15385);
nand U18676 (N_18676,N_15280,N_17309);
or U18677 (N_18677,N_16289,N_15986);
or U18678 (N_18678,N_16250,N_16381);
nand U18679 (N_18679,N_15179,N_16003);
or U18680 (N_18680,N_16844,N_15595);
and U18681 (N_18681,N_15264,N_15614);
and U18682 (N_18682,N_15159,N_16940);
nand U18683 (N_18683,N_15292,N_15237);
nor U18684 (N_18684,N_15112,N_16679);
nor U18685 (N_18685,N_15427,N_17024);
and U18686 (N_18686,N_17250,N_15022);
or U18687 (N_18687,N_17147,N_15511);
or U18688 (N_18688,N_16215,N_16637);
xor U18689 (N_18689,N_15062,N_16659);
xor U18690 (N_18690,N_15027,N_16699);
xnor U18691 (N_18691,N_16009,N_16786);
or U18692 (N_18692,N_16097,N_15928);
or U18693 (N_18693,N_17030,N_15214);
xor U18694 (N_18694,N_16705,N_17268);
or U18695 (N_18695,N_15949,N_16386);
and U18696 (N_18696,N_15046,N_15829);
xor U18697 (N_18697,N_16253,N_15284);
or U18698 (N_18698,N_16329,N_15936);
and U18699 (N_18699,N_17265,N_15863);
nor U18700 (N_18700,N_17451,N_16553);
xnor U18701 (N_18701,N_17040,N_15548);
and U18702 (N_18702,N_17222,N_16869);
nor U18703 (N_18703,N_15191,N_15459);
and U18704 (N_18704,N_15558,N_16175);
and U18705 (N_18705,N_15182,N_16730);
xor U18706 (N_18706,N_16793,N_15414);
or U18707 (N_18707,N_15445,N_15603);
and U18708 (N_18708,N_16952,N_15151);
nor U18709 (N_18709,N_16758,N_15894);
nor U18710 (N_18710,N_17151,N_16400);
or U18711 (N_18711,N_17029,N_16592);
nor U18712 (N_18712,N_17154,N_16485);
or U18713 (N_18713,N_15618,N_16095);
or U18714 (N_18714,N_16523,N_15819);
and U18715 (N_18715,N_16468,N_16040);
or U18716 (N_18716,N_16396,N_16365);
and U18717 (N_18717,N_17480,N_16930);
xnor U18718 (N_18718,N_15328,N_16765);
or U18719 (N_18719,N_17191,N_15542);
or U18720 (N_18720,N_16846,N_16935);
and U18721 (N_18721,N_17065,N_16136);
nand U18722 (N_18722,N_16781,N_16602);
nand U18723 (N_18723,N_17304,N_15893);
and U18724 (N_18724,N_17312,N_15510);
and U18725 (N_18725,N_16484,N_15724);
and U18726 (N_18726,N_16159,N_17101);
xnor U18727 (N_18727,N_16244,N_16397);
or U18728 (N_18728,N_15139,N_15702);
and U18729 (N_18729,N_15634,N_15545);
nand U18730 (N_18730,N_15568,N_17336);
and U18731 (N_18731,N_16998,N_16109);
nor U18732 (N_18732,N_17343,N_16205);
and U18733 (N_18733,N_15646,N_17433);
and U18734 (N_18734,N_15521,N_17481);
or U18735 (N_18735,N_16800,N_15367);
and U18736 (N_18736,N_17140,N_16034);
nand U18737 (N_18737,N_15389,N_15029);
nand U18738 (N_18738,N_17471,N_15659);
and U18739 (N_18739,N_16671,N_15217);
and U18740 (N_18740,N_16182,N_15226);
xnor U18741 (N_18741,N_16140,N_16082);
or U18742 (N_18742,N_17427,N_16366);
or U18743 (N_18743,N_17251,N_17220);
xnor U18744 (N_18744,N_16698,N_15156);
nor U18745 (N_18745,N_16653,N_16451);
nor U18746 (N_18746,N_16172,N_16210);
nor U18747 (N_18747,N_15833,N_16185);
or U18748 (N_18748,N_16452,N_16150);
nor U18749 (N_18749,N_16344,N_15876);
and U18750 (N_18750,N_15470,N_16975);
xnor U18751 (N_18751,N_16090,N_16171);
xor U18752 (N_18752,N_16847,N_17362);
or U18753 (N_18753,N_15732,N_16473);
and U18754 (N_18754,N_16998,N_16524);
and U18755 (N_18755,N_16366,N_16586);
xnor U18756 (N_18756,N_15101,N_16876);
xnor U18757 (N_18757,N_16255,N_17499);
and U18758 (N_18758,N_16329,N_15805);
nand U18759 (N_18759,N_17129,N_16498);
nor U18760 (N_18760,N_16741,N_15041);
or U18761 (N_18761,N_16629,N_15508);
xnor U18762 (N_18762,N_17100,N_16077);
or U18763 (N_18763,N_16648,N_15971);
xnor U18764 (N_18764,N_15734,N_17440);
xnor U18765 (N_18765,N_17301,N_17363);
nand U18766 (N_18766,N_17420,N_15626);
xor U18767 (N_18767,N_17124,N_16984);
xor U18768 (N_18768,N_16207,N_16088);
nor U18769 (N_18769,N_15813,N_17026);
nor U18770 (N_18770,N_15474,N_15861);
or U18771 (N_18771,N_15071,N_16792);
nand U18772 (N_18772,N_17005,N_16078);
nor U18773 (N_18773,N_15718,N_17289);
or U18774 (N_18774,N_16322,N_15228);
nor U18775 (N_18775,N_15974,N_15174);
or U18776 (N_18776,N_17245,N_15163);
nor U18777 (N_18777,N_17370,N_16740);
xnor U18778 (N_18778,N_15172,N_15643);
or U18779 (N_18779,N_16975,N_16459);
or U18780 (N_18780,N_16902,N_16384);
or U18781 (N_18781,N_17441,N_15681);
xnor U18782 (N_18782,N_16566,N_16022);
xor U18783 (N_18783,N_15629,N_15758);
nand U18784 (N_18784,N_15133,N_16898);
or U18785 (N_18785,N_15987,N_16260);
and U18786 (N_18786,N_16565,N_17066);
nor U18787 (N_18787,N_17429,N_15817);
nand U18788 (N_18788,N_16584,N_16621);
nor U18789 (N_18789,N_15583,N_16954);
and U18790 (N_18790,N_16334,N_17160);
xor U18791 (N_18791,N_15789,N_15556);
nand U18792 (N_18792,N_15960,N_16648);
and U18793 (N_18793,N_16062,N_16827);
or U18794 (N_18794,N_15908,N_15201);
nor U18795 (N_18795,N_15432,N_17425);
or U18796 (N_18796,N_17419,N_16775);
or U18797 (N_18797,N_15646,N_16192);
xnor U18798 (N_18798,N_16831,N_15274);
xor U18799 (N_18799,N_15689,N_15471);
nand U18800 (N_18800,N_16056,N_16712);
and U18801 (N_18801,N_17053,N_15769);
and U18802 (N_18802,N_15470,N_16958);
and U18803 (N_18803,N_15086,N_15131);
xor U18804 (N_18804,N_15646,N_15082);
xnor U18805 (N_18805,N_16267,N_16025);
nand U18806 (N_18806,N_16336,N_15063);
nand U18807 (N_18807,N_15584,N_16100);
and U18808 (N_18808,N_15461,N_17313);
nand U18809 (N_18809,N_16858,N_16316);
and U18810 (N_18810,N_17209,N_17054);
nor U18811 (N_18811,N_17195,N_16355);
and U18812 (N_18812,N_17105,N_16504);
nand U18813 (N_18813,N_17213,N_16140);
and U18814 (N_18814,N_15962,N_16899);
and U18815 (N_18815,N_16639,N_16962);
nand U18816 (N_18816,N_15885,N_16551);
nor U18817 (N_18817,N_16852,N_16116);
and U18818 (N_18818,N_16351,N_15962);
or U18819 (N_18819,N_16640,N_15992);
xor U18820 (N_18820,N_15423,N_15270);
and U18821 (N_18821,N_15263,N_17082);
or U18822 (N_18822,N_16186,N_17148);
and U18823 (N_18823,N_16566,N_17333);
xnor U18824 (N_18824,N_15649,N_17169);
xor U18825 (N_18825,N_15670,N_16525);
or U18826 (N_18826,N_15573,N_15280);
xnor U18827 (N_18827,N_15522,N_17015);
or U18828 (N_18828,N_15769,N_17469);
or U18829 (N_18829,N_16873,N_17114);
or U18830 (N_18830,N_15263,N_16573);
nor U18831 (N_18831,N_15593,N_15916);
nand U18832 (N_18832,N_17015,N_16286);
and U18833 (N_18833,N_17132,N_15404);
nand U18834 (N_18834,N_16067,N_15283);
or U18835 (N_18835,N_17193,N_16271);
or U18836 (N_18836,N_16480,N_15857);
or U18837 (N_18837,N_16784,N_17456);
xnor U18838 (N_18838,N_17192,N_15426);
xor U18839 (N_18839,N_17017,N_17051);
or U18840 (N_18840,N_15063,N_15946);
or U18841 (N_18841,N_15335,N_15290);
nand U18842 (N_18842,N_15685,N_16522);
xnor U18843 (N_18843,N_16286,N_15730);
or U18844 (N_18844,N_16416,N_15467);
nand U18845 (N_18845,N_16930,N_16963);
xnor U18846 (N_18846,N_16454,N_16722);
xnor U18847 (N_18847,N_15813,N_16740);
nor U18848 (N_18848,N_15994,N_15394);
nand U18849 (N_18849,N_16847,N_15950);
nand U18850 (N_18850,N_17037,N_15215);
or U18851 (N_18851,N_15305,N_16480);
or U18852 (N_18852,N_16351,N_17435);
or U18853 (N_18853,N_16381,N_17047);
xor U18854 (N_18854,N_15024,N_15480);
nand U18855 (N_18855,N_15060,N_15305);
or U18856 (N_18856,N_16140,N_17461);
and U18857 (N_18857,N_17173,N_17434);
nand U18858 (N_18858,N_15285,N_16456);
xor U18859 (N_18859,N_15258,N_15915);
and U18860 (N_18860,N_16762,N_15500);
and U18861 (N_18861,N_16206,N_15606);
and U18862 (N_18862,N_17096,N_15087);
xor U18863 (N_18863,N_16202,N_16382);
nand U18864 (N_18864,N_16625,N_15218);
nor U18865 (N_18865,N_15689,N_15210);
xor U18866 (N_18866,N_16678,N_15299);
xnor U18867 (N_18867,N_16649,N_16385);
nand U18868 (N_18868,N_16032,N_15575);
nand U18869 (N_18869,N_16238,N_15111);
or U18870 (N_18870,N_15451,N_16085);
nand U18871 (N_18871,N_16419,N_17089);
nand U18872 (N_18872,N_15053,N_17320);
nand U18873 (N_18873,N_16930,N_15804);
nor U18874 (N_18874,N_16788,N_16504);
or U18875 (N_18875,N_16254,N_16480);
xor U18876 (N_18876,N_15156,N_16790);
nand U18877 (N_18877,N_15216,N_17033);
xor U18878 (N_18878,N_16989,N_17155);
or U18879 (N_18879,N_16449,N_15045);
xor U18880 (N_18880,N_17341,N_15848);
nor U18881 (N_18881,N_16275,N_17461);
nand U18882 (N_18882,N_15060,N_15030);
xnor U18883 (N_18883,N_16311,N_16518);
nand U18884 (N_18884,N_15539,N_15383);
nor U18885 (N_18885,N_15997,N_16513);
nor U18886 (N_18886,N_15156,N_16262);
and U18887 (N_18887,N_17280,N_15333);
or U18888 (N_18888,N_15009,N_16409);
nand U18889 (N_18889,N_17274,N_15771);
nor U18890 (N_18890,N_17470,N_16821);
or U18891 (N_18891,N_15616,N_16564);
nor U18892 (N_18892,N_16940,N_16018);
and U18893 (N_18893,N_16315,N_15698);
nor U18894 (N_18894,N_15246,N_16824);
or U18895 (N_18895,N_17204,N_16396);
nor U18896 (N_18896,N_16044,N_16517);
and U18897 (N_18897,N_15769,N_17472);
xor U18898 (N_18898,N_16609,N_16427);
and U18899 (N_18899,N_16930,N_17149);
and U18900 (N_18900,N_15648,N_15370);
xor U18901 (N_18901,N_16582,N_16964);
and U18902 (N_18902,N_16847,N_17231);
nand U18903 (N_18903,N_15805,N_16481);
nand U18904 (N_18904,N_16424,N_15255);
xnor U18905 (N_18905,N_15439,N_16383);
and U18906 (N_18906,N_16332,N_16040);
nor U18907 (N_18907,N_15053,N_15919);
xnor U18908 (N_18908,N_15948,N_17007);
xnor U18909 (N_18909,N_15131,N_16662);
nand U18910 (N_18910,N_16678,N_16299);
or U18911 (N_18911,N_17294,N_16693);
and U18912 (N_18912,N_15627,N_15737);
nand U18913 (N_18913,N_15178,N_15751);
and U18914 (N_18914,N_16836,N_17114);
xnor U18915 (N_18915,N_16733,N_15381);
or U18916 (N_18916,N_17356,N_16482);
or U18917 (N_18917,N_15074,N_17162);
and U18918 (N_18918,N_17258,N_16413);
xnor U18919 (N_18919,N_15930,N_17098);
nand U18920 (N_18920,N_16996,N_15934);
and U18921 (N_18921,N_16785,N_16398);
xnor U18922 (N_18922,N_17127,N_15016);
nor U18923 (N_18923,N_15915,N_15160);
or U18924 (N_18924,N_16240,N_17334);
nor U18925 (N_18925,N_16147,N_15090);
xnor U18926 (N_18926,N_15827,N_17282);
nor U18927 (N_18927,N_16622,N_16400);
and U18928 (N_18928,N_15812,N_15498);
and U18929 (N_18929,N_15153,N_15505);
nand U18930 (N_18930,N_17163,N_16565);
or U18931 (N_18931,N_17454,N_17165);
xor U18932 (N_18932,N_17187,N_17002);
nand U18933 (N_18933,N_15400,N_15015);
nand U18934 (N_18934,N_15208,N_15444);
nor U18935 (N_18935,N_16808,N_16836);
nor U18936 (N_18936,N_16680,N_15364);
xnor U18937 (N_18937,N_17139,N_15438);
and U18938 (N_18938,N_17136,N_15487);
nor U18939 (N_18939,N_17404,N_16007);
or U18940 (N_18940,N_16233,N_15540);
nor U18941 (N_18941,N_15276,N_15105);
and U18942 (N_18942,N_16442,N_16167);
xor U18943 (N_18943,N_17211,N_16446);
nor U18944 (N_18944,N_15349,N_16692);
and U18945 (N_18945,N_16114,N_15569);
xnor U18946 (N_18946,N_15668,N_17161);
xor U18947 (N_18947,N_16759,N_15775);
xor U18948 (N_18948,N_15865,N_16435);
and U18949 (N_18949,N_16021,N_16885);
nor U18950 (N_18950,N_15226,N_15371);
nor U18951 (N_18951,N_15953,N_16447);
nor U18952 (N_18952,N_17287,N_15384);
nor U18953 (N_18953,N_15225,N_16020);
nand U18954 (N_18954,N_16807,N_17056);
nand U18955 (N_18955,N_15028,N_15549);
and U18956 (N_18956,N_17069,N_17106);
or U18957 (N_18957,N_15492,N_15030);
and U18958 (N_18958,N_15958,N_17216);
nor U18959 (N_18959,N_16566,N_15082);
or U18960 (N_18960,N_17224,N_15491);
nor U18961 (N_18961,N_16151,N_16046);
or U18962 (N_18962,N_15426,N_15244);
nand U18963 (N_18963,N_15793,N_16010);
and U18964 (N_18964,N_15076,N_16661);
nand U18965 (N_18965,N_16346,N_17364);
nand U18966 (N_18966,N_16901,N_16895);
xnor U18967 (N_18967,N_15958,N_16366);
xor U18968 (N_18968,N_15171,N_17444);
xnor U18969 (N_18969,N_17254,N_16446);
and U18970 (N_18970,N_15126,N_16934);
xnor U18971 (N_18971,N_15555,N_15439);
or U18972 (N_18972,N_16269,N_17448);
or U18973 (N_18973,N_17076,N_17297);
xnor U18974 (N_18974,N_15494,N_15551);
xor U18975 (N_18975,N_16198,N_16225);
nand U18976 (N_18976,N_16508,N_17264);
or U18977 (N_18977,N_16311,N_17085);
nor U18978 (N_18978,N_15398,N_16222);
nor U18979 (N_18979,N_15728,N_16296);
nand U18980 (N_18980,N_15680,N_17129);
xnor U18981 (N_18981,N_17258,N_15486);
xnor U18982 (N_18982,N_15257,N_15208);
and U18983 (N_18983,N_17487,N_17177);
xor U18984 (N_18984,N_16571,N_16409);
or U18985 (N_18985,N_17125,N_15469);
nand U18986 (N_18986,N_15922,N_15488);
xnor U18987 (N_18987,N_16687,N_16317);
nor U18988 (N_18988,N_15777,N_15451);
and U18989 (N_18989,N_15486,N_16273);
and U18990 (N_18990,N_16933,N_16280);
or U18991 (N_18991,N_15152,N_17086);
nand U18992 (N_18992,N_16513,N_17152);
or U18993 (N_18993,N_16615,N_16977);
nor U18994 (N_18994,N_15436,N_15521);
and U18995 (N_18995,N_17437,N_17352);
or U18996 (N_18996,N_15171,N_17463);
or U18997 (N_18997,N_15378,N_16477);
nand U18998 (N_18998,N_16418,N_17169);
nand U18999 (N_18999,N_15396,N_16772);
nand U19000 (N_19000,N_15713,N_16684);
nor U19001 (N_19001,N_16483,N_16968);
xnor U19002 (N_19002,N_17075,N_15584);
nand U19003 (N_19003,N_15199,N_16700);
or U19004 (N_19004,N_17427,N_16225);
and U19005 (N_19005,N_15689,N_15295);
xnor U19006 (N_19006,N_15384,N_16122);
or U19007 (N_19007,N_15566,N_15380);
nand U19008 (N_19008,N_15420,N_16038);
or U19009 (N_19009,N_16998,N_16525);
and U19010 (N_19010,N_15404,N_15016);
nor U19011 (N_19011,N_16384,N_15123);
and U19012 (N_19012,N_17478,N_15999);
nor U19013 (N_19013,N_15133,N_15263);
or U19014 (N_19014,N_15201,N_15340);
and U19015 (N_19015,N_16982,N_16131);
and U19016 (N_19016,N_16056,N_17188);
and U19017 (N_19017,N_16178,N_17116);
nor U19018 (N_19018,N_16449,N_16347);
or U19019 (N_19019,N_16645,N_16046);
or U19020 (N_19020,N_16021,N_17322);
and U19021 (N_19021,N_17160,N_15139);
nand U19022 (N_19022,N_15630,N_15184);
or U19023 (N_19023,N_16832,N_16955);
xnor U19024 (N_19024,N_16105,N_17187);
and U19025 (N_19025,N_16630,N_15594);
and U19026 (N_19026,N_16647,N_16343);
xnor U19027 (N_19027,N_17455,N_16744);
nor U19028 (N_19028,N_15419,N_17246);
nor U19029 (N_19029,N_17035,N_15219);
nor U19030 (N_19030,N_17467,N_15199);
nand U19031 (N_19031,N_16343,N_17080);
nand U19032 (N_19032,N_16205,N_15424);
xnor U19033 (N_19033,N_16781,N_15780);
xor U19034 (N_19034,N_17350,N_15020);
and U19035 (N_19035,N_15773,N_16232);
xnor U19036 (N_19036,N_16287,N_15128);
or U19037 (N_19037,N_15724,N_16376);
xor U19038 (N_19038,N_16267,N_16138);
nor U19039 (N_19039,N_16890,N_16253);
and U19040 (N_19040,N_16308,N_16010);
nand U19041 (N_19041,N_15770,N_16144);
and U19042 (N_19042,N_17194,N_16854);
or U19043 (N_19043,N_16866,N_16194);
or U19044 (N_19044,N_17297,N_16056);
or U19045 (N_19045,N_16959,N_15069);
nor U19046 (N_19046,N_16635,N_15930);
and U19047 (N_19047,N_16935,N_15499);
or U19048 (N_19048,N_16048,N_16755);
and U19049 (N_19049,N_17189,N_17401);
nor U19050 (N_19050,N_16868,N_16923);
xor U19051 (N_19051,N_15811,N_15787);
and U19052 (N_19052,N_17237,N_17166);
nor U19053 (N_19053,N_15389,N_15576);
nand U19054 (N_19054,N_16024,N_15930);
nor U19055 (N_19055,N_16723,N_17405);
and U19056 (N_19056,N_15920,N_16092);
and U19057 (N_19057,N_17065,N_16564);
or U19058 (N_19058,N_15980,N_15331);
xor U19059 (N_19059,N_16718,N_15425);
nand U19060 (N_19060,N_15332,N_17118);
or U19061 (N_19061,N_15501,N_15405);
and U19062 (N_19062,N_16330,N_15449);
xnor U19063 (N_19063,N_16391,N_16685);
and U19064 (N_19064,N_15317,N_16066);
xnor U19065 (N_19065,N_16775,N_17451);
or U19066 (N_19066,N_15496,N_15960);
nand U19067 (N_19067,N_17153,N_16386);
nand U19068 (N_19068,N_16581,N_16242);
or U19069 (N_19069,N_15442,N_16835);
nor U19070 (N_19070,N_16794,N_15073);
nand U19071 (N_19071,N_16162,N_15879);
and U19072 (N_19072,N_16285,N_17023);
and U19073 (N_19073,N_15170,N_16036);
nand U19074 (N_19074,N_16343,N_16773);
nand U19075 (N_19075,N_17383,N_17364);
nand U19076 (N_19076,N_17283,N_17300);
nand U19077 (N_19077,N_16185,N_15295);
nor U19078 (N_19078,N_16379,N_17485);
nor U19079 (N_19079,N_16880,N_17123);
nor U19080 (N_19080,N_17308,N_15497);
xor U19081 (N_19081,N_17172,N_15671);
nor U19082 (N_19082,N_15019,N_15000);
nand U19083 (N_19083,N_17275,N_16262);
nor U19084 (N_19084,N_15950,N_16531);
nand U19085 (N_19085,N_15643,N_15497);
nor U19086 (N_19086,N_15163,N_15890);
xor U19087 (N_19087,N_15208,N_16953);
nand U19088 (N_19088,N_15475,N_15367);
xor U19089 (N_19089,N_15809,N_15040);
and U19090 (N_19090,N_16576,N_15131);
and U19091 (N_19091,N_16390,N_16208);
nand U19092 (N_19092,N_16255,N_17404);
nor U19093 (N_19093,N_15700,N_15432);
nor U19094 (N_19094,N_15641,N_17026);
nor U19095 (N_19095,N_17165,N_15755);
nand U19096 (N_19096,N_16342,N_16828);
or U19097 (N_19097,N_15068,N_17186);
nor U19098 (N_19098,N_15339,N_16225);
nor U19099 (N_19099,N_15776,N_16435);
nor U19100 (N_19100,N_17349,N_17442);
xor U19101 (N_19101,N_15655,N_15547);
and U19102 (N_19102,N_15189,N_16998);
xor U19103 (N_19103,N_15316,N_15842);
nor U19104 (N_19104,N_16983,N_17471);
or U19105 (N_19105,N_16810,N_16712);
or U19106 (N_19106,N_16590,N_17183);
or U19107 (N_19107,N_17061,N_16310);
nand U19108 (N_19108,N_17395,N_15235);
xnor U19109 (N_19109,N_15645,N_17164);
nor U19110 (N_19110,N_16568,N_16101);
nor U19111 (N_19111,N_16160,N_15668);
or U19112 (N_19112,N_17020,N_17086);
nand U19113 (N_19113,N_16246,N_16998);
nand U19114 (N_19114,N_16389,N_16940);
nand U19115 (N_19115,N_15070,N_17379);
or U19116 (N_19116,N_15029,N_15327);
nand U19117 (N_19117,N_16458,N_17108);
xnor U19118 (N_19118,N_17421,N_16304);
nor U19119 (N_19119,N_16205,N_15492);
or U19120 (N_19120,N_16447,N_15820);
xnor U19121 (N_19121,N_15493,N_15000);
nor U19122 (N_19122,N_15272,N_17421);
xnor U19123 (N_19123,N_17443,N_15121);
nand U19124 (N_19124,N_16620,N_15240);
nand U19125 (N_19125,N_16620,N_15000);
or U19126 (N_19126,N_16837,N_17494);
or U19127 (N_19127,N_16874,N_16347);
xor U19128 (N_19128,N_16763,N_15617);
or U19129 (N_19129,N_15707,N_15613);
or U19130 (N_19130,N_16356,N_17004);
xor U19131 (N_19131,N_15745,N_15367);
nand U19132 (N_19132,N_15402,N_16216);
and U19133 (N_19133,N_16818,N_16784);
nand U19134 (N_19134,N_16189,N_15073);
and U19135 (N_19135,N_16479,N_16524);
or U19136 (N_19136,N_15094,N_16538);
xor U19137 (N_19137,N_15668,N_16413);
nand U19138 (N_19138,N_16979,N_17114);
nor U19139 (N_19139,N_17447,N_16767);
nand U19140 (N_19140,N_16396,N_17154);
nand U19141 (N_19141,N_15944,N_15614);
and U19142 (N_19142,N_15046,N_16715);
nor U19143 (N_19143,N_17499,N_16781);
nand U19144 (N_19144,N_15250,N_16049);
and U19145 (N_19145,N_15622,N_16735);
nor U19146 (N_19146,N_16179,N_15742);
and U19147 (N_19147,N_15991,N_15861);
nor U19148 (N_19148,N_15564,N_17266);
nand U19149 (N_19149,N_17062,N_17389);
or U19150 (N_19150,N_16137,N_16742);
xor U19151 (N_19151,N_16079,N_16483);
or U19152 (N_19152,N_16855,N_16517);
xnor U19153 (N_19153,N_15752,N_17015);
xnor U19154 (N_19154,N_17345,N_16737);
and U19155 (N_19155,N_16857,N_16215);
xnor U19156 (N_19156,N_17494,N_16993);
nand U19157 (N_19157,N_16783,N_16506);
or U19158 (N_19158,N_15995,N_16694);
and U19159 (N_19159,N_16916,N_17252);
nor U19160 (N_19160,N_15605,N_17397);
nand U19161 (N_19161,N_16499,N_15911);
xnor U19162 (N_19162,N_15086,N_15904);
nand U19163 (N_19163,N_17412,N_16132);
or U19164 (N_19164,N_15054,N_15810);
and U19165 (N_19165,N_16741,N_15397);
nand U19166 (N_19166,N_16102,N_15594);
and U19167 (N_19167,N_16788,N_16931);
nand U19168 (N_19168,N_16164,N_15419);
nor U19169 (N_19169,N_16630,N_16515);
nand U19170 (N_19170,N_15183,N_17197);
xnor U19171 (N_19171,N_15764,N_16309);
nand U19172 (N_19172,N_16537,N_17449);
and U19173 (N_19173,N_16754,N_15288);
nor U19174 (N_19174,N_15496,N_16177);
or U19175 (N_19175,N_16755,N_17405);
nor U19176 (N_19176,N_15567,N_16938);
nand U19177 (N_19177,N_16695,N_16419);
and U19178 (N_19178,N_17488,N_16958);
and U19179 (N_19179,N_16392,N_16153);
nand U19180 (N_19180,N_16839,N_15591);
or U19181 (N_19181,N_15298,N_15967);
and U19182 (N_19182,N_17467,N_17051);
nor U19183 (N_19183,N_16404,N_15835);
nand U19184 (N_19184,N_15520,N_17149);
xor U19185 (N_19185,N_17363,N_15813);
and U19186 (N_19186,N_15349,N_15047);
or U19187 (N_19187,N_15341,N_16460);
or U19188 (N_19188,N_17297,N_16387);
or U19189 (N_19189,N_16472,N_17470);
nand U19190 (N_19190,N_16375,N_16192);
xor U19191 (N_19191,N_15728,N_16250);
nand U19192 (N_19192,N_16513,N_16559);
or U19193 (N_19193,N_16162,N_17427);
xnor U19194 (N_19194,N_15636,N_16001);
nand U19195 (N_19195,N_15025,N_17205);
or U19196 (N_19196,N_15290,N_17057);
nand U19197 (N_19197,N_16376,N_15249);
nor U19198 (N_19198,N_15420,N_16745);
and U19199 (N_19199,N_15286,N_17492);
xor U19200 (N_19200,N_15290,N_16142);
or U19201 (N_19201,N_15106,N_16425);
xor U19202 (N_19202,N_16188,N_16294);
xor U19203 (N_19203,N_16085,N_15062);
or U19204 (N_19204,N_15986,N_17077);
or U19205 (N_19205,N_16362,N_15655);
or U19206 (N_19206,N_16594,N_16070);
nand U19207 (N_19207,N_15335,N_15514);
xnor U19208 (N_19208,N_15632,N_17263);
and U19209 (N_19209,N_15286,N_15911);
nor U19210 (N_19210,N_15397,N_17357);
nand U19211 (N_19211,N_17060,N_15557);
xnor U19212 (N_19212,N_15382,N_15179);
xnor U19213 (N_19213,N_16673,N_17428);
xnor U19214 (N_19214,N_16185,N_16514);
and U19215 (N_19215,N_16591,N_16032);
or U19216 (N_19216,N_16491,N_16566);
or U19217 (N_19217,N_16627,N_15655);
xnor U19218 (N_19218,N_15813,N_16373);
and U19219 (N_19219,N_15293,N_15942);
xnor U19220 (N_19220,N_16979,N_15853);
and U19221 (N_19221,N_15827,N_17305);
nor U19222 (N_19222,N_15028,N_16741);
nand U19223 (N_19223,N_15884,N_16885);
and U19224 (N_19224,N_15694,N_15043);
nor U19225 (N_19225,N_16335,N_15412);
nor U19226 (N_19226,N_16553,N_16511);
or U19227 (N_19227,N_15399,N_17208);
and U19228 (N_19228,N_15643,N_15802);
nor U19229 (N_19229,N_17058,N_16772);
and U19230 (N_19230,N_16795,N_15439);
or U19231 (N_19231,N_16389,N_16002);
xor U19232 (N_19232,N_15108,N_15969);
nand U19233 (N_19233,N_16580,N_17044);
nor U19234 (N_19234,N_15998,N_16237);
nand U19235 (N_19235,N_16708,N_16067);
nand U19236 (N_19236,N_15391,N_16571);
and U19237 (N_19237,N_15470,N_16064);
nand U19238 (N_19238,N_15824,N_16339);
xnor U19239 (N_19239,N_16121,N_15390);
and U19240 (N_19240,N_17121,N_16279);
and U19241 (N_19241,N_17230,N_16942);
and U19242 (N_19242,N_16235,N_17136);
xnor U19243 (N_19243,N_15948,N_15865);
and U19244 (N_19244,N_15599,N_16525);
and U19245 (N_19245,N_16599,N_15033);
nand U19246 (N_19246,N_16563,N_16324);
or U19247 (N_19247,N_16710,N_16564);
nor U19248 (N_19248,N_16788,N_16519);
and U19249 (N_19249,N_16647,N_15500);
or U19250 (N_19250,N_15855,N_15907);
or U19251 (N_19251,N_16246,N_15482);
nand U19252 (N_19252,N_15050,N_16404);
nor U19253 (N_19253,N_16665,N_16692);
xor U19254 (N_19254,N_15721,N_16301);
nor U19255 (N_19255,N_16949,N_17470);
or U19256 (N_19256,N_15746,N_16843);
nand U19257 (N_19257,N_16756,N_16646);
nand U19258 (N_19258,N_16922,N_17061);
xnor U19259 (N_19259,N_16231,N_15605);
or U19260 (N_19260,N_15435,N_16033);
or U19261 (N_19261,N_16468,N_16682);
and U19262 (N_19262,N_17191,N_15644);
nand U19263 (N_19263,N_17218,N_16734);
xnor U19264 (N_19264,N_17335,N_15911);
xor U19265 (N_19265,N_15944,N_16957);
and U19266 (N_19266,N_16982,N_17055);
nor U19267 (N_19267,N_15388,N_15777);
xnor U19268 (N_19268,N_15591,N_16995);
xnor U19269 (N_19269,N_17088,N_16331);
or U19270 (N_19270,N_15964,N_15946);
nor U19271 (N_19271,N_15184,N_16319);
xnor U19272 (N_19272,N_17225,N_15407);
and U19273 (N_19273,N_15885,N_17485);
nor U19274 (N_19274,N_17458,N_17459);
xnor U19275 (N_19275,N_15703,N_15101);
nand U19276 (N_19276,N_16961,N_16192);
and U19277 (N_19277,N_17218,N_15641);
nor U19278 (N_19278,N_17282,N_17400);
xor U19279 (N_19279,N_17381,N_15773);
xnor U19280 (N_19280,N_17365,N_17274);
or U19281 (N_19281,N_16121,N_17003);
or U19282 (N_19282,N_17321,N_16753);
nor U19283 (N_19283,N_16898,N_15540);
xnor U19284 (N_19284,N_16714,N_16269);
xnor U19285 (N_19285,N_16700,N_16213);
or U19286 (N_19286,N_15946,N_15100);
nor U19287 (N_19287,N_16205,N_15709);
and U19288 (N_19288,N_16982,N_17374);
nor U19289 (N_19289,N_16103,N_16268);
or U19290 (N_19290,N_15437,N_15572);
nand U19291 (N_19291,N_16059,N_15623);
nor U19292 (N_19292,N_17111,N_17004);
nand U19293 (N_19293,N_16414,N_16574);
xor U19294 (N_19294,N_16251,N_15602);
nand U19295 (N_19295,N_16175,N_16743);
and U19296 (N_19296,N_15947,N_15698);
nor U19297 (N_19297,N_15460,N_17081);
and U19298 (N_19298,N_16407,N_15085);
nor U19299 (N_19299,N_17156,N_15303);
and U19300 (N_19300,N_15790,N_16333);
and U19301 (N_19301,N_16247,N_15707);
or U19302 (N_19302,N_15980,N_16281);
and U19303 (N_19303,N_15621,N_15268);
nand U19304 (N_19304,N_15061,N_16444);
xor U19305 (N_19305,N_15457,N_15109);
xor U19306 (N_19306,N_15798,N_16733);
nand U19307 (N_19307,N_16895,N_17030);
or U19308 (N_19308,N_16938,N_15209);
nor U19309 (N_19309,N_15734,N_16798);
xnor U19310 (N_19310,N_16706,N_15964);
or U19311 (N_19311,N_16707,N_16416);
nand U19312 (N_19312,N_15470,N_15625);
xor U19313 (N_19313,N_17313,N_15579);
nand U19314 (N_19314,N_17388,N_15968);
nor U19315 (N_19315,N_15810,N_16846);
and U19316 (N_19316,N_16635,N_17423);
nor U19317 (N_19317,N_15418,N_16455);
or U19318 (N_19318,N_16394,N_17251);
and U19319 (N_19319,N_16841,N_16913);
nand U19320 (N_19320,N_16407,N_16412);
xnor U19321 (N_19321,N_15395,N_15689);
and U19322 (N_19322,N_15595,N_15017);
nor U19323 (N_19323,N_16253,N_16057);
xnor U19324 (N_19324,N_16189,N_17112);
or U19325 (N_19325,N_15852,N_16992);
nor U19326 (N_19326,N_15799,N_16980);
nand U19327 (N_19327,N_17448,N_16518);
and U19328 (N_19328,N_15757,N_17114);
and U19329 (N_19329,N_15085,N_15434);
nor U19330 (N_19330,N_16016,N_17464);
xor U19331 (N_19331,N_17122,N_17039);
xnor U19332 (N_19332,N_16523,N_16179);
nand U19333 (N_19333,N_16963,N_16532);
xnor U19334 (N_19334,N_15343,N_16565);
or U19335 (N_19335,N_15250,N_17337);
and U19336 (N_19336,N_15098,N_15314);
xor U19337 (N_19337,N_15888,N_15904);
nand U19338 (N_19338,N_15943,N_17391);
xnor U19339 (N_19339,N_17008,N_16507);
and U19340 (N_19340,N_15453,N_15050);
nand U19341 (N_19341,N_16167,N_16194);
xor U19342 (N_19342,N_17454,N_16733);
nor U19343 (N_19343,N_15087,N_15832);
xnor U19344 (N_19344,N_16376,N_17427);
nand U19345 (N_19345,N_15568,N_15089);
nor U19346 (N_19346,N_16601,N_16896);
and U19347 (N_19347,N_15686,N_17389);
xor U19348 (N_19348,N_17466,N_15562);
or U19349 (N_19349,N_15863,N_15223);
nand U19350 (N_19350,N_15512,N_16077);
nor U19351 (N_19351,N_15303,N_16237);
nand U19352 (N_19352,N_15578,N_17348);
nand U19353 (N_19353,N_15988,N_16143);
or U19354 (N_19354,N_16982,N_15208);
xor U19355 (N_19355,N_17234,N_17434);
nand U19356 (N_19356,N_15034,N_17051);
nor U19357 (N_19357,N_17041,N_15683);
and U19358 (N_19358,N_15852,N_15849);
or U19359 (N_19359,N_15727,N_16041);
or U19360 (N_19360,N_15762,N_17080);
nor U19361 (N_19361,N_15669,N_15753);
nor U19362 (N_19362,N_17159,N_15796);
or U19363 (N_19363,N_15520,N_17496);
xnor U19364 (N_19364,N_15057,N_17364);
xor U19365 (N_19365,N_15403,N_16402);
nand U19366 (N_19366,N_15565,N_15906);
xor U19367 (N_19367,N_16645,N_17065);
xor U19368 (N_19368,N_17195,N_17146);
and U19369 (N_19369,N_17299,N_15422);
nor U19370 (N_19370,N_15488,N_15437);
nand U19371 (N_19371,N_16563,N_17260);
xnor U19372 (N_19372,N_15008,N_15260);
and U19373 (N_19373,N_16036,N_17420);
or U19374 (N_19374,N_16991,N_16274);
and U19375 (N_19375,N_15975,N_15897);
or U19376 (N_19376,N_15478,N_16660);
nand U19377 (N_19377,N_15006,N_16821);
xnor U19378 (N_19378,N_16233,N_15234);
nor U19379 (N_19379,N_15849,N_17457);
nand U19380 (N_19380,N_15351,N_16550);
nand U19381 (N_19381,N_17007,N_15983);
and U19382 (N_19382,N_16506,N_17042);
and U19383 (N_19383,N_16402,N_16645);
or U19384 (N_19384,N_17013,N_17193);
xor U19385 (N_19385,N_16482,N_17276);
nor U19386 (N_19386,N_16613,N_15422);
nand U19387 (N_19387,N_15758,N_15391);
and U19388 (N_19388,N_17381,N_16056);
and U19389 (N_19389,N_16029,N_16470);
or U19390 (N_19390,N_17425,N_16923);
and U19391 (N_19391,N_15790,N_16737);
and U19392 (N_19392,N_16640,N_17401);
or U19393 (N_19393,N_16659,N_15209);
or U19394 (N_19394,N_17403,N_17065);
nand U19395 (N_19395,N_17121,N_16904);
nor U19396 (N_19396,N_16561,N_16542);
nor U19397 (N_19397,N_16928,N_15386);
and U19398 (N_19398,N_15465,N_15396);
nand U19399 (N_19399,N_17381,N_16242);
or U19400 (N_19400,N_15175,N_17432);
nor U19401 (N_19401,N_15275,N_15298);
or U19402 (N_19402,N_16959,N_16845);
and U19403 (N_19403,N_15733,N_16267);
and U19404 (N_19404,N_16303,N_16757);
nand U19405 (N_19405,N_16771,N_17062);
nand U19406 (N_19406,N_16027,N_16443);
nor U19407 (N_19407,N_16944,N_16906);
or U19408 (N_19408,N_15732,N_17173);
and U19409 (N_19409,N_17197,N_16362);
or U19410 (N_19410,N_16117,N_16453);
and U19411 (N_19411,N_15546,N_15091);
and U19412 (N_19412,N_16895,N_15862);
xnor U19413 (N_19413,N_15441,N_15876);
nor U19414 (N_19414,N_15658,N_15598);
xor U19415 (N_19415,N_15068,N_17401);
xor U19416 (N_19416,N_15799,N_16220);
and U19417 (N_19417,N_16795,N_15063);
xnor U19418 (N_19418,N_17169,N_15983);
nand U19419 (N_19419,N_15765,N_15221);
nor U19420 (N_19420,N_16038,N_17356);
nor U19421 (N_19421,N_15521,N_16061);
and U19422 (N_19422,N_17085,N_16171);
nand U19423 (N_19423,N_17111,N_15592);
xnor U19424 (N_19424,N_15551,N_17415);
nor U19425 (N_19425,N_15012,N_16443);
or U19426 (N_19426,N_15096,N_15705);
xnor U19427 (N_19427,N_17131,N_16049);
xnor U19428 (N_19428,N_15264,N_16247);
or U19429 (N_19429,N_16763,N_16923);
or U19430 (N_19430,N_17432,N_15984);
xnor U19431 (N_19431,N_17333,N_15375);
or U19432 (N_19432,N_16502,N_15917);
and U19433 (N_19433,N_16366,N_15798);
and U19434 (N_19434,N_16201,N_16049);
or U19435 (N_19435,N_16558,N_17484);
and U19436 (N_19436,N_15054,N_15380);
nand U19437 (N_19437,N_15757,N_16310);
xor U19438 (N_19438,N_16068,N_15848);
or U19439 (N_19439,N_15960,N_15189);
nor U19440 (N_19440,N_15116,N_16746);
nand U19441 (N_19441,N_15722,N_16723);
nand U19442 (N_19442,N_17317,N_16116);
xor U19443 (N_19443,N_15949,N_17175);
and U19444 (N_19444,N_17038,N_17498);
and U19445 (N_19445,N_15992,N_16455);
xnor U19446 (N_19446,N_16810,N_15612);
xor U19447 (N_19447,N_17146,N_16741);
nor U19448 (N_19448,N_17206,N_16950);
nor U19449 (N_19449,N_15942,N_15856);
nor U19450 (N_19450,N_16339,N_15045);
nand U19451 (N_19451,N_17488,N_16951);
and U19452 (N_19452,N_15803,N_17187);
or U19453 (N_19453,N_17103,N_17447);
or U19454 (N_19454,N_16363,N_16970);
xnor U19455 (N_19455,N_16757,N_16693);
nor U19456 (N_19456,N_17057,N_16747);
or U19457 (N_19457,N_17314,N_15463);
and U19458 (N_19458,N_15657,N_16832);
xor U19459 (N_19459,N_15429,N_15282);
or U19460 (N_19460,N_15901,N_16082);
xor U19461 (N_19461,N_15927,N_16858);
or U19462 (N_19462,N_15726,N_15874);
xor U19463 (N_19463,N_15595,N_17366);
xnor U19464 (N_19464,N_17447,N_16136);
and U19465 (N_19465,N_17076,N_17080);
and U19466 (N_19466,N_15407,N_15025);
nand U19467 (N_19467,N_15035,N_15542);
nor U19468 (N_19468,N_16351,N_16928);
xnor U19469 (N_19469,N_16554,N_16679);
nand U19470 (N_19470,N_16133,N_16527);
nand U19471 (N_19471,N_16780,N_17103);
nand U19472 (N_19472,N_15363,N_17389);
or U19473 (N_19473,N_15597,N_16384);
nor U19474 (N_19474,N_17080,N_15487);
and U19475 (N_19475,N_16542,N_16491);
nor U19476 (N_19476,N_15729,N_15408);
or U19477 (N_19477,N_16718,N_17442);
xor U19478 (N_19478,N_16031,N_15471);
nand U19479 (N_19479,N_17402,N_17023);
and U19480 (N_19480,N_16708,N_16732);
nand U19481 (N_19481,N_15939,N_15662);
nand U19482 (N_19482,N_15339,N_15565);
nand U19483 (N_19483,N_16521,N_15408);
nand U19484 (N_19484,N_16134,N_16963);
or U19485 (N_19485,N_16354,N_15548);
xnor U19486 (N_19486,N_16919,N_17229);
or U19487 (N_19487,N_16597,N_16888);
or U19488 (N_19488,N_16934,N_15812);
or U19489 (N_19489,N_15474,N_16833);
nor U19490 (N_19490,N_15072,N_17145);
or U19491 (N_19491,N_17442,N_15775);
or U19492 (N_19492,N_16840,N_15664);
or U19493 (N_19493,N_16031,N_15225);
xor U19494 (N_19494,N_16010,N_15977);
nor U19495 (N_19495,N_16134,N_16575);
xor U19496 (N_19496,N_15631,N_15681);
and U19497 (N_19497,N_15571,N_15449);
nor U19498 (N_19498,N_17115,N_15061);
nor U19499 (N_19499,N_16334,N_16465);
nor U19500 (N_19500,N_17260,N_16091);
and U19501 (N_19501,N_16577,N_15456);
nor U19502 (N_19502,N_17478,N_15752);
nor U19503 (N_19503,N_15237,N_15437);
or U19504 (N_19504,N_16214,N_15353);
or U19505 (N_19505,N_16760,N_15342);
and U19506 (N_19506,N_17216,N_15308);
and U19507 (N_19507,N_17208,N_15123);
xor U19508 (N_19508,N_16155,N_16274);
or U19509 (N_19509,N_15422,N_15976);
nand U19510 (N_19510,N_16823,N_17159);
xnor U19511 (N_19511,N_15077,N_17042);
nor U19512 (N_19512,N_16276,N_15475);
or U19513 (N_19513,N_15657,N_16881);
nand U19514 (N_19514,N_16078,N_16436);
nor U19515 (N_19515,N_16752,N_16446);
nor U19516 (N_19516,N_17431,N_16226);
or U19517 (N_19517,N_16985,N_16376);
and U19518 (N_19518,N_15377,N_15225);
xnor U19519 (N_19519,N_15492,N_16144);
and U19520 (N_19520,N_16292,N_15077);
and U19521 (N_19521,N_17269,N_17053);
nor U19522 (N_19522,N_17139,N_15149);
nand U19523 (N_19523,N_15021,N_17329);
nand U19524 (N_19524,N_16283,N_15050);
or U19525 (N_19525,N_15478,N_17257);
nand U19526 (N_19526,N_16246,N_17195);
or U19527 (N_19527,N_17168,N_16479);
xor U19528 (N_19528,N_16505,N_16442);
nand U19529 (N_19529,N_15756,N_15496);
and U19530 (N_19530,N_17223,N_15128);
or U19531 (N_19531,N_16751,N_16044);
xor U19532 (N_19532,N_16482,N_16223);
nand U19533 (N_19533,N_16373,N_15595);
xor U19534 (N_19534,N_17490,N_15615);
or U19535 (N_19535,N_15613,N_17047);
nor U19536 (N_19536,N_16474,N_16309);
nor U19537 (N_19537,N_15044,N_15133);
xor U19538 (N_19538,N_16471,N_16041);
nor U19539 (N_19539,N_15710,N_16478);
nor U19540 (N_19540,N_15899,N_15157);
or U19541 (N_19541,N_16791,N_15523);
nand U19542 (N_19542,N_15782,N_15578);
and U19543 (N_19543,N_16040,N_15192);
nor U19544 (N_19544,N_15350,N_17116);
nand U19545 (N_19545,N_15789,N_15805);
xnor U19546 (N_19546,N_16649,N_15756);
xor U19547 (N_19547,N_17058,N_17429);
xnor U19548 (N_19548,N_15905,N_15043);
and U19549 (N_19549,N_15799,N_17467);
and U19550 (N_19550,N_16736,N_16902);
or U19551 (N_19551,N_15729,N_16737);
and U19552 (N_19552,N_15440,N_15380);
nor U19553 (N_19553,N_16636,N_17193);
nor U19554 (N_19554,N_15222,N_15125);
or U19555 (N_19555,N_15177,N_16923);
xor U19556 (N_19556,N_15442,N_15672);
nand U19557 (N_19557,N_15511,N_16533);
or U19558 (N_19558,N_15350,N_15897);
xor U19559 (N_19559,N_16500,N_15117);
and U19560 (N_19560,N_16313,N_15747);
or U19561 (N_19561,N_15630,N_15913);
nor U19562 (N_19562,N_17215,N_16378);
or U19563 (N_19563,N_16511,N_15981);
xor U19564 (N_19564,N_17172,N_16282);
and U19565 (N_19565,N_15561,N_16839);
nor U19566 (N_19566,N_16016,N_16622);
xnor U19567 (N_19567,N_16037,N_15500);
or U19568 (N_19568,N_16998,N_16564);
or U19569 (N_19569,N_17030,N_15258);
and U19570 (N_19570,N_16224,N_15246);
xor U19571 (N_19571,N_17426,N_16760);
or U19572 (N_19572,N_15972,N_17168);
nor U19573 (N_19573,N_16214,N_17448);
xor U19574 (N_19574,N_15901,N_15413);
and U19575 (N_19575,N_15787,N_17061);
nand U19576 (N_19576,N_15285,N_16087);
or U19577 (N_19577,N_15286,N_15381);
nor U19578 (N_19578,N_16023,N_16150);
or U19579 (N_19579,N_16850,N_15143);
xor U19580 (N_19580,N_17220,N_16874);
nor U19581 (N_19581,N_16913,N_16050);
xor U19582 (N_19582,N_16050,N_15920);
nor U19583 (N_19583,N_16764,N_16731);
nand U19584 (N_19584,N_17338,N_16235);
xor U19585 (N_19585,N_16805,N_17121);
nand U19586 (N_19586,N_16143,N_15029);
nand U19587 (N_19587,N_17349,N_16488);
nand U19588 (N_19588,N_15617,N_16177);
nor U19589 (N_19589,N_15489,N_17375);
nor U19590 (N_19590,N_16870,N_16167);
nand U19591 (N_19591,N_17364,N_16641);
and U19592 (N_19592,N_16390,N_17026);
or U19593 (N_19593,N_16421,N_16933);
or U19594 (N_19594,N_16026,N_15206);
and U19595 (N_19595,N_17370,N_16022);
nand U19596 (N_19596,N_15703,N_15770);
or U19597 (N_19597,N_15442,N_16212);
nor U19598 (N_19598,N_15753,N_17360);
xor U19599 (N_19599,N_15453,N_15326);
or U19600 (N_19600,N_16623,N_16253);
xnor U19601 (N_19601,N_15830,N_17223);
and U19602 (N_19602,N_16452,N_16799);
or U19603 (N_19603,N_17263,N_16119);
or U19604 (N_19604,N_15918,N_15493);
or U19605 (N_19605,N_16013,N_17004);
nor U19606 (N_19606,N_17291,N_15907);
or U19607 (N_19607,N_15133,N_16765);
nor U19608 (N_19608,N_16299,N_16794);
nand U19609 (N_19609,N_16397,N_17390);
xnor U19610 (N_19610,N_16861,N_17227);
nand U19611 (N_19611,N_15358,N_15521);
nor U19612 (N_19612,N_16815,N_15375);
nor U19613 (N_19613,N_16883,N_17297);
and U19614 (N_19614,N_15760,N_17086);
or U19615 (N_19615,N_16082,N_16174);
nand U19616 (N_19616,N_15844,N_15691);
xnor U19617 (N_19617,N_17375,N_16629);
and U19618 (N_19618,N_16079,N_15265);
nor U19619 (N_19619,N_16819,N_17497);
or U19620 (N_19620,N_17123,N_16713);
and U19621 (N_19621,N_16517,N_15940);
nand U19622 (N_19622,N_16799,N_15680);
or U19623 (N_19623,N_17140,N_17465);
nand U19624 (N_19624,N_15596,N_16929);
xor U19625 (N_19625,N_15568,N_17204);
or U19626 (N_19626,N_17266,N_15700);
or U19627 (N_19627,N_16805,N_15206);
xnor U19628 (N_19628,N_15538,N_16628);
nand U19629 (N_19629,N_16128,N_15371);
nand U19630 (N_19630,N_16972,N_17316);
and U19631 (N_19631,N_15302,N_17254);
or U19632 (N_19632,N_16516,N_17176);
nor U19633 (N_19633,N_17142,N_17127);
and U19634 (N_19634,N_15105,N_15285);
and U19635 (N_19635,N_15451,N_15385);
nor U19636 (N_19636,N_16147,N_16125);
nand U19637 (N_19637,N_15349,N_16583);
xnor U19638 (N_19638,N_17032,N_15072);
and U19639 (N_19639,N_15323,N_16640);
nand U19640 (N_19640,N_16504,N_16930);
xnor U19641 (N_19641,N_17377,N_16942);
and U19642 (N_19642,N_16594,N_16533);
nor U19643 (N_19643,N_15694,N_15938);
nor U19644 (N_19644,N_16946,N_17204);
nor U19645 (N_19645,N_15015,N_15865);
xnor U19646 (N_19646,N_17313,N_17240);
and U19647 (N_19647,N_16468,N_15324);
xnor U19648 (N_19648,N_17196,N_17299);
nor U19649 (N_19649,N_15578,N_17105);
nor U19650 (N_19650,N_15646,N_17339);
nand U19651 (N_19651,N_16283,N_16539);
nand U19652 (N_19652,N_17199,N_16161);
xor U19653 (N_19653,N_16262,N_15692);
nand U19654 (N_19654,N_16046,N_16345);
nand U19655 (N_19655,N_17246,N_17358);
nor U19656 (N_19656,N_16923,N_15879);
and U19657 (N_19657,N_16290,N_15294);
nor U19658 (N_19658,N_15485,N_17088);
and U19659 (N_19659,N_16596,N_15813);
or U19660 (N_19660,N_16178,N_16701);
or U19661 (N_19661,N_15834,N_15745);
or U19662 (N_19662,N_16201,N_15480);
or U19663 (N_19663,N_16784,N_16681);
and U19664 (N_19664,N_16818,N_17052);
or U19665 (N_19665,N_15198,N_15595);
nor U19666 (N_19666,N_15557,N_15729);
and U19667 (N_19667,N_16693,N_16248);
or U19668 (N_19668,N_15250,N_16881);
xnor U19669 (N_19669,N_15192,N_15007);
nor U19670 (N_19670,N_15990,N_16893);
and U19671 (N_19671,N_17036,N_15471);
nand U19672 (N_19672,N_17487,N_17067);
xor U19673 (N_19673,N_16881,N_16247);
nor U19674 (N_19674,N_15552,N_15451);
or U19675 (N_19675,N_17152,N_15318);
nor U19676 (N_19676,N_16973,N_15869);
nand U19677 (N_19677,N_15830,N_17101);
xor U19678 (N_19678,N_15860,N_15222);
xnor U19679 (N_19679,N_16088,N_16411);
nand U19680 (N_19680,N_16195,N_15395);
or U19681 (N_19681,N_16587,N_15848);
nor U19682 (N_19682,N_15419,N_15445);
xnor U19683 (N_19683,N_16888,N_15729);
nor U19684 (N_19684,N_15399,N_15053);
nand U19685 (N_19685,N_16909,N_17169);
nand U19686 (N_19686,N_15177,N_15847);
or U19687 (N_19687,N_15765,N_16069);
nand U19688 (N_19688,N_17142,N_16898);
nand U19689 (N_19689,N_17153,N_15074);
or U19690 (N_19690,N_16875,N_16529);
xnor U19691 (N_19691,N_17070,N_16724);
nor U19692 (N_19692,N_17074,N_16452);
or U19693 (N_19693,N_17175,N_15733);
nand U19694 (N_19694,N_16524,N_15027);
nor U19695 (N_19695,N_16227,N_16815);
nor U19696 (N_19696,N_16428,N_15403);
nand U19697 (N_19697,N_15550,N_15802);
nor U19698 (N_19698,N_17088,N_16731);
xor U19699 (N_19699,N_16257,N_16040);
and U19700 (N_19700,N_15329,N_15781);
nor U19701 (N_19701,N_15899,N_15297);
nor U19702 (N_19702,N_15970,N_16789);
nor U19703 (N_19703,N_15798,N_15543);
and U19704 (N_19704,N_15497,N_16351);
or U19705 (N_19705,N_15605,N_17467);
xnor U19706 (N_19706,N_15962,N_16188);
or U19707 (N_19707,N_15725,N_16327);
nor U19708 (N_19708,N_17103,N_15491);
nor U19709 (N_19709,N_16246,N_16650);
nand U19710 (N_19710,N_16199,N_17183);
nor U19711 (N_19711,N_16537,N_16043);
nand U19712 (N_19712,N_16242,N_16923);
and U19713 (N_19713,N_17268,N_15046);
or U19714 (N_19714,N_15000,N_15631);
nand U19715 (N_19715,N_16842,N_15102);
nand U19716 (N_19716,N_15760,N_17427);
xor U19717 (N_19717,N_15057,N_16547);
nand U19718 (N_19718,N_16676,N_15508);
or U19719 (N_19719,N_17427,N_16867);
nand U19720 (N_19720,N_16363,N_15337);
and U19721 (N_19721,N_16966,N_16639);
nand U19722 (N_19722,N_15235,N_16187);
nor U19723 (N_19723,N_16297,N_15799);
nand U19724 (N_19724,N_16301,N_16694);
and U19725 (N_19725,N_16436,N_15581);
nand U19726 (N_19726,N_17243,N_16785);
xor U19727 (N_19727,N_15741,N_16144);
nor U19728 (N_19728,N_17115,N_16859);
or U19729 (N_19729,N_15458,N_15263);
nor U19730 (N_19730,N_16218,N_15201);
or U19731 (N_19731,N_15781,N_16019);
nand U19732 (N_19732,N_17308,N_15574);
xnor U19733 (N_19733,N_15374,N_15428);
xor U19734 (N_19734,N_16810,N_16481);
nand U19735 (N_19735,N_15295,N_16983);
nor U19736 (N_19736,N_16219,N_15610);
and U19737 (N_19737,N_15387,N_15211);
xnor U19738 (N_19738,N_16959,N_17411);
nand U19739 (N_19739,N_16861,N_15874);
or U19740 (N_19740,N_15033,N_17264);
and U19741 (N_19741,N_16927,N_15521);
nand U19742 (N_19742,N_16447,N_16729);
and U19743 (N_19743,N_15115,N_16857);
nor U19744 (N_19744,N_16694,N_17213);
and U19745 (N_19745,N_17001,N_16888);
and U19746 (N_19746,N_15190,N_15981);
nor U19747 (N_19747,N_16444,N_16251);
nor U19748 (N_19748,N_15561,N_15577);
nor U19749 (N_19749,N_15412,N_16474);
nand U19750 (N_19750,N_15980,N_17414);
xnor U19751 (N_19751,N_16187,N_16850);
and U19752 (N_19752,N_15602,N_15673);
nand U19753 (N_19753,N_17355,N_16356);
or U19754 (N_19754,N_17329,N_17132);
and U19755 (N_19755,N_16452,N_15164);
or U19756 (N_19756,N_17089,N_17361);
xnor U19757 (N_19757,N_15945,N_17149);
or U19758 (N_19758,N_16142,N_16865);
nor U19759 (N_19759,N_15905,N_15527);
or U19760 (N_19760,N_16626,N_15104);
or U19761 (N_19761,N_16823,N_16595);
nor U19762 (N_19762,N_16981,N_15066);
nand U19763 (N_19763,N_17360,N_15659);
and U19764 (N_19764,N_16499,N_16210);
nand U19765 (N_19765,N_16631,N_16930);
and U19766 (N_19766,N_15481,N_15773);
nor U19767 (N_19767,N_17247,N_17062);
nor U19768 (N_19768,N_15746,N_15755);
xnor U19769 (N_19769,N_16563,N_15385);
nand U19770 (N_19770,N_17014,N_16378);
or U19771 (N_19771,N_17367,N_17441);
nor U19772 (N_19772,N_15613,N_16892);
nand U19773 (N_19773,N_16846,N_15087);
or U19774 (N_19774,N_17157,N_15335);
or U19775 (N_19775,N_15742,N_16971);
nand U19776 (N_19776,N_15351,N_17368);
nand U19777 (N_19777,N_15971,N_15588);
and U19778 (N_19778,N_16765,N_17190);
xnor U19779 (N_19779,N_16471,N_16068);
nand U19780 (N_19780,N_15362,N_17065);
nand U19781 (N_19781,N_17364,N_16595);
nor U19782 (N_19782,N_16718,N_15908);
nand U19783 (N_19783,N_15256,N_16132);
and U19784 (N_19784,N_16509,N_16587);
and U19785 (N_19785,N_17075,N_16958);
nor U19786 (N_19786,N_16535,N_15319);
xor U19787 (N_19787,N_16903,N_15657);
and U19788 (N_19788,N_16428,N_17284);
nor U19789 (N_19789,N_16751,N_17123);
xor U19790 (N_19790,N_15798,N_15013);
nor U19791 (N_19791,N_15252,N_15033);
nor U19792 (N_19792,N_15457,N_15773);
nor U19793 (N_19793,N_16098,N_15590);
or U19794 (N_19794,N_16862,N_15733);
nor U19795 (N_19795,N_16300,N_15573);
nor U19796 (N_19796,N_16488,N_15830);
and U19797 (N_19797,N_15725,N_15056);
nand U19798 (N_19798,N_16750,N_15746);
nand U19799 (N_19799,N_16433,N_15372);
and U19800 (N_19800,N_15046,N_16563);
nor U19801 (N_19801,N_16101,N_17219);
and U19802 (N_19802,N_16448,N_16773);
nor U19803 (N_19803,N_15001,N_16078);
nor U19804 (N_19804,N_15407,N_16095);
or U19805 (N_19805,N_15275,N_15514);
or U19806 (N_19806,N_15240,N_15125);
nand U19807 (N_19807,N_17094,N_17462);
nand U19808 (N_19808,N_17472,N_16446);
nor U19809 (N_19809,N_15699,N_15603);
nor U19810 (N_19810,N_17011,N_16447);
and U19811 (N_19811,N_15296,N_17059);
nand U19812 (N_19812,N_17115,N_16149);
and U19813 (N_19813,N_15715,N_16534);
or U19814 (N_19814,N_16384,N_16094);
and U19815 (N_19815,N_15336,N_16896);
xnor U19816 (N_19816,N_15593,N_16646);
xnor U19817 (N_19817,N_15617,N_17219);
and U19818 (N_19818,N_15572,N_17208);
nand U19819 (N_19819,N_16152,N_17300);
or U19820 (N_19820,N_16695,N_17268);
nand U19821 (N_19821,N_17099,N_16774);
xor U19822 (N_19822,N_17375,N_16059);
or U19823 (N_19823,N_15550,N_15975);
nand U19824 (N_19824,N_15756,N_17196);
nand U19825 (N_19825,N_16895,N_15389);
xnor U19826 (N_19826,N_16598,N_16182);
and U19827 (N_19827,N_16739,N_16001);
xor U19828 (N_19828,N_16709,N_16597);
nor U19829 (N_19829,N_16261,N_15610);
and U19830 (N_19830,N_15121,N_17303);
nor U19831 (N_19831,N_15155,N_15003);
nand U19832 (N_19832,N_16179,N_15128);
or U19833 (N_19833,N_16989,N_16175);
nand U19834 (N_19834,N_16091,N_17310);
nand U19835 (N_19835,N_17041,N_16139);
xnor U19836 (N_19836,N_16716,N_16694);
nand U19837 (N_19837,N_15784,N_17494);
and U19838 (N_19838,N_15695,N_15811);
and U19839 (N_19839,N_16079,N_15536);
nand U19840 (N_19840,N_15834,N_17415);
xor U19841 (N_19841,N_17000,N_15655);
and U19842 (N_19842,N_16636,N_17007);
or U19843 (N_19843,N_17472,N_15202);
nor U19844 (N_19844,N_16204,N_16714);
and U19845 (N_19845,N_15733,N_16637);
nor U19846 (N_19846,N_15466,N_16358);
or U19847 (N_19847,N_16523,N_15657);
and U19848 (N_19848,N_16350,N_16593);
or U19849 (N_19849,N_16975,N_15999);
nor U19850 (N_19850,N_16594,N_15207);
or U19851 (N_19851,N_15358,N_17032);
xnor U19852 (N_19852,N_15411,N_15981);
xor U19853 (N_19853,N_16796,N_16277);
nor U19854 (N_19854,N_15137,N_15850);
and U19855 (N_19855,N_16890,N_15885);
xnor U19856 (N_19856,N_16256,N_16257);
xnor U19857 (N_19857,N_17488,N_17256);
xnor U19858 (N_19858,N_15845,N_16361);
and U19859 (N_19859,N_17413,N_16623);
or U19860 (N_19860,N_15432,N_16545);
xnor U19861 (N_19861,N_17405,N_16588);
or U19862 (N_19862,N_17264,N_15038);
and U19863 (N_19863,N_15165,N_17290);
nand U19864 (N_19864,N_17155,N_15610);
nor U19865 (N_19865,N_15214,N_15386);
xor U19866 (N_19866,N_15332,N_16140);
and U19867 (N_19867,N_16657,N_16473);
nor U19868 (N_19868,N_16037,N_16010);
xnor U19869 (N_19869,N_17040,N_16493);
nand U19870 (N_19870,N_15077,N_15080);
nand U19871 (N_19871,N_16850,N_15379);
nor U19872 (N_19872,N_15687,N_15219);
or U19873 (N_19873,N_15631,N_16579);
or U19874 (N_19874,N_15078,N_17195);
nand U19875 (N_19875,N_17113,N_15977);
or U19876 (N_19876,N_15197,N_15270);
or U19877 (N_19877,N_15195,N_16760);
or U19878 (N_19878,N_16176,N_15942);
nor U19879 (N_19879,N_15838,N_15197);
xnor U19880 (N_19880,N_15157,N_16671);
xnor U19881 (N_19881,N_15702,N_15002);
nand U19882 (N_19882,N_15627,N_15891);
nand U19883 (N_19883,N_17494,N_16874);
nand U19884 (N_19884,N_16548,N_16296);
nand U19885 (N_19885,N_16179,N_15950);
and U19886 (N_19886,N_16739,N_17400);
and U19887 (N_19887,N_15093,N_17328);
xnor U19888 (N_19888,N_15487,N_16934);
nand U19889 (N_19889,N_15676,N_16268);
or U19890 (N_19890,N_15173,N_17360);
nor U19891 (N_19891,N_16393,N_16352);
nand U19892 (N_19892,N_15167,N_15647);
or U19893 (N_19893,N_16379,N_16583);
xor U19894 (N_19894,N_15049,N_16131);
nor U19895 (N_19895,N_15549,N_15112);
nor U19896 (N_19896,N_15146,N_16992);
nand U19897 (N_19897,N_15313,N_17312);
or U19898 (N_19898,N_17442,N_17478);
and U19899 (N_19899,N_16649,N_17108);
nand U19900 (N_19900,N_15643,N_15911);
xnor U19901 (N_19901,N_17189,N_16880);
nand U19902 (N_19902,N_15628,N_15675);
and U19903 (N_19903,N_17104,N_16093);
or U19904 (N_19904,N_15610,N_16366);
and U19905 (N_19905,N_16039,N_15635);
nand U19906 (N_19906,N_16180,N_16311);
nand U19907 (N_19907,N_16233,N_16719);
nor U19908 (N_19908,N_15760,N_16195);
nand U19909 (N_19909,N_16597,N_16014);
and U19910 (N_19910,N_16425,N_16539);
nor U19911 (N_19911,N_16109,N_17011);
nor U19912 (N_19912,N_17499,N_16233);
xor U19913 (N_19913,N_16074,N_17477);
nor U19914 (N_19914,N_16937,N_16343);
nor U19915 (N_19915,N_16556,N_16857);
or U19916 (N_19916,N_16739,N_16202);
or U19917 (N_19917,N_16150,N_15688);
nand U19918 (N_19918,N_17178,N_16097);
or U19919 (N_19919,N_16226,N_16977);
xor U19920 (N_19920,N_15225,N_15984);
nor U19921 (N_19921,N_17010,N_17493);
and U19922 (N_19922,N_16791,N_17448);
and U19923 (N_19923,N_16717,N_15878);
and U19924 (N_19924,N_16516,N_15790);
and U19925 (N_19925,N_15896,N_17006);
and U19926 (N_19926,N_16352,N_17097);
nor U19927 (N_19927,N_17492,N_16831);
and U19928 (N_19928,N_15317,N_16863);
nor U19929 (N_19929,N_15531,N_17434);
nand U19930 (N_19930,N_15220,N_17171);
nor U19931 (N_19931,N_16347,N_15722);
xnor U19932 (N_19932,N_16618,N_15524);
nand U19933 (N_19933,N_15479,N_15280);
or U19934 (N_19934,N_16490,N_16099);
xor U19935 (N_19935,N_16112,N_16352);
nor U19936 (N_19936,N_16344,N_16081);
or U19937 (N_19937,N_16119,N_16874);
xor U19938 (N_19938,N_17345,N_16701);
or U19939 (N_19939,N_15135,N_16798);
nor U19940 (N_19940,N_15961,N_16237);
or U19941 (N_19941,N_16866,N_15955);
or U19942 (N_19942,N_17462,N_17214);
nor U19943 (N_19943,N_15648,N_16238);
or U19944 (N_19944,N_16836,N_16082);
xor U19945 (N_19945,N_17013,N_16869);
nor U19946 (N_19946,N_16849,N_16060);
or U19947 (N_19947,N_15924,N_16993);
and U19948 (N_19948,N_15872,N_16059);
or U19949 (N_19949,N_15956,N_16088);
nor U19950 (N_19950,N_17154,N_15986);
nor U19951 (N_19951,N_16951,N_15716);
xnor U19952 (N_19952,N_16769,N_16802);
and U19953 (N_19953,N_17103,N_15359);
or U19954 (N_19954,N_15389,N_15740);
nor U19955 (N_19955,N_15364,N_15872);
and U19956 (N_19956,N_15148,N_15533);
nand U19957 (N_19957,N_15062,N_15507);
or U19958 (N_19958,N_16621,N_16130);
xor U19959 (N_19959,N_16598,N_16737);
nand U19960 (N_19960,N_16878,N_15417);
or U19961 (N_19961,N_17154,N_15194);
or U19962 (N_19962,N_16853,N_16934);
nand U19963 (N_19963,N_15108,N_16334);
nor U19964 (N_19964,N_15833,N_17118);
and U19965 (N_19965,N_16215,N_15927);
nand U19966 (N_19966,N_15386,N_17047);
or U19967 (N_19967,N_16336,N_15917);
xor U19968 (N_19968,N_16698,N_17232);
nand U19969 (N_19969,N_16721,N_15951);
and U19970 (N_19970,N_15459,N_17343);
xor U19971 (N_19971,N_15790,N_16389);
nand U19972 (N_19972,N_16214,N_15488);
nor U19973 (N_19973,N_16231,N_15997);
xor U19974 (N_19974,N_15004,N_16197);
nand U19975 (N_19975,N_15010,N_16677);
xnor U19976 (N_19976,N_15681,N_16529);
xor U19977 (N_19977,N_16383,N_17366);
nand U19978 (N_19978,N_16856,N_17241);
xor U19979 (N_19979,N_15487,N_17317);
xnor U19980 (N_19980,N_17265,N_15774);
nor U19981 (N_19981,N_17204,N_15491);
nor U19982 (N_19982,N_15320,N_17194);
or U19983 (N_19983,N_15734,N_16064);
xnor U19984 (N_19984,N_16091,N_16728);
nand U19985 (N_19985,N_17349,N_16991);
and U19986 (N_19986,N_16390,N_15206);
nor U19987 (N_19987,N_15150,N_16246);
or U19988 (N_19988,N_16890,N_15191);
nand U19989 (N_19989,N_15637,N_16004);
nor U19990 (N_19990,N_15258,N_15158);
nand U19991 (N_19991,N_16297,N_15952);
or U19992 (N_19992,N_15118,N_16624);
xor U19993 (N_19993,N_15905,N_16758);
or U19994 (N_19994,N_15798,N_16294);
and U19995 (N_19995,N_15739,N_16930);
or U19996 (N_19996,N_15705,N_16565);
xnor U19997 (N_19997,N_16080,N_15950);
or U19998 (N_19998,N_16909,N_16513);
and U19999 (N_19999,N_15956,N_16052);
or U20000 (N_20000,N_19647,N_18762);
nor U20001 (N_20001,N_19593,N_19304);
nor U20002 (N_20002,N_17871,N_19709);
and U20003 (N_20003,N_18513,N_19004);
and U20004 (N_20004,N_18764,N_19364);
or U20005 (N_20005,N_18486,N_19118);
and U20006 (N_20006,N_19038,N_18353);
nor U20007 (N_20007,N_19149,N_18897);
nand U20008 (N_20008,N_18859,N_18545);
and U20009 (N_20009,N_19099,N_18450);
nand U20010 (N_20010,N_18958,N_19691);
or U20011 (N_20011,N_18081,N_19505);
xor U20012 (N_20012,N_19035,N_17708);
nor U20013 (N_20013,N_19386,N_19240);
and U20014 (N_20014,N_18084,N_17959);
and U20015 (N_20015,N_17832,N_18993);
xor U20016 (N_20016,N_19881,N_17789);
xor U20017 (N_20017,N_17926,N_19447);
nand U20018 (N_20018,N_18593,N_19820);
or U20019 (N_20019,N_17684,N_19028);
xor U20020 (N_20020,N_19520,N_18594);
nand U20021 (N_20021,N_19581,N_18138);
or U20022 (N_20022,N_19070,N_19419);
xor U20023 (N_20023,N_19341,N_17575);
or U20024 (N_20024,N_18905,N_18273);
and U20025 (N_20025,N_19395,N_19170);
or U20026 (N_20026,N_18526,N_19915);
nor U20027 (N_20027,N_18225,N_18003);
nor U20028 (N_20028,N_18759,N_19237);
and U20029 (N_20029,N_17605,N_19279);
xnor U20030 (N_20030,N_17515,N_18773);
or U20031 (N_20031,N_18504,N_18153);
nor U20032 (N_20032,N_17770,N_19867);
xnor U20033 (N_20033,N_19904,N_19354);
nor U20034 (N_20034,N_18757,N_17991);
xnor U20035 (N_20035,N_19791,N_18396);
nor U20036 (N_20036,N_18063,N_19229);
and U20037 (N_20037,N_18795,N_17651);
nand U20038 (N_20038,N_19834,N_19203);
nor U20039 (N_20039,N_18419,N_18917);
nor U20040 (N_20040,N_17799,N_18567);
nor U20041 (N_20041,N_19734,N_18972);
or U20042 (N_20042,N_19355,N_17960);
or U20043 (N_20043,N_17934,N_17969);
xnor U20044 (N_20044,N_18343,N_19797);
xnor U20045 (N_20045,N_17933,N_19199);
nor U20046 (N_20046,N_18695,N_19625);
and U20047 (N_20047,N_19649,N_19913);
xnor U20048 (N_20048,N_19608,N_17633);
and U20049 (N_20049,N_18840,N_19343);
nor U20050 (N_20050,N_17907,N_19269);
xnor U20051 (N_20051,N_18102,N_18448);
nand U20052 (N_20052,N_18591,N_19227);
or U20053 (N_20053,N_19092,N_18838);
or U20054 (N_20054,N_18914,N_18541);
or U20055 (N_20055,N_17553,N_19376);
nand U20056 (N_20056,N_19214,N_19755);
and U20057 (N_20057,N_18600,N_18103);
and U20058 (N_20058,N_18921,N_17608);
xor U20059 (N_20059,N_19638,N_17796);
nor U20060 (N_20060,N_18203,N_19049);
or U20061 (N_20061,N_18809,N_17518);
and U20062 (N_20062,N_17771,N_19827);
or U20063 (N_20063,N_18888,N_19885);
and U20064 (N_20064,N_19995,N_18324);
nand U20065 (N_20065,N_18024,N_18642);
xnor U20066 (N_20066,N_18853,N_17929);
or U20067 (N_20067,N_18312,N_17635);
and U20068 (N_20068,N_19346,N_19730);
nor U20069 (N_20069,N_17571,N_18633);
nand U20070 (N_20070,N_17587,N_17947);
nor U20071 (N_20071,N_19333,N_17677);
nand U20072 (N_20072,N_18061,N_18575);
and U20073 (N_20073,N_18330,N_17893);
nand U20074 (N_20074,N_19620,N_18099);
or U20075 (N_20075,N_18716,N_19851);
or U20076 (N_20076,N_18604,N_18841);
nand U20077 (N_20077,N_19445,N_17722);
and U20078 (N_20078,N_19598,N_19017);
and U20079 (N_20079,N_19729,N_19935);
nor U20080 (N_20080,N_18756,N_19008);
nor U20081 (N_20081,N_18007,N_18493);
xor U20082 (N_20082,N_18965,N_18667);
nor U20083 (N_20083,N_17631,N_19241);
and U20084 (N_20084,N_18162,N_19921);
xnor U20085 (N_20085,N_19251,N_17646);
or U20086 (N_20086,N_19690,N_18665);
nand U20087 (N_20087,N_19969,N_18498);
or U20088 (N_20088,N_18488,N_19473);
xnor U20089 (N_20089,N_17577,N_19694);
xor U20090 (N_20090,N_19806,N_19781);
nor U20091 (N_20091,N_19145,N_17510);
nor U20092 (N_20092,N_19999,N_18360);
nor U20093 (N_20093,N_19086,N_17639);
xor U20094 (N_20094,N_17804,N_17552);
nand U20095 (N_20095,N_19223,N_18345);
nor U20096 (N_20096,N_19385,N_19786);
xnor U20097 (N_20097,N_17533,N_18868);
and U20098 (N_20098,N_17966,N_18266);
xnor U20099 (N_20099,N_18098,N_19964);
nor U20100 (N_20100,N_17746,N_18248);
nand U20101 (N_20101,N_18967,N_19330);
and U20102 (N_20102,N_17989,N_19809);
nand U20103 (N_20103,N_19011,N_17671);
nor U20104 (N_20104,N_17936,N_19356);
and U20105 (N_20105,N_18984,N_18451);
and U20106 (N_20106,N_17974,N_19607);
and U20107 (N_20107,N_19181,N_19126);
or U20108 (N_20108,N_18160,N_18124);
nand U20109 (N_20109,N_19158,N_19496);
or U20110 (N_20110,N_18246,N_19094);
or U20111 (N_20111,N_19313,N_18692);
xor U20112 (N_20112,N_18672,N_18645);
xnor U20113 (N_20113,N_18707,N_19077);
nor U20114 (N_20114,N_18350,N_17938);
and U20115 (N_20115,N_19772,N_18851);
and U20116 (N_20116,N_17810,N_18915);
nand U20117 (N_20117,N_19048,N_19568);
and U20118 (N_20118,N_19169,N_18318);
nand U20119 (N_20119,N_19225,N_19262);
nor U20120 (N_20120,N_17923,N_17693);
or U20121 (N_20121,N_18104,N_18443);
and U20122 (N_20122,N_19379,N_19538);
nor U20123 (N_20123,N_19483,N_18569);
nor U20124 (N_20124,N_19105,N_19571);
or U20125 (N_20125,N_19578,N_18338);
nor U20126 (N_20126,N_18887,N_19098);
or U20127 (N_20127,N_18306,N_18603);
or U20128 (N_20128,N_18106,N_17738);
nand U20129 (N_20129,N_19308,N_17763);
or U20130 (N_20130,N_19679,N_18482);
nor U20131 (N_20131,N_17852,N_19034);
nor U20132 (N_20132,N_19790,N_18787);
and U20133 (N_20133,N_17669,N_18189);
and U20134 (N_20134,N_19219,N_17697);
and U20135 (N_20135,N_17995,N_19173);
or U20136 (N_20136,N_19479,N_18108);
nor U20137 (N_20137,N_19465,N_19688);
xnor U20138 (N_20138,N_18211,N_17909);
or U20139 (N_20139,N_18854,N_18147);
xor U20140 (N_20140,N_18676,N_18464);
xnor U20141 (N_20141,N_18798,N_19397);
nand U20142 (N_20142,N_19146,N_19622);
nor U20143 (N_20143,N_17534,N_19193);
and U20144 (N_20144,N_18073,N_18959);
or U20145 (N_20145,N_19838,N_18122);
and U20146 (N_20146,N_18332,N_19616);
nor U20147 (N_20147,N_19537,N_19366);
nor U20148 (N_20148,N_18363,N_19165);
and U20149 (N_20149,N_18936,N_18462);
nor U20150 (N_20150,N_18290,N_19114);
and U20151 (N_20151,N_19669,N_19585);
and U20152 (N_20152,N_18060,N_17987);
nand U20153 (N_20153,N_18974,N_19916);
nor U20154 (N_20154,N_17656,N_18932);
nand U20155 (N_20155,N_19026,N_19660);
and U20156 (N_20156,N_19093,N_18496);
nor U20157 (N_20157,N_19492,N_18518);
and U20158 (N_20158,N_17822,N_18207);
or U20159 (N_20159,N_18849,N_19962);
and U20160 (N_20160,N_18085,N_19189);
or U20161 (N_20161,N_19681,N_19221);
xor U20162 (N_20162,N_18348,N_19716);
nand U20163 (N_20163,N_18319,N_18292);
xnor U20164 (N_20164,N_19942,N_17741);
nand U20165 (N_20165,N_18166,N_18521);
xor U20166 (N_20166,N_19176,N_18352);
nand U20167 (N_20167,N_18571,N_18452);
or U20168 (N_20168,N_18572,N_18376);
xor U20169 (N_20169,N_19481,N_18680);
or U20170 (N_20170,N_18337,N_18458);
nor U20171 (N_20171,N_19958,N_18421);
or U20172 (N_20172,N_18816,N_17815);
nor U20173 (N_20173,N_19432,N_17841);
nand U20174 (N_20174,N_19551,N_18922);
and U20175 (N_20175,N_19844,N_19557);
and U20176 (N_20176,N_19287,N_17891);
or U20177 (N_20177,N_19334,N_18322);
xnor U20178 (N_20178,N_17848,N_18815);
and U20179 (N_20179,N_18194,N_18091);
nand U20180 (N_20180,N_17953,N_19980);
nor U20181 (N_20181,N_19052,N_19183);
and U20182 (N_20182,N_17568,N_18725);
or U20183 (N_20183,N_18192,N_18434);
nand U20184 (N_20184,N_19946,N_18274);
or U20185 (N_20185,N_19808,N_19769);
nand U20186 (N_20186,N_17686,N_17823);
xnor U20187 (N_20187,N_18739,N_18430);
nor U20188 (N_20188,N_19847,N_19591);
nor U20189 (N_20189,N_18837,N_19406);
or U20190 (N_20190,N_17973,N_17798);
or U20191 (N_20191,N_17890,N_18694);
nor U20192 (N_20192,N_17692,N_19894);
nand U20193 (N_20193,N_18889,N_19083);
and U20194 (N_20194,N_17759,N_19078);
nand U20195 (N_20195,N_18049,N_18152);
nor U20196 (N_20196,N_18599,N_18528);
nor U20197 (N_20197,N_18018,N_19517);
or U20198 (N_20198,N_18659,N_18782);
nand U20199 (N_20199,N_17522,N_17845);
and U20200 (N_20200,N_18797,N_17607);
nor U20201 (N_20201,N_17531,N_17551);
or U20202 (N_20202,N_19728,N_19140);
and U20203 (N_20203,N_19208,N_19336);
and U20204 (N_20204,N_19668,N_17548);
nand U20205 (N_20205,N_17942,N_17570);
or U20206 (N_20206,N_18856,N_18247);
xnor U20207 (N_20207,N_18015,N_18093);
or U20208 (N_20208,N_19985,N_18052);
nor U20209 (N_20209,N_18503,N_18813);
xor U20210 (N_20210,N_19527,N_18064);
nor U20211 (N_20211,N_19804,N_17831);
and U20212 (N_20212,N_18080,N_18200);
nor U20213 (N_20213,N_18529,N_18260);
and U20214 (N_20214,N_17648,N_19006);
nand U20215 (N_20215,N_19119,N_19878);
and U20216 (N_20216,N_19554,N_18834);
nand U20217 (N_20217,N_19039,N_17644);
nor U20218 (N_20218,N_17743,N_18620);
nand U20219 (N_20219,N_18492,N_18185);
xnor U20220 (N_20220,N_19502,N_18407);
and U20221 (N_20221,N_19375,N_18723);
nor U20222 (N_20222,N_18298,N_18127);
nor U20223 (N_20223,N_17512,N_18953);
nor U20224 (N_20224,N_19320,N_17613);
and U20225 (N_20225,N_19778,N_18997);
or U20226 (N_20226,N_19563,N_18516);
or U20227 (N_20227,N_19053,N_18677);
or U20228 (N_20228,N_19702,N_19205);
nand U20229 (N_20229,N_19139,N_19212);
and U20230 (N_20230,N_17561,N_17598);
nand U20231 (N_20231,N_18955,N_19819);
or U20232 (N_20232,N_18807,N_19795);
or U20233 (N_20233,N_18901,N_17785);
xor U20234 (N_20234,N_19337,N_19978);
xnor U20235 (N_20235,N_18201,N_19949);
xor U20236 (N_20236,N_17961,N_17612);
or U20237 (N_20237,N_18041,N_18611);
xor U20238 (N_20238,N_17970,N_18040);
nor U20239 (N_20239,N_18001,N_19166);
nor U20240 (N_20240,N_17833,N_17526);
or U20241 (N_20241,N_19204,N_19762);
nand U20242 (N_20242,N_19849,N_19384);
xnor U20243 (N_20243,N_18476,N_17630);
and U20244 (N_20244,N_18674,N_19324);
nor U20245 (N_20245,N_19884,N_19986);
or U20246 (N_20246,N_19905,N_19144);
nand U20247 (N_20247,N_18525,N_18562);
nand U20248 (N_20248,N_18708,N_18555);
xor U20249 (N_20249,N_17769,N_18475);
and U20250 (N_20250,N_19388,N_18195);
and U20251 (N_20251,N_19367,N_19218);
nor U20252 (N_20252,N_18923,N_18069);
and U20253 (N_20253,N_19016,N_17728);
or U20254 (N_20254,N_17749,N_19877);
nand U20255 (N_20255,N_19564,N_19007);
xnor U20256 (N_20256,N_19064,N_17811);
nand U20257 (N_20257,N_19464,N_19882);
and U20258 (N_20258,N_19045,N_18497);
or U20259 (N_20259,N_17556,N_17788);
or U20260 (N_20260,N_19518,N_18748);
nor U20261 (N_20261,N_19676,N_17826);
and U20262 (N_20262,N_19233,N_18262);
nor U20263 (N_20263,N_19420,N_18563);
nor U20264 (N_20264,N_18855,N_17589);
or U20265 (N_20265,N_19823,N_18373);
or U20266 (N_20266,N_19689,N_18005);
and U20267 (N_20267,N_19113,N_17886);
and U20268 (N_20268,N_18020,N_18613);
nand U20269 (N_20269,N_18418,N_18654);
xor U20270 (N_20270,N_18301,N_18786);
and U20271 (N_20271,N_18397,N_19899);
and U20272 (N_20272,N_19186,N_17844);
and U20273 (N_20273,N_19135,N_18367);
xor U20274 (N_20274,N_18120,N_18158);
and U20275 (N_20275,N_19010,N_18022);
and U20276 (N_20276,N_18805,N_19635);
nand U20277 (N_20277,N_19238,N_18547);
nor U20278 (N_20278,N_18954,N_18852);
nor U20279 (N_20279,N_18271,N_18589);
and U20280 (N_20280,N_19580,N_19589);
nand U20281 (N_20281,N_18758,N_19658);
nor U20282 (N_20282,N_19352,N_18187);
and U20283 (N_20283,N_19439,N_18011);
nor U20284 (N_20284,N_18414,N_17935);
xnor U20285 (N_20285,N_18025,N_19036);
nor U20286 (N_20286,N_19096,N_19061);
nor U20287 (N_20287,N_19232,N_18232);
or U20288 (N_20288,N_17661,N_19023);
and U20289 (N_20289,N_18255,N_18919);
nand U20290 (N_20290,N_17972,N_18117);
and U20291 (N_20291,N_18027,N_17597);
or U20292 (N_20292,N_19652,N_19091);
and U20293 (N_20293,N_18871,N_19182);
nand U20294 (N_20294,N_17807,N_18895);
and U20295 (N_20295,N_17812,N_17547);
nand U20296 (N_20296,N_18270,N_19046);
nand U20297 (N_20297,N_18754,N_19503);
nor U20298 (N_20298,N_19727,N_19952);
nand U20299 (N_20299,N_17920,N_19879);
and U20300 (N_20300,N_19783,N_19258);
and U20301 (N_20301,N_19714,N_18539);
or U20302 (N_20302,N_18087,N_19471);
nor U20303 (N_20303,N_18426,N_19609);
xor U20304 (N_20304,N_19110,N_19852);
or U20305 (N_20305,N_19903,N_18944);
or U20306 (N_20306,N_19424,N_18487);
and U20307 (N_20307,N_19543,N_17640);
and U20308 (N_20308,N_19531,N_18265);
nor U20309 (N_20309,N_17544,N_19866);
nand U20310 (N_20310,N_19873,N_18438);
or U20311 (N_20311,N_19472,N_19611);
nand U20312 (N_20312,N_17899,N_18622);
or U20313 (N_20313,N_18241,N_19937);
nand U20314 (N_20314,N_19908,N_19216);
nand U20315 (N_20315,N_19850,N_17723);
nand U20316 (N_20316,N_17990,N_18259);
nor U20317 (N_20317,N_19614,N_18808);
xnor U20318 (N_20318,N_19288,N_18258);
and U20319 (N_20319,N_19577,N_18735);
or U20320 (N_20320,N_19927,N_19696);
xnor U20321 (N_20321,N_18245,N_19103);
nand U20322 (N_20322,N_19970,N_19900);
xnor U20323 (N_20323,N_19255,N_18931);
nand U20324 (N_20324,N_17965,N_19357);
or U20325 (N_20325,N_17914,N_19256);
and U20326 (N_20326,N_17932,N_17527);
xor U20327 (N_20327,N_17790,N_18314);
nand U20328 (N_20328,N_18055,N_19111);
and U20329 (N_20329,N_19310,N_19475);
nand U20330 (N_20330,N_18964,N_17637);
xnor U20331 (N_20331,N_18910,N_18962);
or U20332 (N_20332,N_19068,N_19154);
nor U20333 (N_20333,N_19138,N_18721);
nand U20334 (N_20334,N_18354,N_19012);
xnor U20335 (N_20335,N_19009,N_19841);
or U20336 (N_20336,N_18308,N_18862);
xor U20337 (N_20337,N_17817,N_19508);
and U20338 (N_20338,N_18508,N_19121);
nor U20339 (N_20339,N_18199,N_18736);
nand U20340 (N_20340,N_18234,N_18119);
or U20341 (N_20341,N_17501,N_17601);
nor U20342 (N_20342,N_18489,N_18254);
and U20343 (N_20343,N_19041,N_19090);
or U20344 (N_20344,N_17949,N_17869);
nor U20345 (N_20345,N_19044,N_18179);
and U20346 (N_20346,N_18347,N_19329);
xor U20347 (N_20347,N_18926,N_17761);
and U20348 (N_20348,N_19956,N_18644);
nor U20349 (N_20349,N_19236,N_19749);
xor U20350 (N_20350,N_18577,N_17791);
xor U20351 (N_20351,N_18899,N_19559);
nor U20352 (N_20352,N_18941,N_19737);
or U20353 (N_20353,N_17997,N_19360);
xor U20354 (N_20354,N_19271,N_17619);
and U20355 (N_20355,N_17576,N_18067);
or U20356 (N_20356,N_18738,N_18249);
or U20357 (N_20357,N_18357,N_19402);
xor U20358 (N_20358,N_19190,N_17955);
and U20359 (N_20359,N_19686,N_17895);
or U20360 (N_20360,N_19283,N_18453);
xnor U20361 (N_20361,N_19415,N_19639);
nor U20362 (N_20362,N_19678,N_18942);
nor U20363 (N_20363,N_17710,N_18113);
or U20364 (N_20364,N_18131,N_18639);
nor U20365 (N_20365,N_19319,N_19461);
and U20366 (N_20366,N_19859,N_19124);
and U20367 (N_20367,N_18057,N_19861);
nor U20368 (N_20368,N_17540,N_19327);
nand U20369 (N_20369,N_18500,N_17808);
or U20370 (N_20370,N_19756,N_18637);
nand U20371 (N_20371,N_18172,N_18765);
and U20372 (N_20372,N_17611,N_18217);
xor U20373 (N_20373,N_18679,N_19810);
nand U20374 (N_20374,N_17919,N_19477);
xnor U20375 (N_20375,N_17861,N_18750);
nand U20376 (N_20376,N_18802,N_18311);
and U20377 (N_20377,N_18145,N_19440);
nand U20378 (N_20378,N_19513,N_19380);
nor U20379 (N_20379,N_19846,N_19309);
and U20380 (N_20380,N_18075,N_18522);
or U20381 (N_20381,N_19249,N_17504);
xor U20382 (N_20382,N_18356,N_18929);
xor U20383 (N_20383,N_18326,N_17857);
xnor U20384 (N_20384,N_18398,N_18523);
and U20385 (N_20385,N_17560,N_17780);
or U20386 (N_20386,N_17843,N_18641);
xor U20387 (N_20387,N_19944,N_18596);
xnor U20388 (N_20388,N_17979,N_18540);
nor U20389 (N_20389,N_19719,N_18150);
nor U20390 (N_20390,N_18304,N_17657);
xnor U20391 (N_20391,N_19405,N_17873);
or U20392 (N_20392,N_19892,N_18030);
or U20393 (N_20393,N_19939,N_18601);
or U20394 (N_20394,N_18607,N_19742);
nor U20395 (N_20395,N_18874,N_19664);
xnor U20396 (N_20396,N_18714,N_18006);
nand U20397 (N_20397,N_17505,N_19192);
nor U20398 (N_20398,N_17537,N_19316);
and U20399 (N_20399,N_18656,N_18047);
xor U20400 (N_20400,N_18973,N_19632);
or U20401 (N_20401,N_18702,N_19566);
or U20402 (N_20402,N_19315,N_18392);
xnor U20403 (N_20403,N_17580,N_17525);
nand U20404 (N_20404,N_19750,N_18843);
or U20405 (N_20405,N_17839,N_18502);
nand U20406 (N_20406,N_19824,N_18517);
nor U20407 (N_20407,N_18631,N_18191);
xor U20408 (N_20408,N_17529,N_19770);
nand U20409 (N_20409,N_18817,N_19943);
nand U20410 (N_20410,N_18527,N_19383);
or U20411 (N_20411,N_19526,N_19751);
and U20412 (N_20412,N_18902,N_18062);
nor U20413 (N_20413,N_19621,N_17878);
xnor U20414 (N_20414,N_19148,N_17930);
nand U20415 (N_20415,N_18729,N_17666);
xor U20416 (N_20416,N_19230,N_19662);
nand U20417 (N_20417,N_18629,N_18013);
or U20418 (N_20418,N_19997,N_19082);
or U20419 (N_20419,N_18302,N_17765);
and U20420 (N_20420,N_19821,N_19529);
xnor U20421 (N_20421,N_17888,N_19798);
or U20422 (N_20422,N_18740,N_18088);
nand U20423 (N_20423,N_18950,N_18380);
or U20424 (N_20424,N_19276,N_18197);
and U20425 (N_20425,N_18437,N_19080);
nor U20426 (N_20426,N_19188,N_17752);
or U20427 (N_20427,N_18588,N_18114);
xnor U20428 (N_20428,N_19224,N_19371);
nor U20429 (N_20429,N_17818,N_19282);
nand U20430 (N_20430,N_18243,N_19648);
and U20431 (N_20431,N_17800,N_18479);
nand U20432 (N_20432,N_19084,N_19855);
xnor U20433 (N_20433,N_19131,N_18749);
or U20434 (N_20434,N_17764,N_19129);
or U20435 (N_20435,N_18379,N_18580);
or U20436 (N_20436,N_19239,N_19705);
and U20437 (N_20437,N_18351,N_17623);
and U20438 (N_20438,N_17721,N_18385);
nor U20439 (N_20439,N_18130,N_18206);
nand U20440 (N_20440,N_19427,N_19801);
nor U20441 (N_20441,N_18573,N_19839);
and U20442 (N_20442,N_19707,N_17578);
nor U20443 (N_20443,N_19923,N_18945);
nor U20444 (N_20444,N_18193,N_19670);
nand U20445 (N_20445,N_18995,N_17543);
xor U20446 (N_20446,N_18442,N_19579);
and U20447 (N_20447,N_18628,N_19180);
and U20448 (N_20448,N_18157,N_18826);
or U20449 (N_20449,N_18850,N_18515);
nand U20450 (N_20450,N_17829,N_18939);
nand U20451 (N_20451,N_18980,N_18619);
xnor U20452 (N_20452,N_18909,N_18866);
xor U20453 (N_20453,N_18257,N_17588);
nor U20454 (N_20454,N_19914,N_19722);
nor U20455 (N_20455,N_17803,N_18039);
nand U20456 (N_20456,N_19582,N_17582);
nand U20457 (N_20457,N_19274,N_19710);
nand U20458 (N_20458,N_19184,N_17736);
nor U20459 (N_20459,N_17870,N_19072);
or U20460 (N_20460,N_19667,N_19263);
nor U20461 (N_20461,N_19576,N_19700);
nor U20462 (N_20462,N_18724,N_19079);
or U20463 (N_20463,N_18556,N_19156);
and U20464 (N_20464,N_19983,N_18284);
and U20465 (N_20465,N_19553,N_17688);
nand U20466 (N_20466,N_19740,N_18457);
nand U20467 (N_20467,N_19698,N_17549);
xnor U20468 (N_20468,N_19171,N_18038);
xnor U20469 (N_20469,N_19437,N_19717);
nand U20470 (N_20470,N_18956,N_17735);
xor U20471 (N_20471,N_19374,N_18574);
or U20472 (N_20472,N_19209,N_17984);
nand U20473 (N_20473,N_19275,N_19168);
or U20474 (N_20474,N_18144,N_18399);
nand U20475 (N_20475,N_17659,N_19817);
xnor U20476 (N_20476,N_18632,N_18918);
or U20477 (N_20477,N_17680,N_18550);
or U20478 (N_20478,N_19054,N_18638);
and U20479 (N_20479,N_18002,N_19594);
or U20480 (N_20480,N_19711,N_18537);
xor U20481 (N_20481,N_17734,N_19555);
nand U20482 (N_20482,N_18531,N_19252);
or U20483 (N_20483,N_18657,N_18673);
and U20484 (N_20484,N_19488,N_18420);
or U20485 (N_20485,N_18661,N_17517);
or U20486 (N_20486,N_19869,N_17703);
nor U20487 (N_20487,N_18029,N_17977);
nor U20488 (N_20488,N_18658,N_19818);
or U20489 (N_20489,N_19194,N_17528);
xor U20490 (N_20490,N_19501,N_17624);
nand U20491 (N_20491,N_19974,N_18101);
xor U20492 (N_20492,N_19883,N_19491);
nor U20493 (N_20493,N_17539,N_18244);
or U20494 (N_20494,N_18204,N_18021);
and U20495 (N_20495,N_18210,N_18788);
nand U20496 (N_20496,N_18044,N_18263);
nand U20497 (N_20497,N_19998,N_18136);
nor U20498 (N_20498,N_17868,N_19117);
nor U20499 (N_20499,N_18100,N_19947);
nand U20500 (N_20500,N_18783,N_19458);
xnor U20501 (N_20501,N_19550,N_19665);
or U20502 (N_20502,N_19141,N_18986);
and U20503 (N_20503,N_19875,N_17975);
nand U20504 (N_20504,N_19907,N_17634);
nand U20505 (N_20505,N_19112,N_19836);
xor U20506 (N_20506,N_18911,N_18221);
or U20507 (N_20507,N_17720,N_18161);
and U20508 (N_20508,N_18128,N_18461);
or U20509 (N_20509,N_19792,N_18146);
or U20510 (N_20510,N_17879,N_19301);
nand U20511 (N_20511,N_19626,N_17787);
nor U20512 (N_20512,N_18474,N_18096);
or U20513 (N_20513,N_19030,N_19570);
nand U20514 (N_20514,N_18427,N_19215);
or U20515 (N_20515,N_19630,N_19924);
nor U20516 (N_20516,N_18282,N_18176);
or U20517 (N_20517,N_18239,N_19217);
nor U20518 (N_20518,N_19802,N_19246);
nand U20519 (N_20519,N_18801,N_18510);
xor U20520 (N_20520,N_19683,N_18987);
nor U20521 (N_20521,N_17921,N_18937);
or U20522 (N_20522,N_17511,N_19636);
nor U20523 (N_20523,N_18791,N_17779);
nor U20524 (N_20524,N_18804,N_18336);
and U20525 (N_20525,N_19605,N_18829);
nor U20526 (N_20526,N_17711,N_17795);
or U20527 (N_20527,N_18223,N_19462);
xnor U20528 (N_20528,N_17705,N_18960);
xor U20529 (N_20529,N_18690,N_18346);
and U20530 (N_20530,N_18183,N_18032);
nand U20531 (N_20531,N_19687,N_19389);
or U20532 (N_20532,N_18483,N_18220);
xor U20533 (N_20533,N_18307,N_18159);
xor U20534 (N_20534,N_18689,N_19767);
and U20535 (N_20535,N_18325,N_19441);
nand U20536 (N_20536,N_17821,N_19919);
nand U20537 (N_20537,N_18383,N_19785);
nor U20538 (N_20538,N_17753,N_18957);
nand U20539 (N_20539,N_17726,N_19911);
nand U20540 (N_20540,N_18610,N_18703);
nor U20541 (N_20541,N_17647,N_19805);
nor U20542 (N_20542,N_17794,N_19430);
xnor U20543 (N_20543,N_19766,N_19773);
and U20544 (N_20544,N_18137,N_19932);
or U20545 (N_20545,N_18683,N_18751);
nand U20546 (N_20546,N_19452,N_19264);
xor U20547 (N_20547,N_18507,N_19549);
and U20548 (N_20548,N_17892,N_18691);
xnor U20549 (N_20549,N_17913,N_19597);
xor U20550 (N_20550,N_18530,N_18256);
nand U20551 (N_20551,N_19459,N_18700);
nand U20552 (N_20552,N_17658,N_18519);
xnor U20553 (N_20553,N_19993,N_18329);
or U20554 (N_20554,N_19005,N_18916);
and U20555 (N_20555,N_19268,N_19654);
nor U20556 (N_20556,N_17797,N_17632);
nand U20557 (N_20557,N_17963,N_17558);
nor U20558 (N_20558,N_19468,N_17856);
and U20559 (N_20559,N_18818,N_18640);
xnor U20560 (N_20560,N_19069,N_18552);
nand U20561 (N_20561,N_18675,N_19469);
nand U20562 (N_20562,N_17566,N_17766);
and U20563 (N_20563,N_19032,N_19735);
xor U20564 (N_20564,N_18592,N_19401);
and U20565 (N_20565,N_19177,N_18753);
nor U20566 (N_20566,N_18491,N_17653);
and U20567 (N_20567,N_18920,N_17675);
xnor U20568 (N_20568,N_17751,N_18320);
xnor U20569 (N_20569,N_19895,N_19422);
xor U20570 (N_20570,N_18083,N_19901);
and U20571 (N_20571,N_18174,N_18961);
and U20572 (N_20572,N_18963,N_19431);
or U20573 (N_20573,N_17678,N_17816);
xor U20574 (N_20574,N_19507,N_19267);
xnor U20575 (N_20575,N_18092,N_19412);
or U20576 (N_20576,N_17971,N_18026);
and U20577 (N_20577,N_19929,N_17951);
xor U20578 (N_20578,N_19733,N_17875);
and U20579 (N_20579,N_18549,N_18439);
xor U20580 (N_20580,N_19228,N_19590);
and U20581 (N_20581,N_18297,N_19066);
nand U20582 (N_20582,N_18216,N_18303);
nor U20583 (N_20583,N_19033,N_19601);
nor U20584 (N_20584,N_17625,N_19051);
xnor U20585 (N_20585,N_19484,N_19396);
and U20586 (N_20586,N_17636,N_18698);
xor U20587 (N_20587,N_18180,N_19782);
xnor U20588 (N_20588,N_18167,N_18891);
nor U20589 (N_20589,N_19754,N_19934);
and U20590 (N_20590,N_17778,N_19522);
nand U20591 (N_20591,N_19572,N_19021);
nor U20592 (N_20592,N_17682,N_19592);
and U20593 (N_20593,N_17617,N_18940);
or U20594 (N_20594,N_19617,N_17719);
nand U20595 (N_20595,N_18328,N_19387);
nor U20596 (N_20596,N_19443,N_18048);
or U20597 (N_20597,N_18996,N_17604);
nand U20598 (N_20598,N_18317,N_19506);
nand U20599 (N_20599,N_18171,N_19351);
nor U20600 (N_20600,N_18110,N_17904);
nand U20601 (N_20601,N_18881,N_18116);
nor U20602 (N_20602,N_19335,N_18289);
and U20603 (N_20603,N_19470,N_19832);
nor U20604 (N_20604,N_19467,N_18495);
or U20605 (N_20605,N_19936,N_18148);
xnor U20606 (N_20606,N_17696,N_17806);
nor U20607 (N_20607,N_17903,N_19744);
or U20608 (N_20608,N_19788,N_19022);
nor U20609 (N_20609,N_18943,N_17872);
nor U20610 (N_20610,N_19961,N_19515);
xor U20611 (N_20611,N_18533,N_19067);
and U20612 (N_20612,N_19854,N_18669);
nand U20613 (N_20613,N_19331,N_18833);
or U20614 (N_20614,N_19988,N_19708);
xor U20615 (N_20615,N_19497,N_18982);
xnor U20616 (N_20616,N_19556,N_19842);
and U20617 (N_20617,N_19417,N_19774);
and U20618 (N_20618,N_19322,N_19950);
and U20619 (N_20619,N_18228,N_19573);
xnor U20620 (N_20620,N_19989,N_18132);
nor U20621 (N_20621,N_19325,N_18066);
nor U20622 (N_20622,N_19073,N_18907);
xor U20623 (N_20623,N_17707,N_17774);
nand U20624 (N_20624,N_18155,N_19206);
nand U20625 (N_20625,N_18391,N_18863);
nand U20626 (N_20626,N_19574,N_19150);
nand U20627 (N_20627,N_19822,N_18726);
or U20628 (N_20628,N_19957,N_19544);
nor U20629 (N_20629,N_17740,N_17939);
nor U20630 (N_20630,N_18390,N_18512);
nor U20631 (N_20631,N_18004,N_18403);
and U20632 (N_20632,N_18538,N_18283);
nand U20633 (N_20633,N_18701,N_18715);
nor U20634 (N_20634,N_19511,N_19211);
or U20635 (N_20635,N_17900,N_19478);
and U20636 (N_20636,N_18752,N_19725);
nor U20637 (N_20637,N_19106,N_18012);
or U20638 (N_20638,N_19358,N_18717);
xnor U20639 (N_20639,N_18790,N_19906);
xor U20640 (N_20640,N_18214,N_18368);
and U20641 (N_20641,N_18423,N_17742);
or U20642 (N_20642,N_19547,N_19845);
and U20643 (N_20643,N_17700,N_19646);
or U20644 (N_20644,N_19777,N_17563);
and U20645 (N_20645,N_18016,N_18196);
or U20646 (N_20646,N_17737,N_18623);
nand U20647 (N_20647,N_17968,N_17616);
xnor U20648 (N_20648,N_19101,N_18251);
xnor U20649 (N_20649,N_18323,N_19912);
xor U20650 (N_20650,N_19001,N_17660);
nor U20651 (N_20651,N_19741,N_19295);
or U20652 (N_20652,N_18876,N_18618);
nand U20653 (N_20653,N_18381,N_19945);
xnor U20654 (N_20654,N_18409,N_19266);
xor U20655 (N_20655,N_17750,N_19567);
or U20656 (N_20656,N_19816,N_19539);
xnor U20657 (N_20657,N_18864,N_19739);
nand U20658 (N_20658,N_17983,N_19340);
and U20659 (N_20659,N_19813,N_18789);
or U20660 (N_20660,N_18237,N_18485);
xnor U20661 (N_20661,N_19116,N_18660);
and U20662 (N_20662,N_19132,N_19718);
nor U20663 (N_20663,N_18583,N_19382);
xor U20664 (N_20664,N_18779,N_18860);
nand U20665 (N_20665,N_17732,N_18432);
and U20666 (N_20666,N_18361,N_19002);
nand U20667 (N_20667,N_19381,N_19499);
and U20668 (N_20668,N_19037,N_18480);
xnor U20669 (N_20669,N_19243,N_19345);
xnor U20670 (N_20670,N_18177,N_18506);
and U20671 (N_20671,N_19981,N_18267);
nor U20672 (N_20672,N_19444,N_18010);
or U20673 (N_20673,N_18477,N_18666);
nand U20674 (N_20674,N_18828,N_19220);
nor U20675 (N_20675,N_19987,N_18879);
xor U20676 (N_20676,N_18979,N_18230);
and U20677 (N_20677,N_18614,N_19663);
xor U20678 (N_20678,N_17782,N_18869);
nor U20679 (N_20679,N_18938,N_18728);
nor U20680 (N_20680,N_17745,N_19175);
and U20681 (N_20681,N_18468,N_19273);
xor U20682 (N_20682,N_19896,N_18924);
nand U20683 (N_20683,N_17854,N_19732);
nor U20684 (N_20684,N_19361,N_19671);
xor U20685 (N_20685,N_19634,N_19540);
nand U20686 (N_20686,N_19100,N_19446);
and U20687 (N_20687,N_18970,N_18429);
or U20688 (N_20688,N_18845,N_18465);
xnor U20689 (N_20689,N_19565,N_18264);
or U20690 (N_20690,N_19826,N_19272);
or U20691 (N_20691,N_18777,N_18933);
nand U20692 (N_20692,N_18280,N_18878);
nor U20693 (N_20693,N_19344,N_17830);
and U20694 (N_20694,N_17672,N_18431);
nand U20695 (N_20695,N_18218,N_18331);
xnor U20696 (N_20696,N_19074,N_18173);
xnor U20697 (N_20697,N_18579,N_19758);
nor U20698 (N_20698,N_17941,N_18268);
xor U20699 (N_20699,N_18846,N_19759);
xnor U20700 (N_20700,N_19976,N_19793);
or U20701 (N_20701,N_18873,N_18466);
and U20702 (N_20702,N_18374,N_19794);
and U20703 (N_20703,N_19862,N_18704);
nand U20704 (N_20704,N_18710,N_17957);
xnor U20705 (N_20705,N_18976,N_17747);
and U20706 (N_20706,N_19890,N_17849);
nand U20707 (N_20707,N_17864,N_19789);
or U20708 (N_20708,N_19076,N_17645);
nor U20709 (N_20709,N_18647,N_18858);
xnor U20710 (N_20710,N_19147,N_19528);
and U20711 (N_20711,N_19857,N_19153);
and U20712 (N_20712,N_18792,N_19731);
nor U20713 (N_20713,N_18586,N_18576);
or U20714 (N_20714,N_19259,N_19414);
nand U20715 (N_20715,N_19948,N_19682);
nor U20716 (N_20716,N_17565,N_17773);
xnor U20717 (N_20717,N_17727,N_19926);
and U20718 (N_20718,N_19940,N_19257);
nand U20719 (N_20719,N_18561,N_19003);
xnor U20720 (N_20720,N_19680,N_19438);
nor U20721 (N_20721,N_19489,N_19640);
and U20722 (N_20722,N_18235,N_18269);
nand U20723 (N_20723,N_19434,N_19837);
nand U20724 (N_20724,N_17500,N_17889);
nor U20725 (N_20725,N_18985,N_18074);
nand U20726 (N_20726,N_18935,N_17814);
and U20727 (N_20727,N_18170,N_19302);
xor U20728 (N_20728,N_17999,N_17883);
nand U20729 (N_20729,N_19348,N_18410);
nor U20730 (N_20730,N_17945,N_18772);
xor U20731 (N_20731,N_18835,N_18456);
or U20732 (N_20732,N_18181,N_17638);
and U20733 (N_20733,N_19562,N_19661);
nor U20734 (N_20734,N_18017,N_19456);
nor U20735 (N_20735,N_19545,N_18688);
nor U20736 (N_20736,N_17954,N_19599);
nor U20737 (N_20737,N_18422,N_17783);
or U20738 (N_20738,N_19596,N_17673);
or U20739 (N_20739,N_17906,N_19586);
or U20740 (N_20740,N_18371,N_18139);
or U20741 (N_20741,N_19480,N_19699);
and U20742 (N_20742,N_19938,N_19510);
or U20743 (N_20743,N_17687,N_18433);
and U20744 (N_20744,N_18031,N_17988);
nand U20745 (N_20745,N_19931,N_19162);
xnor U20746 (N_20746,N_18565,N_18558);
and U20747 (N_20747,N_17557,N_19656);
nand U20748 (N_20748,N_18310,N_17964);
and U20749 (N_20749,N_17731,N_19403);
xnor U20750 (N_20750,N_19909,N_17801);
and U20751 (N_20751,N_19338,N_18389);
nand U20752 (N_20752,N_19524,N_18077);
nand U20753 (N_20753,N_18394,N_18934);
or U20754 (N_20754,N_18467,N_18992);
nor U20755 (N_20755,N_19874,N_17982);
or U20756 (N_20756,N_19152,N_17825);
nand U20757 (N_20757,N_17690,N_19201);
or U20758 (N_20758,N_18315,N_19102);
and U20759 (N_20759,N_19534,N_18906);
nor U20760 (N_20760,N_18198,N_19748);
or U20761 (N_20761,N_18557,N_19757);
or U20762 (N_20762,N_18884,N_17948);
nor U20763 (N_20763,N_19167,N_18794);
xor U20764 (N_20764,N_17676,N_18165);
nor U20765 (N_20765,N_19285,N_18830);
and U20766 (N_20766,N_18587,N_19532);
xnor U20767 (N_20767,N_18090,N_17981);
nor U20768 (N_20768,N_18156,N_19829);
nor U20769 (N_20769,N_18627,N_18205);
xor U20770 (N_20770,N_17958,N_19745);
nor U20771 (N_20771,N_18288,N_19242);
or U20772 (N_20772,N_18900,N_19454);
xnor U20773 (N_20773,N_18780,N_18570);
and U20774 (N_20774,N_19291,N_18440);
nand U20775 (N_20775,N_18823,N_19128);
xor U20776 (N_20776,N_18226,N_19799);
or U20777 (N_20777,N_19326,N_19474);
or U20778 (N_20778,N_17704,N_19018);
xnor U20779 (N_20779,N_18606,N_18141);
or U20780 (N_20780,N_18339,N_18408);
nand U20781 (N_20781,N_19659,N_17626);
nand U20782 (N_20782,N_19643,N_19058);
and U20783 (N_20783,N_17714,N_17775);
nand U20784 (N_20784,N_19104,N_17996);
nand U20785 (N_20785,N_17842,N_17758);
xnor U20786 (N_20786,N_18544,N_18366);
xor U20787 (N_20787,N_19155,N_17835);
nor U20788 (N_20788,N_19864,N_19843);
nand U20789 (N_20789,N_18542,N_17908);
and U20790 (N_20790,N_18912,N_18295);
nor U20791 (N_20791,N_18509,N_18133);
xnor U20792 (N_20792,N_19040,N_19645);
nor U20793 (N_20793,N_19642,N_18595);
and U20794 (N_20794,N_17725,N_19865);
nand U20795 (N_20795,N_19404,N_17622);
xnor U20796 (N_20796,N_18649,N_19675);
nor U20797 (N_20797,N_18275,N_18819);
nand U20798 (N_20798,N_19050,N_19918);
or U20799 (N_20799,N_18149,N_18781);
and U20800 (N_20800,N_18775,N_18121);
or U20801 (N_20801,N_17917,N_17918);
xor U20802 (N_20802,N_19025,N_18281);
or U20803 (N_20803,N_19600,N_17863);
and U20804 (N_20804,N_19738,N_19546);
nand U20805 (N_20805,N_19724,N_19623);
or U20806 (N_20806,N_19157,N_18272);
and U20807 (N_20807,N_19558,N_18129);
nor U20808 (N_20808,N_18401,N_19455);
nor U20809 (N_20809,N_19253,N_17838);
xnor U20810 (N_20810,N_18402,N_17573);
or U20811 (N_20811,N_18585,N_18898);
xnor U20812 (N_20812,N_17572,N_19095);
nand U20813 (N_20813,N_19311,N_17950);
and U20814 (N_20814,N_19521,N_18597);
nand U20815 (N_20815,N_18634,N_18109);
xnor U20816 (N_20816,N_18242,N_18359);
or U20817 (N_20817,N_19125,N_19265);
or U20818 (N_20818,N_19161,N_19624);
xor U20819 (N_20819,N_17706,N_19000);
nor U20820 (N_20820,N_18553,N_17944);
nand U20821 (N_20821,N_18412,N_19060);
or U20822 (N_20822,N_19323,N_18184);
nand U20823 (N_20823,N_18424,N_19122);
and U20824 (N_20824,N_19089,N_17629);
nand U20825 (N_20825,N_18382,N_17813);
nor U20826 (N_20826,N_19059,N_18625);
nand U20827 (N_20827,N_19971,N_19763);
xor U20828 (N_20828,N_18417,N_17776);
and U20829 (N_20829,N_18341,N_19752);
xnor U20830 (N_20830,N_18023,N_18250);
and U20831 (N_20831,N_19418,N_18990);
xor U20832 (N_20832,N_19871,N_17615);
and U20833 (N_20833,N_19413,N_18411);
or U20834 (N_20834,N_17867,N_18811);
nand U20835 (N_20835,N_19761,N_17599);
nor U20836 (N_20836,N_17685,N_18785);
nand U20837 (N_20837,N_19451,N_18872);
xor U20838 (N_20838,N_18050,N_17784);
and U20839 (N_20839,N_19442,N_19613);
xor U20840 (N_20840,N_18009,N_18584);
nor U20841 (N_20841,N_17670,N_19548);
nor U20842 (N_20842,N_18653,N_17992);
nand U20843 (N_20843,N_19920,N_18105);
xor U20844 (N_20844,N_18999,N_18188);
nand U20845 (N_20845,N_17859,N_17600);
and U20846 (N_20846,N_19020,N_18892);
nand U20847 (N_20847,N_19065,N_19953);
nand U20848 (N_20848,N_17777,N_19109);
xor U20849 (N_20849,N_17652,N_17874);
nand U20850 (N_20850,N_17956,N_18857);
nand U20851 (N_20851,N_18470,N_17910);
nand U20852 (N_20852,N_18971,N_18425);
nand U20853 (N_20853,N_18975,N_18682);
xnor U20854 (N_20854,N_19815,N_19753);
nor U20855 (N_20855,N_18761,N_19179);
or U20856 (N_20856,N_19512,N_17882);
or U20857 (N_20857,N_19298,N_19286);
nand U20858 (N_20858,N_17569,N_19886);
or U20859 (N_20859,N_17860,N_18760);
nor U20860 (N_20860,N_19764,N_17516);
nor U20861 (N_20861,N_17902,N_19828);
xnor U20862 (N_20862,N_17760,N_18643);
and U20863 (N_20863,N_17585,N_19990);
or U20864 (N_20864,N_17937,N_18344);
nor U20865 (N_20865,N_19435,N_18065);
and U20866 (N_20866,N_17717,N_17922);
xor U20867 (N_20867,N_18082,N_18650);
and U20868 (N_20868,N_17668,N_18636);
and U20869 (N_20869,N_19394,N_19250);
xor U20870 (N_20870,N_18333,N_17836);
xnor U20871 (N_20871,N_17819,N_19280);
nor U20872 (N_20872,N_18514,N_19142);
xnor U20873 (N_20873,N_19955,N_18712);
xnor U20874 (N_20874,N_19619,N_19787);
or U20875 (N_20875,N_17986,N_19294);
nand U20876 (N_20876,N_18981,N_19318);
or U20877 (N_20877,N_17594,N_19860);
and U20878 (N_20878,N_17897,N_17562);
nand U20879 (N_20879,N_19160,N_19519);
and U20880 (N_20880,N_19723,N_18186);
xor U20881 (N_20881,N_17665,N_18472);
nand U20882 (N_20882,N_17786,N_18384);
nand U20883 (N_20883,N_17931,N_17993);
nand U20884 (N_20884,N_18112,N_18163);
nand U20885 (N_20885,N_19187,N_18806);
and U20886 (N_20886,N_19504,N_18202);
or U20887 (N_20887,N_19055,N_19587);
nor U20888 (N_20888,N_19870,N_19509);
nand U20889 (N_20889,N_19198,N_19876);
or U20890 (N_20890,N_18037,N_17851);
or U20891 (N_20891,N_17712,N_17618);
nor U20892 (N_20892,N_17730,N_18365);
and U20893 (N_20893,N_19610,N_18070);
nand U20894 (N_20894,N_17564,N_18711);
or U20895 (N_20895,N_17928,N_18276);
nand U20896 (N_20896,N_18164,N_19612);
or U20897 (N_20897,N_17627,N_17985);
xnor U20898 (N_20898,N_18727,N_19136);
or U20899 (N_20899,N_17513,N_17521);
nand U20900 (N_20900,N_19416,N_18617);
or U20901 (N_20901,N_18028,N_18952);
nor U20902 (N_20902,N_17905,N_18499);
and U20903 (N_20903,N_18386,N_18054);
or U20904 (N_20904,N_18635,N_19290);
nor U20905 (N_20905,N_18463,N_18774);
nand U20906 (N_20906,N_19393,N_19692);
and U20907 (N_20907,N_19494,N_18034);
xor U20908 (N_20908,N_19191,N_19042);
nor U20909 (N_20909,N_17967,N_19653);
or U20910 (N_20910,N_18670,N_18178);
and U20911 (N_20911,N_19765,N_19029);
xnor U20912 (N_20912,N_17602,N_19973);
nand U20913 (N_20913,N_19933,N_18294);
nor U20914 (N_20914,N_19858,N_18812);
and U20915 (N_20915,N_19164,N_17649);
and U20916 (N_20916,N_19925,N_17768);
or U20917 (N_20917,N_18405,N_18125);
and U20918 (N_20918,N_17567,N_17716);
nand U20919 (N_20919,N_18615,N_18697);
and U20920 (N_20920,N_17574,N_17744);
nand U20921 (N_20921,N_19466,N_19713);
nand U20922 (N_20922,N_17509,N_18094);
nor U20923 (N_20923,N_19235,N_18947);
xnor U20924 (N_20924,N_18763,N_18454);
nand U20925 (N_20925,N_18994,N_19743);
nor U20926 (N_20926,N_18831,N_17837);
or U20927 (N_20927,N_19715,N_17542);
and U20928 (N_20928,N_18685,N_19127);
or U20929 (N_20929,N_19450,N_18435);
and U20930 (N_20930,N_19677,N_18182);
nor U20931 (N_20931,N_18548,N_18222);
nand U20932 (N_20932,N_19975,N_18441);
xnor U20933 (N_20933,N_19426,N_19893);
or U20934 (N_20934,N_19848,N_19399);
nand U20935 (N_20935,N_19370,N_18053);
and U20936 (N_20936,N_18904,N_19195);
xnor U20937 (N_20937,N_19726,N_19684);
and U20938 (N_20938,N_19423,N_19043);
xnor U20939 (N_20939,N_19982,N_18946);
nor U20940 (N_20940,N_18720,N_18652);
nand U20941 (N_20941,N_19075,N_18968);
and U20942 (N_20942,N_18655,N_19575);
xnor U20943 (N_20943,N_17614,N_19365);
nand U20944 (N_20944,N_18135,N_19207);
nor U20945 (N_20945,N_19172,N_17679);
nor U20946 (N_20946,N_19768,N_19296);
nand U20947 (N_20947,N_19673,N_18746);
nor U20948 (N_20948,N_17887,N_19071);
or U20949 (N_20949,N_18000,N_18209);
and U20950 (N_20950,N_18364,N_18142);
nand U20951 (N_20951,N_18455,N_18928);
or U20952 (N_20952,N_17853,N_18215);
xor U20953 (N_20953,N_19410,N_17911);
nand U20954 (N_20954,N_18799,N_17514);
or U20955 (N_20955,N_17898,N_19321);
and U20956 (N_20956,N_19498,N_18334);
xor U20957 (N_20957,N_19482,N_19307);
xnor U20958 (N_20958,N_19373,N_19666);
or U20959 (N_20959,N_18097,N_17502);
and U20960 (N_20960,N_18755,N_17689);
nand U20961 (N_20961,N_18377,N_18678);
or U20962 (N_20962,N_18822,N_19391);
nor U20963 (N_20963,N_18882,N_18836);
nor U20964 (N_20964,N_17824,N_19651);
xnor U20965 (N_20965,N_18413,N_19476);
and U20966 (N_20966,N_19231,N_18951);
and U20967 (N_20967,N_18231,N_18033);
or U20968 (N_20968,N_19210,N_18086);
or U20969 (N_20969,N_17924,N_19603);
nor U20970 (N_20970,N_19523,N_17709);
xor U20971 (N_20971,N_18844,N_19655);
nor U20972 (N_20972,N_18886,N_19561);
xnor U20973 (N_20973,N_19115,N_19583);
nand U20974 (N_20974,N_18208,N_18800);
or U20975 (N_20975,N_17952,N_18079);
nand U20976 (N_20976,N_17805,N_18894);
or U20977 (N_20977,N_18608,N_17792);
and U20978 (N_20978,N_18778,N_18771);
and U20979 (N_20979,N_17756,N_18893);
and U20980 (N_20980,N_18118,N_18880);
xor U20981 (N_20981,N_17681,N_18664);
and U20982 (N_20982,N_17590,N_18494);
and U20983 (N_20983,N_19984,N_17896);
or U20984 (N_20984,N_19363,N_19151);
or U20985 (N_20985,N_18051,N_19495);
or U20986 (N_20986,N_19487,N_19650);
nor U20987 (N_20987,N_18076,N_17506);
and U20988 (N_20988,N_18154,N_18219);
nor U20989 (N_20989,N_19853,N_18484);
xor U20990 (N_20990,N_18375,N_19378);
and U20991 (N_20991,N_19047,N_19421);
xor U20992 (N_20992,N_18406,N_19019);
xnor U20993 (N_20993,N_18925,N_18285);
and U20994 (N_20994,N_19959,N_18630);
or U20995 (N_20995,N_18568,N_18233);
nand U20996 (N_20996,N_18058,N_18535);
nor U20997 (N_20997,N_18966,N_17702);
xor U20998 (N_20998,N_18605,N_18335);
or U20999 (N_20999,N_17662,N_18663);
nand U21000 (N_21000,N_19457,N_19897);
nor U21001 (N_21001,N_18867,N_19200);
nand U21002 (N_21002,N_17507,N_17858);
xnor U21003 (N_21003,N_18224,N_19779);
xnor U21004 (N_21004,N_18046,N_18651);
nand U21005 (N_21005,N_19339,N_19133);
nand U21006 (N_21006,N_19902,N_17998);
and U21007 (N_21007,N_18019,N_19247);
xnor U21008 (N_21008,N_19359,N_19887);
nor U21009 (N_21009,N_19130,N_18340);
xor U21010 (N_21010,N_19514,N_18278);
nand U21011 (N_21011,N_17976,N_19657);
and U21012 (N_21012,N_18559,N_18089);
or U21013 (N_21013,N_18327,N_18370);
nand U21014 (N_21014,N_18709,N_18803);
nor U21015 (N_21015,N_17621,N_19463);
and U21016 (N_21016,N_19057,N_17535);
nand U21017 (N_21017,N_18473,N_19588);
and U21018 (N_21018,N_19056,N_19163);
and U21019 (N_21019,N_18078,N_17663);
and U21020 (N_21020,N_18977,N_18372);
or U21021 (N_21021,N_18043,N_18989);
and U21022 (N_21022,N_18253,N_17664);
and U21023 (N_21023,N_17603,N_17733);
nor U21024 (N_21024,N_17695,N_17595);
and U21025 (N_21025,N_19803,N_18151);
and U21026 (N_21026,N_17581,N_19278);
xnor U21027 (N_21027,N_19604,N_18705);
nor U21028 (N_21028,N_19196,N_17994);
nor U21029 (N_21029,N_18316,N_18983);
nand U21030 (N_21030,N_17925,N_19024);
and U21031 (N_21031,N_17755,N_19486);
xor U21032 (N_21032,N_19248,N_19917);
xor U21033 (N_21033,N_17809,N_19536);
nor U21034 (N_21034,N_19979,N_18741);
xnor U21035 (N_21035,N_19831,N_19922);
and U21036 (N_21036,N_18168,N_18444);
nor U21037 (N_21037,N_19530,N_18524);
and U21038 (N_21038,N_19108,N_18770);
and U21039 (N_21039,N_19292,N_19780);
nand U21040 (N_21040,N_19013,N_17718);
and U21041 (N_21041,N_19830,N_18240);
xor U21042 (N_21042,N_17980,N_18279);
nor U21043 (N_21043,N_19631,N_19746);
nor U21044 (N_21044,N_18722,N_19428);
or U21045 (N_21045,N_18988,N_19400);
xor U21046 (N_21046,N_19411,N_17655);
nor U21047 (N_21047,N_17545,N_18287);
nand U21048 (N_21048,N_19317,N_17609);
and U21049 (N_21049,N_17583,N_19972);
or U21050 (N_21050,N_19840,N_19433);
nand U21051 (N_21051,N_17915,N_17916);
nand U21052 (N_21052,N_18733,N_19595);
or U21053 (N_21053,N_18998,N_17538);
or U21054 (N_21054,N_17554,N_19535);
and U21055 (N_21055,N_18213,N_18612);
nor U21056 (N_21056,N_18949,N_18229);
and U21057 (N_21057,N_19760,N_18578);
nand U21058 (N_21058,N_19796,N_18393);
xor U21059 (N_21059,N_17586,N_18903);
nor U21060 (N_21060,N_18286,N_18861);
xor U21061 (N_21061,N_18684,N_17748);
nand U21062 (N_21062,N_18143,N_18566);
and U21063 (N_21063,N_18481,N_18564);
xnor U21064 (N_21064,N_19392,N_18768);
and U21065 (N_21065,N_19637,N_19776);
and U21066 (N_21066,N_18766,N_17946);
nand U21067 (N_21067,N_19493,N_17876);
xor U21068 (N_21068,N_18014,N_18732);
or U21069 (N_21069,N_18212,N_19081);
xor U21070 (N_21070,N_18769,N_19453);
or U21071 (N_21071,N_19835,N_18072);
and U21072 (N_21072,N_18511,N_17877);
nor U21073 (N_21073,N_18930,N_19436);
nand U21074 (N_21074,N_19992,N_19811);
and U21075 (N_21075,N_18848,N_19720);
and U21076 (N_21076,N_19289,N_18126);
and U21077 (N_21077,N_18362,N_17523);
and U21078 (N_21078,N_18190,N_19390);
or U21079 (N_21079,N_18662,N_18042);
and U21080 (N_21080,N_18602,N_18490);
or U21081 (N_21081,N_18648,N_18948);
nor U21082 (N_21082,N_19123,N_18668);
xor U21083 (N_21083,N_18696,N_18624);
xor U21084 (N_21084,N_19968,N_18238);
or U21085 (N_21085,N_18832,N_19697);
or U21086 (N_21086,N_17962,N_19087);
or U21087 (N_21087,N_18742,N_18321);
xnor U21088 (N_21088,N_19784,N_18730);
or U21089 (N_21089,N_17524,N_18313);
or U21090 (N_21090,N_18293,N_18400);
nor U21091 (N_21091,N_17503,N_17781);
xor U21092 (N_21092,N_17592,N_17546);
and U21093 (N_21093,N_18388,N_19629);
nor U21094 (N_21094,N_19299,N_17912);
or U21095 (N_21095,N_18445,N_17591);
nand U21096 (N_21096,N_19674,N_19260);
nand U21097 (N_21097,N_17667,N_19872);
nand U21098 (N_21098,N_17593,N_19963);
nand U21099 (N_21099,N_17699,N_19500);
nand U21100 (N_21100,N_17550,N_19693);
xor U21101 (N_21101,N_17683,N_18501);
or U21102 (N_21102,N_19704,N_19485);
and U21103 (N_21103,N_18582,N_17827);
nor U21104 (N_21104,N_19143,N_19014);
nand U21105 (N_21105,N_19965,N_19889);
nand U21106 (N_21106,N_17802,N_19312);
xnor U21107 (N_21107,N_17880,N_18299);
xor U21108 (N_21108,N_18369,N_18745);
and U21109 (N_21109,N_19814,N_19178);
nor U21110 (N_21110,N_19812,N_17850);
or U21111 (N_21111,N_17940,N_17881);
nand U21112 (N_21112,N_18036,N_18908);
nor U21113 (N_21113,N_18227,N_17943);
or U21114 (N_21114,N_19868,N_19159);
nor U21115 (N_21115,N_18646,N_17530);
nand U21116 (N_21116,N_18291,N_18309);
nor U21117 (N_21117,N_19701,N_19347);
or U21118 (N_21118,N_17579,N_19449);
or U21119 (N_21119,N_17650,N_18821);
xnor U21120 (N_21120,N_18609,N_18416);
and U21121 (N_21121,N_19305,N_18686);
nand U21122 (N_21122,N_19490,N_17713);
nand U21123 (N_21123,N_19703,N_18776);
or U21124 (N_21124,N_19977,N_19197);
xor U21125 (N_21125,N_19960,N_19706);
nand U21126 (N_21126,N_18428,N_18978);
nand U21127 (N_21127,N_18616,N_18842);
xor U21128 (N_21128,N_18796,N_19398);
nor U21129 (N_21129,N_18415,N_19185);
and U21130 (N_21130,N_19270,N_18825);
or U21131 (N_21131,N_19015,N_17519);
xor U21132 (N_21132,N_18460,N_18719);
nor U21133 (N_21133,N_19377,N_18883);
or U21134 (N_21134,N_18115,N_18469);
and U21135 (N_21135,N_19314,N_17674);
xor U21136 (N_21136,N_18300,N_17901);
xnor U21137 (N_21137,N_18436,N_17865);
or U21138 (N_21138,N_17596,N_19448);
or U21139 (N_21139,N_18913,N_19991);
and U21140 (N_21140,N_17828,N_19930);
xor U21141 (N_21141,N_17541,N_19584);
nor U21142 (N_21142,N_17694,N_18045);
nor U21143 (N_21143,N_19213,N_19541);
nand U21144 (N_21144,N_19027,N_19031);
and U21145 (N_21145,N_17762,N_19825);
or U21146 (N_21146,N_19303,N_18236);
and U21147 (N_21147,N_18459,N_18059);
nand U21148 (N_21148,N_17698,N_19633);
and U21149 (N_21149,N_18734,N_17654);
nand U21150 (N_21150,N_19888,N_19369);
or U21151 (N_21151,N_19542,N_18877);
and U21152 (N_21152,N_17641,N_18581);
nand U21153 (N_21153,N_19966,N_17866);
or U21154 (N_21154,N_18870,N_18008);
nor U21155 (N_21155,N_17757,N_17715);
nor U21156 (N_21156,N_18814,N_18784);
nor U21157 (N_21157,N_19425,N_18744);
and U21158 (N_21158,N_19569,N_19910);
and U21159 (N_21159,N_18706,N_19775);
or U21160 (N_21160,N_18277,N_19293);
nor U21161 (N_21161,N_18261,N_17691);
or U21162 (N_21162,N_18743,N_19085);
and U21163 (N_21163,N_19641,N_17555);
or U21164 (N_21164,N_17840,N_18713);
or U21165 (N_21165,N_19685,N_18847);
xnor U21166 (N_21166,N_18731,N_18793);
and U21167 (N_21167,N_19062,N_17606);
nor U21168 (N_21168,N_19362,N_18875);
or U21169 (N_21169,N_19300,N_18404);
nor U21170 (N_21170,N_19863,N_19254);
nor U21171 (N_21171,N_19174,N_19736);
or U21172 (N_21172,N_18478,N_19407);
and U21173 (N_21173,N_19429,N_19856);
nor U21174 (N_21174,N_17642,N_18349);
nand U21175 (N_21175,N_17847,N_19994);
nor U21176 (N_21176,N_18471,N_18446);
nor U21177 (N_21177,N_17584,N_18699);
nand U21178 (N_21178,N_19328,N_17559);
nand U21179 (N_21179,N_19137,N_18885);
nor U21180 (N_21180,N_18827,N_18342);
nand U21181 (N_21181,N_17520,N_18551);
xor U21182 (N_21182,N_19097,N_18134);
and U21183 (N_21183,N_19891,N_19712);
and U21184 (N_21184,N_19460,N_19281);
nor U21185 (N_21185,N_17885,N_17855);
and U21186 (N_21186,N_19533,N_19349);
or U21187 (N_21187,N_18355,N_18693);
nand U21188 (N_21188,N_19107,N_18095);
nand U21189 (N_21189,N_19951,N_18554);
or U21190 (N_21190,N_17754,N_17724);
and U21191 (N_21191,N_18687,N_19120);
nand U21192 (N_21192,N_19672,N_19408);
xor U21193 (N_21193,N_18534,N_17739);
xor U21194 (N_21194,N_19284,N_19747);
xnor U21195 (N_21195,N_19134,N_19941);
or U21196 (N_21196,N_17772,N_19928);
or U21197 (N_21197,N_19222,N_17978);
nor U21198 (N_21198,N_19606,N_19297);
or U21199 (N_21199,N_19602,N_19063);
nor U21200 (N_21200,N_19807,N_17894);
xor U21201 (N_21201,N_17862,N_19350);
nor U21202 (N_21202,N_17846,N_18175);
and U21203 (N_21203,N_18810,N_19277);
xor U21204 (N_21204,N_18671,N_18035);
or U21205 (N_21205,N_19833,N_17927);
or U21206 (N_21206,N_18747,N_19332);
nor U21207 (N_21207,N_19721,N_18111);
xnor U21208 (N_21208,N_19644,N_19525);
xnor U21209 (N_21209,N_17643,N_18378);
nand U21210 (N_21210,N_18056,N_19552);
xnor U21211 (N_21211,N_19353,N_18169);
or U21212 (N_21212,N_17536,N_18681);
or U21213 (N_21213,N_18991,N_17820);
xor U21214 (N_21214,N_18447,N_19372);
xnor U21215 (N_21215,N_18820,N_18536);
nand U21216 (N_21216,N_19244,N_18824);
and U21217 (N_21217,N_18068,N_17628);
and U21218 (N_21218,N_18395,N_18590);
xor U21219 (N_21219,N_18140,N_19695);
or U21220 (N_21220,N_17793,N_18927);
nand U21221 (N_21221,N_19628,N_19880);
and U21222 (N_21222,N_19618,N_18718);
and U21223 (N_21223,N_18560,N_18839);
nand U21224 (N_21224,N_19996,N_17532);
and U21225 (N_21225,N_17834,N_19368);
xnor U21226 (N_21226,N_19342,N_18387);
or U21227 (N_21227,N_19967,N_18071);
nor U21228 (N_21228,N_19898,N_18737);
nand U21229 (N_21229,N_17508,N_18107);
and U21230 (N_21230,N_18896,N_18305);
and U21231 (N_21231,N_18767,N_19954);
and U21232 (N_21232,N_17610,N_19306);
xor U21233 (N_21233,N_18969,N_18546);
and U21234 (N_21234,N_19627,N_19800);
or U21235 (N_21235,N_18520,N_18598);
or U21236 (N_21236,N_19245,N_19261);
or U21237 (N_21237,N_19516,N_19088);
nand U21238 (N_21238,N_18543,N_17884);
and U21239 (N_21239,N_18532,N_18865);
or U21240 (N_21240,N_19615,N_18252);
nand U21241 (N_21241,N_18358,N_19771);
nor U21242 (N_21242,N_19226,N_17729);
nor U21243 (N_21243,N_17701,N_18505);
or U21244 (N_21244,N_18123,N_18890);
or U21245 (N_21245,N_19409,N_19560);
or U21246 (N_21246,N_19234,N_18296);
nor U21247 (N_21247,N_18626,N_18621);
or U21248 (N_21248,N_17767,N_17620);
nor U21249 (N_21249,N_19202,N_18449);
or U21250 (N_21250,N_17507,N_19037);
xnor U21251 (N_21251,N_17825,N_18072);
nor U21252 (N_21252,N_18076,N_18002);
or U21253 (N_21253,N_17643,N_17544);
xnor U21254 (N_21254,N_19019,N_17681);
nor U21255 (N_21255,N_19131,N_18258);
and U21256 (N_21256,N_18593,N_19760);
xnor U21257 (N_21257,N_19282,N_17546);
nor U21258 (N_21258,N_19103,N_17528);
xor U21259 (N_21259,N_19958,N_19705);
or U21260 (N_21260,N_19266,N_19661);
and U21261 (N_21261,N_19192,N_18746);
and U21262 (N_21262,N_17765,N_17725);
or U21263 (N_21263,N_19203,N_19226);
nor U21264 (N_21264,N_18238,N_18958);
nor U21265 (N_21265,N_19647,N_18098);
or U21266 (N_21266,N_19961,N_19549);
nor U21267 (N_21267,N_18405,N_19266);
or U21268 (N_21268,N_17697,N_17844);
xnor U21269 (N_21269,N_18660,N_18397);
or U21270 (N_21270,N_17665,N_19174);
and U21271 (N_21271,N_19063,N_18073);
nor U21272 (N_21272,N_17986,N_19902);
and U21273 (N_21273,N_19659,N_17583);
or U21274 (N_21274,N_19525,N_19679);
xor U21275 (N_21275,N_19563,N_19899);
or U21276 (N_21276,N_19160,N_19315);
xor U21277 (N_21277,N_17710,N_19905);
xor U21278 (N_21278,N_19139,N_18280);
xnor U21279 (N_21279,N_18357,N_19769);
nand U21280 (N_21280,N_19163,N_17823);
or U21281 (N_21281,N_18588,N_18086);
xnor U21282 (N_21282,N_19200,N_17880);
or U21283 (N_21283,N_17835,N_19420);
nor U21284 (N_21284,N_19015,N_17560);
xnor U21285 (N_21285,N_19817,N_19602);
xnor U21286 (N_21286,N_18105,N_18638);
or U21287 (N_21287,N_19380,N_18931);
and U21288 (N_21288,N_18783,N_18756);
xor U21289 (N_21289,N_19480,N_17705);
nand U21290 (N_21290,N_18998,N_18130);
nor U21291 (N_21291,N_19041,N_18246);
and U21292 (N_21292,N_19094,N_19365);
and U21293 (N_21293,N_18870,N_19915);
or U21294 (N_21294,N_18573,N_19245);
or U21295 (N_21295,N_18606,N_19630);
xor U21296 (N_21296,N_18730,N_18244);
nand U21297 (N_21297,N_18915,N_19914);
or U21298 (N_21298,N_19366,N_19083);
or U21299 (N_21299,N_19341,N_18035);
nand U21300 (N_21300,N_17953,N_19697);
xor U21301 (N_21301,N_19660,N_19383);
xor U21302 (N_21302,N_17782,N_17988);
nor U21303 (N_21303,N_18330,N_19704);
or U21304 (N_21304,N_18114,N_18486);
or U21305 (N_21305,N_18515,N_17826);
or U21306 (N_21306,N_18622,N_17645);
nand U21307 (N_21307,N_19449,N_18105);
nor U21308 (N_21308,N_18294,N_19315);
and U21309 (N_21309,N_18050,N_18178);
or U21310 (N_21310,N_19697,N_17712);
nor U21311 (N_21311,N_17735,N_19402);
xor U21312 (N_21312,N_17519,N_18418);
or U21313 (N_21313,N_17639,N_18947);
or U21314 (N_21314,N_17525,N_17716);
nor U21315 (N_21315,N_19407,N_19604);
or U21316 (N_21316,N_19699,N_17711);
nand U21317 (N_21317,N_17681,N_18875);
nor U21318 (N_21318,N_17827,N_18888);
nand U21319 (N_21319,N_19709,N_17662);
and U21320 (N_21320,N_19454,N_17568);
nor U21321 (N_21321,N_19625,N_19308);
and U21322 (N_21322,N_17542,N_18610);
or U21323 (N_21323,N_19551,N_19465);
nand U21324 (N_21324,N_17559,N_17753);
and U21325 (N_21325,N_19387,N_19504);
or U21326 (N_21326,N_19411,N_18659);
xor U21327 (N_21327,N_19254,N_18411);
nand U21328 (N_21328,N_17706,N_19060);
and U21329 (N_21329,N_17811,N_19887);
and U21330 (N_21330,N_19895,N_18021);
nor U21331 (N_21331,N_17525,N_19335);
or U21332 (N_21332,N_19307,N_17829);
and U21333 (N_21333,N_18373,N_18193);
or U21334 (N_21334,N_19740,N_18936);
xor U21335 (N_21335,N_18494,N_18917);
xor U21336 (N_21336,N_19989,N_18260);
and U21337 (N_21337,N_18766,N_18965);
nand U21338 (N_21338,N_18181,N_17973);
nand U21339 (N_21339,N_19095,N_17744);
nor U21340 (N_21340,N_19570,N_18187);
nor U21341 (N_21341,N_18544,N_19580);
or U21342 (N_21342,N_19926,N_18299);
nor U21343 (N_21343,N_19908,N_19446);
and U21344 (N_21344,N_18334,N_18282);
xor U21345 (N_21345,N_19374,N_19286);
and U21346 (N_21346,N_19688,N_19690);
nor U21347 (N_21347,N_18556,N_17520);
xnor U21348 (N_21348,N_17771,N_17824);
and U21349 (N_21349,N_17614,N_18204);
nor U21350 (N_21350,N_18176,N_18016);
and U21351 (N_21351,N_17549,N_19381);
xor U21352 (N_21352,N_19249,N_18031);
nor U21353 (N_21353,N_19477,N_19109);
xor U21354 (N_21354,N_18294,N_18613);
and U21355 (N_21355,N_19407,N_19817);
or U21356 (N_21356,N_18185,N_19688);
or U21357 (N_21357,N_18709,N_19129);
or U21358 (N_21358,N_18949,N_17851);
nand U21359 (N_21359,N_18529,N_19964);
nand U21360 (N_21360,N_18798,N_19491);
nand U21361 (N_21361,N_19151,N_19257);
xnor U21362 (N_21362,N_18115,N_19402);
nor U21363 (N_21363,N_18043,N_18345);
nor U21364 (N_21364,N_18183,N_19199);
and U21365 (N_21365,N_18528,N_18409);
xnor U21366 (N_21366,N_19045,N_18800);
or U21367 (N_21367,N_19246,N_18273);
and U21368 (N_21368,N_18269,N_19768);
nand U21369 (N_21369,N_19372,N_19359);
nand U21370 (N_21370,N_18627,N_17935);
and U21371 (N_21371,N_18933,N_18863);
nor U21372 (N_21372,N_18047,N_18254);
nand U21373 (N_21373,N_17840,N_18074);
nand U21374 (N_21374,N_17685,N_17831);
or U21375 (N_21375,N_18917,N_19077);
or U21376 (N_21376,N_18246,N_17686);
and U21377 (N_21377,N_19752,N_18952);
xor U21378 (N_21378,N_19350,N_17919);
and U21379 (N_21379,N_18139,N_18844);
xnor U21380 (N_21380,N_18164,N_19248);
and U21381 (N_21381,N_19800,N_19547);
nand U21382 (N_21382,N_19572,N_18268);
xnor U21383 (N_21383,N_18725,N_17741);
nor U21384 (N_21384,N_19911,N_17982);
xnor U21385 (N_21385,N_18341,N_19241);
nand U21386 (N_21386,N_19826,N_18226);
nand U21387 (N_21387,N_18921,N_19107);
nor U21388 (N_21388,N_19668,N_18618);
nand U21389 (N_21389,N_19018,N_18499);
or U21390 (N_21390,N_17842,N_19183);
nor U21391 (N_21391,N_18116,N_18583);
and U21392 (N_21392,N_19567,N_19928);
nor U21393 (N_21393,N_19897,N_19252);
xor U21394 (N_21394,N_17743,N_19164);
xnor U21395 (N_21395,N_18514,N_18089);
or U21396 (N_21396,N_17966,N_18394);
or U21397 (N_21397,N_17997,N_18623);
nor U21398 (N_21398,N_17981,N_18941);
and U21399 (N_21399,N_17593,N_19259);
and U21400 (N_21400,N_18912,N_18065);
xor U21401 (N_21401,N_18518,N_17920);
nand U21402 (N_21402,N_18148,N_18564);
xnor U21403 (N_21403,N_18677,N_19560);
nor U21404 (N_21404,N_17615,N_18029);
or U21405 (N_21405,N_19157,N_17999);
nand U21406 (N_21406,N_17954,N_18372);
nor U21407 (N_21407,N_18846,N_19998);
nand U21408 (N_21408,N_17675,N_18601);
nor U21409 (N_21409,N_18582,N_17553);
or U21410 (N_21410,N_18756,N_18445);
nor U21411 (N_21411,N_19676,N_19160);
and U21412 (N_21412,N_17514,N_19371);
xnor U21413 (N_21413,N_19888,N_19331);
nand U21414 (N_21414,N_18612,N_19579);
nand U21415 (N_21415,N_18017,N_19086);
nand U21416 (N_21416,N_18230,N_19736);
nor U21417 (N_21417,N_18770,N_17983);
nor U21418 (N_21418,N_17960,N_17921);
xor U21419 (N_21419,N_17605,N_18142);
or U21420 (N_21420,N_18763,N_19712);
and U21421 (N_21421,N_19374,N_18213);
or U21422 (N_21422,N_19192,N_19823);
nand U21423 (N_21423,N_19160,N_18555);
and U21424 (N_21424,N_19016,N_19185);
or U21425 (N_21425,N_19882,N_19244);
or U21426 (N_21426,N_17549,N_18847);
nand U21427 (N_21427,N_18267,N_17905);
nor U21428 (N_21428,N_18587,N_19843);
nand U21429 (N_21429,N_19535,N_18289);
xnor U21430 (N_21430,N_18568,N_18407);
xnor U21431 (N_21431,N_18510,N_19388);
nor U21432 (N_21432,N_18258,N_19196);
nand U21433 (N_21433,N_18659,N_19497);
xor U21434 (N_21434,N_17709,N_18878);
xnor U21435 (N_21435,N_19948,N_18655);
xnor U21436 (N_21436,N_18175,N_19024);
and U21437 (N_21437,N_19687,N_19242);
and U21438 (N_21438,N_19297,N_18711);
and U21439 (N_21439,N_18576,N_18606);
xnor U21440 (N_21440,N_17689,N_18480);
xnor U21441 (N_21441,N_19144,N_17998);
nand U21442 (N_21442,N_18560,N_18334);
nor U21443 (N_21443,N_19843,N_17890);
nand U21444 (N_21444,N_18023,N_19199);
and U21445 (N_21445,N_18450,N_19397);
nor U21446 (N_21446,N_19365,N_19384);
or U21447 (N_21447,N_18313,N_19958);
nor U21448 (N_21448,N_19581,N_18424);
and U21449 (N_21449,N_18342,N_19935);
and U21450 (N_21450,N_18620,N_17793);
or U21451 (N_21451,N_17744,N_18205);
or U21452 (N_21452,N_17524,N_17798);
nor U21453 (N_21453,N_19548,N_19756);
and U21454 (N_21454,N_19790,N_18749);
xnor U21455 (N_21455,N_18817,N_18117);
nor U21456 (N_21456,N_17589,N_19059);
nand U21457 (N_21457,N_19247,N_18592);
and U21458 (N_21458,N_18101,N_19495);
nand U21459 (N_21459,N_18471,N_18637);
or U21460 (N_21460,N_19363,N_19490);
and U21461 (N_21461,N_19357,N_18821);
nand U21462 (N_21462,N_19054,N_18366);
xnor U21463 (N_21463,N_18143,N_18677);
and U21464 (N_21464,N_18650,N_19572);
nand U21465 (N_21465,N_19692,N_17881);
xor U21466 (N_21466,N_18582,N_18790);
and U21467 (N_21467,N_18113,N_18857);
nand U21468 (N_21468,N_18705,N_18946);
xnor U21469 (N_21469,N_19949,N_18522);
nand U21470 (N_21470,N_18595,N_18522);
nand U21471 (N_21471,N_19236,N_19613);
nor U21472 (N_21472,N_18615,N_19479);
xnor U21473 (N_21473,N_19345,N_19015);
xnor U21474 (N_21474,N_17850,N_17518);
or U21475 (N_21475,N_19338,N_17632);
nand U21476 (N_21476,N_18230,N_18307);
and U21477 (N_21477,N_18695,N_19508);
xor U21478 (N_21478,N_18039,N_18251);
nor U21479 (N_21479,N_18698,N_19783);
nor U21480 (N_21480,N_17510,N_18440);
nand U21481 (N_21481,N_19490,N_18100);
nor U21482 (N_21482,N_19733,N_19043);
and U21483 (N_21483,N_18961,N_18345);
and U21484 (N_21484,N_19937,N_17670);
nand U21485 (N_21485,N_18507,N_19575);
and U21486 (N_21486,N_18595,N_17848);
nor U21487 (N_21487,N_19248,N_18605);
nand U21488 (N_21488,N_17600,N_18742);
nand U21489 (N_21489,N_19963,N_17993);
and U21490 (N_21490,N_17778,N_18709);
or U21491 (N_21491,N_19512,N_18343);
and U21492 (N_21492,N_18225,N_18592);
xor U21493 (N_21493,N_17532,N_18231);
nand U21494 (N_21494,N_18921,N_18884);
or U21495 (N_21495,N_19292,N_19220);
and U21496 (N_21496,N_18094,N_17994);
and U21497 (N_21497,N_18847,N_18171);
nand U21498 (N_21498,N_19856,N_18193);
nand U21499 (N_21499,N_19649,N_17918);
or U21500 (N_21500,N_19739,N_19718);
and U21501 (N_21501,N_19790,N_18654);
or U21502 (N_21502,N_18460,N_19463);
xnor U21503 (N_21503,N_18541,N_17871);
or U21504 (N_21504,N_18723,N_18027);
nand U21505 (N_21505,N_18485,N_18280);
nand U21506 (N_21506,N_18686,N_18554);
or U21507 (N_21507,N_17937,N_19322);
xor U21508 (N_21508,N_17690,N_18673);
and U21509 (N_21509,N_18634,N_19146);
nand U21510 (N_21510,N_17793,N_18575);
nor U21511 (N_21511,N_17578,N_17737);
nor U21512 (N_21512,N_19313,N_18675);
nor U21513 (N_21513,N_18845,N_18907);
nand U21514 (N_21514,N_19136,N_18421);
and U21515 (N_21515,N_18956,N_18070);
or U21516 (N_21516,N_19407,N_19730);
nor U21517 (N_21517,N_18609,N_19502);
nand U21518 (N_21518,N_19925,N_19333);
and U21519 (N_21519,N_18511,N_17894);
xnor U21520 (N_21520,N_17570,N_17723);
nor U21521 (N_21521,N_17682,N_19534);
or U21522 (N_21522,N_18617,N_17512);
and U21523 (N_21523,N_18176,N_18615);
and U21524 (N_21524,N_17532,N_19412);
or U21525 (N_21525,N_17932,N_18696);
and U21526 (N_21526,N_18766,N_17686);
nor U21527 (N_21527,N_18786,N_17985);
nor U21528 (N_21528,N_18111,N_19811);
nor U21529 (N_21529,N_17900,N_17742);
and U21530 (N_21530,N_19154,N_18823);
or U21531 (N_21531,N_18159,N_18853);
xnor U21532 (N_21532,N_19245,N_18306);
nand U21533 (N_21533,N_18896,N_18319);
nor U21534 (N_21534,N_19505,N_19162);
and U21535 (N_21535,N_17884,N_18845);
xnor U21536 (N_21536,N_19142,N_17750);
or U21537 (N_21537,N_17897,N_18562);
nor U21538 (N_21538,N_19409,N_18118);
xor U21539 (N_21539,N_19333,N_19922);
and U21540 (N_21540,N_18868,N_19301);
nand U21541 (N_21541,N_18974,N_19559);
and U21542 (N_21542,N_19228,N_18333);
or U21543 (N_21543,N_18173,N_19440);
nor U21544 (N_21544,N_18055,N_17905);
nor U21545 (N_21545,N_18711,N_19362);
nand U21546 (N_21546,N_19679,N_19057);
or U21547 (N_21547,N_19260,N_18831);
or U21548 (N_21548,N_19506,N_19945);
nand U21549 (N_21549,N_17543,N_17976);
xnor U21550 (N_21550,N_18736,N_17926);
xor U21551 (N_21551,N_19004,N_19206);
xnor U21552 (N_21552,N_18037,N_19599);
or U21553 (N_21553,N_17939,N_18620);
and U21554 (N_21554,N_18603,N_19433);
nand U21555 (N_21555,N_18573,N_18045);
or U21556 (N_21556,N_18634,N_18087);
xor U21557 (N_21557,N_17526,N_18412);
nand U21558 (N_21558,N_18763,N_18122);
xnor U21559 (N_21559,N_17671,N_18535);
nor U21560 (N_21560,N_18867,N_19752);
and U21561 (N_21561,N_19791,N_19151);
nor U21562 (N_21562,N_17660,N_18277);
nand U21563 (N_21563,N_17526,N_18606);
nor U21564 (N_21564,N_19069,N_18133);
nor U21565 (N_21565,N_17519,N_18737);
nor U21566 (N_21566,N_18551,N_17990);
or U21567 (N_21567,N_19374,N_18680);
xor U21568 (N_21568,N_18114,N_19318);
nand U21569 (N_21569,N_19282,N_18611);
nand U21570 (N_21570,N_18073,N_17711);
nor U21571 (N_21571,N_18481,N_17726);
nand U21572 (N_21572,N_18309,N_19649);
nor U21573 (N_21573,N_18449,N_18728);
nor U21574 (N_21574,N_18952,N_17765);
nand U21575 (N_21575,N_19297,N_18923);
xor U21576 (N_21576,N_18323,N_17569);
nand U21577 (N_21577,N_19108,N_19856);
nor U21578 (N_21578,N_18519,N_19996);
nor U21579 (N_21579,N_19449,N_19660);
xor U21580 (N_21580,N_18220,N_19687);
and U21581 (N_21581,N_18106,N_19380);
xor U21582 (N_21582,N_18582,N_18011);
and U21583 (N_21583,N_19593,N_18114);
nand U21584 (N_21584,N_17677,N_19210);
nor U21585 (N_21585,N_18987,N_18900);
or U21586 (N_21586,N_19940,N_18790);
or U21587 (N_21587,N_18809,N_18682);
nor U21588 (N_21588,N_18917,N_19711);
and U21589 (N_21589,N_18375,N_17762);
nand U21590 (N_21590,N_18145,N_19420);
xor U21591 (N_21591,N_19592,N_19918);
or U21592 (N_21592,N_18320,N_19304);
nor U21593 (N_21593,N_19877,N_17979);
nor U21594 (N_21594,N_18528,N_19663);
xor U21595 (N_21595,N_18661,N_18433);
nand U21596 (N_21596,N_18685,N_19823);
and U21597 (N_21597,N_18533,N_18234);
nor U21598 (N_21598,N_19952,N_17883);
xor U21599 (N_21599,N_19195,N_19898);
nand U21600 (N_21600,N_19755,N_17672);
and U21601 (N_21601,N_18845,N_18755);
or U21602 (N_21602,N_18458,N_18702);
nand U21603 (N_21603,N_17737,N_17625);
nand U21604 (N_21604,N_18766,N_18277);
nor U21605 (N_21605,N_18474,N_19765);
xnor U21606 (N_21606,N_18389,N_19536);
nand U21607 (N_21607,N_18288,N_17922);
xor U21608 (N_21608,N_18342,N_17549);
xnor U21609 (N_21609,N_19641,N_19191);
nor U21610 (N_21610,N_18847,N_18053);
nand U21611 (N_21611,N_19940,N_19733);
or U21612 (N_21612,N_17510,N_18057);
nor U21613 (N_21613,N_18933,N_19262);
or U21614 (N_21614,N_19860,N_17798);
and U21615 (N_21615,N_18424,N_17921);
xor U21616 (N_21616,N_18125,N_19256);
nor U21617 (N_21617,N_19248,N_18442);
xor U21618 (N_21618,N_18361,N_19850);
and U21619 (N_21619,N_19698,N_19891);
or U21620 (N_21620,N_18209,N_18391);
nor U21621 (N_21621,N_18754,N_17652);
xor U21622 (N_21622,N_18403,N_17937);
nor U21623 (N_21623,N_19916,N_17737);
nor U21624 (N_21624,N_18618,N_18333);
and U21625 (N_21625,N_17744,N_18344);
and U21626 (N_21626,N_19813,N_19867);
nor U21627 (N_21627,N_19114,N_17977);
xnor U21628 (N_21628,N_19608,N_19366);
nand U21629 (N_21629,N_19219,N_19867);
nand U21630 (N_21630,N_17810,N_18785);
nor U21631 (N_21631,N_17906,N_18828);
and U21632 (N_21632,N_19978,N_17931);
or U21633 (N_21633,N_18270,N_19675);
or U21634 (N_21634,N_19918,N_18937);
xnor U21635 (N_21635,N_18486,N_17933);
or U21636 (N_21636,N_18100,N_19916);
xor U21637 (N_21637,N_18072,N_17770);
nand U21638 (N_21638,N_18392,N_18644);
nor U21639 (N_21639,N_18180,N_17632);
or U21640 (N_21640,N_19590,N_19314);
nand U21641 (N_21641,N_18017,N_17812);
and U21642 (N_21642,N_17569,N_18247);
nand U21643 (N_21643,N_19357,N_18405);
nand U21644 (N_21644,N_17575,N_18969);
nor U21645 (N_21645,N_18456,N_18959);
or U21646 (N_21646,N_18762,N_18770);
and U21647 (N_21647,N_17924,N_18373);
nand U21648 (N_21648,N_19929,N_19562);
or U21649 (N_21649,N_17909,N_18862);
xor U21650 (N_21650,N_18328,N_19963);
and U21651 (N_21651,N_18850,N_19141);
or U21652 (N_21652,N_19824,N_19641);
and U21653 (N_21653,N_18289,N_17990);
or U21654 (N_21654,N_18187,N_18720);
or U21655 (N_21655,N_18337,N_19129);
xnor U21656 (N_21656,N_19915,N_19199);
and U21657 (N_21657,N_19583,N_18301);
nor U21658 (N_21658,N_19399,N_17645);
and U21659 (N_21659,N_17583,N_19579);
and U21660 (N_21660,N_19172,N_18305);
or U21661 (N_21661,N_17964,N_18872);
nor U21662 (N_21662,N_18504,N_19781);
xnor U21663 (N_21663,N_18066,N_19698);
nor U21664 (N_21664,N_18054,N_19340);
and U21665 (N_21665,N_19940,N_17637);
and U21666 (N_21666,N_17864,N_19204);
and U21667 (N_21667,N_19550,N_19415);
and U21668 (N_21668,N_18784,N_18551);
and U21669 (N_21669,N_19745,N_17962);
and U21670 (N_21670,N_17737,N_19321);
or U21671 (N_21671,N_18916,N_19336);
xnor U21672 (N_21672,N_17793,N_18829);
nand U21673 (N_21673,N_17686,N_18564);
nor U21674 (N_21674,N_19822,N_18312);
nand U21675 (N_21675,N_19620,N_17996);
nand U21676 (N_21676,N_17769,N_19750);
and U21677 (N_21677,N_19201,N_19219);
nor U21678 (N_21678,N_18090,N_19765);
xnor U21679 (N_21679,N_19548,N_19393);
or U21680 (N_21680,N_18915,N_17803);
and U21681 (N_21681,N_18283,N_17829);
and U21682 (N_21682,N_18873,N_17991);
xor U21683 (N_21683,N_17971,N_19160);
xor U21684 (N_21684,N_17942,N_18314);
xnor U21685 (N_21685,N_18264,N_17970);
and U21686 (N_21686,N_17909,N_18829);
or U21687 (N_21687,N_18032,N_19464);
or U21688 (N_21688,N_18826,N_19602);
xor U21689 (N_21689,N_19103,N_19970);
and U21690 (N_21690,N_18015,N_18888);
xor U21691 (N_21691,N_18055,N_19738);
nor U21692 (N_21692,N_18368,N_19681);
or U21693 (N_21693,N_18664,N_18563);
or U21694 (N_21694,N_19637,N_19356);
nand U21695 (N_21695,N_18614,N_18989);
or U21696 (N_21696,N_19349,N_19535);
or U21697 (N_21697,N_17757,N_19026);
nor U21698 (N_21698,N_19268,N_17513);
xnor U21699 (N_21699,N_19146,N_17984);
nor U21700 (N_21700,N_19196,N_17857);
nand U21701 (N_21701,N_18033,N_18271);
or U21702 (N_21702,N_18380,N_18085);
or U21703 (N_21703,N_19696,N_19388);
nor U21704 (N_21704,N_18372,N_18122);
and U21705 (N_21705,N_18397,N_17704);
nand U21706 (N_21706,N_18422,N_18697);
nor U21707 (N_21707,N_19148,N_18372);
nand U21708 (N_21708,N_18718,N_19919);
and U21709 (N_21709,N_18288,N_19384);
xnor U21710 (N_21710,N_19768,N_17737);
or U21711 (N_21711,N_17523,N_18371);
nor U21712 (N_21712,N_19591,N_19432);
nor U21713 (N_21713,N_18856,N_19937);
nor U21714 (N_21714,N_18726,N_18442);
and U21715 (N_21715,N_19082,N_17783);
nor U21716 (N_21716,N_19765,N_19068);
xor U21717 (N_21717,N_19090,N_19281);
xor U21718 (N_21718,N_18541,N_19764);
nand U21719 (N_21719,N_18002,N_18673);
nand U21720 (N_21720,N_19169,N_17948);
xor U21721 (N_21721,N_19293,N_19860);
nand U21722 (N_21722,N_19891,N_18232);
and U21723 (N_21723,N_18555,N_19284);
nand U21724 (N_21724,N_18285,N_18138);
nor U21725 (N_21725,N_18683,N_18183);
or U21726 (N_21726,N_18777,N_19995);
xor U21727 (N_21727,N_18226,N_19146);
or U21728 (N_21728,N_19356,N_18031);
nand U21729 (N_21729,N_18123,N_19332);
nand U21730 (N_21730,N_19984,N_18260);
xor U21731 (N_21731,N_19469,N_19635);
nor U21732 (N_21732,N_19289,N_19328);
and U21733 (N_21733,N_18580,N_17877);
and U21734 (N_21734,N_19129,N_19880);
xor U21735 (N_21735,N_19088,N_18255);
nor U21736 (N_21736,N_19396,N_19158);
nand U21737 (N_21737,N_19261,N_18672);
nand U21738 (N_21738,N_19923,N_19125);
and U21739 (N_21739,N_19457,N_17776);
or U21740 (N_21740,N_19110,N_19010);
and U21741 (N_21741,N_19656,N_19186);
and U21742 (N_21742,N_19051,N_18787);
nor U21743 (N_21743,N_19491,N_19809);
and U21744 (N_21744,N_18843,N_19936);
nor U21745 (N_21745,N_18025,N_18664);
xor U21746 (N_21746,N_18050,N_18953);
nor U21747 (N_21747,N_19213,N_17601);
xnor U21748 (N_21748,N_17680,N_18650);
nor U21749 (N_21749,N_17666,N_19052);
xor U21750 (N_21750,N_19203,N_18188);
nand U21751 (N_21751,N_18639,N_17615);
nand U21752 (N_21752,N_17545,N_18401);
nand U21753 (N_21753,N_19952,N_18041);
and U21754 (N_21754,N_18239,N_17544);
nor U21755 (N_21755,N_19406,N_19440);
or U21756 (N_21756,N_18044,N_19405);
xor U21757 (N_21757,N_18585,N_18744);
nor U21758 (N_21758,N_18635,N_17645);
nor U21759 (N_21759,N_18037,N_17875);
nor U21760 (N_21760,N_19054,N_18521);
and U21761 (N_21761,N_18142,N_18377);
xnor U21762 (N_21762,N_19055,N_19042);
and U21763 (N_21763,N_17926,N_19193);
and U21764 (N_21764,N_19303,N_18125);
or U21765 (N_21765,N_18836,N_19875);
or U21766 (N_21766,N_17641,N_18612);
and U21767 (N_21767,N_18166,N_19444);
and U21768 (N_21768,N_19565,N_19299);
or U21769 (N_21769,N_17832,N_19130);
nand U21770 (N_21770,N_18435,N_19064);
nand U21771 (N_21771,N_18413,N_19941);
or U21772 (N_21772,N_18837,N_18889);
or U21773 (N_21773,N_18138,N_17957);
or U21774 (N_21774,N_18040,N_18611);
xor U21775 (N_21775,N_17757,N_19385);
nand U21776 (N_21776,N_18035,N_19294);
nand U21777 (N_21777,N_19112,N_17998);
xnor U21778 (N_21778,N_19392,N_18533);
xor U21779 (N_21779,N_19432,N_19779);
xnor U21780 (N_21780,N_19253,N_18003);
nand U21781 (N_21781,N_17970,N_19137);
or U21782 (N_21782,N_19194,N_19176);
nor U21783 (N_21783,N_19743,N_19923);
nand U21784 (N_21784,N_19192,N_19704);
and U21785 (N_21785,N_18903,N_19247);
nand U21786 (N_21786,N_18964,N_19911);
and U21787 (N_21787,N_17950,N_19571);
nand U21788 (N_21788,N_18395,N_18183);
nand U21789 (N_21789,N_18309,N_17500);
and U21790 (N_21790,N_19966,N_19636);
and U21791 (N_21791,N_19193,N_19138);
nor U21792 (N_21792,N_19975,N_18898);
xnor U21793 (N_21793,N_18001,N_17577);
nand U21794 (N_21794,N_17916,N_18102);
nor U21795 (N_21795,N_18593,N_19087);
xor U21796 (N_21796,N_19291,N_18068);
nor U21797 (N_21797,N_19750,N_17536);
and U21798 (N_21798,N_19191,N_18842);
or U21799 (N_21799,N_18449,N_17679);
xnor U21800 (N_21800,N_17742,N_18051);
and U21801 (N_21801,N_18381,N_17777);
nand U21802 (N_21802,N_17505,N_19657);
or U21803 (N_21803,N_19560,N_19091);
or U21804 (N_21804,N_19337,N_18603);
or U21805 (N_21805,N_18952,N_18736);
xor U21806 (N_21806,N_17645,N_18191);
nand U21807 (N_21807,N_17815,N_18235);
or U21808 (N_21808,N_17694,N_18933);
xor U21809 (N_21809,N_17801,N_18118);
nand U21810 (N_21810,N_19502,N_18665);
nor U21811 (N_21811,N_17531,N_19971);
xnor U21812 (N_21812,N_17680,N_18270);
nand U21813 (N_21813,N_18281,N_19125);
and U21814 (N_21814,N_18376,N_19233);
nand U21815 (N_21815,N_17552,N_19413);
xnor U21816 (N_21816,N_19007,N_19028);
or U21817 (N_21817,N_19239,N_17649);
xor U21818 (N_21818,N_17918,N_17600);
nor U21819 (N_21819,N_17593,N_18163);
nor U21820 (N_21820,N_17770,N_18284);
xnor U21821 (N_21821,N_19907,N_19522);
nor U21822 (N_21822,N_19937,N_18894);
or U21823 (N_21823,N_18594,N_18302);
and U21824 (N_21824,N_19877,N_18846);
xnor U21825 (N_21825,N_19332,N_17737);
or U21826 (N_21826,N_18664,N_19493);
nor U21827 (N_21827,N_17773,N_18888);
or U21828 (N_21828,N_18991,N_18427);
or U21829 (N_21829,N_17783,N_17542);
nor U21830 (N_21830,N_18013,N_19213);
nor U21831 (N_21831,N_18420,N_19485);
nand U21832 (N_21832,N_19216,N_19405);
nand U21833 (N_21833,N_18888,N_18351);
nand U21834 (N_21834,N_18803,N_19808);
and U21835 (N_21835,N_19465,N_19905);
xor U21836 (N_21836,N_17712,N_19595);
or U21837 (N_21837,N_19410,N_17652);
or U21838 (N_21838,N_18060,N_19909);
and U21839 (N_21839,N_17957,N_19980);
or U21840 (N_21840,N_19782,N_19513);
nor U21841 (N_21841,N_19730,N_18512);
or U21842 (N_21842,N_17724,N_18436);
nor U21843 (N_21843,N_19297,N_17987);
nand U21844 (N_21844,N_18199,N_17689);
and U21845 (N_21845,N_19292,N_17751);
xnor U21846 (N_21846,N_19876,N_17919);
nand U21847 (N_21847,N_17673,N_17893);
nor U21848 (N_21848,N_19133,N_18397);
nor U21849 (N_21849,N_19282,N_17978);
nor U21850 (N_21850,N_17652,N_19478);
nand U21851 (N_21851,N_18220,N_18074);
nor U21852 (N_21852,N_17895,N_18795);
nor U21853 (N_21853,N_19141,N_17935);
nand U21854 (N_21854,N_18990,N_18279);
nor U21855 (N_21855,N_19323,N_18820);
xor U21856 (N_21856,N_19938,N_17517);
or U21857 (N_21857,N_18973,N_19771);
nor U21858 (N_21858,N_19612,N_19025);
or U21859 (N_21859,N_17740,N_17585);
or U21860 (N_21860,N_17857,N_18396);
and U21861 (N_21861,N_18382,N_19100);
nor U21862 (N_21862,N_19344,N_18036);
nand U21863 (N_21863,N_19126,N_19529);
nand U21864 (N_21864,N_18503,N_18358);
xor U21865 (N_21865,N_18939,N_19507);
nand U21866 (N_21866,N_19491,N_19234);
nand U21867 (N_21867,N_18905,N_18479);
and U21868 (N_21868,N_18893,N_19920);
xor U21869 (N_21869,N_19575,N_18166);
nor U21870 (N_21870,N_19268,N_18692);
nor U21871 (N_21871,N_19737,N_18636);
and U21872 (N_21872,N_19323,N_18922);
nand U21873 (N_21873,N_18672,N_19291);
nor U21874 (N_21874,N_19108,N_17931);
and U21875 (N_21875,N_17642,N_18306);
xnor U21876 (N_21876,N_17581,N_18254);
or U21877 (N_21877,N_18921,N_18664);
or U21878 (N_21878,N_17582,N_19519);
xnor U21879 (N_21879,N_19898,N_18202);
and U21880 (N_21880,N_19773,N_18218);
or U21881 (N_21881,N_19265,N_18011);
xnor U21882 (N_21882,N_17616,N_17629);
nand U21883 (N_21883,N_18453,N_19034);
nand U21884 (N_21884,N_19032,N_19321);
xor U21885 (N_21885,N_19518,N_19145);
xnor U21886 (N_21886,N_18676,N_18202);
and U21887 (N_21887,N_19199,N_18975);
or U21888 (N_21888,N_18673,N_18128);
nand U21889 (N_21889,N_18778,N_19556);
xnor U21890 (N_21890,N_19769,N_17603);
and U21891 (N_21891,N_18600,N_17596);
xnor U21892 (N_21892,N_18484,N_17751);
nor U21893 (N_21893,N_18094,N_18419);
nand U21894 (N_21894,N_18445,N_18423);
xnor U21895 (N_21895,N_17956,N_19119);
nand U21896 (N_21896,N_18509,N_19740);
or U21897 (N_21897,N_18184,N_17863);
xor U21898 (N_21898,N_18482,N_18266);
and U21899 (N_21899,N_19572,N_17830);
nor U21900 (N_21900,N_18115,N_19458);
nor U21901 (N_21901,N_18070,N_18987);
nand U21902 (N_21902,N_18403,N_18585);
nand U21903 (N_21903,N_19721,N_17608);
and U21904 (N_21904,N_18333,N_17523);
nor U21905 (N_21905,N_17677,N_19920);
or U21906 (N_21906,N_17684,N_18730);
xor U21907 (N_21907,N_19251,N_17659);
xor U21908 (N_21908,N_19869,N_19445);
or U21909 (N_21909,N_18636,N_19953);
xor U21910 (N_21910,N_19638,N_17621);
nand U21911 (N_21911,N_18831,N_17687);
xnor U21912 (N_21912,N_18722,N_18763);
nand U21913 (N_21913,N_17824,N_18509);
nor U21914 (N_21914,N_17971,N_18096);
xnor U21915 (N_21915,N_18895,N_18723);
and U21916 (N_21916,N_19880,N_18146);
and U21917 (N_21917,N_19133,N_19485);
and U21918 (N_21918,N_19578,N_18123);
nand U21919 (N_21919,N_19798,N_19633);
and U21920 (N_21920,N_18008,N_18464);
xor U21921 (N_21921,N_17755,N_18869);
nand U21922 (N_21922,N_19190,N_18612);
xnor U21923 (N_21923,N_18529,N_17816);
nor U21924 (N_21924,N_19263,N_18778);
xnor U21925 (N_21925,N_19136,N_19637);
nor U21926 (N_21926,N_17654,N_19883);
and U21927 (N_21927,N_19156,N_19449);
nand U21928 (N_21928,N_18348,N_19405);
nand U21929 (N_21929,N_19336,N_19031);
nor U21930 (N_21930,N_18908,N_18510);
xor U21931 (N_21931,N_19407,N_19749);
nor U21932 (N_21932,N_19829,N_17751);
xnor U21933 (N_21933,N_19633,N_19505);
and U21934 (N_21934,N_19319,N_18586);
nor U21935 (N_21935,N_18798,N_17967);
and U21936 (N_21936,N_17531,N_18905);
or U21937 (N_21937,N_18933,N_18017);
nor U21938 (N_21938,N_19198,N_17886);
nor U21939 (N_21939,N_19435,N_19941);
xor U21940 (N_21940,N_19578,N_19747);
xnor U21941 (N_21941,N_18359,N_18177);
or U21942 (N_21942,N_19869,N_19837);
xor U21943 (N_21943,N_17993,N_19821);
nand U21944 (N_21944,N_18496,N_19760);
and U21945 (N_21945,N_18043,N_19020);
and U21946 (N_21946,N_19940,N_19018);
nor U21947 (N_21947,N_18149,N_18640);
nor U21948 (N_21948,N_18529,N_18965);
nor U21949 (N_21949,N_17856,N_18936);
nand U21950 (N_21950,N_18830,N_18583);
xnor U21951 (N_21951,N_18790,N_19872);
nand U21952 (N_21952,N_19287,N_19266);
and U21953 (N_21953,N_19386,N_18302);
nand U21954 (N_21954,N_19552,N_19739);
xor U21955 (N_21955,N_19849,N_17797);
nand U21956 (N_21956,N_19931,N_18347);
and U21957 (N_21957,N_17611,N_17620);
or U21958 (N_21958,N_17532,N_18240);
nor U21959 (N_21959,N_19965,N_18001);
nand U21960 (N_21960,N_18423,N_19149);
nor U21961 (N_21961,N_17639,N_18891);
nand U21962 (N_21962,N_19274,N_19992);
xor U21963 (N_21963,N_18121,N_17778);
xor U21964 (N_21964,N_18459,N_18331);
nand U21965 (N_21965,N_18637,N_19043);
xnor U21966 (N_21966,N_19861,N_19820);
and U21967 (N_21967,N_18473,N_19927);
or U21968 (N_21968,N_18016,N_17877);
nor U21969 (N_21969,N_18974,N_18807);
xnor U21970 (N_21970,N_18819,N_18400);
nand U21971 (N_21971,N_18362,N_19901);
nand U21972 (N_21972,N_19636,N_19415);
and U21973 (N_21973,N_19362,N_19251);
or U21974 (N_21974,N_18485,N_19309);
and U21975 (N_21975,N_19715,N_18812);
and U21976 (N_21976,N_19699,N_18599);
nor U21977 (N_21977,N_17734,N_18420);
nand U21978 (N_21978,N_18281,N_17959);
and U21979 (N_21979,N_18567,N_19630);
nand U21980 (N_21980,N_19198,N_17924);
nor U21981 (N_21981,N_19902,N_18793);
and U21982 (N_21982,N_18681,N_19080);
nand U21983 (N_21983,N_18748,N_18270);
and U21984 (N_21984,N_17999,N_18927);
and U21985 (N_21985,N_19945,N_18836);
nor U21986 (N_21986,N_18730,N_19331);
or U21987 (N_21987,N_18048,N_19319);
or U21988 (N_21988,N_18844,N_18689);
nand U21989 (N_21989,N_18424,N_19983);
nor U21990 (N_21990,N_18513,N_17655);
nor U21991 (N_21991,N_18708,N_18796);
nor U21992 (N_21992,N_18685,N_18604);
nor U21993 (N_21993,N_18679,N_19212);
nand U21994 (N_21994,N_17633,N_18904);
and U21995 (N_21995,N_19872,N_19410);
and U21996 (N_21996,N_18216,N_19839);
nand U21997 (N_21997,N_17910,N_19803);
xnor U21998 (N_21998,N_19769,N_18221);
or U21999 (N_21999,N_19363,N_17879);
and U22000 (N_22000,N_19164,N_19585);
nand U22001 (N_22001,N_18536,N_18940);
nand U22002 (N_22002,N_17701,N_19044);
xnor U22003 (N_22003,N_18737,N_19262);
or U22004 (N_22004,N_18808,N_19554);
or U22005 (N_22005,N_19868,N_19979);
nand U22006 (N_22006,N_17906,N_18956);
nand U22007 (N_22007,N_19609,N_19345);
nand U22008 (N_22008,N_19358,N_19857);
xnor U22009 (N_22009,N_19125,N_17861);
and U22010 (N_22010,N_18007,N_18802);
xor U22011 (N_22011,N_18572,N_17619);
nor U22012 (N_22012,N_18418,N_19742);
or U22013 (N_22013,N_17960,N_18734);
and U22014 (N_22014,N_19007,N_19599);
nand U22015 (N_22015,N_18088,N_18626);
xor U22016 (N_22016,N_17976,N_18747);
and U22017 (N_22017,N_19948,N_19769);
xor U22018 (N_22018,N_19070,N_19065);
xnor U22019 (N_22019,N_19403,N_18778);
and U22020 (N_22020,N_18560,N_18804);
xnor U22021 (N_22021,N_18739,N_17677);
nor U22022 (N_22022,N_19291,N_18408);
nor U22023 (N_22023,N_17826,N_18064);
and U22024 (N_22024,N_18162,N_19032);
nand U22025 (N_22025,N_18100,N_18246);
nor U22026 (N_22026,N_19825,N_17937);
and U22027 (N_22027,N_17546,N_19537);
xor U22028 (N_22028,N_18819,N_18060);
or U22029 (N_22029,N_17680,N_19125);
xor U22030 (N_22030,N_18891,N_19062);
or U22031 (N_22031,N_19687,N_17608);
nor U22032 (N_22032,N_18399,N_17876);
or U22033 (N_22033,N_19742,N_19461);
or U22034 (N_22034,N_19522,N_17624);
or U22035 (N_22035,N_18365,N_18887);
xnor U22036 (N_22036,N_18832,N_19981);
xor U22037 (N_22037,N_18129,N_19687);
and U22038 (N_22038,N_19479,N_17782);
or U22039 (N_22039,N_19629,N_18281);
or U22040 (N_22040,N_18006,N_19242);
nor U22041 (N_22041,N_18931,N_19191);
and U22042 (N_22042,N_19860,N_19690);
and U22043 (N_22043,N_19788,N_18564);
nor U22044 (N_22044,N_18367,N_18386);
nand U22045 (N_22045,N_17782,N_18662);
or U22046 (N_22046,N_19745,N_19627);
nor U22047 (N_22047,N_19483,N_19103);
and U22048 (N_22048,N_18508,N_19159);
nand U22049 (N_22049,N_18759,N_19826);
nand U22050 (N_22050,N_19406,N_19634);
xor U22051 (N_22051,N_17571,N_19694);
xnor U22052 (N_22052,N_19489,N_17708);
xor U22053 (N_22053,N_18339,N_19352);
or U22054 (N_22054,N_18325,N_17780);
and U22055 (N_22055,N_18679,N_18136);
nand U22056 (N_22056,N_18442,N_19982);
and U22057 (N_22057,N_17947,N_19813);
xor U22058 (N_22058,N_18325,N_17824);
nor U22059 (N_22059,N_19271,N_19976);
nor U22060 (N_22060,N_19513,N_18691);
and U22061 (N_22061,N_18861,N_19764);
xor U22062 (N_22062,N_19454,N_19250);
and U22063 (N_22063,N_19620,N_18062);
nand U22064 (N_22064,N_19579,N_18506);
nor U22065 (N_22065,N_19129,N_19402);
and U22066 (N_22066,N_19991,N_17871);
nor U22067 (N_22067,N_18008,N_19663);
nor U22068 (N_22068,N_17904,N_18774);
nand U22069 (N_22069,N_19473,N_19443);
nand U22070 (N_22070,N_17606,N_18438);
or U22071 (N_22071,N_19571,N_18399);
xnor U22072 (N_22072,N_18806,N_19749);
nor U22073 (N_22073,N_19829,N_19561);
or U22074 (N_22074,N_19633,N_18740);
nor U22075 (N_22075,N_17645,N_19866);
and U22076 (N_22076,N_17926,N_18654);
nor U22077 (N_22077,N_17711,N_18461);
xor U22078 (N_22078,N_19401,N_17885);
nor U22079 (N_22079,N_18568,N_18307);
xor U22080 (N_22080,N_19606,N_18940);
nand U22081 (N_22081,N_18899,N_19093);
or U22082 (N_22082,N_18476,N_18116);
nor U22083 (N_22083,N_18612,N_18472);
nand U22084 (N_22084,N_18862,N_19087);
nand U22085 (N_22085,N_18145,N_17809);
and U22086 (N_22086,N_17606,N_19893);
nor U22087 (N_22087,N_18397,N_19820);
or U22088 (N_22088,N_19944,N_19590);
nand U22089 (N_22089,N_18573,N_18289);
nor U22090 (N_22090,N_19902,N_18896);
xor U22091 (N_22091,N_18673,N_18434);
nand U22092 (N_22092,N_19071,N_18361);
xor U22093 (N_22093,N_17915,N_18401);
xor U22094 (N_22094,N_18005,N_19914);
and U22095 (N_22095,N_19367,N_19659);
xor U22096 (N_22096,N_19244,N_19467);
nor U22097 (N_22097,N_18661,N_19178);
or U22098 (N_22098,N_18974,N_18203);
nor U22099 (N_22099,N_18852,N_19241);
nand U22100 (N_22100,N_17952,N_18690);
nand U22101 (N_22101,N_19556,N_19400);
or U22102 (N_22102,N_18582,N_17922);
and U22103 (N_22103,N_19106,N_19907);
nor U22104 (N_22104,N_17749,N_18862);
xor U22105 (N_22105,N_18262,N_17723);
and U22106 (N_22106,N_19537,N_18624);
nor U22107 (N_22107,N_18239,N_18840);
and U22108 (N_22108,N_17763,N_17573);
nor U22109 (N_22109,N_19255,N_19536);
nor U22110 (N_22110,N_19179,N_17845);
nand U22111 (N_22111,N_18014,N_17557);
xor U22112 (N_22112,N_19940,N_18121);
nand U22113 (N_22113,N_18700,N_18319);
nor U22114 (N_22114,N_18004,N_18176);
xor U22115 (N_22115,N_19940,N_18894);
xor U22116 (N_22116,N_17791,N_18093);
and U22117 (N_22117,N_17776,N_18955);
and U22118 (N_22118,N_19487,N_18586);
or U22119 (N_22119,N_18726,N_19569);
and U22120 (N_22120,N_19843,N_19780);
and U22121 (N_22121,N_17603,N_19604);
nor U22122 (N_22122,N_18685,N_18369);
xnor U22123 (N_22123,N_19948,N_19980);
nand U22124 (N_22124,N_18052,N_18692);
xor U22125 (N_22125,N_19221,N_17853);
or U22126 (N_22126,N_19183,N_18402);
nor U22127 (N_22127,N_19843,N_19890);
or U22128 (N_22128,N_18478,N_19811);
or U22129 (N_22129,N_19076,N_19996);
and U22130 (N_22130,N_18305,N_19942);
nor U22131 (N_22131,N_18512,N_17638);
nor U22132 (N_22132,N_19704,N_18481);
nand U22133 (N_22133,N_18227,N_19016);
nor U22134 (N_22134,N_18895,N_17852);
xor U22135 (N_22135,N_19775,N_18175);
nand U22136 (N_22136,N_19673,N_19720);
and U22137 (N_22137,N_18324,N_19247);
nor U22138 (N_22138,N_18649,N_18045);
and U22139 (N_22139,N_18534,N_19496);
nor U22140 (N_22140,N_19670,N_18226);
nand U22141 (N_22141,N_19619,N_18947);
and U22142 (N_22142,N_19732,N_17557);
or U22143 (N_22143,N_18040,N_17528);
or U22144 (N_22144,N_18189,N_18377);
xnor U22145 (N_22145,N_19522,N_19175);
nand U22146 (N_22146,N_18380,N_19933);
or U22147 (N_22147,N_19728,N_18261);
xnor U22148 (N_22148,N_17691,N_19845);
and U22149 (N_22149,N_18283,N_18417);
nand U22150 (N_22150,N_17799,N_18676);
or U22151 (N_22151,N_19657,N_17614);
or U22152 (N_22152,N_17752,N_17584);
xor U22153 (N_22153,N_18047,N_18060);
xnor U22154 (N_22154,N_19822,N_18617);
nor U22155 (N_22155,N_19351,N_19445);
xnor U22156 (N_22156,N_19106,N_18378);
xnor U22157 (N_22157,N_19770,N_19101);
nand U22158 (N_22158,N_18148,N_18302);
nand U22159 (N_22159,N_19863,N_19275);
nor U22160 (N_22160,N_18426,N_19712);
nand U22161 (N_22161,N_19133,N_19915);
nand U22162 (N_22162,N_17838,N_18296);
or U22163 (N_22163,N_18426,N_18811);
xnor U22164 (N_22164,N_18662,N_17857);
or U22165 (N_22165,N_19847,N_19774);
nor U22166 (N_22166,N_18531,N_18960);
nor U22167 (N_22167,N_18572,N_18175);
or U22168 (N_22168,N_18134,N_18736);
or U22169 (N_22169,N_18132,N_18553);
nor U22170 (N_22170,N_19939,N_18668);
and U22171 (N_22171,N_18254,N_18993);
nand U22172 (N_22172,N_18412,N_18485);
nand U22173 (N_22173,N_19626,N_19647);
nor U22174 (N_22174,N_18284,N_19633);
and U22175 (N_22175,N_18438,N_18682);
xnor U22176 (N_22176,N_19383,N_17892);
nor U22177 (N_22177,N_19257,N_18056);
xnor U22178 (N_22178,N_19668,N_17786);
nor U22179 (N_22179,N_19297,N_19846);
nand U22180 (N_22180,N_18524,N_18545);
nor U22181 (N_22181,N_19019,N_19464);
or U22182 (N_22182,N_18806,N_18105);
or U22183 (N_22183,N_19677,N_18691);
nor U22184 (N_22184,N_18970,N_19808);
nor U22185 (N_22185,N_18758,N_19020);
xor U22186 (N_22186,N_18897,N_18466);
or U22187 (N_22187,N_19752,N_18586);
xor U22188 (N_22188,N_17791,N_19157);
nor U22189 (N_22189,N_19638,N_19408);
nand U22190 (N_22190,N_18365,N_17935);
or U22191 (N_22191,N_18492,N_19516);
nand U22192 (N_22192,N_18754,N_19494);
and U22193 (N_22193,N_18859,N_19081);
xnor U22194 (N_22194,N_19722,N_18241);
or U22195 (N_22195,N_19573,N_18761);
nand U22196 (N_22196,N_19234,N_19416);
xnor U22197 (N_22197,N_19551,N_18428);
and U22198 (N_22198,N_18086,N_19361);
xnor U22199 (N_22199,N_19557,N_18240);
and U22200 (N_22200,N_19434,N_19548);
or U22201 (N_22201,N_18223,N_17818);
nor U22202 (N_22202,N_18891,N_18254);
nand U22203 (N_22203,N_18235,N_17853);
xor U22204 (N_22204,N_18888,N_18796);
nand U22205 (N_22205,N_18052,N_17801);
nand U22206 (N_22206,N_18279,N_19144);
xnor U22207 (N_22207,N_18134,N_18515);
and U22208 (N_22208,N_18051,N_19297);
nand U22209 (N_22209,N_17678,N_18324);
or U22210 (N_22210,N_17656,N_19332);
and U22211 (N_22211,N_18685,N_18319);
nand U22212 (N_22212,N_18078,N_18245);
nand U22213 (N_22213,N_18788,N_18679);
nor U22214 (N_22214,N_18551,N_19407);
nor U22215 (N_22215,N_19925,N_18789);
or U22216 (N_22216,N_19780,N_18587);
xnor U22217 (N_22217,N_19345,N_18098);
xnor U22218 (N_22218,N_19229,N_19211);
nand U22219 (N_22219,N_19247,N_18766);
xor U22220 (N_22220,N_17988,N_19735);
and U22221 (N_22221,N_17596,N_18866);
or U22222 (N_22222,N_18955,N_19805);
nor U22223 (N_22223,N_19009,N_19351);
and U22224 (N_22224,N_19371,N_19589);
xor U22225 (N_22225,N_18639,N_18900);
and U22226 (N_22226,N_19532,N_18314);
and U22227 (N_22227,N_18193,N_18444);
nand U22228 (N_22228,N_18907,N_18566);
nor U22229 (N_22229,N_18183,N_18250);
xor U22230 (N_22230,N_18963,N_19332);
nor U22231 (N_22231,N_19335,N_18447);
xnor U22232 (N_22232,N_17656,N_17535);
and U22233 (N_22233,N_19066,N_18255);
or U22234 (N_22234,N_18624,N_19856);
nor U22235 (N_22235,N_18557,N_19957);
and U22236 (N_22236,N_18730,N_17780);
or U22237 (N_22237,N_19209,N_17828);
xnor U22238 (N_22238,N_19904,N_17570);
and U22239 (N_22239,N_17706,N_19383);
nor U22240 (N_22240,N_19728,N_18881);
nor U22241 (N_22241,N_19553,N_19990);
nand U22242 (N_22242,N_18472,N_19320);
and U22243 (N_22243,N_17970,N_19771);
or U22244 (N_22244,N_17857,N_18671);
nor U22245 (N_22245,N_17879,N_17799);
nand U22246 (N_22246,N_18350,N_17792);
nand U22247 (N_22247,N_17782,N_19494);
nand U22248 (N_22248,N_17786,N_19600);
nor U22249 (N_22249,N_18183,N_19729);
nor U22250 (N_22250,N_17865,N_17606);
and U22251 (N_22251,N_19936,N_19493);
xnor U22252 (N_22252,N_18011,N_18302);
and U22253 (N_22253,N_18806,N_18901);
nor U22254 (N_22254,N_18520,N_17867);
or U22255 (N_22255,N_17631,N_18902);
and U22256 (N_22256,N_19665,N_19242);
nor U22257 (N_22257,N_19600,N_18158);
nor U22258 (N_22258,N_18178,N_19772);
nand U22259 (N_22259,N_19597,N_18342);
and U22260 (N_22260,N_19329,N_18317);
xnor U22261 (N_22261,N_19828,N_18666);
xor U22262 (N_22262,N_17510,N_19725);
or U22263 (N_22263,N_17899,N_19570);
nor U22264 (N_22264,N_17803,N_19872);
nor U22265 (N_22265,N_18610,N_19328);
nand U22266 (N_22266,N_19144,N_19162);
xor U22267 (N_22267,N_18895,N_17835);
nand U22268 (N_22268,N_18938,N_18126);
nand U22269 (N_22269,N_17662,N_18930);
and U22270 (N_22270,N_19330,N_18520);
xnor U22271 (N_22271,N_17773,N_17755);
and U22272 (N_22272,N_17657,N_19073);
xnor U22273 (N_22273,N_17856,N_19309);
nor U22274 (N_22274,N_17554,N_19784);
and U22275 (N_22275,N_17547,N_19389);
xnor U22276 (N_22276,N_19128,N_18595);
nand U22277 (N_22277,N_18046,N_17830);
nor U22278 (N_22278,N_18766,N_19402);
nand U22279 (N_22279,N_19149,N_17732);
nand U22280 (N_22280,N_18322,N_17860);
nand U22281 (N_22281,N_19720,N_18864);
and U22282 (N_22282,N_18891,N_18031);
nor U22283 (N_22283,N_18059,N_18321);
nor U22284 (N_22284,N_18927,N_18847);
nand U22285 (N_22285,N_18524,N_18889);
or U22286 (N_22286,N_18028,N_19251);
nand U22287 (N_22287,N_19384,N_19297);
xnor U22288 (N_22288,N_19624,N_18602);
and U22289 (N_22289,N_19283,N_19406);
nand U22290 (N_22290,N_17923,N_17836);
or U22291 (N_22291,N_17863,N_18838);
xor U22292 (N_22292,N_19694,N_18864);
nand U22293 (N_22293,N_19113,N_19342);
or U22294 (N_22294,N_19561,N_18446);
nor U22295 (N_22295,N_18317,N_18144);
nand U22296 (N_22296,N_19285,N_17543);
nand U22297 (N_22297,N_18525,N_19280);
nand U22298 (N_22298,N_19326,N_19549);
or U22299 (N_22299,N_17770,N_19654);
or U22300 (N_22300,N_18446,N_18541);
xnor U22301 (N_22301,N_17659,N_18513);
or U22302 (N_22302,N_19946,N_19755);
xor U22303 (N_22303,N_19433,N_17753);
xor U22304 (N_22304,N_17988,N_17880);
xnor U22305 (N_22305,N_18824,N_19771);
and U22306 (N_22306,N_19691,N_19500);
or U22307 (N_22307,N_19004,N_18997);
and U22308 (N_22308,N_19161,N_19869);
or U22309 (N_22309,N_19902,N_17875);
nand U22310 (N_22310,N_18727,N_18438);
or U22311 (N_22311,N_19237,N_19361);
xor U22312 (N_22312,N_17781,N_19344);
xor U22313 (N_22313,N_17519,N_18112);
and U22314 (N_22314,N_18592,N_19940);
or U22315 (N_22315,N_19468,N_17629);
nor U22316 (N_22316,N_18901,N_19268);
xnor U22317 (N_22317,N_19028,N_18198);
nand U22318 (N_22318,N_18040,N_17990);
xnor U22319 (N_22319,N_18512,N_18270);
nor U22320 (N_22320,N_18148,N_19122);
xnor U22321 (N_22321,N_17642,N_19103);
or U22322 (N_22322,N_19049,N_19408);
and U22323 (N_22323,N_17775,N_17967);
or U22324 (N_22324,N_19420,N_18163);
and U22325 (N_22325,N_17642,N_18407);
nand U22326 (N_22326,N_18163,N_18040);
nor U22327 (N_22327,N_18470,N_18048);
nand U22328 (N_22328,N_17639,N_18139);
nand U22329 (N_22329,N_18149,N_18218);
nor U22330 (N_22330,N_18392,N_18250);
xnor U22331 (N_22331,N_19259,N_19849);
nand U22332 (N_22332,N_19721,N_19198);
and U22333 (N_22333,N_17959,N_17674);
xor U22334 (N_22334,N_18017,N_18685);
nor U22335 (N_22335,N_18856,N_18929);
xor U22336 (N_22336,N_17656,N_19204);
or U22337 (N_22337,N_18705,N_17767);
nand U22338 (N_22338,N_18846,N_18260);
nor U22339 (N_22339,N_19279,N_18315);
nand U22340 (N_22340,N_18944,N_19730);
nor U22341 (N_22341,N_19359,N_18918);
xor U22342 (N_22342,N_18295,N_18337);
xor U22343 (N_22343,N_18763,N_19256);
xnor U22344 (N_22344,N_17828,N_19216);
or U22345 (N_22345,N_17855,N_18751);
or U22346 (N_22346,N_19621,N_19789);
nor U22347 (N_22347,N_19451,N_17663);
nor U22348 (N_22348,N_18311,N_18606);
nand U22349 (N_22349,N_17830,N_18348);
nor U22350 (N_22350,N_19507,N_18142);
nor U22351 (N_22351,N_18504,N_18207);
nand U22352 (N_22352,N_18076,N_17998);
and U22353 (N_22353,N_18625,N_19784);
and U22354 (N_22354,N_19108,N_18807);
or U22355 (N_22355,N_19435,N_19900);
nor U22356 (N_22356,N_18619,N_18128);
and U22357 (N_22357,N_18471,N_19884);
nor U22358 (N_22358,N_17835,N_18934);
nor U22359 (N_22359,N_19096,N_18422);
nand U22360 (N_22360,N_18816,N_18973);
nor U22361 (N_22361,N_17502,N_18891);
xnor U22362 (N_22362,N_19817,N_19941);
xnor U22363 (N_22363,N_19945,N_19987);
and U22364 (N_22364,N_19700,N_18837);
or U22365 (N_22365,N_18566,N_18911);
nor U22366 (N_22366,N_18137,N_18087);
nand U22367 (N_22367,N_19919,N_19467);
nor U22368 (N_22368,N_19423,N_17791);
or U22369 (N_22369,N_19079,N_19642);
xnor U22370 (N_22370,N_18864,N_19522);
nand U22371 (N_22371,N_18662,N_18381);
nor U22372 (N_22372,N_19140,N_18842);
xnor U22373 (N_22373,N_19607,N_19327);
nand U22374 (N_22374,N_17932,N_18015);
xor U22375 (N_22375,N_18793,N_19624);
and U22376 (N_22376,N_19094,N_19132);
nand U22377 (N_22377,N_18257,N_17647);
and U22378 (N_22378,N_18512,N_17688);
nor U22379 (N_22379,N_18870,N_19785);
xor U22380 (N_22380,N_19173,N_18725);
or U22381 (N_22381,N_19844,N_19536);
nor U22382 (N_22382,N_19475,N_18515);
nand U22383 (N_22383,N_18445,N_18499);
xnor U22384 (N_22384,N_18855,N_19934);
nor U22385 (N_22385,N_19131,N_19816);
and U22386 (N_22386,N_17917,N_19694);
nand U22387 (N_22387,N_18312,N_17764);
xnor U22388 (N_22388,N_17544,N_19863);
nor U22389 (N_22389,N_18154,N_18072);
xnor U22390 (N_22390,N_19802,N_19386);
and U22391 (N_22391,N_18036,N_18896);
xor U22392 (N_22392,N_17692,N_18455);
xnor U22393 (N_22393,N_18155,N_18225);
and U22394 (N_22394,N_17836,N_18112);
and U22395 (N_22395,N_17695,N_18743);
nor U22396 (N_22396,N_19520,N_17932);
or U22397 (N_22397,N_19499,N_19526);
xnor U22398 (N_22398,N_18493,N_19300);
and U22399 (N_22399,N_19852,N_17784);
or U22400 (N_22400,N_18927,N_18292);
nor U22401 (N_22401,N_18822,N_18009);
xnor U22402 (N_22402,N_17507,N_17908);
or U22403 (N_22403,N_17521,N_19589);
and U22404 (N_22404,N_19111,N_19099);
or U22405 (N_22405,N_19914,N_19297);
nor U22406 (N_22406,N_19007,N_19779);
or U22407 (N_22407,N_18753,N_19451);
xnor U22408 (N_22408,N_18458,N_17611);
nor U22409 (N_22409,N_18555,N_18705);
nor U22410 (N_22410,N_17809,N_17791);
nor U22411 (N_22411,N_19922,N_19895);
xnor U22412 (N_22412,N_18444,N_17794);
nor U22413 (N_22413,N_19895,N_17698);
nand U22414 (N_22414,N_19877,N_18568);
nand U22415 (N_22415,N_19567,N_19140);
or U22416 (N_22416,N_19145,N_19236);
nor U22417 (N_22417,N_19161,N_19964);
nand U22418 (N_22418,N_19389,N_19092);
nand U22419 (N_22419,N_18698,N_18018);
xnor U22420 (N_22420,N_19092,N_19539);
and U22421 (N_22421,N_18154,N_19728);
nor U22422 (N_22422,N_19417,N_19326);
nand U22423 (N_22423,N_19684,N_17692);
or U22424 (N_22424,N_19370,N_19288);
and U22425 (N_22425,N_17590,N_18465);
or U22426 (N_22426,N_18930,N_19928);
nand U22427 (N_22427,N_17664,N_19132);
or U22428 (N_22428,N_19698,N_19842);
or U22429 (N_22429,N_19384,N_18430);
or U22430 (N_22430,N_19172,N_17819);
or U22431 (N_22431,N_19457,N_18357);
nor U22432 (N_22432,N_18384,N_18546);
nor U22433 (N_22433,N_17600,N_17750);
or U22434 (N_22434,N_18084,N_18899);
nor U22435 (N_22435,N_17716,N_19885);
nor U22436 (N_22436,N_19865,N_18064);
nand U22437 (N_22437,N_18612,N_18946);
nand U22438 (N_22438,N_18629,N_18356);
or U22439 (N_22439,N_18825,N_18779);
nor U22440 (N_22440,N_19770,N_19743);
and U22441 (N_22441,N_18251,N_18500);
nor U22442 (N_22442,N_19162,N_18994);
nand U22443 (N_22443,N_17571,N_18276);
or U22444 (N_22444,N_18868,N_17728);
and U22445 (N_22445,N_18833,N_19092);
nand U22446 (N_22446,N_19632,N_18668);
or U22447 (N_22447,N_17753,N_18744);
nand U22448 (N_22448,N_18827,N_17925);
and U22449 (N_22449,N_17723,N_19544);
nor U22450 (N_22450,N_17810,N_18693);
or U22451 (N_22451,N_19399,N_18235);
or U22452 (N_22452,N_17785,N_19209);
or U22453 (N_22453,N_18887,N_17993);
and U22454 (N_22454,N_18029,N_18933);
xnor U22455 (N_22455,N_19338,N_19739);
or U22456 (N_22456,N_17932,N_19837);
and U22457 (N_22457,N_18873,N_19788);
and U22458 (N_22458,N_18872,N_18359);
and U22459 (N_22459,N_19211,N_18439);
nand U22460 (N_22460,N_19194,N_18321);
nor U22461 (N_22461,N_19676,N_18716);
xnor U22462 (N_22462,N_17628,N_19736);
and U22463 (N_22463,N_17731,N_19895);
or U22464 (N_22464,N_18412,N_18131);
nor U22465 (N_22465,N_19567,N_17844);
nand U22466 (N_22466,N_18925,N_18451);
or U22467 (N_22467,N_18697,N_17874);
or U22468 (N_22468,N_19232,N_18195);
nand U22469 (N_22469,N_19424,N_17526);
xnor U22470 (N_22470,N_19959,N_18099);
xnor U22471 (N_22471,N_18009,N_19303);
nand U22472 (N_22472,N_17522,N_18820);
or U22473 (N_22473,N_19771,N_17950);
or U22474 (N_22474,N_17745,N_19809);
xnor U22475 (N_22475,N_19908,N_19179);
nor U22476 (N_22476,N_19741,N_18788);
nand U22477 (N_22477,N_18301,N_19706);
nand U22478 (N_22478,N_18282,N_19363);
nand U22479 (N_22479,N_18981,N_19996);
or U22480 (N_22480,N_19585,N_18330);
nor U22481 (N_22481,N_19474,N_18798);
and U22482 (N_22482,N_18140,N_18190);
xor U22483 (N_22483,N_19821,N_19994);
or U22484 (N_22484,N_18234,N_18069);
nor U22485 (N_22485,N_19240,N_19459);
and U22486 (N_22486,N_19403,N_19502);
nor U22487 (N_22487,N_19785,N_18677);
nor U22488 (N_22488,N_19582,N_18552);
xor U22489 (N_22489,N_19134,N_19963);
nor U22490 (N_22490,N_19666,N_18927);
and U22491 (N_22491,N_18110,N_19705);
and U22492 (N_22492,N_18348,N_19435);
or U22493 (N_22493,N_17761,N_19332);
and U22494 (N_22494,N_17523,N_18829);
and U22495 (N_22495,N_17684,N_17826);
nor U22496 (N_22496,N_19256,N_19508);
xor U22497 (N_22497,N_19144,N_18143);
and U22498 (N_22498,N_19111,N_17950);
or U22499 (N_22499,N_18100,N_19321);
nand U22500 (N_22500,N_20422,N_22397);
nor U22501 (N_22501,N_21946,N_21655);
and U22502 (N_22502,N_21939,N_22233);
xor U22503 (N_22503,N_20269,N_20672);
xor U22504 (N_22504,N_21198,N_20618);
and U22505 (N_22505,N_21706,N_22066);
or U22506 (N_22506,N_22483,N_21312);
nand U22507 (N_22507,N_22421,N_20669);
or U22508 (N_22508,N_20121,N_21614);
and U22509 (N_22509,N_21897,N_20727);
xor U22510 (N_22510,N_20325,N_20335);
or U22511 (N_22511,N_20675,N_22193);
and U22512 (N_22512,N_20459,N_20909);
and U22513 (N_22513,N_20319,N_20446);
nor U22514 (N_22514,N_21020,N_21698);
or U22515 (N_22515,N_22032,N_21018);
or U22516 (N_22516,N_22383,N_21699);
nor U22517 (N_22517,N_21628,N_22191);
xor U22518 (N_22518,N_21039,N_20592);
nor U22519 (N_22519,N_21543,N_20509);
nand U22520 (N_22520,N_21675,N_20685);
nand U22521 (N_22521,N_20706,N_20186);
and U22522 (N_22522,N_20972,N_20808);
nor U22523 (N_22523,N_20893,N_20390);
nand U22524 (N_22524,N_20031,N_21566);
xor U22525 (N_22525,N_20845,N_21272);
nor U22526 (N_22526,N_21152,N_21284);
nand U22527 (N_22527,N_22247,N_21650);
nor U22528 (N_22528,N_22123,N_22456);
or U22529 (N_22529,N_20160,N_21777);
or U22530 (N_22530,N_22122,N_21804);
and U22531 (N_22531,N_21762,N_22455);
and U22532 (N_22532,N_21883,N_21890);
xor U22533 (N_22533,N_21214,N_20869);
nand U22534 (N_22534,N_22102,N_20700);
nor U22535 (N_22535,N_20698,N_20671);
nand U22536 (N_22536,N_20169,N_20066);
or U22537 (N_22537,N_20064,N_20769);
or U22538 (N_22538,N_21941,N_22293);
nor U22539 (N_22539,N_20109,N_22109);
nand U22540 (N_22540,N_22317,N_21831);
and U22541 (N_22541,N_20384,N_20484);
or U22542 (N_22542,N_21058,N_20326);
xor U22543 (N_22543,N_21345,N_21665);
nand U22544 (N_22544,N_20681,N_21686);
and U22545 (N_22545,N_21639,N_21783);
xor U22546 (N_22546,N_21501,N_22003);
nor U22547 (N_22547,N_22140,N_20217);
nand U22548 (N_22548,N_22257,N_22352);
or U22549 (N_22549,N_21603,N_22221);
and U22550 (N_22550,N_20890,N_21500);
nor U22551 (N_22551,N_21949,N_21182);
xor U22552 (N_22552,N_21926,N_20960);
nand U22553 (N_22553,N_21256,N_20417);
or U22554 (N_22554,N_20880,N_20818);
nand U22555 (N_22555,N_22062,N_20265);
and U22556 (N_22556,N_20765,N_20070);
xnor U22557 (N_22557,N_21649,N_20842);
or U22558 (N_22558,N_20154,N_20615);
nor U22559 (N_22559,N_21143,N_20099);
or U22560 (N_22560,N_21746,N_21659);
nor U22561 (N_22561,N_20493,N_20737);
xnor U22562 (N_22562,N_20807,N_20918);
xnor U22563 (N_22563,N_21979,N_21134);
xor U22564 (N_22564,N_22313,N_20044);
or U22565 (N_22565,N_21451,N_22112);
xnor U22566 (N_22566,N_21768,N_20133);
nor U22567 (N_22567,N_22400,N_20521);
nand U22568 (N_22568,N_22145,N_21903);
nand U22569 (N_22569,N_22342,N_21110);
xor U22570 (N_22570,N_20771,N_20789);
and U22571 (N_22571,N_22127,N_20014);
nor U22572 (N_22572,N_21732,N_21327);
and U22573 (N_22573,N_20891,N_22038);
or U22574 (N_22574,N_21269,N_20474);
xor U22575 (N_22575,N_22085,N_22196);
and U22576 (N_22576,N_20917,N_20910);
or U22577 (N_22577,N_21412,N_20806);
and U22578 (N_22578,N_21499,N_20187);
and U22579 (N_22579,N_20831,N_20522);
and U22580 (N_22580,N_20043,N_20879);
xnor U22581 (N_22581,N_20013,N_20196);
and U22582 (N_22582,N_21785,N_22101);
and U22583 (N_22583,N_21991,N_21227);
nor U22584 (N_22584,N_21402,N_21995);
nand U22585 (N_22585,N_22154,N_22220);
xor U22586 (N_22586,N_20676,N_21733);
and U22587 (N_22587,N_20191,N_21021);
and U22588 (N_22588,N_20504,N_22250);
nor U22589 (N_22589,N_20429,N_22280);
xor U22590 (N_22590,N_22451,N_21672);
nand U22591 (N_22591,N_20110,N_20627);
or U22592 (N_22592,N_21988,N_20206);
nor U22593 (N_22593,N_21881,N_21094);
nor U22594 (N_22594,N_20209,N_21385);
xnor U22595 (N_22595,N_20858,N_20132);
nand U22596 (N_22596,N_21563,N_22105);
nor U22597 (N_22597,N_22449,N_21488);
xnor U22598 (N_22598,N_22419,N_21537);
xor U22599 (N_22599,N_22244,N_20621);
xnor U22600 (N_22600,N_21679,N_22039);
or U22601 (N_22601,N_20796,N_21942);
or U22602 (N_22602,N_20298,N_20297);
and U22603 (N_22603,N_22016,N_20886);
xor U22604 (N_22604,N_21474,N_20510);
nand U22605 (N_22605,N_21719,N_20995);
xor U22606 (N_22606,N_21476,N_21260);
xnor U22607 (N_22607,N_21888,N_20666);
nor U22608 (N_22608,N_20365,N_22000);
nor U22609 (N_22609,N_22186,N_22231);
xor U22610 (N_22610,N_20002,N_22010);
or U22611 (N_22611,N_20553,N_20825);
or U22612 (N_22612,N_20904,N_21159);
and U22613 (N_22613,N_20799,N_20358);
xor U22614 (N_22614,N_20409,N_21645);
nor U22615 (N_22615,N_20738,N_22442);
and U22616 (N_22616,N_21800,N_22019);
or U22617 (N_22617,N_21992,N_22033);
nor U22618 (N_22618,N_21641,N_20740);
nor U22619 (N_22619,N_22143,N_22319);
and U22620 (N_22620,N_21265,N_21169);
nand U22621 (N_22621,N_21360,N_21258);
xor U22622 (N_22622,N_21075,N_20866);
and U22623 (N_22623,N_21723,N_20035);
or U22624 (N_22624,N_21811,N_21290);
and U22625 (N_22625,N_20673,N_20076);
xnor U22626 (N_22626,N_21190,N_21299);
xnor U22627 (N_22627,N_21849,N_20084);
xnor U22628 (N_22628,N_22359,N_21388);
or U22629 (N_22629,N_20134,N_21502);
nor U22630 (N_22630,N_21183,N_20688);
and U22631 (N_22631,N_22264,N_21009);
and U22632 (N_22632,N_20660,N_21173);
or U22633 (N_22633,N_21821,N_20571);
xnor U22634 (N_22634,N_20913,N_21782);
and U22635 (N_22635,N_20585,N_20711);
nor U22636 (N_22636,N_21487,N_22391);
and U22637 (N_22637,N_21635,N_21450);
nor U22638 (N_22638,N_22173,N_20457);
nand U22639 (N_22639,N_21670,N_21709);
or U22640 (N_22640,N_22165,N_21736);
nand U22641 (N_22641,N_20603,N_21088);
nor U22642 (N_22642,N_21423,N_20752);
or U22643 (N_22643,N_21036,N_21370);
and U22644 (N_22644,N_20968,N_22229);
nand U22645 (N_22645,N_20235,N_20466);
or U22646 (N_22646,N_21186,N_21779);
or U22647 (N_22647,N_20231,N_22188);
nor U22648 (N_22648,N_20956,N_20392);
nor U22649 (N_22649,N_20742,N_20227);
or U22650 (N_22650,N_20993,N_20216);
nor U22651 (N_22651,N_21973,N_21323);
or U22652 (N_22652,N_20140,N_21396);
xnor U22653 (N_22653,N_21393,N_21765);
and U22654 (N_22654,N_21205,N_21100);
xor U22655 (N_22655,N_20363,N_21264);
xor U22656 (N_22656,N_21914,N_22457);
and U22657 (N_22657,N_22492,N_20868);
nor U22658 (N_22658,N_22096,N_21781);
xor U22659 (N_22659,N_21271,N_20939);
nor U22660 (N_22660,N_21122,N_21063);
or U22661 (N_22661,N_20884,N_20381);
xor U22662 (N_22662,N_22373,N_22026);
nor U22663 (N_22663,N_21507,N_22118);
or U22664 (N_22664,N_21523,N_20533);
and U22665 (N_22665,N_20017,N_20586);
nor U22666 (N_22666,N_21911,N_21262);
and U22667 (N_22667,N_21985,N_21998);
xor U22668 (N_22668,N_20844,N_22163);
and U22669 (N_22669,N_20357,N_20515);
nor U22670 (N_22670,N_20116,N_20096);
nand U22671 (N_22671,N_22476,N_20911);
nor U22672 (N_22672,N_21763,N_22015);
nand U22673 (N_22673,N_20130,N_21405);
nor U22674 (N_22674,N_21105,N_20104);
nand U22675 (N_22675,N_20239,N_21987);
or U22676 (N_22676,N_20835,N_21278);
nand U22677 (N_22677,N_21623,N_21825);
xnor U22678 (N_22678,N_21947,N_22242);
nand U22679 (N_22679,N_22226,N_20667);
nor U22680 (N_22680,N_21443,N_21163);
nor U22681 (N_22681,N_21232,N_20458);
nand U22682 (N_22682,N_21661,N_20237);
nand U22683 (N_22683,N_21336,N_20683);
and U22684 (N_22684,N_21644,N_22360);
nand U22685 (N_22685,N_20559,N_22422);
or U22686 (N_22686,N_20170,N_20261);
nand U22687 (N_22687,N_21933,N_20470);
nand U22688 (N_22688,N_20026,N_20949);
and U22689 (N_22689,N_22098,N_20963);
nor U22690 (N_22690,N_20920,N_21626);
and U22691 (N_22691,N_20285,N_20996);
nor U22692 (N_22692,N_21715,N_20090);
or U22693 (N_22693,N_20003,N_21150);
nand U22694 (N_22694,N_20577,N_20287);
xor U22695 (N_22695,N_20185,N_20425);
nor U22696 (N_22696,N_22368,N_20593);
nor U22697 (N_22697,N_20848,N_20992);
nor U22698 (N_22698,N_22023,N_21695);
and U22699 (N_22699,N_21960,N_20094);
and U22700 (N_22700,N_20950,N_21213);
nor U22701 (N_22701,N_20469,N_22069);
xor U22702 (N_22702,N_21442,N_21878);
and U22703 (N_22703,N_21786,N_22322);
or U22704 (N_22704,N_21330,N_21744);
nor U22705 (N_22705,N_20128,N_21229);
xnor U22706 (N_22706,N_20755,N_20408);
or U22707 (N_22707,N_20455,N_22050);
and U22708 (N_22708,N_21238,N_20946);
and U22709 (N_22709,N_21351,N_21352);
nor U22710 (N_22710,N_22286,N_21206);
nand U22711 (N_22711,N_21701,N_21652);
or U22712 (N_22712,N_22114,N_21592);
nor U22713 (N_22713,N_20346,N_20964);
nor U22714 (N_22714,N_20940,N_21480);
and U22715 (N_22715,N_20980,N_21165);
or U22716 (N_22716,N_20350,N_21703);
nor U22717 (N_22717,N_20641,N_20106);
or U22718 (N_22718,N_21617,N_20514);
and U22719 (N_22719,N_20307,N_21452);
nor U22720 (N_22720,N_20612,N_20888);
nor U22721 (N_22721,N_22487,N_20453);
xnor U22722 (N_22722,N_20611,N_22413);
nand U22723 (N_22723,N_21550,N_20756);
xor U22724 (N_22724,N_21092,N_21924);
nor U22725 (N_22725,N_20108,N_21432);
nor U22726 (N_22726,N_21195,N_21717);
or U22727 (N_22727,N_21439,N_22262);
nand U22728 (N_22728,N_21399,N_21710);
nand U22729 (N_22729,N_22281,N_21819);
nor U22730 (N_22730,N_21448,N_21742);
nand U22731 (N_22731,N_21207,N_20811);
nor U22732 (N_22732,N_21671,N_21851);
nand U22733 (N_22733,N_20403,N_20967);
nand U22734 (N_22734,N_21216,N_20887);
nor U22735 (N_22735,N_21688,N_20780);
xor U22736 (N_22736,N_21052,N_21918);
and U22737 (N_22737,N_20062,N_20933);
nand U22738 (N_22738,N_20941,N_21263);
and U22739 (N_22739,N_20012,N_21339);
nand U22740 (N_22740,N_21820,N_20855);
xor U22741 (N_22741,N_21721,N_21463);
nand U22742 (N_22742,N_22327,N_20473);
and U22743 (N_22743,N_20784,N_21016);
xnor U22744 (N_22744,N_22110,N_20924);
and U22745 (N_22745,N_21266,N_22007);
nor U22746 (N_22746,N_20863,N_20220);
nand U22747 (N_22747,N_22454,N_20304);
xor U22748 (N_22748,N_22309,N_22387);
nand U22749 (N_22749,N_20311,N_20822);
nor U22750 (N_22750,N_21589,N_21683);
and U22751 (N_22751,N_21362,N_21072);
nor U22752 (N_22752,N_21981,N_21254);
and U22753 (N_22753,N_20150,N_20814);
or U22754 (N_22754,N_22399,N_22377);
xor U22755 (N_22755,N_20545,N_20411);
and U22756 (N_22756,N_21656,N_21752);
xor U22757 (N_22757,N_20147,N_20800);
and U22758 (N_22758,N_20063,N_22170);
and U22759 (N_22759,N_20397,N_21775);
nor U22760 (N_22760,N_21251,N_21066);
or U22761 (N_22761,N_20481,N_20720);
nand U22762 (N_22762,N_21001,N_21139);
or U22763 (N_22763,N_21615,N_21404);
or U22764 (N_22764,N_21113,N_22304);
or U22765 (N_22765,N_20291,N_20762);
nand U22766 (N_22766,N_20229,N_20337);
nor U22767 (N_22767,N_20230,N_20399);
nand U22768 (N_22768,N_22357,N_20450);
nor U22769 (N_22769,N_21731,N_20065);
or U22770 (N_22770,N_21877,N_21261);
or U22771 (N_22771,N_21974,N_21347);
nor U22772 (N_22772,N_21417,N_20146);
xnor U22773 (N_22773,N_20826,N_20373);
or U22774 (N_22774,N_21803,N_22084);
nand U22775 (N_22775,N_20749,N_20345);
and U22776 (N_22776,N_21040,N_20573);
xnor U22777 (N_22777,N_22292,N_22031);
nor U22778 (N_22778,N_20754,N_21335);
and U22779 (N_22779,N_21607,N_21243);
or U22780 (N_22780,N_22215,N_21189);
nor U22781 (N_22781,N_22372,N_21303);
nor U22782 (N_22782,N_20344,N_21793);
nand U22783 (N_22783,N_21891,N_22022);
and U22784 (N_22784,N_21031,N_22208);
nor U22785 (N_22785,N_21253,N_20174);
or U22786 (N_22786,N_22395,N_20334);
or U22787 (N_22787,N_20744,N_22040);
and U22788 (N_22788,N_21747,N_22300);
or U22789 (N_22789,N_21904,N_22356);
xnor U22790 (N_22790,N_21632,N_21167);
or U22791 (N_22791,N_20783,N_22273);
xor U22792 (N_22792,N_22049,N_22432);
and U22793 (N_22793,N_22241,N_20439);
and U22794 (N_22794,N_21149,N_22494);
nor U22795 (N_22795,N_22008,N_21753);
xnor U22796 (N_22796,N_21575,N_21226);
nor U22797 (N_22797,N_21449,N_21522);
xnor U22798 (N_22798,N_20902,N_21776);
xnor U22799 (N_22799,N_22094,N_20208);
xnor U22800 (N_22800,N_20016,N_20562);
or U22801 (N_22801,N_20085,N_21468);
nor U22802 (N_22802,N_21527,N_21944);
xor U22803 (N_22803,N_21922,N_20678);
nand U22804 (N_22804,N_20854,N_21220);
and U22805 (N_22805,N_22447,N_22271);
or U22806 (N_22806,N_22222,N_22498);
nor U22807 (N_22807,N_20323,N_22401);
nor U22808 (N_22808,N_20029,N_20308);
nor U22809 (N_22809,N_20316,N_21048);
or U22810 (N_22810,N_22219,N_22336);
nor U22811 (N_22811,N_20341,N_20802);
or U22812 (N_22812,N_21029,N_20978);
and U22813 (N_22813,N_22329,N_21797);
xor U22814 (N_22814,N_21204,N_22128);
nor U22815 (N_22815,N_20772,N_21757);
xor U22816 (N_22816,N_21869,N_21239);
and U22817 (N_22817,N_20629,N_20088);
xnor U22818 (N_22818,N_21491,N_21799);
nand U22819 (N_22819,N_20240,N_21551);
nor U22820 (N_22820,N_22197,N_21095);
or U22821 (N_22821,N_20735,N_21937);
or U22822 (N_22822,N_21473,N_20376);
and U22823 (N_22823,N_22474,N_22305);
and U22824 (N_22824,N_20382,N_21861);
or U22825 (N_22825,N_20351,N_21305);
and U22826 (N_22826,N_21394,N_20489);
xnor U22827 (N_22827,N_20233,N_21334);
xor U22828 (N_22828,N_21267,N_20374);
xor U22829 (N_22829,N_20536,N_22296);
xor U22830 (N_22830,N_20353,N_22048);
or U22831 (N_22831,N_21879,N_21787);
nor U22832 (N_22832,N_21544,N_21378);
or U22833 (N_22833,N_21123,N_20644);
nand U22834 (N_22834,N_21983,N_20194);
nand U22835 (N_22835,N_21140,N_21276);
xor U22836 (N_22836,N_21244,N_20111);
and U22837 (N_22837,N_21125,N_22137);
and U22838 (N_22838,N_21745,N_22497);
nor U22839 (N_22839,N_20253,N_20004);
nor U22840 (N_22840,N_21677,N_22328);
nor U22841 (N_22841,N_21807,N_21430);
nor U22842 (N_22842,N_22130,N_20404);
nor U22843 (N_22843,N_21618,N_21465);
or U22844 (N_22844,N_20386,N_20159);
nand U22845 (N_22845,N_21761,N_21587);
xor U22846 (N_22846,N_21136,N_21837);
nand U22847 (N_22847,N_20268,N_21651);
or U22848 (N_22848,N_21792,N_21069);
or U22849 (N_22849,N_20300,N_20182);
xnor U22850 (N_22850,N_22210,N_20100);
or U22851 (N_22851,N_21602,N_20072);
or U22852 (N_22852,N_21886,N_20916);
or U22853 (N_22853,N_20077,N_20637);
and U22854 (N_22854,N_22083,N_21221);
nand U22855 (N_22855,N_20200,N_20605);
and U22856 (N_22856,N_21564,N_21045);
and U22857 (N_22857,N_21087,N_20616);
xor U22858 (N_22858,N_20258,N_20471);
nand U22859 (N_22859,N_20383,N_20856);
nor U22860 (N_22860,N_22429,N_20418);
nor U22861 (N_22861,N_21726,N_20490);
or U22862 (N_22862,N_22072,N_20028);
or U22863 (N_22863,N_22071,N_20103);
or U22864 (N_22864,N_20677,N_21673);
or U22865 (N_22865,N_20785,N_22174);
and U22866 (N_22866,N_20375,N_22423);
or U22867 (N_22867,N_21364,N_22124);
and U22868 (N_22868,N_21823,N_21311);
or U22869 (N_22869,N_20640,N_21872);
xnor U22870 (N_22870,N_20999,N_20694);
nand U22871 (N_22871,N_22389,N_20565);
nand U22872 (N_22872,N_21466,N_21958);
xor U22873 (N_22873,N_20460,N_21026);
nand U22874 (N_22874,N_21454,N_22473);
and U22875 (N_22875,N_22435,N_20338);
and U22876 (N_22876,N_20056,N_21520);
or U22877 (N_22877,N_20018,N_21498);
nor U22878 (N_22878,N_20168,N_21309);
nor U22879 (N_22879,N_20985,N_22158);
xor U22880 (N_22880,N_20943,N_21322);
xor U22881 (N_22881,N_20944,N_22459);
xor U22882 (N_22882,N_21300,N_21633);
nand U22883 (N_22883,N_21676,N_21383);
and U22884 (N_22884,N_20263,N_21222);
nand U22885 (N_22885,N_20689,N_21078);
xor U22886 (N_22886,N_22164,N_20367);
and U22887 (N_22887,N_21714,N_20867);
xor U22888 (N_22888,N_21556,N_21047);
nand U22889 (N_22889,N_22018,N_21577);
xor U22890 (N_22890,N_20540,N_20039);
nor U22891 (N_22891,N_20480,N_20751);
nand U22892 (N_22892,N_20779,N_21546);
or U22893 (N_22893,N_22346,N_20279);
or U22894 (N_22894,N_21805,N_21156);
and U22895 (N_22895,N_21978,N_20850);
xor U22896 (N_22896,N_20256,N_21489);
nand U22897 (N_22897,N_20511,N_21080);
or U22898 (N_22898,N_20809,N_20274);
nor U22899 (N_22899,N_21737,N_21490);
nand U22900 (N_22900,N_22375,N_20589);
xor U22901 (N_22901,N_20803,N_21464);
xnor U22902 (N_22902,N_21693,N_22180);
nand U22903 (N_22903,N_22020,N_20050);
nand U22904 (N_22904,N_21038,N_21193);
nor U22905 (N_22905,N_22035,N_21539);
nand U22906 (N_22906,N_20712,N_22445);
nand U22907 (N_22907,N_21350,N_21839);
nor U22908 (N_22908,N_20576,N_21774);
nor U22909 (N_22909,N_22479,N_22266);
and U22910 (N_22910,N_20042,N_21606);
nand U22911 (N_22911,N_20402,N_20501);
nor U22912 (N_22912,N_20982,N_21492);
nand U22913 (N_22913,N_21621,N_22200);
or U22914 (N_22914,N_20597,N_22161);
and U22915 (N_22915,N_22464,N_20655);
and U22916 (N_22916,N_21282,N_21735);
and U22917 (N_22917,N_21873,N_21814);
nor U22918 (N_22918,N_22070,N_22082);
xnor U22919 (N_22919,N_20120,N_20927);
and U22920 (N_22920,N_20267,N_20380);
nor U22921 (N_22921,N_20477,N_21482);
nand U22922 (N_22922,N_20000,N_21410);
nor U22923 (N_22923,N_21608,N_20966);
xor U22924 (N_22924,N_21508,N_21209);
nor U22925 (N_22925,N_20859,N_21542);
and U22926 (N_22926,N_22028,N_20984);
nor U22927 (N_22927,N_20183,N_21056);
xor U22928 (N_22928,N_20288,N_21532);
nand U22929 (N_22929,N_21188,N_20262);
xor U22930 (N_22930,N_20391,N_22225);
or U22931 (N_22931,N_21376,N_21840);
or U22932 (N_22932,N_21061,N_22198);
xnor U22933 (N_22933,N_21653,N_21479);
nor U22934 (N_22934,N_22338,N_21916);
nor U22935 (N_22935,N_20219,N_20981);
and U22936 (N_22936,N_22472,N_21711);
or U22937 (N_22937,N_20563,N_21197);
nand U22938 (N_22938,N_22478,N_21912);
nor U22939 (N_22939,N_20878,N_20733);
xor U22940 (N_22940,N_22092,N_21503);
xor U22941 (N_22941,N_20360,N_21977);
xor U22942 (N_22942,N_20622,N_20841);
nand U22943 (N_22943,N_21750,N_20033);
nand U22944 (N_22944,N_21319,N_20036);
nor U22945 (N_22945,N_20937,N_22254);
and U22946 (N_22946,N_21554,N_22162);
xnor U22947 (N_22947,N_21103,N_22149);
xor U22948 (N_22948,N_20584,N_20317);
nor U22949 (N_22949,N_20630,N_21836);
xnor U22950 (N_22950,N_22111,N_21925);
nor U22951 (N_22951,N_20609,N_22404);
and U22952 (N_22952,N_21462,N_22171);
or U22953 (N_22953,N_20221,N_21636);
xor U22954 (N_22954,N_22234,N_22403);
xor U22955 (N_22955,N_20979,N_21091);
nand U22956 (N_22956,N_20770,N_22441);
nor U22957 (N_22957,N_20575,N_22224);
xnor U22958 (N_22958,N_20086,N_22320);
and U22959 (N_22959,N_21344,N_20152);
nand U22960 (N_22960,N_22298,N_21363);
and U22961 (N_22961,N_20158,N_20596);
xor U22962 (N_22962,N_20554,N_20273);
xor U22963 (N_22963,N_22211,N_21860);
or U22964 (N_22964,N_22202,N_22267);
xnor U22965 (N_22965,N_20889,N_21484);
xnor U22966 (N_22966,N_21403,N_22284);
and U22967 (N_22967,N_20899,N_21968);
nand U22968 (N_22968,N_20687,N_20530);
nor U22969 (N_22969,N_21033,N_20122);
xnor U22970 (N_22970,N_20624,N_20447);
or U22971 (N_22971,N_22260,N_20746);
xnor U22972 (N_22972,N_21601,N_21855);
or U22973 (N_22973,N_21014,N_22121);
and U22974 (N_22974,N_22408,N_20024);
xnor U22975 (N_22975,N_21098,N_20327);
xor U22976 (N_22976,N_21822,N_20732);
or U22977 (N_22977,N_20517,N_20025);
or U22978 (N_22978,N_20781,N_20777);
xor U22979 (N_22979,N_21286,N_20923);
nor U22980 (N_22980,N_20872,N_21441);
xnor U22981 (N_22981,N_21023,N_22374);
and U22982 (N_22982,N_20894,N_20815);
and U22983 (N_22983,N_20449,N_21081);
nor U22984 (N_22984,N_21982,N_21905);
nor U22985 (N_22985,N_20652,N_21340);
xnor U22986 (N_22986,N_20415,N_21953);
nor U22987 (N_22987,N_20468,N_22378);
nand U22988 (N_22988,N_20582,N_21758);
nand U22989 (N_22989,N_21177,N_20567);
nor U22990 (N_22990,N_20606,N_22079);
nand U22991 (N_22991,N_21060,N_20843);
and U22992 (N_22992,N_20936,N_21510);
nand U22993 (N_22993,N_21841,N_21371);
xnor U22994 (N_22994,N_21863,N_20177);
xor U22995 (N_22995,N_21852,N_20723);
and U22996 (N_22996,N_20820,N_22351);
and U22997 (N_22997,N_21691,N_20531);
nand U22998 (N_22998,N_21109,N_20734);
xnor U22999 (N_22999,N_20019,N_20275);
or U23000 (N_23000,N_20117,N_22269);
nor U23001 (N_23001,N_21333,N_21610);
xor U23002 (N_23002,N_20551,N_21273);
nand U23003 (N_23003,N_22141,N_20349);
xor U23004 (N_23004,N_20503,N_21730);
nand U23005 (N_23005,N_20527,N_20211);
nor U23006 (N_23006,N_21921,N_20895);
xnor U23007 (N_23007,N_20234,N_20921);
nand U23008 (N_23008,N_20252,N_21684);
and U23009 (N_23009,N_21416,N_22064);
nand U23010 (N_23010,N_21218,N_22347);
nor U23011 (N_23011,N_20143,N_22063);
xor U23012 (N_23012,N_20015,N_20741);
nor U23013 (N_23013,N_20729,N_20714);
or U23014 (N_23014,N_22136,N_20142);
nand U23015 (N_23015,N_20876,N_21337);
and U23016 (N_23016,N_20883,N_20436);
xor U23017 (N_23017,N_20102,N_21838);
and U23018 (N_23018,N_20764,N_20974);
or U23019 (N_23019,N_20310,N_20225);
or U23020 (N_23020,N_21240,N_21808);
xor U23021 (N_23021,N_21538,N_21071);
or U23022 (N_23022,N_21421,N_20707);
nand U23023 (N_23023,N_22424,N_22480);
xnor U23024 (N_23024,N_21086,N_20739);
and U23025 (N_23025,N_21660,N_20587);
nand U23026 (N_23026,N_21434,N_21917);
nand U23027 (N_23027,N_20162,N_21475);
nor U23028 (N_23028,N_20997,N_21980);
nand U23029 (N_23029,N_21935,N_22376);
xor U23030 (N_23030,N_20126,N_20054);
nand U23031 (N_23031,N_20849,N_20544);
and U23032 (N_23032,N_20074,N_21697);
and U23033 (N_23033,N_21366,N_22394);
or U23034 (N_23034,N_21516,N_20724);
nand U23035 (N_23035,N_20634,N_21077);
xnor U23036 (N_23036,N_20362,N_21591);
nand U23037 (N_23037,N_21131,N_20433);
nor U23038 (N_23038,N_22153,N_21984);
and U23039 (N_23039,N_22446,N_20314);
or U23040 (N_23040,N_21749,N_20476);
nor U23041 (N_23041,N_20271,N_20405);
nor U23042 (N_23042,N_22418,N_21354);
nor U23043 (N_23043,N_21959,N_22443);
and U23044 (N_23044,N_21096,N_20670);
xnor U23045 (N_23045,N_20333,N_20479);
nand U23046 (N_23046,N_21348,N_22306);
or U23047 (N_23047,N_21630,N_20846);
and U23048 (N_23048,N_21248,N_20564);
nand U23049 (N_23049,N_20931,N_22243);
nand U23050 (N_23050,N_20073,N_21798);
nand U23051 (N_23051,N_22312,N_20601);
nor U23052 (N_23052,N_20788,N_21826);
nor U23053 (N_23053,N_22055,N_22076);
nor U23054 (N_23054,N_20801,N_20512);
nand U23055 (N_23055,N_21338,N_21514);
and U23056 (N_23056,N_22183,N_20148);
or U23057 (N_23057,N_20199,N_20976);
or U23058 (N_23058,N_21114,N_22425);
and U23059 (N_23059,N_21329,N_21034);
and U23060 (N_23060,N_20614,N_21424);
nand U23061 (N_23061,N_20797,N_21724);
and U23062 (N_23062,N_20197,N_22006);
nand U23063 (N_23063,N_20038,N_20368);
xnor U23064 (N_23064,N_21164,N_20590);
xnor U23065 (N_23065,N_20994,N_21124);
nand U23066 (N_23066,N_22179,N_21318);
or U23067 (N_23067,N_21358,N_21064);
nor U23068 (N_23068,N_20549,N_21874);
and U23069 (N_23069,N_20773,N_20041);
or U23070 (N_23070,N_21574,N_20226);
or U23071 (N_23071,N_21000,N_20176);
xnor U23072 (N_23072,N_21494,N_21241);
xnor U23073 (N_23073,N_21413,N_21082);
xor U23074 (N_23074,N_21611,N_21127);
xor U23075 (N_23075,N_20516,N_20786);
xor U23076 (N_23076,N_20692,N_22393);
nand U23077 (N_23077,N_21233,N_22024);
nand U23078 (N_23078,N_22496,N_21485);
and U23079 (N_23079,N_21157,N_20581);
nor U23080 (N_23080,N_21553,N_20912);
nor U23081 (N_23081,N_21547,N_20149);
nor U23082 (N_23082,N_22235,N_20804);
xnor U23083 (N_23083,N_21862,N_20875);
or U23084 (N_23084,N_20173,N_21549);
and U23085 (N_23085,N_20715,N_22061);
or U23086 (N_23086,N_20205,N_21024);
and U23087 (N_23087,N_22406,N_21155);
nor U23088 (N_23088,N_20900,N_20975);
nor U23089 (N_23089,N_21766,N_20926);
and U23090 (N_23090,N_22147,N_21093);
or U23091 (N_23091,N_20705,N_21495);
nor U23092 (N_23092,N_20830,N_21631);
nor U23093 (N_23093,N_21268,N_20628);
and U23094 (N_23094,N_21853,N_21280);
nand U23095 (N_23095,N_21687,N_22427);
nor U23096 (N_23096,N_21512,N_21887);
xnor U23097 (N_23097,N_21927,N_22189);
and U23098 (N_23098,N_20699,N_20608);
and U23099 (N_23099,N_22482,N_20874);
nand U23100 (N_23100,N_22288,N_20928);
or U23101 (N_23101,N_20969,N_22277);
and U23102 (N_23102,N_21812,N_21062);
and U23103 (N_23103,N_22282,N_21669);
and U23104 (N_23104,N_21325,N_22236);
or U23105 (N_23105,N_22278,N_20659);
xor U23106 (N_23106,N_20767,N_20882);
xnor U23107 (N_23107,N_20278,N_21097);
or U23108 (N_23108,N_20745,N_21576);
and U23109 (N_23109,N_21307,N_21289);
xor U23110 (N_23110,N_20428,N_20454);
xor U23111 (N_23111,N_21046,N_21647);
and U23112 (N_23112,N_20427,N_21902);
nand U23113 (N_23113,N_20091,N_22086);
nor U23114 (N_23114,N_20834,N_21993);
xor U23115 (N_23115,N_20561,N_21896);
xnor U23116 (N_23116,N_21552,N_20312);
nand U23117 (N_23117,N_21705,N_21971);
nor U23118 (N_23118,N_22316,N_22420);
nor U23119 (N_23119,N_20339,N_21854);
nor U23120 (N_23120,N_20286,N_22100);
xnor U23121 (N_23121,N_21605,N_21919);
xnor U23122 (N_23122,N_22139,N_21590);
nor U23123 (N_23123,N_21535,N_22465);
and U23124 (N_23124,N_20726,N_20343);
nor U23125 (N_23125,N_22001,N_21943);
nand U23126 (N_23126,N_22287,N_21531);
and U23127 (N_23127,N_21788,N_21324);
or U23128 (N_23128,N_22333,N_21108);
or U23129 (N_23129,N_20332,N_21297);
xnor U23130 (N_23130,N_21331,N_22245);
and U23131 (N_23131,N_21252,N_21042);
nor U23132 (N_23132,N_22485,N_21012);
or U23133 (N_23133,N_20195,N_21145);
nor U23134 (N_23134,N_21210,N_20617);
nor U23135 (N_23135,N_21237,N_21832);
nand U23136 (N_23136,N_21357,N_21936);
nor U23137 (N_23137,N_22057,N_21524);
and U23138 (N_23138,N_21445,N_22103);
xnor U23139 (N_23139,N_21754,N_20172);
nor U23140 (N_23140,N_21528,N_20294);
nor U23141 (N_23141,N_21940,N_21966);
and U23142 (N_23142,N_20990,N_21578);
nor U23143 (N_23143,N_22017,N_21249);
xnor U23144 (N_23144,N_20068,N_22195);
or U23145 (N_23145,N_20289,N_22259);
and U23146 (N_23146,N_21461,N_21435);
xnor U23147 (N_23147,N_20594,N_21079);
xor U23148 (N_23148,N_21409,N_20212);
or U23149 (N_23149,N_22059,N_22047);
nand U23150 (N_23150,N_21864,N_20218);
or U23151 (N_23151,N_20060,N_22067);
and U23152 (N_23152,N_21277,N_20697);
or U23153 (N_23153,N_22261,N_21868);
nand U23154 (N_23154,N_21681,N_20535);
nor U23155 (N_23155,N_20426,N_21217);
nand U23156 (N_23156,N_22438,N_20708);
nand U23157 (N_23157,N_20491,N_21882);
or U23158 (N_23158,N_21037,N_20961);
and U23159 (N_23159,N_21596,N_21569);
and U23160 (N_23160,N_20574,N_21562);
and U23161 (N_23161,N_21469,N_21418);
or U23162 (N_23162,N_20620,N_20423);
nor U23163 (N_23163,N_21612,N_20721);
nand U23164 (N_23164,N_22152,N_22157);
xnor U23165 (N_23165,N_22046,N_20682);
nand U23166 (N_23166,N_21530,N_20684);
nor U23167 (N_23167,N_20548,N_22358);
nand U23168 (N_23168,N_22237,N_20580);
nor U23169 (N_23169,N_22392,N_21595);
or U23170 (N_23170,N_20812,N_22354);
nand U23171 (N_23171,N_21467,N_20184);
or U23172 (N_23172,N_22251,N_21778);
and U23173 (N_23173,N_20171,N_22407);
and U23174 (N_23174,N_20255,N_20602);
or U23175 (N_23175,N_20435,N_20276);
xnor U23176 (N_23176,N_21743,N_21712);
nand U23177 (N_23177,N_21898,N_22444);
or U23178 (N_23178,N_21089,N_20761);
nor U23179 (N_23179,N_20853,N_22081);
xor U23180 (N_23180,N_20301,N_21722);
nor U23181 (N_23181,N_20011,N_20523);
or U23182 (N_23182,N_21208,N_21906);
nor U23183 (N_23183,N_20758,N_20824);
nor U23184 (N_23184,N_20328,N_20541);
xor U23185 (N_23185,N_20862,N_21521);
nor U23186 (N_23186,N_20400,N_21901);
nand U23187 (N_23187,N_21184,N_22213);
nand U23188 (N_23188,N_20166,N_21773);
xor U23189 (N_23189,N_21954,N_20371);
and U23190 (N_23190,N_20005,N_21585);
nor U23191 (N_23191,N_21457,N_20970);
nand U23192 (N_23192,N_20556,N_22248);
nor U23193 (N_23193,N_20626,N_21567);
nand U23194 (N_23194,N_20579,N_21809);
nand U23195 (N_23195,N_20896,N_20095);
nor U23196 (N_23196,N_22021,N_21308);
nor U23197 (N_23197,N_20753,N_21477);
nand U23198 (N_23198,N_22415,N_20915);
xnor U23199 (N_23199,N_21022,N_20600);
xor U23200 (N_23200,N_22012,N_21497);
or U23201 (N_23201,N_21583,N_20925);
or U23202 (N_23202,N_21972,N_21967);
nor U23203 (N_23203,N_20293,N_21291);
or U23204 (N_23204,N_21767,N_20865);
nor U23205 (N_23205,N_22205,N_20922);
nand U23206 (N_23206,N_20204,N_21420);
nor U23207 (N_23207,N_20465,N_20494);
or U23208 (N_23208,N_21304,N_21200);
nand U23209 (N_23209,N_20290,N_21880);
nand U23210 (N_23210,N_21440,N_21894);
nand U23211 (N_23211,N_20040,N_21433);
xnor U23212 (N_23212,N_21201,N_22434);
and U23213 (N_23213,N_20977,N_20986);
xor U23214 (N_23214,N_20656,N_20055);
and U23215 (N_23215,N_21784,N_20693);
nor U23216 (N_23216,N_22364,N_22150);
or U23217 (N_23217,N_22499,N_21076);
nand U23218 (N_23218,N_20053,N_20914);
and U23219 (N_23219,N_21437,N_22272);
and U23220 (N_23220,N_20817,N_21035);
or U23221 (N_23221,N_20813,N_21178);
nor U23222 (N_23222,N_22053,N_21142);
and U23223 (N_23223,N_21456,N_22177);
and U23224 (N_23224,N_21956,N_21909);
nor U23225 (N_23225,N_22462,N_20759);
xor U23226 (N_23226,N_20663,N_20164);
or U23227 (N_23227,N_20324,N_22240);
or U23228 (N_23228,N_20354,N_21342);
nand U23229 (N_23229,N_21830,N_20161);
and U23230 (N_23230,N_22468,N_20089);
nand U23231 (N_23231,N_21640,N_21884);
nor U23232 (N_23232,N_21288,N_21115);
or U23233 (N_23233,N_21422,N_22290);
xor U23234 (N_23234,N_22253,N_20636);
nand U23235 (N_23235,N_20958,N_21375);
or U23236 (N_23236,N_20760,N_20305);
nor U23237 (N_23237,N_21622,N_22371);
or U23238 (N_23238,N_21728,N_20898);
or U23239 (N_23239,N_21126,N_21006);
and U23240 (N_23240,N_20047,N_22117);
and U23241 (N_23241,N_21525,N_22002);
xor U23242 (N_23242,N_20837,N_20020);
and U23243 (N_23243,N_21316,N_21381);
nand U23244 (N_23244,N_22396,N_20547);
and U23245 (N_23245,N_20080,N_22310);
and U23246 (N_23246,N_22239,N_21148);
nor U23247 (N_23247,N_21073,N_20736);
or U23248 (N_23248,N_20847,N_22009);
nand U23249 (N_23249,N_21613,N_20078);
nand U23250 (N_23250,N_21361,N_21051);
and U23251 (N_23251,N_22343,N_20139);
nand U23252 (N_23252,N_22151,N_21380);
xor U23253 (N_23253,N_21568,N_20082);
nor U23254 (N_23254,N_21815,N_20058);
nor U23255 (N_23255,N_21624,N_21314);
nor U23256 (N_23256,N_21386,N_22142);
or U23257 (N_23257,N_21739,N_21196);
nand U23258 (N_23258,N_20897,N_20665);
and U23259 (N_23259,N_22388,N_21274);
or U23260 (N_23260,N_20248,N_20988);
nand U23261 (N_23261,N_21395,N_21121);
xnor U23262 (N_23262,N_21584,N_22276);
or U23263 (N_23263,N_20647,N_21938);
and U23264 (N_23264,N_21930,N_21321);
or U23265 (N_23265,N_22439,N_20125);
xnor U23266 (N_23266,N_20558,N_20244);
nand U23267 (N_23267,N_21230,N_21050);
nor U23268 (N_23268,N_22365,N_20821);
nand U23269 (N_23269,N_21740,N_21281);
or U23270 (N_23270,N_21453,N_21147);
nand U23271 (N_23271,N_20599,N_20555);
and U23272 (N_23272,N_21638,N_21704);
or U23273 (N_23273,N_21970,N_21828);
or U23274 (N_23274,N_20881,N_20008);
nor U23275 (N_23275,N_20827,N_20387);
or U23276 (N_23276,N_22275,N_20377);
nor U23277 (N_23277,N_22192,N_20816);
nand U23278 (N_23278,N_21306,N_21455);
or U23279 (N_23279,N_20467,N_20492);
or U23280 (N_23280,N_20953,N_20696);
and U23281 (N_23281,N_21794,N_20651);
nand U23282 (N_23282,N_22133,N_21192);
or U23283 (N_23283,N_20081,N_20942);
nand U23284 (N_23284,N_20438,N_21680);
nand U23285 (N_23285,N_22175,N_20416);
or U23286 (N_23286,N_21975,N_21509);
xor U23287 (N_23287,N_21425,N_21725);
nand U23288 (N_23288,N_20989,N_21242);
and U23289 (N_23289,N_20215,N_20475);
and U23290 (N_23290,N_21459,N_22058);
nand U23291 (N_23291,N_20658,N_21802);
nor U23292 (N_23292,N_21824,N_20938);
nor U23293 (N_23293,N_20097,N_20462);
nor U23294 (N_23294,N_20568,N_22185);
and U23295 (N_23295,N_20270,N_20497);
xnor U23296 (N_23296,N_20052,N_22314);
xnor U23297 (N_23297,N_20691,N_21162);
or U23298 (N_23298,N_21856,N_21962);
nand U23299 (N_23299,N_20610,N_20839);
xor U23300 (N_23300,N_21326,N_22030);
xor U23301 (N_23301,N_22489,N_22380);
and U23302 (N_23302,N_21472,N_22348);
or U23303 (N_23303,N_20635,N_21866);
nor U23304 (N_23304,N_21663,N_22052);
or U23305 (N_23305,N_21573,N_20569);
nor U23306 (N_23306,N_20165,N_20525);
and U23307 (N_23307,N_21689,N_21438);
xnor U23308 (N_23308,N_21171,N_22088);
or U23309 (N_23309,N_22493,N_20538);
xor U23310 (N_23310,N_20232,N_22416);
nor U23311 (N_23311,N_21827,N_21460);
xor U23312 (N_23312,N_22477,N_21604);
xor U23313 (N_23313,N_20710,N_21102);
and U23314 (N_23314,N_21845,N_20355);
nor U23315 (N_23315,N_21257,N_21414);
nor U23316 (N_23316,N_22176,N_20657);
and U23317 (N_23317,N_21629,N_20101);
nand U23318 (N_23318,N_22044,N_21382);
or U23319 (N_23319,N_20249,N_21945);
or U23320 (N_23320,N_22056,N_21019);
nor U23321 (N_23321,N_20075,N_20372);
nor U23322 (N_23322,N_20124,N_20242);
nor U23323 (N_23323,N_21764,N_21328);
or U23324 (N_23324,N_22249,N_22051);
or U23325 (N_23325,N_21481,N_21203);
nand U23326 (N_23326,N_21368,N_20442);
nor U23327 (N_23327,N_21002,N_21548);
nor U23328 (N_23328,N_21707,N_21493);
nand U23329 (N_23329,N_21225,N_20137);
nand U23330 (N_23330,N_20406,N_20649);
xnor U23331 (N_23331,N_22037,N_22402);
nand U23332 (N_23332,N_20991,N_20959);
xor U23333 (N_23333,N_20524,N_22379);
nor U23334 (N_23334,N_22426,N_21969);
xor U23335 (N_23335,N_21398,N_21951);
or U23336 (N_23336,N_20010,N_22108);
or U23337 (N_23337,N_22054,N_20034);
xnor U23338 (N_23338,N_22323,N_21829);
nand U23339 (N_23339,N_20069,N_22385);
and U23340 (N_23340,N_20421,N_20532);
nor U23341 (N_23341,N_20793,N_20190);
xnor U23342 (N_23342,N_20828,N_20864);
and U23343 (N_23343,N_21343,N_20546);
nor U23344 (N_23344,N_22467,N_22078);
or U23345 (N_23345,N_20303,N_20045);
and U23346 (N_23346,N_21146,N_22471);
or U23347 (N_23347,N_22097,N_21700);
nand U23348 (N_23348,N_20145,N_22349);
nor U23349 (N_23349,N_21835,N_21555);
and U23350 (N_23350,N_21160,N_21598);
xnor U23351 (N_23351,N_21401,N_20619);
nand U23352 (N_23352,N_21990,N_21294);
xnor U23353 (N_23353,N_20543,N_20722);
nor U23354 (N_23354,N_20604,N_20901);
and U23355 (N_23355,N_21070,N_21847);
nand U23356 (N_23356,N_21099,N_22113);
and U23357 (N_23357,N_20983,N_21074);
or U23358 (N_23358,N_20163,N_20407);
nor U23359 (N_23359,N_21892,N_20264);
nand U23360 (N_23360,N_20437,N_21408);
xnor U23361 (N_23361,N_21920,N_20131);
nor U23362 (N_23362,N_21646,N_21144);
or U23363 (N_23363,N_20236,N_21907);
xor U23364 (N_23364,N_20507,N_21118);
xor U23365 (N_23365,N_21561,N_21374);
or U23366 (N_23366,N_20023,N_21317);
xor U23367 (N_23367,N_20370,N_21053);
nor U23368 (N_23368,N_22475,N_21228);
nand U23369 (N_23369,N_21250,N_20228);
or U23370 (N_23370,N_22324,N_21729);
and U23371 (N_23371,N_21392,N_21030);
nand U23372 (N_23372,N_21580,N_21513);
nand U23373 (N_23373,N_22431,N_21994);
xnor U23374 (N_23374,N_21172,N_20118);
or U23375 (N_23375,N_22453,N_21471);
nand U23376 (N_23376,N_20623,N_21895);
xnor U23377 (N_23377,N_20266,N_21285);
xor U23378 (N_23378,N_22065,N_22138);
nand U23379 (N_23379,N_21961,N_21428);
nand U23380 (N_23380,N_20318,N_20907);
nor U23381 (N_23381,N_20445,N_20001);
xor U23382 (N_23382,N_20643,N_21526);
nand U23383 (N_23383,N_20537,N_22209);
nand U23384 (N_23384,N_21519,N_22340);
nor U23385 (N_23385,N_20852,N_20595);
or U23386 (N_23386,N_21356,N_22263);
and U23387 (N_23387,N_22367,N_21637);
nand U23388 (N_23388,N_20908,N_20434);
or U23389 (N_23389,N_21234,N_20356);
nand U23390 (N_23390,N_20775,N_21682);
nor U23391 (N_23391,N_21529,N_22204);
nor U23392 (N_23392,N_21359,N_21795);
or U23393 (N_23393,N_21270,N_21727);
nand U23394 (N_23394,N_20790,N_22430);
nand U23395 (N_23395,N_21120,N_20948);
xor U23396 (N_23396,N_21834,N_20284);
nor U23397 (N_23397,N_21135,N_20798);
and U23398 (N_23398,N_21161,N_22325);
and U23399 (N_23399,N_22217,N_22246);
xor U23400 (N_23400,N_22436,N_22410);
xnor U23401 (N_23401,N_21486,N_22448);
nand U23402 (N_23402,N_20478,N_21017);
nor U23403 (N_23403,N_20393,N_20728);
nand U23404 (N_23404,N_20342,N_20135);
and U23405 (N_23405,N_20782,N_21390);
nor U23406 (N_23406,N_21511,N_21315);
nand U23407 (N_23407,N_22042,N_20520);
nor U23408 (N_23408,N_22469,N_21560);
or U23409 (N_23409,N_20987,N_20155);
xnor U23410 (N_23410,N_20379,N_21236);
and U23411 (N_23411,N_21406,N_21557);
and U23412 (N_23412,N_20792,N_20935);
xnor U23413 (N_23413,N_22014,N_21130);
nor U23414 (N_23414,N_20713,N_20795);
and U23415 (N_23415,N_20247,N_22169);
or U23416 (N_23416,N_20389,N_20743);
nand U23417 (N_23417,N_20838,N_21734);
xor U23418 (N_23418,N_20251,N_22181);
nand U23419 (N_23419,N_21180,N_21426);
nor U23420 (N_23420,N_20528,N_22207);
xor U23421 (N_23421,N_22461,N_22034);
xor U23422 (N_23422,N_22299,N_21153);
nor U23423 (N_23423,N_22172,N_22486);
or U23424 (N_23424,N_21027,N_20550);
and U23425 (N_23425,N_21609,N_21215);
nand U23426 (N_23426,N_21373,N_21885);
and U23427 (N_23427,N_22074,N_22089);
nand U23428 (N_23428,N_20500,N_20093);
or U23429 (N_23429,N_21844,N_20296);
nand U23430 (N_23430,N_20105,N_22361);
and U23431 (N_23431,N_22295,N_21003);
and U23432 (N_23432,N_20552,N_20578);
xor U23433 (N_23433,N_20701,N_20513);
xnor U23434 (N_23434,N_21154,N_20250);
xnor U23435 (N_23435,N_21310,N_20934);
nor U23436 (N_23436,N_21211,N_21769);
nor U23437 (N_23437,N_22491,N_22381);
or U23438 (N_23438,N_20420,N_21067);
xnor U23439 (N_23439,N_20486,N_21597);
nand U23440 (N_23440,N_20716,N_21964);
nand U23441 (N_23441,N_21372,N_20747);
xor U23442 (N_23442,N_22452,N_21559);
xor U23443 (N_23443,N_20607,N_21168);
or U23444 (N_23444,N_20071,N_21049);
and U23445 (N_23445,N_21101,N_21349);
xor U23446 (N_23446,N_21848,N_20870);
or U23447 (N_23447,N_21117,N_20138);
or U23448 (N_23448,N_21235,N_22160);
nand U23449 (N_23449,N_21111,N_20410);
xor U23450 (N_23450,N_20181,N_21558);
or U23451 (N_23451,N_20030,N_20763);
nor U23452 (N_23452,N_20719,N_20153);
nand U23453 (N_23453,N_22187,N_22095);
nor U23454 (N_23454,N_21287,N_21107);
or U23455 (N_23455,N_20329,N_21059);
or U23456 (N_23456,N_20819,N_20718);
nor U23457 (N_23457,N_22119,N_20369);
or U23458 (N_23458,N_20810,N_22307);
nand U23459 (N_23459,N_21976,N_21643);
or U23460 (N_23460,N_20107,N_21948);
or U23461 (N_23461,N_21104,N_21893);
nand U23462 (N_23462,N_20022,N_20905);
nand U23463 (N_23463,N_21582,N_20906);
xor U23464 (N_23464,N_20321,N_20113);
nor U23465 (N_23465,N_20115,N_21843);
nand U23466 (N_23466,N_22227,N_21738);
xor U23467 (N_23467,N_20295,N_21119);
or U23468 (N_23468,N_21713,N_20452);
or U23469 (N_23469,N_22252,N_21332);
xnor U23470 (N_23470,N_21518,N_21586);
xnor U23471 (N_23471,N_20526,N_21279);
or U23472 (N_23472,N_22087,N_20046);
xnor U23473 (N_23473,N_22330,N_20441);
and U23474 (N_23474,N_21379,N_21870);
and U23475 (N_23475,N_21816,N_21504);
and U23476 (N_23476,N_21889,N_20260);
or U23477 (N_23477,N_20189,N_21044);
nor U23478 (N_23478,N_20957,N_21899);
nor U23479 (N_23479,N_21957,N_21541);
nor U23480 (N_23480,N_21313,N_20087);
and U23481 (N_23481,N_22450,N_20583);
nor U23482 (N_23482,N_21255,N_21065);
xor U23483 (N_23483,N_22466,N_21875);
or U23484 (N_23484,N_21355,N_21565);
and U23485 (N_23485,N_20464,N_22218);
xor U23486 (N_23486,N_21791,N_21185);
nor U23487 (N_23487,N_20413,N_20787);
xor U23488 (N_23488,N_20222,N_21090);
xnor U23489 (N_23489,N_21588,N_22004);
nor U23490 (N_23490,N_22488,N_20330);
or U23491 (N_23491,N_22182,N_20193);
and U23492 (N_23492,N_20645,N_20566);
or U23493 (N_23493,N_22326,N_22256);
xnor U23494 (N_23494,N_21224,N_20049);
xor U23495 (N_23495,N_21642,N_21858);
and U23496 (N_23496,N_21259,N_21129);
nor U23497 (N_23497,N_21634,N_20309);
or U23498 (N_23498,N_21212,N_21085);
xnor U23499 (N_23499,N_20591,N_22265);
xnor U23500 (N_23500,N_20306,N_20557);
nand U23501 (N_23501,N_22411,N_22386);
xor U23502 (N_23502,N_22334,N_21708);
nor U23503 (N_23503,N_20654,N_21692);
and U23504 (N_23504,N_22134,N_22129);
nand U23505 (N_23505,N_20998,N_21068);
and U23506 (N_23506,N_21579,N_22178);
nor U23507 (N_23507,N_21806,N_21517);
or U23508 (N_23508,N_20067,N_20871);
and U23509 (N_23509,N_20861,N_21986);
and U23510 (N_23510,N_20588,N_21013);
and U23511 (N_23511,N_20954,N_22409);
xor U23512 (N_23512,N_21295,N_20331);
nand U23513 (N_23513,N_21690,N_20487);
nor U23514 (N_23514,N_20009,N_22043);
nor U23515 (N_23515,N_22311,N_21600);
nand U23516 (N_23516,N_22027,N_21415);
or U23517 (N_23517,N_22350,N_20774);
nor U23518 (N_23518,N_22238,N_22011);
nand U23519 (N_23519,N_22045,N_20823);
nand U23520 (N_23520,N_21857,N_22332);
xnor U23521 (N_23521,N_21400,N_22068);
nand U23522 (N_23522,N_22390,N_21187);
nand U23523 (N_23523,N_21702,N_20424);
or U23524 (N_23524,N_20430,N_20506);
and U23525 (N_23525,N_20680,N_22363);
xor U23526 (N_23526,N_20207,N_22495);
nor U23527 (N_23527,N_20347,N_22206);
or U23528 (N_23528,N_21545,N_20129);
nand U23529 (N_23529,N_21572,N_20348);
or U23530 (N_23530,N_20833,N_20495);
xnor U23531 (N_23531,N_20027,N_20151);
nand U23532 (N_23532,N_20725,N_22148);
or U23533 (N_23533,N_21116,N_22166);
and U23534 (N_23534,N_21540,N_20570);
nand U23535 (N_23535,N_21932,N_20451);
nand U23536 (N_23536,N_22291,N_22077);
and U23537 (N_23537,N_22398,N_20560);
and U23538 (N_23538,N_22125,N_22115);
xnor U23539 (N_23539,N_20167,N_21771);
nand U23540 (N_23540,N_21593,N_21900);
and U23541 (N_23541,N_22104,N_20704);
nor U23542 (N_23542,N_22369,N_20456);
nor U23543 (N_23543,N_20947,N_20542);
or U23544 (N_23544,N_22428,N_20061);
nand U23545 (N_23545,N_20114,N_20007);
and U23546 (N_23546,N_22041,N_20254);
or U23547 (N_23547,N_20282,N_22144);
or U23548 (N_23548,N_21929,N_20112);
or U23549 (N_23549,N_21353,N_20836);
nand U23550 (N_23550,N_20748,N_21231);
nor U23551 (N_23551,N_22460,N_20805);
xnor U23552 (N_23552,N_20971,N_20179);
xnor U23553 (N_23553,N_21174,N_22308);
nand U23554 (N_23554,N_21367,N_20829);
xor U23555 (N_23555,N_21483,N_21015);
nor U23556 (N_23556,N_21458,N_21341);
nor U23557 (N_23557,N_20083,N_22303);
xor U23558 (N_23558,N_21055,N_22366);
nand U23559 (N_23559,N_22362,N_20299);
and U23560 (N_23560,N_22184,N_22289);
and U23561 (N_23561,N_21772,N_20973);
or U23562 (N_23562,N_20791,N_21181);
and U23563 (N_23563,N_22463,N_21674);
nor U23564 (N_23564,N_20648,N_20572);
and U23565 (N_23565,N_21627,N_21718);
nand U23566 (N_23566,N_20778,N_21246);
nor U23567 (N_23567,N_21429,N_22297);
nor U23568 (N_23568,N_22458,N_20127);
nand U23569 (N_23569,N_22159,N_20539);
nand U23570 (N_23570,N_22255,N_20245);
nor U23571 (N_23571,N_20048,N_20962);
nor U23572 (N_23572,N_22339,N_20951);
nor U23573 (N_23573,N_20440,N_20092);
nand U23574 (N_23574,N_20488,N_21846);
and U23575 (N_23575,N_21427,N_21032);
xor U23576 (N_23576,N_21817,N_20443);
xor U23577 (N_23577,N_20302,N_21619);
nand U23578 (N_23578,N_21446,N_21755);
or U23579 (N_23579,N_20180,N_22470);
and U23580 (N_23580,N_21025,N_21298);
nand U23581 (N_23581,N_22120,N_20703);
nand U23582 (N_23582,N_20598,N_21908);
or U23583 (N_23583,N_22135,N_21694);
or U23584 (N_23584,N_20892,N_20679);
nand U23585 (N_23585,N_20932,N_20750);
nor U23586 (N_23586,N_21028,N_22230);
nor U23587 (N_23587,N_20059,N_20945);
xnor U23588 (N_23588,N_20246,N_20098);
or U23589 (N_23589,N_22036,N_22132);
xor U23590 (N_23590,N_21365,N_20534);
and U23591 (N_23591,N_20840,N_21447);
or U23592 (N_23592,N_21751,N_21859);
nor U23593 (N_23593,N_20674,N_20178);
xnor U23594 (N_23594,N_22270,N_22331);
or U23595 (N_23595,N_20461,N_22199);
or U23596 (N_23596,N_22091,N_22384);
nor U23597 (N_23597,N_20203,N_22490);
nand U23598 (N_23598,N_20519,N_20717);
xor U23599 (N_23599,N_20877,N_22345);
nand U23600 (N_23600,N_20483,N_20776);
nor U23601 (N_23601,N_20668,N_22212);
nor U23602 (N_23602,N_21112,N_20259);
and U23603 (N_23603,N_21293,N_21008);
xnor U23604 (N_23604,N_21151,N_21369);
xor U23605 (N_23605,N_20198,N_20224);
xor U23606 (N_23606,N_22433,N_20272);
or U23607 (N_23607,N_21057,N_20632);
nand U23608 (N_23608,N_20315,N_22029);
nand U23609 (N_23609,N_22194,N_20156);
and U23610 (N_23610,N_20730,N_21054);
and U23611 (N_23611,N_22025,N_22073);
and U23612 (N_23612,N_22302,N_21989);
xor U23613 (N_23613,N_20631,N_20766);
nor U23614 (N_23614,N_21923,N_20320);
nor U23615 (N_23615,N_21871,N_20432);
and U23616 (N_23616,N_22301,N_21275);
and U23617 (N_23617,N_21411,N_20496);
xnor U23618 (N_23618,N_20690,N_22268);
nand U23619 (N_23619,N_20832,N_21515);
or U23620 (N_23620,N_20518,N_20340);
nor U23621 (N_23621,N_21138,N_21005);
nand U23622 (N_23622,N_20873,N_20395);
xnor U23623 (N_23623,N_22167,N_22337);
nand U23624 (N_23624,N_21867,N_21478);
or U23625 (N_23625,N_22131,N_22116);
or U23626 (N_23626,N_20385,N_20157);
nand U23627 (N_23627,N_21789,N_22274);
and U23628 (N_23628,N_20280,N_20277);
or U23629 (N_23629,N_20175,N_21292);
nand U23630 (N_23630,N_20188,N_21007);
nand U23631 (N_23631,N_22146,N_21419);
or U23632 (N_23632,N_21302,N_21245);
and U23633 (N_23633,N_21397,N_21770);
and U23634 (N_23634,N_21759,N_20223);
or U23635 (N_23635,N_20952,N_21796);
nor U23636 (N_23636,N_21658,N_22353);
or U23637 (N_23637,N_21170,N_20731);
or U23638 (N_23638,N_22417,N_21950);
and U23639 (N_23639,N_21760,N_20401);
xor U23640 (N_23640,N_21668,N_22341);
xor U23641 (N_23641,N_21219,N_21581);
xor U23642 (N_23642,N_21534,N_22107);
or U23643 (N_23643,N_20366,N_20650);
nand U23644 (N_23644,N_22156,N_20021);
nand U23645 (N_23645,N_20006,N_20419);
or U23646 (N_23646,N_22440,N_20613);
and U23647 (N_23647,N_21928,N_20192);
nor U23648 (N_23648,N_21436,N_20364);
nand U23649 (N_23649,N_20322,N_21377);
and U23650 (N_23650,N_20388,N_21137);
and U23651 (N_23651,N_22335,N_21833);
or U23652 (N_23652,N_21915,N_20394);
xor U23653 (N_23653,N_21720,N_22279);
xnor U23654 (N_23654,N_20051,N_20210);
and U23655 (N_23655,N_21391,N_20359);
and U23656 (N_23656,N_22318,N_20079);
and U23657 (N_23657,N_21801,N_22060);
nor U23658 (N_23658,N_21571,N_20757);
or U23659 (N_23659,N_21685,N_22414);
or U23660 (N_23660,N_21842,N_21505);
xor U23661 (N_23661,N_21570,N_20057);
nand U23662 (N_23662,N_20499,N_22484);
and U23663 (N_23663,N_21952,N_20281);
xor U23664 (N_23664,N_21997,N_21041);
or U23665 (N_23665,N_21011,N_21913);
and U23666 (N_23666,N_21654,N_20412);
and U23667 (N_23667,N_21133,N_20498);
nand U23668 (N_23668,N_21179,N_20930);
or U23669 (N_23669,N_22090,N_20144);
xnor U23670 (N_23670,N_21470,N_21166);
and U23671 (N_23671,N_21506,N_22190);
and U23672 (N_23672,N_21790,N_20431);
nand U23673 (N_23673,N_20123,N_22344);
nor U23674 (N_23674,N_21191,N_20292);
nand U23675 (N_23675,N_20664,N_20639);
or U23676 (N_23676,N_21666,N_20448);
xnor U23677 (N_23677,N_22214,N_21296);
xnor U23678 (N_23678,N_20243,N_21083);
nand U23679 (N_23679,N_21223,N_20336);
xnor U23680 (N_23680,N_20686,N_20485);
nor U23681 (N_23681,N_21696,N_21158);
nand U23682 (N_23682,N_21965,N_21931);
nand U23683 (N_23683,N_21741,N_21599);
nor U23684 (N_23684,N_21850,N_20646);
xor U23685 (N_23685,N_21283,N_21662);
nor U23686 (N_23686,N_21616,N_21141);
and U23687 (N_23687,N_21043,N_21407);
nand U23688 (N_23688,N_20505,N_20661);
xnor U23689 (N_23689,N_20633,N_22382);
and U23690 (N_23690,N_22232,N_21004);
nor U23691 (N_23691,N_20214,N_20201);
nor U23692 (N_23692,N_21876,N_21810);
and U23693 (N_23693,N_21748,N_21301);
or U23694 (N_23694,N_22370,N_21084);
and U23695 (N_23695,N_21106,N_22315);
nor U23696 (N_23696,N_20283,N_20136);
nor U23697 (N_23697,N_20141,N_22155);
nand U23698 (N_23698,N_20885,N_22355);
or U23699 (N_23699,N_21431,N_21194);
nand U23700 (N_23700,N_22405,N_21387);
or U23701 (N_23701,N_21625,N_21780);
xnor U23702 (N_23702,N_22013,N_20502);
and U23703 (N_23703,N_21128,N_22228);
xnor U23704 (N_23704,N_22437,N_20508);
and U23705 (N_23705,N_20398,N_22283);
and U23706 (N_23706,N_20119,N_22126);
nor U23707 (N_23707,N_21202,N_22216);
xnor U23708 (N_23708,N_21955,N_22223);
xnor U23709 (N_23709,N_20361,N_21657);
nand U23710 (N_23710,N_22093,N_21444);
or U23711 (N_23711,N_22412,N_21620);
or U23712 (N_23712,N_20444,N_21389);
xor U23713 (N_23713,N_20794,N_21999);
nand U23714 (N_23714,N_22285,N_20860);
or U23715 (N_23715,N_21865,N_22005);
nand U23716 (N_23716,N_20257,N_22168);
or U23717 (N_23717,N_21648,N_20709);
and U23718 (N_23718,N_22294,N_21963);
xnor U23719 (N_23719,N_21813,N_21678);
xor U23720 (N_23720,N_20482,N_21818);
nand U23721 (N_23721,N_21132,N_20768);
or U23722 (N_23722,N_20213,N_20625);
nor U23723 (N_23723,N_21176,N_22106);
and U23724 (N_23724,N_20702,N_22075);
xor U23725 (N_23725,N_22201,N_22258);
xnor U23726 (N_23726,N_20037,N_21667);
and U23727 (N_23727,N_20919,N_20313);
nor U23728 (N_23728,N_21756,N_21996);
xnor U23729 (N_23729,N_22321,N_20396);
or U23730 (N_23730,N_20695,N_21175);
xor U23731 (N_23731,N_20929,N_20414);
nor U23732 (N_23732,N_20238,N_22481);
xnor U23733 (N_23733,N_22080,N_20241);
xor U23734 (N_23734,N_20851,N_20202);
nand U23735 (N_23735,N_21536,N_21533);
and U23736 (N_23736,N_21664,N_20955);
nor U23737 (N_23737,N_21716,N_21934);
xnor U23738 (N_23738,N_21346,N_20638);
or U23739 (N_23739,N_20529,N_20662);
xor U23740 (N_23740,N_20378,N_20965);
nor U23741 (N_23741,N_20463,N_20653);
xor U23742 (N_23742,N_20903,N_22099);
xor U23743 (N_23743,N_21247,N_20857);
xor U23744 (N_23744,N_20642,N_20352);
or U23745 (N_23745,N_21320,N_21496);
or U23746 (N_23746,N_21594,N_21910);
nand U23747 (N_23747,N_21199,N_22203);
xnor U23748 (N_23748,N_20032,N_20472);
xor U23749 (N_23749,N_21010,N_21384);
nor U23750 (N_23750,N_21307,N_20750);
or U23751 (N_23751,N_20661,N_22195);
nand U23752 (N_23752,N_22028,N_22358);
xor U23753 (N_23753,N_21024,N_20882);
or U23754 (N_23754,N_21297,N_22342);
nand U23755 (N_23755,N_20520,N_22418);
or U23756 (N_23756,N_21203,N_21431);
and U23757 (N_23757,N_20377,N_22060);
nand U23758 (N_23758,N_20907,N_20853);
nand U23759 (N_23759,N_21827,N_20652);
nor U23760 (N_23760,N_21549,N_22248);
nand U23761 (N_23761,N_20005,N_21969);
and U23762 (N_23762,N_22193,N_21639);
nand U23763 (N_23763,N_20214,N_20384);
and U23764 (N_23764,N_20582,N_21410);
nor U23765 (N_23765,N_21554,N_20936);
nor U23766 (N_23766,N_20241,N_20575);
and U23767 (N_23767,N_20029,N_22085);
nand U23768 (N_23768,N_21018,N_20430);
or U23769 (N_23769,N_20365,N_21800);
or U23770 (N_23770,N_20768,N_21363);
nor U23771 (N_23771,N_22332,N_21825);
or U23772 (N_23772,N_22326,N_21825);
and U23773 (N_23773,N_21418,N_20783);
nor U23774 (N_23774,N_21925,N_21810);
xnor U23775 (N_23775,N_21266,N_20359);
and U23776 (N_23776,N_20620,N_20008);
nand U23777 (N_23777,N_20269,N_21112);
or U23778 (N_23778,N_20890,N_21682);
nand U23779 (N_23779,N_20733,N_21564);
xor U23780 (N_23780,N_22466,N_20124);
or U23781 (N_23781,N_20000,N_22335);
and U23782 (N_23782,N_21107,N_20205);
xnor U23783 (N_23783,N_22341,N_20288);
xnor U23784 (N_23784,N_21708,N_21278);
and U23785 (N_23785,N_22146,N_21399);
xnor U23786 (N_23786,N_21959,N_22476);
or U23787 (N_23787,N_21478,N_20219);
or U23788 (N_23788,N_21154,N_22037);
or U23789 (N_23789,N_21314,N_20289);
and U23790 (N_23790,N_20796,N_20028);
nor U23791 (N_23791,N_20451,N_20645);
nor U23792 (N_23792,N_22481,N_20195);
nor U23793 (N_23793,N_20154,N_21613);
and U23794 (N_23794,N_21220,N_20903);
nor U23795 (N_23795,N_21457,N_20411);
xor U23796 (N_23796,N_20748,N_20750);
nand U23797 (N_23797,N_21284,N_21148);
xor U23798 (N_23798,N_20724,N_22107);
xor U23799 (N_23799,N_22122,N_22488);
xnor U23800 (N_23800,N_20116,N_21707);
nor U23801 (N_23801,N_21868,N_21030);
or U23802 (N_23802,N_22119,N_21685);
nand U23803 (N_23803,N_21202,N_20690);
xnor U23804 (N_23804,N_20134,N_21031);
nand U23805 (N_23805,N_20170,N_22151);
or U23806 (N_23806,N_22369,N_21605);
or U23807 (N_23807,N_22285,N_21070);
xor U23808 (N_23808,N_20646,N_21248);
nand U23809 (N_23809,N_21978,N_21088);
nor U23810 (N_23810,N_20052,N_20669);
nor U23811 (N_23811,N_21984,N_20308);
nor U23812 (N_23812,N_21732,N_20638);
nand U23813 (N_23813,N_21834,N_21797);
nand U23814 (N_23814,N_21825,N_22059);
nor U23815 (N_23815,N_20881,N_20986);
nor U23816 (N_23816,N_20607,N_20547);
xor U23817 (N_23817,N_20822,N_20662);
xnor U23818 (N_23818,N_20161,N_22244);
nor U23819 (N_23819,N_21295,N_21227);
nor U23820 (N_23820,N_20573,N_22265);
nor U23821 (N_23821,N_20509,N_20083);
nor U23822 (N_23822,N_21924,N_20896);
and U23823 (N_23823,N_20040,N_22416);
and U23824 (N_23824,N_21821,N_21287);
or U23825 (N_23825,N_20507,N_22483);
nand U23826 (N_23826,N_22199,N_22291);
or U23827 (N_23827,N_21158,N_22175);
xor U23828 (N_23828,N_22387,N_21331);
xor U23829 (N_23829,N_21020,N_20919);
or U23830 (N_23830,N_20904,N_20212);
or U23831 (N_23831,N_21948,N_21899);
or U23832 (N_23832,N_20362,N_21997);
or U23833 (N_23833,N_21442,N_20371);
or U23834 (N_23834,N_20189,N_20817);
or U23835 (N_23835,N_21328,N_22044);
xor U23836 (N_23836,N_22405,N_20530);
xnor U23837 (N_23837,N_20654,N_20562);
nor U23838 (N_23838,N_21903,N_22306);
nand U23839 (N_23839,N_22430,N_21797);
nand U23840 (N_23840,N_20814,N_20491);
nand U23841 (N_23841,N_21898,N_20888);
xnor U23842 (N_23842,N_21561,N_20097);
nand U23843 (N_23843,N_21606,N_21998);
and U23844 (N_23844,N_21514,N_20524);
and U23845 (N_23845,N_20762,N_20142);
nand U23846 (N_23846,N_22348,N_20286);
or U23847 (N_23847,N_20660,N_21021);
xor U23848 (N_23848,N_22342,N_21195);
nand U23849 (N_23849,N_21237,N_20026);
nand U23850 (N_23850,N_20736,N_20622);
nor U23851 (N_23851,N_20049,N_21894);
nor U23852 (N_23852,N_20891,N_21566);
xnor U23853 (N_23853,N_21753,N_21654);
xnor U23854 (N_23854,N_21052,N_21810);
nand U23855 (N_23855,N_20400,N_20185);
or U23856 (N_23856,N_22429,N_21373);
xor U23857 (N_23857,N_21399,N_20196);
or U23858 (N_23858,N_21282,N_21240);
nor U23859 (N_23859,N_20525,N_20565);
xor U23860 (N_23860,N_20000,N_20756);
or U23861 (N_23861,N_20732,N_21562);
nand U23862 (N_23862,N_22341,N_22265);
or U23863 (N_23863,N_22171,N_21756);
xnor U23864 (N_23864,N_22401,N_20276);
nor U23865 (N_23865,N_21698,N_21370);
nand U23866 (N_23866,N_22435,N_22168);
or U23867 (N_23867,N_22213,N_21251);
nor U23868 (N_23868,N_20881,N_20052);
and U23869 (N_23869,N_21681,N_20781);
or U23870 (N_23870,N_21363,N_20545);
or U23871 (N_23871,N_21925,N_20174);
xnor U23872 (N_23872,N_20803,N_21443);
nand U23873 (N_23873,N_22403,N_20749);
xnor U23874 (N_23874,N_20211,N_20741);
and U23875 (N_23875,N_21663,N_20695);
xor U23876 (N_23876,N_22176,N_20229);
xnor U23877 (N_23877,N_22425,N_20958);
xor U23878 (N_23878,N_20969,N_21911);
or U23879 (N_23879,N_21251,N_21340);
and U23880 (N_23880,N_21944,N_20876);
or U23881 (N_23881,N_21749,N_21775);
xnor U23882 (N_23882,N_21548,N_21150);
nand U23883 (N_23883,N_21741,N_21710);
nor U23884 (N_23884,N_22418,N_21063);
and U23885 (N_23885,N_20228,N_20599);
nand U23886 (N_23886,N_20113,N_20287);
nor U23887 (N_23887,N_20147,N_20409);
nor U23888 (N_23888,N_20622,N_20618);
or U23889 (N_23889,N_20218,N_20547);
xnor U23890 (N_23890,N_20960,N_20181);
nor U23891 (N_23891,N_20725,N_20285);
xor U23892 (N_23892,N_21214,N_20002);
xor U23893 (N_23893,N_20564,N_20732);
xnor U23894 (N_23894,N_20328,N_21926);
nand U23895 (N_23895,N_20742,N_21277);
nand U23896 (N_23896,N_22334,N_21147);
and U23897 (N_23897,N_21689,N_21941);
nand U23898 (N_23898,N_20832,N_20741);
and U23899 (N_23899,N_20628,N_20401);
xnor U23900 (N_23900,N_21738,N_20717);
xor U23901 (N_23901,N_21617,N_20142);
xor U23902 (N_23902,N_22414,N_20160);
and U23903 (N_23903,N_21001,N_20600);
nand U23904 (N_23904,N_21184,N_20936);
nand U23905 (N_23905,N_22061,N_20189);
or U23906 (N_23906,N_20785,N_20193);
and U23907 (N_23907,N_22322,N_20617);
and U23908 (N_23908,N_22190,N_21368);
nand U23909 (N_23909,N_22306,N_21511);
xor U23910 (N_23910,N_22301,N_20220);
xnor U23911 (N_23911,N_20434,N_22094);
xor U23912 (N_23912,N_20917,N_21929);
or U23913 (N_23913,N_21764,N_21445);
or U23914 (N_23914,N_21734,N_21534);
xor U23915 (N_23915,N_21280,N_20811);
and U23916 (N_23916,N_20501,N_21719);
nor U23917 (N_23917,N_20327,N_20525);
nor U23918 (N_23918,N_21651,N_22153);
nor U23919 (N_23919,N_21452,N_21859);
nor U23920 (N_23920,N_20376,N_20721);
nand U23921 (N_23921,N_21851,N_20239);
nor U23922 (N_23922,N_20645,N_20337);
or U23923 (N_23923,N_20743,N_22471);
nand U23924 (N_23924,N_22430,N_21588);
and U23925 (N_23925,N_21037,N_21777);
xor U23926 (N_23926,N_22373,N_22170);
nand U23927 (N_23927,N_21011,N_21705);
or U23928 (N_23928,N_21671,N_20855);
and U23929 (N_23929,N_22092,N_20173);
nand U23930 (N_23930,N_21804,N_20933);
nand U23931 (N_23931,N_21300,N_20882);
or U23932 (N_23932,N_20001,N_20645);
nand U23933 (N_23933,N_21509,N_21987);
and U23934 (N_23934,N_20948,N_20371);
nor U23935 (N_23935,N_21637,N_21383);
nand U23936 (N_23936,N_20174,N_21190);
xor U23937 (N_23937,N_20749,N_22060);
or U23938 (N_23938,N_21254,N_21728);
xnor U23939 (N_23939,N_21264,N_20154);
nand U23940 (N_23940,N_22304,N_20503);
nor U23941 (N_23941,N_20134,N_21135);
or U23942 (N_23942,N_21661,N_22177);
and U23943 (N_23943,N_21978,N_20495);
xnor U23944 (N_23944,N_20989,N_22129);
and U23945 (N_23945,N_22122,N_21966);
or U23946 (N_23946,N_20781,N_20682);
xor U23947 (N_23947,N_20580,N_20980);
nor U23948 (N_23948,N_21630,N_20133);
nand U23949 (N_23949,N_20012,N_21432);
and U23950 (N_23950,N_20677,N_20601);
nor U23951 (N_23951,N_20692,N_22016);
and U23952 (N_23952,N_22399,N_22255);
xor U23953 (N_23953,N_21624,N_21841);
nand U23954 (N_23954,N_20021,N_22098);
or U23955 (N_23955,N_22393,N_22468);
nor U23956 (N_23956,N_21674,N_22390);
nor U23957 (N_23957,N_22051,N_21729);
nor U23958 (N_23958,N_22347,N_20943);
or U23959 (N_23959,N_21753,N_22185);
nand U23960 (N_23960,N_21282,N_21302);
nand U23961 (N_23961,N_21549,N_22251);
or U23962 (N_23962,N_21212,N_21994);
and U23963 (N_23963,N_20554,N_20052);
nand U23964 (N_23964,N_22404,N_21748);
xnor U23965 (N_23965,N_21420,N_20869);
nand U23966 (N_23966,N_20190,N_22468);
nor U23967 (N_23967,N_21039,N_22305);
xnor U23968 (N_23968,N_21380,N_21927);
nor U23969 (N_23969,N_21810,N_20011);
xor U23970 (N_23970,N_21757,N_20643);
nand U23971 (N_23971,N_21976,N_20722);
and U23972 (N_23972,N_22018,N_21283);
nor U23973 (N_23973,N_20706,N_20985);
nor U23974 (N_23974,N_20699,N_20724);
nand U23975 (N_23975,N_20736,N_21810);
and U23976 (N_23976,N_22013,N_21885);
xor U23977 (N_23977,N_20295,N_20138);
and U23978 (N_23978,N_22301,N_20654);
xnor U23979 (N_23979,N_20192,N_21242);
xor U23980 (N_23980,N_20031,N_20868);
nor U23981 (N_23981,N_20351,N_21046);
nor U23982 (N_23982,N_22476,N_21006);
xor U23983 (N_23983,N_21594,N_21069);
nor U23984 (N_23984,N_21080,N_21415);
and U23985 (N_23985,N_21326,N_20858);
or U23986 (N_23986,N_21147,N_22266);
nor U23987 (N_23987,N_21916,N_20509);
nor U23988 (N_23988,N_20543,N_22142);
nor U23989 (N_23989,N_22028,N_20800);
or U23990 (N_23990,N_21603,N_21525);
and U23991 (N_23991,N_20174,N_22231);
nand U23992 (N_23992,N_22160,N_21028);
or U23993 (N_23993,N_22498,N_21077);
xor U23994 (N_23994,N_21755,N_20236);
nor U23995 (N_23995,N_22336,N_21827);
nor U23996 (N_23996,N_22452,N_22353);
or U23997 (N_23997,N_21743,N_22105);
and U23998 (N_23998,N_21062,N_20851);
or U23999 (N_23999,N_21646,N_21616);
or U24000 (N_24000,N_22159,N_20374);
nand U24001 (N_24001,N_21257,N_20796);
nor U24002 (N_24002,N_21275,N_21167);
nand U24003 (N_24003,N_21205,N_20115);
xnor U24004 (N_24004,N_20354,N_22112);
nand U24005 (N_24005,N_20862,N_20023);
xnor U24006 (N_24006,N_21283,N_21832);
and U24007 (N_24007,N_21214,N_20772);
and U24008 (N_24008,N_20889,N_22225);
xor U24009 (N_24009,N_21501,N_20857);
and U24010 (N_24010,N_22321,N_21162);
xnor U24011 (N_24011,N_21022,N_22345);
xor U24012 (N_24012,N_21700,N_21376);
nor U24013 (N_24013,N_21803,N_21105);
nand U24014 (N_24014,N_22043,N_22457);
nor U24015 (N_24015,N_22369,N_21589);
and U24016 (N_24016,N_21884,N_20698);
xnor U24017 (N_24017,N_20885,N_21495);
xnor U24018 (N_24018,N_20920,N_22052);
xnor U24019 (N_24019,N_21709,N_21298);
and U24020 (N_24020,N_21036,N_22018);
nand U24021 (N_24021,N_21347,N_20675);
nor U24022 (N_24022,N_20994,N_20219);
nand U24023 (N_24023,N_20583,N_21521);
nand U24024 (N_24024,N_21439,N_22455);
nor U24025 (N_24025,N_21386,N_21814);
and U24026 (N_24026,N_22448,N_21839);
nand U24027 (N_24027,N_20432,N_21213);
or U24028 (N_24028,N_21148,N_22309);
or U24029 (N_24029,N_21461,N_22346);
nand U24030 (N_24030,N_20628,N_20073);
and U24031 (N_24031,N_22191,N_21631);
nor U24032 (N_24032,N_20899,N_21291);
or U24033 (N_24033,N_21758,N_20042);
nor U24034 (N_24034,N_21255,N_22174);
xnor U24035 (N_24035,N_22325,N_21214);
and U24036 (N_24036,N_21762,N_20548);
nor U24037 (N_24037,N_21033,N_21168);
nand U24038 (N_24038,N_20364,N_21304);
and U24039 (N_24039,N_20139,N_22113);
nor U24040 (N_24040,N_20304,N_21904);
and U24041 (N_24041,N_22176,N_21956);
nor U24042 (N_24042,N_22285,N_21057);
xor U24043 (N_24043,N_21095,N_20502);
nor U24044 (N_24044,N_21475,N_21448);
or U24045 (N_24045,N_20001,N_21816);
or U24046 (N_24046,N_22121,N_21281);
and U24047 (N_24047,N_20441,N_22125);
or U24048 (N_24048,N_20850,N_21297);
and U24049 (N_24049,N_22106,N_20188);
or U24050 (N_24050,N_21243,N_20714);
or U24051 (N_24051,N_20021,N_20263);
and U24052 (N_24052,N_20821,N_22298);
and U24053 (N_24053,N_20602,N_21989);
xor U24054 (N_24054,N_20069,N_20860);
and U24055 (N_24055,N_20000,N_21700);
xnor U24056 (N_24056,N_20047,N_20719);
or U24057 (N_24057,N_22186,N_22005);
nor U24058 (N_24058,N_21892,N_22144);
and U24059 (N_24059,N_20267,N_22148);
nand U24060 (N_24060,N_20925,N_21354);
and U24061 (N_24061,N_20945,N_20295);
and U24062 (N_24062,N_22019,N_20206);
and U24063 (N_24063,N_21884,N_21873);
or U24064 (N_24064,N_21645,N_21466);
nor U24065 (N_24065,N_20520,N_22321);
nand U24066 (N_24066,N_22361,N_20319);
nand U24067 (N_24067,N_21230,N_22123);
nor U24068 (N_24068,N_20312,N_22114);
nand U24069 (N_24069,N_21996,N_20171);
nor U24070 (N_24070,N_20184,N_20649);
nand U24071 (N_24071,N_21826,N_20517);
xnor U24072 (N_24072,N_21752,N_22382);
nand U24073 (N_24073,N_20280,N_21747);
or U24074 (N_24074,N_21992,N_21920);
or U24075 (N_24075,N_20654,N_21920);
xnor U24076 (N_24076,N_22473,N_20461);
xor U24077 (N_24077,N_21867,N_22137);
nand U24078 (N_24078,N_21216,N_20783);
and U24079 (N_24079,N_20301,N_21968);
nand U24080 (N_24080,N_21897,N_20392);
xnor U24081 (N_24081,N_20831,N_21093);
xor U24082 (N_24082,N_20536,N_21996);
xor U24083 (N_24083,N_21731,N_22242);
or U24084 (N_24084,N_21268,N_20055);
nor U24085 (N_24085,N_20108,N_20299);
nand U24086 (N_24086,N_21953,N_20865);
nor U24087 (N_24087,N_21715,N_21949);
and U24088 (N_24088,N_20081,N_21811);
or U24089 (N_24089,N_20367,N_21529);
xnor U24090 (N_24090,N_20866,N_20368);
nor U24091 (N_24091,N_20026,N_22373);
xnor U24092 (N_24092,N_21951,N_20574);
nand U24093 (N_24093,N_20944,N_22486);
and U24094 (N_24094,N_22004,N_20669);
xnor U24095 (N_24095,N_21200,N_22343);
or U24096 (N_24096,N_20239,N_21829);
xor U24097 (N_24097,N_20483,N_20413);
nor U24098 (N_24098,N_21601,N_20397);
and U24099 (N_24099,N_21069,N_21331);
and U24100 (N_24100,N_20522,N_22139);
nand U24101 (N_24101,N_20051,N_21293);
xnor U24102 (N_24102,N_21296,N_22010);
nand U24103 (N_24103,N_21550,N_20846);
or U24104 (N_24104,N_20305,N_20810);
xnor U24105 (N_24105,N_22494,N_22224);
xor U24106 (N_24106,N_21834,N_20106);
xor U24107 (N_24107,N_20455,N_21033);
and U24108 (N_24108,N_20311,N_21561);
or U24109 (N_24109,N_20030,N_22261);
nor U24110 (N_24110,N_21895,N_20257);
or U24111 (N_24111,N_21651,N_20106);
xnor U24112 (N_24112,N_21501,N_22450);
or U24113 (N_24113,N_22051,N_21499);
and U24114 (N_24114,N_22190,N_22085);
xor U24115 (N_24115,N_20940,N_21459);
and U24116 (N_24116,N_21095,N_20349);
nor U24117 (N_24117,N_20954,N_21665);
or U24118 (N_24118,N_21432,N_21506);
nand U24119 (N_24119,N_20627,N_21345);
nor U24120 (N_24120,N_21999,N_20961);
or U24121 (N_24121,N_20274,N_20452);
and U24122 (N_24122,N_20371,N_22373);
xnor U24123 (N_24123,N_22471,N_20034);
xnor U24124 (N_24124,N_21440,N_22164);
nand U24125 (N_24125,N_22447,N_20409);
xor U24126 (N_24126,N_21885,N_22179);
or U24127 (N_24127,N_22033,N_20286);
or U24128 (N_24128,N_20600,N_20592);
nand U24129 (N_24129,N_20208,N_21932);
and U24130 (N_24130,N_20886,N_22296);
xor U24131 (N_24131,N_21591,N_20675);
xor U24132 (N_24132,N_20318,N_20387);
xor U24133 (N_24133,N_20460,N_20475);
nor U24134 (N_24134,N_20517,N_21580);
nor U24135 (N_24135,N_20937,N_21930);
or U24136 (N_24136,N_21872,N_21750);
and U24137 (N_24137,N_20795,N_22216);
or U24138 (N_24138,N_22204,N_22176);
nor U24139 (N_24139,N_22190,N_20990);
or U24140 (N_24140,N_21024,N_20400);
or U24141 (N_24141,N_21791,N_21266);
nand U24142 (N_24142,N_21868,N_21434);
nand U24143 (N_24143,N_22103,N_21120);
or U24144 (N_24144,N_21547,N_20088);
nor U24145 (N_24145,N_20542,N_21980);
nand U24146 (N_24146,N_21520,N_21403);
nand U24147 (N_24147,N_20686,N_20755);
nand U24148 (N_24148,N_20726,N_21574);
nor U24149 (N_24149,N_20226,N_22074);
and U24150 (N_24150,N_21400,N_20795);
xor U24151 (N_24151,N_21466,N_21680);
or U24152 (N_24152,N_22408,N_20959);
xnor U24153 (N_24153,N_20884,N_20317);
and U24154 (N_24154,N_20447,N_21741);
and U24155 (N_24155,N_21410,N_20362);
xor U24156 (N_24156,N_20615,N_21761);
or U24157 (N_24157,N_20887,N_21611);
nand U24158 (N_24158,N_20749,N_21246);
and U24159 (N_24159,N_20227,N_21455);
nand U24160 (N_24160,N_21378,N_21092);
nand U24161 (N_24161,N_20056,N_20468);
nor U24162 (N_24162,N_21128,N_20579);
or U24163 (N_24163,N_22373,N_20568);
or U24164 (N_24164,N_20374,N_20895);
or U24165 (N_24165,N_20666,N_20216);
xnor U24166 (N_24166,N_21646,N_21499);
xor U24167 (N_24167,N_21452,N_20225);
or U24168 (N_24168,N_22191,N_21305);
nor U24169 (N_24169,N_21157,N_20471);
xnor U24170 (N_24170,N_21001,N_21864);
and U24171 (N_24171,N_20710,N_20684);
xor U24172 (N_24172,N_20036,N_21168);
or U24173 (N_24173,N_21625,N_21518);
nand U24174 (N_24174,N_20890,N_22003);
xnor U24175 (N_24175,N_21342,N_22003);
nor U24176 (N_24176,N_21246,N_20523);
nor U24177 (N_24177,N_20121,N_22151);
xor U24178 (N_24178,N_20263,N_20609);
nand U24179 (N_24179,N_22446,N_20394);
or U24180 (N_24180,N_20842,N_20290);
nand U24181 (N_24181,N_22053,N_21358);
or U24182 (N_24182,N_22108,N_22128);
or U24183 (N_24183,N_21922,N_20861);
nand U24184 (N_24184,N_20625,N_20793);
nor U24185 (N_24185,N_21342,N_21038);
or U24186 (N_24186,N_20750,N_21740);
xnor U24187 (N_24187,N_22071,N_20577);
xnor U24188 (N_24188,N_21478,N_20139);
nor U24189 (N_24189,N_21996,N_21241);
xor U24190 (N_24190,N_22124,N_20734);
nor U24191 (N_24191,N_20276,N_21361);
and U24192 (N_24192,N_21120,N_21220);
and U24193 (N_24193,N_20661,N_20786);
nor U24194 (N_24194,N_20039,N_22354);
nor U24195 (N_24195,N_21363,N_22181);
nand U24196 (N_24196,N_22358,N_21236);
or U24197 (N_24197,N_21620,N_22364);
xnor U24198 (N_24198,N_21080,N_21251);
and U24199 (N_24199,N_22001,N_20059);
and U24200 (N_24200,N_20177,N_22404);
and U24201 (N_24201,N_22087,N_21402);
nor U24202 (N_24202,N_20388,N_20985);
or U24203 (N_24203,N_21460,N_22251);
nand U24204 (N_24204,N_21375,N_22217);
nor U24205 (N_24205,N_22132,N_20696);
or U24206 (N_24206,N_20253,N_20456);
nand U24207 (N_24207,N_21082,N_20495);
xnor U24208 (N_24208,N_20274,N_21231);
nand U24209 (N_24209,N_22013,N_21299);
or U24210 (N_24210,N_20191,N_22465);
or U24211 (N_24211,N_21933,N_22410);
xnor U24212 (N_24212,N_21749,N_22451);
nand U24213 (N_24213,N_21789,N_21921);
xnor U24214 (N_24214,N_21919,N_21302);
nor U24215 (N_24215,N_22005,N_22366);
and U24216 (N_24216,N_20860,N_21578);
xnor U24217 (N_24217,N_21499,N_22460);
nand U24218 (N_24218,N_22350,N_20415);
or U24219 (N_24219,N_21616,N_20439);
and U24220 (N_24220,N_20322,N_22090);
nor U24221 (N_24221,N_20904,N_22388);
or U24222 (N_24222,N_22242,N_21465);
or U24223 (N_24223,N_22175,N_22294);
nor U24224 (N_24224,N_20841,N_21148);
nor U24225 (N_24225,N_20079,N_21551);
nand U24226 (N_24226,N_21212,N_20793);
or U24227 (N_24227,N_22417,N_20687);
and U24228 (N_24228,N_22006,N_20472);
nor U24229 (N_24229,N_20674,N_20761);
and U24230 (N_24230,N_21664,N_20234);
nor U24231 (N_24231,N_20965,N_20225);
xor U24232 (N_24232,N_20910,N_20264);
nand U24233 (N_24233,N_20741,N_20715);
nor U24234 (N_24234,N_22037,N_20137);
and U24235 (N_24235,N_21803,N_20569);
nand U24236 (N_24236,N_21864,N_20164);
nand U24237 (N_24237,N_22275,N_20780);
or U24238 (N_24238,N_20062,N_21723);
nor U24239 (N_24239,N_20309,N_20474);
or U24240 (N_24240,N_21554,N_21680);
and U24241 (N_24241,N_20917,N_20858);
nor U24242 (N_24242,N_20767,N_21185);
or U24243 (N_24243,N_21203,N_22357);
and U24244 (N_24244,N_22264,N_21405);
or U24245 (N_24245,N_21275,N_20834);
nor U24246 (N_24246,N_22293,N_22299);
xor U24247 (N_24247,N_21986,N_20316);
nand U24248 (N_24248,N_20421,N_22325);
and U24249 (N_24249,N_21879,N_20383);
xnor U24250 (N_24250,N_21176,N_21977);
xor U24251 (N_24251,N_21588,N_22343);
xor U24252 (N_24252,N_22186,N_21367);
nor U24253 (N_24253,N_22039,N_22443);
nand U24254 (N_24254,N_21241,N_22075);
and U24255 (N_24255,N_22325,N_21401);
and U24256 (N_24256,N_21602,N_22289);
and U24257 (N_24257,N_21341,N_20155);
xor U24258 (N_24258,N_21888,N_20465);
and U24259 (N_24259,N_21564,N_20314);
nand U24260 (N_24260,N_21861,N_21780);
and U24261 (N_24261,N_21717,N_21375);
and U24262 (N_24262,N_21466,N_21485);
or U24263 (N_24263,N_20783,N_20233);
or U24264 (N_24264,N_20749,N_20807);
or U24265 (N_24265,N_21046,N_21654);
nand U24266 (N_24266,N_20368,N_20196);
nand U24267 (N_24267,N_20385,N_22275);
or U24268 (N_24268,N_20252,N_21722);
or U24269 (N_24269,N_21536,N_21125);
xnor U24270 (N_24270,N_20023,N_20737);
xor U24271 (N_24271,N_20065,N_21713);
nand U24272 (N_24272,N_20738,N_20302);
xor U24273 (N_24273,N_21179,N_21479);
or U24274 (N_24274,N_21838,N_21476);
nor U24275 (N_24275,N_21670,N_20444);
nor U24276 (N_24276,N_22201,N_21374);
xor U24277 (N_24277,N_21937,N_20414);
xor U24278 (N_24278,N_21248,N_22373);
and U24279 (N_24279,N_21223,N_20995);
xor U24280 (N_24280,N_21695,N_21783);
xor U24281 (N_24281,N_21938,N_20813);
nand U24282 (N_24282,N_20723,N_20579);
nor U24283 (N_24283,N_20510,N_21582);
nor U24284 (N_24284,N_20729,N_22242);
xnor U24285 (N_24285,N_21582,N_20642);
xnor U24286 (N_24286,N_20759,N_21404);
and U24287 (N_24287,N_20085,N_20138);
nand U24288 (N_24288,N_20058,N_21544);
nand U24289 (N_24289,N_20250,N_20162);
nand U24290 (N_24290,N_22069,N_20697);
or U24291 (N_24291,N_20371,N_22089);
nand U24292 (N_24292,N_22166,N_20264);
nor U24293 (N_24293,N_20116,N_20326);
xor U24294 (N_24294,N_20435,N_20623);
nor U24295 (N_24295,N_21600,N_20806);
nand U24296 (N_24296,N_22286,N_20970);
or U24297 (N_24297,N_22128,N_21715);
nor U24298 (N_24298,N_21310,N_20028);
or U24299 (N_24299,N_21403,N_20593);
nor U24300 (N_24300,N_21965,N_20780);
or U24301 (N_24301,N_20280,N_20598);
nor U24302 (N_24302,N_22247,N_20515);
and U24303 (N_24303,N_20772,N_21612);
xnor U24304 (N_24304,N_21968,N_21260);
nor U24305 (N_24305,N_22288,N_22491);
or U24306 (N_24306,N_21526,N_21833);
or U24307 (N_24307,N_21812,N_21004);
and U24308 (N_24308,N_20782,N_22375);
xnor U24309 (N_24309,N_22495,N_22228);
and U24310 (N_24310,N_22058,N_22402);
xnor U24311 (N_24311,N_21505,N_21467);
xor U24312 (N_24312,N_20114,N_21669);
nor U24313 (N_24313,N_21361,N_22106);
nand U24314 (N_24314,N_21423,N_21320);
xor U24315 (N_24315,N_20902,N_22357);
or U24316 (N_24316,N_21853,N_21924);
nand U24317 (N_24317,N_20375,N_20750);
nor U24318 (N_24318,N_20105,N_20479);
nand U24319 (N_24319,N_20333,N_21350);
and U24320 (N_24320,N_21750,N_21370);
nand U24321 (N_24321,N_22167,N_21479);
and U24322 (N_24322,N_20570,N_21669);
and U24323 (N_24323,N_21260,N_21472);
and U24324 (N_24324,N_20606,N_20481);
or U24325 (N_24325,N_22361,N_21639);
xor U24326 (N_24326,N_22116,N_20570);
and U24327 (N_24327,N_21745,N_20044);
and U24328 (N_24328,N_20853,N_20075);
and U24329 (N_24329,N_20120,N_22373);
or U24330 (N_24330,N_20668,N_22161);
nand U24331 (N_24331,N_21580,N_22423);
nor U24332 (N_24332,N_21438,N_20441);
or U24333 (N_24333,N_22403,N_22241);
xor U24334 (N_24334,N_21289,N_21992);
nand U24335 (N_24335,N_21529,N_20818);
or U24336 (N_24336,N_20766,N_20237);
or U24337 (N_24337,N_20707,N_20916);
nor U24338 (N_24338,N_22116,N_20608);
nand U24339 (N_24339,N_20286,N_21474);
nand U24340 (N_24340,N_22333,N_20823);
nor U24341 (N_24341,N_21784,N_21230);
nand U24342 (N_24342,N_20120,N_21072);
and U24343 (N_24343,N_20049,N_20703);
nor U24344 (N_24344,N_21944,N_20827);
xor U24345 (N_24345,N_20295,N_20053);
xor U24346 (N_24346,N_21483,N_22461);
or U24347 (N_24347,N_20846,N_20709);
nor U24348 (N_24348,N_20381,N_20184);
and U24349 (N_24349,N_20135,N_22269);
nand U24350 (N_24350,N_20005,N_20389);
xnor U24351 (N_24351,N_21201,N_22372);
xnor U24352 (N_24352,N_20226,N_20507);
or U24353 (N_24353,N_22374,N_20400);
nor U24354 (N_24354,N_20345,N_21555);
or U24355 (N_24355,N_20613,N_21135);
nor U24356 (N_24356,N_22307,N_21004);
or U24357 (N_24357,N_21287,N_22217);
nor U24358 (N_24358,N_20728,N_20523);
and U24359 (N_24359,N_20887,N_20731);
nor U24360 (N_24360,N_22124,N_22222);
xnor U24361 (N_24361,N_21511,N_20922);
xnor U24362 (N_24362,N_21852,N_20120);
xor U24363 (N_24363,N_21191,N_21416);
nor U24364 (N_24364,N_20515,N_20490);
nor U24365 (N_24365,N_22116,N_21507);
and U24366 (N_24366,N_21451,N_21606);
and U24367 (N_24367,N_22233,N_21246);
xnor U24368 (N_24368,N_20854,N_20698);
and U24369 (N_24369,N_21898,N_20753);
nand U24370 (N_24370,N_21765,N_20272);
nor U24371 (N_24371,N_22393,N_22442);
nor U24372 (N_24372,N_21005,N_21963);
and U24373 (N_24373,N_20330,N_22276);
and U24374 (N_24374,N_21162,N_21775);
and U24375 (N_24375,N_21508,N_20801);
nand U24376 (N_24376,N_21511,N_20242);
and U24377 (N_24377,N_21315,N_20911);
xnor U24378 (N_24378,N_20683,N_20622);
or U24379 (N_24379,N_21792,N_20426);
and U24380 (N_24380,N_21608,N_21543);
nand U24381 (N_24381,N_20821,N_21304);
nand U24382 (N_24382,N_22410,N_21227);
and U24383 (N_24383,N_22027,N_20479);
and U24384 (N_24384,N_20404,N_22027);
nand U24385 (N_24385,N_20386,N_22460);
xnor U24386 (N_24386,N_20529,N_21738);
or U24387 (N_24387,N_20033,N_21008);
or U24388 (N_24388,N_21945,N_22435);
or U24389 (N_24389,N_21907,N_21924);
or U24390 (N_24390,N_21494,N_22067);
xor U24391 (N_24391,N_21697,N_22152);
nand U24392 (N_24392,N_20504,N_20991);
or U24393 (N_24393,N_20734,N_21170);
xor U24394 (N_24394,N_20594,N_21034);
nor U24395 (N_24395,N_21903,N_21333);
nor U24396 (N_24396,N_21752,N_22483);
nand U24397 (N_24397,N_21843,N_20395);
nand U24398 (N_24398,N_20056,N_20785);
nand U24399 (N_24399,N_21482,N_21085);
nor U24400 (N_24400,N_22412,N_20620);
xor U24401 (N_24401,N_20745,N_21415);
and U24402 (N_24402,N_21722,N_22447);
xor U24403 (N_24403,N_22305,N_22443);
and U24404 (N_24404,N_20864,N_21464);
nor U24405 (N_24405,N_20723,N_21988);
nand U24406 (N_24406,N_21367,N_21728);
or U24407 (N_24407,N_20715,N_21100);
or U24408 (N_24408,N_20344,N_20472);
nor U24409 (N_24409,N_20911,N_21476);
or U24410 (N_24410,N_22153,N_21486);
or U24411 (N_24411,N_21335,N_20711);
and U24412 (N_24412,N_21353,N_20044);
nor U24413 (N_24413,N_20722,N_21795);
nor U24414 (N_24414,N_20911,N_21488);
nand U24415 (N_24415,N_20595,N_21955);
or U24416 (N_24416,N_20560,N_22130);
nand U24417 (N_24417,N_22146,N_20493);
nor U24418 (N_24418,N_20794,N_21058);
and U24419 (N_24419,N_20268,N_20438);
nor U24420 (N_24420,N_21352,N_22323);
nor U24421 (N_24421,N_22233,N_20522);
nand U24422 (N_24422,N_21054,N_22234);
xnor U24423 (N_24423,N_20994,N_20917);
or U24424 (N_24424,N_20609,N_21917);
or U24425 (N_24425,N_21409,N_20882);
xor U24426 (N_24426,N_20732,N_22344);
nand U24427 (N_24427,N_21220,N_21635);
or U24428 (N_24428,N_22195,N_20509);
nor U24429 (N_24429,N_20685,N_21287);
nand U24430 (N_24430,N_20755,N_22073);
xnor U24431 (N_24431,N_20414,N_20937);
and U24432 (N_24432,N_22235,N_20617);
and U24433 (N_24433,N_21357,N_20397);
xor U24434 (N_24434,N_21132,N_22445);
xor U24435 (N_24435,N_22276,N_20176);
nand U24436 (N_24436,N_22155,N_21573);
nor U24437 (N_24437,N_21885,N_20561);
and U24438 (N_24438,N_21773,N_22134);
or U24439 (N_24439,N_21954,N_21295);
xor U24440 (N_24440,N_22076,N_21568);
nor U24441 (N_24441,N_20785,N_20673);
xor U24442 (N_24442,N_20541,N_22244);
or U24443 (N_24443,N_20071,N_21705);
and U24444 (N_24444,N_21717,N_22153);
nor U24445 (N_24445,N_22348,N_20418);
or U24446 (N_24446,N_21621,N_20173);
nor U24447 (N_24447,N_21496,N_21010);
and U24448 (N_24448,N_21670,N_21065);
or U24449 (N_24449,N_21845,N_21503);
and U24450 (N_24450,N_22350,N_21443);
xor U24451 (N_24451,N_22293,N_20467);
xor U24452 (N_24452,N_20599,N_22306);
or U24453 (N_24453,N_21944,N_21161);
and U24454 (N_24454,N_21998,N_22257);
or U24455 (N_24455,N_20757,N_20384);
nor U24456 (N_24456,N_22379,N_20159);
nand U24457 (N_24457,N_20324,N_20784);
xor U24458 (N_24458,N_21929,N_21453);
xnor U24459 (N_24459,N_21268,N_22113);
nor U24460 (N_24460,N_21814,N_21133);
nand U24461 (N_24461,N_21276,N_20802);
nor U24462 (N_24462,N_21793,N_20543);
or U24463 (N_24463,N_21931,N_20097);
nor U24464 (N_24464,N_22400,N_20472);
nor U24465 (N_24465,N_20632,N_20307);
nand U24466 (N_24466,N_20357,N_20297);
or U24467 (N_24467,N_21246,N_21142);
or U24468 (N_24468,N_21021,N_21310);
or U24469 (N_24469,N_20466,N_20583);
nand U24470 (N_24470,N_20470,N_21198);
nor U24471 (N_24471,N_20612,N_20687);
or U24472 (N_24472,N_20352,N_21428);
and U24473 (N_24473,N_20967,N_22037);
xor U24474 (N_24474,N_20829,N_20115);
xnor U24475 (N_24475,N_20231,N_22334);
and U24476 (N_24476,N_20851,N_21777);
nor U24477 (N_24477,N_22303,N_20205);
and U24478 (N_24478,N_22214,N_20433);
xnor U24479 (N_24479,N_21545,N_21889);
or U24480 (N_24480,N_20628,N_21781);
and U24481 (N_24481,N_21215,N_20701);
xor U24482 (N_24482,N_21740,N_21953);
nor U24483 (N_24483,N_20418,N_21832);
nor U24484 (N_24484,N_21405,N_21459);
xnor U24485 (N_24485,N_20906,N_20681);
or U24486 (N_24486,N_20236,N_21705);
and U24487 (N_24487,N_22015,N_21225);
nand U24488 (N_24488,N_21524,N_21420);
or U24489 (N_24489,N_20442,N_21879);
xor U24490 (N_24490,N_22462,N_21395);
xor U24491 (N_24491,N_20982,N_22158);
xnor U24492 (N_24492,N_20212,N_20275);
and U24493 (N_24493,N_20181,N_20223);
and U24494 (N_24494,N_21359,N_21767);
nand U24495 (N_24495,N_21454,N_20359);
and U24496 (N_24496,N_20230,N_21492);
or U24497 (N_24497,N_21863,N_20683);
nor U24498 (N_24498,N_21621,N_20289);
or U24499 (N_24499,N_21212,N_21582);
or U24500 (N_24500,N_20453,N_22495);
and U24501 (N_24501,N_20268,N_20033);
or U24502 (N_24502,N_20940,N_22026);
nor U24503 (N_24503,N_22401,N_21537);
nor U24504 (N_24504,N_20560,N_20166);
nand U24505 (N_24505,N_21887,N_20109);
nand U24506 (N_24506,N_20436,N_21678);
xor U24507 (N_24507,N_21810,N_20404);
nand U24508 (N_24508,N_21705,N_21972);
or U24509 (N_24509,N_21383,N_21374);
nor U24510 (N_24510,N_20525,N_20161);
and U24511 (N_24511,N_21133,N_20610);
xnor U24512 (N_24512,N_22381,N_21526);
nand U24513 (N_24513,N_20770,N_21421);
nor U24514 (N_24514,N_20028,N_21674);
nand U24515 (N_24515,N_21193,N_21561);
and U24516 (N_24516,N_20083,N_22274);
and U24517 (N_24517,N_20374,N_21282);
nor U24518 (N_24518,N_20051,N_20738);
or U24519 (N_24519,N_21422,N_20699);
xnor U24520 (N_24520,N_21174,N_20542);
nor U24521 (N_24521,N_22176,N_20128);
and U24522 (N_24522,N_21289,N_20556);
nand U24523 (N_24523,N_20265,N_20338);
and U24524 (N_24524,N_20420,N_21750);
nand U24525 (N_24525,N_20826,N_21716);
nand U24526 (N_24526,N_22062,N_20571);
nand U24527 (N_24527,N_20622,N_22274);
or U24528 (N_24528,N_20546,N_22435);
or U24529 (N_24529,N_21145,N_21886);
nor U24530 (N_24530,N_22064,N_21040);
or U24531 (N_24531,N_21797,N_20401);
nand U24532 (N_24532,N_20747,N_20410);
or U24533 (N_24533,N_22337,N_22296);
nand U24534 (N_24534,N_21127,N_21192);
nor U24535 (N_24535,N_20598,N_21565);
nor U24536 (N_24536,N_20062,N_20055);
and U24537 (N_24537,N_20485,N_21342);
xnor U24538 (N_24538,N_20709,N_22023);
and U24539 (N_24539,N_22046,N_21186);
and U24540 (N_24540,N_22357,N_21182);
nand U24541 (N_24541,N_21762,N_22358);
and U24542 (N_24542,N_22133,N_20495);
and U24543 (N_24543,N_21584,N_20042);
xnor U24544 (N_24544,N_21620,N_20541);
or U24545 (N_24545,N_20030,N_21369);
or U24546 (N_24546,N_21645,N_20732);
nor U24547 (N_24547,N_21262,N_20259);
nand U24548 (N_24548,N_20716,N_21819);
nor U24549 (N_24549,N_21905,N_22408);
nor U24550 (N_24550,N_21956,N_20236);
or U24551 (N_24551,N_21177,N_21951);
or U24552 (N_24552,N_20907,N_21989);
and U24553 (N_24553,N_21390,N_20548);
nand U24554 (N_24554,N_22228,N_22374);
nand U24555 (N_24555,N_21734,N_21979);
and U24556 (N_24556,N_22417,N_21081);
nand U24557 (N_24557,N_20597,N_21810);
or U24558 (N_24558,N_20334,N_22034);
nor U24559 (N_24559,N_20141,N_20347);
xor U24560 (N_24560,N_21158,N_20979);
or U24561 (N_24561,N_20506,N_21390);
nand U24562 (N_24562,N_21802,N_20222);
or U24563 (N_24563,N_20824,N_22019);
and U24564 (N_24564,N_20296,N_21486);
or U24565 (N_24565,N_21298,N_22339);
nor U24566 (N_24566,N_20155,N_22430);
and U24567 (N_24567,N_20570,N_21505);
xor U24568 (N_24568,N_20152,N_20343);
or U24569 (N_24569,N_20870,N_20684);
xnor U24570 (N_24570,N_22208,N_20311);
nor U24571 (N_24571,N_21886,N_21543);
nor U24572 (N_24572,N_21303,N_20096);
nand U24573 (N_24573,N_21140,N_21631);
and U24574 (N_24574,N_21902,N_22193);
and U24575 (N_24575,N_20639,N_22338);
xnor U24576 (N_24576,N_20487,N_20602);
or U24577 (N_24577,N_21490,N_20382);
and U24578 (N_24578,N_21405,N_20083);
nand U24579 (N_24579,N_20961,N_22219);
or U24580 (N_24580,N_21383,N_21468);
and U24581 (N_24581,N_20541,N_20734);
or U24582 (N_24582,N_22010,N_21437);
xnor U24583 (N_24583,N_22251,N_22056);
nor U24584 (N_24584,N_22311,N_20714);
nor U24585 (N_24585,N_20062,N_21271);
nor U24586 (N_24586,N_21102,N_21436);
nor U24587 (N_24587,N_20776,N_20658);
nor U24588 (N_24588,N_22330,N_22377);
and U24589 (N_24589,N_20646,N_21208);
and U24590 (N_24590,N_20230,N_22160);
nor U24591 (N_24591,N_21922,N_20263);
or U24592 (N_24592,N_22440,N_21952);
nor U24593 (N_24593,N_21619,N_20817);
nor U24594 (N_24594,N_20710,N_20821);
nor U24595 (N_24595,N_20037,N_21067);
and U24596 (N_24596,N_20656,N_20282);
nor U24597 (N_24597,N_21086,N_21570);
nand U24598 (N_24598,N_22046,N_22133);
xnor U24599 (N_24599,N_20475,N_21214);
and U24600 (N_24600,N_21102,N_21658);
nand U24601 (N_24601,N_21486,N_20771);
nand U24602 (N_24602,N_21081,N_22271);
and U24603 (N_24603,N_21217,N_20831);
or U24604 (N_24604,N_20045,N_22325);
and U24605 (N_24605,N_20542,N_20840);
or U24606 (N_24606,N_20845,N_21837);
xor U24607 (N_24607,N_20130,N_20542);
and U24608 (N_24608,N_20892,N_21229);
xor U24609 (N_24609,N_21643,N_20518);
xnor U24610 (N_24610,N_21869,N_20207);
nor U24611 (N_24611,N_22325,N_21056);
and U24612 (N_24612,N_22014,N_21964);
nand U24613 (N_24613,N_21005,N_20901);
nor U24614 (N_24614,N_20984,N_20612);
or U24615 (N_24615,N_21708,N_20096);
nor U24616 (N_24616,N_21849,N_20717);
or U24617 (N_24617,N_20471,N_22339);
nand U24618 (N_24618,N_22204,N_21985);
xnor U24619 (N_24619,N_21443,N_22221);
or U24620 (N_24620,N_21519,N_21863);
nor U24621 (N_24621,N_20355,N_21425);
or U24622 (N_24622,N_20025,N_21084);
nand U24623 (N_24623,N_20663,N_21473);
or U24624 (N_24624,N_21991,N_20000);
nor U24625 (N_24625,N_20717,N_20609);
nand U24626 (N_24626,N_21705,N_21549);
and U24627 (N_24627,N_21264,N_20473);
and U24628 (N_24628,N_22276,N_22470);
nor U24629 (N_24629,N_20353,N_20012);
nor U24630 (N_24630,N_20741,N_21888);
or U24631 (N_24631,N_21705,N_21178);
and U24632 (N_24632,N_20457,N_20030);
or U24633 (N_24633,N_21304,N_21549);
nand U24634 (N_24634,N_20715,N_21158);
and U24635 (N_24635,N_20409,N_22434);
and U24636 (N_24636,N_20486,N_21942);
and U24637 (N_24637,N_21668,N_20035);
xor U24638 (N_24638,N_20955,N_21092);
and U24639 (N_24639,N_22417,N_21854);
or U24640 (N_24640,N_20765,N_20598);
and U24641 (N_24641,N_22347,N_22288);
or U24642 (N_24642,N_22497,N_21347);
nand U24643 (N_24643,N_20916,N_20686);
nor U24644 (N_24644,N_20870,N_22398);
nand U24645 (N_24645,N_21332,N_20220);
nor U24646 (N_24646,N_20592,N_20079);
xnor U24647 (N_24647,N_20073,N_20483);
nor U24648 (N_24648,N_21253,N_21566);
and U24649 (N_24649,N_21011,N_22037);
and U24650 (N_24650,N_20103,N_20051);
or U24651 (N_24651,N_21977,N_22406);
and U24652 (N_24652,N_22230,N_21458);
xor U24653 (N_24653,N_20908,N_22172);
xnor U24654 (N_24654,N_21241,N_21345);
xor U24655 (N_24655,N_22053,N_22313);
nor U24656 (N_24656,N_21431,N_20235);
and U24657 (N_24657,N_21582,N_20942);
nor U24658 (N_24658,N_22293,N_21535);
nor U24659 (N_24659,N_22099,N_20958);
nand U24660 (N_24660,N_20238,N_20279);
nand U24661 (N_24661,N_22408,N_20745);
nor U24662 (N_24662,N_21687,N_22031);
xnor U24663 (N_24663,N_21508,N_20601);
and U24664 (N_24664,N_21562,N_20460);
or U24665 (N_24665,N_21811,N_20240);
or U24666 (N_24666,N_21613,N_21565);
nand U24667 (N_24667,N_21483,N_22140);
nand U24668 (N_24668,N_21053,N_22019);
nand U24669 (N_24669,N_22215,N_22143);
and U24670 (N_24670,N_21718,N_21699);
nand U24671 (N_24671,N_20740,N_22230);
or U24672 (N_24672,N_21416,N_20493);
nor U24673 (N_24673,N_21954,N_21373);
nand U24674 (N_24674,N_21352,N_22217);
nor U24675 (N_24675,N_21142,N_21833);
and U24676 (N_24676,N_21065,N_21944);
nor U24677 (N_24677,N_21712,N_21598);
or U24678 (N_24678,N_21130,N_20328);
and U24679 (N_24679,N_21869,N_21209);
nor U24680 (N_24680,N_21227,N_20855);
xor U24681 (N_24681,N_20377,N_22214);
nor U24682 (N_24682,N_22477,N_21568);
nor U24683 (N_24683,N_22142,N_21238);
nand U24684 (N_24684,N_20127,N_20225);
nand U24685 (N_24685,N_20012,N_20415);
or U24686 (N_24686,N_20838,N_21749);
and U24687 (N_24687,N_22092,N_21493);
nand U24688 (N_24688,N_20932,N_20859);
nand U24689 (N_24689,N_20882,N_20691);
nand U24690 (N_24690,N_21031,N_20767);
xnor U24691 (N_24691,N_21047,N_20303);
and U24692 (N_24692,N_20478,N_21746);
nand U24693 (N_24693,N_21637,N_20495);
nor U24694 (N_24694,N_21714,N_22122);
and U24695 (N_24695,N_20794,N_21170);
xnor U24696 (N_24696,N_20255,N_20027);
xnor U24697 (N_24697,N_22392,N_22162);
nor U24698 (N_24698,N_21212,N_20261);
nor U24699 (N_24699,N_21746,N_21900);
or U24700 (N_24700,N_22145,N_20731);
nand U24701 (N_24701,N_22020,N_21503);
nor U24702 (N_24702,N_22096,N_21224);
nand U24703 (N_24703,N_20012,N_20796);
or U24704 (N_24704,N_22008,N_21877);
and U24705 (N_24705,N_21667,N_22252);
nand U24706 (N_24706,N_21131,N_21149);
nor U24707 (N_24707,N_20502,N_21642);
and U24708 (N_24708,N_20892,N_21480);
nor U24709 (N_24709,N_21583,N_21856);
xnor U24710 (N_24710,N_21544,N_21188);
nor U24711 (N_24711,N_20104,N_20793);
xor U24712 (N_24712,N_20573,N_20399);
or U24713 (N_24713,N_20557,N_22157);
xor U24714 (N_24714,N_21445,N_20968);
nand U24715 (N_24715,N_22085,N_21160);
or U24716 (N_24716,N_21851,N_20967);
and U24717 (N_24717,N_21694,N_21736);
nand U24718 (N_24718,N_20148,N_21617);
xnor U24719 (N_24719,N_21669,N_22176);
or U24720 (N_24720,N_22035,N_20330);
xnor U24721 (N_24721,N_21097,N_21320);
xor U24722 (N_24722,N_20503,N_21074);
and U24723 (N_24723,N_21389,N_22089);
and U24724 (N_24724,N_20592,N_20411);
or U24725 (N_24725,N_22082,N_22187);
or U24726 (N_24726,N_22013,N_22240);
or U24727 (N_24727,N_21182,N_21887);
nand U24728 (N_24728,N_21771,N_21934);
or U24729 (N_24729,N_21187,N_21048);
xnor U24730 (N_24730,N_20539,N_20468);
nor U24731 (N_24731,N_20276,N_21463);
xor U24732 (N_24732,N_20124,N_21626);
nand U24733 (N_24733,N_20978,N_21481);
nor U24734 (N_24734,N_22485,N_20834);
and U24735 (N_24735,N_20266,N_22441);
nand U24736 (N_24736,N_22457,N_20446);
xnor U24737 (N_24737,N_22460,N_21190);
nor U24738 (N_24738,N_21496,N_20814);
xnor U24739 (N_24739,N_20746,N_21951);
and U24740 (N_24740,N_21743,N_21924);
or U24741 (N_24741,N_21523,N_22055);
nand U24742 (N_24742,N_20795,N_21392);
and U24743 (N_24743,N_21482,N_22092);
or U24744 (N_24744,N_21709,N_21352);
nand U24745 (N_24745,N_21529,N_20027);
and U24746 (N_24746,N_20410,N_21958);
nand U24747 (N_24747,N_21878,N_20250);
nand U24748 (N_24748,N_21072,N_20533);
nand U24749 (N_24749,N_20848,N_20181);
or U24750 (N_24750,N_20852,N_20048);
nor U24751 (N_24751,N_22412,N_21109);
nor U24752 (N_24752,N_20547,N_22239);
or U24753 (N_24753,N_21145,N_21797);
and U24754 (N_24754,N_20850,N_20011);
or U24755 (N_24755,N_21164,N_21053);
nor U24756 (N_24756,N_20728,N_22471);
and U24757 (N_24757,N_20834,N_20443);
nor U24758 (N_24758,N_22448,N_21550);
nand U24759 (N_24759,N_20927,N_21730);
and U24760 (N_24760,N_20049,N_21085);
nand U24761 (N_24761,N_22306,N_21236);
or U24762 (N_24762,N_21780,N_21145);
or U24763 (N_24763,N_21396,N_22396);
nor U24764 (N_24764,N_21187,N_20963);
xnor U24765 (N_24765,N_22388,N_22256);
xnor U24766 (N_24766,N_22332,N_20389);
and U24767 (N_24767,N_22053,N_20627);
nand U24768 (N_24768,N_20433,N_21135);
or U24769 (N_24769,N_21829,N_20237);
and U24770 (N_24770,N_22022,N_21166);
xnor U24771 (N_24771,N_22225,N_22142);
and U24772 (N_24772,N_20482,N_21683);
nand U24773 (N_24773,N_22197,N_22355);
and U24774 (N_24774,N_22247,N_21051);
or U24775 (N_24775,N_22491,N_20710);
and U24776 (N_24776,N_20229,N_20814);
nand U24777 (N_24777,N_22191,N_21323);
xor U24778 (N_24778,N_22105,N_20814);
and U24779 (N_24779,N_20198,N_22398);
xnor U24780 (N_24780,N_21229,N_21921);
nand U24781 (N_24781,N_20557,N_21340);
and U24782 (N_24782,N_20108,N_21742);
xnor U24783 (N_24783,N_22044,N_21326);
xnor U24784 (N_24784,N_20827,N_22391);
nand U24785 (N_24785,N_21356,N_21397);
nand U24786 (N_24786,N_20214,N_21043);
nor U24787 (N_24787,N_21467,N_20238);
nand U24788 (N_24788,N_20462,N_22321);
xor U24789 (N_24789,N_21096,N_20598);
and U24790 (N_24790,N_22381,N_21358);
xor U24791 (N_24791,N_21821,N_22073);
xor U24792 (N_24792,N_21412,N_21555);
or U24793 (N_24793,N_20397,N_22237);
xnor U24794 (N_24794,N_20010,N_21844);
or U24795 (N_24795,N_22066,N_20807);
or U24796 (N_24796,N_22039,N_20294);
and U24797 (N_24797,N_21341,N_22077);
nor U24798 (N_24798,N_20354,N_21345);
or U24799 (N_24799,N_21313,N_20347);
xnor U24800 (N_24800,N_22494,N_21814);
nand U24801 (N_24801,N_20058,N_21540);
and U24802 (N_24802,N_21944,N_20751);
or U24803 (N_24803,N_22074,N_20935);
and U24804 (N_24804,N_22487,N_20288);
and U24805 (N_24805,N_20653,N_20896);
and U24806 (N_24806,N_21928,N_20854);
nor U24807 (N_24807,N_22493,N_21028);
or U24808 (N_24808,N_21349,N_21295);
nand U24809 (N_24809,N_20941,N_22459);
or U24810 (N_24810,N_20232,N_22202);
or U24811 (N_24811,N_21030,N_22169);
nand U24812 (N_24812,N_21039,N_22486);
nand U24813 (N_24813,N_21487,N_22315);
nand U24814 (N_24814,N_22145,N_20457);
xor U24815 (N_24815,N_21763,N_21510);
nor U24816 (N_24816,N_20479,N_22462);
xnor U24817 (N_24817,N_20249,N_21832);
xnor U24818 (N_24818,N_20631,N_22208);
nand U24819 (N_24819,N_21865,N_22315);
nand U24820 (N_24820,N_22402,N_21750);
xor U24821 (N_24821,N_20407,N_21018);
and U24822 (N_24822,N_20485,N_20812);
and U24823 (N_24823,N_20459,N_20628);
nand U24824 (N_24824,N_20228,N_22263);
or U24825 (N_24825,N_21196,N_22218);
xnor U24826 (N_24826,N_21843,N_21955);
nor U24827 (N_24827,N_20882,N_21336);
nand U24828 (N_24828,N_21802,N_21364);
nand U24829 (N_24829,N_21853,N_21089);
xor U24830 (N_24830,N_20466,N_21913);
nor U24831 (N_24831,N_20343,N_21997);
and U24832 (N_24832,N_21119,N_21968);
nand U24833 (N_24833,N_22179,N_20078);
nand U24834 (N_24834,N_21196,N_21154);
nor U24835 (N_24835,N_21118,N_22273);
xor U24836 (N_24836,N_21407,N_21861);
nor U24837 (N_24837,N_20019,N_20631);
nor U24838 (N_24838,N_21385,N_21968);
xnor U24839 (N_24839,N_22479,N_20828);
nor U24840 (N_24840,N_21920,N_21485);
and U24841 (N_24841,N_20367,N_21113);
xnor U24842 (N_24842,N_21310,N_21947);
nand U24843 (N_24843,N_20620,N_20817);
nand U24844 (N_24844,N_22499,N_21170);
or U24845 (N_24845,N_21671,N_21118);
nor U24846 (N_24846,N_22006,N_21500);
and U24847 (N_24847,N_22333,N_20573);
xnor U24848 (N_24848,N_20044,N_20005);
nand U24849 (N_24849,N_21928,N_20840);
nand U24850 (N_24850,N_21938,N_21569);
or U24851 (N_24851,N_21022,N_22118);
or U24852 (N_24852,N_20884,N_22174);
nor U24853 (N_24853,N_20416,N_22064);
nor U24854 (N_24854,N_20508,N_21873);
nor U24855 (N_24855,N_22175,N_21120);
xor U24856 (N_24856,N_20787,N_22315);
nor U24857 (N_24857,N_21788,N_21872);
or U24858 (N_24858,N_20304,N_21088);
nand U24859 (N_24859,N_22493,N_22093);
and U24860 (N_24860,N_21673,N_20938);
or U24861 (N_24861,N_21472,N_21566);
or U24862 (N_24862,N_22023,N_21575);
and U24863 (N_24863,N_22258,N_20111);
nor U24864 (N_24864,N_22383,N_22001);
and U24865 (N_24865,N_21157,N_20539);
or U24866 (N_24866,N_21943,N_21006);
nand U24867 (N_24867,N_20678,N_20818);
nor U24868 (N_24868,N_21649,N_21519);
nor U24869 (N_24869,N_21500,N_22144);
xor U24870 (N_24870,N_20557,N_21046);
or U24871 (N_24871,N_21930,N_20696);
xor U24872 (N_24872,N_20690,N_21976);
nand U24873 (N_24873,N_22444,N_21228);
nor U24874 (N_24874,N_20401,N_21734);
nor U24875 (N_24875,N_20100,N_22001);
and U24876 (N_24876,N_20465,N_20681);
nand U24877 (N_24877,N_21601,N_20879);
or U24878 (N_24878,N_22199,N_20418);
and U24879 (N_24879,N_21374,N_21462);
nor U24880 (N_24880,N_21566,N_20728);
nor U24881 (N_24881,N_22273,N_22317);
or U24882 (N_24882,N_21699,N_21269);
nand U24883 (N_24883,N_21855,N_20823);
or U24884 (N_24884,N_21407,N_21829);
and U24885 (N_24885,N_20835,N_20626);
and U24886 (N_24886,N_20640,N_20672);
or U24887 (N_24887,N_21651,N_20674);
nor U24888 (N_24888,N_20523,N_21618);
xor U24889 (N_24889,N_20826,N_21831);
nor U24890 (N_24890,N_20988,N_22157);
or U24891 (N_24891,N_22246,N_20185);
xor U24892 (N_24892,N_21179,N_20564);
nand U24893 (N_24893,N_21284,N_20364);
nand U24894 (N_24894,N_21552,N_21492);
nand U24895 (N_24895,N_21142,N_20260);
and U24896 (N_24896,N_21353,N_21548);
nor U24897 (N_24897,N_20299,N_22204);
nor U24898 (N_24898,N_22392,N_20243);
and U24899 (N_24899,N_22112,N_21798);
and U24900 (N_24900,N_22364,N_21252);
nor U24901 (N_24901,N_20606,N_21034);
and U24902 (N_24902,N_21219,N_20981);
nor U24903 (N_24903,N_22398,N_21725);
nor U24904 (N_24904,N_22109,N_21730);
or U24905 (N_24905,N_22310,N_21315);
xnor U24906 (N_24906,N_20048,N_20657);
and U24907 (N_24907,N_21652,N_22495);
or U24908 (N_24908,N_21454,N_20521);
xnor U24909 (N_24909,N_20073,N_20833);
xor U24910 (N_24910,N_22339,N_21017);
nor U24911 (N_24911,N_22059,N_22183);
nor U24912 (N_24912,N_21014,N_22387);
nand U24913 (N_24913,N_21230,N_21408);
or U24914 (N_24914,N_21491,N_22067);
nand U24915 (N_24915,N_20775,N_21657);
nand U24916 (N_24916,N_21732,N_21286);
and U24917 (N_24917,N_20192,N_20705);
nor U24918 (N_24918,N_21582,N_21380);
nor U24919 (N_24919,N_20717,N_20838);
xnor U24920 (N_24920,N_21356,N_20146);
xnor U24921 (N_24921,N_20237,N_22063);
and U24922 (N_24922,N_21422,N_21708);
and U24923 (N_24923,N_21780,N_21829);
nand U24924 (N_24924,N_21143,N_20254);
xor U24925 (N_24925,N_20537,N_20809);
nor U24926 (N_24926,N_21577,N_20719);
nor U24927 (N_24927,N_20642,N_20000);
and U24928 (N_24928,N_20356,N_20416);
or U24929 (N_24929,N_20088,N_21638);
or U24930 (N_24930,N_20939,N_22455);
or U24931 (N_24931,N_20777,N_20344);
and U24932 (N_24932,N_22428,N_21115);
or U24933 (N_24933,N_20832,N_22140);
and U24934 (N_24934,N_20896,N_20670);
nor U24935 (N_24935,N_20287,N_21877);
xor U24936 (N_24936,N_20203,N_20170);
or U24937 (N_24937,N_20789,N_22327);
nor U24938 (N_24938,N_21937,N_21926);
nor U24939 (N_24939,N_21077,N_20026);
xnor U24940 (N_24940,N_20216,N_20369);
nor U24941 (N_24941,N_22488,N_20592);
xnor U24942 (N_24942,N_21555,N_21832);
nand U24943 (N_24943,N_22164,N_22137);
or U24944 (N_24944,N_22401,N_20857);
xnor U24945 (N_24945,N_20918,N_20943);
nand U24946 (N_24946,N_20629,N_21813);
nor U24947 (N_24947,N_20895,N_21730);
and U24948 (N_24948,N_21787,N_20201);
or U24949 (N_24949,N_20803,N_20813);
nor U24950 (N_24950,N_21454,N_22369);
and U24951 (N_24951,N_21437,N_20471);
xor U24952 (N_24952,N_22450,N_20053);
xor U24953 (N_24953,N_20546,N_22132);
or U24954 (N_24954,N_21016,N_20088);
or U24955 (N_24955,N_21974,N_21940);
xnor U24956 (N_24956,N_22059,N_21516);
nand U24957 (N_24957,N_22337,N_21749);
nor U24958 (N_24958,N_20796,N_20281);
xor U24959 (N_24959,N_21420,N_22475);
nor U24960 (N_24960,N_22188,N_20111);
nor U24961 (N_24961,N_20794,N_21154);
and U24962 (N_24962,N_20393,N_20350);
or U24963 (N_24963,N_20177,N_22271);
xor U24964 (N_24964,N_20620,N_20862);
and U24965 (N_24965,N_20622,N_20668);
xnor U24966 (N_24966,N_21992,N_21591);
xor U24967 (N_24967,N_20482,N_22252);
and U24968 (N_24968,N_20089,N_22335);
or U24969 (N_24969,N_21970,N_21625);
xnor U24970 (N_24970,N_20722,N_22479);
nor U24971 (N_24971,N_22047,N_21560);
xnor U24972 (N_24972,N_20610,N_22175);
xnor U24973 (N_24973,N_22026,N_20621);
and U24974 (N_24974,N_20528,N_21926);
or U24975 (N_24975,N_20485,N_20332);
or U24976 (N_24976,N_21446,N_21081);
and U24977 (N_24977,N_22486,N_22075);
or U24978 (N_24978,N_21379,N_22167);
xnor U24979 (N_24979,N_21856,N_20161);
xor U24980 (N_24980,N_21771,N_22034);
xor U24981 (N_24981,N_20317,N_21052);
and U24982 (N_24982,N_22216,N_22014);
nor U24983 (N_24983,N_22351,N_20065);
xnor U24984 (N_24984,N_20478,N_20172);
nor U24985 (N_24985,N_21022,N_21294);
and U24986 (N_24986,N_21882,N_21808);
and U24987 (N_24987,N_21476,N_21578);
or U24988 (N_24988,N_20169,N_20010);
nand U24989 (N_24989,N_20162,N_21174);
nand U24990 (N_24990,N_20904,N_20429);
and U24991 (N_24991,N_20900,N_20603);
and U24992 (N_24992,N_20373,N_22042);
nor U24993 (N_24993,N_20066,N_21094);
xor U24994 (N_24994,N_20632,N_20859);
nand U24995 (N_24995,N_22369,N_21146);
or U24996 (N_24996,N_20599,N_20856);
nor U24997 (N_24997,N_21128,N_20183);
xor U24998 (N_24998,N_21745,N_20136);
xnor U24999 (N_24999,N_20062,N_21648);
nand U25000 (N_25000,N_24839,N_23613);
nand U25001 (N_25001,N_23815,N_22872);
xor U25002 (N_25002,N_22793,N_24545);
nor U25003 (N_25003,N_23761,N_23789);
xor U25004 (N_25004,N_22920,N_24803);
nand U25005 (N_25005,N_23132,N_24102);
xor U25006 (N_25006,N_24166,N_24665);
or U25007 (N_25007,N_24008,N_22982);
nor U25008 (N_25008,N_24368,N_24666);
xor U25009 (N_25009,N_23906,N_23072);
or U25010 (N_25010,N_22785,N_23721);
nand U25011 (N_25011,N_24083,N_23223);
or U25012 (N_25012,N_24825,N_24869);
or U25013 (N_25013,N_24196,N_23590);
and U25014 (N_25014,N_24997,N_22968);
and U25015 (N_25015,N_24721,N_23288);
nor U25016 (N_25016,N_24565,N_24964);
and U25017 (N_25017,N_22877,N_24677);
nor U25018 (N_25018,N_24408,N_23491);
and U25019 (N_25019,N_24375,N_23099);
xor U25020 (N_25020,N_23151,N_24880);
xor U25021 (N_25021,N_24920,N_24608);
and U25022 (N_25022,N_23283,N_24082);
nand U25023 (N_25023,N_24468,N_23543);
or U25024 (N_25024,N_23946,N_23429);
nor U25025 (N_25025,N_23193,N_24984);
and U25026 (N_25026,N_22909,N_22811);
nor U25027 (N_25027,N_23595,N_22572);
nor U25028 (N_25028,N_24830,N_22706);
nor U25029 (N_25029,N_23125,N_24999);
or U25030 (N_25030,N_23292,N_24541);
or U25031 (N_25031,N_23790,N_23091);
and U25032 (N_25032,N_23920,N_22542);
nand U25033 (N_25033,N_24135,N_23318);
xor U25034 (N_25034,N_22721,N_23402);
or U25035 (N_25035,N_23059,N_23123);
xnor U25036 (N_25036,N_23286,N_23069);
nor U25037 (N_25037,N_23084,N_23976);
or U25038 (N_25038,N_24316,N_24497);
nor U25039 (N_25039,N_24722,N_24584);
nor U25040 (N_25040,N_24380,N_23020);
nor U25041 (N_25041,N_24042,N_22611);
nor U25042 (N_25042,N_24851,N_24988);
nor U25043 (N_25043,N_24471,N_23396);
xor U25044 (N_25044,N_23332,N_23531);
nand U25045 (N_25045,N_22635,N_24965);
nand U25046 (N_25046,N_23948,N_22709);
nand U25047 (N_25047,N_23350,N_23953);
or U25048 (N_25048,N_24615,N_24759);
xor U25049 (N_25049,N_22955,N_23664);
or U25050 (N_25050,N_23743,N_23235);
and U25051 (N_25051,N_24208,N_24342);
or U25052 (N_25052,N_24566,N_24612);
nor U25053 (N_25053,N_24231,N_24694);
nand U25054 (N_25054,N_24774,N_23588);
or U25055 (N_25055,N_23724,N_24801);
xnor U25056 (N_25056,N_23453,N_22832);
nor U25057 (N_25057,N_23206,N_24422);
or U25058 (N_25058,N_22645,N_24872);
nor U25059 (N_25059,N_24621,N_24922);
and U25060 (N_25060,N_23931,N_23044);
xnor U25061 (N_25061,N_24732,N_23498);
nand U25062 (N_25062,N_24619,N_23347);
and U25063 (N_25063,N_22949,N_24059);
nand U25064 (N_25064,N_24553,N_23477);
nor U25065 (N_25065,N_22505,N_23984);
nor U25066 (N_25066,N_22613,N_23112);
nand U25067 (N_25067,N_22624,N_24815);
and U25068 (N_25068,N_23582,N_24601);
and U25069 (N_25069,N_24182,N_22500);
xor U25070 (N_25070,N_22735,N_23136);
nor U25071 (N_25071,N_24288,N_23162);
or U25072 (N_25072,N_24167,N_23969);
nand U25073 (N_25073,N_24210,N_23506);
and U25074 (N_25074,N_24117,N_24644);
or U25075 (N_25075,N_22555,N_24020);
xor U25076 (N_25076,N_22634,N_24290);
or U25077 (N_25077,N_24053,N_23379);
xor U25078 (N_25078,N_23488,N_23010);
and U25079 (N_25079,N_22599,N_23441);
nand U25080 (N_25080,N_22797,N_23267);
and U25081 (N_25081,N_24409,N_22775);
and U25082 (N_25082,N_24670,N_23312);
nand U25083 (N_25083,N_24360,N_23266);
nor U25084 (N_25084,N_23411,N_24578);
or U25085 (N_25085,N_22529,N_22743);
nor U25086 (N_25086,N_22547,N_24533);
and U25087 (N_25087,N_24482,N_24931);
xnor U25088 (N_25088,N_24884,N_23601);
nor U25089 (N_25089,N_22571,N_24646);
nand U25090 (N_25090,N_22621,N_23179);
nand U25091 (N_25091,N_23509,N_23838);
nor U25092 (N_25092,N_22586,N_22890);
and U25093 (N_25093,N_23591,N_24241);
nand U25094 (N_25094,N_23363,N_24847);
nor U25095 (N_25095,N_24357,N_23034);
or U25096 (N_25096,N_22615,N_24456);
or U25097 (N_25097,N_24430,N_23291);
nand U25098 (N_25098,N_24831,N_24087);
nor U25099 (N_25099,N_23188,N_23698);
and U25100 (N_25100,N_24770,N_22892);
and U25101 (N_25101,N_24443,N_24900);
or U25102 (N_25102,N_24274,N_23598);
nor U25103 (N_25103,N_23416,N_22759);
nor U25104 (N_25104,N_23476,N_24558);
and U25105 (N_25105,N_24062,N_24433);
xor U25106 (N_25106,N_24969,N_23997);
nor U25107 (N_25107,N_24729,N_22703);
nand U25108 (N_25108,N_24188,N_23225);
xnor U25109 (N_25109,N_23460,N_23515);
nor U25110 (N_25110,N_23327,N_24426);
xor U25111 (N_25111,N_24664,N_23618);
xor U25112 (N_25112,N_24377,N_23690);
and U25113 (N_25113,N_23486,N_23699);
or U25114 (N_25114,N_24286,N_24275);
nor U25115 (N_25115,N_23321,N_24001);
or U25116 (N_25116,N_24459,N_24628);
and U25117 (N_25117,N_22847,N_22679);
nor U25118 (N_25118,N_24346,N_23454);
nand U25119 (N_25119,N_24766,N_23541);
nor U25120 (N_25120,N_23717,N_24516);
nand U25121 (N_25121,N_22819,N_24014);
xor U25122 (N_25122,N_23804,N_24779);
nor U25123 (N_25123,N_23482,N_23102);
nand U25124 (N_25124,N_23787,N_23759);
xor U25125 (N_25125,N_23277,N_24473);
and U25126 (N_25126,N_23417,N_22822);
nand U25127 (N_25127,N_24239,N_22535);
nor U25128 (N_25128,N_22975,N_22526);
nor U25129 (N_25129,N_24325,N_22821);
or U25130 (N_25130,N_23234,N_24760);
or U25131 (N_25131,N_24451,N_23280);
or U25132 (N_25132,N_23819,N_23957);
or U25133 (N_25133,N_22928,N_24370);
xor U25134 (N_25134,N_23144,N_23974);
nor U25135 (N_25135,N_24777,N_22812);
and U25136 (N_25136,N_24324,N_22708);
xor U25137 (N_25137,N_23782,N_22632);
xnor U25138 (N_25138,N_23923,N_23097);
nor U25139 (N_25139,N_24273,N_24054);
nand U25140 (N_25140,N_24101,N_24491);
and U25141 (N_25141,N_24199,N_24667);
xnor U25142 (N_25142,N_24414,N_23424);
or U25143 (N_25143,N_24149,N_24662);
and U25144 (N_25144,N_23092,N_24121);
and U25145 (N_25145,N_23085,N_24023);
nand U25146 (N_25146,N_24725,N_22844);
nor U25147 (N_25147,N_23461,N_23547);
nand U25148 (N_25148,N_22995,N_24356);
and U25149 (N_25149,N_22864,N_23192);
nor U25150 (N_25150,N_23539,N_22715);
nor U25151 (N_25151,N_22751,N_23552);
xor U25152 (N_25152,N_24189,N_23557);
xnor U25153 (N_25153,N_24844,N_22673);
xnor U25154 (N_25154,N_22963,N_24962);
and U25155 (N_25155,N_22912,N_23051);
xnor U25156 (N_25156,N_23258,N_23875);
nor U25157 (N_25157,N_23121,N_23302);
nand U25158 (N_25158,N_24030,N_23777);
xor U25159 (N_25159,N_23571,N_24379);
nor U25160 (N_25160,N_24950,N_22697);
xor U25161 (N_25161,N_23653,N_24994);
xor U25162 (N_25162,N_23968,N_23130);
nand U25163 (N_25163,N_23232,N_24811);
nor U25164 (N_25164,N_23306,N_23849);
or U25165 (N_25165,N_22591,N_22704);
and U25166 (N_25166,N_23304,N_24604);
and U25167 (N_25167,N_24095,N_23154);
xnor U25168 (N_25168,N_24319,N_23928);
xor U25169 (N_25169,N_23471,N_24376);
and U25170 (N_25170,N_24484,N_23317);
nor U25171 (N_25171,N_22910,N_22658);
nand U25172 (N_25172,N_24685,N_23328);
nand U25173 (N_25173,N_24944,N_24209);
nand U25174 (N_25174,N_22630,N_23702);
xnor U25175 (N_25175,N_24778,N_24192);
xnor U25176 (N_25176,N_24501,N_24133);
or U25177 (N_25177,N_24855,N_23855);
xnor U25178 (N_25178,N_23432,N_23750);
nor U25179 (N_25179,N_24036,N_24983);
and U25180 (N_25180,N_23636,N_23854);
nor U25181 (N_25181,N_24879,N_22998);
xor U25182 (N_25182,N_23683,N_23269);
and U25183 (N_25183,N_22727,N_23391);
or U25184 (N_25184,N_22923,N_23722);
xnor U25185 (N_25185,N_23894,N_23305);
nor U25186 (N_25186,N_23061,N_24183);
or U25187 (N_25187,N_23585,N_24048);
nor U25188 (N_25188,N_24589,N_23958);
nand U25189 (N_25189,N_23298,N_24554);
or U25190 (N_25190,N_24603,N_24049);
and U25191 (N_25191,N_22807,N_23848);
nor U25192 (N_25192,N_23274,N_24650);
nor U25193 (N_25193,N_23988,N_24898);
xnor U25194 (N_25194,N_24986,N_24509);
xor U25195 (N_25195,N_23314,N_23459);
nand U25196 (N_25196,N_24098,N_24245);
nor U25197 (N_25197,N_24306,N_24906);
nor U25198 (N_25198,N_22986,N_23129);
nand U25199 (N_25199,N_23325,N_23510);
nor U25200 (N_25200,N_23368,N_24613);
or U25201 (N_25201,N_23555,N_22941);
xor U25202 (N_25202,N_24493,N_23545);
nand U25203 (N_25203,N_23261,N_23430);
nand U25204 (N_25204,N_23190,N_24506);
xor U25205 (N_25205,N_22991,N_23201);
nor U25206 (N_25206,N_23898,N_22809);
and U25207 (N_25207,N_24918,N_23117);
or U25208 (N_25208,N_23995,N_23043);
and U25209 (N_25209,N_23271,N_22659);
nand U25210 (N_25210,N_24293,N_22996);
nor U25211 (N_25211,N_24849,N_24436);
or U25212 (N_25212,N_23310,N_24873);
nor U25213 (N_25213,N_24405,N_24576);
xor U25214 (N_25214,N_23566,N_23633);
xor U25215 (N_25215,N_23927,N_24452);
and U25216 (N_25216,N_23670,N_23941);
xnor U25217 (N_25217,N_23666,N_22929);
and U25218 (N_25218,N_23297,N_22707);
nor U25219 (N_25219,N_22870,N_22947);
nor U25220 (N_25220,N_23727,N_24065);
and U25221 (N_25221,N_22712,N_24386);
nand U25222 (N_25222,N_24534,N_23448);
xor U25223 (N_25223,N_23446,N_24713);
nor U25224 (N_25224,N_24462,N_22728);
and U25225 (N_25225,N_22800,N_23285);
nor U25226 (N_25226,N_24934,N_24258);
nor U25227 (N_25227,N_23248,N_23165);
xor U25228 (N_25228,N_24201,N_23548);
nand U25229 (N_25229,N_24442,N_23518);
nand U25230 (N_25230,N_24763,N_23352);
or U25231 (N_25231,N_22560,N_22590);
or U25232 (N_25232,N_23290,N_24141);
and U25233 (N_25233,N_23829,N_23975);
nor U25234 (N_25234,N_23167,N_23684);
nor U25235 (N_25235,N_23216,N_24846);
nor U25236 (N_25236,N_24792,N_23888);
and U25237 (N_25237,N_23977,N_24315);
nand U25238 (N_25238,N_23646,N_24094);
and U25239 (N_25239,N_24009,N_23853);
and U25240 (N_25240,N_24622,N_24546);
nor U25241 (N_25241,N_23542,N_22738);
and U25242 (N_25242,N_23361,N_23103);
nor U25243 (N_25243,N_24813,N_23532);
nand U25244 (N_25244,N_23115,N_24013);
nor U25245 (N_25245,N_22579,N_24798);
nand U25246 (N_25246,N_24060,N_22852);
or U25247 (N_25247,N_24657,N_24365);
nand U25248 (N_25248,N_24384,N_24397);
xor U25249 (N_25249,N_22898,N_22965);
or U25250 (N_25250,N_24215,N_24543);
and U25251 (N_25251,N_23611,N_22772);
or U25252 (N_25252,N_24431,N_24564);
and U25253 (N_25253,N_23281,N_22519);
xnor U25254 (N_25254,N_23708,N_24161);
and U25255 (N_25255,N_23839,N_23282);
xor U25256 (N_25256,N_23457,N_24282);
nand U25257 (N_25257,N_22696,N_23315);
or U25258 (N_25258,N_23648,N_22960);
xor U25259 (N_25259,N_23249,N_23307);
and U25260 (N_25260,N_22845,N_24096);
nor U25261 (N_25261,N_22680,N_24720);
and U25262 (N_25262,N_24861,N_23870);
or U25263 (N_25263,N_22565,N_22976);
or U25264 (N_25264,N_24883,N_22527);
nor U25265 (N_25265,N_23578,N_24814);
nor U25266 (N_25266,N_22989,N_24416);
and U25267 (N_25267,N_22858,N_23983);
or U25268 (N_25268,N_22918,N_23148);
nor U25269 (N_25269,N_22914,N_22665);
and U25270 (N_25270,N_23109,N_24887);
nand U25271 (N_25271,N_22523,N_23039);
or U25272 (N_25272,N_24595,N_23828);
xor U25273 (N_25273,N_24382,N_24304);
xor U25274 (N_25274,N_23407,N_24527);
xnor U25275 (N_25275,N_24015,N_24842);
xor U25276 (N_25276,N_24289,N_24047);
xor U25277 (N_25277,N_24206,N_22574);
and U25278 (N_25278,N_23512,N_24165);
or U25279 (N_25279,N_23651,N_22862);
nor U25280 (N_25280,N_23577,N_22808);
nor U25281 (N_25281,N_22810,N_24785);
and U25282 (N_25282,N_22924,N_24993);
or U25283 (N_25283,N_23279,N_23824);
and U25284 (N_25284,N_23268,N_22552);
xor U25285 (N_25285,N_23674,N_22512);
or U25286 (N_25286,N_23354,N_24061);
nor U25287 (N_25287,N_23233,N_22532);
or U25288 (N_25288,N_22884,N_23326);
xnor U25289 (N_25289,N_23047,N_23776);
and U25290 (N_25290,N_23987,N_22753);
xor U25291 (N_25291,N_22863,N_22806);
or U25292 (N_25292,N_24281,N_24904);
nor U25293 (N_25293,N_23319,N_24810);
and U25294 (N_25294,N_23348,N_23623);
or U25295 (N_25295,N_24418,N_24413);
and U25296 (N_25296,N_22652,N_23944);
nand U25297 (N_25297,N_24871,N_24753);
and U25298 (N_25298,N_24594,N_23676);
nand U25299 (N_25299,N_23796,N_23821);
nand U25300 (N_25300,N_23001,N_24629);
nor U25301 (N_25301,N_24560,N_22602);
and U25302 (N_25302,N_24929,N_23871);
and U25303 (N_25303,N_23514,N_24140);
and U25304 (N_25304,N_22685,N_22776);
nand U25305 (N_25305,N_23800,N_24874);
and U25306 (N_25306,N_24264,N_23746);
or U25307 (N_25307,N_22618,N_23309);
nor U25308 (N_25308,N_23823,N_24562);
nand U25309 (N_25309,N_24152,N_22643);
nor U25310 (N_25310,N_22691,N_23925);
xor U25311 (N_25311,N_22952,N_22961);
nor U25312 (N_25312,N_24772,N_24512);
nor U25313 (N_25313,N_23797,N_22916);
or U25314 (N_25314,N_23140,N_24794);
nor U25315 (N_25315,N_23608,N_23924);
or U25316 (N_25316,N_23035,N_24691);
nor U25317 (N_25317,N_24446,N_23600);
nor U25318 (N_25318,N_24859,N_22663);
and U25319 (N_25319,N_24817,N_24336);
xnor U25320 (N_25320,N_23351,N_23709);
xor U25321 (N_25321,N_22631,N_24321);
or U25322 (N_25322,N_24947,N_23986);
xnor U25323 (N_25323,N_23067,N_24756);
nor U25324 (N_25324,N_23852,N_23264);
and U25325 (N_25325,N_24498,N_24795);
nor U25326 (N_25326,N_23626,N_23970);
nor U25327 (N_25327,N_24585,N_22686);
or U25328 (N_25328,N_23023,N_23725);
xor U25329 (N_25329,N_22554,N_24132);
nand U25330 (N_25330,N_24190,N_22622);
or U25331 (N_25331,N_23414,N_22550);
or U25332 (N_25332,N_24178,N_24051);
xor U25333 (N_25333,N_24109,N_24806);
xnor U25334 (N_25334,N_24742,N_24067);
or U25335 (N_25335,N_23889,N_24353);
and U25336 (N_25336,N_22860,N_23723);
nor U25337 (N_25337,N_24122,N_23998);
and U25338 (N_25338,N_24521,N_22623);
xnor U25339 (N_25339,N_23805,N_23745);
nand U25340 (N_25340,N_24461,N_22661);
nand U25341 (N_25341,N_23570,N_22689);
xnor U25342 (N_25342,N_24680,N_24039);
nand U25343 (N_25343,N_23668,N_24428);
xor U25344 (N_25344,N_23138,N_22873);
xor U25345 (N_25345,N_23594,N_22829);
xnor U25346 (N_25346,N_23816,N_22805);
or U25347 (N_25347,N_24998,N_24513);
xnor U25348 (N_25348,N_23388,N_22934);
nand U25349 (N_25349,N_24676,N_23330);
nand U25350 (N_25350,N_24186,N_22700);
nor U25351 (N_25351,N_24262,N_23141);
nand U25352 (N_25352,N_23357,N_24526);
nand U25353 (N_25353,N_23916,N_22839);
and U25354 (N_25354,N_23753,N_23041);
xnor U25355 (N_25355,N_24157,N_24385);
xor U25356 (N_25356,N_22504,N_24181);
and U25357 (N_25357,N_24099,N_23873);
and U25358 (N_25358,N_24507,N_24352);
or U25359 (N_25359,N_24727,N_23569);
nand U25360 (N_25360,N_23134,N_23949);
and U25361 (N_25361,N_24388,N_23730);
and U25362 (N_25362,N_23485,N_22931);
nand U25363 (N_25363,N_22945,N_23042);
nor U25364 (N_25364,N_23226,N_23250);
or U25365 (N_25365,N_23341,N_23857);
xor U25366 (N_25366,N_23086,N_23003);
xor U25367 (N_25367,N_24271,N_24848);
and U25368 (N_25368,N_23803,N_24710);
nor U25369 (N_25369,N_22939,N_22940);
and U25370 (N_25370,N_23369,N_24320);
or U25371 (N_25371,N_24230,N_22857);
xor U25372 (N_25372,N_22840,N_24755);
xor U25373 (N_25373,N_23869,N_23886);
nor U25374 (N_25374,N_24125,N_23647);
nand U25375 (N_25375,N_24953,N_24350);
or U25376 (N_25376,N_23468,N_22980);
nand U25377 (N_25377,N_22951,N_24466);
nor U25378 (N_25378,N_24715,N_23996);
and U25379 (N_25379,N_22551,N_23101);
or U25380 (N_25380,N_24055,N_24228);
or U25381 (N_25381,N_23016,N_24309);
nand U25382 (N_25382,N_23435,N_22693);
and U25383 (N_25383,N_24735,N_23398);
nor U25384 (N_25384,N_24620,N_22978);
and U25385 (N_25385,N_24706,N_23574);
or U25386 (N_25386,N_22506,N_23519);
and U25387 (N_25387,N_23386,N_24464);
and U25388 (N_25388,N_24338,N_22593);
nand U25389 (N_25389,N_23170,N_22786);
xor U25390 (N_25390,N_22541,N_23781);
xor U25391 (N_25391,N_24651,N_22831);
xor U25392 (N_25392,N_24723,N_23385);
nand U25393 (N_25393,N_22606,N_24951);
xnor U25394 (N_25394,N_23877,N_23644);
xor U25395 (N_25395,N_22990,N_23456);
nor U25396 (N_25396,N_22647,N_22695);
xnor U25397 (N_25397,N_22641,N_22654);
nor U25398 (N_25398,N_22792,N_22734);
or U25399 (N_25399,N_24441,N_23169);
xor U25400 (N_25400,N_23556,N_23525);
xor U25401 (N_25401,N_23544,N_23173);
and U25402 (N_25402,N_23239,N_23015);
or U25403 (N_25403,N_23529,N_23198);
and U25404 (N_25404,N_23667,N_24640);
or U25405 (N_25405,N_23716,N_24475);
xnor U25406 (N_25406,N_23846,N_22798);
nor U25407 (N_25407,N_24439,N_23056);
nand U25408 (N_25408,N_22770,N_24635);
nand U25409 (N_25409,N_23495,N_24658);
and U25410 (N_25410,N_22617,N_24420);
nand U25411 (N_25411,N_23194,N_24040);
or U25412 (N_25412,N_24177,N_23697);
and U25413 (N_25413,N_23632,N_24679);
xnor U25414 (N_25414,N_23891,N_24381);
nor U25415 (N_25415,N_23534,N_24016);
xnor U25416 (N_25416,N_22773,N_24536);
nand U25417 (N_25417,N_23712,N_24238);
xor U25418 (N_25418,N_24791,N_24295);
and U25419 (N_25419,N_24236,N_24378);
or U25420 (N_25420,N_24519,N_23246);
nor U25421 (N_25421,N_22724,N_23436);
nor U25422 (N_25422,N_24764,N_22537);
nand U25423 (N_25423,N_24556,N_24302);
nand U25424 (N_25424,N_24624,N_23410);
or U25425 (N_25425,N_22531,N_23114);
and U25426 (N_25426,N_22886,N_23622);
or U25427 (N_25427,N_22678,N_24347);
nor U25428 (N_25428,N_24100,N_22999);
and U25429 (N_25429,N_24686,N_23858);
or U25430 (N_25430,N_23550,N_23019);
or U25431 (N_25431,N_22889,N_23247);
nor U25432 (N_25432,N_23224,N_22660);
and U25433 (N_25433,N_23580,N_23994);
xor U25434 (N_25434,N_22666,N_24311);
nor U25435 (N_25435,N_24063,N_24392);
nor U25436 (N_25436,N_23660,N_24250);
and U25437 (N_25437,N_22609,N_23675);
or U25438 (N_25438,N_24124,N_24728);
nor U25439 (N_25439,N_22903,N_22592);
or U25440 (N_25440,N_24470,N_24463);
or U25441 (N_25441,N_24073,N_23265);
xnor U25442 (N_25442,N_24028,N_22874);
and U25443 (N_25443,N_24033,N_22824);
and U25444 (N_25444,N_24411,N_24818);
or U25445 (N_25445,N_24276,N_23419);
and U25446 (N_25446,N_23473,N_23238);
or U25447 (N_25447,N_22901,N_23657);
nor U25448 (N_25448,N_22777,N_24899);
or U25449 (N_25449,N_22736,N_24359);
xnor U25450 (N_25450,N_22675,N_23054);
nor U25451 (N_25451,N_22752,N_24233);
or U25452 (N_25452,N_22534,N_23037);
nand U25453 (N_25453,N_23489,N_22783);
or U25454 (N_25454,N_24467,N_23340);
nand U25455 (N_25455,N_24642,N_23494);
nand U25456 (N_25456,N_22705,N_23336);
xnor U25457 (N_25457,N_23935,N_23775);
nand U25458 (N_25458,N_22917,N_22699);
nand U25459 (N_25459,N_24652,N_22508);
and U25460 (N_25460,N_23017,N_23972);
xnor U25461 (N_25461,N_24398,N_24623);
nand U25462 (N_25462,N_23287,N_23820);
or U25463 (N_25463,N_24614,N_23911);
and U25464 (N_25464,N_24277,N_22754);
nor U25465 (N_25465,N_22984,N_24910);
nand U25466 (N_25466,N_22970,N_22813);
nor U25467 (N_25467,N_24675,N_24116);
nor U25468 (N_25468,N_24719,N_22637);
or U25469 (N_25469,N_24674,N_23863);
nor U25470 (N_25470,N_22546,N_24896);
xnor U25471 (N_25471,N_22842,N_24695);
or U25472 (N_25472,N_24972,N_24809);
or U25473 (N_25473,N_23767,N_22900);
nand U25474 (N_25474,N_23905,N_23449);
or U25475 (N_25475,N_23126,N_23989);
nand U25476 (N_25476,N_23499,N_24151);
and U25477 (N_25477,N_24007,N_23401);
xnor U25478 (N_25478,N_24502,N_24911);
nand U25479 (N_25479,N_22878,N_24169);
nand U25480 (N_25480,N_23062,N_23367);
nand U25481 (N_25481,N_23562,N_22973);
and U25482 (N_25482,N_24399,N_22578);
and U25483 (N_25483,N_23762,N_24348);
or U25484 (N_25484,N_24632,N_24943);
xnor U25485 (N_25485,N_23526,N_24592);
xor U25486 (N_25486,N_23758,N_24607);
xor U25487 (N_25487,N_24307,N_24574);
nand U25488 (N_25488,N_23784,N_24410);
nor U25489 (N_25489,N_24294,N_24750);
xnor U25490 (N_25490,N_22883,N_23474);
nand U25491 (N_25491,N_24137,N_22854);
nand U25492 (N_25492,N_24888,N_24862);
nor U25493 (N_25493,N_23000,N_22642);
or U25494 (N_25494,N_24265,N_23908);
nor U25495 (N_25495,N_23719,N_24396);
and U25496 (N_25496,N_23389,N_23741);
nand U25497 (N_25497,N_24415,N_23813);
or U25498 (N_25498,N_24481,N_23962);
nor U25499 (N_25499,N_24200,N_23842);
xor U25500 (N_25500,N_24003,N_23910);
nand U25501 (N_25501,N_23581,N_24130);
nand U25502 (N_25502,N_23006,N_24902);
nand U25503 (N_25503,N_23253,N_24148);
or U25504 (N_25504,N_23596,N_24726);
nor U25505 (N_25505,N_23458,N_24021);
nand U25506 (N_25506,N_23720,N_24477);
or U25507 (N_25507,N_23812,N_23096);
and U25508 (N_25508,N_24106,N_24826);
nor U25509 (N_25509,N_23237,N_24333);
xnor U25510 (N_25510,N_24598,N_24211);
and U25511 (N_25511,N_24789,N_24852);
and U25512 (N_25512,N_23353,N_24089);
xor U25513 (N_25513,N_24226,N_23152);
xor U25514 (N_25514,N_22802,N_23979);
nor U25515 (N_25515,N_24138,N_23175);
xor U25516 (N_25516,N_22740,N_23936);
nor U25517 (N_25517,N_22894,N_23404);
nor U25518 (N_25518,N_24793,N_22530);
nor U25519 (N_25519,N_22627,N_23625);
nand U25520 (N_25520,N_24240,N_24559);
and U25521 (N_25521,N_24634,N_24864);
or U25522 (N_25522,N_23252,N_23090);
nor U25523 (N_25523,N_24026,N_24268);
and U25524 (N_25524,N_24401,N_23256);
or U25525 (N_25525,N_22790,N_24427);
nor U25526 (N_25526,N_24668,N_23892);
xnor U25527 (N_25527,N_23959,N_24510);
and U25528 (N_25528,N_23832,N_24682);
nor U25529 (N_25529,N_22573,N_24191);
nor U25530 (N_25530,N_24697,N_24834);
xnor U25531 (N_25531,N_22967,N_24542);
nand U25532 (N_25532,N_23573,N_23887);
and U25533 (N_25533,N_24078,N_24771);
and U25534 (N_25534,N_24606,N_23769);
and U25535 (N_25535,N_24828,N_24454);
nand U25536 (N_25536,N_23046,N_23502);
nor U25537 (N_25537,N_22714,N_24701);
nor U25538 (N_25538,N_24123,N_24212);
and U25539 (N_25539,N_23145,N_22969);
and U25540 (N_25540,N_23025,N_23364);
nand U25541 (N_25541,N_23293,N_23158);
nor U25542 (N_25542,N_22742,N_24853);
xor U25543 (N_25543,N_22762,N_23926);
or U25544 (N_25544,N_23100,N_24748);
nor U25545 (N_25545,N_24423,N_22997);
nor U25546 (N_25546,N_22667,N_23742);
nor U25547 (N_25547,N_24229,N_23940);
nor U25548 (N_25548,N_23189,N_23549);
nor U25549 (N_25549,N_22972,N_23747);
nand U25550 (N_25550,N_24158,N_23628);
and U25551 (N_25551,N_24248,N_24091);
nand U25552 (N_25552,N_22992,N_22616);
nor U25553 (N_25553,N_22871,N_24361);
nor U25554 (N_25554,N_23013,N_23211);
and U25555 (N_25555,N_23560,N_22876);
and U25556 (N_25556,N_23786,N_23440);
or U25557 (N_25557,N_23005,N_22887);
or U25558 (N_25558,N_22853,N_22644);
and U25559 (N_25559,N_22778,N_24932);
nand U25560 (N_25560,N_24237,N_24903);
nand U25561 (N_25561,N_24284,N_24979);
nand U25562 (N_25562,N_24362,N_23203);
xor U25563 (N_25563,N_24194,N_22769);
nand U25564 (N_25564,N_23113,N_24909);
xor U25565 (N_25565,N_23075,N_23275);
nand U25566 (N_25566,N_23501,N_23466);
and U25567 (N_25567,N_23415,N_22719);
or U25568 (N_25568,N_24119,N_24981);
nor U25569 (N_25569,N_24499,N_24548);
nor U25570 (N_25570,N_23294,N_24090);
and U25571 (N_25571,N_24256,N_24845);
xor U25572 (N_25572,N_22672,N_24569);
xnor U25573 (N_25573,N_24429,N_22522);
nand U25574 (N_25574,N_23929,N_24034);
nor U25575 (N_25575,N_22942,N_24503);
nor U25576 (N_25576,N_22683,N_23465);
xnor U25577 (N_25577,N_22801,N_24730);
xnor U25578 (N_25578,N_24808,N_24866);
nand U25579 (N_25579,N_24741,N_24086);
and U25580 (N_25580,N_24220,N_23881);
or U25581 (N_25581,N_23068,N_24967);
xnor U25582 (N_25582,N_23692,N_24305);
xnor U25583 (N_25583,N_24247,N_22885);
and U25584 (N_25584,N_22581,N_24908);
xnor U25585 (N_25585,N_23859,N_23426);
and U25586 (N_25586,N_24949,N_22979);
nor U25587 (N_25587,N_24417,N_23359);
nand U25588 (N_25588,N_23847,N_23187);
or U25589 (N_25589,N_23686,N_24025);
xor U25590 (N_25590,N_24630,N_23738);
xnor U25591 (N_25591,N_23654,N_24479);
nor U25592 (N_25592,N_23026,N_24114);
and U25593 (N_25593,N_23358,N_22981);
nor U25594 (N_25594,N_22758,N_24504);
nor U25595 (N_25595,N_23785,N_23659);
nor U25596 (N_25596,N_23553,N_23833);
or U25597 (N_25597,N_23752,N_22690);
or U25598 (N_25598,N_24978,N_24103);
nand U25599 (N_25599,N_24261,N_23083);
and U25600 (N_25600,N_24689,N_22936);
and U25601 (N_25601,N_22922,N_24126);
or U25602 (N_25602,N_23729,N_24591);
and U25603 (N_25603,N_22716,N_24637);
xnor U25604 (N_25604,N_22545,N_22974);
or U25605 (N_25605,N_24337,N_24575);
nor U25606 (N_25606,N_24913,N_23930);
nor U25607 (N_25607,N_22650,N_24093);
and U25608 (N_25608,N_23751,N_22825);
nand U25609 (N_25609,N_24530,N_22958);
or U25610 (N_25610,N_23965,N_24786);
nor U25611 (N_25611,N_24460,N_23893);
nor U25612 (N_25612,N_23011,N_24837);
nor U25613 (N_25613,N_24968,N_23561);
nor U25614 (N_25614,N_22959,N_23434);
xnor U25615 (N_25615,N_23757,N_23445);
and U25616 (N_25616,N_23040,N_23007);
or U25617 (N_25617,N_22653,N_23397);
or U25618 (N_25618,N_23375,N_23262);
xor U25619 (N_25619,N_23323,N_22556);
and U25620 (N_25620,N_23943,N_23810);
or U25621 (N_25621,N_23642,N_24299);
xor U25622 (N_25622,N_24970,N_22726);
nand U25623 (N_25623,N_23807,N_23663);
and U25624 (N_25624,N_24633,N_24364);
and U25625 (N_25625,N_24782,N_22562);
xor U25626 (N_25626,N_23687,N_22760);
and U25627 (N_25627,N_24249,N_22925);
and U25628 (N_25628,N_23685,N_22843);
or U25629 (N_25629,N_23728,N_22838);
xor U25630 (N_25630,N_22649,N_24469);
xor U25631 (N_25631,N_23879,N_23373);
nor U25632 (N_25632,N_24921,N_23120);
nand U25633 (N_25633,N_23004,N_24074);
nand U25634 (N_25634,N_23074,N_23827);
and U25635 (N_25635,N_23381,N_23587);
xnor U25636 (N_25636,N_24625,N_24653);
or U25637 (N_25637,N_23313,N_22766);
nor U25638 (N_25638,N_22533,N_24222);
nand U25639 (N_25639,N_24490,N_23524);
nand U25640 (N_25640,N_23616,N_23655);
and U25641 (N_25641,N_23568,N_23658);
or U25642 (N_25642,N_24163,N_22865);
xnor U25643 (N_25643,N_24129,N_23423);
nand U25644 (N_25644,N_24214,N_23428);
xnor U25645 (N_25645,N_24525,N_22564);
nand U25646 (N_25646,N_22520,N_22629);
nor U25647 (N_25647,N_23210,N_24537);
nor U25648 (N_25648,N_24492,N_23058);
or U25649 (N_25649,N_23022,N_23778);
or U25650 (N_25650,N_22729,N_24954);
nand U25651 (N_25651,N_24941,N_23993);
and U25652 (N_25652,N_24709,N_24816);
xnor U25653 (N_25653,N_23128,N_24843);
nor U25654 (N_25654,N_22732,N_23980);
and U25655 (N_25655,N_23339,N_24681);
and U25656 (N_25656,N_24531,N_22636);
and U25657 (N_25657,N_22646,N_24660);
or U25658 (N_25658,N_24649,N_24586);
and U25659 (N_25659,N_23093,N_23830);
nand U25660 (N_25660,N_24757,N_23071);
xnor U25661 (N_25661,N_24010,N_23094);
or U25662 (N_25662,N_23029,N_24850);
nand U25663 (N_25663,N_22604,N_24627);
nor U25664 (N_25664,N_23740,N_23551);
and U25665 (N_25665,N_22781,N_23376);
nand U25666 (N_25666,N_23146,N_23770);
nor U25667 (N_25667,N_22861,N_22656);
or U25668 (N_25668,N_23221,N_24363);
or U25669 (N_25669,N_24259,N_24802);
xnor U25670 (N_25670,N_23731,N_24907);
or U25671 (N_25671,N_23982,N_22668);
nor U25672 (N_25672,N_24821,N_23774);
xnor U25673 (N_25673,N_24407,N_24982);
or U25674 (N_25674,N_24232,N_23133);
nand U25675 (N_25675,N_22639,N_23338);
nor U25676 (N_25676,N_22834,N_23480);
nand U25677 (N_25677,N_24656,N_24734);
or U25678 (N_25678,N_22702,N_23300);
nor U25679 (N_25679,N_24334,N_23157);
or U25680 (N_25680,N_24547,N_24805);
or U25681 (N_25681,N_24391,N_24204);
and U25682 (N_25682,N_24804,N_24580);
or U25683 (N_25683,N_24110,N_24996);
and U25684 (N_25684,N_23967,N_22588);
nor U25685 (N_25685,N_22515,N_24739);
nand U25686 (N_25686,N_24618,N_24942);
xor U25687 (N_25687,N_23137,N_23033);
xor U25688 (N_25688,N_24581,N_24367);
or U25689 (N_25689,N_24308,N_24128);
or U25690 (N_25690,N_23567,N_23228);
xor U25691 (N_25691,N_23384,N_22717);
xnor U25692 (N_25692,N_23078,N_23345);
and U25693 (N_25693,N_23793,N_23606);
nand U25694 (N_25694,N_23024,N_24648);
nand U25695 (N_25695,N_22569,N_22779);
xnor U25696 (N_25696,N_24303,N_24390);
nor U25697 (N_25697,N_24494,N_23073);
and U25698 (N_25698,N_23672,N_24115);
xor U25699 (N_25699,N_24974,N_24780);
nor U25700 (N_25700,N_23272,N_22730);
nand U25701 (N_25701,N_23118,N_23334);
and U25702 (N_25702,N_23904,N_24437);
xor U25703 (N_25703,N_23641,N_24616);
nor U25704 (N_25704,N_24077,N_23124);
or U25705 (N_25705,N_24912,N_24955);
xor U25706 (N_25706,N_24072,N_24963);
nor U25707 (N_25707,N_23865,N_23079);
xor U25708 (N_25708,N_22513,N_23795);
nor U25709 (N_25709,N_22919,N_24692);
nand U25710 (N_25710,N_23615,N_23469);
nor U25711 (N_25711,N_22835,N_23030);
and U25712 (N_25712,N_23181,N_24980);
nor U25713 (N_25713,N_23656,N_24254);
and U25714 (N_25714,N_23903,N_24995);
and U25715 (N_25715,N_24659,N_22605);
xnor U25716 (N_25716,N_24478,N_22688);
and U25717 (N_25717,N_24079,N_22746);
xor U25718 (N_25718,N_24221,N_23183);
and U25719 (N_25719,N_24744,N_24854);
or U25720 (N_25720,N_24876,N_23909);
xnor U25721 (N_25721,N_24219,N_24823);
xor U25722 (N_25722,N_24312,N_23950);
and U25723 (N_25723,N_24251,N_24297);
and U25724 (N_25724,N_24332,N_24945);
xor U25725 (N_25725,N_24322,N_24762);
xnor U25726 (N_25726,N_23270,N_22962);
nor U25727 (N_25727,N_23450,N_24296);
nand U25728 (N_25728,N_24643,N_24142);
xor U25729 (N_25729,N_22638,N_24024);
or U25730 (N_25730,N_24693,N_23303);
nor U25731 (N_25731,N_24926,N_24435);
nor U25732 (N_25732,N_24263,N_24860);
nand U25733 (N_25733,N_23185,N_23105);
nor U25734 (N_25734,N_23693,N_24528);
or U25735 (N_25735,N_23604,N_24310);
nor U25736 (N_25736,N_22953,N_23490);
or U25737 (N_25737,N_23934,N_22795);
and U25738 (N_25738,N_24164,N_22507);
nand U25739 (N_25739,N_23431,N_23661);
nand U25740 (N_25740,N_23408,N_23245);
and U25741 (N_25741,N_23008,N_23222);
nor U25742 (N_25742,N_22748,N_23371);
and U25743 (N_25743,N_24938,N_24919);
and U25744 (N_25744,N_24933,N_23081);
nor U25745 (N_25745,N_24895,N_23082);
or U25746 (N_25746,N_24787,N_24572);
nor U25747 (N_25747,N_23260,N_23484);
xnor U25748 (N_25748,N_23344,N_23572);
and U25749 (N_25749,N_24318,N_24202);
nand U25750 (N_25750,N_24923,N_24754);
nand U25751 (N_25751,N_23603,N_22755);
nor U25752 (N_25752,N_24878,N_23299);
nand U25753 (N_25753,N_22908,N_23496);
nand U25754 (N_25754,N_22791,N_24520);
and U25755 (N_25755,N_24841,N_23992);
nand U25756 (N_25756,N_24561,N_24654);
or U25757 (N_25757,N_24781,N_24989);
or U25758 (N_25758,N_24776,N_23901);
nor U25759 (N_25759,N_24535,N_23726);
and U25760 (N_25760,N_24940,N_24455);
xnor U25761 (N_25761,N_24369,N_23143);
or U25762 (N_25762,N_24071,N_23220);
nand U25763 (N_25763,N_22589,N_24004);
nor U25764 (N_25764,N_22587,N_23467);
nor U25765 (N_25765,N_23447,N_23050);
nand U25766 (N_25766,N_23939,N_23942);
nor U25767 (N_25767,N_23536,N_23400);
or U25768 (N_25768,N_23214,N_24889);
or U25769 (N_25769,N_24505,N_23841);
nand U25770 (N_25770,N_23749,N_23320);
nor U25771 (N_25771,N_22600,N_23346);
and U25772 (N_25772,N_24326,N_23900);
nor U25773 (N_25773,N_23772,N_23878);
xnor U25774 (N_25774,N_23912,N_23172);
nand U25775 (N_25775,N_24571,N_22561);
and U25776 (N_25776,N_22662,N_24075);
xor U25777 (N_25777,N_24699,N_24877);
xor U25778 (N_25778,N_24266,N_24291);
nor U25779 (N_25779,N_24393,N_22803);
or U25780 (N_25780,N_23497,N_24154);
or U25781 (N_25781,N_22608,N_23890);
nand U25782 (N_25782,N_23760,N_23421);
nor U25783 (N_25783,N_22902,N_22880);
xor U25784 (N_25784,N_22946,N_23018);
nand U25785 (N_25785,N_22948,N_24875);
nand U25786 (N_25786,N_24387,N_23665);
nor U25787 (N_25787,N_24716,N_23200);
or U25788 (N_25788,N_23337,N_23296);
or U25789 (N_25789,N_24143,N_23991);
xnor U25790 (N_25790,N_22625,N_24458);
nand U25791 (N_25791,N_23918,N_22514);
and U25792 (N_25792,N_22739,N_24022);
xnor U25793 (N_25793,N_23696,N_24403);
or U25794 (N_25794,N_23131,N_24961);
nand U25795 (N_25795,N_23263,N_22682);
nor U25796 (N_25796,N_24928,N_23403);
xor U25797 (N_25797,N_23856,N_24833);
and U25798 (N_25798,N_24609,N_23324);
nand U25799 (N_25799,N_24205,N_23479);
nor U25800 (N_25800,N_24434,N_24136);
or U25801 (N_25801,N_24936,N_24465);
or U25802 (N_25802,N_23802,N_24819);
or U25803 (N_25803,N_23107,N_22502);
nand U25804 (N_25804,N_22620,N_23718);
or U25805 (N_25805,N_22796,N_24400);
xnor U25806 (N_25806,N_24031,N_23897);
and U25807 (N_25807,N_23522,N_23076);
xnor U25808 (N_25808,N_23662,N_23012);
and U25809 (N_25809,N_23885,N_23554);
xor U25810 (N_25810,N_23215,N_24550);
and U25811 (N_25811,N_23342,N_22741);
nand U25812 (N_25812,N_23433,N_24168);
nor U25813 (N_25813,N_24663,N_22567);
xor U25814 (N_25814,N_24577,N_22856);
and U25815 (N_25815,N_23963,N_23243);
or U25816 (N_25816,N_24567,N_23227);
xnor U25817 (N_25817,N_22684,N_23254);
and U25818 (N_25818,N_24225,N_23511);
nand U25819 (N_25819,N_22899,N_23392);
nand U25820 (N_25820,N_23844,N_24487);
nor U25821 (N_25821,N_24472,N_24882);
nor U25822 (N_25822,N_23945,N_24946);
xor U25823 (N_25823,N_24684,N_24145);
nand U25824 (N_25824,N_22750,N_22789);
and U25825 (N_25825,N_24349,N_23316);
and U25826 (N_25826,N_22610,N_22548);
and U25827 (N_25827,N_23060,N_23405);
or U25828 (N_25828,N_22681,N_23837);
nand U25829 (N_25829,N_23575,N_24731);
nor U25830 (N_25830,N_23736,N_23610);
and U25831 (N_25831,N_23475,N_24870);
nand U25832 (N_25832,N_24582,N_23009);
nor U25833 (N_25833,N_24006,N_22756);
xnor U25834 (N_25834,N_24108,N_23799);
and U25835 (N_25835,N_24402,N_22503);
and U25836 (N_25836,N_23883,N_23938);
nand U25837 (N_25837,N_24863,N_22904);
nor U25838 (N_25838,N_23689,N_24704);
xnor U25839 (N_25839,N_24081,N_23231);
nor U25840 (N_25840,N_24743,N_24517);
and U25841 (N_25841,N_24767,N_24523);
xnor U25842 (N_25842,N_23990,N_24856);
xnor U25843 (N_25843,N_23558,N_24406);
and U25844 (N_25844,N_23106,N_24092);
and U25845 (N_25845,N_22669,N_22628);
or U25846 (N_25846,N_23418,N_22582);
and U25847 (N_25847,N_22851,N_22720);
and U25848 (N_25848,N_24661,N_24323);
and U25849 (N_25849,N_22782,N_22761);
or U25850 (N_25850,N_24147,N_22869);
or U25851 (N_25851,N_23481,N_22619);
and U25852 (N_25852,N_24924,N_24588);
or U25853 (N_25853,N_22640,N_23624);
or U25854 (N_25854,N_24894,N_24104);
nor U25855 (N_25855,N_24736,N_23027);
nor U25856 (N_25856,N_23365,N_23639);
nand U25857 (N_25857,N_22875,N_23360);
and U25858 (N_25858,N_22927,N_24737);
nor U25859 (N_25859,N_23649,N_23301);
or U25860 (N_25860,N_23150,N_22501);
nand U25861 (N_25861,N_23500,N_22788);
xor U25862 (N_25862,N_24207,N_24179);
or U25863 (N_25863,N_23840,N_23808);
xnor U25864 (N_25864,N_23612,N_24488);
or U25865 (N_25865,N_24579,N_23240);
or U25866 (N_25866,N_23864,N_23617);
nand U25867 (N_25867,N_23559,N_23217);
nor U25868 (N_25868,N_22597,N_23956);
and U25869 (N_25869,N_22517,N_22818);
xnor U25870 (N_25870,N_22895,N_23241);
nand U25871 (N_25871,N_24118,N_23116);
nand U25872 (N_25872,N_24987,N_23383);
nand U25873 (N_25873,N_23202,N_22817);
and U25874 (N_25874,N_23251,N_23439);
and U25875 (N_25875,N_23153,N_22670);
nor U25876 (N_25876,N_24807,N_24820);
xor U25877 (N_25877,N_22977,N_22557);
nand U25878 (N_25878,N_23064,N_24673);
xor U25879 (N_25879,N_24752,N_24703);
and U25880 (N_25880,N_24761,N_24474);
or U25881 (N_25881,N_23966,N_24389);
nor U25882 (N_25882,N_23806,N_24893);
xnor U25883 (N_25883,N_24252,N_24002);
xnor U25884 (N_25884,N_24975,N_24610);
and U25885 (N_25885,N_23196,N_24253);
or U25886 (N_25886,N_24027,N_23095);
nor U25887 (N_25887,N_22749,N_24897);
nor U25888 (N_25888,N_24184,N_23412);
nor U25889 (N_25889,N_23289,N_23546);
or U25890 (N_25890,N_24840,N_24038);
or U25891 (N_25891,N_23695,N_24070);
and U25892 (N_25892,N_24645,N_24544);
and U25893 (N_25893,N_23631,N_22598);
or U25894 (N_25894,N_22518,N_24702);
and U25895 (N_25895,N_22827,N_24783);
nand U25896 (N_25896,N_23492,N_23399);
nand U25897 (N_25897,N_23902,N_23895);
nand U25898 (N_25898,N_23565,N_24111);
nand U25899 (N_25899,N_24394,N_24599);
nor U25900 (N_25900,N_22559,N_24937);
nand U25901 (N_25901,N_24971,N_24515);
nor U25902 (N_25902,N_23826,N_23932);
nand U25903 (N_25903,N_24966,N_22767);
xnor U25904 (N_25904,N_23191,N_22544);
or U25905 (N_25905,N_23349,N_23119);
nand U25906 (N_25906,N_24868,N_23527);
and U25907 (N_25907,N_23438,N_22826);
nor U25908 (N_25908,N_24043,N_24977);
and U25909 (N_25909,N_23635,N_22983);
and U25910 (N_25910,N_24724,N_23209);
xor U25911 (N_25911,N_24341,N_23861);
nand U25912 (N_25912,N_24084,N_23444);
and U25913 (N_25913,N_24374,N_23703);
or U25914 (N_25914,N_23207,N_22855);
or U25915 (N_25915,N_22576,N_24203);
xor U25916 (N_25916,N_24812,N_24000);
and U25917 (N_25917,N_23915,N_24583);
nand U25918 (N_25918,N_24538,N_23333);
nor U25919 (N_25919,N_24636,N_24218);
nor U25920 (N_25920,N_24672,N_24244);
nand U25921 (N_25921,N_24838,N_24351);
nand U25922 (N_25922,N_23504,N_22954);
nand U25923 (N_25923,N_24524,N_22694);
and U25924 (N_25924,N_23147,N_22511);
or U25925 (N_25925,N_23168,N_23487);
or U25926 (N_25926,N_23576,N_24867);
nor U25927 (N_25927,N_22525,N_23589);
nand U25928 (N_25928,N_23516,N_24959);
or U25929 (N_25929,N_24836,N_22828);
xnor U25930 (N_25930,N_24796,N_23788);
nand U25931 (N_25931,N_23537,N_24383);
nor U25932 (N_25932,N_23679,N_24960);
nor U25933 (N_25933,N_23701,N_24080);
xor U25934 (N_25934,N_23754,N_23362);
nand U25935 (N_25935,N_24195,N_24335);
xnor U25936 (N_25936,N_23048,N_22879);
nor U25937 (N_25937,N_22780,N_23732);
nor U25938 (N_25938,N_24056,N_22911);
xor U25939 (N_25939,N_23180,N_23443);
nand U25940 (N_25940,N_23442,N_24085);
nor U25941 (N_25941,N_23308,N_24563);
or U25942 (N_25942,N_23077,N_24768);
nand U25943 (N_25943,N_22897,N_23380);
or U25944 (N_25944,N_24508,N_24829);
xnor U25945 (N_25945,N_24150,N_23135);
nand U25946 (N_25946,N_22633,N_23706);
xnor U25947 (N_25947,N_24597,N_22583);
xor U25948 (N_25948,N_24448,N_24176);
xnor U25949 (N_25949,N_23765,N_24985);
nand U25950 (N_25950,N_23704,N_24990);
nor U25951 (N_25951,N_22558,N_23229);
and U25952 (N_25952,N_22932,N_23186);
nor U25953 (N_25953,N_24738,N_23387);
nor U25954 (N_25954,N_23032,N_24824);
nand U25955 (N_25955,N_23184,N_24097);
xor U25956 (N_25956,N_23052,N_23508);
nand U25957 (N_25957,N_23744,N_22859);
and U25958 (N_25958,N_24255,N_22570);
xnor U25959 (N_25959,N_23142,N_23329);
and U25960 (N_25960,N_24917,N_22585);
and U25961 (N_25961,N_24300,N_24330);
or U25962 (N_25962,N_22882,N_23650);
nand U25963 (N_25963,N_23425,N_22836);
xor U25964 (N_25964,N_24799,N_23978);
or U25965 (N_25965,N_23836,N_24213);
nor U25966 (N_25966,N_23951,N_24425);
xnor U25967 (N_25967,N_22763,N_24617);
xnor U25968 (N_25968,N_23098,N_23917);
nor U25969 (N_25969,N_24865,N_22538);
or U25970 (N_25970,N_23614,N_24160);
nor U25971 (N_25971,N_23834,N_23452);
or U25972 (N_25972,N_24712,N_23159);
nand U25973 (N_25973,N_24930,N_24162);
nor U25974 (N_25974,N_23862,N_22987);
or U25975 (N_25975,N_24279,N_23705);
xor U25976 (N_25976,N_24557,N_22692);
nor U25977 (N_25977,N_23700,N_23356);
nor U25978 (N_25978,N_22849,N_24444);
and U25979 (N_25979,N_23764,N_24373);
and U25980 (N_25980,N_24480,N_22744);
xnor U25981 (N_25981,N_22577,N_24881);
nor U25982 (N_25982,N_23593,N_22655);
nand U25983 (N_25983,N_24301,N_23605);
and U25984 (N_25984,N_24438,N_23586);
nor U25985 (N_25985,N_24717,N_22648);
and U25986 (N_25986,N_23197,N_23505);
nor U25987 (N_25987,N_23630,N_24485);
or U25988 (N_25988,N_24242,N_22771);
xnor U25989 (N_25989,N_23850,N_24746);
xnor U25990 (N_25990,N_23579,N_23971);
or U25991 (N_25991,N_24029,N_24857);
xor U25992 (N_25992,N_24952,N_23707);
nor U25993 (N_25993,N_23933,N_24885);
or U25994 (N_25994,N_24916,N_23876);
nor U25995 (N_25995,N_22881,N_24283);
or U25996 (N_25996,N_24678,N_23609);
nor U25997 (N_25997,N_24711,N_22804);
or U25998 (N_25998,N_23874,N_23427);
nand U25999 (N_25999,N_23178,N_24496);
nand U26000 (N_26000,N_23236,N_24453);
xor U26001 (N_26001,N_24718,N_22594);
or U26002 (N_26002,N_23049,N_22787);
xnor U26003 (N_26003,N_22713,N_24011);
and U26004 (N_26004,N_24058,N_24790);
and U26005 (N_26005,N_23538,N_23734);
xor U26006 (N_26006,N_22677,N_24827);
xnor U26007 (N_26007,N_23814,N_22626);
or U26008 (N_26008,N_24172,N_23599);
or U26009 (N_26009,N_24068,N_23783);
and U26010 (N_26010,N_22536,N_24555);
xor U26011 (N_26011,N_23366,N_24956);
or U26012 (N_26012,N_24113,N_24050);
nand U26013 (N_26013,N_23255,N_24355);
xnor U26014 (N_26014,N_23780,N_23540);
or U26015 (N_26015,N_24747,N_22905);
nor U26016 (N_26016,N_24146,N_23156);
nand U26017 (N_26017,N_24171,N_23028);
or U26018 (N_26018,N_23592,N_23295);
nor U26019 (N_26019,N_22921,N_23370);
xnor U26020 (N_26020,N_23374,N_23464);
nand U26021 (N_26021,N_22601,N_23331);
xor U26022 (N_26022,N_24835,N_24549);
and U26023 (N_26023,N_22718,N_23080);
nand U26024 (N_26024,N_24298,N_22774);
nor U26025 (N_26025,N_22607,N_22509);
nand U26026 (N_26026,N_23451,N_22614);
nand U26027 (N_26027,N_22528,N_23278);
nor U26028 (N_26028,N_22757,N_22540);
nand U26029 (N_26029,N_23166,N_22850);
nand U26030 (N_26030,N_24216,N_23164);
nand U26031 (N_26031,N_23176,N_24450);
xnor U26032 (N_26032,N_24600,N_22988);
xnor U26033 (N_26033,N_24522,N_23688);
nand U26034 (N_26034,N_23677,N_24647);
nand U26035 (N_26035,N_24532,N_23843);
nor U26036 (N_26036,N_23638,N_24235);
nand U26037 (N_26037,N_23066,N_24751);
and U26038 (N_26038,N_24626,N_23478);
and U26039 (N_26039,N_24331,N_24139);
and U26040 (N_26040,N_23089,N_23621);
or U26041 (N_26041,N_24593,N_23163);
xnor U26042 (N_26042,N_24696,N_23535);
nor U26043 (N_26043,N_23208,N_23242);
nand U26044 (N_26044,N_23669,N_23634);
and U26045 (N_26045,N_22814,N_22510);
nand U26046 (N_26046,N_24775,N_24939);
and U26047 (N_26047,N_23715,N_23204);
xnor U26048 (N_26048,N_23160,N_24915);
or U26049 (N_26049,N_23880,N_24698);
nor U26050 (N_26050,N_22674,N_24345);
xnor U26051 (N_26051,N_24976,N_23507);
or U26052 (N_26052,N_23564,N_24690);
and U26053 (N_26053,N_22765,N_24683);
nand U26054 (N_26054,N_23860,N_23645);
xnor U26055 (N_26055,N_22747,N_24905);
xnor U26056 (N_26056,N_24707,N_24957);
and U26057 (N_26057,N_23673,N_24749);
and U26058 (N_26058,N_23563,N_23756);
nand U26059 (N_26059,N_22891,N_24057);
nor U26060 (N_26060,N_24486,N_22687);
nor U26061 (N_26061,N_24655,N_23811);
and U26062 (N_26062,N_24858,N_23681);
or U26063 (N_26063,N_24708,N_22820);
nor U26064 (N_26064,N_24339,N_23637);
and U26065 (N_26065,N_22731,N_23766);
and U26066 (N_26066,N_24144,N_23682);
xor U26067 (N_26067,N_24105,N_24234);
or U26068 (N_26068,N_23219,N_24327);
xnor U26069 (N_26069,N_24287,N_24925);
and U26070 (N_26070,N_23922,N_24590);
or U26071 (N_26071,N_24539,N_24120);
or U26072 (N_26072,N_23867,N_24173);
nor U26073 (N_26073,N_23884,N_22563);
xor U26074 (N_26074,N_23913,N_23961);
or U26075 (N_26075,N_24270,N_23413);
nand U26076 (N_26076,N_24892,N_22723);
nand U26077 (N_26077,N_24551,N_22913);
xor U26078 (N_26078,N_23108,N_23831);
nand U26079 (N_26079,N_23528,N_23031);
or U26080 (N_26080,N_24570,N_23919);
and U26081 (N_26081,N_23377,N_23244);
xor U26082 (N_26082,N_23053,N_24224);
or U26083 (N_26083,N_24611,N_24153);
xor U26084 (N_26084,N_24107,N_23463);
xor U26085 (N_26085,N_24412,N_24639);
and U26086 (N_26086,N_23355,N_23409);
xnor U26087 (N_26087,N_23406,N_24269);
nor U26088 (N_26088,N_22701,N_24784);
nand U26089 (N_26089,N_24890,N_23896);
and U26090 (N_26090,N_24447,N_23393);
nor U26091 (N_26091,N_24568,N_22841);
or U26092 (N_26092,N_23735,N_22816);
or U26093 (N_26093,N_22966,N_24260);
and U26094 (N_26094,N_23973,N_24529);
or U26095 (N_26095,N_24602,N_24540);
or U26096 (N_26096,N_24193,N_23809);
nor U26097 (N_26097,N_23057,N_22539);
nand U26098 (N_26098,N_24822,N_23483);
xor U26099 (N_26099,N_23619,N_22926);
and U26100 (N_26100,N_22580,N_23127);
or U26101 (N_26101,N_23104,N_24159);
or U26102 (N_26102,N_23755,N_22794);
and U26103 (N_26103,N_23763,N_24631);
nor U26104 (N_26104,N_23174,N_24032);
and U26105 (N_26105,N_23899,N_24243);
nand U26106 (N_26106,N_24155,N_23710);
nand U26107 (N_26107,N_23652,N_22722);
nor U26108 (N_26108,N_24197,N_22915);
and U26109 (N_26109,N_24198,N_24669);
or U26110 (N_26110,N_22568,N_22710);
xnor U26111 (N_26111,N_24511,N_23739);
and U26112 (N_26112,N_23985,N_22935);
nand U26113 (N_26113,N_22993,N_22725);
nor U26114 (N_26114,N_24280,N_24797);
nor U26115 (N_26115,N_22799,N_24733);
nor U26116 (N_26116,N_24267,N_24958);
and U26117 (N_26117,N_23737,N_24700);
xor U26118 (N_26118,N_24041,N_24076);
nor U26119 (N_26119,N_22933,N_24317);
xor U26120 (N_26120,N_22612,N_23014);
nand U26121 (N_26121,N_22676,N_24272);
or U26122 (N_26122,N_22596,N_23629);
nor U26123 (N_26123,N_23230,N_23394);
nand U26124 (N_26124,N_23177,N_23372);
nor U26125 (N_26125,N_23851,N_22575);
xnor U26126 (N_26126,N_23065,N_23947);
nand U26127 (N_26127,N_22837,N_23343);
xor U26128 (N_26128,N_22657,N_24112);
and U26129 (N_26129,N_23420,N_24495);
nor U26130 (N_26130,N_24340,N_24404);
and U26131 (N_26131,N_23110,N_24066);
and U26132 (N_26132,N_23087,N_23779);
nand U26133 (N_26133,N_23964,N_23284);
nor U26134 (N_26134,N_22956,N_23021);
and U26135 (N_26135,N_24489,N_22764);
xor U26136 (N_26136,N_24419,N_24705);
nor U26137 (N_26137,N_22906,N_23835);
nor U26138 (N_26138,N_22745,N_22524);
and U26139 (N_26139,N_23002,N_23872);
and U26140 (N_26140,N_22549,N_23955);
nor U26141 (N_26141,N_23530,N_24714);
nand U26142 (N_26142,N_24687,N_23493);
nor U26143 (N_26143,N_24891,N_23773);
nor U26144 (N_26144,N_24914,N_24641);
or U26145 (N_26145,N_23273,N_23620);
nor U26146 (N_26146,N_24424,N_23513);
nor U26147 (N_26147,N_24476,N_22866);
or U26148 (N_26148,N_24329,N_23914);
or U26149 (N_26149,N_22543,N_23205);
and U26150 (N_26150,N_22664,N_22737);
nor U26151 (N_26151,N_22698,N_24769);
nand U26152 (N_26152,N_24343,N_24788);
xnor U26153 (N_26153,N_23597,N_23045);
nand U26154 (N_26154,N_23798,N_24992);
nor U26155 (N_26155,N_24052,N_22815);
and U26156 (N_26156,N_23792,N_24012);
nor U26157 (N_26157,N_23999,N_22971);
and U26158 (N_26158,N_23382,N_23070);
nor U26159 (N_26159,N_24223,N_24358);
and U26160 (N_26160,N_24587,N_22985);
nor U26161 (N_26161,N_23937,N_24372);
nor U26162 (N_26162,N_23583,N_23733);
nor U26163 (N_26163,N_22603,N_24180);
nor U26164 (N_26164,N_23503,N_24217);
xor U26165 (N_26165,N_23088,N_23627);
xor U26166 (N_26166,N_24134,N_22711);
xor U26167 (N_26167,N_23607,N_22566);
and U26168 (N_26168,N_22944,N_24131);
xnor U26169 (N_26169,N_23825,N_24573);
nor U26170 (N_26170,N_24758,N_24800);
or U26171 (N_26171,N_24156,N_23036);
xor U26172 (N_26172,N_23276,N_22516);
or U26173 (N_26173,N_23981,N_24457);
or U26174 (N_26174,N_23680,N_24638);
nor U26175 (N_26175,N_24037,N_22595);
or U26176 (N_26176,N_24017,N_24285);
xor U26177 (N_26177,N_23714,N_24045);
or U26178 (N_26178,N_23584,N_23818);
xnor U26179 (N_26179,N_23378,N_23794);
xnor U26180 (N_26180,N_22830,N_23521);
nand U26181 (N_26181,N_23678,N_24371);
nand U26182 (N_26182,N_23952,N_24185);
nor U26183 (N_26183,N_23155,N_23335);
or U26184 (N_26184,N_24018,N_24973);
nor U26185 (N_26185,N_23395,N_23161);
xor U26186 (N_26186,N_24064,N_22768);
xor U26187 (N_26187,N_24671,N_24175);
and U26188 (N_26188,N_22833,N_23523);
nand U26189 (N_26189,N_24366,N_24449);
nand U26190 (N_26190,N_23713,N_23311);
nor U26191 (N_26191,N_24314,N_23748);
xor U26192 (N_26192,N_24440,N_23771);
nand U26193 (N_26193,N_22888,N_23866);
xnor U26194 (N_26194,N_23768,N_24991);
and U26195 (N_26195,N_23691,N_23212);
xnor U26196 (N_26196,N_22823,N_24035);
nor U26197 (N_26197,N_22994,N_23694);
or U26198 (N_26198,N_24773,N_24927);
nand U26199 (N_26199,N_23257,N_23845);
nand U26200 (N_26200,N_23671,N_23149);
nor U26201 (N_26201,N_23437,N_23472);
xor U26202 (N_26202,N_24005,N_24605);
or U26203 (N_26203,N_24069,N_24552);
and U26204 (N_26204,N_23868,N_22846);
nor U26205 (N_26205,N_24886,N_23960);
nor U26206 (N_26206,N_23322,N_22521);
and U26207 (N_26207,N_24257,N_23711);
xor U26208 (N_26208,N_22957,N_23921);
nand U26209 (N_26209,N_23817,N_23791);
nand U26210 (N_26210,N_22651,N_24518);
and U26211 (N_26211,N_24044,N_23390);
and U26212 (N_26212,N_22733,N_23882);
xor U26213 (N_26213,N_24432,N_24483);
and U26214 (N_26214,N_24170,N_22784);
and U26215 (N_26215,N_24445,N_24088);
nand U26216 (N_26216,N_23139,N_23954);
nand U26217 (N_26217,N_23199,N_24187);
and U26218 (N_26218,N_23801,N_24740);
nor U26219 (N_26219,N_22896,N_24596);
nor U26220 (N_26220,N_24935,N_23470);
xor U26221 (N_26221,N_24745,N_23218);
nand U26222 (N_26222,N_22867,N_23602);
xnor U26223 (N_26223,N_24313,N_24046);
and U26224 (N_26224,N_23171,N_23822);
xor U26225 (N_26225,N_22938,N_24514);
and U26226 (N_26226,N_23422,N_23259);
and U26227 (N_26227,N_22848,N_22907);
nand U26228 (N_26228,N_22671,N_24688);
or U26229 (N_26229,N_23111,N_24344);
xor U26230 (N_26230,N_24292,N_23520);
nor U26231 (N_26231,N_24227,N_24765);
nor U26232 (N_26232,N_22553,N_24328);
nand U26233 (N_26233,N_23517,N_24421);
xnor U26234 (N_26234,N_23055,N_24395);
nor U26235 (N_26235,N_22943,N_24127);
nor U26236 (N_26236,N_24354,N_22950);
nor U26237 (N_26237,N_23907,N_22893);
or U26238 (N_26238,N_22868,N_24948);
nor U26239 (N_26239,N_23533,N_22964);
xor U26240 (N_26240,N_22930,N_24278);
nor U26241 (N_26241,N_23122,N_22584);
nor U26242 (N_26242,N_24500,N_23455);
nand U26243 (N_26243,N_23182,N_23195);
nor U26244 (N_26244,N_23038,N_23643);
nor U26245 (N_26245,N_24246,N_24832);
nor U26246 (N_26246,N_23063,N_23462);
nand U26247 (N_26247,N_24901,N_23640);
xnor U26248 (N_26248,N_23213,N_24174);
or U26249 (N_26249,N_22937,N_24019);
or U26250 (N_26250,N_23926,N_23948);
and U26251 (N_26251,N_22910,N_22922);
xnor U26252 (N_26252,N_22939,N_22820);
nand U26253 (N_26253,N_22719,N_23960);
xnor U26254 (N_26254,N_24743,N_23047);
xnor U26255 (N_26255,N_23895,N_22548);
or U26256 (N_26256,N_24495,N_24317);
xnor U26257 (N_26257,N_23285,N_22662);
nand U26258 (N_26258,N_24893,N_23648);
and U26259 (N_26259,N_23448,N_24263);
xor U26260 (N_26260,N_24955,N_22607);
nand U26261 (N_26261,N_23614,N_23339);
or U26262 (N_26262,N_22665,N_22825);
and U26263 (N_26263,N_24238,N_23757);
xor U26264 (N_26264,N_22866,N_23309);
xor U26265 (N_26265,N_24743,N_24273);
and U26266 (N_26266,N_22919,N_24600);
or U26267 (N_26267,N_24839,N_23799);
or U26268 (N_26268,N_24786,N_24168);
and U26269 (N_26269,N_23155,N_22896);
nor U26270 (N_26270,N_23750,N_24571);
and U26271 (N_26271,N_24057,N_22595);
and U26272 (N_26272,N_23767,N_23808);
xnor U26273 (N_26273,N_23416,N_24153);
xor U26274 (N_26274,N_24905,N_23003);
nor U26275 (N_26275,N_24662,N_24961);
or U26276 (N_26276,N_24739,N_24204);
nor U26277 (N_26277,N_23308,N_24167);
and U26278 (N_26278,N_22745,N_23702);
nor U26279 (N_26279,N_23940,N_23401);
xnor U26280 (N_26280,N_22741,N_24158);
and U26281 (N_26281,N_24474,N_23950);
and U26282 (N_26282,N_24091,N_23330);
and U26283 (N_26283,N_22680,N_23624);
or U26284 (N_26284,N_24150,N_23560);
and U26285 (N_26285,N_23223,N_23668);
xnor U26286 (N_26286,N_24948,N_24498);
xor U26287 (N_26287,N_22950,N_23498);
or U26288 (N_26288,N_24300,N_23293);
and U26289 (N_26289,N_24792,N_23889);
xor U26290 (N_26290,N_22582,N_23636);
xor U26291 (N_26291,N_23473,N_22517);
nor U26292 (N_26292,N_24630,N_22827);
nand U26293 (N_26293,N_22528,N_23178);
xnor U26294 (N_26294,N_23217,N_23010);
or U26295 (N_26295,N_22597,N_24650);
and U26296 (N_26296,N_23492,N_23148);
and U26297 (N_26297,N_23306,N_23928);
and U26298 (N_26298,N_24083,N_22603);
xor U26299 (N_26299,N_24398,N_23350);
and U26300 (N_26300,N_24519,N_24797);
xnor U26301 (N_26301,N_23703,N_24799);
nand U26302 (N_26302,N_22590,N_23790);
and U26303 (N_26303,N_23365,N_23475);
nand U26304 (N_26304,N_24024,N_24363);
and U26305 (N_26305,N_24971,N_24289);
nor U26306 (N_26306,N_23537,N_23692);
and U26307 (N_26307,N_24383,N_24718);
nor U26308 (N_26308,N_23902,N_23486);
or U26309 (N_26309,N_24676,N_23307);
nor U26310 (N_26310,N_22999,N_23767);
nor U26311 (N_26311,N_24211,N_24967);
nor U26312 (N_26312,N_24675,N_24063);
xor U26313 (N_26313,N_24943,N_24014);
xor U26314 (N_26314,N_23285,N_23907);
or U26315 (N_26315,N_23467,N_22515);
xnor U26316 (N_26316,N_24371,N_24288);
or U26317 (N_26317,N_22674,N_23953);
nor U26318 (N_26318,N_22982,N_22695);
or U26319 (N_26319,N_23529,N_22802);
and U26320 (N_26320,N_22839,N_23684);
and U26321 (N_26321,N_22777,N_24741);
xor U26322 (N_26322,N_24071,N_24237);
nor U26323 (N_26323,N_22583,N_23820);
nor U26324 (N_26324,N_24041,N_22969);
and U26325 (N_26325,N_24972,N_24883);
nor U26326 (N_26326,N_23052,N_23235);
nand U26327 (N_26327,N_23416,N_24115);
and U26328 (N_26328,N_22818,N_23905);
nand U26329 (N_26329,N_24515,N_24942);
nor U26330 (N_26330,N_23772,N_24696);
nand U26331 (N_26331,N_23406,N_24050);
nand U26332 (N_26332,N_23395,N_22863);
nor U26333 (N_26333,N_23484,N_24998);
nor U26334 (N_26334,N_24473,N_24024);
nor U26335 (N_26335,N_23590,N_23496);
nand U26336 (N_26336,N_24086,N_24083);
or U26337 (N_26337,N_23792,N_22685);
and U26338 (N_26338,N_23695,N_24739);
and U26339 (N_26339,N_24306,N_23590);
nor U26340 (N_26340,N_22858,N_24437);
or U26341 (N_26341,N_24460,N_23605);
xor U26342 (N_26342,N_22677,N_24208);
xor U26343 (N_26343,N_24085,N_24439);
xnor U26344 (N_26344,N_24366,N_24597);
nor U26345 (N_26345,N_24734,N_22995);
nand U26346 (N_26346,N_23328,N_23219);
or U26347 (N_26347,N_23261,N_23791);
or U26348 (N_26348,N_23157,N_23988);
or U26349 (N_26349,N_23827,N_23094);
xor U26350 (N_26350,N_23040,N_22563);
and U26351 (N_26351,N_24640,N_22544);
nand U26352 (N_26352,N_24381,N_23649);
xor U26353 (N_26353,N_24176,N_24101);
nand U26354 (N_26354,N_23463,N_23443);
and U26355 (N_26355,N_24965,N_23433);
nor U26356 (N_26356,N_24988,N_24173);
or U26357 (N_26357,N_24908,N_23190);
nand U26358 (N_26358,N_24226,N_23613);
nor U26359 (N_26359,N_22620,N_23610);
xnor U26360 (N_26360,N_24925,N_22551);
xnor U26361 (N_26361,N_22754,N_22847);
nor U26362 (N_26362,N_24209,N_22768);
and U26363 (N_26363,N_24329,N_24079);
nor U26364 (N_26364,N_24511,N_24371);
nor U26365 (N_26365,N_23609,N_24789);
and U26366 (N_26366,N_23857,N_23843);
nor U26367 (N_26367,N_23851,N_23621);
nor U26368 (N_26368,N_23995,N_23774);
nand U26369 (N_26369,N_22609,N_24478);
nor U26370 (N_26370,N_22916,N_23065);
xor U26371 (N_26371,N_23167,N_23159);
xnor U26372 (N_26372,N_23031,N_23867);
nor U26373 (N_26373,N_22604,N_24989);
nand U26374 (N_26374,N_24856,N_23412);
nand U26375 (N_26375,N_23102,N_23594);
xnor U26376 (N_26376,N_24144,N_22867);
nor U26377 (N_26377,N_22805,N_24921);
or U26378 (N_26378,N_24222,N_23358);
nor U26379 (N_26379,N_23890,N_23611);
nand U26380 (N_26380,N_24866,N_23614);
nand U26381 (N_26381,N_23438,N_24679);
nor U26382 (N_26382,N_22690,N_24141);
xor U26383 (N_26383,N_23607,N_24505);
or U26384 (N_26384,N_24530,N_23964);
nand U26385 (N_26385,N_22956,N_24244);
and U26386 (N_26386,N_23637,N_24511);
nor U26387 (N_26387,N_22594,N_24198);
xor U26388 (N_26388,N_23196,N_23563);
xor U26389 (N_26389,N_23575,N_23098);
or U26390 (N_26390,N_23263,N_24285);
xor U26391 (N_26391,N_23265,N_23129);
xor U26392 (N_26392,N_24010,N_24480);
or U26393 (N_26393,N_24370,N_23560);
nand U26394 (N_26394,N_24618,N_22604);
nand U26395 (N_26395,N_24291,N_22759);
nand U26396 (N_26396,N_24306,N_23442);
nor U26397 (N_26397,N_23629,N_23395);
nor U26398 (N_26398,N_23808,N_23229);
nor U26399 (N_26399,N_23776,N_23622);
nor U26400 (N_26400,N_23586,N_22818);
and U26401 (N_26401,N_23161,N_22576);
nor U26402 (N_26402,N_22635,N_23753);
xnor U26403 (N_26403,N_24001,N_23913);
nand U26404 (N_26404,N_24707,N_23915);
xnor U26405 (N_26405,N_23119,N_24258);
or U26406 (N_26406,N_24683,N_24362);
nand U26407 (N_26407,N_22927,N_22948);
and U26408 (N_26408,N_24413,N_23075);
nor U26409 (N_26409,N_22803,N_24347);
nor U26410 (N_26410,N_22782,N_24689);
xor U26411 (N_26411,N_24096,N_22699);
nor U26412 (N_26412,N_22794,N_24262);
nor U26413 (N_26413,N_22828,N_22890);
xor U26414 (N_26414,N_23523,N_23477);
nand U26415 (N_26415,N_22762,N_24376);
or U26416 (N_26416,N_24763,N_24631);
and U26417 (N_26417,N_23255,N_22761);
or U26418 (N_26418,N_22686,N_24640);
nand U26419 (N_26419,N_23400,N_23781);
xor U26420 (N_26420,N_24644,N_23311);
nor U26421 (N_26421,N_23791,N_22888);
nand U26422 (N_26422,N_22829,N_22740);
nand U26423 (N_26423,N_24933,N_22500);
xor U26424 (N_26424,N_24142,N_24939);
xor U26425 (N_26425,N_24825,N_22710);
or U26426 (N_26426,N_24555,N_23236);
nand U26427 (N_26427,N_23488,N_23523);
and U26428 (N_26428,N_23800,N_22768);
and U26429 (N_26429,N_22869,N_23496);
or U26430 (N_26430,N_24397,N_24458);
and U26431 (N_26431,N_24025,N_24902);
xnor U26432 (N_26432,N_23089,N_24906);
nor U26433 (N_26433,N_23458,N_23185);
nand U26434 (N_26434,N_24505,N_23765);
and U26435 (N_26435,N_23892,N_23881);
nand U26436 (N_26436,N_23418,N_24200);
nor U26437 (N_26437,N_23285,N_23591);
and U26438 (N_26438,N_23427,N_24667);
and U26439 (N_26439,N_23442,N_22594);
nor U26440 (N_26440,N_24127,N_24818);
or U26441 (N_26441,N_24171,N_24533);
nor U26442 (N_26442,N_24897,N_22992);
nor U26443 (N_26443,N_22718,N_23897);
xor U26444 (N_26444,N_24563,N_24253);
and U26445 (N_26445,N_24781,N_23653);
or U26446 (N_26446,N_22824,N_22771);
nor U26447 (N_26447,N_23209,N_23179);
nor U26448 (N_26448,N_22822,N_23029);
or U26449 (N_26449,N_22801,N_23038);
nand U26450 (N_26450,N_22512,N_23437);
or U26451 (N_26451,N_23382,N_23991);
nor U26452 (N_26452,N_23050,N_23626);
or U26453 (N_26453,N_22759,N_22836);
xor U26454 (N_26454,N_22697,N_23917);
nand U26455 (N_26455,N_23394,N_22767);
and U26456 (N_26456,N_22956,N_23337);
xnor U26457 (N_26457,N_22930,N_23957);
nor U26458 (N_26458,N_22872,N_22550);
xor U26459 (N_26459,N_23289,N_24646);
nand U26460 (N_26460,N_23638,N_24451);
nor U26461 (N_26461,N_24939,N_23280);
and U26462 (N_26462,N_23167,N_24982);
nor U26463 (N_26463,N_22879,N_24411);
and U26464 (N_26464,N_22969,N_23657);
and U26465 (N_26465,N_24394,N_24118);
xor U26466 (N_26466,N_23941,N_22863);
or U26467 (N_26467,N_24117,N_23494);
nand U26468 (N_26468,N_22667,N_24076);
xor U26469 (N_26469,N_24321,N_23625);
nand U26470 (N_26470,N_24963,N_22562);
xor U26471 (N_26471,N_24288,N_24752);
xor U26472 (N_26472,N_23977,N_24237);
xor U26473 (N_26473,N_24529,N_23110);
nand U26474 (N_26474,N_23140,N_22671);
nor U26475 (N_26475,N_23077,N_23081);
nand U26476 (N_26476,N_23045,N_22600);
or U26477 (N_26477,N_24166,N_22554);
and U26478 (N_26478,N_23383,N_24142);
nor U26479 (N_26479,N_23952,N_22978);
or U26480 (N_26480,N_24941,N_22815);
or U26481 (N_26481,N_23957,N_22713);
or U26482 (N_26482,N_23781,N_24826);
xor U26483 (N_26483,N_22820,N_23289);
or U26484 (N_26484,N_23827,N_24362);
and U26485 (N_26485,N_23247,N_24458);
nor U26486 (N_26486,N_23124,N_22750);
xor U26487 (N_26487,N_24067,N_24266);
and U26488 (N_26488,N_22528,N_24390);
nor U26489 (N_26489,N_24128,N_22779);
nand U26490 (N_26490,N_24989,N_23122);
nand U26491 (N_26491,N_23443,N_23366);
xnor U26492 (N_26492,N_22536,N_24422);
and U26493 (N_26493,N_24842,N_22632);
and U26494 (N_26494,N_24417,N_24039);
xnor U26495 (N_26495,N_24226,N_22842);
nor U26496 (N_26496,N_24937,N_24051);
or U26497 (N_26497,N_23146,N_24139);
and U26498 (N_26498,N_23649,N_23150);
nor U26499 (N_26499,N_24252,N_23777);
and U26500 (N_26500,N_24437,N_24434);
nand U26501 (N_26501,N_24263,N_24927);
nor U26502 (N_26502,N_23544,N_24130);
and U26503 (N_26503,N_23936,N_22890);
nor U26504 (N_26504,N_24003,N_23271);
nor U26505 (N_26505,N_24467,N_23164);
nor U26506 (N_26506,N_23442,N_24225);
and U26507 (N_26507,N_24052,N_23796);
nand U26508 (N_26508,N_23636,N_24420);
nor U26509 (N_26509,N_24875,N_23955);
nor U26510 (N_26510,N_23605,N_23844);
xor U26511 (N_26511,N_23084,N_22991);
xnor U26512 (N_26512,N_23528,N_22636);
or U26513 (N_26513,N_24166,N_23523);
xnor U26514 (N_26514,N_23625,N_24941);
nand U26515 (N_26515,N_23986,N_23271);
and U26516 (N_26516,N_24159,N_24795);
or U26517 (N_26517,N_23503,N_22805);
nor U26518 (N_26518,N_23765,N_23499);
nor U26519 (N_26519,N_24421,N_24522);
xnor U26520 (N_26520,N_24429,N_24284);
or U26521 (N_26521,N_22829,N_23241);
and U26522 (N_26522,N_22526,N_24972);
and U26523 (N_26523,N_23089,N_23660);
and U26524 (N_26524,N_24636,N_22587);
nor U26525 (N_26525,N_24807,N_23759);
or U26526 (N_26526,N_23418,N_22775);
nor U26527 (N_26527,N_23546,N_24230);
xor U26528 (N_26528,N_23132,N_23746);
nand U26529 (N_26529,N_23388,N_22886);
nor U26530 (N_26530,N_24964,N_22616);
or U26531 (N_26531,N_23417,N_24474);
and U26532 (N_26532,N_23786,N_24404);
nor U26533 (N_26533,N_24324,N_22663);
xor U26534 (N_26534,N_23633,N_24696);
nor U26535 (N_26535,N_23249,N_24059);
and U26536 (N_26536,N_23668,N_23881);
nor U26537 (N_26537,N_22828,N_24767);
or U26538 (N_26538,N_22553,N_24223);
xnor U26539 (N_26539,N_22577,N_23395);
nor U26540 (N_26540,N_24633,N_23906);
nor U26541 (N_26541,N_24300,N_22656);
xor U26542 (N_26542,N_22733,N_24881);
nor U26543 (N_26543,N_24221,N_24288);
nor U26544 (N_26544,N_23217,N_24958);
or U26545 (N_26545,N_24370,N_23260);
nor U26546 (N_26546,N_23813,N_24125);
xor U26547 (N_26547,N_23540,N_24821);
nor U26548 (N_26548,N_24285,N_23017);
nor U26549 (N_26549,N_24642,N_23223);
nand U26550 (N_26550,N_23699,N_23850);
nor U26551 (N_26551,N_23882,N_24049);
xor U26552 (N_26552,N_23967,N_23545);
xor U26553 (N_26553,N_24586,N_24322);
and U26554 (N_26554,N_24403,N_23468);
xor U26555 (N_26555,N_24774,N_22609);
or U26556 (N_26556,N_24018,N_22799);
and U26557 (N_26557,N_23455,N_24612);
or U26558 (N_26558,N_23368,N_24688);
nand U26559 (N_26559,N_22902,N_24157);
or U26560 (N_26560,N_24492,N_23106);
and U26561 (N_26561,N_24932,N_23654);
or U26562 (N_26562,N_22613,N_23788);
and U26563 (N_26563,N_22751,N_22815);
nand U26564 (N_26564,N_22615,N_22627);
xor U26565 (N_26565,N_24394,N_23788);
xnor U26566 (N_26566,N_24877,N_22978);
and U26567 (N_26567,N_23278,N_22859);
nand U26568 (N_26568,N_23372,N_24759);
nor U26569 (N_26569,N_22737,N_23518);
and U26570 (N_26570,N_23981,N_22988);
nand U26571 (N_26571,N_23168,N_22613);
or U26572 (N_26572,N_23879,N_22886);
and U26573 (N_26573,N_24053,N_24879);
nand U26574 (N_26574,N_23068,N_22960);
xnor U26575 (N_26575,N_24813,N_23811);
xor U26576 (N_26576,N_23548,N_22886);
nand U26577 (N_26577,N_24681,N_24449);
xor U26578 (N_26578,N_24023,N_23419);
xnor U26579 (N_26579,N_23815,N_22823);
nand U26580 (N_26580,N_23784,N_24798);
xnor U26581 (N_26581,N_24815,N_23490);
nor U26582 (N_26582,N_24210,N_23734);
nor U26583 (N_26583,N_22521,N_24064);
xor U26584 (N_26584,N_23152,N_22989);
nor U26585 (N_26585,N_24062,N_23561);
nand U26586 (N_26586,N_24706,N_23013);
or U26587 (N_26587,N_22809,N_23846);
nand U26588 (N_26588,N_23569,N_22719);
nand U26589 (N_26589,N_23682,N_24683);
and U26590 (N_26590,N_23307,N_22816);
and U26591 (N_26591,N_24691,N_24298);
and U26592 (N_26592,N_22701,N_24751);
nand U26593 (N_26593,N_22889,N_23644);
or U26594 (N_26594,N_24324,N_22597);
nand U26595 (N_26595,N_22835,N_24372);
or U26596 (N_26596,N_23788,N_24336);
nand U26597 (N_26597,N_22763,N_24800);
and U26598 (N_26598,N_22934,N_23254);
nand U26599 (N_26599,N_23103,N_24837);
xor U26600 (N_26600,N_24982,N_23793);
or U26601 (N_26601,N_24955,N_22989);
and U26602 (N_26602,N_24722,N_23498);
or U26603 (N_26603,N_23655,N_22884);
or U26604 (N_26604,N_24004,N_23317);
and U26605 (N_26605,N_22539,N_24420);
xnor U26606 (N_26606,N_24588,N_24868);
nand U26607 (N_26607,N_23060,N_24764);
or U26608 (N_26608,N_23484,N_23122);
or U26609 (N_26609,N_22848,N_22787);
nand U26610 (N_26610,N_24580,N_23426);
xnor U26611 (N_26611,N_24036,N_22840);
and U26612 (N_26612,N_24405,N_23126);
nor U26613 (N_26613,N_23902,N_24585);
xor U26614 (N_26614,N_23728,N_24762);
nor U26615 (N_26615,N_24388,N_24288);
and U26616 (N_26616,N_22649,N_23487);
and U26617 (N_26617,N_23407,N_24919);
nor U26618 (N_26618,N_24622,N_24099);
nand U26619 (N_26619,N_23342,N_23960);
and U26620 (N_26620,N_23814,N_23630);
or U26621 (N_26621,N_24682,N_22800);
or U26622 (N_26622,N_23267,N_23432);
or U26623 (N_26623,N_23339,N_22524);
or U26624 (N_26624,N_23589,N_24426);
nor U26625 (N_26625,N_22612,N_22682);
and U26626 (N_26626,N_23598,N_23983);
xnor U26627 (N_26627,N_23669,N_23451);
nand U26628 (N_26628,N_24437,N_23258);
xnor U26629 (N_26629,N_23634,N_23196);
and U26630 (N_26630,N_23340,N_24502);
and U26631 (N_26631,N_22979,N_24525);
nor U26632 (N_26632,N_24847,N_24985);
or U26633 (N_26633,N_23384,N_24926);
xnor U26634 (N_26634,N_22937,N_22690);
and U26635 (N_26635,N_23641,N_23830);
nor U26636 (N_26636,N_23042,N_24238);
and U26637 (N_26637,N_22613,N_23098);
nand U26638 (N_26638,N_23341,N_22794);
nand U26639 (N_26639,N_24875,N_24618);
or U26640 (N_26640,N_24743,N_23562);
xor U26641 (N_26641,N_24444,N_22561);
and U26642 (N_26642,N_23215,N_23417);
xnor U26643 (N_26643,N_22928,N_24122);
xor U26644 (N_26644,N_24716,N_22722);
xnor U26645 (N_26645,N_22696,N_24030);
xor U26646 (N_26646,N_23081,N_24363);
and U26647 (N_26647,N_23535,N_24888);
nand U26648 (N_26648,N_24445,N_23659);
nor U26649 (N_26649,N_24010,N_23167);
nand U26650 (N_26650,N_23343,N_22865);
and U26651 (N_26651,N_24954,N_24636);
and U26652 (N_26652,N_23230,N_23941);
xnor U26653 (N_26653,N_22728,N_24013);
xnor U26654 (N_26654,N_22669,N_23196);
and U26655 (N_26655,N_24365,N_23726);
nand U26656 (N_26656,N_23138,N_24741);
and U26657 (N_26657,N_23571,N_23568);
nor U26658 (N_26658,N_24129,N_23174);
or U26659 (N_26659,N_24386,N_24967);
nand U26660 (N_26660,N_24270,N_22638);
nand U26661 (N_26661,N_24503,N_24805);
or U26662 (N_26662,N_24401,N_22734);
and U26663 (N_26663,N_23593,N_24833);
nor U26664 (N_26664,N_24374,N_23447);
xnor U26665 (N_26665,N_22540,N_22665);
xnor U26666 (N_26666,N_24958,N_24848);
or U26667 (N_26667,N_24326,N_24389);
nor U26668 (N_26668,N_24422,N_23058);
or U26669 (N_26669,N_22702,N_23880);
nor U26670 (N_26670,N_23075,N_24965);
xnor U26671 (N_26671,N_24887,N_23975);
and U26672 (N_26672,N_23403,N_23909);
or U26673 (N_26673,N_24366,N_23270);
nor U26674 (N_26674,N_24339,N_24120);
nor U26675 (N_26675,N_24581,N_22699);
nor U26676 (N_26676,N_24136,N_23672);
xnor U26677 (N_26677,N_22744,N_22730);
nand U26678 (N_26678,N_22675,N_24643);
nor U26679 (N_26679,N_22954,N_24038);
nand U26680 (N_26680,N_24497,N_23254);
and U26681 (N_26681,N_23467,N_22915);
or U26682 (N_26682,N_24572,N_22541);
or U26683 (N_26683,N_23683,N_23821);
nand U26684 (N_26684,N_23439,N_24389);
and U26685 (N_26685,N_23428,N_22696);
and U26686 (N_26686,N_23279,N_23219);
nor U26687 (N_26687,N_24224,N_24513);
or U26688 (N_26688,N_23971,N_24924);
xnor U26689 (N_26689,N_23333,N_23943);
and U26690 (N_26690,N_23057,N_24106);
xor U26691 (N_26691,N_22916,N_23043);
nor U26692 (N_26692,N_23337,N_24088);
nor U26693 (N_26693,N_24655,N_23666);
nand U26694 (N_26694,N_23348,N_24538);
nand U26695 (N_26695,N_24053,N_24793);
nand U26696 (N_26696,N_24410,N_24238);
nand U26697 (N_26697,N_24053,N_23929);
and U26698 (N_26698,N_24353,N_23752);
or U26699 (N_26699,N_23171,N_22876);
or U26700 (N_26700,N_22779,N_23911);
or U26701 (N_26701,N_24326,N_22636);
nand U26702 (N_26702,N_23206,N_23049);
nor U26703 (N_26703,N_24173,N_24567);
nand U26704 (N_26704,N_24933,N_24879);
xor U26705 (N_26705,N_23809,N_24800);
and U26706 (N_26706,N_24858,N_24026);
or U26707 (N_26707,N_23221,N_23668);
nand U26708 (N_26708,N_23103,N_23459);
nand U26709 (N_26709,N_23390,N_23459);
nor U26710 (N_26710,N_24380,N_24903);
nor U26711 (N_26711,N_24127,N_22871);
and U26712 (N_26712,N_23411,N_22534);
nor U26713 (N_26713,N_23634,N_24826);
nor U26714 (N_26714,N_24821,N_23596);
or U26715 (N_26715,N_23459,N_23669);
nand U26716 (N_26716,N_22814,N_24851);
xor U26717 (N_26717,N_24956,N_24720);
and U26718 (N_26718,N_24759,N_24963);
nand U26719 (N_26719,N_23763,N_24238);
xnor U26720 (N_26720,N_23545,N_24341);
xnor U26721 (N_26721,N_22689,N_23759);
or U26722 (N_26722,N_23065,N_24637);
or U26723 (N_26723,N_24369,N_22729);
xor U26724 (N_26724,N_22623,N_22877);
nand U26725 (N_26725,N_24174,N_23913);
nor U26726 (N_26726,N_24288,N_22821);
nor U26727 (N_26727,N_23205,N_23210);
xor U26728 (N_26728,N_24308,N_24133);
and U26729 (N_26729,N_24930,N_22852);
nand U26730 (N_26730,N_23447,N_24710);
nand U26731 (N_26731,N_23861,N_23190);
or U26732 (N_26732,N_23324,N_24722);
and U26733 (N_26733,N_23221,N_22521);
xor U26734 (N_26734,N_24925,N_24800);
nand U26735 (N_26735,N_23903,N_24278);
nor U26736 (N_26736,N_24948,N_23937);
nand U26737 (N_26737,N_23563,N_24568);
xor U26738 (N_26738,N_22876,N_24386);
nand U26739 (N_26739,N_22657,N_23285);
nor U26740 (N_26740,N_24927,N_24509);
or U26741 (N_26741,N_22597,N_23571);
nand U26742 (N_26742,N_23160,N_23380);
and U26743 (N_26743,N_23564,N_24935);
nor U26744 (N_26744,N_24896,N_23050);
nand U26745 (N_26745,N_23324,N_24704);
nor U26746 (N_26746,N_23491,N_24061);
or U26747 (N_26747,N_23202,N_22677);
nor U26748 (N_26748,N_24463,N_24236);
nand U26749 (N_26749,N_23419,N_23347);
nor U26750 (N_26750,N_24694,N_22551);
and U26751 (N_26751,N_23725,N_23684);
nor U26752 (N_26752,N_23690,N_22502);
nand U26753 (N_26753,N_24418,N_23563);
or U26754 (N_26754,N_24577,N_24019);
nand U26755 (N_26755,N_24788,N_24114);
and U26756 (N_26756,N_23310,N_23779);
nor U26757 (N_26757,N_23758,N_24104);
and U26758 (N_26758,N_24305,N_24573);
or U26759 (N_26759,N_23969,N_23153);
xor U26760 (N_26760,N_23379,N_22906);
xor U26761 (N_26761,N_24706,N_23323);
nor U26762 (N_26762,N_24058,N_22591);
nor U26763 (N_26763,N_23816,N_23456);
nand U26764 (N_26764,N_22510,N_22857);
and U26765 (N_26765,N_23557,N_23440);
xnor U26766 (N_26766,N_23864,N_22795);
nor U26767 (N_26767,N_23980,N_22928);
nand U26768 (N_26768,N_22636,N_24327);
nand U26769 (N_26769,N_24936,N_23233);
nor U26770 (N_26770,N_22644,N_23311);
nor U26771 (N_26771,N_24859,N_23774);
xnor U26772 (N_26772,N_24905,N_22797);
or U26773 (N_26773,N_23061,N_22650);
xor U26774 (N_26774,N_24685,N_23924);
or U26775 (N_26775,N_24005,N_24276);
nor U26776 (N_26776,N_24476,N_22891);
nor U26777 (N_26777,N_23868,N_22795);
nand U26778 (N_26778,N_24790,N_24583);
nand U26779 (N_26779,N_23220,N_24723);
and U26780 (N_26780,N_24716,N_24872);
nor U26781 (N_26781,N_24528,N_24913);
xor U26782 (N_26782,N_23511,N_22981);
and U26783 (N_26783,N_23246,N_24632);
nand U26784 (N_26784,N_22524,N_23154);
nor U26785 (N_26785,N_23245,N_22856);
nor U26786 (N_26786,N_24075,N_23844);
xnor U26787 (N_26787,N_22769,N_24226);
and U26788 (N_26788,N_23794,N_23463);
nand U26789 (N_26789,N_22600,N_24664);
or U26790 (N_26790,N_24578,N_22719);
xnor U26791 (N_26791,N_24538,N_24384);
nor U26792 (N_26792,N_23644,N_24565);
nand U26793 (N_26793,N_23146,N_24541);
or U26794 (N_26794,N_22705,N_22698);
nand U26795 (N_26795,N_23199,N_23443);
nand U26796 (N_26796,N_24757,N_23633);
and U26797 (N_26797,N_23319,N_23647);
xnor U26798 (N_26798,N_23670,N_23974);
nand U26799 (N_26799,N_24623,N_23104);
xor U26800 (N_26800,N_23376,N_22706);
nor U26801 (N_26801,N_22521,N_22993);
xor U26802 (N_26802,N_23127,N_24805);
xnor U26803 (N_26803,N_24143,N_24138);
xnor U26804 (N_26804,N_22905,N_24030);
xor U26805 (N_26805,N_22793,N_24441);
or U26806 (N_26806,N_23736,N_22662);
and U26807 (N_26807,N_22873,N_23020);
or U26808 (N_26808,N_24738,N_22701);
and U26809 (N_26809,N_23594,N_24958);
and U26810 (N_26810,N_23915,N_23806);
and U26811 (N_26811,N_22850,N_22930);
nand U26812 (N_26812,N_24298,N_24105);
xnor U26813 (N_26813,N_23184,N_23076);
or U26814 (N_26814,N_24907,N_23749);
xnor U26815 (N_26815,N_23076,N_23477);
or U26816 (N_26816,N_23861,N_22847);
nor U26817 (N_26817,N_23409,N_23207);
and U26818 (N_26818,N_22676,N_23782);
nor U26819 (N_26819,N_23029,N_22745);
xnor U26820 (N_26820,N_24001,N_23130);
nor U26821 (N_26821,N_24298,N_24931);
or U26822 (N_26822,N_23284,N_24228);
or U26823 (N_26823,N_23194,N_24815);
nand U26824 (N_26824,N_23725,N_24330);
xnor U26825 (N_26825,N_22624,N_22947);
nand U26826 (N_26826,N_24874,N_23905);
or U26827 (N_26827,N_24814,N_24715);
or U26828 (N_26828,N_23493,N_23263);
or U26829 (N_26829,N_23347,N_22688);
nand U26830 (N_26830,N_23472,N_23380);
xnor U26831 (N_26831,N_23264,N_24165);
and U26832 (N_26832,N_22929,N_22936);
nand U26833 (N_26833,N_22886,N_23085);
nand U26834 (N_26834,N_23295,N_24461);
nand U26835 (N_26835,N_22863,N_23623);
and U26836 (N_26836,N_23829,N_22946);
and U26837 (N_26837,N_23428,N_24893);
or U26838 (N_26838,N_22827,N_24039);
or U26839 (N_26839,N_24058,N_23886);
nor U26840 (N_26840,N_24593,N_24829);
xnor U26841 (N_26841,N_23312,N_24729);
or U26842 (N_26842,N_23831,N_22711);
nand U26843 (N_26843,N_23561,N_24075);
or U26844 (N_26844,N_23302,N_22695);
xor U26845 (N_26845,N_22628,N_24622);
xor U26846 (N_26846,N_24933,N_24323);
nor U26847 (N_26847,N_24958,N_23471);
nor U26848 (N_26848,N_23709,N_23386);
nor U26849 (N_26849,N_24632,N_23596);
nor U26850 (N_26850,N_24379,N_22973);
or U26851 (N_26851,N_22698,N_22978);
nor U26852 (N_26852,N_23814,N_23899);
nor U26853 (N_26853,N_24052,N_24064);
nor U26854 (N_26854,N_23779,N_24292);
nand U26855 (N_26855,N_23788,N_24868);
xor U26856 (N_26856,N_24237,N_22703);
and U26857 (N_26857,N_24521,N_24691);
nand U26858 (N_26858,N_23757,N_22532);
or U26859 (N_26859,N_23347,N_22698);
and U26860 (N_26860,N_23366,N_24778);
nor U26861 (N_26861,N_23299,N_24729);
nand U26862 (N_26862,N_23533,N_22506);
and U26863 (N_26863,N_23898,N_24333);
or U26864 (N_26864,N_22512,N_23263);
nand U26865 (N_26865,N_24547,N_24223);
and U26866 (N_26866,N_22819,N_23629);
xnor U26867 (N_26867,N_22515,N_24725);
nor U26868 (N_26868,N_24519,N_23517);
xnor U26869 (N_26869,N_23106,N_24742);
nor U26870 (N_26870,N_23748,N_24283);
nor U26871 (N_26871,N_23489,N_24795);
nand U26872 (N_26872,N_23852,N_22725);
or U26873 (N_26873,N_22866,N_23241);
or U26874 (N_26874,N_23800,N_23310);
nand U26875 (N_26875,N_24731,N_23602);
or U26876 (N_26876,N_24143,N_23287);
xor U26877 (N_26877,N_23144,N_23957);
and U26878 (N_26878,N_23893,N_24249);
and U26879 (N_26879,N_22786,N_23705);
and U26880 (N_26880,N_24466,N_24979);
nand U26881 (N_26881,N_23790,N_24468);
xor U26882 (N_26882,N_23718,N_22601);
nand U26883 (N_26883,N_24823,N_23198);
or U26884 (N_26884,N_23394,N_24371);
or U26885 (N_26885,N_23561,N_24011);
nor U26886 (N_26886,N_24790,N_22762);
nor U26887 (N_26887,N_23302,N_24661);
nor U26888 (N_26888,N_24561,N_23481);
and U26889 (N_26889,N_23585,N_24228);
or U26890 (N_26890,N_24439,N_22848);
and U26891 (N_26891,N_24479,N_23428);
nor U26892 (N_26892,N_22863,N_24081);
and U26893 (N_26893,N_22787,N_24341);
nand U26894 (N_26894,N_23932,N_23447);
nor U26895 (N_26895,N_24906,N_23869);
xnor U26896 (N_26896,N_22519,N_23686);
and U26897 (N_26897,N_24799,N_23296);
and U26898 (N_26898,N_23181,N_22986);
xor U26899 (N_26899,N_22586,N_23734);
and U26900 (N_26900,N_23526,N_23779);
nand U26901 (N_26901,N_22871,N_23122);
nand U26902 (N_26902,N_23143,N_24120);
or U26903 (N_26903,N_24938,N_23786);
and U26904 (N_26904,N_22966,N_23406);
nor U26905 (N_26905,N_22722,N_22955);
nor U26906 (N_26906,N_23743,N_23574);
nor U26907 (N_26907,N_23195,N_22872);
or U26908 (N_26908,N_22511,N_24639);
or U26909 (N_26909,N_23878,N_22936);
and U26910 (N_26910,N_23414,N_24585);
and U26911 (N_26911,N_23776,N_24005);
and U26912 (N_26912,N_22535,N_24287);
nand U26913 (N_26913,N_24538,N_22724);
xnor U26914 (N_26914,N_24527,N_24496);
nor U26915 (N_26915,N_23402,N_24299);
or U26916 (N_26916,N_24845,N_22792);
nand U26917 (N_26917,N_22681,N_23291);
xor U26918 (N_26918,N_24866,N_22690);
nor U26919 (N_26919,N_22973,N_24478);
or U26920 (N_26920,N_24470,N_22872);
nand U26921 (N_26921,N_22900,N_22938);
nand U26922 (N_26922,N_23554,N_24500);
and U26923 (N_26923,N_23642,N_23619);
xnor U26924 (N_26924,N_24753,N_24622);
nand U26925 (N_26925,N_22722,N_24319);
nand U26926 (N_26926,N_22986,N_23872);
or U26927 (N_26927,N_24955,N_23334);
nand U26928 (N_26928,N_23877,N_24591);
nand U26929 (N_26929,N_23861,N_23144);
nand U26930 (N_26930,N_22522,N_23872);
and U26931 (N_26931,N_22930,N_23735);
nor U26932 (N_26932,N_22582,N_23994);
xnor U26933 (N_26933,N_23294,N_23209);
or U26934 (N_26934,N_24621,N_24294);
xor U26935 (N_26935,N_24768,N_24316);
nand U26936 (N_26936,N_24138,N_23341);
and U26937 (N_26937,N_24159,N_23880);
nand U26938 (N_26938,N_23206,N_23863);
xor U26939 (N_26939,N_23015,N_23497);
xor U26940 (N_26940,N_22888,N_24316);
or U26941 (N_26941,N_22536,N_24774);
nand U26942 (N_26942,N_24268,N_24656);
or U26943 (N_26943,N_24758,N_24793);
nor U26944 (N_26944,N_23349,N_23986);
xor U26945 (N_26945,N_22824,N_24854);
nand U26946 (N_26946,N_24331,N_23014);
xor U26947 (N_26947,N_24232,N_24907);
xnor U26948 (N_26948,N_23324,N_23511);
or U26949 (N_26949,N_24081,N_23274);
or U26950 (N_26950,N_23036,N_23514);
nand U26951 (N_26951,N_24952,N_24908);
nand U26952 (N_26952,N_24317,N_24199);
nor U26953 (N_26953,N_22848,N_23217);
and U26954 (N_26954,N_23552,N_23647);
or U26955 (N_26955,N_23680,N_23691);
and U26956 (N_26956,N_23957,N_24661);
or U26957 (N_26957,N_22734,N_22648);
xor U26958 (N_26958,N_23985,N_22958);
or U26959 (N_26959,N_24915,N_23132);
or U26960 (N_26960,N_23571,N_24919);
and U26961 (N_26961,N_22910,N_23491);
nand U26962 (N_26962,N_23804,N_23861);
nor U26963 (N_26963,N_24827,N_23412);
nand U26964 (N_26964,N_24960,N_24217);
nand U26965 (N_26965,N_24445,N_23639);
and U26966 (N_26966,N_24677,N_23151);
and U26967 (N_26967,N_23182,N_24959);
or U26968 (N_26968,N_22681,N_22979);
or U26969 (N_26969,N_24425,N_24823);
xor U26970 (N_26970,N_24553,N_22923);
nand U26971 (N_26971,N_24935,N_24749);
xnor U26972 (N_26972,N_24402,N_24288);
nor U26973 (N_26973,N_23654,N_23034);
and U26974 (N_26974,N_24095,N_24487);
and U26975 (N_26975,N_24985,N_23159);
nor U26976 (N_26976,N_24440,N_22662);
or U26977 (N_26977,N_23290,N_23046);
nor U26978 (N_26978,N_24587,N_23905);
nand U26979 (N_26979,N_24071,N_24749);
or U26980 (N_26980,N_22677,N_24780);
and U26981 (N_26981,N_23537,N_23402);
or U26982 (N_26982,N_23342,N_24354);
nand U26983 (N_26983,N_24979,N_22841);
nor U26984 (N_26984,N_23690,N_24399);
and U26985 (N_26985,N_23885,N_24306);
nand U26986 (N_26986,N_24237,N_22985);
and U26987 (N_26987,N_22631,N_22574);
nand U26988 (N_26988,N_22619,N_23102);
nand U26989 (N_26989,N_22946,N_24101);
and U26990 (N_26990,N_24626,N_23694);
or U26991 (N_26991,N_23837,N_23485);
and U26992 (N_26992,N_23535,N_22778);
and U26993 (N_26993,N_23969,N_23965);
xor U26994 (N_26994,N_23701,N_24071);
nor U26995 (N_26995,N_24718,N_24315);
nand U26996 (N_26996,N_23565,N_24291);
nand U26997 (N_26997,N_24506,N_22851);
or U26998 (N_26998,N_24654,N_22729);
nand U26999 (N_26999,N_24093,N_24641);
nor U27000 (N_27000,N_23257,N_23857);
xnor U27001 (N_27001,N_22776,N_24724);
nand U27002 (N_27002,N_23594,N_22543);
xor U27003 (N_27003,N_23559,N_24872);
nor U27004 (N_27004,N_22742,N_24582);
xnor U27005 (N_27005,N_22686,N_22567);
or U27006 (N_27006,N_23928,N_22691);
nand U27007 (N_27007,N_23315,N_22660);
xnor U27008 (N_27008,N_24264,N_23870);
nand U27009 (N_27009,N_23202,N_24847);
xor U27010 (N_27010,N_24402,N_24708);
xor U27011 (N_27011,N_22948,N_24823);
and U27012 (N_27012,N_23326,N_23738);
xnor U27013 (N_27013,N_22734,N_23255);
nor U27014 (N_27014,N_24169,N_24205);
nand U27015 (N_27015,N_23117,N_22914);
xor U27016 (N_27016,N_22759,N_24227);
nand U27017 (N_27017,N_24348,N_23350);
xnor U27018 (N_27018,N_24702,N_24163);
xor U27019 (N_27019,N_22742,N_23848);
nand U27020 (N_27020,N_22798,N_24905);
nor U27021 (N_27021,N_23705,N_24806);
xor U27022 (N_27022,N_24700,N_24113);
nand U27023 (N_27023,N_24161,N_23298);
nor U27024 (N_27024,N_24797,N_24848);
or U27025 (N_27025,N_24739,N_22695);
nor U27026 (N_27026,N_22578,N_24133);
nand U27027 (N_27027,N_22522,N_24218);
xor U27028 (N_27028,N_23027,N_22967);
nor U27029 (N_27029,N_23928,N_24262);
or U27030 (N_27030,N_24658,N_24067);
and U27031 (N_27031,N_23718,N_23891);
and U27032 (N_27032,N_24648,N_23311);
xor U27033 (N_27033,N_24090,N_24698);
or U27034 (N_27034,N_24366,N_23914);
nand U27035 (N_27035,N_23573,N_23264);
xor U27036 (N_27036,N_23274,N_23027);
and U27037 (N_27037,N_23268,N_23748);
or U27038 (N_27038,N_24510,N_24461);
nand U27039 (N_27039,N_23687,N_23801);
or U27040 (N_27040,N_23014,N_23947);
nand U27041 (N_27041,N_22851,N_23055);
nor U27042 (N_27042,N_23275,N_24817);
and U27043 (N_27043,N_24988,N_24545);
or U27044 (N_27044,N_24760,N_23585);
xor U27045 (N_27045,N_24362,N_23228);
and U27046 (N_27046,N_24886,N_24298);
or U27047 (N_27047,N_24330,N_24827);
nand U27048 (N_27048,N_23543,N_24613);
nand U27049 (N_27049,N_24336,N_22752);
and U27050 (N_27050,N_24773,N_23450);
xnor U27051 (N_27051,N_24532,N_24373);
xor U27052 (N_27052,N_23763,N_24869);
xor U27053 (N_27053,N_23222,N_24072);
nand U27054 (N_27054,N_23767,N_24938);
and U27055 (N_27055,N_24212,N_23586);
nor U27056 (N_27056,N_23296,N_22831);
and U27057 (N_27057,N_24090,N_24494);
nand U27058 (N_27058,N_23580,N_22659);
nor U27059 (N_27059,N_24717,N_22655);
nor U27060 (N_27060,N_24487,N_23761);
xor U27061 (N_27061,N_24136,N_22931);
nand U27062 (N_27062,N_24051,N_22962);
nand U27063 (N_27063,N_22581,N_23029);
and U27064 (N_27064,N_23423,N_24633);
or U27065 (N_27065,N_23556,N_23185);
nand U27066 (N_27066,N_24081,N_23442);
or U27067 (N_27067,N_24796,N_24166);
xor U27068 (N_27068,N_23746,N_24796);
xnor U27069 (N_27069,N_24274,N_22513);
or U27070 (N_27070,N_23244,N_23153);
xnor U27071 (N_27071,N_23140,N_24099);
nand U27072 (N_27072,N_24071,N_23690);
or U27073 (N_27073,N_23640,N_23007);
nand U27074 (N_27074,N_24519,N_23388);
or U27075 (N_27075,N_23816,N_22964);
nand U27076 (N_27076,N_24573,N_23119);
and U27077 (N_27077,N_24833,N_23817);
and U27078 (N_27078,N_22608,N_23635);
nand U27079 (N_27079,N_23991,N_23206);
and U27080 (N_27080,N_24432,N_24134);
and U27081 (N_27081,N_23802,N_24331);
nor U27082 (N_27082,N_24314,N_23227);
and U27083 (N_27083,N_22677,N_22980);
nor U27084 (N_27084,N_24838,N_23355);
and U27085 (N_27085,N_23851,N_24476);
nand U27086 (N_27086,N_24948,N_23158);
xnor U27087 (N_27087,N_22625,N_23743);
nand U27088 (N_27088,N_22794,N_24840);
and U27089 (N_27089,N_24974,N_23868);
xor U27090 (N_27090,N_23259,N_22627);
nand U27091 (N_27091,N_24301,N_23846);
nor U27092 (N_27092,N_24815,N_22949);
and U27093 (N_27093,N_22604,N_24882);
xnor U27094 (N_27094,N_23446,N_24776);
or U27095 (N_27095,N_22541,N_24523);
nor U27096 (N_27096,N_24730,N_22765);
and U27097 (N_27097,N_22537,N_24513);
xnor U27098 (N_27098,N_22827,N_22806);
nand U27099 (N_27099,N_23816,N_22829);
nor U27100 (N_27100,N_24760,N_23936);
xor U27101 (N_27101,N_23671,N_24995);
or U27102 (N_27102,N_23126,N_22934);
nand U27103 (N_27103,N_23044,N_24531);
xor U27104 (N_27104,N_23869,N_23263);
nor U27105 (N_27105,N_22713,N_23818);
or U27106 (N_27106,N_24485,N_24926);
and U27107 (N_27107,N_24462,N_22720);
or U27108 (N_27108,N_23733,N_24915);
or U27109 (N_27109,N_22572,N_23545);
nor U27110 (N_27110,N_22532,N_23348);
xor U27111 (N_27111,N_23943,N_23852);
xnor U27112 (N_27112,N_24904,N_23847);
and U27113 (N_27113,N_24349,N_23044);
and U27114 (N_27114,N_23839,N_24658);
xor U27115 (N_27115,N_24300,N_24445);
nor U27116 (N_27116,N_23873,N_24432);
and U27117 (N_27117,N_24452,N_23861);
or U27118 (N_27118,N_24563,N_23234);
and U27119 (N_27119,N_23530,N_22587);
or U27120 (N_27120,N_23903,N_24296);
or U27121 (N_27121,N_24451,N_24385);
xnor U27122 (N_27122,N_23886,N_24315);
and U27123 (N_27123,N_24231,N_23589);
and U27124 (N_27124,N_24393,N_24067);
xnor U27125 (N_27125,N_22672,N_24872);
xnor U27126 (N_27126,N_24216,N_24605);
and U27127 (N_27127,N_23562,N_24411);
and U27128 (N_27128,N_24658,N_23231);
xor U27129 (N_27129,N_24868,N_23596);
or U27130 (N_27130,N_22563,N_23780);
nor U27131 (N_27131,N_24703,N_24046);
and U27132 (N_27132,N_24093,N_24961);
xor U27133 (N_27133,N_24753,N_24108);
nor U27134 (N_27134,N_24541,N_23933);
nand U27135 (N_27135,N_24120,N_22957);
nand U27136 (N_27136,N_23648,N_23121);
and U27137 (N_27137,N_24669,N_23790);
nand U27138 (N_27138,N_24375,N_22683);
nand U27139 (N_27139,N_22630,N_24174);
nor U27140 (N_27140,N_23515,N_23102);
or U27141 (N_27141,N_23392,N_24290);
xnor U27142 (N_27142,N_22556,N_23837);
and U27143 (N_27143,N_24311,N_23766);
nor U27144 (N_27144,N_24125,N_24424);
nand U27145 (N_27145,N_23025,N_22882);
and U27146 (N_27146,N_23834,N_24622);
nor U27147 (N_27147,N_24803,N_23026);
nor U27148 (N_27148,N_24543,N_23289);
nor U27149 (N_27149,N_23924,N_24129);
xor U27150 (N_27150,N_23913,N_24769);
and U27151 (N_27151,N_24003,N_24799);
or U27152 (N_27152,N_24949,N_23696);
xnor U27153 (N_27153,N_23815,N_24391);
nor U27154 (N_27154,N_23857,N_24620);
or U27155 (N_27155,N_23199,N_23953);
or U27156 (N_27156,N_24225,N_23449);
or U27157 (N_27157,N_23504,N_24856);
nor U27158 (N_27158,N_22908,N_23640);
nor U27159 (N_27159,N_24273,N_23909);
nand U27160 (N_27160,N_24931,N_24337);
nor U27161 (N_27161,N_24844,N_23293);
nor U27162 (N_27162,N_23149,N_22947);
or U27163 (N_27163,N_23563,N_22557);
nor U27164 (N_27164,N_24069,N_23303);
and U27165 (N_27165,N_23958,N_24625);
nor U27166 (N_27166,N_24099,N_23544);
xor U27167 (N_27167,N_24433,N_23869);
xnor U27168 (N_27168,N_23444,N_22614);
nand U27169 (N_27169,N_23464,N_24587);
nand U27170 (N_27170,N_24750,N_22842);
nor U27171 (N_27171,N_22883,N_23745);
nand U27172 (N_27172,N_23478,N_24510);
and U27173 (N_27173,N_23780,N_23969);
or U27174 (N_27174,N_24871,N_24713);
nand U27175 (N_27175,N_23954,N_24170);
nand U27176 (N_27176,N_23183,N_22711);
nor U27177 (N_27177,N_24042,N_23457);
nand U27178 (N_27178,N_24875,N_24303);
nor U27179 (N_27179,N_22532,N_23810);
and U27180 (N_27180,N_22511,N_24180);
nand U27181 (N_27181,N_22549,N_23112);
nand U27182 (N_27182,N_24732,N_23048);
or U27183 (N_27183,N_24707,N_24180);
nor U27184 (N_27184,N_23131,N_22855);
or U27185 (N_27185,N_22867,N_24737);
or U27186 (N_27186,N_22656,N_24671);
xor U27187 (N_27187,N_23481,N_23932);
and U27188 (N_27188,N_24749,N_22646);
nor U27189 (N_27189,N_24714,N_23529);
nand U27190 (N_27190,N_23353,N_24501);
or U27191 (N_27191,N_22816,N_23984);
or U27192 (N_27192,N_23416,N_22779);
nor U27193 (N_27193,N_23482,N_24770);
and U27194 (N_27194,N_24232,N_24902);
xor U27195 (N_27195,N_23296,N_24044);
nor U27196 (N_27196,N_23627,N_23132);
xnor U27197 (N_27197,N_23899,N_23102);
or U27198 (N_27198,N_23633,N_23961);
nand U27199 (N_27199,N_23997,N_23955);
xor U27200 (N_27200,N_24393,N_24257);
xor U27201 (N_27201,N_24899,N_23806);
nor U27202 (N_27202,N_24590,N_23377);
and U27203 (N_27203,N_23603,N_23135);
and U27204 (N_27204,N_24568,N_24212);
nand U27205 (N_27205,N_23032,N_24452);
nor U27206 (N_27206,N_24505,N_23204);
nand U27207 (N_27207,N_24376,N_24002);
and U27208 (N_27208,N_24666,N_23873);
nand U27209 (N_27209,N_23079,N_24430);
xor U27210 (N_27210,N_24820,N_23239);
nand U27211 (N_27211,N_22849,N_24795);
xor U27212 (N_27212,N_24503,N_22623);
xnor U27213 (N_27213,N_24444,N_23672);
xor U27214 (N_27214,N_24262,N_24276);
nor U27215 (N_27215,N_24925,N_24966);
or U27216 (N_27216,N_24504,N_23090);
nand U27217 (N_27217,N_23467,N_23166);
nor U27218 (N_27218,N_24566,N_23955);
xnor U27219 (N_27219,N_24074,N_24686);
or U27220 (N_27220,N_24654,N_24852);
and U27221 (N_27221,N_24177,N_23998);
and U27222 (N_27222,N_24796,N_22847);
and U27223 (N_27223,N_22815,N_23896);
nand U27224 (N_27224,N_22711,N_24831);
or U27225 (N_27225,N_24841,N_24468);
xnor U27226 (N_27226,N_23017,N_24055);
or U27227 (N_27227,N_22811,N_23179);
and U27228 (N_27228,N_24182,N_24801);
or U27229 (N_27229,N_23787,N_23728);
xnor U27230 (N_27230,N_22998,N_22835);
xor U27231 (N_27231,N_24888,N_24027);
xor U27232 (N_27232,N_24208,N_23070);
xnor U27233 (N_27233,N_24023,N_22629);
or U27234 (N_27234,N_22660,N_23286);
or U27235 (N_27235,N_23804,N_23694);
nor U27236 (N_27236,N_23296,N_22840);
or U27237 (N_27237,N_24797,N_24396);
and U27238 (N_27238,N_23286,N_24900);
and U27239 (N_27239,N_23519,N_23008);
nand U27240 (N_27240,N_22884,N_24393);
nor U27241 (N_27241,N_23280,N_22923);
xor U27242 (N_27242,N_24507,N_23602);
or U27243 (N_27243,N_24575,N_23253);
nor U27244 (N_27244,N_23549,N_23163);
nor U27245 (N_27245,N_24483,N_22561);
nor U27246 (N_27246,N_24968,N_24114);
xnor U27247 (N_27247,N_23660,N_24156);
nor U27248 (N_27248,N_24006,N_24946);
and U27249 (N_27249,N_23239,N_24495);
nand U27250 (N_27250,N_24350,N_22839);
or U27251 (N_27251,N_24363,N_24446);
and U27252 (N_27252,N_23300,N_23967);
nor U27253 (N_27253,N_24220,N_22815);
or U27254 (N_27254,N_22945,N_24769);
xor U27255 (N_27255,N_23302,N_24431);
nor U27256 (N_27256,N_22780,N_22540);
or U27257 (N_27257,N_23260,N_24672);
and U27258 (N_27258,N_22883,N_24912);
or U27259 (N_27259,N_24287,N_23241);
nand U27260 (N_27260,N_24471,N_22791);
or U27261 (N_27261,N_24128,N_24951);
or U27262 (N_27262,N_23944,N_22991);
xor U27263 (N_27263,N_22921,N_22837);
nor U27264 (N_27264,N_23825,N_22622);
and U27265 (N_27265,N_24205,N_23023);
nor U27266 (N_27266,N_24136,N_23416);
and U27267 (N_27267,N_24415,N_24417);
and U27268 (N_27268,N_24307,N_23513);
nor U27269 (N_27269,N_24186,N_22926);
and U27270 (N_27270,N_24153,N_24431);
and U27271 (N_27271,N_23178,N_23843);
xor U27272 (N_27272,N_24864,N_22998);
xor U27273 (N_27273,N_23600,N_24330);
and U27274 (N_27274,N_23527,N_23479);
nand U27275 (N_27275,N_22866,N_24701);
nand U27276 (N_27276,N_24330,N_23068);
nor U27277 (N_27277,N_22954,N_23913);
or U27278 (N_27278,N_23098,N_22677);
xnor U27279 (N_27279,N_22990,N_24179);
nor U27280 (N_27280,N_24733,N_23022);
and U27281 (N_27281,N_24273,N_24105);
nor U27282 (N_27282,N_23471,N_22890);
and U27283 (N_27283,N_22687,N_22719);
and U27284 (N_27284,N_24273,N_23354);
and U27285 (N_27285,N_22981,N_23977);
or U27286 (N_27286,N_23929,N_24615);
nand U27287 (N_27287,N_24267,N_23340);
nand U27288 (N_27288,N_23561,N_23843);
nor U27289 (N_27289,N_24465,N_24381);
or U27290 (N_27290,N_24278,N_22525);
nand U27291 (N_27291,N_23705,N_23200);
nand U27292 (N_27292,N_23089,N_22924);
nor U27293 (N_27293,N_24751,N_23586);
nor U27294 (N_27294,N_24295,N_24936);
and U27295 (N_27295,N_23450,N_24692);
nor U27296 (N_27296,N_24881,N_22820);
nor U27297 (N_27297,N_24794,N_24379);
or U27298 (N_27298,N_23005,N_22560);
nand U27299 (N_27299,N_22550,N_23060);
xor U27300 (N_27300,N_24009,N_23605);
or U27301 (N_27301,N_22889,N_24875);
and U27302 (N_27302,N_24136,N_22940);
or U27303 (N_27303,N_22775,N_24614);
nor U27304 (N_27304,N_24404,N_24325);
or U27305 (N_27305,N_24632,N_23855);
and U27306 (N_27306,N_24910,N_24194);
and U27307 (N_27307,N_24274,N_23534);
nor U27308 (N_27308,N_24749,N_24435);
xnor U27309 (N_27309,N_24828,N_24839);
and U27310 (N_27310,N_24001,N_22928);
nand U27311 (N_27311,N_23250,N_22934);
and U27312 (N_27312,N_23064,N_22967);
nand U27313 (N_27313,N_23702,N_22767);
nor U27314 (N_27314,N_23857,N_22833);
nand U27315 (N_27315,N_23571,N_23041);
or U27316 (N_27316,N_24133,N_23324);
or U27317 (N_27317,N_22890,N_23772);
or U27318 (N_27318,N_22718,N_24627);
xnor U27319 (N_27319,N_23249,N_22723);
and U27320 (N_27320,N_23985,N_24651);
xnor U27321 (N_27321,N_22739,N_24102);
or U27322 (N_27322,N_24935,N_23592);
or U27323 (N_27323,N_23338,N_23116);
xnor U27324 (N_27324,N_24684,N_24269);
nand U27325 (N_27325,N_24640,N_24888);
or U27326 (N_27326,N_24738,N_24885);
or U27327 (N_27327,N_23376,N_23360);
and U27328 (N_27328,N_22989,N_22610);
nand U27329 (N_27329,N_23825,N_23869);
nor U27330 (N_27330,N_22970,N_24802);
nor U27331 (N_27331,N_24798,N_23630);
xnor U27332 (N_27332,N_24372,N_22567);
xor U27333 (N_27333,N_23119,N_23898);
nor U27334 (N_27334,N_23297,N_24376);
nor U27335 (N_27335,N_23460,N_24357);
xor U27336 (N_27336,N_24995,N_23602);
xnor U27337 (N_27337,N_24701,N_22539);
xor U27338 (N_27338,N_24373,N_23066);
and U27339 (N_27339,N_22501,N_24802);
or U27340 (N_27340,N_23937,N_24705);
xnor U27341 (N_27341,N_24438,N_24832);
or U27342 (N_27342,N_23406,N_23350);
or U27343 (N_27343,N_24822,N_23261);
xnor U27344 (N_27344,N_24055,N_23423);
xor U27345 (N_27345,N_22969,N_22593);
nand U27346 (N_27346,N_23988,N_22990);
or U27347 (N_27347,N_24006,N_24453);
xnor U27348 (N_27348,N_23693,N_23468);
or U27349 (N_27349,N_24005,N_22928);
nand U27350 (N_27350,N_24146,N_22781);
nor U27351 (N_27351,N_22667,N_23514);
xnor U27352 (N_27352,N_24842,N_23890);
or U27353 (N_27353,N_22753,N_24741);
nor U27354 (N_27354,N_23601,N_24999);
and U27355 (N_27355,N_23583,N_23268);
nand U27356 (N_27356,N_23248,N_23636);
or U27357 (N_27357,N_24580,N_24528);
and U27358 (N_27358,N_23555,N_23678);
and U27359 (N_27359,N_24424,N_24650);
nand U27360 (N_27360,N_24397,N_24130);
nand U27361 (N_27361,N_24431,N_22507);
nand U27362 (N_27362,N_22619,N_24468);
nand U27363 (N_27363,N_24338,N_24199);
nand U27364 (N_27364,N_22629,N_24598);
nand U27365 (N_27365,N_23417,N_24999);
or U27366 (N_27366,N_23230,N_24294);
and U27367 (N_27367,N_22779,N_23983);
or U27368 (N_27368,N_24927,N_24527);
nor U27369 (N_27369,N_24570,N_24555);
nand U27370 (N_27370,N_22874,N_23869);
or U27371 (N_27371,N_23997,N_24367);
xor U27372 (N_27372,N_24547,N_23811);
nand U27373 (N_27373,N_24829,N_22527);
or U27374 (N_27374,N_24248,N_24578);
xnor U27375 (N_27375,N_23894,N_23787);
xnor U27376 (N_27376,N_22706,N_24726);
and U27377 (N_27377,N_22895,N_24940);
xor U27378 (N_27378,N_23396,N_23271);
or U27379 (N_27379,N_24060,N_24237);
nand U27380 (N_27380,N_23086,N_24897);
nor U27381 (N_27381,N_24194,N_22949);
and U27382 (N_27382,N_22514,N_22644);
xor U27383 (N_27383,N_24509,N_24905);
xor U27384 (N_27384,N_24261,N_22511);
and U27385 (N_27385,N_23592,N_24821);
nand U27386 (N_27386,N_23235,N_22564);
xnor U27387 (N_27387,N_23010,N_24397);
nor U27388 (N_27388,N_24000,N_22900);
or U27389 (N_27389,N_23270,N_24770);
xor U27390 (N_27390,N_23637,N_24856);
xnor U27391 (N_27391,N_23788,N_24089);
or U27392 (N_27392,N_24299,N_23541);
or U27393 (N_27393,N_24270,N_24726);
and U27394 (N_27394,N_23672,N_23233);
or U27395 (N_27395,N_24363,N_23417);
nand U27396 (N_27396,N_24756,N_23160);
nor U27397 (N_27397,N_23765,N_24869);
nor U27398 (N_27398,N_23926,N_24905);
nand U27399 (N_27399,N_23231,N_23654);
nor U27400 (N_27400,N_23953,N_24531);
and U27401 (N_27401,N_24152,N_24001);
or U27402 (N_27402,N_23458,N_23429);
and U27403 (N_27403,N_23566,N_24469);
xnor U27404 (N_27404,N_23753,N_24038);
nand U27405 (N_27405,N_23451,N_24005);
and U27406 (N_27406,N_22543,N_23378);
nor U27407 (N_27407,N_22772,N_24594);
and U27408 (N_27408,N_23770,N_24889);
xnor U27409 (N_27409,N_24906,N_22795);
and U27410 (N_27410,N_23004,N_23892);
and U27411 (N_27411,N_22842,N_24181);
and U27412 (N_27412,N_24855,N_23238);
or U27413 (N_27413,N_24963,N_22629);
nand U27414 (N_27414,N_24865,N_24875);
nand U27415 (N_27415,N_23811,N_22852);
xor U27416 (N_27416,N_23055,N_23004);
xnor U27417 (N_27417,N_24059,N_24089);
nand U27418 (N_27418,N_23626,N_24785);
nor U27419 (N_27419,N_24980,N_24683);
xor U27420 (N_27420,N_22542,N_23029);
nor U27421 (N_27421,N_24008,N_24387);
nand U27422 (N_27422,N_22911,N_24748);
nand U27423 (N_27423,N_24621,N_23672);
or U27424 (N_27424,N_23513,N_22756);
or U27425 (N_27425,N_23991,N_24747);
xor U27426 (N_27426,N_23136,N_24719);
xor U27427 (N_27427,N_24044,N_22637);
nand U27428 (N_27428,N_22870,N_23266);
xor U27429 (N_27429,N_24111,N_23997);
or U27430 (N_27430,N_22596,N_23485);
or U27431 (N_27431,N_23593,N_22796);
nor U27432 (N_27432,N_22848,N_24151);
xor U27433 (N_27433,N_23847,N_23153);
or U27434 (N_27434,N_23175,N_24783);
nand U27435 (N_27435,N_24274,N_23302);
or U27436 (N_27436,N_22688,N_23554);
and U27437 (N_27437,N_23517,N_24484);
nand U27438 (N_27438,N_23676,N_23777);
nor U27439 (N_27439,N_23359,N_22961);
nor U27440 (N_27440,N_23229,N_23969);
nand U27441 (N_27441,N_22658,N_24787);
and U27442 (N_27442,N_24536,N_23902);
nor U27443 (N_27443,N_24326,N_24010);
nand U27444 (N_27444,N_23346,N_24056);
and U27445 (N_27445,N_24098,N_22508);
or U27446 (N_27446,N_22843,N_23896);
or U27447 (N_27447,N_22761,N_22859);
nand U27448 (N_27448,N_24331,N_24748);
xor U27449 (N_27449,N_22647,N_22524);
nand U27450 (N_27450,N_23358,N_23252);
xnor U27451 (N_27451,N_24981,N_23967);
xor U27452 (N_27452,N_23231,N_24966);
xnor U27453 (N_27453,N_22758,N_24512);
nor U27454 (N_27454,N_23873,N_24642);
nor U27455 (N_27455,N_24974,N_24089);
nor U27456 (N_27456,N_22812,N_23009);
nand U27457 (N_27457,N_23494,N_24725);
nand U27458 (N_27458,N_24019,N_23963);
or U27459 (N_27459,N_24624,N_22687);
nand U27460 (N_27460,N_24645,N_22653);
and U27461 (N_27461,N_22790,N_23836);
nor U27462 (N_27462,N_22887,N_23466);
and U27463 (N_27463,N_24423,N_23808);
and U27464 (N_27464,N_23607,N_23806);
nand U27465 (N_27465,N_23361,N_23584);
and U27466 (N_27466,N_22559,N_24350);
nor U27467 (N_27467,N_24087,N_22850);
and U27468 (N_27468,N_24245,N_23408);
nor U27469 (N_27469,N_23711,N_23681);
xnor U27470 (N_27470,N_24215,N_24393);
and U27471 (N_27471,N_23311,N_24826);
nand U27472 (N_27472,N_23388,N_23812);
or U27473 (N_27473,N_23920,N_24867);
nand U27474 (N_27474,N_23931,N_23202);
or U27475 (N_27475,N_23743,N_24478);
xnor U27476 (N_27476,N_23371,N_24687);
nor U27477 (N_27477,N_24360,N_24656);
or U27478 (N_27478,N_23282,N_22861);
or U27479 (N_27479,N_22928,N_24922);
xnor U27480 (N_27480,N_24762,N_24687);
nand U27481 (N_27481,N_24650,N_23954);
and U27482 (N_27482,N_24002,N_23079);
or U27483 (N_27483,N_23765,N_22556);
nand U27484 (N_27484,N_24585,N_23827);
xor U27485 (N_27485,N_23792,N_22932);
and U27486 (N_27486,N_22655,N_24464);
nor U27487 (N_27487,N_24327,N_23806);
xor U27488 (N_27488,N_24575,N_23124);
nand U27489 (N_27489,N_24200,N_24837);
xor U27490 (N_27490,N_23720,N_23773);
nor U27491 (N_27491,N_22958,N_23282);
nand U27492 (N_27492,N_24859,N_22650);
nand U27493 (N_27493,N_23797,N_23309);
and U27494 (N_27494,N_23952,N_23991);
xor U27495 (N_27495,N_24537,N_22991);
or U27496 (N_27496,N_22552,N_23387);
nor U27497 (N_27497,N_22741,N_24840);
nor U27498 (N_27498,N_22919,N_23339);
and U27499 (N_27499,N_23817,N_23130);
xor U27500 (N_27500,N_25316,N_25909);
nor U27501 (N_27501,N_27385,N_25177);
nand U27502 (N_27502,N_25254,N_27457);
or U27503 (N_27503,N_27083,N_25566);
or U27504 (N_27504,N_26986,N_27002);
and U27505 (N_27505,N_25619,N_25621);
xnor U27506 (N_27506,N_25752,N_26699);
xnor U27507 (N_27507,N_26329,N_26852);
or U27508 (N_27508,N_25387,N_26269);
nand U27509 (N_27509,N_27360,N_26761);
nor U27510 (N_27510,N_27373,N_25609);
xor U27511 (N_27511,N_25979,N_25668);
xor U27512 (N_27512,N_27172,N_26088);
nor U27513 (N_27513,N_25069,N_27053);
xor U27514 (N_27514,N_25150,N_25038);
xor U27515 (N_27515,N_27036,N_27283);
or U27516 (N_27516,N_26407,N_25685);
and U27517 (N_27517,N_25964,N_26502);
nor U27518 (N_27518,N_25191,N_25902);
or U27519 (N_27519,N_25246,N_26194);
and U27520 (N_27520,N_27104,N_27334);
xor U27521 (N_27521,N_26948,N_26819);
nand U27522 (N_27522,N_26432,N_25414);
nand U27523 (N_27523,N_25644,N_27446);
or U27524 (N_27524,N_25986,N_25989);
nand U27525 (N_27525,N_25791,N_25946);
xor U27526 (N_27526,N_26289,N_25125);
xor U27527 (N_27527,N_26863,N_25420);
or U27528 (N_27528,N_25981,N_26633);
nand U27529 (N_27529,N_26987,N_25289);
nand U27530 (N_27530,N_26008,N_25808);
or U27531 (N_27531,N_26672,N_27115);
xor U27532 (N_27532,N_26443,N_25443);
xnor U27533 (N_27533,N_26702,N_27153);
nor U27534 (N_27534,N_27157,N_27009);
xnor U27535 (N_27535,N_25825,N_25733);
nor U27536 (N_27536,N_26964,N_25449);
or U27537 (N_27537,N_25140,N_27482);
nor U27538 (N_27538,N_27177,N_26656);
xor U27539 (N_27539,N_25336,N_27465);
nor U27540 (N_27540,N_25804,N_25624);
or U27541 (N_27541,N_26306,N_27393);
xor U27542 (N_27542,N_26249,N_25592);
or U27543 (N_27543,N_25014,N_25035);
or U27544 (N_27544,N_25811,N_25867);
nand U27545 (N_27545,N_25994,N_25085);
or U27546 (N_27546,N_25232,N_25798);
and U27547 (N_27547,N_26158,N_26052);
xor U27548 (N_27548,N_26757,N_25090);
nand U27549 (N_27549,N_26366,N_26775);
xnor U27550 (N_27550,N_25724,N_25192);
and U27551 (N_27551,N_25375,N_26530);
nor U27552 (N_27552,N_26114,N_26477);
nor U27553 (N_27553,N_25091,N_26940);
and U27554 (N_27554,N_26063,N_26189);
nor U27555 (N_27555,N_26983,N_26186);
nand U27556 (N_27556,N_25359,N_26591);
or U27557 (N_27557,N_25755,N_26414);
nor U27558 (N_27558,N_25153,N_25215);
and U27559 (N_27559,N_25862,N_27026);
nor U27560 (N_27560,N_26913,N_26452);
nand U27561 (N_27561,N_26939,N_25655);
xor U27562 (N_27562,N_26625,N_26092);
nand U27563 (N_27563,N_27391,N_27378);
xor U27564 (N_27564,N_25747,N_25834);
xnor U27565 (N_27565,N_25250,N_26685);
xor U27566 (N_27566,N_25425,N_26365);
and U27567 (N_27567,N_27021,N_27377);
nor U27568 (N_27568,N_26406,N_27357);
nand U27569 (N_27569,N_25880,N_27249);
nand U27570 (N_27570,N_25923,N_25123);
and U27571 (N_27571,N_25794,N_25661);
and U27572 (N_27572,N_25866,N_25918);
or U27573 (N_27573,N_27062,N_25228);
xnor U27574 (N_27574,N_26715,N_27178);
nand U27575 (N_27575,N_27440,N_25380);
or U27576 (N_27576,N_26420,N_26442);
nor U27577 (N_27577,N_26455,N_26816);
and U27578 (N_27578,N_26547,N_27302);
nand U27579 (N_27579,N_25006,N_26730);
nand U27580 (N_27580,N_25002,N_27164);
or U27581 (N_27581,N_26815,N_27354);
or U27582 (N_27582,N_26473,N_26509);
xnor U27583 (N_27583,N_26479,N_25486);
and U27584 (N_27584,N_25714,N_25552);
or U27585 (N_27585,N_25429,N_25824);
xnor U27586 (N_27586,N_25141,N_26229);
or U27587 (N_27587,N_26586,N_27282);
nand U27588 (N_27588,N_27067,N_26155);
or U27589 (N_27589,N_25721,N_27049);
xor U27590 (N_27590,N_27098,N_26760);
and U27591 (N_27591,N_25487,N_27093);
and U27592 (N_27592,N_26051,N_26776);
nor U27593 (N_27593,N_26043,N_25026);
nand U27594 (N_27594,N_26830,N_26894);
nand U27595 (N_27595,N_27278,N_25188);
nand U27596 (N_27596,N_26943,N_26756);
and U27597 (N_27597,N_26202,N_26603);
nor U27598 (N_27598,N_26972,N_25819);
and U27599 (N_27599,N_25996,N_27027);
xor U27600 (N_27600,N_27312,N_26826);
nor U27601 (N_27601,N_26118,N_25746);
nand U27602 (N_27602,N_25813,N_26977);
xnor U27603 (N_27603,N_26572,N_25110);
xnor U27604 (N_27604,N_27347,N_25353);
or U27605 (N_27605,N_27409,N_26230);
xor U27606 (N_27606,N_25405,N_26682);
and U27607 (N_27607,N_26431,N_25692);
or U27608 (N_27608,N_26480,N_26352);
xor U27609 (N_27609,N_26521,N_25501);
nand U27610 (N_27610,N_26347,N_25585);
or U27611 (N_27611,N_27056,N_26267);
xnor U27612 (N_27612,N_26887,N_26005);
or U27613 (N_27613,N_25271,N_25182);
nand U27614 (N_27614,N_26742,N_26303);
nor U27615 (N_27615,N_25442,N_26214);
nor U27616 (N_27616,N_26778,N_26000);
xor U27617 (N_27617,N_26271,N_25324);
or U27618 (N_27618,N_25753,N_26951);
nor U27619 (N_27619,N_27116,N_26218);
and U27620 (N_27620,N_25312,N_26526);
and U27621 (N_27621,N_25659,N_25897);
or U27622 (N_27622,N_26478,N_25985);
or U27623 (N_27623,N_26388,N_27291);
nand U27624 (N_27624,N_26143,N_27316);
nor U27625 (N_27625,N_25213,N_27007);
and U27626 (N_27626,N_27102,N_25635);
or U27627 (N_27627,N_26927,N_26313);
or U27628 (N_27628,N_25265,N_25974);
nand U27629 (N_27629,N_25533,N_26401);
or U27630 (N_27630,N_26213,N_26963);
xor U27631 (N_27631,N_25596,N_26093);
nor U27632 (N_27632,N_25664,N_26305);
nand U27633 (N_27633,N_25251,N_25383);
nand U27634 (N_27634,N_26227,N_26332);
nand U27635 (N_27635,N_25745,N_26032);
and U27636 (N_27636,N_25593,N_27095);
nand U27637 (N_27637,N_25190,N_26378);
or U27638 (N_27638,N_26930,N_25666);
and U27639 (N_27639,N_25597,N_25730);
or U27640 (N_27640,N_25194,N_27339);
xnor U27641 (N_27641,N_25317,N_26693);
nor U27642 (N_27642,N_25079,N_27017);
and U27643 (N_27643,N_26483,N_25308);
nor U27644 (N_27644,N_25831,N_27111);
nand U27645 (N_27645,N_25339,N_27081);
nor U27646 (N_27646,N_26689,N_26680);
nand U27647 (N_27647,N_25990,N_25588);
nor U27648 (N_27648,N_26708,N_25602);
and U27649 (N_27649,N_26884,N_25853);
nand U27650 (N_27650,N_26866,N_25537);
and U27651 (N_27651,N_26112,N_27154);
xnor U27652 (N_27652,N_25842,N_26706);
nand U27653 (N_27653,N_27311,N_25444);
or U27654 (N_27654,N_26212,N_26241);
and U27655 (N_27655,N_26827,N_26619);
nor U27656 (N_27656,N_25476,N_27078);
nor U27657 (N_27657,N_25896,N_27080);
xnor U27658 (N_27658,N_27025,N_26833);
or U27659 (N_27659,N_25446,N_27043);
nand U27660 (N_27660,N_25800,N_26037);
nand U27661 (N_27661,N_27486,N_26512);
and U27662 (N_27662,N_25473,N_26135);
xor U27663 (N_27663,N_26027,N_25895);
or U27664 (N_27664,N_26127,N_27314);
xnor U27665 (N_27665,N_27193,N_26518);
xor U27666 (N_27666,N_27287,N_26598);
or U27667 (N_27667,N_27308,N_26817);
nand U27668 (N_27668,N_25484,N_25796);
nor U27669 (N_27669,N_25663,N_27472);
nor U27670 (N_27670,N_27134,N_27030);
nor U27671 (N_27671,N_27034,N_27085);
or U27672 (N_27672,N_26322,N_26500);
nor U27673 (N_27673,N_25623,N_25482);
xnor U27674 (N_27674,N_27270,N_25175);
xnor U27675 (N_27675,N_26028,N_27481);
and U27676 (N_27676,N_25882,N_25843);
and U27677 (N_27677,N_26176,N_27417);
nor U27678 (N_27678,N_25421,N_26272);
or U27679 (N_27679,N_26872,N_27369);
nand U27680 (N_27680,N_25977,N_27069);
and U27681 (N_27681,N_25224,N_27408);
and U27682 (N_27682,N_25894,N_25419);
nand U27683 (N_27683,N_25314,N_27000);
and U27684 (N_27684,N_26446,N_25822);
nor U27685 (N_27685,N_25416,N_26980);
nor U27686 (N_27686,N_27431,N_26735);
nand U27687 (N_27687,N_26075,N_27267);
nand U27688 (N_27688,N_25066,N_25269);
and U27689 (N_27689,N_26565,N_27439);
nand U27690 (N_27690,N_26601,N_26101);
xnor U27691 (N_27691,N_25195,N_25517);
and U27692 (N_27692,N_26221,N_26015);
or U27693 (N_27693,N_26408,N_26487);
xnor U27694 (N_27694,N_25680,N_26797);
or U27695 (N_27695,N_26179,N_26159);
nand U27696 (N_27696,N_26599,N_27169);
nand U27697 (N_27697,N_27075,N_27336);
or U27698 (N_27698,N_25058,N_26589);
xnor U27699 (N_27699,N_26783,N_26224);
and U27700 (N_27700,N_25017,N_26920);
or U27701 (N_27701,N_27054,N_26361);
and U27702 (N_27702,N_26721,N_25385);
and U27703 (N_27703,N_27253,N_25741);
and U27704 (N_27704,N_25530,N_25435);
nor U27705 (N_27705,N_25292,N_26558);
nor U27706 (N_27706,N_26880,N_26837);
xnor U27707 (N_27707,N_27264,N_26279);
or U27708 (N_27708,N_25954,N_26009);
and U27709 (N_27709,N_25710,N_27045);
and U27710 (N_27710,N_25172,N_26497);
xor U27711 (N_27711,N_25935,N_25179);
nor U27712 (N_27712,N_25737,N_26191);
or U27713 (N_27713,N_25382,N_27269);
xor U27714 (N_27714,N_26704,N_27129);
and U27715 (N_27715,N_27242,N_27361);
nor U27716 (N_27716,N_26768,N_26461);
or U27717 (N_27717,N_25720,N_25860);
xnor U27718 (N_27718,N_25313,N_27458);
nor U27719 (N_27719,N_26942,N_27497);
or U27720 (N_27720,N_26377,N_26834);
nor U27721 (N_27721,N_26206,N_25402);
xor U27722 (N_27722,N_26353,N_25957);
nor U27723 (N_27723,N_25526,N_25000);
nand U27724 (N_27724,N_26412,N_26785);
nor U27725 (N_27725,N_27418,N_25539);
xor U27726 (N_27726,N_26163,N_25829);
nor U27727 (N_27727,N_25071,N_25433);
nand U27728 (N_27728,N_25950,N_25163);
nor U27729 (N_27729,N_26198,N_25560);
nor U27730 (N_27730,N_26083,N_26383);
and U27731 (N_27731,N_27171,N_27149);
or U27732 (N_27732,N_25916,N_25891);
nor U27733 (N_27733,N_25589,N_25936);
nor U27734 (N_27734,N_26391,N_26304);
and U27735 (N_27735,N_26885,N_25726);
xor U27736 (N_27736,N_26758,N_26338);
xor U27737 (N_27737,N_25260,N_27490);
nand U27738 (N_27738,N_25396,N_25003);
nand U27739 (N_27739,N_27107,N_25638);
nand U27740 (N_27740,N_25052,N_26307);
or U27741 (N_27741,N_25927,N_26533);
or U27742 (N_27742,N_26843,N_26277);
or U27743 (N_27743,N_25158,N_25478);
nand U27744 (N_27744,N_26720,N_27322);
and U27745 (N_27745,N_25047,N_25756);
nor U27746 (N_27746,N_27212,N_26319);
nor U27747 (N_27747,N_26362,N_27271);
nand U27748 (N_27748,N_26892,N_26808);
nand U27749 (N_27749,N_27175,N_26190);
and U27750 (N_27750,N_26566,N_25493);
xnor U27751 (N_27751,N_26275,N_26038);
and U27752 (N_27752,N_26968,N_25032);
nand U27753 (N_27753,N_27342,N_25529);
or U27754 (N_27754,N_25516,N_26626);
xnor U27755 (N_27755,N_25681,N_25912);
xnor U27756 (N_27756,N_25827,N_27100);
and U27757 (N_27757,N_26934,N_27252);
and U27758 (N_27758,N_25817,N_27162);
nand U27759 (N_27759,N_25321,N_27241);
nor U27760 (N_27760,N_27443,N_26635);
nand U27761 (N_27761,N_27261,N_26284);
or U27762 (N_27762,N_25112,N_25976);
xor U27763 (N_27763,N_27407,N_25341);
or U27764 (N_27764,N_27170,N_26255);
xnor U27765 (N_27765,N_27304,N_26099);
nand U27766 (N_27766,N_26354,N_27018);
nand U27767 (N_27767,N_25427,N_26136);
and U27768 (N_27768,N_25454,N_27106);
xor U27769 (N_27769,N_27079,N_25972);
and U27770 (N_27770,N_26749,N_27213);
and U27771 (N_27771,N_27065,N_26936);
nor U27772 (N_27772,N_25392,N_26281);
or U27773 (N_27773,N_26138,N_25379);
or U27774 (N_27774,N_26301,N_26596);
nor U27775 (N_27775,N_25543,N_27276);
and U27776 (N_27776,N_25766,N_25147);
xor U27777 (N_27777,N_25226,N_25709);
nand U27778 (N_27778,N_25101,N_26430);
or U27779 (N_27779,N_26851,N_26926);
nor U27780 (N_27780,N_25471,N_26748);
or U27781 (N_27781,N_26949,N_26703);
nor U27782 (N_27782,N_25143,N_26839);
xor U27783 (N_27783,N_25403,N_26197);
or U27784 (N_27784,N_26091,N_27295);
and U27785 (N_27785,N_26450,N_25291);
or U27786 (N_27786,N_25915,N_25610);
and U27787 (N_27787,N_26771,N_25126);
xnor U27788 (N_27788,N_26723,N_27084);
xor U27789 (N_27789,N_25634,N_26899);
nor U27790 (N_27790,N_27097,N_25691);
or U27791 (N_27791,N_26342,N_27415);
xor U27792 (N_27792,N_25013,N_25485);
nor U27793 (N_27793,N_26979,N_26288);
xor U27794 (N_27794,N_25459,N_27478);
nand U27795 (N_27795,N_26489,N_25719);
or U27796 (N_27796,N_26929,N_25470);
xnor U27797 (N_27797,N_26121,N_26587);
nor U27798 (N_27798,N_25281,N_26781);
xor U27799 (N_27799,N_27058,N_27413);
nor U27800 (N_27800,N_27037,N_25969);
xnor U27801 (N_27801,N_25045,N_25508);
xor U27802 (N_27802,N_25279,N_26064);
xnor U27803 (N_27803,N_25388,N_26650);
and U27804 (N_27804,N_26139,N_25278);
or U27805 (N_27805,N_26261,N_25348);
and U27806 (N_27806,N_27112,N_26459);
nand U27807 (N_27807,N_27210,N_26046);
or U27808 (N_27808,N_27023,N_25735);
or U27809 (N_27809,N_25189,N_26078);
and U27810 (N_27810,N_26335,N_26346);
and U27811 (N_27811,N_26130,N_25648);
nand U27812 (N_27812,N_25333,N_25650);
nor U27813 (N_27813,N_25542,N_26759);
and U27814 (N_27814,N_26096,N_25601);
xor U27815 (N_27815,N_26593,N_25049);
nor U27816 (N_27816,N_25285,N_27425);
nor U27817 (N_27817,N_26517,N_26178);
and U27818 (N_27818,N_25948,N_25582);
and U27819 (N_27819,N_25113,N_25305);
or U27820 (N_27820,N_25165,N_26103);
and U27821 (N_27821,N_26004,N_25039);
nand U27822 (N_27822,N_25315,N_25641);
nor U27823 (N_27823,N_26310,N_25608);
nand U27824 (N_27824,N_27281,N_25234);
nand U27825 (N_27825,N_25577,N_25792);
nor U27826 (N_27826,N_26247,N_25103);
nor U27827 (N_27827,N_25247,N_27118);
nand U27828 (N_27828,N_27370,N_25932);
nand U27829 (N_27829,N_26974,N_27142);
or U27830 (N_27830,N_25378,N_26597);
nor U27831 (N_27831,N_26829,N_26813);
and U27832 (N_27832,N_26505,N_26413);
xor U27833 (N_27833,N_25318,N_25335);
or U27834 (N_27834,N_25795,N_26766);
and U27835 (N_27835,N_27195,N_26617);
and U27836 (N_27836,N_27484,N_26035);
and U27837 (N_27837,N_25465,N_25157);
xor U27838 (N_27838,N_25077,N_25080);
or U27839 (N_27839,N_25227,N_26490);
or U27840 (N_27840,N_26888,N_26527);
xor U27841 (N_27841,N_25061,N_25706);
nor U27842 (N_27842,N_26034,N_26950);
nor U27843 (N_27843,N_26540,N_26171);
nand U27844 (N_27844,N_27426,N_27392);
nand U27845 (N_27845,N_26546,N_27127);
nor U27846 (N_27846,N_25391,N_27070);
nor U27847 (N_27847,N_25220,N_26510);
nand U27848 (N_27848,N_26256,N_26330);
nand U27849 (N_27849,N_25105,N_26832);
nand U27850 (N_27850,N_27255,N_25642);
xor U27851 (N_27851,N_26321,N_26800);
and U27852 (N_27852,N_25092,N_26696);
and U27853 (N_27853,N_25358,N_26793);
xor U27854 (N_27854,N_26665,N_27217);
nand U27855 (N_27855,N_25073,N_27248);
and U27856 (N_27856,N_26339,N_25288);
and U27857 (N_27857,N_25629,N_25674);
xor U27858 (N_27858,N_26196,N_25196);
xor U27859 (N_27859,N_25261,N_26554);
or U27860 (N_27860,N_25009,N_25697);
xnor U27861 (N_27861,N_27327,N_27186);
or U27862 (N_27862,N_26645,N_25369);
nand U27863 (N_27863,N_26690,N_26327);
xnor U27864 (N_27864,N_26410,N_26909);
and U27865 (N_27865,N_27404,N_25612);
nand U27866 (N_27866,N_25980,N_25970);
nand U27867 (N_27867,N_26999,N_26678);
or U27868 (N_27868,N_25469,N_26020);
nor U27869 (N_27869,N_25447,N_26111);
or U27870 (N_27870,N_26368,N_27235);
nand U27871 (N_27871,N_25776,N_25750);
xor U27872 (N_27872,N_26867,N_26337);
nor U27873 (N_27873,N_25397,N_25764);
and U27874 (N_27874,N_26157,N_25239);
nor U27875 (N_27875,N_26454,N_25249);
and U27876 (N_27876,N_26782,N_26804);
nor U27877 (N_27877,N_25836,N_26891);
xnor U27878 (N_27878,N_25332,N_25043);
xor U27879 (N_27879,N_26550,N_26613);
xor U27880 (N_27880,N_25576,N_25214);
and U27881 (N_27881,N_25100,N_26711);
nand U27882 (N_27882,N_25283,N_26873);
or U27883 (N_27883,N_25893,N_26294);
and U27884 (N_27884,N_26393,N_25276);
and U27885 (N_27885,N_26795,N_27236);
xnor U27886 (N_27886,N_25005,N_27135);
or U27887 (N_27887,N_25803,N_25743);
xor U27888 (N_27888,N_26567,N_25877);
xnor U27889 (N_27889,N_26799,N_27284);
nor U27890 (N_27890,N_26059,N_26753);
and U27891 (N_27891,N_26396,N_25708);
nor U27892 (N_27892,N_25694,N_26007);
and U27893 (N_27893,N_25488,N_25183);
or U27894 (N_27894,N_26541,N_26146);
nand U27895 (N_27895,N_27485,N_26745);
nor U27896 (N_27896,N_26283,N_27207);
nand U27897 (N_27897,N_26369,N_26405);
nand U27898 (N_27898,N_26719,N_27468);
nand U27899 (N_27899,N_26955,N_27216);
and U27900 (N_27900,N_26148,N_25164);
or U27901 (N_27901,N_26150,N_25928);
nand U27902 (N_27902,N_26636,N_27405);
and U27903 (N_27903,N_26246,N_25657);
and U27904 (N_27904,N_27279,N_25181);
and U27905 (N_27905,N_26810,N_25633);
xor U27906 (N_27906,N_25068,N_26675);
xor U27907 (N_27907,N_26382,N_26925);
nor U27908 (N_27908,N_25581,N_26710);
xor U27909 (N_27909,N_25952,N_27200);
and U27910 (N_27910,N_25170,N_25472);
xor U27911 (N_27911,N_27320,N_27341);
xor U27912 (N_27912,N_25084,N_26055);
or U27913 (N_27913,N_25684,N_27187);
xnor U27914 (N_27914,N_27325,N_27437);
nor U27915 (N_27915,N_25607,N_27019);
nor U27916 (N_27916,N_27300,N_25761);
nand U27917 (N_27917,N_25807,N_25769);
or U27918 (N_27918,N_25578,N_25240);
and U27919 (N_27919,N_26060,N_25622);
or U27920 (N_27920,N_26110,N_25546);
and U27921 (N_27921,N_25127,N_26661);
nand U27922 (N_27922,N_27233,N_26850);
or U27923 (N_27923,N_25778,N_25152);
or U27924 (N_27924,N_27087,N_25738);
or U27925 (N_27925,N_26156,N_25330);
or U27926 (N_27926,N_25672,N_26724);
nor U27927 (N_27927,N_26491,N_25587);
nor U27928 (N_27928,N_26309,N_27167);
or U27929 (N_27929,N_26595,N_26142);
nand U27930 (N_27930,N_25225,N_26298);
xnor U27931 (N_27931,N_26002,N_25266);
nand U27932 (N_27932,N_25137,N_26688);
nand U27933 (N_27933,N_27372,N_25280);
or U27934 (N_27934,N_26504,N_27318);
xnor U27935 (N_27935,N_25949,N_25413);
or U27936 (N_27936,N_25430,N_25490);
or U27937 (N_27937,N_25857,N_25089);
and U27938 (N_27938,N_26580,N_26411);
xnor U27939 (N_27939,N_27203,N_25604);
xor U27940 (N_27940,N_26425,N_25222);
nor U27941 (N_27941,N_27332,N_26258);
and U27942 (N_27942,N_26080,N_26054);
nor U27943 (N_27943,N_27411,N_26903);
and U27944 (N_27944,N_26462,N_27324);
nor U27945 (N_27945,N_26215,N_25975);
nand U27946 (N_27946,N_25171,N_27113);
xnor U27947 (N_27947,N_25632,N_25984);
xor U27948 (N_27948,N_25620,N_25572);
or U27949 (N_27949,N_26209,N_25108);
and U27950 (N_27950,N_25540,N_27161);
nor U27951 (N_27951,N_26622,N_25565);
nand U27952 (N_27952,N_25828,N_26583);
nand U27953 (N_27953,N_25945,N_26875);
xor U27954 (N_27954,N_26707,N_27368);
or U27955 (N_27955,N_26528,N_26219);
or U27956 (N_27956,N_26564,N_25723);
nand U27957 (N_27957,N_26278,N_25799);
or U27958 (N_27958,N_25329,N_26845);
or U27959 (N_27959,N_27277,N_25094);
nand U27960 (N_27960,N_26824,N_25739);
or U27961 (N_27961,N_25018,N_26529);
nand U27962 (N_27962,N_26422,N_25740);
and U27963 (N_27963,N_27428,N_26097);
and U27964 (N_27964,N_27032,N_25489);
xor U27965 (N_27965,N_27001,N_25368);
xor U27966 (N_27966,N_27362,N_26652);
nand U27967 (N_27967,N_26831,N_27401);
nand U27968 (N_27968,N_27382,N_25216);
or U27969 (N_27969,N_25114,N_26575);
nor U27970 (N_27970,N_25699,N_25931);
or U27971 (N_27971,N_26344,N_25168);
nand U27972 (N_27972,N_26117,N_25233);
and U27973 (N_27973,N_25645,N_26068);
or U27974 (N_27974,N_25599,N_26961);
nand U27975 (N_27975,N_25051,N_25614);
nor U27976 (N_27976,N_25784,N_25423);
nand U27977 (N_27977,N_27310,N_25956);
nor U27978 (N_27978,N_26058,N_27495);
nand U27979 (N_27979,N_25781,N_25628);
nor U27980 (N_27980,N_27143,N_27003);
nor U27981 (N_27981,N_26225,N_26686);
or U27982 (N_27982,N_25404,N_25744);
and U27983 (N_27983,N_25426,N_25921);
nor U27984 (N_27984,N_25410,N_26390);
nand U27985 (N_27985,N_26772,N_26553);
nor U27986 (N_27986,N_26578,N_25217);
nand U27987 (N_27987,N_26025,N_25673);
nor U27988 (N_27988,N_25892,N_25671);
and U27989 (N_27989,N_26475,N_26276);
nor U27990 (N_27990,N_26809,N_25257);
nor U27991 (N_27991,N_26416,N_26081);
or U27992 (N_27992,N_25218,N_25630);
and U27993 (N_27993,N_26013,N_25512);
xnor U27994 (N_27994,N_27338,N_26147);
xnor U27995 (N_27995,N_26610,N_25497);
nand U27996 (N_27996,N_25509,N_26729);
nor U27997 (N_27997,N_26042,N_26513);
nor U27998 (N_27998,N_25545,N_26556);
nor U27999 (N_27999,N_25826,N_27356);
and U28000 (N_28000,N_25906,N_25056);
nand U28001 (N_28001,N_26835,N_25480);
and U28002 (N_28002,N_25751,N_26287);
nand U28003 (N_28003,N_27121,N_26854);
nor U28004 (N_28004,N_26592,N_26095);
nor U28005 (N_28005,N_27303,N_27293);
or U28006 (N_28006,N_27317,N_25498);
or U28007 (N_28007,N_25728,N_27289);
or U28008 (N_28008,N_26644,N_27487);
nor U28009 (N_28009,N_26838,N_25809);
xor U28010 (N_28010,N_25406,N_26474);
or U28011 (N_28011,N_26265,N_25351);
xor U28012 (N_28012,N_25337,N_26902);
nand U28013 (N_28013,N_27052,N_25564);
nor U28014 (N_28014,N_27456,N_25145);
xnor U28015 (N_28015,N_26655,N_27346);
or U28016 (N_28016,N_25504,N_25371);
and U28017 (N_28017,N_26988,N_25046);
xnor U28018 (N_28018,N_25010,N_27496);
nand U28019 (N_28019,N_27273,N_25676);
nand U28020 (N_28020,N_25982,N_26030);
or U28021 (N_28021,N_26632,N_26286);
and U28022 (N_28022,N_25463,N_26982);
nor U28023 (N_28023,N_27453,N_27060);
nand U28024 (N_28024,N_25967,N_26254);
nor U28025 (N_28025,N_26577,N_26666);
xor U28026 (N_28026,N_26788,N_27449);
nor U28027 (N_28027,N_27180,N_25322);
and U28028 (N_28028,N_25944,N_26801);
or U28029 (N_28029,N_26300,N_25357);
nand U28030 (N_28030,N_25722,N_26228);
xnor U28031 (N_28031,N_26923,N_26372);
nor U28032 (N_28032,N_25422,N_27463);
and U28033 (N_28033,N_26021,N_26789);
nor U28034 (N_28034,N_27124,N_25788);
and U28035 (N_28035,N_26188,N_27064);
or U28036 (N_28036,N_25771,N_26714);
xnor U28037 (N_28037,N_26360,N_26177);
and U28038 (N_28038,N_26394,N_27321);
or U28039 (N_28039,N_25643,N_25028);
xor U28040 (N_28040,N_25107,N_25262);
nand U28041 (N_28041,N_25373,N_25919);
or U28042 (N_28042,N_26498,N_25991);
nand U28043 (N_28043,N_25186,N_26876);
xnor U28044 (N_28044,N_25849,N_26175);
and U28045 (N_28045,N_25787,N_25524);
or U28046 (N_28046,N_25119,N_26898);
nor U28047 (N_28047,N_25538,N_27451);
or U28048 (N_28048,N_26798,N_27375);
nor U28049 (N_28049,N_25015,N_25268);
xor U28050 (N_28050,N_26609,N_26399);
nor U28051 (N_28051,N_27197,N_25683);
nand U28052 (N_28052,N_25120,N_26011);
and U28053 (N_28053,N_25639,N_26791);
and U28054 (N_28054,N_27268,N_25023);
nand U28055 (N_28055,N_25729,N_26089);
and U28056 (N_28056,N_25611,N_27454);
xnor U28057 (N_28057,N_25208,N_27272);
or U28058 (N_28058,N_26435,N_26123);
nor U28059 (N_28059,N_26944,N_26722);
nor U28060 (N_28060,N_26812,N_25559);
and U28061 (N_28061,N_26743,N_26419);
or U28062 (N_28062,N_25765,N_26663);
nand U28063 (N_28063,N_27266,N_26242);
xnor U28064 (N_28064,N_27299,N_25193);
nor U28065 (N_28065,N_26555,N_26174);
xor U28066 (N_28066,N_25525,N_26879);
or U28067 (N_28067,N_26741,N_26585);
or U28068 (N_28068,N_26915,N_26681);
or U28069 (N_28069,N_26010,N_26251);
and U28070 (N_28070,N_26822,N_25059);
nand U28071 (N_28071,N_26297,N_25377);
nand U28072 (N_28072,N_25088,N_27145);
xnor U28073 (N_28073,N_25275,N_25965);
or U28074 (N_28074,N_25670,N_26193);
nor U28075 (N_28075,N_25903,N_26260);
nor U28076 (N_28076,N_25557,N_26226);
xor U28077 (N_28077,N_26536,N_27138);
nand U28078 (N_28078,N_26886,N_26557);
xnor U28079 (N_28079,N_25338,N_25782);
or U28080 (N_28080,N_25924,N_26239);
xor U28081 (N_28081,N_25631,N_26869);
nor U28082 (N_28082,N_27351,N_27250);
and U28083 (N_28083,N_25400,N_25617);
xor U28084 (N_28084,N_26180,N_27215);
and U28085 (N_28085,N_26145,N_25282);
nor U28086 (N_28086,N_26340,N_27035);
xnor U28087 (N_28087,N_26253,N_27459);
nand U28088 (N_28088,N_25310,N_25255);
xor U28089 (N_28089,N_25349,N_25693);
nor U28090 (N_28090,N_26460,N_25832);
or U28091 (N_28091,N_26713,N_25647);
or U28092 (N_28092,N_26559,N_25354);
nor U28093 (N_28093,N_26223,N_25570);
nor U28094 (N_28094,N_26752,N_25492);
xnor U28095 (N_28095,N_26992,N_27220);
or U28096 (N_28096,N_27051,N_26700);
xor U28097 (N_28097,N_26847,N_26434);
and U28098 (N_28098,N_25252,N_27384);
xnor U28099 (N_28099,N_25197,N_25245);
xnor U28100 (N_28100,N_27345,N_25941);
and U28101 (N_28101,N_25839,N_26954);
or U28102 (N_28102,N_25838,N_27390);
nand U28103 (N_28103,N_27191,N_25139);
xor U28104 (N_28104,N_25284,N_26731);
nor U28105 (N_28105,N_25131,N_25815);
xor U28106 (N_28106,N_27168,N_26836);
nor U28107 (N_28107,N_27126,N_25995);
nand U28108 (N_28108,N_25762,N_27038);
nand U28109 (N_28109,N_26238,N_25238);
or U28110 (N_28110,N_27114,N_27004);
nor U28111 (N_28111,N_25591,N_26668);
and U28112 (N_28112,N_25615,N_27315);
or U28113 (N_28113,N_26893,N_26417);
nor U28114 (N_28114,N_25342,N_25389);
nand U28115 (N_28115,N_26170,N_26821);
xor U28116 (N_28116,N_25528,N_25507);
or U28117 (N_28117,N_27011,N_25865);
and U28118 (N_28118,N_26119,N_25888);
and U28119 (N_28119,N_25869,N_27227);
and U28120 (N_28120,N_26094,N_26744);
nor U28121 (N_28121,N_27447,N_25095);
nand U28122 (N_28122,N_26065,N_25812);
and U28123 (N_28123,N_27194,N_27476);
nand U28124 (N_28124,N_26323,N_27189);
and U28125 (N_28125,N_26698,N_26849);
xor U28126 (N_28126,N_25445,N_27343);
or U28127 (N_28127,N_26216,N_25759);
xnor U28128 (N_28128,N_26090,N_26203);
xor U28129 (N_28129,N_27159,N_26908);
nor U28130 (N_28130,N_25142,N_26029);
nor U28131 (N_28131,N_26076,N_26662);
or U28132 (N_28132,N_26349,N_25922);
or U28133 (N_28133,N_27442,N_27290);
xor U28134 (N_28134,N_25598,N_25267);
or U28135 (N_28135,N_25072,N_27286);
xnor U28136 (N_28136,N_26165,N_26328);
or U28137 (N_28137,N_25198,N_25558);
or U28138 (N_28138,N_26642,N_25549);
nand U28139 (N_28139,N_26590,N_26457);
nand U28140 (N_28140,N_25253,N_25868);
nor U28141 (N_28141,N_25102,N_26493);
nand U28142 (N_28142,N_25082,N_26024);
nor U28143 (N_28143,N_27258,N_25063);
nor U28144 (N_28144,N_26786,N_25551);
and U28145 (N_28145,N_26331,N_27139);
and U28146 (N_28146,N_26631,N_25534);
or U28147 (N_28147,N_27128,N_27329);
and U28148 (N_28148,N_25651,N_26794);
xnor U28149 (N_28149,N_25675,N_25658);
nand U28150 (N_28150,N_25129,N_25412);
and U28151 (N_28151,N_26608,N_26701);
and U28152 (N_28152,N_25797,N_26853);
nand U28153 (N_28153,N_25370,N_27298);
or U28154 (N_28154,N_25627,N_26857);
nand U28155 (N_28155,N_26131,N_25178);
xor U28156 (N_28156,N_26240,N_25115);
xnor U28157 (N_28157,N_26439,N_27108);
nand U28158 (N_28158,N_25019,N_26074);
or U28159 (N_28159,N_26115,N_26315);
or U28160 (N_28160,N_27256,N_27110);
or U28161 (N_28161,N_26440,N_27123);
or U28162 (N_28162,N_26100,N_27165);
nand U28163 (N_28163,N_26506,N_26048);
nand U28164 (N_28164,N_26981,N_25793);
nor U28165 (N_28165,N_27119,N_27074);
xor U28166 (N_28166,N_27148,N_27441);
or U28167 (N_28167,N_26195,N_27288);
and U28168 (N_28168,N_25758,N_26334);
or U28169 (N_28169,N_25287,N_27173);
and U28170 (N_28170,N_26922,N_25259);
and U28171 (N_28171,N_26268,N_26210);
xnor U28172 (N_28172,N_26379,N_25098);
nor U28173 (N_28173,N_27474,N_27101);
or U28174 (N_28174,N_25054,N_27020);
and U28175 (N_28175,N_27262,N_27328);
nand U28176 (N_28176,N_27246,N_25754);
xnor U28177 (N_28177,N_25180,N_26077);
xnor U28178 (N_28178,N_25987,N_26576);
and U28179 (N_28179,N_25340,N_25616);
xor U28180 (N_28180,N_26933,N_26784);
or U28181 (N_28181,N_26581,N_26105);
and U28182 (N_28182,N_25522,N_25012);
nand U28183 (N_28183,N_26499,N_26144);
and U28184 (N_28184,N_25520,N_25149);
or U28185 (N_28185,N_27444,N_25665);
nor U28186 (N_28186,N_25686,N_25742);
nor U28187 (N_28187,N_26451,N_25978);
and U28188 (N_28188,N_25513,N_27358);
and U28189 (N_28189,N_25160,N_25374);
nand U28190 (N_28190,N_25715,N_26400);
and U28191 (N_28191,N_27414,N_27181);
and U28192 (N_28192,N_27306,N_26947);
nor U28193 (N_28193,N_25106,N_26616);
nor U28194 (N_28194,N_25030,N_25304);
nor U28195 (N_28195,N_26201,N_26990);
nand U28196 (N_28196,N_27424,N_26485);
and U28197 (N_28197,N_25025,N_27410);
and U28198 (N_28198,N_26767,N_25942);
xnor U28199 (N_28199,N_25503,N_26259);
nor U28200 (N_28200,N_26897,N_27179);
nor U28201 (N_28201,N_26856,N_26161);
or U28202 (N_28202,N_26436,N_25161);
or U28203 (N_28203,N_27419,N_26252);
and U28204 (N_28204,N_26124,N_25230);
or U28205 (N_28205,N_25311,N_25875);
xor U28206 (N_28206,N_26725,N_26780);
or U28207 (N_28207,N_25855,N_27082);
xnor U28208 (N_28208,N_25835,N_26120);
nor U28209 (N_28209,N_25117,N_26257);
nor U28210 (N_28210,N_27462,N_26200);
or U28211 (N_28211,N_25494,N_25394);
and U28212 (N_28212,N_25235,N_27344);
nor U28213 (N_28213,N_25555,N_25097);
xor U28214 (N_28214,N_26709,N_27218);
nand U28215 (N_28215,N_27006,N_25122);
nand U28216 (N_28216,N_26594,N_25236);
and U28217 (N_28217,N_26364,N_26989);
nand U28218 (N_28218,N_25859,N_26295);
xnor U28219 (N_28219,N_25256,N_25514);
nor U28220 (N_28220,N_26660,N_25460);
nor U28221 (N_28221,N_25983,N_25515);
nor U28222 (N_28222,N_26848,N_27491);
xnor U28223 (N_28223,N_25688,N_27445);
and U28224 (N_28224,N_27319,N_26790);
nor U28225 (N_28225,N_27105,N_26871);
nand U28226 (N_28226,N_26270,N_26840);
nor U28227 (N_28227,N_25858,N_25133);
nand U28228 (N_28228,N_26343,N_25847);
and U28229 (N_28229,N_26185,N_26890);
nor U28230 (N_28230,N_26233,N_25968);
xnor U28231 (N_28231,N_26673,N_27090);
or U28232 (N_28232,N_25136,N_26946);
xor U28233 (N_28233,N_26445,N_26082);
nor U28234 (N_28234,N_27430,N_27479);
or U28235 (N_28235,N_26984,N_25652);
nand U28236 (N_28236,N_25992,N_26423);
or U28237 (N_28237,N_26584,N_27202);
nand U28238 (N_28238,N_27387,N_25569);
and U28239 (N_28239,N_25801,N_25810);
nand U28240 (N_28240,N_25901,N_26629);
and U28241 (N_28241,N_27150,N_26472);
nor U28242 (N_28242,N_26073,N_27480);
nor U28243 (N_28243,N_26066,N_25034);
nand U28244 (N_28244,N_27452,N_26905);
or U28245 (N_28245,N_27251,N_26859);
xor U28246 (N_28246,N_27136,N_26820);
nand U28247 (N_28247,N_26542,N_25532);
and U28248 (N_28248,N_25062,N_26814);
xnor U28249 (N_28249,N_26779,N_26481);
nand U28250 (N_28250,N_26363,N_27475);
xor U28251 (N_28251,N_25096,N_25571);
nor U28252 (N_28252,N_26311,N_27103);
nor U28253 (N_28253,N_26965,N_25907);
or U28254 (N_28254,N_25364,N_25083);
nand U28255 (N_28255,N_25971,N_26003);
xor U28256 (N_28256,N_26033,N_27130);
nor U28257 (N_28257,N_25736,N_25355);
or U28258 (N_28258,N_26916,N_25258);
nor U28259 (N_28259,N_27471,N_25625);
and U28260 (N_28260,N_27265,N_27436);
xor U28261 (N_28261,N_25086,N_27188);
nand U28262 (N_28262,N_25879,N_27348);
and U28263 (N_28263,N_26324,N_25206);
nand U28264 (N_28264,N_27381,N_26918);
nor U28265 (N_28265,N_26733,N_27323);
or U28266 (N_28266,N_27063,N_26878);
or U28267 (N_28267,N_27089,N_27400);
nand U28268 (N_28268,N_26966,N_27209);
nand U28269 (N_28269,N_27305,N_27039);
nor U28270 (N_28270,N_25210,N_26667);
nor U28271 (N_28271,N_27092,N_26691);
xnor U28272 (N_28272,N_25124,N_27015);
nand U28273 (N_28273,N_26385,N_27048);
nand U28274 (N_28274,N_26630,N_25134);
nand U28275 (N_28275,N_25461,N_26716);
nor U28276 (N_28276,N_27066,N_25911);
xnor U28277 (N_28277,N_25033,N_26151);
or U28278 (N_28278,N_26648,N_25687);
or U28279 (N_28279,N_26910,N_27055);
nand U28280 (N_28280,N_25074,N_26825);
and U28281 (N_28281,N_26604,N_25527);
or U28282 (N_28282,N_26326,N_27155);
xor U28283 (N_28283,N_26736,N_25519);
and U28284 (N_28284,N_25649,N_25500);
xor U28285 (N_28285,N_26359,N_25201);
nor U28286 (N_28286,N_25099,N_26523);
xnor U28287 (N_28287,N_25732,N_26960);
or U28288 (N_28288,N_25148,N_25821);
nor U28289 (N_28289,N_25966,N_26102);
nand U28290 (N_28290,N_26348,N_27137);
nor U28291 (N_28291,N_25554,N_26548);
xor U28292 (N_28292,N_27467,N_26792);
and U28293 (N_28293,N_26222,N_25048);
and U28294 (N_28294,N_27132,N_27352);
and U28295 (N_28295,N_25904,N_26970);
nand U28296 (N_28296,N_26488,N_25556);
or U28297 (N_28297,N_26409,N_27033);
or U28298 (N_28298,N_25307,N_25169);
or U28299 (N_28299,N_26674,N_25702);
and U28300 (N_28300,N_25438,N_25908);
nand U28301 (N_28301,N_25135,N_25457);
or U28302 (N_28302,N_27309,N_27260);
and U28303 (N_28303,N_27420,N_25042);
nor U28304 (N_28304,N_26991,N_26803);
nand U28305 (N_28305,N_25913,N_26621);
and U28306 (N_28306,N_25568,N_27229);
nand U28307 (N_28307,N_26402,N_25943);
and U28308 (N_28308,N_25362,N_26726);
nand U28309 (N_28309,N_25499,N_26524);
xor U28310 (N_28310,N_26107,N_27301);
nand U28311 (N_28311,N_25763,N_26469);
or U28312 (N_28312,N_25231,N_25293);
xnor U28313 (N_28313,N_26519,N_27469);
or U28314 (N_28314,N_26628,N_26071);
nand U28315 (N_28315,N_25646,N_25899);
and U28316 (N_28316,N_27192,N_25352);
nor U28317 (N_28317,N_25346,N_26732);
xnor U28318 (N_28318,N_26679,N_26494);
nor U28319 (N_28319,N_27333,N_27224);
and U28320 (N_28320,N_26292,N_27012);
nand U28321 (N_28321,N_26106,N_25690);
xnor U28322 (N_28322,N_25777,N_25244);
nand U28323 (N_28323,N_27247,N_25786);
xor U28324 (N_28324,N_25081,N_26187);
xor U28325 (N_28325,N_25704,N_25154);
nor U28326 (N_28326,N_25887,N_25848);
xnor U28327 (N_28327,N_26373,N_26978);
and U28328 (N_28328,N_25725,N_26122);
and U28329 (N_28329,N_26570,N_25237);
xnor U28330 (N_28330,N_25187,N_26012);
nand U28331 (N_28331,N_26600,N_25613);
nand U28332 (N_28332,N_27403,N_25951);
and U28333 (N_28333,N_26612,N_26486);
nor U28334 (N_28334,N_25219,N_25820);
or U28335 (N_28335,N_25483,N_25041);
xnor U28336 (N_28336,N_27190,N_25398);
nor U28337 (N_28337,N_26921,N_27184);
nor U28338 (N_28338,N_26568,N_26858);
xor U28339 (N_28339,N_26415,N_25852);
and U28340 (N_28340,N_25040,N_26746);
nand U28341 (N_28341,N_27374,N_25331);
xor U28342 (N_28342,N_26770,N_25550);
and U28343 (N_28343,N_27402,N_25656);
nor U28344 (N_28344,N_25345,N_25938);
and U28345 (N_28345,N_25481,N_26466);
nand U28346 (N_28346,N_27259,N_26314);
xnor U28347 (N_28347,N_25343,N_26371);
nand U28348 (N_28348,N_26079,N_26456);
nand U28349 (N_28349,N_26868,N_25518);
nor U28350 (N_28350,N_27450,N_27394);
and U28351 (N_28351,N_26649,N_25850);
xnor U28352 (N_28352,N_26560,N_25409);
xor U28353 (N_28353,N_25401,N_26865);
nand U28354 (N_28354,N_26958,N_25440);
xor U28355 (N_28355,N_25886,N_27363);
and U28356 (N_28356,N_26484,N_25833);
and U28357 (N_28357,N_25151,N_26511);
nand U28358 (N_28358,N_25361,N_25521);
or U28359 (N_28359,N_26173,N_27359);
and U28360 (N_28360,N_27163,N_25562);
nor U28361 (N_28361,N_27047,N_26312);
nor U28362 (N_28362,N_26182,N_26356);
or U28363 (N_28363,N_26881,N_25606);
nor U28364 (N_28364,N_26168,N_25076);
xor U28365 (N_28365,N_26014,N_25050);
xnor U28366 (N_28366,N_26467,N_27072);
and U28367 (N_28367,N_26676,N_27239);
nand U28368 (N_28368,N_26067,N_25814);
xnor U28369 (N_28369,N_26172,N_27198);
or U28370 (N_28370,N_26877,N_26160);
or U28371 (N_28371,N_27016,N_26734);
or U28372 (N_28372,N_25677,N_26448);
nor U28373 (N_28373,N_26358,N_26657);
nand U28374 (N_28374,N_25679,N_27204);
and U28375 (N_28375,N_27206,N_27196);
xor U28376 (N_28376,N_27435,N_26205);
or U28377 (N_28377,N_25805,N_26006);
or U28378 (N_28378,N_26217,N_25434);
or U28379 (N_28379,N_25689,N_27146);
xor U28380 (N_28380,N_26282,N_26468);
xor U28381 (N_28381,N_25036,N_27488);
nand U28382 (N_28382,N_25431,N_26614);
nand U28383 (N_28383,N_25707,N_25209);
nor U28384 (N_28384,N_26039,N_27061);
nor U28385 (N_28385,N_26532,N_26762);
or U28386 (N_28386,N_25479,N_26424);
or U28387 (N_28387,N_25301,N_26291);
nand U28388 (N_28388,N_25573,N_25411);
nor U28389 (N_28389,N_27340,N_26846);
xor U28390 (N_28390,N_26263,N_26647);
xnor U28391 (N_28391,N_26520,N_27174);
or U28392 (N_28392,N_27010,N_25159);
nand U28393 (N_28393,N_26333,N_27144);
nand U28394 (N_28394,N_25823,N_25156);
xor U28395 (N_28395,N_26428,N_26973);
or U28396 (N_28396,N_26274,N_26152);
xnor U28397 (N_28397,N_25958,N_25248);
xor U28398 (N_28398,N_26634,N_25731);
and U28399 (N_28399,N_27330,N_25955);
or U28400 (N_28400,N_26844,N_26199);
nor U28401 (N_28401,N_25505,N_26551);
xnor U28402 (N_28402,N_27244,N_27254);
nand U28403 (N_28403,N_26245,N_26664);
nand U28404 (N_28404,N_26697,N_25243);
nand U28405 (N_28405,N_25873,N_25594);
and U28406 (N_28406,N_26086,N_25789);
and U28407 (N_28407,N_26398,N_26862);
nor U28408 (N_28408,N_25636,N_25856);
xnor U28409 (N_28409,N_26941,N_26184);
or U28410 (N_28410,N_26874,N_26427);
xor U28411 (N_28411,N_25390,N_25111);
or U28412 (N_28412,N_26754,N_27158);
nor U28413 (N_28413,N_26380,N_26207);
and U28414 (N_28414,N_26705,N_25898);
and U28415 (N_28415,N_26640,N_27028);
nand U28416 (N_28416,N_26739,N_25712);
or U28417 (N_28417,N_25678,N_27275);
or U28418 (N_28418,N_25027,N_25696);
or U28419 (N_28419,N_26952,N_26418);
and U28420 (N_28420,N_25933,N_25011);
and U28421 (N_28421,N_26273,N_25415);
xor U28422 (N_28422,N_25779,N_25128);
or U28423 (N_28423,N_27086,N_26108);
nand U28424 (N_28424,N_25185,N_26962);
nand U28425 (N_28425,N_25466,N_26237);
and U28426 (N_28426,N_27088,N_25439);
xor U28427 (N_28427,N_25347,N_27031);
or U28428 (N_28428,N_26140,N_25075);
nor U28429 (N_28429,N_25070,N_27029);
nand U28430 (N_28430,N_27238,N_25567);
nand U28431 (N_28431,N_26618,N_25204);
nor U28432 (N_28432,N_25325,N_26811);
nor U28433 (N_28433,N_27140,N_26769);
nor U28434 (N_28434,N_25840,N_25146);
and U28435 (N_28435,N_26387,N_25109);
nand U28436 (N_28436,N_26883,N_27460);
xnor U28437 (N_28437,N_26308,N_27466);
xor U28438 (N_28438,N_26109,N_26266);
nand U28439 (N_28439,N_27470,N_27223);
nor U28440 (N_28440,N_26386,N_26220);
or U28441 (N_28441,N_26935,N_25001);
or U28442 (N_28442,N_27008,N_26906);
or U28443 (N_28443,N_26740,N_27096);
or U28444 (N_28444,N_26501,N_26471);
or U28445 (N_28445,N_27399,N_27263);
or U28446 (N_28446,N_26860,N_25700);
xnor U28447 (N_28447,N_26765,N_25806);
nor U28448 (N_28448,N_25785,N_27331);
xor U28449 (N_28449,N_25365,N_26750);
nor U28450 (N_28450,N_27350,N_26620);
nand U28451 (N_28451,N_27160,N_26116);
nor U28452 (N_28452,N_27477,N_25455);
xnor U28453 (N_28453,N_25603,N_26403);
nand U28454 (N_28454,N_26842,N_27243);
nor U28455 (N_28455,N_26737,N_26318);
nor U28456 (N_28456,N_25273,N_26374);
xnor U28457 (N_28457,N_26465,N_26985);
and U28458 (N_28458,N_26516,N_26539);
and U28459 (N_28459,N_25184,N_25428);
or U28460 (N_28460,N_25078,N_25060);
nand U28461 (N_28461,N_25930,N_25727);
xnor U28462 (N_28462,N_27208,N_26728);
nand U28463 (N_28463,N_26098,N_25093);
nor U28464 (N_28464,N_26235,N_25768);
nand U28465 (N_28465,N_27201,N_26084);
xnor U28466 (N_28466,N_26169,N_26061);
or U28467 (N_28467,N_26316,N_27396);
nor U28468 (N_28468,N_25277,N_27379);
xor U28469 (N_28469,N_25790,N_27448);
or U28470 (N_28470,N_26805,N_25999);
nor U28471 (N_28471,N_27335,N_27046);
nor U28472 (N_28472,N_25960,N_26602);
xnor U28473 (N_28473,N_25437,N_25008);
or U28474 (N_28474,N_25695,N_27296);
nor U28475 (N_28475,N_26381,N_27499);
or U28476 (N_28476,N_26953,N_25523);
nor U28477 (N_28477,N_26476,N_25876);
and U28478 (N_28478,N_27040,N_25775);
and U28479 (N_28479,N_25874,N_25698);
nand U28480 (N_28480,N_26470,N_26677);
xor U28481 (N_28481,N_26912,N_25547);
nand U28482 (N_28482,N_27398,N_25864);
xnor U28483 (N_28483,N_26574,N_27228);
xnor U28484 (N_28484,N_27349,N_25536);
or U28485 (N_28485,N_26104,N_26615);
nor U28486 (N_28486,N_26376,N_26534);
nor U28487 (N_28487,N_26192,N_26796);
nor U28488 (N_28488,N_26895,N_26134);
nor U28489 (N_28489,N_25016,N_26543);
and U28490 (N_28490,N_25130,N_26514);
nand U28491 (N_28491,N_26293,N_26350);
and U28492 (N_28492,N_27219,N_25883);
xor U28493 (N_28493,N_26040,N_26137);
nor U28494 (N_28494,N_25579,N_25386);
and U28495 (N_28495,N_27423,N_26384);
nand U28496 (N_28496,N_25176,N_27226);
or U28497 (N_28497,N_25925,N_25436);
or U28498 (N_28498,N_26458,N_26924);
or U28499 (N_28499,N_26280,N_26969);
xnor U28500 (N_28500,N_25863,N_27050);
or U28501 (N_28501,N_27376,N_25973);
nand U28502 (N_28502,N_27433,N_27141);
nor U28503 (N_28503,N_25780,N_25300);
xnor U28504 (N_28504,N_26569,N_25575);
nand U28505 (N_28505,N_25205,N_27014);
and U28506 (N_28506,N_26956,N_26264);
nand U28507 (N_28507,N_25174,N_26738);
xnor U28508 (N_28508,N_25669,N_25334);
nor U28509 (N_28509,N_25272,N_26654);
nand U28510 (N_28510,N_25701,N_25878);
nor U28511 (N_28511,N_27222,N_26507);
nand U28512 (N_28512,N_26901,N_25711);
and U28513 (N_28513,N_27099,N_25242);
nor U28514 (N_28514,N_27422,N_26049);
and U28515 (N_28515,N_26085,N_26646);
or U28516 (N_28516,N_26367,N_26262);
nand U28517 (N_28517,N_27245,N_26823);
nor U28518 (N_28518,N_25920,N_26669);
xnor U28519 (N_28519,N_25477,N_25963);
and U28520 (N_28520,N_25713,N_26204);
nand U28521 (N_28521,N_27211,N_26607);
xnor U28522 (N_28522,N_25748,N_26641);
nand U28523 (N_28523,N_26044,N_26167);
nor U28524 (N_28524,N_25846,N_25211);
nand U28525 (N_28525,N_25393,N_27438);
xor U28526 (N_28526,N_26031,N_27274);
nor U28527 (N_28527,N_26375,N_26882);
nor U28528 (N_28528,N_25845,N_27416);
nand U28529 (N_28529,N_26132,N_26453);
and U28530 (N_28530,N_25144,N_25718);
nand U28531 (N_28531,N_26433,N_26290);
nor U28532 (N_28532,N_25929,N_25757);
and U28533 (N_28533,N_27230,N_26996);
xor U28534 (N_28534,N_26659,N_25841);
xor U28535 (N_28535,N_25937,N_27432);
nand U28536 (N_28536,N_25770,N_25366);
and U28537 (N_28537,N_25132,N_25626);
and U28538 (N_28538,N_25212,N_25830);
or U28539 (N_28539,N_27307,N_25553);
nor U28540 (N_28540,N_27091,N_25221);
or U28541 (N_28541,N_25309,N_26317);
nand U28542 (N_28542,N_26695,N_25959);
nor U28543 (N_28543,N_27071,N_27337);
nor U28544 (N_28544,N_25531,N_26125);
or U28545 (N_28545,N_25660,N_25044);
xor U28546 (N_28546,N_26522,N_26959);
and U28547 (N_28547,N_26997,N_25462);
and U28548 (N_28548,N_27498,N_26606);
nor U28549 (N_28549,N_26643,N_27455);
nand U28550 (N_28550,N_26932,N_27383);
nor U28551 (N_28551,N_27109,N_26900);
or U28552 (N_28552,N_25053,N_26302);
nand U28553 (N_28553,N_27152,N_26164);
and U28554 (N_28554,N_27380,N_26684);
and U28555 (N_28555,N_27117,N_25029);
nor U28556 (N_28556,N_25384,N_27013);
nor U28557 (N_28557,N_26777,N_25356);
and U28558 (N_28558,N_25417,N_25510);
nor U28559 (N_28559,N_26126,N_26429);
or U28560 (N_28560,N_25166,N_27492);
nand U28561 (N_28561,N_25871,N_25653);
xor U28562 (N_28562,N_27297,N_25274);
nor U28563 (N_28563,N_27122,N_26727);
nor U28564 (N_28564,N_26149,N_25087);
nand U28565 (N_28565,N_27473,N_25202);
or U28566 (N_28566,N_25024,N_25456);
nor U28567 (N_28567,N_26166,N_27494);
nand U28568 (N_28568,N_25917,N_26582);
nor U28569 (N_28569,N_25716,N_25495);
or U28570 (N_28570,N_25424,N_26019);
nand U28571 (N_28571,N_26552,N_27156);
or U28572 (N_28572,N_25350,N_26588);
xor U28573 (N_28573,N_25263,N_26773);
or U28574 (N_28574,N_25851,N_25376);
xnor U28575 (N_28575,N_26404,N_27421);
and U28576 (N_28576,N_26658,N_26976);
or U28577 (N_28577,N_26056,N_27240);
or U28578 (N_28578,N_27234,N_26397);
or U28579 (N_28579,N_26573,N_25962);
or U28580 (N_28580,N_25328,N_26069);
and U28581 (N_28581,N_26579,N_26153);
or U28582 (N_28582,N_25993,N_25057);
nand U28583 (N_28583,N_26181,N_26023);
or U28584 (N_28584,N_25367,N_26016);
and U28585 (N_28585,N_26026,N_26967);
or U28586 (N_28586,N_26563,N_26624);
and U28587 (N_28587,N_25326,N_25605);
nor U28588 (N_28588,N_26841,N_27371);
or U28589 (N_28589,N_27386,N_26802);
xor U28590 (N_28590,N_25749,N_26755);
nand U28591 (N_28591,N_25200,N_25451);
or U28592 (N_28592,N_25116,N_25682);
nor U28593 (N_28593,N_27389,N_25468);
nor U28594 (N_28594,N_27199,N_25870);
and U28595 (N_28595,N_27493,N_26861);
xnor U28596 (N_28596,N_25055,N_26904);
and U28597 (N_28597,N_26605,N_25298);
nand U28598 (N_28598,N_26444,N_26208);
nor U28599 (N_28599,N_25448,N_25381);
and U28600 (N_28600,N_27353,N_26183);
xnor U28601 (N_28601,N_26250,N_26561);
and U28602 (N_28602,N_27285,N_26447);
nand U28603 (N_28603,N_25065,N_25583);
and U28604 (N_28604,N_26495,N_26496);
nor U28605 (N_28605,N_25703,N_27280);
nor U28606 (N_28606,N_26243,N_27313);
nand U28607 (N_28607,N_26001,N_27434);
nand U28608 (N_28608,N_27094,N_27388);
xor U28609 (N_28609,N_27044,N_26503);
xor U28610 (N_28610,N_26392,N_25535);
xor U28611 (N_28611,N_26623,N_25600);
nand U28612 (N_28612,N_26911,N_25037);
nor U28613 (N_28613,N_26531,N_25900);
and U28614 (N_28614,N_26763,N_27185);
nand U28615 (N_28615,N_27427,N_25772);
xnor U28616 (N_28616,N_26537,N_27257);
and U28617 (N_28617,N_25961,N_26244);
nor U28618 (N_28618,N_27125,N_26712);
and U28619 (N_28619,N_27005,N_25502);
nand U28620 (N_28620,N_27397,N_25241);
nand U28621 (N_28621,N_26345,N_25760);
nand U28622 (N_28622,N_25773,N_26482);
nor U28623 (N_28623,N_27237,N_26441);
and U28624 (N_28624,N_27205,N_26062);
or U28625 (N_28625,N_25464,N_25299);
xor U28626 (N_28626,N_27429,N_26395);
xnor U28627 (N_28627,N_26914,N_27041);
and U28628 (N_28628,N_27412,N_25199);
or U28629 (N_28629,N_27176,N_26889);
xnor U28630 (N_28630,N_25294,N_25327);
nor U28631 (N_28631,N_25458,N_26022);
nor U28632 (N_28632,N_27131,N_26231);
nand U28633 (N_28633,N_27059,N_27077);
nand U28634 (N_28634,N_26508,N_26919);
xnor U28635 (N_28635,N_25173,N_27489);
xnor U28636 (N_28636,N_25323,N_25872);
or U28637 (N_28637,N_26357,N_27147);
nor U28638 (N_28638,N_26045,N_26694);
nand U28639 (N_28639,N_27294,N_25561);
xor U28640 (N_28640,N_25548,N_27406);
and U28641 (N_28641,N_25286,N_25618);
and U28642 (N_28642,N_27221,N_25997);
nand U28643 (N_28643,N_25496,N_25306);
or U28644 (N_28644,N_25837,N_25910);
xnor U28645 (N_28645,N_26928,N_26957);
nor U28646 (N_28646,N_27365,N_25167);
nor U28647 (N_28647,N_25302,N_26907);
or U28648 (N_28648,N_25885,N_26538);
or U28649 (N_28649,N_25104,N_26807);
and U28650 (N_28650,N_25432,N_25491);
xor U28651 (N_28651,N_26971,N_27367);
xor U28652 (N_28652,N_26571,N_25890);
nor U28653 (N_28653,N_26047,N_26053);
or U28654 (N_28654,N_26320,N_26018);
nand U28655 (N_28655,N_25207,N_25475);
xnor U28656 (N_28656,N_25914,N_26896);
nor U28657 (N_28657,N_25574,N_25320);
or U28658 (N_28658,N_26070,N_27461);
nand U28659 (N_28659,N_26525,N_25264);
nand U28660 (N_28660,N_25408,N_27151);
nand U28661 (N_28661,N_26774,N_25290);
nor U28662 (N_28662,N_25203,N_25884);
nor U28663 (N_28663,N_26355,N_25450);
nand U28664 (N_28664,N_27464,N_25506);
nor U28665 (N_28665,N_25734,N_26937);
and U28666 (N_28666,N_25344,N_25138);
nor U28667 (N_28667,N_26545,N_25654);
xnor U28668 (N_28668,N_26917,N_27231);
or U28669 (N_28669,N_26236,N_26747);
nand U28670 (N_28670,N_25988,N_25953);
or U28671 (N_28671,N_27214,N_25998);
nand U28672 (N_28672,N_26017,N_26072);
nand U28673 (N_28673,N_25767,N_25229);
xnor U28674 (N_28674,N_25541,N_26141);
nor U28675 (N_28675,N_25418,N_27292);
nand U28676 (N_28676,N_27024,N_25303);
xor U28677 (N_28677,N_26437,N_25270);
xor U28678 (N_28678,N_26162,N_27120);
xor U28679 (N_28679,N_26945,N_26764);
and U28680 (N_28680,N_25595,N_26370);
nor U28681 (N_28681,N_27326,N_25705);
nor U28682 (N_28682,N_25121,N_25453);
and U28683 (N_28683,N_26544,N_26670);
nor U28684 (N_28684,N_25441,N_26036);
or U28685 (N_28685,N_25818,N_25934);
nor U28686 (N_28686,N_26998,N_25395);
nor U28687 (N_28687,N_25854,N_25399);
and U28688 (N_28688,N_26535,N_26651);
xor U28689 (N_28689,N_26683,N_26975);
nand U28690 (N_28690,N_25363,N_26806);
nand U28691 (N_28691,N_25020,N_25296);
nor U28692 (N_28692,N_26299,N_27182);
nand U28693 (N_28693,N_26627,N_25474);
nor U28694 (N_28694,N_27483,N_25580);
xnor U28695 (N_28695,N_26296,N_25004);
or U28696 (N_28696,N_27042,N_27183);
xnor U28697 (N_28697,N_26637,N_26818);
or U28698 (N_28698,N_26438,N_26351);
and U28699 (N_28699,N_27076,N_25881);
and U28700 (N_28700,N_26993,N_25667);
nor U28701 (N_28701,N_25947,N_25662);
nor U28702 (N_28702,N_25064,N_25544);
and U28703 (N_28703,N_25155,N_25031);
or U28704 (N_28704,N_27232,N_26931);
xor U28705 (N_28705,N_26389,N_26717);
xor U28706 (N_28706,N_26687,N_26870);
and U28707 (N_28707,N_26129,N_26611);
and U28708 (N_28708,N_26087,N_25022);
or U28709 (N_28709,N_25360,N_26133);
nand U28710 (N_28710,N_26787,N_26464);
and U28711 (N_28711,N_25774,N_25223);
xor U28712 (N_28712,N_26341,N_25467);
nand U28713 (N_28713,N_26211,N_26041);
nand U28714 (N_28714,N_25118,N_25590);
nor U28715 (N_28715,N_26638,N_25717);
and U28716 (N_28716,N_26426,N_26248);
and U28717 (N_28717,N_25563,N_26492);
or U28718 (N_28718,N_26449,N_26515);
and U28719 (N_28719,N_25905,N_25861);
xor U28720 (N_28720,N_25844,N_26864);
xnor U28721 (N_28721,N_26285,N_27166);
or U28722 (N_28722,N_25511,N_26421);
or U28723 (N_28723,N_27364,N_26938);
nand U28724 (N_28724,N_27395,N_26995);
or U28725 (N_28725,N_26232,N_25162);
nor U28726 (N_28726,N_25007,N_25452);
nor U28727 (N_28727,N_25372,N_26718);
nand U28728 (N_28728,N_26692,N_25783);
or U28729 (N_28729,N_26671,N_26549);
nand U28730 (N_28730,N_26057,N_26751);
and U28731 (N_28731,N_25067,N_25297);
nor U28732 (N_28732,N_26113,N_25319);
or U28733 (N_28733,N_25584,N_25926);
nor U28734 (N_28734,N_26562,N_25939);
and U28735 (N_28735,N_25889,N_27073);
or U28736 (N_28736,N_26653,N_25586);
nand U28737 (N_28737,N_27355,N_26855);
or U28738 (N_28738,N_26325,N_25295);
nor U28739 (N_28739,N_26994,N_27068);
or U28740 (N_28740,N_25940,N_26234);
xor U28741 (N_28741,N_25407,N_26336);
and U28742 (N_28742,N_25640,N_26828);
xnor U28743 (N_28743,N_26128,N_26639);
nand U28744 (N_28744,N_25816,N_26463);
and U28745 (N_28745,N_25637,N_26050);
nand U28746 (N_28746,N_26154,N_25802);
and U28747 (N_28747,N_25021,N_27366);
nor U28748 (N_28748,N_27133,N_27057);
xnor U28749 (N_28749,N_27225,N_27022);
xnor U28750 (N_28750,N_26354,N_25840);
nand U28751 (N_28751,N_25834,N_26316);
and U28752 (N_28752,N_26314,N_25766);
or U28753 (N_28753,N_26083,N_26597);
and U28754 (N_28754,N_25000,N_26042);
nor U28755 (N_28755,N_25740,N_26995);
nor U28756 (N_28756,N_27453,N_26273);
and U28757 (N_28757,N_25197,N_25776);
nand U28758 (N_28758,N_26817,N_27494);
and U28759 (N_28759,N_26429,N_25201);
nor U28760 (N_28760,N_26129,N_27043);
or U28761 (N_28761,N_27174,N_26853);
xnor U28762 (N_28762,N_25018,N_25586);
and U28763 (N_28763,N_27421,N_25904);
and U28764 (N_28764,N_26963,N_27354);
nand U28765 (N_28765,N_26764,N_26729);
nor U28766 (N_28766,N_26837,N_25515);
xor U28767 (N_28767,N_26572,N_26756);
nor U28768 (N_28768,N_26350,N_27385);
nand U28769 (N_28769,N_26042,N_26653);
or U28770 (N_28770,N_25613,N_26842);
nor U28771 (N_28771,N_25235,N_25872);
nand U28772 (N_28772,N_25280,N_26649);
nor U28773 (N_28773,N_25453,N_25310);
and U28774 (N_28774,N_27457,N_25108);
xnor U28775 (N_28775,N_26263,N_25076);
nand U28776 (N_28776,N_25521,N_26034);
or U28777 (N_28777,N_27091,N_26060);
and U28778 (N_28778,N_26673,N_25064);
or U28779 (N_28779,N_25816,N_25219);
nor U28780 (N_28780,N_26127,N_25004);
nand U28781 (N_28781,N_25796,N_26753);
nor U28782 (N_28782,N_26614,N_27260);
or U28783 (N_28783,N_25927,N_26267);
xnor U28784 (N_28784,N_26019,N_27165);
nor U28785 (N_28785,N_25639,N_25312);
nand U28786 (N_28786,N_26155,N_25893);
nor U28787 (N_28787,N_26434,N_25749);
and U28788 (N_28788,N_25450,N_26382);
or U28789 (N_28789,N_26774,N_26239);
nand U28790 (N_28790,N_26042,N_25471);
nor U28791 (N_28791,N_26733,N_27034);
nor U28792 (N_28792,N_27001,N_25190);
or U28793 (N_28793,N_25132,N_26347);
and U28794 (N_28794,N_25090,N_27176);
or U28795 (N_28795,N_25529,N_25229);
nor U28796 (N_28796,N_26646,N_25537);
or U28797 (N_28797,N_27163,N_25175);
nor U28798 (N_28798,N_26786,N_25848);
nand U28799 (N_28799,N_26070,N_26482);
and U28800 (N_28800,N_25342,N_27074);
nor U28801 (N_28801,N_27219,N_26852);
nor U28802 (N_28802,N_26654,N_26755);
xor U28803 (N_28803,N_25992,N_26286);
or U28804 (N_28804,N_26392,N_26631);
and U28805 (N_28805,N_26064,N_25782);
or U28806 (N_28806,N_26424,N_27419);
xnor U28807 (N_28807,N_25690,N_25295);
xor U28808 (N_28808,N_26397,N_25232);
or U28809 (N_28809,N_26995,N_25490);
xnor U28810 (N_28810,N_25418,N_26125);
xor U28811 (N_28811,N_26365,N_26317);
and U28812 (N_28812,N_27208,N_26295);
or U28813 (N_28813,N_26041,N_25709);
nand U28814 (N_28814,N_26678,N_25570);
nand U28815 (N_28815,N_25702,N_25556);
nand U28816 (N_28816,N_26989,N_25257);
xor U28817 (N_28817,N_26134,N_26462);
or U28818 (N_28818,N_26981,N_26071);
nor U28819 (N_28819,N_26115,N_27319);
or U28820 (N_28820,N_27398,N_27059);
or U28821 (N_28821,N_25995,N_25139);
nor U28822 (N_28822,N_25067,N_27404);
xor U28823 (N_28823,N_25927,N_26973);
nor U28824 (N_28824,N_27418,N_26092);
or U28825 (N_28825,N_26143,N_26464);
xor U28826 (N_28826,N_25724,N_25831);
nand U28827 (N_28827,N_27269,N_25731);
nand U28828 (N_28828,N_25475,N_27325);
and U28829 (N_28829,N_26564,N_27048);
nor U28830 (N_28830,N_26433,N_25653);
and U28831 (N_28831,N_27143,N_26018);
and U28832 (N_28832,N_26301,N_25398);
nor U28833 (N_28833,N_25776,N_26619);
or U28834 (N_28834,N_26440,N_25374);
nand U28835 (N_28835,N_25671,N_25862);
nand U28836 (N_28836,N_26177,N_25692);
nor U28837 (N_28837,N_26736,N_25123);
nand U28838 (N_28838,N_26796,N_26887);
nand U28839 (N_28839,N_25212,N_26623);
nor U28840 (N_28840,N_25286,N_27377);
nor U28841 (N_28841,N_26199,N_25804);
xor U28842 (N_28842,N_27054,N_27446);
nor U28843 (N_28843,N_26345,N_25820);
xor U28844 (N_28844,N_26895,N_25903);
nand U28845 (N_28845,N_25755,N_25924);
or U28846 (N_28846,N_25983,N_26040);
nand U28847 (N_28847,N_26019,N_26458);
or U28848 (N_28848,N_26198,N_27283);
nand U28849 (N_28849,N_26664,N_26460);
or U28850 (N_28850,N_26183,N_26968);
and U28851 (N_28851,N_27085,N_25762);
and U28852 (N_28852,N_26483,N_25679);
or U28853 (N_28853,N_26559,N_26224);
xor U28854 (N_28854,N_26767,N_25919);
xor U28855 (N_28855,N_25581,N_27053);
nand U28856 (N_28856,N_25473,N_25608);
or U28857 (N_28857,N_26410,N_25188);
xor U28858 (N_28858,N_25006,N_26962);
and U28859 (N_28859,N_26825,N_26045);
or U28860 (N_28860,N_26884,N_26932);
and U28861 (N_28861,N_25654,N_25396);
and U28862 (N_28862,N_25851,N_25951);
xnor U28863 (N_28863,N_26153,N_26897);
nor U28864 (N_28864,N_25157,N_27416);
and U28865 (N_28865,N_26580,N_25657);
nand U28866 (N_28866,N_26028,N_27182);
and U28867 (N_28867,N_25826,N_26123);
or U28868 (N_28868,N_26852,N_26295);
nand U28869 (N_28869,N_25585,N_26898);
xnor U28870 (N_28870,N_25007,N_25857);
or U28871 (N_28871,N_27020,N_25991);
nor U28872 (N_28872,N_25748,N_26159);
nand U28873 (N_28873,N_25487,N_25439);
nor U28874 (N_28874,N_26424,N_26602);
nor U28875 (N_28875,N_26773,N_26117);
xnor U28876 (N_28876,N_25767,N_27239);
xor U28877 (N_28877,N_25374,N_25742);
xor U28878 (N_28878,N_26569,N_25396);
nor U28879 (N_28879,N_27404,N_26041);
xor U28880 (N_28880,N_27163,N_25587);
or U28881 (N_28881,N_25721,N_25478);
and U28882 (N_28882,N_26945,N_25785);
xor U28883 (N_28883,N_27301,N_25514);
and U28884 (N_28884,N_26228,N_25118);
nand U28885 (N_28885,N_26284,N_25094);
nor U28886 (N_28886,N_26296,N_27130);
nor U28887 (N_28887,N_26844,N_25686);
nand U28888 (N_28888,N_27344,N_26062);
or U28889 (N_28889,N_27399,N_25722);
or U28890 (N_28890,N_25045,N_25604);
and U28891 (N_28891,N_27049,N_26526);
nand U28892 (N_28892,N_26709,N_26016);
nor U28893 (N_28893,N_26871,N_25276);
nor U28894 (N_28894,N_26697,N_25800);
nor U28895 (N_28895,N_25195,N_27149);
nand U28896 (N_28896,N_25808,N_26009);
and U28897 (N_28897,N_26358,N_27379);
nor U28898 (N_28898,N_26461,N_27429);
or U28899 (N_28899,N_26935,N_25407);
xnor U28900 (N_28900,N_26782,N_26897);
and U28901 (N_28901,N_26739,N_26463);
nand U28902 (N_28902,N_26059,N_25067);
xnor U28903 (N_28903,N_26553,N_25068);
nor U28904 (N_28904,N_27280,N_25982);
and U28905 (N_28905,N_27100,N_25063);
nor U28906 (N_28906,N_27325,N_27032);
nand U28907 (N_28907,N_26908,N_26801);
xor U28908 (N_28908,N_27270,N_25317);
nor U28909 (N_28909,N_27309,N_26368);
or U28910 (N_28910,N_26618,N_25515);
or U28911 (N_28911,N_26129,N_26619);
xor U28912 (N_28912,N_25147,N_26529);
or U28913 (N_28913,N_26532,N_26461);
xnor U28914 (N_28914,N_26476,N_26712);
and U28915 (N_28915,N_27206,N_26897);
nand U28916 (N_28916,N_25517,N_27185);
or U28917 (N_28917,N_26582,N_25226);
nor U28918 (N_28918,N_26937,N_25422);
or U28919 (N_28919,N_26533,N_27319);
xor U28920 (N_28920,N_26115,N_26991);
xor U28921 (N_28921,N_25304,N_26891);
nand U28922 (N_28922,N_26097,N_26093);
or U28923 (N_28923,N_26633,N_26397);
nand U28924 (N_28924,N_27146,N_27385);
or U28925 (N_28925,N_26060,N_27200);
nor U28926 (N_28926,N_27050,N_26386);
xor U28927 (N_28927,N_25307,N_26851);
nand U28928 (N_28928,N_25085,N_26630);
and U28929 (N_28929,N_26671,N_26112);
and U28930 (N_28930,N_27214,N_27050);
nor U28931 (N_28931,N_25910,N_26311);
xnor U28932 (N_28932,N_27151,N_26766);
xor U28933 (N_28933,N_27453,N_26723);
nand U28934 (N_28934,N_25192,N_25630);
and U28935 (N_28935,N_27110,N_25063);
or U28936 (N_28936,N_25239,N_26985);
or U28937 (N_28937,N_25807,N_25268);
or U28938 (N_28938,N_26705,N_26784);
xor U28939 (N_28939,N_26739,N_26716);
or U28940 (N_28940,N_25958,N_25781);
or U28941 (N_28941,N_26676,N_25315);
or U28942 (N_28942,N_25110,N_26275);
nand U28943 (N_28943,N_25018,N_26843);
or U28944 (N_28944,N_25126,N_25657);
xor U28945 (N_28945,N_25812,N_27086);
xor U28946 (N_28946,N_26295,N_27227);
xor U28947 (N_28947,N_25995,N_26229);
and U28948 (N_28948,N_26771,N_25286);
or U28949 (N_28949,N_25196,N_25737);
nand U28950 (N_28950,N_26831,N_26675);
nor U28951 (N_28951,N_25681,N_25790);
xor U28952 (N_28952,N_25672,N_26162);
or U28953 (N_28953,N_27479,N_25571);
xor U28954 (N_28954,N_26895,N_25357);
or U28955 (N_28955,N_27162,N_25743);
and U28956 (N_28956,N_25900,N_25240);
or U28957 (N_28957,N_26235,N_27318);
nor U28958 (N_28958,N_25333,N_26676);
nand U28959 (N_28959,N_27119,N_26008);
xor U28960 (N_28960,N_26520,N_25925);
nor U28961 (N_28961,N_27018,N_27460);
and U28962 (N_28962,N_25102,N_26351);
and U28963 (N_28963,N_27343,N_25269);
and U28964 (N_28964,N_26470,N_26632);
nor U28965 (N_28965,N_26121,N_25446);
and U28966 (N_28966,N_27077,N_25496);
or U28967 (N_28967,N_25918,N_26427);
xnor U28968 (N_28968,N_25247,N_25127);
or U28969 (N_28969,N_25196,N_27209);
nor U28970 (N_28970,N_27436,N_26970);
or U28971 (N_28971,N_25162,N_25988);
and U28972 (N_28972,N_26546,N_26461);
or U28973 (N_28973,N_26903,N_26410);
nand U28974 (N_28974,N_25564,N_26689);
nor U28975 (N_28975,N_25347,N_25982);
xnor U28976 (N_28976,N_26461,N_26055);
and U28977 (N_28977,N_25258,N_26064);
xor U28978 (N_28978,N_26623,N_25779);
and U28979 (N_28979,N_26439,N_25391);
xor U28980 (N_28980,N_27417,N_25204);
xnor U28981 (N_28981,N_26393,N_26186);
nor U28982 (N_28982,N_25045,N_25968);
nand U28983 (N_28983,N_25193,N_26782);
xor U28984 (N_28984,N_26803,N_27246);
xor U28985 (N_28985,N_25188,N_26738);
xnor U28986 (N_28986,N_26442,N_25853);
nor U28987 (N_28987,N_25646,N_26407);
or U28988 (N_28988,N_26464,N_26564);
nand U28989 (N_28989,N_27166,N_26603);
or U28990 (N_28990,N_25536,N_26572);
nand U28991 (N_28991,N_25986,N_26964);
and U28992 (N_28992,N_27184,N_27337);
and U28993 (N_28993,N_26248,N_25362);
and U28994 (N_28994,N_26541,N_26936);
and U28995 (N_28995,N_26998,N_26667);
nand U28996 (N_28996,N_25607,N_26777);
nor U28997 (N_28997,N_27402,N_25825);
and U28998 (N_28998,N_25213,N_25315);
nand U28999 (N_28999,N_27460,N_26143);
xor U29000 (N_29000,N_27481,N_26842);
or U29001 (N_29001,N_27125,N_27473);
or U29002 (N_29002,N_26531,N_26122);
nor U29003 (N_29003,N_25359,N_26188);
nor U29004 (N_29004,N_26931,N_25730);
and U29005 (N_29005,N_26082,N_26552);
nor U29006 (N_29006,N_26409,N_27250);
or U29007 (N_29007,N_26996,N_25076);
xnor U29008 (N_29008,N_25991,N_27241);
or U29009 (N_29009,N_25396,N_26450);
nor U29010 (N_29010,N_26655,N_26415);
and U29011 (N_29011,N_26162,N_25660);
xnor U29012 (N_29012,N_26681,N_25224);
nor U29013 (N_29013,N_26079,N_27077);
nand U29014 (N_29014,N_26350,N_27232);
nor U29015 (N_29015,N_25833,N_26724);
and U29016 (N_29016,N_27150,N_25762);
and U29017 (N_29017,N_26017,N_25246);
and U29018 (N_29018,N_25693,N_26294);
or U29019 (N_29019,N_25933,N_25724);
or U29020 (N_29020,N_26909,N_26959);
xnor U29021 (N_29021,N_26616,N_25423);
or U29022 (N_29022,N_25394,N_26223);
or U29023 (N_29023,N_26320,N_25706);
nor U29024 (N_29024,N_25535,N_25176);
and U29025 (N_29025,N_27420,N_27314);
or U29026 (N_29026,N_26734,N_27424);
and U29027 (N_29027,N_25064,N_25698);
and U29028 (N_29028,N_26275,N_25133);
nand U29029 (N_29029,N_27133,N_25167);
or U29030 (N_29030,N_25311,N_26604);
xnor U29031 (N_29031,N_26355,N_26369);
and U29032 (N_29032,N_25958,N_25773);
or U29033 (N_29033,N_26195,N_27150);
or U29034 (N_29034,N_25257,N_25144);
nand U29035 (N_29035,N_27003,N_25209);
and U29036 (N_29036,N_25446,N_25978);
nand U29037 (N_29037,N_25970,N_25365);
or U29038 (N_29038,N_25433,N_27282);
and U29039 (N_29039,N_27158,N_26096);
or U29040 (N_29040,N_25140,N_25151);
nand U29041 (N_29041,N_27050,N_26414);
or U29042 (N_29042,N_25794,N_25825);
or U29043 (N_29043,N_27062,N_26406);
and U29044 (N_29044,N_25737,N_27039);
nor U29045 (N_29045,N_25992,N_26231);
or U29046 (N_29046,N_26155,N_26448);
and U29047 (N_29047,N_25593,N_26944);
nor U29048 (N_29048,N_25155,N_27320);
and U29049 (N_29049,N_26954,N_25939);
xnor U29050 (N_29050,N_26524,N_27345);
xor U29051 (N_29051,N_25964,N_26190);
and U29052 (N_29052,N_25703,N_26937);
nor U29053 (N_29053,N_27243,N_25210);
nor U29054 (N_29054,N_26866,N_27209);
nand U29055 (N_29055,N_25350,N_25151);
and U29056 (N_29056,N_26717,N_26321);
or U29057 (N_29057,N_27470,N_26252);
or U29058 (N_29058,N_25973,N_26872);
xnor U29059 (N_29059,N_25950,N_26159);
xor U29060 (N_29060,N_26195,N_27220);
nand U29061 (N_29061,N_25061,N_26178);
xor U29062 (N_29062,N_26051,N_26189);
or U29063 (N_29063,N_25122,N_25700);
nor U29064 (N_29064,N_25038,N_27157);
xnor U29065 (N_29065,N_27259,N_26751);
and U29066 (N_29066,N_27247,N_25912);
nand U29067 (N_29067,N_25711,N_25394);
nor U29068 (N_29068,N_26744,N_26266);
nand U29069 (N_29069,N_25578,N_27233);
and U29070 (N_29070,N_25318,N_25463);
nand U29071 (N_29071,N_26270,N_26894);
nand U29072 (N_29072,N_25557,N_25564);
nor U29073 (N_29073,N_26943,N_26004);
or U29074 (N_29074,N_25498,N_26786);
or U29075 (N_29075,N_26631,N_27247);
xnor U29076 (N_29076,N_27482,N_26399);
nand U29077 (N_29077,N_25944,N_25613);
nand U29078 (N_29078,N_27298,N_26999);
nor U29079 (N_29079,N_25318,N_26740);
nand U29080 (N_29080,N_26505,N_26465);
nor U29081 (N_29081,N_25669,N_27137);
and U29082 (N_29082,N_25484,N_25653);
xnor U29083 (N_29083,N_25747,N_25154);
nand U29084 (N_29084,N_27377,N_26505);
and U29085 (N_29085,N_26349,N_26860);
and U29086 (N_29086,N_25416,N_25841);
nor U29087 (N_29087,N_25547,N_26817);
nand U29088 (N_29088,N_26012,N_27405);
and U29089 (N_29089,N_26720,N_26578);
nand U29090 (N_29090,N_26623,N_27175);
and U29091 (N_29091,N_25844,N_25561);
nand U29092 (N_29092,N_26090,N_26636);
nor U29093 (N_29093,N_26988,N_25884);
or U29094 (N_29094,N_26587,N_25460);
nand U29095 (N_29095,N_26942,N_26377);
and U29096 (N_29096,N_26503,N_26284);
and U29097 (N_29097,N_25666,N_26664);
or U29098 (N_29098,N_25884,N_25322);
xnor U29099 (N_29099,N_25655,N_25875);
and U29100 (N_29100,N_25274,N_25023);
or U29101 (N_29101,N_25266,N_26351);
and U29102 (N_29102,N_27235,N_25101);
nor U29103 (N_29103,N_25973,N_27284);
and U29104 (N_29104,N_26292,N_26352);
or U29105 (N_29105,N_25436,N_25420);
nor U29106 (N_29106,N_26014,N_26128);
and U29107 (N_29107,N_25020,N_26103);
nor U29108 (N_29108,N_26389,N_26913);
nand U29109 (N_29109,N_26154,N_25636);
nor U29110 (N_29110,N_25360,N_25790);
nand U29111 (N_29111,N_25628,N_26729);
nand U29112 (N_29112,N_25193,N_25244);
nor U29113 (N_29113,N_25369,N_25499);
nand U29114 (N_29114,N_27013,N_25541);
nor U29115 (N_29115,N_25240,N_27353);
and U29116 (N_29116,N_26073,N_26943);
nor U29117 (N_29117,N_27425,N_26590);
nor U29118 (N_29118,N_27366,N_26404);
nand U29119 (N_29119,N_25074,N_26184);
nand U29120 (N_29120,N_26584,N_26644);
and U29121 (N_29121,N_26304,N_26501);
or U29122 (N_29122,N_26038,N_25024);
nand U29123 (N_29123,N_26499,N_25468);
nor U29124 (N_29124,N_26715,N_25449);
nand U29125 (N_29125,N_26334,N_25113);
nand U29126 (N_29126,N_26221,N_26874);
and U29127 (N_29127,N_25317,N_26280);
nand U29128 (N_29128,N_26095,N_26116);
nor U29129 (N_29129,N_26458,N_27085);
and U29130 (N_29130,N_26722,N_25294);
or U29131 (N_29131,N_26309,N_25142);
and U29132 (N_29132,N_27039,N_25741);
xnor U29133 (N_29133,N_26972,N_26193);
and U29134 (N_29134,N_27047,N_27241);
or U29135 (N_29135,N_25405,N_25622);
or U29136 (N_29136,N_26342,N_25925);
nor U29137 (N_29137,N_25896,N_26864);
xnor U29138 (N_29138,N_26164,N_25742);
or U29139 (N_29139,N_25036,N_26211);
and U29140 (N_29140,N_26305,N_26302);
or U29141 (N_29141,N_26665,N_25333);
nand U29142 (N_29142,N_25234,N_27391);
nor U29143 (N_29143,N_26213,N_26900);
or U29144 (N_29144,N_27152,N_26898);
or U29145 (N_29145,N_25862,N_25469);
nor U29146 (N_29146,N_26875,N_25773);
xor U29147 (N_29147,N_27376,N_26181);
and U29148 (N_29148,N_25224,N_26725);
and U29149 (N_29149,N_25594,N_25372);
or U29150 (N_29150,N_26371,N_26202);
nor U29151 (N_29151,N_26928,N_26846);
or U29152 (N_29152,N_26910,N_26666);
xor U29153 (N_29153,N_25532,N_27034);
and U29154 (N_29154,N_26040,N_25736);
xnor U29155 (N_29155,N_26717,N_26401);
and U29156 (N_29156,N_25713,N_27399);
xnor U29157 (N_29157,N_25684,N_25727);
nand U29158 (N_29158,N_26547,N_26927);
and U29159 (N_29159,N_25458,N_26024);
xor U29160 (N_29160,N_25860,N_27052);
and U29161 (N_29161,N_27116,N_26925);
or U29162 (N_29162,N_25501,N_26815);
nor U29163 (N_29163,N_26130,N_27451);
nand U29164 (N_29164,N_25215,N_26800);
or U29165 (N_29165,N_25865,N_26638);
or U29166 (N_29166,N_26737,N_26806);
nor U29167 (N_29167,N_25486,N_25980);
and U29168 (N_29168,N_25223,N_25504);
xor U29169 (N_29169,N_25852,N_27331);
and U29170 (N_29170,N_26250,N_26010);
nand U29171 (N_29171,N_25329,N_26851);
or U29172 (N_29172,N_25520,N_26830);
xnor U29173 (N_29173,N_25959,N_25643);
and U29174 (N_29174,N_25459,N_25268);
xnor U29175 (N_29175,N_25591,N_27263);
and U29176 (N_29176,N_26527,N_25515);
and U29177 (N_29177,N_25700,N_26815);
xnor U29178 (N_29178,N_26041,N_27067);
or U29179 (N_29179,N_25455,N_26843);
nand U29180 (N_29180,N_25151,N_25489);
or U29181 (N_29181,N_26408,N_25978);
nor U29182 (N_29182,N_26187,N_27028);
or U29183 (N_29183,N_26756,N_26713);
and U29184 (N_29184,N_25147,N_25343);
nand U29185 (N_29185,N_27113,N_25742);
and U29186 (N_29186,N_26674,N_25004);
nor U29187 (N_29187,N_26764,N_25642);
or U29188 (N_29188,N_27360,N_27292);
and U29189 (N_29189,N_25634,N_25519);
or U29190 (N_29190,N_25033,N_26796);
nand U29191 (N_29191,N_27173,N_26239);
or U29192 (N_29192,N_25563,N_26864);
nor U29193 (N_29193,N_27330,N_26552);
or U29194 (N_29194,N_27370,N_25547);
xnor U29195 (N_29195,N_27379,N_26947);
and U29196 (N_29196,N_25134,N_25394);
xnor U29197 (N_29197,N_25463,N_25620);
nand U29198 (N_29198,N_25821,N_27113);
xnor U29199 (N_29199,N_26176,N_26202);
nor U29200 (N_29200,N_26939,N_26440);
nand U29201 (N_29201,N_27412,N_26137);
and U29202 (N_29202,N_26516,N_25188);
nand U29203 (N_29203,N_26627,N_25071);
or U29204 (N_29204,N_25519,N_27230);
nand U29205 (N_29205,N_27258,N_26079);
nor U29206 (N_29206,N_25770,N_27455);
and U29207 (N_29207,N_25283,N_25909);
nor U29208 (N_29208,N_26281,N_26770);
and U29209 (N_29209,N_26039,N_27471);
xor U29210 (N_29210,N_25417,N_27443);
nor U29211 (N_29211,N_25757,N_26475);
nor U29212 (N_29212,N_25654,N_26892);
xor U29213 (N_29213,N_25859,N_26792);
or U29214 (N_29214,N_25653,N_27497);
nor U29215 (N_29215,N_27374,N_25742);
nor U29216 (N_29216,N_27153,N_26900);
nor U29217 (N_29217,N_25670,N_25306);
and U29218 (N_29218,N_25412,N_26968);
or U29219 (N_29219,N_26635,N_26664);
xnor U29220 (N_29220,N_26613,N_26041);
and U29221 (N_29221,N_26063,N_26737);
nor U29222 (N_29222,N_27057,N_27402);
or U29223 (N_29223,N_26941,N_25885);
or U29224 (N_29224,N_25458,N_26030);
or U29225 (N_29225,N_26408,N_25187);
nor U29226 (N_29226,N_25552,N_25470);
xnor U29227 (N_29227,N_26598,N_26484);
nand U29228 (N_29228,N_25821,N_26249);
xor U29229 (N_29229,N_26417,N_26326);
or U29230 (N_29230,N_25725,N_25127);
nand U29231 (N_29231,N_26567,N_26721);
nor U29232 (N_29232,N_25751,N_26354);
and U29233 (N_29233,N_26440,N_26818);
nor U29234 (N_29234,N_25573,N_26179);
nor U29235 (N_29235,N_27080,N_26374);
or U29236 (N_29236,N_25208,N_25656);
nand U29237 (N_29237,N_25200,N_26061);
and U29238 (N_29238,N_27373,N_27071);
nor U29239 (N_29239,N_25976,N_25137);
and U29240 (N_29240,N_25802,N_25307);
and U29241 (N_29241,N_25617,N_26867);
nand U29242 (N_29242,N_27078,N_25924);
xnor U29243 (N_29243,N_26669,N_26281);
nand U29244 (N_29244,N_25088,N_27479);
nand U29245 (N_29245,N_27316,N_25788);
xor U29246 (N_29246,N_25234,N_25265);
or U29247 (N_29247,N_25689,N_27439);
nand U29248 (N_29248,N_26405,N_25507);
xor U29249 (N_29249,N_26966,N_25892);
nand U29250 (N_29250,N_25143,N_25781);
xor U29251 (N_29251,N_27307,N_25236);
nand U29252 (N_29252,N_25915,N_25168);
or U29253 (N_29253,N_27055,N_26356);
xor U29254 (N_29254,N_25498,N_26385);
and U29255 (N_29255,N_25169,N_27088);
or U29256 (N_29256,N_26033,N_26751);
xnor U29257 (N_29257,N_26274,N_27332);
xor U29258 (N_29258,N_25215,N_25105);
and U29259 (N_29259,N_25463,N_25526);
xor U29260 (N_29260,N_26554,N_26743);
nor U29261 (N_29261,N_25199,N_26530);
or U29262 (N_29262,N_26039,N_26550);
and U29263 (N_29263,N_25284,N_26515);
or U29264 (N_29264,N_25714,N_27383);
and U29265 (N_29265,N_25156,N_25411);
xnor U29266 (N_29266,N_26760,N_25287);
nand U29267 (N_29267,N_25179,N_25246);
nor U29268 (N_29268,N_26217,N_27423);
nor U29269 (N_29269,N_25441,N_27167);
nor U29270 (N_29270,N_25477,N_25991);
nor U29271 (N_29271,N_26769,N_25934);
nor U29272 (N_29272,N_26584,N_26539);
nand U29273 (N_29273,N_26269,N_26406);
nor U29274 (N_29274,N_26464,N_26011);
and U29275 (N_29275,N_26090,N_26784);
xnor U29276 (N_29276,N_26523,N_27057);
nor U29277 (N_29277,N_26980,N_26985);
nor U29278 (N_29278,N_25972,N_26283);
xor U29279 (N_29279,N_26011,N_26045);
or U29280 (N_29280,N_25738,N_25949);
nor U29281 (N_29281,N_26869,N_26886);
nor U29282 (N_29282,N_26024,N_27091);
nor U29283 (N_29283,N_27392,N_26577);
or U29284 (N_29284,N_25693,N_27304);
xor U29285 (N_29285,N_25341,N_27466);
or U29286 (N_29286,N_25563,N_26971);
nor U29287 (N_29287,N_27239,N_27154);
nand U29288 (N_29288,N_26343,N_27081);
xor U29289 (N_29289,N_26399,N_26208);
and U29290 (N_29290,N_26745,N_26833);
nand U29291 (N_29291,N_25070,N_26935);
or U29292 (N_29292,N_25852,N_27438);
xnor U29293 (N_29293,N_25098,N_26281);
xnor U29294 (N_29294,N_27252,N_25271);
and U29295 (N_29295,N_27091,N_26578);
and U29296 (N_29296,N_26229,N_27120);
xnor U29297 (N_29297,N_25043,N_26141);
nor U29298 (N_29298,N_25005,N_27171);
xnor U29299 (N_29299,N_26572,N_26407);
xor U29300 (N_29300,N_26044,N_26568);
and U29301 (N_29301,N_26765,N_26835);
nor U29302 (N_29302,N_25673,N_26490);
nor U29303 (N_29303,N_26605,N_26494);
nand U29304 (N_29304,N_26131,N_27455);
xor U29305 (N_29305,N_25092,N_25782);
nand U29306 (N_29306,N_27460,N_26272);
nand U29307 (N_29307,N_26347,N_26170);
xor U29308 (N_29308,N_26594,N_27284);
nand U29309 (N_29309,N_25728,N_26590);
nor U29310 (N_29310,N_26695,N_25376);
and U29311 (N_29311,N_25727,N_26376);
or U29312 (N_29312,N_26079,N_26044);
and U29313 (N_29313,N_27338,N_27058);
or U29314 (N_29314,N_26801,N_26516);
nand U29315 (N_29315,N_25460,N_27202);
nor U29316 (N_29316,N_25602,N_27251);
xnor U29317 (N_29317,N_25819,N_27271);
and U29318 (N_29318,N_27295,N_25609);
nor U29319 (N_29319,N_25870,N_27473);
xor U29320 (N_29320,N_26870,N_26024);
nor U29321 (N_29321,N_25101,N_27294);
or U29322 (N_29322,N_25271,N_27015);
and U29323 (N_29323,N_27435,N_26177);
or U29324 (N_29324,N_25982,N_25411);
nand U29325 (N_29325,N_25838,N_27253);
nand U29326 (N_29326,N_25160,N_25375);
nor U29327 (N_29327,N_27128,N_25760);
and U29328 (N_29328,N_25813,N_25605);
nor U29329 (N_29329,N_26312,N_25761);
or U29330 (N_29330,N_25474,N_26120);
and U29331 (N_29331,N_26783,N_26928);
or U29332 (N_29332,N_25994,N_27258);
and U29333 (N_29333,N_26548,N_25319);
xnor U29334 (N_29334,N_26909,N_25399);
and U29335 (N_29335,N_25684,N_25130);
nor U29336 (N_29336,N_26102,N_26152);
or U29337 (N_29337,N_26527,N_25780);
and U29338 (N_29338,N_26904,N_26774);
xnor U29339 (N_29339,N_26439,N_26809);
and U29340 (N_29340,N_26376,N_25988);
and U29341 (N_29341,N_25736,N_27135);
nor U29342 (N_29342,N_27372,N_25803);
xor U29343 (N_29343,N_25117,N_26133);
xnor U29344 (N_29344,N_27178,N_27129);
xor U29345 (N_29345,N_27249,N_25175);
or U29346 (N_29346,N_26400,N_26893);
or U29347 (N_29347,N_27491,N_26709);
nor U29348 (N_29348,N_27037,N_27076);
and U29349 (N_29349,N_26633,N_25041);
nor U29350 (N_29350,N_25631,N_26724);
xor U29351 (N_29351,N_25262,N_25665);
and U29352 (N_29352,N_26812,N_25154);
nor U29353 (N_29353,N_26988,N_26875);
and U29354 (N_29354,N_26501,N_26756);
or U29355 (N_29355,N_26065,N_25708);
xor U29356 (N_29356,N_27140,N_26432);
xnor U29357 (N_29357,N_26976,N_25260);
nand U29358 (N_29358,N_25898,N_26404);
and U29359 (N_29359,N_25527,N_26330);
xor U29360 (N_29360,N_25790,N_26957);
nor U29361 (N_29361,N_27470,N_27198);
and U29362 (N_29362,N_26019,N_25814);
and U29363 (N_29363,N_26937,N_26855);
nand U29364 (N_29364,N_25728,N_26770);
nand U29365 (N_29365,N_26499,N_26695);
nand U29366 (N_29366,N_25457,N_25992);
or U29367 (N_29367,N_26473,N_26001);
xnor U29368 (N_29368,N_25470,N_27404);
nor U29369 (N_29369,N_26049,N_27308);
and U29370 (N_29370,N_26311,N_27222);
nand U29371 (N_29371,N_26590,N_25015);
xor U29372 (N_29372,N_25652,N_26694);
nand U29373 (N_29373,N_26553,N_26638);
or U29374 (N_29374,N_27099,N_25990);
nor U29375 (N_29375,N_26925,N_27468);
nand U29376 (N_29376,N_26089,N_26151);
xnor U29377 (N_29377,N_26806,N_26587);
or U29378 (N_29378,N_26747,N_26694);
nand U29379 (N_29379,N_27404,N_27373);
and U29380 (N_29380,N_25801,N_26035);
or U29381 (N_29381,N_27358,N_25752);
xnor U29382 (N_29382,N_25411,N_25180);
nor U29383 (N_29383,N_25637,N_27021);
and U29384 (N_29384,N_26365,N_25252);
or U29385 (N_29385,N_27136,N_25109);
xnor U29386 (N_29386,N_27088,N_26632);
or U29387 (N_29387,N_27496,N_25194);
xnor U29388 (N_29388,N_25380,N_26898);
nor U29389 (N_29389,N_25112,N_25611);
and U29390 (N_29390,N_27233,N_27474);
or U29391 (N_29391,N_26893,N_26870);
and U29392 (N_29392,N_25724,N_27256);
or U29393 (N_29393,N_27411,N_25756);
nor U29394 (N_29394,N_25019,N_26035);
and U29395 (N_29395,N_26103,N_25149);
nor U29396 (N_29396,N_25997,N_26545);
or U29397 (N_29397,N_25507,N_25384);
and U29398 (N_29398,N_26842,N_26984);
or U29399 (N_29399,N_25272,N_26902);
or U29400 (N_29400,N_26364,N_25264);
xnor U29401 (N_29401,N_25406,N_26369);
xor U29402 (N_29402,N_26887,N_27062);
nor U29403 (N_29403,N_25779,N_26698);
xor U29404 (N_29404,N_25649,N_26595);
xor U29405 (N_29405,N_27275,N_26946);
xnor U29406 (N_29406,N_25375,N_25711);
or U29407 (N_29407,N_25957,N_26378);
nand U29408 (N_29408,N_26358,N_25547);
nand U29409 (N_29409,N_25116,N_26969);
nand U29410 (N_29410,N_25045,N_26634);
nand U29411 (N_29411,N_27498,N_26646);
nor U29412 (N_29412,N_27005,N_26991);
nor U29413 (N_29413,N_27231,N_26199);
nor U29414 (N_29414,N_25198,N_26881);
and U29415 (N_29415,N_25229,N_26091);
xnor U29416 (N_29416,N_25782,N_25242);
nor U29417 (N_29417,N_26780,N_25645);
nand U29418 (N_29418,N_26793,N_27113);
nand U29419 (N_29419,N_25456,N_25318);
or U29420 (N_29420,N_25363,N_26746);
nor U29421 (N_29421,N_25133,N_27394);
xnor U29422 (N_29422,N_27027,N_26385);
or U29423 (N_29423,N_27285,N_26588);
or U29424 (N_29424,N_26921,N_26101);
and U29425 (N_29425,N_25999,N_25004);
xor U29426 (N_29426,N_26790,N_26358);
nand U29427 (N_29427,N_26113,N_26935);
or U29428 (N_29428,N_27149,N_25313);
and U29429 (N_29429,N_25552,N_25138);
or U29430 (N_29430,N_25576,N_25457);
nor U29431 (N_29431,N_26166,N_25599);
and U29432 (N_29432,N_25572,N_25502);
and U29433 (N_29433,N_25153,N_26646);
nand U29434 (N_29434,N_26271,N_25947);
or U29435 (N_29435,N_26784,N_25806);
and U29436 (N_29436,N_25248,N_26202);
xnor U29437 (N_29437,N_26547,N_25689);
nor U29438 (N_29438,N_25741,N_26338);
xnor U29439 (N_29439,N_25933,N_25422);
xor U29440 (N_29440,N_26805,N_25522);
xor U29441 (N_29441,N_26964,N_26757);
nand U29442 (N_29442,N_26087,N_25095);
nand U29443 (N_29443,N_27127,N_26516);
nand U29444 (N_29444,N_25625,N_27149);
xnor U29445 (N_29445,N_26787,N_25760);
nand U29446 (N_29446,N_25478,N_26498);
or U29447 (N_29447,N_25701,N_27121);
xor U29448 (N_29448,N_27367,N_27420);
nor U29449 (N_29449,N_25745,N_25545);
nor U29450 (N_29450,N_26009,N_26018);
nand U29451 (N_29451,N_27353,N_25071);
and U29452 (N_29452,N_26380,N_26039);
nand U29453 (N_29453,N_27270,N_26707);
and U29454 (N_29454,N_26022,N_25525);
xor U29455 (N_29455,N_26228,N_25285);
or U29456 (N_29456,N_25311,N_25774);
nand U29457 (N_29457,N_27283,N_26071);
xnor U29458 (N_29458,N_26038,N_25428);
and U29459 (N_29459,N_26852,N_26387);
and U29460 (N_29460,N_26256,N_26231);
or U29461 (N_29461,N_25838,N_26017);
nand U29462 (N_29462,N_25123,N_27326);
or U29463 (N_29463,N_27447,N_25175);
nor U29464 (N_29464,N_26606,N_25265);
or U29465 (N_29465,N_25297,N_25907);
nand U29466 (N_29466,N_25400,N_26152);
and U29467 (N_29467,N_26368,N_26694);
or U29468 (N_29468,N_26861,N_25900);
or U29469 (N_29469,N_25368,N_25694);
nor U29470 (N_29470,N_25010,N_26358);
nand U29471 (N_29471,N_27005,N_27135);
nand U29472 (N_29472,N_25266,N_25397);
and U29473 (N_29473,N_25321,N_26876);
nor U29474 (N_29474,N_26304,N_25335);
or U29475 (N_29475,N_26629,N_27194);
nor U29476 (N_29476,N_27389,N_25544);
and U29477 (N_29477,N_26189,N_27093);
nor U29478 (N_29478,N_26237,N_27101);
nand U29479 (N_29479,N_26888,N_26495);
xnor U29480 (N_29480,N_26969,N_26414);
nand U29481 (N_29481,N_25631,N_27233);
nor U29482 (N_29482,N_27107,N_25711);
nor U29483 (N_29483,N_25147,N_26201);
xor U29484 (N_29484,N_27315,N_27405);
xor U29485 (N_29485,N_26344,N_26357);
or U29486 (N_29486,N_25818,N_25763);
and U29487 (N_29487,N_27408,N_26453);
nand U29488 (N_29488,N_26450,N_25208);
nor U29489 (N_29489,N_25402,N_26809);
or U29490 (N_29490,N_27484,N_26642);
and U29491 (N_29491,N_27490,N_26787);
nor U29492 (N_29492,N_26858,N_26828);
and U29493 (N_29493,N_27478,N_26623);
and U29494 (N_29494,N_25703,N_27298);
nor U29495 (N_29495,N_26049,N_25028);
or U29496 (N_29496,N_26215,N_25059);
or U29497 (N_29497,N_26101,N_26143);
xor U29498 (N_29498,N_25218,N_26696);
nand U29499 (N_29499,N_26320,N_26288);
or U29500 (N_29500,N_26032,N_27028);
nor U29501 (N_29501,N_25105,N_26429);
or U29502 (N_29502,N_25362,N_26501);
or U29503 (N_29503,N_25296,N_25971);
nor U29504 (N_29504,N_27416,N_25139);
nor U29505 (N_29505,N_27429,N_25916);
or U29506 (N_29506,N_25560,N_27381);
and U29507 (N_29507,N_25737,N_27468);
nand U29508 (N_29508,N_26691,N_26982);
nand U29509 (N_29509,N_26408,N_27294);
and U29510 (N_29510,N_25169,N_26275);
nand U29511 (N_29511,N_25987,N_26244);
xor U29512 (N_29512,N_26308,N_25186);
or U29513 (N_29513,N_26553,N_27295);
or U29514 (N_29514,N_25740,N_27229);
nand U29515 (N_29515,N_26571,N_27436);
xor U29516 (N_29516,N_26707,N_27333);
xor U29517 (N_29517,N_26185,N_27436);
and U29518 (N_29518,N_25485,N_25982);
nor U29519 (N_29519,N_26889,N_26408);
xor U29520 (N_29520,N_25918,N_27409);
nor U29521 (N_29521,N_26571,N_25433);
or U29522 (N_29522,N_25584,N_25175);
and U29523 (N_29523,N_27164,N_26873);
xor U29524 (N_29524,N_25455,N_25204);
nor U29525 (N_29525,N_27120,N_27068);
nand U29526 (N_29526,N_25609,N_25403);
and U29527 (N_29527,N_26180,N_27406);
and U29528 (N_29528,N_25190,N_25575);
and U29529 (N_29529,N_25096,N_25264);
nand U29530 (N_29530,N_25977,N_26477);
nand U29531 (N_29531,N_25402,N_25351);
and U29532 (N_29532,N_25752,N_26811);
or U29533 (N_29533,N_25332,N_25695);
xor U29534 (N_29534,N_27379,N_27352);
or U29535 (N_29535,N_25062,N_27379);
and U29536 (N_29536,N_25929,N_27256);
nand U29537 (N_29537,N_26582,N_26265);
nor U29538 (N_29538,N_27198,N_26207);
xnor U29539 (N_29539,N_26153,N_26054);
nor U29540 (N_29540,N_26508,N_26379);
nand U29541 (N_29541,N_26848,N_25277);
nor U29542 (N_29542,N_25807,N_26066);
nor U29543 (N_29543,N_27198,N_25630);
nand U29544 (N_29544,N_25253,N_25166);
nor U29545 (N_29545,N_27357,N_25579);
nor U29546 (N_29546,N_27356,N_26418);
nor U29547 (N_29547,N_25649,N_26340);
nor U29548 (N_29548,N_25246,N_26474);
nand U29549 (N_29549,N_26077,N_26625);
or U29550 (N_29550,N_25801,N_25250);
nand U29551 (N_29551,N_26766,N_26752);
and U29552 (N_29552,N_25865,N_27377);
nand U29553 (N_29553,N_25921,N_26347);
and U29554 (N_29554,N_27494,N_26185);
xor U29555 (N_29555,N_26794,N_26521);
nand U29556 (N_29556,N_27312,N_26839);
or U29557 (N_29557,N_25466,N_27359);
nor U29558 (N_29558,N_26853,N_26250);
or U29559 (N_29559,N_26215,N_25675);
and U29560 (N_29560,N_27496,N_26216);
xor U29561 (N_29561,N_26480,N_26005);
nand U29562 (N_29562,N_25183,N_26244);
or U29563 (N_29563,N_26899,N_25620);
xor U29564 (N_29564,N_26356,N_25651);
and U29565 (N_29565,N_26588,N_25568);
and U29566 (N_29566,N_25431,N_26112);
and U29567 (N_29567,N_25497,N_25344);
xnor U29568 (N_29568,N_27471,N_26246);
xor U29569 (N_29569,N_26585,N_27235);
nor U29570 (N_29570,N_26685,N_26511);
nand U29571 (N_29571,N_26436,N_26367);
xnor U29572 (N_29572,N_25704,N_25538);
nor U29573 (N_29573,N_26891,N_26998);
or U29574 (N_29574,N_27022,N_25369);
nor U29575 (N_29575,N_26303,N_27141);
or U29576 (N_29576,N_26884,N_26969);
or U29577 (N_29577,N_26073,N_27235);
nand U29578 (N_29578,N_26533,N_26891);
and U29579 (N_29579,N_27053,N_25147);
nor U29580 (N_29580,N_25786,N_26458);
and U29581 (N_29581,N_26275,N_27385);
xor U29582 (N_29582,N_26989,N_25155);
nand U29583 (N_29583,N_25908,N_27464);
xnor U29584 (N_29584,N_26509,N_26077);
nor U29585 (N_29585,N_25439,N_26165);
nand U29586 (N_29586,N_26002,N_25056);
nand U29587 (N_29587,N_25377,N_26064);
and U29588 (N_29588,N_27036,N_27137);
xor U29589 (N_29589,N_27385,N_26519);
and U29590 (N_29590,N_27166,N_25223);
nor U29591 (N_29591,N_26311,N_25689);
and U29592 (N_29592,N_26593,N_25814);
nor U29593 (N_29593,N_25142,N_25256);
xor U29594 (N_29594,N_26075,N_27238);
nand U29595 (N_29595,N_25125,N_26475);
nand U29596 (N_29596,N_25018,N_26998);
nand U29597 (N_29597,N_26003,N_26681);
and U29598 (N_29598,N_25002,N_25122);
and U29599 (N_29599,N_27107,N_25210);
or U29600 (N_29600,N_26725,N_27388);
nor U29601 (N_29601,N_25929,N_25364);
or U29602 (N_29602,N_27495,N_27470);
xor U29603 (N_29603,N_26900,N_26106);
nor U29604 (N_29604,N_25159,N_25146);
and U29605 (N_29605,N_27010,N_25430);
nand U29606 (N_29606,N_26232,N_25973);
or U29607 (N_29607,N_25573,N_25770);
xnor U29608 (N_29608,N_25475,N_26354);
and U29609 (N_29609,N_26950,N_26060);
or U29610 (N_29610,N_25270,N_25708);
and U29611 (N_29611,N_27361,N_25529);
nand U29612 (N_29612,N_26432,N_27489);
xor U29613 (N_29613,N_25369,N_27310);
xnor U29614 (N_29614,N_26305,N_27307);
or U29615 (N_29615,N_25066,N_26656);
nand U29616 (N_29616,N_26237,N_27267);
xor U29617 (N_29617,N_27015,N_27355);
nand U29618 (N_29618,N_26310,N_26457);
and U29619 (N_29619,N_25571,N_26063);
and U29620 (N_29620,N_25373,N_27169);
nor U29621 (N_29621,N_26380,N_25481);
and U29622 (N_29622,N_27281,N_25552);
nor U29623 (N_29623,N_27493,N_27161);
nor U29624 (N_29624,N_26351,N_26650);
nor U29625 (N_29625,N_26649,N_25118);
nor U29626 (N_29626,N_26905,N_26043);
and U29627 (N_29627,N_25335,N_27219);
nor U29628 (N_29628,N_25143,N_26248);
nor U29629 (N_29629,N_26847,N_27344);
nor U29630 (N_29630,N_27488,N_25174);
or U29631 (N_29631,N_25731,N_27459);
nand U29632 (N_29632,N_25429,N_25154);
nand U29633 (N_29633,N_26182,N_25051);
nor U29634 (N_29634,N_25360,N_25842);
xor U29635 (N_29635,N_25403,N_25469);
xor U29636 (N_29636,N_25723,N_27228);
nor U29637 (N_29637,N_25934,N_25929);
nand U29638 (N_29638,N_26151,N_27337);
and U29639 (N_29639,N_25072,N_25070);
or U29640 (N_29640,N_27039,N_26133);
xnor U29641 (N_29641,N_26453,N_25274);
nor U29642 (N_29642,N_26591,N_25737);
xnor U29643 (N_29643,N_26668,N_26975);
xnor U29644 (N_29644,N_26494,N_25696);
xor U29645 (N_29645,N_25239,N_26848);
nor U29646 (N_29646,N_25996,N_25682);
xor U29647 (N_29647,N_26152,N_26778);
nor U29648 (N_29648,N_27037,N_27224);
xnor U29649 (N_29649,N_27408,N_26647);
xor U29650 (N_29650,N_25689,N_27243);
nor U29651 (N_29651,N_25916,N_27145);
nor U29652 (N_29652,N_25879,N_26632);
nand U29653 (N_29653,N_25800,N_25156);
and U29654 (N_29654,N_26184,N_26150);
nor U29655 (N_29655,N_25157,N_25758);
nor U29656 (N_29656,N_26987,N_26303);
and U29657 (N_29657,N_26749,N_27367);
nand U29658 (N_29658,N_25995,N_25820);
or U29659 (N_29659,N_27481,N_25706);
and U29660 (N_29660,N_25700,N_27483);
xnor U29661 (N_29661,N_26115,N_25852);
or U29662 (N_29662,N_25223,N_26029);
or U29663 (N_29663,N_25510,N_26545);
nor U29664 (N_29664,N_26424,N_26945);
nor U29665 (N_29665,N_26700,N_26494);
or U29666 (N_29666,N_26391,N_27324);
nand U29667 (N_29667,N_26808,N_26058);
and U29668 (N_29668,N_25715,N_26544);
nand U29669 (N_29669,N_27091,N_26288);
xor U29670 (N_29670,N_26966,N_26283);
xnor U29671 (N_29671,N_26440,N_25745);
or U29672 (N_29672,N_25207,N_26785);
or U29673 (N_29673,N_26852,N_26977);
xor U29674 (N_29674,N_26769,N_26307);
nor U29675 (N_29675,N_26916,N_25067);
or U29676 (N_29676,N_25642,N_25475);
or U29677 (N_29677,N_25079,N_26670);
or U29678 (N_29678,N_25041,N_25587);
xor U29679 (N_29679,N_25696,N_27088);
and U29680 (N_29680,N_26193,N_26582);
nand U29681 (N_29681,N_25492,N_26298);
nor U29682 (N_29682,N_25403,N_26241);
xor U29683 (N_29683,N_26481,N_25656);
nand U29684 (N_29684,N_27016,N_25561);
and U29685 (N_29685,N_25217,N_26469);
nand U29686 (N_29686,N_27422,N_26787);
nand U29687 (N_29687,N_26211,N_25429);
nand U29688 (N_29688,N_26051,N_25224);
or U29689 (N_29689,N_25894,N_25511);
and U29690 (N_29690,N_25236,N_25439);
or U29691 (N_29691,N_26134,N_26432);
and U29692 (N_29692,N_25973,N_25699);
nor U29693 (N_29693,N_26186,N_27020);
xor U29694 (N_29694,N_27040,N_26432);
or U29695 (N_29695,N_27019,N_26843);
or U29696 (N_29696,N_25207,N_26981);
nand U29697 (N_29697,N_26567,N_27015);
or U29698 (N_29698,N_25995,N_25264);
nor U29699 (N_29699,N_26142,N_27032);
nor U29700 (N_29700,N_25914,N_25269);
nor U29701 (N_29701,N_27494,N_25889);
xor U29702 (N_29702,N_26574,N_26591);
xnor U29703 (N_29703,N_25871,N_26202);
nand U29704 (N_29704,N_27192,N_25607);
nor U29705 (N_29705,N_25106,N_26758);
nand U29706 (N_29706,N_26826,N_26069);
xnor U29707 (N_29707,N_27415,N_25097);
nand U29708 (N_29708,N_25008,N_25573);
nor U29709 (N_29709,N_25941,N_26660);
or U29710 (N_29710,N_25762,N_26304);
xor U29711 (N_29711,N_25452,N_25482);
and U29712 (N_29712,N_25897,N_25209);
or U29713 (N_29713,N_25756,N_26424);
nor U29714 (N_29714,N_26563,N_26987);
and U29715 (N_29715,N_26073,N_26740);
or U29716 (N_29716,N_26109,N_27347);
xor U29717 (N_29717,N_27407,N_27249);
nand U29718 (N_29718,N_25271,N_27343);
nor U29719 (N_29719,N_25792,N_25676);
xor U29720 (N_29720,N_25718,N_26277);
xor U29721 (N_29721,N_25730,N_25786);
and U29722 (N_29722,N_25100,N_25936);
nand U29723 (N_29723,N_27149,N_27130);
xor U29724 (N_29724,N_25826,N_26652);
xnor U29725 (N_29725,N_26917,N_26798);
nor U29726 (N_29726,N_26847,N_27317);
or U29727 (N_29727,N_26964,N_27148);
xor U29728 (N_29728,N_27295,N_25760);
nand U29729 (N_29729,N_26163,N_26889);
nand U29730 (N_29730,N_25448,N_25512);
nand U29731 (N_29731,N_26153,N_25783);
xor U29732 (N_29732,N_25972,N_25348);
and U29733 (N_29733,N_27498,N_25307);
nor U29734 (N_29734,N_25998,N_27332);
xor U29735 (N_29735,N_25745,N_25857);
or U29736 (N_29736,N_27119,N_27428);
nand U29737 (N_29737,N_25654,N_26880);
or U29738 (N_29738,N_25044,N_26656);
nand U29739 (N_29739,N_25481,N_27300);
xnor U29740 (N_29740,N_25975,N_26597);
nor U29741 (N_29741,N_25042,N_25581);
xor U29742 (N_29742,N_25614,N_26765);
nor U29743 (N_29743,N_25178,N_26206);
nand U29744 (N_29744,N_27201,N_27395);
or U29745 (N_29745,N_25400,N_25651);
nor U29746 (N_29746,N_27086,N_25938);
nand U29747 (N_29747,N_25298,N_27173);
and U29748 (N_29748,N_26031,N_26280);
xor U29749 (N_29749,N_26250,N_26137);
nand U29750 (N_29750,N_25109,N_26620);
or U29751 (N_29751,N_25478,N_25562);
nor U29752 (N_29752,N_26552,N_25704);
nor U29753 (N_29753,N_25350,N_26343);
and U29754 (N_29754,N_26059,N_25575);
and U29755 (N_29755,N_25654,N_25913);
and U29756 (N_29756,N_26272,N_25699);
nand U29757 (N_29757,N_25375,N_26241);
nand U29758 (N_29758,N_25658,N_26839);
nor U29759 (N_29759,N_26533,N_25936);
nand U29760 (N_29760,N_26970,N_26459);
nand U29761 (N_29761,N_26942,N_27087);
xnor U29762 (N_29762,N_26411,N_26364);
nand U29763 (N_29763,N_27193,N_27270);
xor U29764 (N_29764,N_27419,N_27227);
nand U29765 (N_29765,N_26816,N_25103);
xor U29766 (N_29766,N_26528,N_25030);
xor U29767 (N_29767,N_25543,N_25396);
nand U29768 (N_29768,N_25877,N_25197);
and U29769 (N_29769,N_27096,N_25132);
xor U29770 (N_29770,N_25749,N_27023);
or U29771 (N_29771,N_26283,N_26695);
nor U29772 (N_29772,N_27332,N_27480);
xor U29773 (N_29773,N_26359,N_26148);
xnor U29774 (N_29774,N_25861,N_26445);
nand U29775 (N_29775,N_25261,N_25826);
nand U29776 (N_29776,N_26735,N_26149);
nand U29777 (N_29777,N_26242,N_27297);
and U29778 (N_29778,N_25456,N_26184);
nand U29779 (N_29779,N_26854,N_25599);
and U29780 (N_29780,N_26942,N_26395);
nand U29781 (N_29781,N_26260,N_27085);
xor U29782 (N_29782,N_27427,N_25214);
nand U29783 (N_29783,N_27476,N_25392);
xor U29784 (N_29784,N_25491,N_26555);
nor U29785 (N_29785,N_25534,N_26406);
and U29786 (N_29786,N_27397,N_26608);
and U29787 (N_29787,N_25924,N_26827);
or U29788 (N_29788,N_25653,N_25173);
and U29789 (N_29789,N_26320,N_25229);
xor U29790 (N_29790,N_25334,N_26862);
nand U29791 (N_29791,N_26040,N_25597);
and U29792 (N_29792,N_25068,N_27398);
nor U29793 (N_29793,N_26423,N_27454);
xor U29794 (N_29794,N_27072,N_25286);
nand U29795 (N_29795,N_26909,N_27093);
and U29796 (N_29796,N_26111,N_26247);
and U29797 (N_29797,N_26796,N_25293);
or U29798 (N_29798,N_26496,N_26266);
nand U29799 (N_29799,N_25940,N_27482);
nand U29800 (N_29800,N_25549,N_26360);
nand U29801 (N_29801,N_25388,N_25003);
nand U29802 (N_29802,N_26980,N_27063);
nor U29803 (N_29803,N_26151,N_27378);
xor U29804 (N_29804,N_26076,N_26994);
xnor U29805 (N_29805,N_25150,N_25186);
nor U29806 (N_29806,N_26133,N_26052);
or U29807 (N_29807,N_25229,N_26974);
nand U29808 (N_29808,N_27014,N_26591);
nor U29809 (N_29809,N_25088,N_25669);
or U29810 (N_29810,N_27094,N_26394);
xnor U29811 (N_29811,N_25583,N_27380);
and U29812 (N_29812,N_27271,N_26136);
and U29813 (N_29813,N_25943,N_26389);
nand U29814 (N_29814,N_27155,N_26963);
or U29815 (N_29815,N_26889,N_26685);
nor U29816 (N_29816,N_25997,N_26348);
or U29817 (N_29817,N_27283,N_26907);
or U29818 (N_29818,N_26415,N_25451);
nand U29819 (N_29819,N_25473,N_27324);
nor U29820 (N_29820,N_25460,N_26547);
or U29821 (N_29821,N_27370,N_25535);
xor U29822 (N_29822,N_26250,N_25661);
or U29823 (N_29823,N_25004,N_26234);
or U29824 (N_29824,N_25922,N_25995);
nand U29825 (N_29825,N_25717,N_26083);
or U29826 (N_29826,N_25087,N_26813);
or U29827 (N_29827,N_25011,N_25630);
nor U29828 (N_29828,N_25007,N_27264);
nor U29829 (N_29829,N_26373,N_27183);
and U29830 (N_29830,N_27492,N_26806);
or U29831 (N_29831,N_25066,N_27052);
nor U29832 (N_29832,N_25051,N_27127);
nor U29833 (N_29833,N_26430,N_25623);
xor U29834 (N_29834,N_25398,N_26977);
nand U29835 (N_29835,N_26088,N_26882);
and U29836 (N_29836,N_27492,N_25737);
or U29837 (N_29837,N_27254,N_26089);
nand U29838 (N_29838,N_25443,N_26120);
nand U29839 (N_29839,N_27413,N_25892);
xnor U29840 (N_29840,N_26145,N_26264);
or U29841 (N_29841,N_25243,N_27079);
and U29842 (N_29842,N_25737,N_27104);
or U29843 (N_29843,N_25664,N_25758);
nand U29844 (N_29844,N_27335,N_26238);
nor U29845 (N_29845,N_25399,N_26023);
nor U29846 (N_29846,N_25416,N_27035);
nand U29847 (N_29847,N_26048,N_26835);
nand U29848 (N_29848,N_26529,N_25276);
and U29849 (N_29849,N_25384,N_26428);
nor U29850 (N_29850,N_26123,N_25856);
nand U29851 (N_29851,N_27053,N_25707);
nor U29852 (N_29852,N_27268,N_25535);
nor U29853 (N_29853,N_27272,N_26245);
or U29854 (N_29854,N_25423,N_26553);
or U29855 (N_29855,N_25621,N_26002);
nand U29856 (N_29856,N_25769,N_26056);
nand U29857 (N_29857,N_26203,N_26123);
nor U29858 (N_29858,N_25255,N_25385);
xnor U29859 (N_29859,N_27440,N_26956);
nor U29860 (N_29860,N_26723,N_27321);
nor U29861 (N_29861,N_25083,N_26131);
nand U29862 (N_29862,N_25504,N_25857);
xor U29863 (N_29863,N_27148,N_25741);
xnor U29864 (N_29864,N_25031,N_27201);
nor U29865 (N_29865,N_27036,N_25577);
nor U29866 (N_29866,N_27339,N_25870);
or U29867 (N_29867,N_25875,N_25402);
and U29868 (N_29868,N_26431,N_26056);
or U29869 (N_29869,N_25980,N_25989);
or U29870 (N_29870,N_26354,N_26670);
xor U29871 (N_29871,N_26045,N_25685);
xnor U29872 (N_29872,N_26500,N_26624);
nand U29873 (N_29873,N_25958,N_26264);
and U29874 (N_29874,N_25244,N_26676);
or U29875 (N_29875,N_27047,N_27013);
xnor U29876 (N_29876,N_26201,N_27043);
nand U29877 (N_29877,N_27360,N_27249);
and U29878 (N_29878,N_25736,N_27423);
or U29879 (N_29879,N_26724,N_26165);
nand U29880 (N_29880,N_25634,N_26465);
or U29881 (N_29881,N_26876,N_25990);
and U29882 (N_29882,N_27300,N_26347);
and U29883 (N_29883,N_26131,N_26197);
or U29884 (N_29884,N_25237,N_26416);
xor U29885 (N_29885,N_26784,N_25389);
xnor U29886 (N_29886,N_26925,N_26277);
xnor U29887 (N_29887,N_25874,N_27123);
or U29888 (N_29888,N_26741,N_26732);
nor U29889 (N_29889,N_25516,N_25190);
nand U29890 (N_29890,N_27477,N_25248);
and U29891 (N_29891,N_25911,N_25196);
or U29892 (N_29892,N_25377,N_25345);
or U29893 (N_29893,N_26679,N_26601);
nor U29894 (N_29894,N_26895,N_25781);
nand U29895 (N_29895,N_26665,N_26029);
xor U29896 (N_29896,N_27340,N_25189);
xnor U29897 (N_29897,N_26469,N_25344);
and U29898 (N_29898,N_27237,N_27353);
nand U29899 (N_29899,N_26279,N_27181);
xor U29900 (N_29900,N_26260,N_26085);
or U29901 (N_29901,N_27187,N_26448);
nand U29902 (N_29902,N_25217,N_26634);
or U29903 (N_29903,N_27459,N_25421);
nor U29904 (N_29904,N_26043,N_26781);
or U29905 (N_29905,N_27291,N_25792);
nor U29906 (N_29906,N_27231,N_26587);
xnor U29907 (N_29907,N_26323,N_25175);
nor U29908 (N_29908,N_27225,N_26044);
nand U29909 (N_29909,N_27484,N_25143);
nand U29910 (N_29910,N_26922,N_25545);
nand U29911 (N_29911,N_26235,N_25633);
nand U29912 (N_29912,N_25016,N_25513);
and U29913 (N_29913,N_26862,N_27122);
nand U29914 (N_29914,N_27134,N_25961);
and U29915 (N_29915,N_25336,N_25108);
nor U29916 (N_29916,N_27221,N_25459);
nand U29917 (N_29917,N_26575,N_26991);
xnor U29918 (N_29918,N_26249,N_27444);
nor U29919 (N_29919,N_26812,N_27458);
and U29920 (N_29920,N_25314,N_26385);
and U29921 (N_29921,N_25244,N_26103);
or U29922 (N_29922,N_26493,N_25908);
nand U29923 (N_29923,N_26200,N_26519);
and U29924 (N_29924,N_27185,N_26376);
or U29925 (N_29925,N_26175,N_26611);
or U29926 (N_29926,N_26306,N_26048);
or U29927 (N_29927,N_27021,N_26863);
and U29928 (N_29928,N_26431,N_27066);
and U29929 (N_29929,N_26637,N_25827);
nor U29930 (N_29930,N_25042,N_26772);
nor U29931 (N_29931,N_25919,N_26305);
nor U29932 (N_29932,N_26517,N_25243);
nor U29933 (N_29933,N_27068,N_27019);
and U29934 (N_29934,N_27239,N_25800);
nand U29935 (N_29935,N_27406,N_26885);
xor U29936 (N_29936,N_27283,N_26006);
xnor U29937 (N_29937,N_26385,N_25180);
and U29938 (N_29938,N_25728,N_26589);
xnor U29939 (N_29939,N_26923,N_25635);
and U29940 (N_29940,N_26821,N_26427);
nor U29941 (N_29941,N_27443,N_26438);
nor U29942 (N_29942,N_26525,N_26843);
nand U29943 (N_29943,N_26649,N_26421);
and U29944 (N_29944,N_26887,N_25740);
and U29945 (N_29945,N_25543,N_25149);
and U29946 (N_29946,N_25460,N_26625);
nor U29947 (N_29947,N_26101,N_27111);
xnor U29948 (N_29948,N_27498,N_26452);
nor U29949 (N_29949,N_26570,N_27245);
nor U29950 (N_29950,N_25402,N_26627);
xnor U29951 (N_29951,N_27193,N_26014);
nand U29952 (N_29952,N_26272,N_25640);
and U29953 (N_29953,N_26866,N_25127);
and U29954 (N_29954,N_26914,N_27319);
or U29955 (N_29955,N_25944,N_25407);
xor U29956 (N_29956,N_25746,N_26716);
or U29957 (N_29957,N_25595,N_25751);
xnor U29958 (N_29958,N_27090,N_27186);
nor U29959 (N_29959,N_25781,N_25978);
nand U29960 (N_29960,N_25263,N_25959);
and U29961 (N_29961,N_26517,N_25559);
nand U29962 (N_29962,N_26794,N_25321);
or U29963 (N_29963,N_27154,N_27438);
and U29964 (N_29964,N_27167,N_27249);
and U29965 (N_29965,N_26741,N_26266);
nor U29966 (N_29966,N_25695,N_27419);
and U29967 (N_29967,N_26997,N_27208);
xnor U29968 (N_29968,N_26301,N_26258);
and U29969 (N_29969,N_25924,N_26415);
nand U29970 (N_29970,N_26095,N_25058);
xor U29971 (N_29971,N_25922,N_25059);
and U29972 (N_29972,N_25525,N_26233);
and U29973 (N_29973,N_25367,N_26752);
nand U29974 (N_29974,N_26138,N_26568);
and U29975 (N_29975,N_25442,N_26807);
xnor U29976 (N_29976,N_25817,N_25170);
xnor U29977 (N_29977,N_26335,N_25893);
or U29978 (N_29978,N_25469,N_26814);
and U29979 (N_29979,N_26908,N_25398);
nand U29980 (N_29980,N_26071,N_25664);
xor U29981 (N_29981,N_26347,N_26210);
nand U29982 (N_29982,N_25803,N_25842);
xnor U29983 (N_29983,N_27243,N_26904);
nor U29984 (N_29984,N_27279,N_25676);
or U29985 (N_29985,N_25717,N_26946);
nor U29986 (N_29986,N_26597,N_27137);
nand U29987 (N_29987,N_26115,N_26011);
and U29988 (N_29988,N_27354,N_27420);
nor U29989 (N_29989,N_27370,N_26477);
or U29990 (N_29990,N_25342,N_27016);
or U29991 (N_29991,N_27411,N_25614);
nand U29992 (N_29992,N_26703,N_26064);
nor U29993 (N_29993,N_26286,N_25271);
xor U29994 (N_29994,N_26106,N_25742);
nor U29995 (N_29995,N_25572,N_25526);
nor U29996 (N_29996,N_26281,N_25242);
nor U29997 (N_29997,N_25837,N_26465);
nor U29998 (N_29998,N_25650,N_27189);
or U29999 (N_29999,N_25246,N_26169);
xnor U30000 (N_30000,N_28290,N_29762);
or U30001 (N_30001,N_27968,N_27681);
nand U30002 (N_30002,N_29784,N_28927);
xnor U30003 (N_30003,N_29840,N_28673);
nand U30004 (N_30004,N_29754,N_28850);
nand U30005 (N_30005,N_28041,N_28883);
and U30006 (N_30006,N_29594,N_29978);
xnor U30007 (N_30007,N_28768,N_28536);
and U30008 (N_30008,N_29715,N_28879);
nor U30009 (N_30009,N_29801,N_29935);
xor U30010 (N_30010,N_27874,N_29134);
nand U30011 (N_30011,N_29422,N_29703);
or U30012 (N_30012,N_27908,N_27522);
and U30013 (N_30013,N_29753,N_28366);
nand U30014 (N_30014,N_28208,N_29377);
xnor U30015 (N_30015,N_28378,N_28990);
or U30016 (N_30016,N_28655,N_28097);
and U30017 (N_30017,N_28310,N_29323);
or U30018 (N_30018,N_29729,N_27887);
xnor U30019 (N_30019,N_29218,N_28389);
xor U30020 (N_30020,N_28585,N_29354);
and U30021 (N_30021,N_27628,N_29358);
xor U30022 (N_30022,N_28452,N_29999);
nor U30023 (N_30023,N_28816,N_28792);
nor U30024 (N_30024,N_27899,N_29239);
or U30025 (N_30025,N_27748,N_29448);
or U30026 (N_30026,N_28151,N_27745);
and U30027 (N_30027,N_27756,N_28566);
and U30028 (N_30028,N_28147,N_27867);
and U30029 (N_30029,N_27790,N_29351);
and U30030 (N_30030,N_29771,N_28004);
and U30031 (N_30031,N_28778,N_29327);
and U30032 (N_30032,N_28257,N_28034);
and U30033 (N_30033,N_27610,N_29603);
or U30034 (N_30034,N_28423,N_29975);
xor U30035 (N_30035,N_28739,N_29251);
nor U30036 (N_30036,N_27843,N_29942);
nand U30037 (N_30037,N_29770,N_29882);
nor U30038 (N_30038,N_28613,N_27783);
nand U30039 (N_30039,N_27836,N_28232);
nand U30040 (N_30040,N_28849,N_27816);
nand U30041 (N_30041,N_29020,N_27923);
nand U30042 (N_30042,N_28973,N_28829);
nand U30043 (N_30043,N_29839,N_29936);
or U30044 (N_30044,N_29657,N_28149);
xor U30045 (N_30045,N_27630,N_29705);
or U30046 (N_30046,N_27654,N_28909);
xnor U30047 (N_30047,N_27655,N_29044);
or U30048 (N_30048,N_29699,N_28868);
xor U30049 (N_30049,N_29930,N_29141);
nand U30050 (N_30050,N_29662,N_28709);
nand U30051 (N_30051,N_28839,N_29332);
and U30052 (N_30052,N_27729,N_29062);
nor U30053 (N_30053,N_29861,N_28334);
or U30054 (N_30054,N_28763,N_29056);
and U30055 (N_30055,N_27549,N_28193);
and U30056 (N_30056,N_28002,N_29099);
or U30057 (N_30057,N_29996,N_28790);
or U30058 (N_30058,N_29535,N_28560);
nor U30059 (N_30059,N_27513,N_29842);
nand U30060 (N_30060,N_29880,N_28797);
nor U30061 (N_30061,N_28029,N_28450);
xor U30062 (N_30062,N_28157,N_28510);
nand U30063 (N_30063,N_29819,N_29776);
nand U30064 (N_30064,N_27953,N_28307);
or U30065 (N_30065,N_28812,N_29916);
nor U30066 (N_30066,N_28710,N_28602);
and U30067 (N_30067,N_27632,N_29574);
or U30068 (N_30068,N_29871,N_28210);
xor U30069 (N_30069,N_28875,N_29960);
nand U30070 (N_30070,N_29234,N_28730);
and U30071 (N_30071,N_29410,N_28220);
and U30072 (N_30072,N_29449,N_28747);
or U30073 (N_30073,N_29441,N_29206);
xor U30074 (N_30074,N_29627,N_29115);
nand U30075 (N_30075,N_29273,N_27502);
nand U30076 (N_30076,N_29922,N_28171);
and U30077 (N_30077,N_28779,N_28652);
and U30078 (N_30078,N_29797,N_28793);
xor U30079 (N_30079,N_29809,N_29287);
and U30080 (N_30080,N_29268,N_28644);
nor U30081 (N_30081,N_28794,N_27557);
nand U30082 (N_30082,N_27539,N_28016);
nor U30083 (N_30083,N_28174,N_28687);
nand U30084 (N_30084,N_29944,N_27798);
and U30085 (N_30085,N_27944,N_29101);
nand U30086 (N_30086,N_29676,N_29479);
nand U30087 (N_30087,N_27648,N_29624);
or U30088 (N_30088,N_29411,N_28375);
nand U30089 (N_30089,N_29316,N_28876);
or U30090 (N_30090,N_29154,N_28035);
or U30091 (N_30091,N_29976,N_28489);
nand U30092 (N_30092,N_29367,N_28825);
or U30093 (N_30093,N_28328,N_27730);
nor U30094 (N_30094,N_29997,N_29275);
or U30095 (N_30095,N_28444,N_29238);
xor U30096 (N_30096,N_29046,N_29526);
or U30097 (N_30097,N_29029,N_29602);
and U30098 (N_30098,N_29290,N_28425);
nor U30099 (N_30099,N_29910,N_29897);
xor U30100 (N_30100,N_27869,N_28067);
or U30101 (N_30101,N_28595,N_29734);
and U30102 (N_30102,N_29452,N_27698);
nand U30103 (N_30103,N_28482,N_28531);
xor U30104 (N_30104,N_28690,N_29051);
nor U30105 (N_30105,N_29660,N_29952);
nor U30106 (N_30106,N_28660,N_29259);
and U30107 (N_30107,N_28820,N_29277);
and U30108 (N_30108,N_29274,N_28640);
or U30109 (N_30109,N_27870,N_29878);
nand U30110 (N_30110,N_28507,N_28350);
xor U30111 (N_30111,N_29236,N_27823);
or U30112 (N_30112,N_27863,N_27937);
xor U30113 (N_30113,N_29262,N_28718);
nand U30114 (N_30114,N_29495,N_28442);
or U30115 (N_30115,N_27709,N_29249);
nor U30116 (N_30116,N_27677,N_27912);
and U30117 (N_30117,N_29061,N_29445);
nand U30118 (N_30118,N_28471,N_28961);
nor U30119 (N_30119,N_28209,N_29844);
xor U30120 (N_30120,N_28217,N_28700);
or U30121 (N_30121,N_28024,N_29924);
or U30122 (N_30122,N_29356,N_29196);
xor U30123 (N_30123,N_28873,N_27845);
xor U30124 (N_30124,N_29565,N_28649);
nor U30125 (N_30125,N_28132,N_29625);
or U30126 (N_30126,N_27857,N_28242);
and U30127 (N_30127,N_28666,N_29832);
nor U30128 (N_30128,N_29547,N_28126);
nand U30129 (N_30129,N_29352,N_29836);
and U30130 (N_30130,N_28661,N_27743);
xor U30131 (N_30131,N_28871,N_28179);
nor U30132 (N_30132,N_27533,N_29483);
or U30133 (N_30133,N_28827,N_29132);
nand U30134 (N_30134,N_29938,N_28413);
nor U30135 (N_30135,N_28599,N_27925);
xnor U30136 (N_30136,N_28196,N_28060);
nor U30137 (N_30137,N_27515,N_28087);
or U30138 (N_30138,N_28459,N_28299);
xnor U30139 (N_30139,N_27639,N_28971);
and U30140 (N_30140,N_27817,N_28386);
nand U30141 (N_30141,N_28059,N_29900);
or U30142 (N_30142,N_28913,N_28994);
or U30143 (N_30143,N_29515,N_28705);
nand U30144 (N_30144,N_28924,N_29455);
xor U30145 (N_30145,N_29429,N_27560);
nor U30146 (N_30146,N_27651,N_28456);
and U30147 (N_30147,N_27961,N_29042);
nor U30148 (N_30148,N_29641,N_27771);
nor U30149 (N_30149,N_27517,N_29623);
nand U30150 (N_30150,N_29747,N_29365);
or U30151 (N_30151,N_27693,N_29962);
nand U30152 (N_30152,N_28601,N_29985);
nor U30153 (N_30153,N_27896,N_28997);
nand U30154 (N_30154,N_27721,N_29025);
xnor U30155 (N_30155,N_27919,N_28582);
or U30156 (N_30156,N_27852,N_28108);
and U30157 (N_30157,N_28771,N_28751);
or U30158 (N_30158,N_29873,N_29718);
or U30159 (N_30159,N_28342,N_28250);
or U30160 (N_30160,N_29690,N_28504);
and U30161 (N_30161,N_29125,N_29442);
xnor U30162 (N_30162,N_28557,N_28055);
or U30163 (N_30163,N_29870,N_27685);
nand U30164 (N_30164,N_29570,N_29851);
nand U30165 (N_30165,N_27956,N_28317);
or U30166 (N_30166,N_28499,N_28138);
xor U30167 (N_30167,N_27930,N_29482);
xor U30168 (N_30168,N_29189,N_29163);
nand U30169 (N_30169,N_29988,N_28937);
xor U30170 (N_30170,N_28623,N_29925);
nand U30171 (N_30171,N_29970,N_28239);
nor U30172 (N_30172,N_28866,N_29263);
or U30173 (N_30173,N_27580,N_29566);
and U30174 (N_30174,N_28096,N_29890);
or U30175 (N_30175,N_29955,N_29773);
xor U30176 (N_30176,N_28720,N_29158);
xnor U30177 (N_30177,N_29689,N_27650);
or U30178 (N_30178,N_29194,N_29473);
xnor U30179 (N_30179,N_28135,N_28934);
or U30180 (N_30180,N_28134,N_29853);
nor U30181 (N_30181,N_29629,N_29752);
nand U30182 (N_30182,N_28194,N_29255);
and U30183 (N_30183,N_28611,N_29301);
nor U30184 (N_30184,N_29685,N_29708);
or U30185 (N_30185,N_28983,N_28010);
nand U30186 (N_30186,N_28339,N_29270);
nor U30187 (N_30187,N_28956,N_28119);
nand U30188 (N_30188,N_29169,N_29510);
nor U30189 (N_30189,N_28938,N_29122);
nor U30190 (N_30190,N_28026,N_29959);
and U30191 (N_30191,N_28648,N_29611);
or U30192 (N_30192,N_28515,N_28377);
nand U30193 (N_30193,N_28053,N_29898);
nand U30194 (N_30194,N_28206,N_28363);
and U30195 (N_30195,N_29070,N_27747);
and U30196 (N_30196,N_28335,N_27744);
nor U30197 (N_30197,N_29181,N_29892);
nor U30198 (N_30198,N_28033,N_28270);
nor U30199 (N_30199,N_29427,N_28845);
xor U30200 (N_30200,N_28619,N_28943);
nor U30201 (N_30201,N_27775,N_29969);
xor U30202 (N_30202,N_29133,N_27605);
or U30203 (N_30203,N_28449,N_29039);
nand U30204 (N_30204,N_29179,N_28926);
or U30205 (N_30205,N_27976,N_29912);
or U30206 (N_30206,N_28104,N_29655);
and U30207 (N_30207,N_28214,N_29100);
and U30208 (N_30208,N_27678,N_28609);
and U30209 (N_30209,N_27931,N_29310);
nand U30210 (N_30210,N_28738,N_28650);
xor U30211 (N_30211,N_27621,N_29644);
or U30212 (N_30212,N_29469,N_29406);
nand U30213 (N_30213,N_29972,N_28732);
nor U30214 (N_30214,N_28929,N_29027);
nand U30215 (N_30215,N_27697,N_28397);
nor U30216 (N_30216,N_29011,N_29185);
nor U30217 (N_30217,N_28205,N_27584);
nor U30218 (N_30218,N_29470,N_28407);
nand U30219 (N_30219,N_29030,N_28524);
xor U30220 (N_30220,N_27773,N_28427);
and U30221 (N_30221,N_29383,N_28184);
nand U30222 (N_30222,N_29137,N_29545);
nand U30223 (N_30223,N_28643,N_29531);
nand U30224 (N_30224,N_29764,N_29738);
nor U30225 (N_30225,N_29360,N_27609);
nor U30226 (N_30226,N_29182,N_29775);
nand U30227 (N_30227,N_27914,N_27714);
nor U30228 (N_30228,N_28384,N_27544);
nand U30229 (N_30229,N_29394,N_28505);
xor U30230 (N_30230,N_27703,N_28548);
nand U30231 (N_30231,N_28562,N_29845);
or U30232 (N_30232,N_29677,N_28360);
or U30233 (N_30233,N_28908,N_29084);
nor U30234 (N_30234,N_29678,N_29331);
or U30235 (N_30235,N_28767,N_28326);
and U30236 (N_30236,N_27971,N_29079);
nor U30237 (N_30237,N_29034,N_28960);
or U30238 (N_30238,N_29405,N_27757);
or U30239 (N_30239,N_28392,N_27599);
xnor U30240 (N_30240,N_29369,N_28600);
and U30241 (N_30241,N_29297,N_28668);
or U30242 (N_30242,N_27873,N_29119);
nor U30243 (N_30243,N_29060,N_28563);
or U30244 (N_30244,N_27841,N_29103);
or U30245 (N_30245,N_29608,N_29437);
nor U30246 (N_30246,N_29192,N_28857);
and U30247 (N_30247,N_28261,N_28945);
or U30248 (N_30248,N_28109,N_29187);
xnor U30249 (N_30249,N_29457,N_28801);
or U30250 (N_30250,N_29120,N_27543);
nor U30251 (N_30251,N_27905,N_29626);
xnor U30252 (N_30252,N_27601,N_29081);
nand U30253 (N_30253,N_28914,N_28021);
nand U30254 (N_30254,N_28882,N_28915);
xnor U30255 (N_30255,N_28382,N_28519);
and U30256 (N_30256,N_27571,N_27928);
nand U30257 (N_30257,N_28251,N_29830);
nand U30258 (N_30258,N_28796,N_29386);
xnor U30259 (N_30259,N_27789,N_29471);
or U30260 (N_30260,N_29589,N_29013);
or U30261 (N_30261,N_27797,N_29325);
nor U30262 (N_30262,N_28224,N_29697);
xnor U30263 (N_30263,N_28967,N_27606);
xnor U30264 (N_30264,N_27828,N_29211);
and U30265 (N_30265,N_29069,N_29344);
nor U30266 (N_30266,N_28745,N_28725);
and U30267 (N_30267,N_28786,N_29146);
nand U30268 (N_30268,N_29083,N_28461);
nor U30269 (N_30269,N_28852,N_29663);
xor U30270 (N_30270,N_28300,N_28361);
xnor U30271 (N_30271,N_29649,N_28422);
and U30272 (N_30272,N_29711,N_28155);
nor U30273 (N_30273,N_27746,N_29478);
nor U30274 (N_30274,N_28030,N_27766);
nand U30275 (N_30275,N_27786,N_29907);
and U30276 (N_30276,N_28818,N_29906);
nand U30277 (N_30277,N_27694,N_29739);
or U30278 (N_30278,N_29981,N_29317);
nand U30279 (N_30279,N_29281,N_28981);
nor U30280 (N_30280,N_28586,N_28991);
and U30281 (N_30281,N_29090,N_28588);
or U30282 (N_30282,N_28365,N_29528);
nand U30283 (N_30283,N_28027,N_28735);
or U30284 (N_30284,N_28932,N_29516);
and U30285 (N_30285,N_28176,N_29347);
or U30286 (N_30286,N_28003,N_29184);
nand U30287 (N_30287,N_29918,N_27612);
nor U30288 (N_30288,N_28127,N_28410);
nor U30289 (N_30289,N_29229,N_29186);
nand U30290 (N_30290,N_29698,N_28547);
and U30291 (N_30291,N_28411,N_29476);
nand U30292 (N_30292,N_29917,N_29064);
or U30293 (N_30293,N_28530,N_29859);
nor U30294 (N_30294,N_28780,N_27827);
nand U30295 (N_30295,N_28085,N_28417);
nand U30296 (N_30296,N_27634,N_29811);
and U30297 (N_30297,N_28851,N_28014);
nor U30298 (N_30298,N_29214,N_28736);
nor U30299 (N_30299,N_28574,N_29459);
nand U30300 (N_30300,N_29901,N_28729);
nand U30301 (N_30301,N_28216,N_27755);
nor U30302 (N_30302,N_29203,N_29195);
nand U30303 (N_30303,N_27615,N_27734);
or U30304 (N_30304,N_28697,N_28128);
and U30305 (N_30305,N_29709,N_29760);
or U30306 (N_30306,N_28597,N_29140);
xnor U30307 (N_30307,N_28589,N_29884);
and U30308 (N_30308,N_27529,N_27579);
nor U30309 (N_30309,N_27578,N_28102);
and U30310 (N_30310,N_29318,N_28570);
nor U30311 (N_30311,N_28789,N_28090);
nor U30312 (N_30312,N_28269,N_27569);
or U30313 (N_30313,N_28698,N_28150);
nor U30314 (N_30314,N_28762,N_28869);
or U30315 (N_30315,N_28841,N_27988);
xor U30316 (N_30316,N_27531,N_28190);
and U30317 (N_30317,N_29105,N_29075);
and U30318 (N_30318,N_27687,N_27715);
nand U30319 (N_30319,N_27565,N_28374);
nand U30320 (N_30320,N_28722,N_29648);
xor U30321 (N_30321,N_28884,N_28169);
xnor U30322 (N_30322,N_27717,N_28670);
nor U30323 (N_30323,N_29393,N_29583);
nand U30324 (N_30324,N_28188,N_28110);
or U30325 (N_30325,N_28622,N_27812);
nand U30326 (N_30326,N_29491,N_28520);
and U30327 (N_30327,N_27883,N_28187);
and U30328 (N_30328,N_28291,N_27970);
xor U30329 (N_30329,N_29587,N_29359);
nand U30330 (N_30330,N_28833,N_29050);
nor U30331 (N_30331,N_28688,N_27768);
nand U30332 (N_30332,N_29379,N_29043);
nor U30333 (N_30333,N_29706,N_29235);
xnor U30334 (N_30334,N_29872,N_29823);
nor U30335 (N_30335,N_29951,N_29364);
xor U30336 (N_30336,N_28100,N_28592);
or U30337 (N_30337,N_28322,N_29191);
and U30338 (N_30338,N_28741,N_28638);
nand U30339 (N_30339,N_28508,N_28534);
and U30340 (N_30340,N_27758,N_28606);
nor U30341 (N_30341,N_28153,N_29588);
or U30342 (N_30342,N_28996,N_28432);
or U30343 (N_30343,N_29803,N_29201);
nand U30344 (N_30344,N_27826,N_29756);
and U30345 (N_30345,N_29131,N_28404);
or U30346 (N_30346,N_28254,N_29399);
nand U30347 (N_30347,N_28440,N_29554);
xor U30348 (N_30348,N_28754,N_28921);
nand U30349 (N_30349,N_29835,N_27975);
nand U30350 (N_30350,N_29487,N_27573);
xor U30351 (N_30351,N_28861,N_29546);
or U30352 (N_30352,N_29597,N_27538);
xnor U30353 (N_30353,N_28028,N_29401);
and U30354 (N_30354,N_29593,N_29374);
and U30355 (N_30355,N_28313,N_28941);
xnor U30356 (N_30356,N_29544,N_27951);
or U30357 (N_30357,N_28364,N_29642);
or U30358 (N_30358,N_28145,N_29609);
nand U30359 (N_30359,N_27878,N_27851);
xor U30360 (N_30360,N_28158,N_29102);
nand U30361 (N_30361,N_29048,N_29923);
or U30362 (N_30362,N_27680,N_29205);
xnor U30363 (N_30363,N_27889,N_28554);
nor U30364 (N_30364,N_29741,N_29866);
xnor U30365 (N_30365,N_28315,N_28703);
and U30366 (N_30366,N_29643,N_28071);
xnor U30367 (N_30367,N_28910,N_27804);
xor U30368 (N_30368,N_29646,N_28620);
nor U30369 (N_30369,N_29885,N_27591);
nor U30370 (N_30370,N_28864,N_28788);
or U30371 (N_30371,N_28704,N_29382);
nor U30372 (N_30372,N_29926,N_27737);
nand U30373 (N_30373,N_29390,N_27646);
nor U30374 (N_30374,N_28509,N_28618);
xor U30375 (N_30375,N_27722,N_27659);
or U30376 (N_30376,N_29311,N_28830);
nor U30377 (N_30377,N_29717,N_29765);
nand U30378 (N_30378,N_27991,N_29578);
nand U30379 (N_30379,N_28347,N_29232);
or U30380 (N_30380,N_29198,N_28069);
xor U30381 (N_30381,N_27770,N_29296);
and U30382 (N_30382,N_28180,N_29078);
or U30383 (N_30383,N_27710,N_27589);
xor U30384 (N_30384,N_29782,N_29108);
nor U30385 (N_30385,N_28823,N_29568);
nor U30386 (N_30386,N_28162,N_29984);
xnor U30387 (N_30387,N_29306,N_28419);
nand U30388 (N_30388,N_28354,N_29571);
and U30389 (N_30389,N_28918,N_28919);
and U30390 (N_30390,N_28634,N_28498);
nand U30391 (N_30391,N_28175,N_28603);
nor U30392 (N_30392,N_28222,N_27563);
nor U30393 (N_30393,N_28072,N_27832);
nor U30394 (N_30394,N_29336,N_28874);
and U30395 (N_30395,N_28266,N_28332);
nand U30396 (N_30396,N_28486,N_28737);
nand U30397 (N_30397,N_28327,N_29855);
nor U30398 (N_30398,N_28658,N_28048);
nor U30399 (N_30399,N_28112,N_27566);
and U30400 (N_30400,N_27927,N_28324);
or U30401 (N_30401,N_27506,N_29204);
nand U30402 (N_30402,N_29053,N_28713);
and U30403 (N_30403,N_28063,N_27752);
or U30404 (N_30404,N_29126,N_28795);
nand U30405 (N_30405,N_28296,N_28716);
nor U30406 (N_30406,N_28993,N_29990);
nand U30407 (N_30407,N_28409,N_28744);
nor U30408 (N_30408,N_27625,N_27787);
or U30409 (N_30409,N_27886,N_29421);
xor U30410 (N_30410,N_27683,N_28541);
xor U30411 (N_30411,N_28939,N_27906);
or U30412 (N_30412,N_27781,N_29438);
nand U30413 (N_30413,N_28159,N_28715);
xnor U30414 (N_30414,N_28646,N_28931);
nor U30415 (N_30415,N_29014,N_29927);
nor U30416 (N_30416,N_29291,N_28408);
nor U30417 (N_30417,N_29914,N_28316);
nor U30418 (N_30418,N_29233,N_29921);
or U30419 (N_30419,N_28944,N_27933);
and U30420 (N_30420,N_28312,N_28942);
nor U30421 (N_30421,N_29564,N_28107);
and U30422 (N_30422,N_28974,N_29790);
nand U30423 (N_30423,N_28799,N_27893);
or U30424 (N_30424,N_29726,N_28154);
or U30425 (N_30425,N_27884,N_29054);
nand U30426 (N_30426,N_29414,N_29856);
nand U30427 (N_30427,N_27809,N_28032);
nand U30428 (N_30428,N_29142,N_29400);
nand U30429 (N_30429,N_29579,N_29831);
and U30430 (N_30430,N_27728,N_29742);
nand U30431 (N_30431,N_27969,N_29007);
nand U30432 (N_30432,N_28936,N_28353);
and U30433 (N_30433,N_27846,N_28044);
xor U30434 (N_30434,N_28359,N_28479);
xor U30435 (N_30435,N_27830,N_28630);
and U30436 (N_30436,N_27963,N_28228);
or U30437 (N_30437,N_29017,N_29431);
xnor U30438 (N_30438,N_27541,N_28051);
xnor U30439 (N_30439,N_27540,N_27686);
xor U30440 (N_30440,N_27998,N_29197);
nor U30441 (N_30441,N_28679,N_27725);
nor U30442 (N_30442,N_28947,N_28962);
nand U30443 (N_30443,N_28772,N_29439);
xor U30444 (N_30444,N_29504,N_27922);
and U30445 (N_30445,N_28262,N_29658);
xor U30446 (N_30446,N_27920,N_27695);
or U30447 (N_30447,N_28237,N_28278);
nand U30448 (N_30448,N_28441,N_29692);
nor U30449 (N_30449,N_29006,N_29964);
xnor U30450 (N_30450,N_27972,N_28989);
nand U30451 (N_30451,N_27911,N_28572);
nand U30452 (N_30452,N_28241,N_28529);
xnor U30453 (N_30453,N_28707,N_29049);
nand U30454 (N_30454,N_29622,N_28629);
nor U30455 (N_30455,N_28007,N_29143);
nand U30456 (N_30456,N_28084,N_27572);
xnor U30457 (N_30457,N_28822,N_29063);
xnor U30458 (N_30458,N_28966,N_29758);
and U30459 (N_30459,N_28766,N_29569);
xnor U30460 (N_30460,N_29932,N_27716);
and U30461 (N_30461,N_28682,N_28678);
xor U30462 (N_30462,N_29633,N_29465);
xor U30463 (N_30463,N_29877,N_27806);
or U30464 (N_30464,N_27800,N_28231);
nand U30465 (N_30465,N_29059,N_29228);
xnor U30466 (N_30466,N_28500,N_29598);
or U30467 (N_30467,N_29313,N_28587);
and U30468 (N_30468,N_29168,N_27759);
xnor U30469 (N_30469,N_28046,N_27608);
nor U30470 (N_30470,N_27818,N_29869);
and U30471 (N_30471,N_28274,N_29072);
nand U30472 (N_30472,N_29580,N_29177);
nor U30473 (N_30473,N_28975,N_28211);
and U30474 (N_30474,N_27568,N_27967);
xor U30475 (N_30475,N_29695,N_28683);
and U30476 (N_30476,N_29787,N_29763);
and U30477 (N_30477,N_29493,N_29982);
or U30478 (N_30478,N_28140,N_28118);
nor U30479 (N_30479,N_28819,N_29434);
nand U30480 (N_30480,N_29389,N_28267);
nand U30481 (N_30481,N_28746,N_29650);
xor U30482 (N_30482,N_28385,N_29794);
nor U30483 (N_30483,N_28433,N_29761);
or U30484 (N_30484,N_28025,N_27973);
nor U30485 (N_30485,N_28197,N_28170);
nand U30486 (N_30486,N_28593,N_27671);
and U30487 (N_30487,N_29664,N_29616);
and U30488 (N_30488,N_29555,N_28412);
nor U30489 (N_30489,N_28052,N_28391);
nand U30490 (N_30490,N_29208,N_28474);
nor U30491 (N_30491,N_27949,N_29328);
nor U30492 (N_30492,N_29601,N_29019);
nand U30493 (N_30493,N_27624,N_27880);
xnor U30494 (N_30494,N_28284,N_28415);
nand U30495 (N_30495,N_29973,N_28259);
xor U30496 (N_30496,N_28495,N_28305);
or U30497 (N_30497,N_29857,N_27892);
nor U30498 (N_30498,N_28659,N_27704);
and U30499 (N_30499,N_28785,N_29582);
xor U30500 (N_30500,N_28828,N_29968);
and U30501 (N_30501,N_28058,N_29303);
and U30502 (N_30502,N_28577,N_27813);
nor U30503 (N_30503,N_28447,N_27966);
nor U30504 (N_30504,N_28526,N_29684);
nor U30505 (N_30505,N_29654,N_29418);
and U30506 (N_30506,N_29333,N_28293);
nand U30507 (N_30507,N_29378,N_27801);
nor U30508 (N_30508,N_28020,N_28692);
nand U30509 (N_30509,N_29710,N_29826);
or U30510 (N_30510,N_29501,N_29507);
xor U30511 (N_30511,N_29004,N_29802);
xor U30512 (N_30512,N_28632,N_28677);
and U30513 (N_30513,N_28596,N_28331);
nor U30514 (N_30514,N_29145,N_28068);
nand U30515 (N_30515,N_28846,N_29221);
nor U30516 (N_30516,N_29852,N_29505);
or U30517 (N_30517,N_29796,N_27888);
and U30518 (N_30518,N_27633,N_29575);
or U30519 (N_30519,N_29606,N_29326);
nand U30520 (N_30520,N_28393,N_29879);
nand U30521 (N_30521,N_29675,N_29118);
or U30522 (N_30522,N_27850,N_29159);
nor U30523 (N_30523,N_28949,N_27640);
or U30524 (N_30524,N_29097,N_27611);
or U30525 (N_30525,N_29180,N_28418);
nor U30526 (N_30526,N_28635,N_28164);
and U30527 (N_30527,N_28213,N_27751);
nor U30528 (N_30528,N_28287,N_29392);
and U30529 (N_30529,N_29243,N_28755);
nor U30530 (N_30530,N_28605,N_27712);
xor U30531 (N_30531,N_27838,N_29015);
or U30532 (N_30532,N_27731,N_27629);
and U30533 (N_30533,N_29402,N_27957);
and U30534 (N_30534,N_29702,N_28985);
xor U30535 (N_30535,N_28776,N_29965);
and U30536 (N_30536,N_27807,N_29462);
xor U30537 (N_30537,N_29966,N_29451);
nor U30538 (N_30538,N_29634,N_28093);
nand U30539 (N_30539,N_28379,N_29943);
or U30540 (N_30540,N_27932,N_28598);
xor U30541 (N_30541,N_28223,N_29368);
xnor U30542 (N_30542,N_27727,N_29160);
nor U30543 (N_30543,N_29267,N_29357);
and U30544 (N_30544,N_28528,N_29172);
nor U30545 (N_30545,N_28240,N_27581);
nor U30546 (N_30546,N_29903,N_28693);
nor U30547 (N_30547,N_28146,N_27943);
xnor U30548 (N_30548,N_28922,N_27637);
nand U30549 (N_30549,N_29928,N_29166);
and U30550 (N_30550,N_29604,N_28463);
nor U30551 (N_30551,N_28856,N_27987);
and U30552 (N_30552,N_27992,N_28064);
xor U30553 (N_30553,N_29319,N_29147);
nand U30554 (N_30554,N_27576,N_29456);
or U30555 (N_30555,N_29216,N_27954);
nor U30556 (N_30556,N_28920,N_29686);
and U30557 (N_30557,N_29018,N_27959);
or U30558 (N_30558,N_29315,N_28338);
and U30559 (N_30559,N_28626,N_28544);
and U30560 (N_30560,N_28079,N_28674);
xnor U30561 (N_30561,N_28472,N_28610);
nand U30562 (N_30562,N_29033,N_28901);
and U30563 (N_30563,N_29241,N_29798);
or U30564 (N_30564,N_27736,N_28302);
and U30565 (N_30565,N_28621,N_28724);
nor U30566 (N_30566,N_29110,N_27985);
or U30567 (N_30567,N_29176,N_28198);
xnor U30568 (N_30568,N_28457,N_29212);
and U30569 (N_30569,N_29888,N_28923);
or U30570 (N_30570,N_29735,N_28708);
nand U30571 (N_30571,N_29614,N_27519);
or U30572 (N_30572,N_28466,N_28464);
xnor U30573 (N_30573,N_29638,N_29816);
or U30574 (N_30574,N_29577,N_27950);
or U30575 (N_30575,N_29058,N_28912);
xnor U30576 (N_30576,N_28428,N_29785);
or U30577 (N_30577,N_29111,N_29672);
nand U30578 (N_30578,N_28847,N_29227);
or U30579 (N_30579,N_29149,N_29789);
nor U30580 (N_30580,N_27670,N_28243);
nand U30581 (N_30581,N_29993,N_27501);
and U30582 (N_30582,N_29373,N_27718);
xnor U30583 (N_30583,N_29444,N_28834);
nand U30584 (N_30584,N_28401,N_29783);
nor U30585 (N_30585,N_29428,N_29939);
nand U30586 (N_30586,N_29067,N_29671);
nand U30587 (N_30587,N_28897,N_27512);
nand U30588 (N_30588,N_27616,N_28383);
and U30589 (N_30589,N_29745,N_27891);
or U30590 (N_30590,N_28639,N_28191);
or U30591 (N_30591,N_29862,N_27649);
nand U30592 (N_30592,N_28821,N_28054);
nand U30593 (N_30593,N_29355,N_29586);
nand U30594 (N_30594,N_28671,N_29694);
xor U30595 (N_30595,N_27839,N_28227);
nand U30596 (N_30596,N_27780,N_28657);
xnor U30597 (N_30597,N_29696,N_29971);
nor U30598 (N_30598,N_27929,N_29276);
or U30599 (N_30599,N_28022,N_27772);
or U30600 (N_30600,N_27527,N_27849);
nor U30601 (N_30601,N_28131,N_27511);
and U30602 (N_30602,N_28451,N_29635);
and U30603 (N_30603,N_28402,N_28694);
or U30604 (N_30604,N_28455,N_29631);
or U30605 (N_30605,N_29256,N_28764);
or U30606 (N_30606,N_28229,N_29781);
and U30607 (N_30607,N_29723,N_29945);
xor U30608 (N_30608,N_28236,N_28283);
nor U30609 (N_30609,N_27674,N_29213);
nand U30610 (N_30610,N_28935,N_29460);
or U30611 (N_30611,N_29065,N_28045);
nor U30612 (N_30612,N_29512,N_29237);
nand U30613 (N_30613,N_28731,N_29931);
nand U30614 (N_30614,N_28832,N_29525);
xor U30615 (N_30615,N_28759,N_29534);
nor U30616 (N_30616,N_29911,N_27915);
nand U30617 (N_30617,N_29028,N_28000);
xor U30618 (N_30618,N_28802,N_28387);
nand U30619 (N_30619,N_28750,N_28902);
xnor U30620 (N_30620,N_29559,N_29562);
xor U30621 (N_30621,N_27618,N_28454);
or U30622 (N_30622,N_28123,N_29584);
xor U30623 (N_30623,N_28089,N_28065);
nor U30624 (N_30624,N_28578,N_27794);
and U30625 (N_30625,N_29052,N_28181);
and U30626 (N_30626,N_28323,N_28273);
or U30627 (N_30627,N_28406,N_29161);
and U30628 (N_30628,N_28523,N_28113);
nand U30629 (N_30629,N_28928,N_28614);
nand U30630 (N_30630,N_29596,N_28120);
xnor U30631 (N_30631,N_29813,N_29958);
and U30632 (N_30632,N_28564,N_27530);
nor U30633 (N_30633,N_29324,N_28341);
or U30634 (N_30634,N_28311,N_28483);
or U30635 (N_30635,N_29541,N_27877);
nand U30636 (N_30636,N_29138,N_28761);
nor U30637 (N_30637,N_29810,N_27622);
and U30638 (N_30638,N_28448,N_29308);
nand U30639 (N_30639,N_27776,N_28245);
nor U30640 (N_30640,N_28781,N_28421);
nand U30641 (N_30641,N_29388,N_29808);
nor U30642 (N_30642,N_28314,N_29489);
and U30643 (N_30643,N_27795,N_28867);
xor U30644 (N_30644,N_29834,N_28556);
nand U30645 (N_30645,N_29337,N_28878);
or U30646 (N_30646,N_28047,N_29567);
nand U30647 (N_30647,N_27941,N_29155);
nor U30648 (N_30648,N_29755,N_29223);
or U30649 (N_30649,N_29674,N_27881);
nand U30650 (N_30650,N_28330,N_27982);
or U30651 (N_30651,N_29843,N_27577);
nand U30652 (N_30652,N_28318,N_28163);
and U30653 (N_30653,N_28414,N_28512);
nor U30654 (N_30654,N_29795,N_27868);
nor U30655 (N_30655,N_28809,N_27567);
and U30656 (N_30656,N_28142,N_27667);
nand U30657 (N_30657,N_27684,N_28189);
xnor U30658 (N_30658,N_29381,N_29557);
xor U30659 (N_30659,N_29563,N_28695);
and U30660 (N_30660,N_28437,N_27754);
nand U30661 (N_30661,N_28552,N_29467);
or U30662 (N_30662,N_28105,N_29961);
nand U30663 (N_30663,N_27814,N_28980);
nor U30664 (N_30664,N_27521,N_27672);
xor U30665 (N_30665,N_27871,N_29659);
or U30666 (N_30666,N_29037,N_29751);
or U30667 (N_30667,N_29165,N_27641);
or U30668 (N_30668,N_29009,N_28995);
nor U30669 (N_30669,N_29095,N_28977);
nor U30670 (N_30670,N_28168,N_27894);
or U30671 (N_30671,N_28465,N_28824);
nand U30672 (N_30672,N_28031,N_28631);
or U30673 (N_30673,N_29068,N_28039);
xnor U30674 (N_30674,N_28775,N_29524);
nand U30675 (N_30675,N_29670,N_27810);
nand U30676 (N_30676,N_27902,N_28309);
or U30677 (N_30677,N_27844,N_29265);
nand U30678 (N_30678,N_29591,N_29940);
and U30679 (N_30679,N_28356,N_29704);
nor U30680 (N_30680,N_28485,N_28854);
nor U30681 (N_30681,N_28037,N_28185);
and U30682 (N_30682,N_29117,N_27924);
nand U30683 (N_30683,N_29613,N_27983);
nand U30684 (N_30684,N_29683,N_27948);
or U30685 (N_30685,N_28271,N_29934);
or U30686 (N_30686,N_28742,N_29980);
and U30687 (N_30687,N_29391,N_28667);
and U30688 (N_30688,N_29883,N_27854);
xnor U30689 (N_30689,N_29701,N_27926);
nor U30690 (N_30690,N_27864,N_29335);
nor U30691 (N_30691,N_27815,N_28487);
nor U30692 (N_30692,N_29886,N_28049);
xor U30693 (N_30693,N_28445,N_29610);
nand U30694 (N_30694,N_29730,N_27829);
nand U30695 (N_30695,N_27575,N_27546);
nor U30696 (N_30696,N_29219,N_27520);
nor U30697 (N_30697,N_28351,N_28320);
or U30698 (N_30698,N_28358,N_29620);
or U30699 (N_30699,N_28279,N_28958);
or U30700 (N_30700,N_29987,N_29653);
nand U30701 (N_30701,N_29736,N_27668);
or U30702 (N_30702,N_27947,N_28207);
nand U30703 (N_30703,N_27981,N_27960);
or U30704 (N_30704,N_29466,N_29248);
nor U30705 (N_30705,N_27675,N_27696);
or U30706 (N_30706,N_28013,N_27890);
xor U30707 (N_30707,N_28172,N_28800);
nand U30708 (N_30708,N_28686,N_28911);
or U30709 (N_30709,N_27700,N_27711);
nand U30710 (N_30710,N_27993,N_29094);
and U30711 (N_30711,N_29016,N_27613);
or U30712 (N_30712,N_29271,N_27825);
and U30713 (N_30713,N_29330,N_28858);
or U30714 (N_30714,N_29074,N_29714);
nand U30715 (N_30715,N_27514,N_29908);
nand U30716 (N_30716,N_27861,N_27562);
nand U30717 (N_30717,N_29136,N_28984);
and U30718 (N_30718,N_27750,N_28062);
nor U30719 (N_30719,N_29778,N_28390);
xnor U30720 (N_30720,N_28581,N_28545);
nor U30721 (N_30721,N_27765,N_28787);
nor U30722 (N_30722,N_28247,N_29423);
nand U30723 (N_30723,N_28019,N_28853);
xor U30724 (N_30724,N_28855,N_29384);
or U30725 (N_30725,N_29385,N_27647);
and U30726 (N_30726,N_28651,N_28805);
or U30727 (N_30727,N_29419,N_27962);
nand U30728 (N_30728,N_28798,N_29225);
or U30729 (N_30729,N_29342,N_28702);
xor U30730 (N_30730,N_29494,N_29986);
or U30731 (N_30731,N_27936,N_27834);
or U30732 (N_30732,N_29114,N_28804);
xnor U30733 (N_30733,N_28144,N_28352);
nand U30734 (N_30734,N_29250,N_27691);
nand U30735 (N_30735,N_29055,N_28439);
nand U30736 (N_30736,N_29600,N_29791);
xnor U30737 (N_30737,N_29523,N_28865);
and U30738 (N_30738,N_28183,N_28001);
and U30739 (N_30739,N_29639,N_29837);
or U30740 (N_30740,N_27824,N_29086);
or U30741 (N_30741,N_28916,N_27767);
and U30742 (N_30742,N_29948,N_29967);
nand U30743 (N_30743,N_29891,N_29314);
nand U30744 (N_30744,N_27600,N_29849);
nor U30745 (N_30745,N_29599,N_28357);
nor U30746 (N_30746,N_27921,N_28496);
xnor U30747 (N_30747,N_29066,N_28959);
and U30748 (N_30748,N_29957,N_29759);
and U30749 (N_30749,N_29403,N_29107);
and U30750 (N_30750,N_29680,N_28612);
nor U30751 (N_30751,N_28607,N_27741);
nor U30752 (N_30752,N_28116,N_27708);
nor U30753 (N_30753,N_29170,N_28098);
and U30754 (N_30754,N_29230,N_27623);
xnor U30755 (N_30755,N_29109,N_28399);
nor U30756 (N_30756,N_29687,N_28723);
nor U30757 (N_30757,N_28863,N_29553);
xnor U30758 (N_30758,N_28543,N_29498);
nand U30759 (N_30759,N_29135,N_29130);
nand U30760 (N_30760,N_29630,N_27733);
xor U30761 (N_30761,N_29521,N_29619);
and U30762 (N_30762,N_28717,N_29171);
xor U30763 (N_30763,N_29889,N_28337);
nand U30764 (N_30764,N_27532,N_28280);
nand U30765 (N_30765,N_28125,N_29397);
nor U30766 (N_30766,N_29533,N_29148);
nor U30767 (N_30767,N_27554,N_27500);
and U30768 (N_30768,N_29963,N_28156);
and U30769 (N_30769,N_29607,N_27631);
and U30770 (N_30770,N_29731,N_28182);
nand U30771 (N_30771,N_28838,N_28148);
and U30772 (N_30772,N_29417,N_28129);
or U30773 (N_30773,N_28009,N_29651);
nand U30774 (N_30774,N_29278,N_27597);
nor U30775 (N_30775,N_29800,N_28576);
xor U30776 (N_30776,N_29707,N_28438);
nor U30777 (N_30777,N_29991,N_28617);
nor U30778 (N_30778,N_27535,N_29804);
or U30779 (N_30779,N_29026,N_28734);
nand U30780 (N_30780,N_29345,N_28757);
or U30781 (N_30781,N_27935,N_28301);
nand U30782 (N_30782,N_27796,N_29652);
nor U30783 (N_30783,N_29284,N_27586);
and U30784 (N_30784,N_29157,N_27587);
xnor U30785 (N_30785,N_29175,N_28950);
or U30786 (N_30786,N_29209,N_28518);
nand U30787 (N_30787,N_29618,N_27552);
nand U30788 (N_30788,N_29590,N_29838);
xor U30789 (N_30789,N_28553,N_29280);
and U30790 (N_30790,N_27661,N_29300);
nor U30791 (N_30791,N_29261,N_27652);
nor U30792 (N_30792,N_28369,N_28538);
and U30793 (N_30793,N_28376,N_29244);
or U30794 (N_30794,N_27688,N_29612);
and U30795 (N_30795,N_27910,N_27989);
xor U30796 (N_30796,N_29304,N_29003);
and U30797 (N_30797,N_27862,N_28468);
nor U30798 (N_30798,N_28549,N_28542);
nor U30799 (N_30799,N_28292,N_28740);
or U30800 (N_30800,N_28195,N_27763);
and U30801 (N_30801,N_27853,N_28532);
nand U30802 (N_30802,N_28130,N_27882);
nand U30803 (N_30803,N_27875,N_28573);
xnor U30804 (N_30804,N_29665,N_29749);
nor U30805 (N_30805,N_29661,N_28711);
nand U30806 (N_30806,N_29713,N_28685);
nor U30807 (N_30807,N_27555,N_29436);
or U30808 (N_30808,N_28862,N_29502);
or U30809 (N_30809,N_28405,N_28264);
and U30810 (N_30810,N_27833,N_28083);
nor U30811 (N_30811,N_29121,N_29092);
nand U30812 (N_30812,N_29164,N_29412);
nand U30813 (N_30813,N_29468,N_29766);
nand U30814 (N_30814,N_29581,N_28281);
nor U30815 (N_30815,N_29520,N_27561);
xnor U30816 (N_30816,N_29288,N_28050);
or U30817 (N_30817,N_28616,N_28388);
nor U30818 (N_30818,N_29572,N_27505);
nor U30819 (N_30819,N_28891,N_29833);
or U30820 (N_30820,N_29363,N_28590);
nor U30821 (N_30821,N_28712,N_28040);
or U30822 (N_30822,N_28807,N_29071);
or U30823 (N_30823,N_29712,N_28551);
xnor U30824 (N_30824,N_27822,N_28645);
nand U30825 (N_30825,N_28770,N_28727);
or U30826 (N_30826,N_27986,N_28304);
nor U30827 (N_30827,N_28372,N_29874);
nor U30828 (N_30828,N_28699,N_27821);
nand U30829 (N_30829,N_28691,N_29461);
nor U30830 (N_30830,N_27627,N_28511);
nand U30831 (N_30831,N_28462,N_29002);
xnor U30832 (N_30832,N_29517,N_29350);
nand U30833 (N_30833,N_28066,N_27916);
nand U30834 (N_30834,N_28167,N_28880);
xor U30835 (N_30835,N_29031,N_28430);
and U30836 (N_30836,N_28558,N_29091);
nor U30837 (N_30837,N_28579,N_28680);
and U30838 (N_30838,N_28870,N_28077);
or U30839 (N_30839,N_29190,N_27707);
nand U30840 (N_30840,N_28760,N_28346);
and U30841 (N_30841,N_28092,N_28061);
xor U30842 (N_30842,N_28753,N_29700);
nor U30843 (N_30843,N_27588,N_28057);
xor U30844 (N_30844,N_29681,N_28380);
xnor U30845 (N_30845,N_28978,N_27663);
nand U30846 (N_30846,N_27979,N_29539);
or U30847 (N_30847,N_28490,N_28056);
nand U30848 (N_30848,N_27556,N_28396);
and U30849 (N_30849,N_28111,N_28080);
or U30850 (N_30850,N_29899,N_29724);
nor U30851 (N_30851,N_29812,N_28636);
xnor U30852 (N_30852,N_28743,N_28426);
nor U30853 (N_30853,N_27900,N_29113);
and U30854 (N_30854,N_28905,N_28591);
nand U30855 (N_30855,N_29032,N_28319);
and U30856 (N_30856,N_28888,N_29777);
nand U30857 (N_30857,N_29343,N_29561);
nand U30858 (N_30858,N_29258,N_27799);
nor U30859 (N_30859,N_29519,N_29104);
and U30860 (N_30860,N_29983,N_28235);
or U30861 (N_30861,N_29408,N_27699);
nand U30862 (N_30862,N_29041,N_27779);
or U30863 (N_30863,N_29640,N_27673);
nand U30864 (N_30864,N_29500,N_28748);
nor U30865 (N_30865,N_28416,N_27996);
and U30866 (N_30866,N_29302,N_29780);
nor U30867 (N_30867,N_29127,N_28791);
or U30868 (N_30868,N_27848,N_29371);
nand U30869 (N_30869,N_28238,N_29806);
nor U30870 (N_30870,N_29173,N_29788);
or U30871 (N_30871,N_29088,N_28204);
nand U30872 (N_30872,N_27598,N_29518);
nor U30873 (N_30873,N_28953,N_28349);
or U30874 (N_30874,N_29024,N_29224);
xnor U30875 (N_30875,N_27895,N_29824);
nor U30876 (N_30876,N_29484,N_29740);
nand U30877 (N_30877,N_27666,N_28783);
nand U30878 (N_30878,N_29820,N_27545);
xor U30879 (N_30879,N_27534,N_28446);
nand U30880 (N_30880,N_29321,N_28933);
and U30881 (N_30881,N_28899,N_27676);
or U30882 (N_30882,N_28212,N_28895);
and U30883 (N_30883,N_27604,N_27701);
and U30884 (N_30884,N_29721,N_29667);
xor U30885 (N_30885,N_28308,N_29617);
xor U30886 (N_30886,N_27990,N_27551);
nand U30887 (N_30887,N_27999,N_29279);
nor U30888 (N_30888,N_28963,N_28930);
or U30889 (N_30889,N_27885,N_29576);
nand U30890 (N_30890,N_28663,N_28215);
nand U30891 (N_30891,N_28329,N_29669);
nand U30892 (N_30892,N_27958,N_29691);
or U30893 (N_30893,N_29772,N_29424);
and U30894 (N_30894,N_29450,N_28886);
or U30895 (N_30895,N_29266,N_28469);
and U30896 (N_30896,N_28202,N_29503);
xnor U30897 (N_30897,N_28256,N_29786);
xnor U30898 (N_30898,N_27753,N_29492);
or U30899 (N_30899,N_27713,N_28493);
nor U30900 (N_30900,N_29226,N_28782);
nand U30901 (N_30901,N_27620,N_28954);
or U30902 (N_30902,N_29294,N_28070);
nor U30903 (N_30903,N_29481,N_29949);
xnor U30904 (N_30904,N_27645,N_28917);
xor U30905 (N_30905,N_28970,N_27855);
or U30906 (N_30906,N_28263,N_27917);
nor U30907 (N_30907,N_29454,N_28494);
and U30908 (N_30908,N_29010,N_27574);
and U30909 (N_30909,N_29953,N_29286);
nand U30910 (N_30910,N_27516,N_28719);
xor U30911 (N_30911,N_29396,N_29472);
nor U30912 (N_30912,N_27508,N_28073);
nor U30913 (N_30913,N_29375,N_28403);
nand U30914 (N_30914,N_29035,N_28647);
nand U30915 (N_30915,N_29905,N_28103);
and U30916 (N_30916,N_27811,N_27723);
nand U30917 (N_30917,N_27974,N_28628);
xnor U30918 (N_30918,N_29757,N_28594);
or U30919 (N_30919,N_27792,N_29497);
nor U30920 (N_30920,N_28252,N_28343);
nor U30921 (N_30921,N_27547,N_29021);
xor U30922 (N_30922,N_28294,N_29348);
nand U30923 (N_30923,N_29252,N_28230);
or U30924 (N_30924,N_28896,N_28475);
xor U30925 (N_30925,N_29038,N_29413);
nor U30926 (N_30926,N_28481,N_27784);
nand U30927 (N_30927,N_28583,N_27720);
or U30928 (N_30928,N_28831,N_27558);
nand U30929 (N_30929,N_29805,N_29864);
or U30930 (N_30930,N_28460,N_27945);
nor U30931 (N_30931,N_29913,N_28166);
xnor U30932 (N_30932,N_28124,N_27706);
nor U30933 (N_30933,N_29254,N_27682);
nand U30934 (N_30934,N_27657,N_29199);
xor U30935 (N_30935,N_28844,N_29769);
nand U30936 (N_30936,N_28840,N_29919);
nor U30937 (N_30937,N_29240,N_29283);
nor U30938 (N_30938,N_27719,N_28203);
nand U30939 (N_30939,N_29174,N_27643);
xor U30940 (N_30940,N_27803,N_28199);
nand U30941 (N_30941,N_29152,N_29719);
and U30942 (N_30942,N_27542,N_27550);
nor U30943 (N_30943,N_29666,N_29085);
or U30944 (N_30944,N_29339,N_28139);
nor U30945 (N_30945,N_28076,N_28749);
nand U30946 (N_30946,N_28435,N_29814);
and U30947 (N_30947,N_28952,N_29464);
or U30948 (N_30948,N_29693,N_29902);
xor U30949 (N_30949,N_27980,N_27965);
nor U30950 (N_30950,N_29779,N_27984);
xor U30951 (N_30951,N_29846,N_28503);
nand U30952 (N_30952,N_29298,N_29728);
or U30953 (N_30953,N_28774,N_28999);
nand U30954 (N_30954,N_29615,N_29128);
nor U30955 (N_30955,N_28675,N_28018);
and U30956 (N_30956,N_29727,N_29167);
nand U30957 (N_30957,N_29430,N_29994);
nor U30958 (N_30958,N_28615,N_27653);
and U30959 (N_30959,N_29881,N_28453);
and U30960 (N_30960,N_27977,N_29477);
xnor U30961 (N_30961,N_29380,N_27802);
and U30962 (N_30962,N_29867,N_29305);
nand U30963 (N_30963,N_28470,N_29123);
nand U30964 (N_30964,N_27596,N_29822);
xor U30965 (N_30965,N_28122,N_27669);
and U30966 (N_30966,N_27664,N_28492);
and U30967 (N_30967,N_27865,N_29679);
xnor U30968 (N_30968,N_29001,N_28502);
and U30969 (N_30969,N_28826,N_29527);
nand U30970 (N_30970,N_28161,N_29047);
nor U30971 (N_30971,N_28373,N_28141);
nand U30972 (N_30972,N_27918,N_29552);
xor U30973 (N_30973,N_28484,N_27837);
nor U30974 (N_30974,N_28561,N_28303);
and U30975 (N_30975,N_29904,N_28811);
or U30976 (N_30976,N_29605,N_29320);
nor U30977 (N_30977,N_29496,N_28081);
xnor U30978 (N_30978,N_27978,N_28584);
or U30979 (N_30979,N_29933,N_29376);
and U30980 (N_30980,N_28728,N_28137);
xnor U30981 (N_30981,N_28226,N_29220);
or U30982 (N_30982,N_29875,N_28260);
nand U30983 (N_30983,N_29909,N_29807);
xor U30984 (N_30984,N_28525,N_29372);
xnor U30985 (N_30985,N_27738,N_28367);
nand U30986 (N_30986,N_28539,N_27840);
nand U30987 (N_30987,N_29341,N_28082);
and U30988 (N_30988,N_29817,N_29946);
or U30989 (N_30989,N_29511,N_28976);
nand U30990 (N_30990,N_28306,N_27898);
nor U30991 (N_30991,N_27689,N_29012);
and U30992 (N_30992,N_28815,N_27583);
xnor U30993 (N_30993,N_29089,N_29860);
or U30994 (N_30994,N_29329,N_28681);
nor U30995 (N_30995,N_29257,N_29895);
nor U30996 (N_30996,N_27872,N_27964);
xor U30997 (N_30997,N_27724,N_28992);
and U30998 (N_30998,N_27594,N_27507);
and U30999 (N_30999,N_27791,N_28756);
and U31000 (N_31000,N_27997,N_28522);
xor U31001 (N_31001,N_28516,N_29139);
and U31002 (N_31002,N_29950,N_28143);
and U31003 (N_31003,N_27548,N_29551);
or U31004 (N_31004,N_29036,N_28043);
nor U31005 (N_31005,N_27774,N_29475);
or U31006 (N_31006,N_27656,N_27582);
nor U31007 (N_31007,N_28881,N_29370);
xor U31008 (N_31008,N_28276,N_28368);
xnor U31009 (N_31009,N_29792,N_28925);
xnor U31010 (N_31010,N_28042,N_28769);
and U31011 (N_31011,N_28488,N_28642);
or U31012 (N_31012,N_28117,N_28443);
nand U31013 (N_31013,N_28192,N_29941);
nor U31014 (N_31014,N_28624,N_29876);
nor U31015 (N_31015,N_28400,N_29894);
nand U31016 (N_31016,N_27570,N_29560);
xnor U31017 (N_31017,N_28477,N_29242);
xnor U31018 (N_31018,N_29178,N_27907);
nor U31019 (N_31019,N_28398,N_29992);
nor U31020 (N_31020,N_28219,N_27858);
nor U31021 (N_31021,N_27994,N_29144);
or U31022 (N_31022,N_29989,N_28177);
or U31023 (N_31023,N_28808,N_29847);
nor U31024 (N_31024,N_28817,N_28608);
nand U31025 (N_31025,N_28604,N_29621);
nand U31026 (N_31026,N_29282,N_29150);
nor U31027 (N_31027,N_28654,N_28969);
or U31028 (N_31028,N_28903,N_27820);
and U31029 (N_31029,N_29977,N_29420);
xnor U31030 (N_31030,N_28458,N_28957);
xor U31031 (N_31031,N_29542,N_27847);
xnor U31032 (N_31032,N_28706,N_28012);
and U31033 (N_31033,N_28546,N_28355);
nand U31034 (N_31034,N_29744,N_28672);
and U31035 (N_31035,N_29536,N_27842);
xnor U31036 (N_31036,N_29737,N_28773);
and U31037 (N_31037,N_28806,N_28165);
or U31038 (N_31038,N_28848,N_28633);
and U31039 (N_31039,N_28265,N_29954);
nand U31040 (N_31040,N_29293,N_28894);
nand U31041 (N_31041,N_29260,N_28656);
xor U31042 (N_31042,N_29513,N_29887);
and U31043 (N_31043,N_29156,N_28892);
and U31044 (N_31044,N_28288,N_28258);
nor U31045 (N_31045,N_29264,N_28431);
nor U31046 (N_31046,N_28424,N_28095);
nand U31047 (N_31047,N_28434,N_28955);
and U31048 (N_31048,N_27879,N_29415);
nand U31049 (N_31049,N_28491,N_29509);
xor U31050 (N_31050,N_29285,N_29463);
nand U31051 (N_31051,N_29443,N_29682);
nand U31052 (N_31052,N_28765,N_28420);
xor U31053 (N_31053,N_29312,N_29543);
or U31054 (N_31054,N_27602,N_29480);
xor U31055 (N_31055,N_27702,N_29558);
or U31056 (N_31056,N_29040,N_28835);
or U31057 (N_31057,N_27679,N_29748);
xor U31058 (N_31058,N_29116,N_29956);
xnor U31059 (N_31059,N_28664,N_28115);
or U31060 (N_31060,N_28381,N_29947);
nor U31061 (N_31061,N_29404,N_29995);
or U31062 (N_31062,N_28289,N_29433);
nand U31063 (N_31063,N_27904,N_29124);
xor U31064 (N_31064,N_29750,N_27705);
nand U31065 (N_31065,N_28571,N_29829);
or U31066 (N_31066,N_28075,N_29863);
nor U31067 (N_31067,N_28133,N_29722);
or U31068 (N_31068,N_29767,N_28429);
or U31069 (N_31069,N_28565,N_27595);
nand U31070 (N_31070,N_28803,N_29338);
and U31071 (N_31071,N_27860,N_29499);
and U31072 (N_31072,N_28979,N_28467);
or U31073 (N_31073,N_29409,N_28965);
nand U31074 (N_31074,N_29151,N_29082);
or U31075 (N_31075,N_28814,N_28298);
or U31076 (N_31076,N_29425,N_29362);
nand U31077 (N_31077,N_28336,N_28218);
and U31078 (N_31078,N_27553,N_27537);
nand U31079 (N_31079,N_29854,N_29077);
nor U31080 (N_31080,N_29207,N_29446);
nor U31081 (N_31081,N_27636,N_29096);
or U31082 (N_31082,N_28178,N_28998);
nor U31083 (N_31083,N_29474,N_28889);
or U31084 (N_31084,N_28842,N_28906);
or U31085 (N_31085,N_28275,N_28005);
nor U31086 (N_31086,N_28653,N_29508);
and U31087 (N_31087,N_29087,N_28669);
nand U31088 (N_31088,N_28497,N_29057);
or U31089 (N_31089,N_29349,N_27509);
or U31090 (N_31090,N_28988,N_29269);
xnor U31091 (N_31091,N_29720,N_28255);
nor U31092 (N_31092,N_28885,N_29538);
nor U31093 (N_31093,N_28837,N_28784);
or U31094 (N_31094,N_27503,N_29307);
xor U31095 (N_31095,N_27536,N_29825);
and U31096 (N_31096,N_27564,N_28186);
or U31097 (N_31097,N_28282,N_29080);
nor U31098 (N_31098,N_28836,N_29548);
nand U31099 (N_31099,N_28810,N_28714);
nor U31100 (N_31100,N_27660,N_27617);
nand U31101 (N_31101,N_29929,N_29000);
nor U31102 (N_31102,N_27866,N_28940);
or U31103 (N_31103,N_29628,N_27585);
or U31104 (N_31104,N_28676,N_29743);
xor U31105 (N_31105,N_28907,N_27638);
and U31106 (N_31106,N_28555,N_27805);
nor U31107 (N_31107,N_29129,N_27518);
nor U31108 (N_31108,N_29073,N_29896);
and U31109 (N_31109,N_28086,N_28501);
nor U31110 (N_31110,N_28733,N_27749);
or U31111 (N_31111,N_27626,N_27510);
xnor U31112 (N_31112,N_29868,N_28964);
nand U31113 (N_31113,N_28244,N_27740);
or U31114 (N_31114,N_29022,N_28106);
or U31115 (N_31115,N_29556,N_27690);
nand U31116 (N_31116,N_29716,N_27939);
and U31117 (N_31117,N_29295,N_29529);
xnor U31118 (N_31118,N_29416,N_27658);
nor U31119 (N_31119,N_29632,N_29595);
and U31120 (N_31120,N_27739,N_28559);
nor U31121 (N_31121,N_27955,N_29246);
nand U31122 (N_31122,N_28568,N_28696);
and U31123 (N_31123,N_28550,N_28344);
nand U31124 (N_31124,N_29645,N_29112);
and U31125 (N_31125,N_29387,N_29215);
nor U31126 (N_31126,N_29733,N_29045);
nor U31127 (N_31127,N_28887,N_28535);
or U31128 (N_31128,N_28225,N_28099);
or U31129 (N_31129,N_27614,N_28843);
and U31130 (N_31130,N_29398,N_27764);
xnor U31131 (N_31131,N_29106,N_29202);
nor U31132 (N_31132,N_28091,N_27619);
xor U31133 (N_31133,N_28234,N_28517);
xnor U31134 (N_31134,N_28567,N_29153);
nor U31135 (N_31135,N_27742,N_29793);
nor U31136 (N_31136,N_28982,N_28627);
and U31137 (N_31137,N_28114,N_29725);
xnor U31138 (N_31138,N_29023,N_28684);
or U31139 (N_31139,N_27946,N_28394);
nand U31140 (N_31140,N_29231,N_29407);
or U31141 (N_31141,N_29093,N_28637);
nor U31142 (N_31142,N_29937,N_28752);
or U31143 (N_31143,N_27793,N_29309);
nand U31144 (N_31144,N_28537,N_27859);
or U31145 (N_31145,N_28362,N_28286);
nand U31146 (N_31146,N_29893,N_28898);
nor U31147 (N_31147,N_27735,N_29289);
nor U31148 (N_31148,N_28689,N_29076);
and U31149 (N_31149,N_29573,N_28023);
and U31150 (N_31150,N_28272,N_29162);
xor U31151 (N_31151,N_29200,N_28038);
nand U31152 (N_31152,N_28348,N_28860);
nand U31153 (N_31153,N_29668,N_29486);
or U31154 (N_31154,N_28268,N_29532);
xnor U31155 (N_31155,N_29636,N_28580);
nand U31156 (N_31156,N_28987,N_28521);
nand U31157 (N_31157,N_28011,N_27504);
or U31158 (N_31158,N_29768,N_27603);
nand U31159 (N_31159,N_28527,N_27903);
xor U31160 (N_31160,N_27635,N_28074);
or U31161 (N_31161,N_27785,N_28904);
and U31162 (N_31162,N_29292,N_29827);
nor U31163 (N_31163,N_29183,N_29818);
nor U31164 (N_31164,N_28478,N_28008);
or U31165 (N_31165,N_29490,N_28721);
xnor U31166 (N_31166,N_27909,N_29647);
nand U31167 (N_31167,N_27761,N_29815);
and U31168 (N_31168,N_27940,N_28948);
xor U31169 (N_31169,N_28859,N_29828);
or U31170 (N_31170,N_29732,N_29299);
or U31171 (N_31171,N_28036,N_27662);
and U31172 (N_31172,N_28370,N_28777);
and U31173 (N_31173,N_27835,N_29637);
xnor U31174 (N_31174,N_28701,N_29530);
and U31175 (N_31175,N_29488,N_28249);
nor U31176 (N_31176,N_29550,N_28946);
and U31177 (N_31177,N_29585,N_29453);
nand U31178 (N_31178,N_29920,N_27808);
or U31179 (N_31179,N_27876,N_28533);
and U31180 (N_31180,N_27665,N_28088);
nor U31181 (N_31181,N_29322,N_29253);
or U31182 (N_31182,N_27524,N_28395);
nand U31183 (N_31183,N_29673,N_28662);
xor U31184 (N_31184,N_28893,N_29361);
nor U31185 (N_31185,N_27607,N_28872);
xnor U31186 (N_31186,N_29440,N_28877);
nor U31187 (N_31187,N_28986,N_27769);
nor U31188 (N_31188,N_28152,N_27523);
nand U31189 (N_31189,N_27593,N_29247);
xor U31190 (N_31190,N_28248,N_28201);
nand U31191 (N_31191,N_28371,N_29850);
nand U31192 (N_31192,N_29865,N_28160);
and U31193 (N_31193,N_27778,N_29098);
nor U31194 (N_31194,N_28078,N_28285);
nor U31195 (N_31195,N_29746,N_27726);
or U31196 (N_31196,N_27526,N_28321);
nand U31197 (N_31197,N_29979,N_27592);
nand U31198 (N_31198,N_28625,N_29506);
or U31199 (N_31199,N_28514,N_29799);
or U31200 (N_31200,N_29549,N_28136);
xor U31201 (N_31201,N_29217,N_29210);
nor U31202 (N_31202,N_29353,N_29821);
nor U31203 (N_31203,N_27901,N_27897);
nand U31204 (N_31204,N_27782,N_28345);
xnor U31205 (N_31205,N_29537,N_28513);
nand U31206 (N_31206,N_29008,N_27528);
nand U31207 (N_31207,N_28200,N_29188);
nand U31208 (N_31208,N_28575,N_27760);
or U31209 (N_31209,N_28758,N_29656);
and U31210 (N_31210,N_29395,N_27642);
nor U31211 (N_31211,N_28813,N_27913);
nor U31212 (N_31212,N_28325,N_29592);
and U31213 (N_31213,N_28006,N_28173);
and U31214 (N_31214,N_29858,N_27692);
or U31215 (N_31215,N_29522,N_27938);
xnor U31216 (N_31216,N_29998,N_27942);
nand U31217 (N_31217,N_28726,N_29447);
and U31218 (N_31218,N_28101,N_29915);
xor U31219 (N_31219,N_28665,N_28641);
xor U31220 (N_31220,N_29688,N_29340);
and U31221 (N_31221,N_29485,N_28253);
xor U31222 (N_31222,N_28017,N_28951);
nor U31223 (N_31223,N_29193,N_28972);
and U31224 (N_31224,N_28221,N_28569);
or U31225 (N_31225,N_27559,N_28015);
xnor U31226 (N_31226,N_29272,N_28295);
nand U31227 (N_31227,N_28540,N_27788);
nor U31228 (N_31228,N_28506,N_29435);
nand U31229 (N_31229,N_27831,N_27590);
xnor U31230 (N_31230,N_28436,N_27644);
and U31231 (N_31231,N_29774,N_29346);
xor U31232 (N_31232,N_27934,N_28297);
nor U31233 (N_31233,N_28121,N_28277);
nor U31234 (N_31234,N_28473,N_29005);
xnor U31235 (N_31235,N_28333,N_29245);
and U31236 (N_31236,N_29426,N_28246);
nor U31237 (N_31237,N_29334,N_28480);
nor U31238 (N_31238,N_27952,N_27525);
and U31239 (N_31239,N_29432,N_29458);
nand U31240 (N_31240,N_29540,N_28968);
xor U31241 (N_31241,N_27762,N_27995);
nor U31242 (N_31242,N_27819,N_29514);
or U31243 (N_31243,N_29366,N_29974);
or U31244 (N_31244,N_28094,N_27856);
and U31245 (N_31245,N_29848,N_27777);
nand U31246 (N_31246,N_28900,N_28890);
and U31247 (N_31247,N_29222,N_28476);
xnor U31248 (N_31248,N_28340,N_29841);
and U31249 (N_31249,N_27732,N_28233);
nor U31250 (N_31250,N_28366,N_27822);
or U31251 (N_31251,N_28082,N_29278);
or U31252 (N_31252,N_28569,N_28875);
or U31253 (N_31253,N_27964,N_28312);
nand U31254 (N_31254,N_29371,N_28007);
or U31255 (N_31255,N_29405,N_29638);
and U31256 (N_31256,N_27703,N_29858);
or U31257 (N_31257,N_27510,N_27501);
or U31258 (N_31258,N_28603,N_29011);
nand U31259 (N_31259,N_29117,N_28865);
and U31260 (N_31260,N_29614,N_29386);
and U31261 (N_31261,N_27602,N_27765);
nor U31262 (N_31262,N_29467,N_29729);
xnor U31263 (N_31263,N_28219,N_28921);
nor U31264 (N_31264,N_27614,N_28428);
or U31265 (N_31265,N_28088,N_28260);
xor U31266 (N_31266,N_29520,N_29803);
nand U31267 (N_31267,N_28510,N_28794);
or U31268 (N_31268,N_29014,N_29007);
nand U31269 (N_31269,N_28559,N_29832);
nor U31270 (N_31270,N_29374,N_28858);
nor U31271 (N_31271,N_29954,N_27895);
or U31272 (N_31272,N_27643,N_29963);
or U31273 (N_31273,N_29711,N_29609);
nor U31274 (N_31274,N_28561,N_28015);
nor U31275 (N_31275,N_29843,N_29525);
nand U31276 (N_31276,N_28821,N_28280);
xor U31277 (N_31277,N_29537,N_28495);
nor U31278 (N_31278,N_28952,N_29933);
and U31279 (N_31279,N_28995,N_29038);
nor U31280 (N_31280,N_28671,N_29961);
xor U31281 (N_31281,N_28885,N_28432);
xor U31282 (N_31282,N_28178,N_28852);
and U31283 (N_31283,N_29608,N_29612);
xnor U31284 (N_31284,N_28907,N_28804);
nor U31285 (N_31285,N_28244,N_29622);
nand U31286 (N_31286,N_27548,N_29757);
and U31287 (N_31287,N_28742,N_28307);
and U31288 (N_31288,N_29935,N_27505);
xor U31289 (N_31289,N_28737,N_29279);
or U31290 (N_31290,N_29129,N_29211);
nor U31291 (N_31291,N_27607,N_27903);
and U31292 (N_31292,N_29679,N_29042);
nand U31293 (N_31293,N_28537,N_27689);
xor U31294 (N_31294,N_28010,N_29837);
and U31295 (N_31295,N_29784,N_28474);
nor U31296 (N_31296,N_28049,N_27831);
nand U31297 (N_31297,N_28316,N_29193);
or U31298 (N_31298,N_27898,N_27799);
nor U31299 (N_31299,N_28989,N_29821);
nor U31300 (N_31300,N_29557,N_29103);
or U31301 (N_31301,N_28944,N_29744);
xor U31302 (N_31302,N_29201,N_29872);
or U31303 (N_31303,N_28126,N_27933);
xnor U31304 (N_31304,N_27797,N_29005);
or U31305 (N_31305,N_28904,N_29098);
xnor U31306 (N_31306,N_29293,N_27543);
nor U31307 (N_31307,N_28804,N_28732);
nand U31308 (N_31308,N_27729,N_28453);
nand U31309 (N_31309,N_28510,N_28223);
nor U31310 (N_31310,N_29695,N_28546);
or U31311 (N_31311,N_29904,N_28045);
xor U31312 (N_31312,N_29491,N_28409);
xnor U31313 (N_31313,N_28555,N_27837);
xor U31314 (N_31314,N_28034,N_29820);
and U31315 (N_31315,N_28835,N_28467);
nor U31316 (N_31316,N_29415,N_28682);
nor U31317 (N_31317,N_28910,N_29581);
and U31318 (N_31318,N_29148,N_29469);
and U31319 (N_31319,N_29168,N_28917);
or U31320 (N_31320,N_28949,N_28745);
or U31321 (N_31321,N_27630,N_27520);
nor U31322 (N_31322,N_28409,N_27560);
or U31323 (N_31323,N_27634,N_28295);
nand U31324 (N_31324,N_28458,N_28640);
or U31325 (N_31325,N_29497,N_28558);
and U31326 (N_31326,N_29289,N_29901);
and U31327 (N_31327,N_28955,N_27687);
and U31328 (N_31328,N_27726,N_27532);
nor U31329 (N_31329,N_29013,N_27510);
xnor U31330 (N_31330,N_28937,N_28835);
nor U31331 (N_31331,N_29160,N_28360);
or U31332 (N_31332,N_27653,N_29578);
and U31333 (N_31333,N_29606,N_29268);
xor U31334 (N_31334,N_27955,N_29481);
nand U31335 (N_31335,N_28842,N_29680);
nor U31336 (N_31336,N_29922,N_27654);
xor U31337 (N_31337,N_29631,N_28865);
and U31338 (N_31338,N_28448,N_28724);
nand U31339 (N_31339,N_29254,N_27775);
or U31340 (N_31340,N_29547,N_27826);
nor U31341 (N_31341,N_28476,N_27941);
or U31342 (N_31342,N_28152,N_29775);
xor U31343 (N_31343,N_28259,N_28647);
nand U31344 (N_31344,N_29744,N_28581);
or U31345 (N_31345,N_28481,N_29012);
nand U31346 (N_31346,N_28087,N_29890);
xor U31347 (N_31347,N_29437,N_29866);
nor U31348 (N_31348,N_27534,N_28425);
and U31349 (N_31349,N_29017,N_28102);
nor U31350 (N_31350,N_29655,N_29173);
nor U31351 (N_31351,N_29454,N_28854);
nor U31352 (N_31352,N_29675,N_29667);
nand U31353 (N_31353,N_29418,N_27903);
nand U31354 (N_31354,N_29079,N_27985);
xnor U31355 (N_31355,N_29542,N_29438);
xnor U31356 (N_31356,N_28417,N_29545);
or U31357 (N_31357,N_29925,N_29040);
nor U31358 (N_31358,N_29574,N_27743);
nand U31359 (N_31359,N_28840,N_28356);
and U31360 (N_31360,N_29607,N_29802);
and U31361 (N_31361,N_27526,N_28332);
xnor U31362 (N_31362,N_28899,N_28700);
and U31363 (N_31363,N_28735,N_28410);
and U31364 (N_31364,N_28830,N_29295);
or U31365 (N_31365,N_27830,N_29137);
nor U31366 (N_31366,N_29237,N_27666);
or U31367 (N_31367,N_29766,N_28538);
nor U31368 (N_31368,N_29175,N_29414);
and U31369 (N_31369,N_29404,N_27943);
xor U31370 (N_31370,N_27955,N_27684);
xor U31371 (N_31371,N_27978,N_28717);
nor U31372 (N_31372,N_28436,N_28420);
xor U31373 (N_31373,N_28227,N_28729);
and U31374 (N_31374,N_28619,N_29232);
or U31375 (N_31375,N_29281,N_28659);
nor U31376 (N_31376,N_29282,N_28240);
nor U31377 (N_31377,N_29995,N_29871);
xor U31378 (N_31378,N_28595,N_28874);
nand U31379 (N_31379,N_28256,N_28493);
or U31380 (N_31380,N_29709,N_29673);
nor U31381 (N_31381,N_27936,N_28161);
nand U31382 (N_31382,N_28722,N_29813);
or U31383 (N_31383,N_29662,N_28417);
or U31384 (N_31384,N_28717,N_29661);
xor U31385 (N_31385,N_28154,N_29859);
nand U31386 (N_31386,N_29409,N_29976);
and U31387 (N_31387,N_29965,N_29399);
nor U31388 (N_31388,N_29728,N_28105);
and U31389 (N_31389,N_29351,N_28751);
and U31390 (N_31390,N_29795,N_28969);
and U31391 (N_31391,N_27559,N_29994);
nand U31392 (N_31392,N_28347,N_27571);
or U31393 (N_31393,N_27557,N_28974);
and U31394 (N_31394,N_29771,N_28808);
xor U31395 (N_31395,N_29275,N_27510);
nand U31396 (N_31396,N_28559,N_28425);
or U31397 (N_31397,N_28846,N_27943);
nand U31398 (N_31398,N_29992,N_29399);
xnor U31399 (N_31399,N_29142,N_27579);
and U31400 (N_31400,N_28046,N_28154);
nand U31401 (N_31401,N_28910,N_29266);
nand U31402 (N_31402,N_28833,N_28474);
and U31403 (N_31403,N_27821,N_29888);
nand U31404 (N_31404,N_29547,N_28031);
nand U31405 (N_31405,N_27593,N_28250);
or U31406 (N_31406,N_28731,N_29187);
nand U31407 (N_31407,N_29555,N_27587);
nor U31408 (N_31408,N_27537,N_29537);
or U31409 (N_31409,N_29316,N_29834);
nor U31410 (N_31410,N_28870,N_29729);
xor U31411 (N_31411,N_28988,N_29503);
nand U31412 (N_31412,N_27575,N_27591);
nor U31413 (N_31413,N_27912,N_29531);
or U31414 (N_31414,N_29011,N_29942);
and U31415 (N_31415,N_29653,N_29736);
and U31416 (N_31416,N_29597,N_27526);
xor U31417 (N_31417,N_28257,N_28263);
xor U31418 (N_31418,N_27791,N_29498);
xor U31419 (N_31419,N_28695,N_27667);
or U31420 (N_31420,N_29966,N_28935);
xor U31421 (N_31421,N_28440,N_27886);
or U31422 (N_31422,N_28492,N_28884);
nor U31423 (N_31423,N_28908,N_28378);
nor U31424 (N_31424,N_28678,N_28263);
or U31425 (N_31425,N_28448,N_29645);
nand U31426 (N_31426,N_27569,N_28993);
and U31427 (N_31427,N_29420,N_27966);
nand U31428 (N_31428,N_29424,N_29037);
or U31429 (N_31429,N_28276,N_28630);
or U31430 (N_31430,N_27932,N_27568);
and U31431 (N_31431,N_28164,N_29774);
xor U31432 (N_31432,N_27983,N_27787);
or U31433 (N_31433,N_28123,N_28830);
or U31434 (N_31434,N_29556,N_28935);
xor U31435 (N_31435,N_29948,N_29847);
xnor U31436 (N_31436,N_28619,N_28560);
or U31437 (N_31437,N_28574,N_27931);
xor U31438 (N_31438,N_27608,N_27556);
nand U31439 (N_31439,N_28286,N_29288);
nor U31440 (N_31440,N_27832,N_29613);
and U31441 (N_31441,N_29538,N_28178);
or U31442 (N_31442,N_28384,N_27980);
or U31443 (N_31443,N_28155,N_27565);
and U31444 (N_31444,N_27597,N_28424);
xor U31445 (N_31445,N_29464,N_29985);
nor U31446 (N_31446,N_28151,N_28082);
or U31447 (N_31447,N_28771,N_29010);
or U31448 (N_31448,N_29783,N_27975);
xor U31449 (N_31449,N_29743,N_27586);
nand U31450 (N_31450,N_29142,N_28998);
nor U31451 (N_31451,N_29390,N_28363);
and U31452 (N_31452,N_28767,N_29449);
or U31453 (N_31453,N_29289,N_28743);
xor U31454 (N_31454,N_28871,N_27501);
xor U31455 (N_31455,N_28600,N_27584);
xnor U31456 (N_31456,N_29267,N_29791);
or U31457 (N_31457,N_28952,N_29243);
nand U31458 (N_31458,N_29419,N_29412);
nor U31459 (N_31459,N_28654,N_28026);
and U31460 (N_31460,N_28825,N_28142);
nor U31461 (N_31461,N_29316,N_29758);
nand U31462 (N_31462,N_29634,N_28897);
or U31463 (N_31463,N_27520,N_29741);
xnor U31464 (N_31464,N_29501,N_28624);
and U31465 (N_31465,N_29856,N_27931);
or U31466 (N_31466,N_28209,N_27947);
nand U31467 (N_31467,N_29249,N_29630);
nor U31468 (N_31468,N_28065,N_28279);
nor U31469 (N_31469,N_29274,N_29497);
nor U31470 (N_31470,N_28744,N_28501);
nand U31471 (N_31471,N_29482,N_28235);
or U31472 (N_31472,N_29701,N_28601);
nor U31473 (N_31473,N_27678,N_28800);
and U31474 (N_31474,N_29157,N_27915);
xor U31475 (N_31475,N_28632,N_28394);
and U31476 (N_31476,N_28419,N_29151);
or U31477 (N_31477,N_27678,N_27746);
and U31478 (N_31478,N_29707,N_28707);
xor U31479 (N_31479,N_28485,N_29716);
nand U31480 (N_31480,N_27574,N_28412);
nor U31481 (N_31481,N_29271,N_28387);
nor U31482 (N_31482,N_29778,N_28085);
nor U31483 (N_31483,N_29331,N_28970);
nor U31484 (N_31484,N_28876,N_28518);
nor U31485 (N_31485,N_28363,N_29579);
or U31486 (N_31486,N_28406,N_29031);
and U31487 (N_31487,N_28214,N_29140);
nor U31488 (N_31488,N_29884,N_27832);
or U31489 (N_31489,N_28780,N_28534);
or U31490 (N_31490,N_29929,N_28328);
or U31491 (N_31491,N_29936,N_29010);
xor U31492 (N_31492,N_29628,N_29616);
nor U31493 (N_31493,N_29328,N_29021);
nor U31494 (N_31494,N_29130,N_27754);
nor U31495 (N_31495,N_28045,N_28679);
or U31496 (N_31496,N_28961,N_27650);
xor U31497 (N_31497,N_29366,N_29961);
and U31498 (N_31498,N_29332,N_28878);
nand U31499 (N_31499,N_29559,N_29143);
xor U31500 (N_31500,N_28199,N_27532);
nor U31501 (N_31501,N_28141,N_27690);
and U31502 (N_31502,N_28729,N_27786);
nand U31503 (N_31503,N_28781,N_28410);
nor U31504 (N_31504,N_28715,N_28401);
nand U31505 (N_31505,N_27917,N_29731);
nor U31506 (N_31506,N_27889,N_28411);
or U31507 (N_31507,N_29057,N_28561);
nand U31508 (N_31508,N_28807,N_29454);
or U31509 (N_31509,N_29227,N_27846);
nand U31510 (N_31510,N_28439,N_29441);
nand U31511 (N_31511,N_29478,N_27523);
nand U31512 (N_31512,N_28380,N_28481);
nor U31513 (N_31513,N_27625,N_29820);
or U31514 (N_31514,N_27745,N_28155);
nor U31515 (N_31515,N_29099,N_28549);
nand U31516 (N_31516,N_29480,N_28957);
nand U31517 (N_31517,N_29741,N_29079);
nor U31518 (N_31518,N_28353,N_29805);
xor U31519 (N_31519,N_28748,N_29092);
and U31520 (N_31520,N_29915,N_29545);
and U31521 (N_31521,N_29849,N_28927);
or U31522 (N_31522,N_28677,N_29127);
xnor U31523 (N_31523,N_27814,N_29417);
nor U31524 (N_31524,N_28210,N_28844);
nor U31525 (N_31525,N_28193,N_28760);
or U31526 (N_31526,N_29268,N_27920);
and U31527 (N_31527,N_28462,N_27914);
xor U31528 (N_31528,N_28873,N_29915);
nor U31529 (N_31529,N_29189,N_29877);
nand U31530 (N_31530,N_28826,N_29192);
xor U31531 (N_31531,N_29662,N_28341);
or U31532 (N_31532,N_27547,N_27965);
nor U31533 (N_31533,N_28100,N_29675);
nand U31534 (N_31534,N_29967,N_29931);
nand U31535 (N_31535,N_28104,N_29177);
nand U31536 (N_31536,N_27830,N_28466);
and U31537 (N_31537,N_28406,N_27984);
and U31538 (N_31538,N_27983,N_28892);
nand U31539 (N_31539,N_27627,N_29705);
and U31540 (N_31540,N_28574,N_28757);
xor U31541 (N_31541,N_29620,N_28802);
nor U31542 (N_31542,N_28289,N_29655);
and U31543 (N_31543,N_28776,N_28964);
nor U31544 (N_31544,N_29466,N_28516);
nand U31545 (N_31545,N_27603,N_28979);
and U31546 (N_31546,N_28114,N_29858);
nor U31547 (N_31547,N_27622,N_29367);
or U31548 (N_31548,N_27580,N_28637);
or U31549 (N_31549,N_29851,N_29026);
nor U31550 (N_31550,N_29682,N_29904);
nand U31551 (N_31551,N_28730,N_28573);
or U31552 (N_31552,N_28494,N_29746);
or U31553 (N_31553,N_28856,N_28590);
nand U31554 (N_31554,N_29532,N_28723);
nand U31555 (N_31555,N_27688,N_28150);
nand U31556 (N_31556,N_28672,N_28239);
xor U31557 (N_31557,N_27678,N_29360);
or U31558 (N_31558,N_28924,N_28572);
and U31559 (N_31559,N_28486,N_27917);
and U31560 (N_31560,N_28871,N_27527);
xnor U31561 (N_31561,N_28791,N_27694);
or U31562 (N_31562,N_27574,N_29828);
xnor U31563 (N_31563,N_29646,N_28472);
nand U31564 (N_31564,N_27889,N_28807);
nor U31565 (N_31565,N_27529,N_28833);
or U31566 (N_31566,N_29260,N_28906);
and U31567 (N_31567,N_29733,N_29152);
or U31568 (N_31568,N_28227,N_27551);
or U31569 (N_31569,N_29852,N_27832);
and U31570 (N_31570,N_29819,N_29964);
and U31571 (N_31571,N_27931,N_29112);
nor U31572 (N_31572,N_28827,N_29528);
or U31573 (N_31573,N_29744,N_29421);
nand U31574 (N_31574,N_29382,N_29227);
nor U31575 (N_31575,N_28320,N_28890);
or U31576 (N_31576,N_27917,N_29216);
or U31577 (N_31577,N_28661,N_28758);
or U31578 (N_31578,N_28893,N_29719);
nand U31579 (N_31579,N_29359,N_29898);
or U31580 (N_31580,N_28586,N_28292);
nor U31581 (N_31581,N_27797,N_29988);
xnor U31582 (N_31582,N_27888,N_27605);
or U31583 (N_31583,N_29197,N_27626);
and U31584 (N_31584,N_28207,N_27513);
or U31585 (N_31585,N_27506,N_29523);
nand U31586 (N_31586,N_28772,N_28479);
and U31587 (N_31587,N_27816,N_28765);
nand U31588 (N_31588,N_27849,N_28550);
nand U31589 (N_31589,N_28858,N_29660);
or U31590 (N_31590,N_28937,N_29132);
or U31591 (N_31591,N_28125,N_28929);
or U31592 (N_31592,N_28101,N_27766);
or U31593 (N_31593,N_29661,N_27803);
or U31594 (N_31594,N_29834,N_29151);
and U31595 (N_31595,N_28384,N_28843);
and U31596 (N_31596,N_28339,N_27627);
nor U31597 (N_31597,N_27537,N_28630);
and U31598 (N_31598,N_28566,N_28304);
or U31599 (N_31599,N_28626,N_27974);
nand U31600 (N_31600,N_28083,N_27982);
xnor U31601 (N_31601,N_28722,N_29484);
and U31602 (N_31602,N_29032,N_29921);
nor U31603 (N_31603,N_28274,N_29458);
nor U31604 (N_31604,N_28721,N_29664);
nor U31605 (N_31605,N_27884,N_29100);
and U31606 (N_31606,N_29792,N_28257);
nor U31607 (N_31607,N_29950,N_28641);
nand U31608 (N_31608,N_29544,N_28389);
nand U31609 (N_31609,N_28100,N_28818);
and U31610 (N_31610,N_29821,N_28699);
nand U31611 (N_31611,N_28455,N_28174);
nor U31612 (N_31612,N_29835,N_28451);
or U31613 (N_31613,N_28930,N_29105);
and U31614 (N_31614,N_28653,N_28003);
xor U31615 (N_31615,N_28096,N_29130);
or U31616 (N_31616,N_29541,N_27729);
xnor U31617 (N_31617,N_29214,N_28178);
nor U31618 (N_31618,N_27750,N_29772);
and U31619 (N_31619,N_29255,N_28843);
xor U31620 (N_31620,N_29536,N_28470);
or U31621 (N_31621,N_28859,N_29780);
nor U31622 (N_31622,N_29600,N_27892);
or U31623 (N_31623,N_27674,N_28801);
xor U31624 (N_31624,N_28972,N_29766);
nor U31625 (N_31625,N_29043,N_28313);
nor U31626 (N_31626,N_27581,N_28455);
and U31627 (N_31627,N_29820,N_27503);
or U31628 (N_31628,N_28339,N_28467);
nor U31629 (N_31629,N_29327,N_29770);
xnor U31630 (N_31630,N_29011,N_28421);
nor U31631 (N_31631,N_29806,N_29397);
xnor U31632 (N_31632,N_29649,N_29467);
and U31633 (N_31633,N_27897,N_27621);
or U31634 (N_31634,N_27786,N_28575);
nor U31635 (N_31635,N_29552,N_28594);
and U31636 (N_31636,N_28929,N_27965);
and U31637 (N_31637,N_28916,N_29007);
nor U31638 (N_31638,N_29270,N_29701);
and U31639 (N_31639,N_27683,N_28921);
nand U31640 (N_31640,N_29879,N_27782);
nor U31641 (N_31641,N_29816,N_27990);
or U31642 (N_31642,N_28252,N_28439);
or U31643 (N_31643,N_29415,N_28083);
or U31644 (N_31644,N_28938,N_29432);
and U31645 (N_31645,N_27725,N_29614);
xnor U31646 (N_31646,N_28428,N_28237);
nor U31647 (N_31647,N_28529,N_28202);
or U31648 (N_31648,N_27906,N_27902);
or U31649 (N_31649,N_29297,N_29356);
or U31650 (N_31650,N_29915,N_28535);
xor U31651 (N_31651,N_29600,N_29625);
nor U31652 (N_31652,N_27669,N_27788);
xor U31653 (N_31653,N_27612,N_27589);
or U31654 (N_31654,N_27616,N_29449);
nand U31655 (N_31655,N_29116,N_29179);
nand U31656 (N_31656,N_27702,N_29768);
or U31657 (N_31657,N_28196,N_27570);
nor U31658 (N_31658,N_27937,N_28124);
and U31659 (N_31659,N_28852,N_28359);
or U31660 (N_31660,N_29962,N_27916);
and U31661 (N_31661,N_28028,N_29565);
and U31662 (N_31662,N_27869,N_29868);
nor U31663 (N_31663,N_28742,N_28788);
or U31664 (N_31664,N_28571,N_29701);
xor U31665 (N_31665,N_28350,N_29355);
nor U31666 (N_31666,N_28975,N_27922);
or U31667 (N_31667,N_28722,N_27829);
and U31668 (N_31668,N_27669,N_28204);
xnor U31669 (N_31669,N_29017,N_29952);
and U31670 (N_31670,N_29465,N_28995);
or U31671 (N_31671,N_28604,N_29254);
nand U31672 (N_31672,N_28394,N_28320);
and U31673 (N_31673,N_28318,N_28726);
nand U31674 (N_31674,N_29521,N_28113);
nand U31675 (N_31675,N_28035,N_28177);
and U31676 (N_31676,N_28641,N_28513);
or U31677 (N_31677,N_27883,N_28780);
nand U31678 (N_31678,N_28028,N_29771);
nor U31679 (N_31679,N_28966,N_28499);
or U31680 (N_31680,N_28231,N_28815);
xor U31681 (N_31681,N_29691,N_27718);
xor U31682 (N_31682,N_28643,N_28504);
xor U31683 (N_31683,N_29952,N_29091);
nand U31684 (N_31684,N_29184,N_28699);
nand U31685 (N_31685,N_27817,N_29861);
xnor U31686 (N_31686,N_28580,N_27917);
nand U31687 (N_31687,N_29521,N_28860);
xor U31688 (N_31688,N_28898,N_29105);
nor U31689 (N_31689,N_28751,N_28293);
nand U31690 (N_31690,N_28957,N_29088);
or U31691 (N_31691,N_28270,N_29534);
xnor U31692 (N_31692,N_27794,N_28504);
xor U31693 (N_31693,N_27796,N_29784);
xor U31694 (N_31694,N_27644,N_27972);
nor U31695 (N_31695,N_27598,N_29873);
xor U31696 (N_31696,N_27698,N_29795);
xnor U31697 (N_31697,N_27776,N_27894);
nor U31698 (N_31698,N_28290,N_29615);
and U31699 (N_31699,N_28424,N_28622);
xnor U31700 (N_31700,N_27682,N_28675);
nor U31701 (N_31701,N_28032,N_29031);
xnor U31702 (N_31702,N_27635,N_28777);
xor U31703 (N_31703,N_27713,N_27966);
xor U31704 (N_31704,N_28957,N_29463);
nand U31705 (N_31705,N_28508,N_28498);
nor U31706 (N_31706,N_28951,N_27851);
xnor U31707 (N_31707,N_29066,N_27572);
or U31708 (N_31708,N_27673,N_28488);
nand U31709 (N_31709,N_27605,N_28992);
xor U31710 (N_31710,N_29848,N_27814);
nor U31711 (N_31711,N_28266,N_28922);
xnor U31712 (N_31712,N_27956,N_28586);
nor U31713 (N_31713,N_27601,N_29257);
or U31714 (N_31714,N_28631,N_29291);
nand U31715 (N_31715,N_28457,N_28674);
and U31716 (N_31716,N_29533,N_29617);
and U31717 (N_31717,N_27581,N_29181);
nand U31718 (N_31718,N_27739,N_29346);
or U31719 (N_31719,N_27928,N_29609);
xnor U31720 (N_31720,N_28739,N_29721);
xor U31721 (N_31721,N_28113,N_29075);
and U31722 (N_31722,N_29788,N_28146);
nand U31723 (N_31723,N_27748,N_28822);
nand U31724 (N_31724,N_29739,N_28801);
xor U31725 (N_31725,N_29001,N_28000);
xnor U31726 (N_31726,N_27797,N_28780);
or U31727 (N_31727,N_29691,N_27797);
xor U31728 (N_31728,N_29689,N_29470);
xnor U31729 (N_31729,N_27509,N_28740);
and U31730 (N_31730,N_28293,N_27943);
nand U31731 (N_31731,N_27774,N_28067);
nand U31732 (N_31732,N_28510,N_29079);
nor U31733 (N_31733,N_27898,N_28300);
and U31734 (N_31734,N_29121,N_27878);
nand U31735 (N_31735,N_28380,N_29195);
xor U31736 (N_31736,N_29989,N_28762);
or U31737 (N_31737,N_29491,N_28148);
xor U31738 (N_31738,N_29869,N_29807);
xnor U31739 (N_31739,N_29766,N_29298);
and U31740 (N_31740,N_29370,N_29558);
xnor U31741 (N_31741,N_27869,N_28884);
and U31742 (N_31742,N_28772,N_28429);
nand U31743 (N_31743,N_29181,N_28279);
nor U31744 (N_31744,N_28626,N_29982);
and U31745 (N_31745,N_29054,N_28651);
and U31746 (N_31746,N_29525,N_28306);
nand U31747 (N_31747,N_29106,N_29975);
and U31748 (N_31748,N_28848,N_29845);
xnor U31749 (N_31749,N_28029,N_29566);
and U31750 (N_31750,N_29060,N_28379);
nand U31751 (N_31751,N_29361,N_29310);
nor U31752 (N_31752,N_29651,N_27596);
and U31753 (N_31753,N_28113,N_29686);
nor U31754 (N_31754,N_28689,N_28100);
and U31755 (N_31755,N_27875,N_27821);
and U31756 (N_31756,N_29321,N_28178);
nor U31757 (N_31757,N_28700,N_27610);
and U31758 (N_31758,N_29399,N_28203);
xnor U31759 (N_31759,N_29340,N_29601);
xnor U31760 (N_31760,N_28682,N_29428);
nand U31761 (N_31761,N_28987,N_28545);
xor U31762 (N_31762,N_29834,N_28130);
xnor U31763 (N_31763,N_28444,N_29470);
nand U31764 (N_31764,N_29362,N_28486);
or U31765 (N_31765,N_29877,N_28469);
xor U31766 (N_31766,N_29385,N_28328);
and U31767 (N_31767,N_28397,N_27757);
and U31768 (N_31768,N_27584,N_28479);
nand U31769 (N_31769,N_28874,N_28951);
and U31770 (N_31770,N_29919,N_29972);
nor U31771 (N_31771,N_29178,N_29155);
or U31772 (N_31772,N_27703,N_27594);
nand U31773 (N_31773,N_29323,N_29166);
nand U31774 (N_31774,N_27654,N_27915);
or U31775 (N_31775,N_28214,N_29149);
and U31776 (N_31776,N_28945,N_28937);
nor U31777 (N_31777,N_29617,N_29994);
nand U31778 (N_31778,N_27769,N_29749);
or U31779 (N_31779,N_28339,N_29333);
and U31780 (N_31780,N_29210,N_27863);
xnor U31781 (N_31781,N_28736,N_29374);
xor U31782 (N_31782,N_27823,N_27838);
or U31783 (N_31783,N_28671,N_29000);
and U31784 (N_31784,N_27513,N_28432);
or U31785 (N_31785,N_28380,N_29626);
nand U31786 (N_31786,N_29902,N_29512);
or U31787 (N_31787,N_28546,N_29859);
or U31788 (N_31788,N_29352,N_27810);
xor U31789 (N_31789,N_29676,N_28327);
xor U31790 (N_31790,N_29346,N_27843);
nor U31791 (N_31791,N_28395,N_29007);
xnor U31792 (N_31792,N_29243,N_28869);
nor U31793 (N_31793,N_27889,N_29528);
and U31794 (N_31794,N_29278,N_28363);
and U31795 (N_31795,N_27929,N_28775);
nand U31796 (N_31796,N_28318,N_29109);
or U31797 (N_31797,N_29264,N_29936);
nor U31798 (N_31798,N_28694,N_29064);
xor U31799 (N_31799,N_27800,N_29460);
and U31800 (N_31800,N_28967,N_29597);
or U31801 (N_31801,N_29101,N_28071);
xnor U31802 (N_31802,N_28265,N_28766);
nand U31803 (N_31803,N_28720,N_28401);
or U31804 (N_31804,N_29601,N_28881);
nor U31805 (N_31805,N_29613,N_28909);
xnor U31806 (N_31806,N_29437,N_28916);
and U31807 (N_31807,N_28216,N_28394);
nand U31808 (N_31808,N_28999,N_28364);
and U31809 (N_31809,N_29795,N_28792);
or U31810 (N_31810,N_28383,N_29801);
xnor U31811 (N_31811,N_27593,N_29907);
nor U31812 (N_31812,N_27885,N_28734);
xor U31813 (N_31813,N_28044,N_27565);
xnor U31814 (N_31814,N_28093,N_28508);
or U31815 (N_31815,N_28840,N_28691);
or U31816 (N_31816,N_27701,N_28786);
nor U31817 (N_31817,N_28689,N_29503);
or U31818 (N_31818,N_27795,N_28937);
nand U31819 (N_31819,N_29414,N_27923);
or U31820 (N_31820,N_28509,N_27995);
nor U31821 (N_31821,N_28089,N_27693);
xor U31822 (N_31822,N_29281,N_28429);
xor U31823 (N_31823,N_27748,N_27612);
nor U31824 (N_31824,N_28985,N_29549);
nor U31825 (N_31825,N_27814,N_29440);
or U31826 (N_31826,N_29055,N_29941);
or U31827 (N_31827,N_27527,N_29846);
and U31828 (N_31828,N_29997,N_29937);
nand U31829 (N_31829,N_28124,N_29934);
and U31830 (N_31830,N_27677,N_27765);
nand U31831 (N_31831,N_29813,N_29207);
nand U31832 (N_31832,N_28815,N_28461);
and U31833 (N_31833,N_29750,N_29305);
or U31834 (N_31834,N_27827,N_29773);
and U31835 (N_31835,N_28211,N_27685);
nand U31836 (N_31836,N_28872,N_29717);
or U31837 (N_31837,N_27565,N_27554);
xnor U31838 (N_31838,N_29627,N_29044);
or U31839 (N_31839,N_28943,N_29846);
and U31840 (N_31840,N_29459,N_28737);
xor U31841 (N_31841,N_28938,N_28075);
nor U31842 (N_31842,N_29180,N_29628);
nand U31843 (N_31843,N_29452,N_28515);
or U31844 (N_31844,N_29616,N_28222);
nand U31845 (N_31845,N_28860,N_29803);
nand U31846 (N_31846,N_27534,N_29835);
or U31847 (N_31847,N_27901,N_29167);
nor U31848 (N_31848,N_28522,N_28406);
xnor U31849 (N_31849,N_28087,N_28218);
or U31850 (N_31850,N_29728,N_27887);
nand U31851 (N_31851,N_27571,N_29816);
xnor U31852 (N_31852,N_29538,N_28206);
xor U31853 (N_31853,N_29205,N_29838);
nand U31854 (N_31854,N_28027,N_27534);
and U31855 (N_31855,N_28391,N_28565);
or U31856 (N_31856,N_27613,N_28231);
nor U31857 (N_31857,N_28405,N_29774);
nand U31858 (N_31858,N_29589,N_27502);
and U31859 (N_31859,N_27862,N_28779);
nand U31860 (N_31860,N_27944,N_29807);
or U31861 (N_31861,N_27810,N_29577);
xor U31862 (N_31862,N_27709,N_29186);
nor U31863 (N_31863,N_28170,N_27538);
and U31864 (N_31864,N_29546,N_28105);
nor U31865 (N_31865,N_29713,N_29417);
xor U31866 (N_31866,N_28391,N_29460);
and U31867 (N_31867,N_29245,N_27971);
nand U31868 (N_31868,N_27744,N_29354);
and U31869 (N_31869,N_28948,N_28664);
nor U31870 (N_31870,N_27607,N_28207);
or U31871 (N_31871,N_29362,N_29931);
and U31872 (N_31872,N_29412,N_28706);
nor U31873 (N_31873,N_28799,N_28764);
nor U31874 (N_31874,N_28774,N_29443);
xnor U31875 (N_31875,N_27992,N_27926);
or U31876 (N_31876,N_28752,N_28772);
and U31877 (N_31877,N_27998,N_28590);
and U31878 (N_31878,N_28880,N_28685);
and U31879 (N_31879,N_29317,N_29100);
nand U31880 (N_31880,N_29495,N_28099);
or U31881 (N_31881,N_29155,N_27914);
and U31882 (N_31882,N_29975,N_28077);
nand U31883 (N_31883,N_29687,N_27667);
or U31884 (N_31884,N_28711,N_29073);
nand U31885 (N_31885,N_29699,N_27908);
xor U31886 (N_31886,N_28433,N_28823);
xor U31887 (N_31887,N_27774,N_29044);
xor U31888 (N_31888,N_28880,N_29286);
and U31889 (N_31889,N_29790,N_29107);
nand U31890 (N_31890,N_28553,N_29329);
or U31891 (N_31891,N_28732,N_29715);
nand U31892 (N_31892,N_28287,N_29169);
or U31893 (N_31893,N_29392,N_27558);
and U31894 (N_31894,N_28458,N_28080);
and U31895 (N_31895,N_28515,N_29150);
nand U31896 (N_31896,N_28384,N_28550);
and U31897 (N_31897,N_29856,N_28069);
nor U31898 (N_31898,N_29281,N_27863);
nor U31899 (N_31899,N_28715,N_28411);
or U31900 (N_31900,N_28396,N_28437);
nor U31901 (N_31901,N_28797,N_28822);
nor U31902 (N_31902,N_29160,N_28931);
or U31903 (N_31903,N_29747,N_29954);
and U31904 (N_31904,N_29950,N_29584);
and U31905 (N_31905,N_28869,N_29283);
or U31906 (N_31906,N_28328,N_29009);
nand U31907 (N_31907,N_28999,N_28512);
nand U31908 (N_31908,N_29628,N_29348);
and U31909 (N_31909,N_29001,N_28942);
nand U31910 (N_31910,N_27643,N_27799);
nor U31911 (N_31911,N_28617,N_29773);
nor U31912 (N_31912,N_29466,N_29170);
xor U31913 (N_31913,N_27791,N_28546);
nor U31914 (N_31914,N_28376,N_28830);
xnor U31915 (N_31915,N_29777,N_29796);
or U31916 (N_31916,N_29066,N_29704);
and U31917 (N_31917,N_29521,N_29131);
or U31918 (N_31918,N_27822,N_28290);
or U31919 (N_31919,N_28202,N_27968);
nor U31920 (N_31920,N_29223,N_29624);
or U31921 (N_31921,N_28642,N_27975);
or U31922 (N_31922,N_28217,N_29338);
nor U31923 (N_31923,N_29171,N_28979);
and U31924 (N_31924,N_28837,N_29989);
xor U31925 (N_31925,N_27887,N_27814);
nor U31926 (N_31926,N_28758,N_28510);
nor U31927 (N_31927,N_29797,N_29209);
nand U31928 (N_31928,N_29999,N_27934);
xor U31929 (N_31929,N_28671,N_28159);
xor U31930 (N_31930,N_29351,N_29311);
xor U31931 (N_31931,N_27997,N_27902);
xor U31932 (N_31932,N_27538,N_27649);
or U31933 (N_31933,N_29196,N_29014);
nand U31934 (N_31934,N_29015,N_28054);
xor U31935 (N_31935,N_29909,N_29960);
or U31936 (N_31936,N_27635,N_29939);
xnor U31937 (N_31937,N_28524,N_28098);
or U31938 (N_31938,N_28411,N_27945);
nor U31939 (N_31939,N_29770,N_27568);
nand U31940 (N_31940,N_27881,N_29700);
nand U31941 (N_31941,N_27571,N_29613);
nor U31942 (N_31942,N_29967,N_27960);
xnor U31943 (N_31943,N_28258,N_29391);
nor U31944 (N_31944,N_27992,N_29624);
nor U31945 (N_31945,N_27666,N_28671);
nand U31946 (N_31946,N_28895,N_28656);
and U31947 (N_31947,N_27656,N_28000);
nor U31948 (N_31948,N_29398,N_28877);
and U31949 (N_31949,N_29304,N_28214);
nor U31950 (N_31950,N_29783,N_28023);
nand U31951 (N_31951,N_29926,N_27805);
nand U31952 (N_31952,N_29979,N_27501);
and U31953 (N_31953,N_28287,N_28323);
xnor U31954 (N_31954,N_27647,N_29334);
or U31955 (N_31955,N_28369,N_28309);
nand U31956 (N_31956,N_28243,N_29141);
and U31957 (N_31957,N_29335,N_28452);
or U31958 (N_31958,N_29413,N_29513);
nand U31959 (N_31959,N_29662,N_29205);
xnor U31960 (N_31960,N_27798,N_27765);
or U31961 (N_31961,N_29875,N_27513);
and U31962 (N_31962,N_28864,N_28225);
xnor U31963 (N_31963,N_27979,N_29767);
nand U31964 (N_31964,N_28095,N_28114);
nor U31965 (N_31965,N_28783,N_29713);
nand U31966 (N_31966,N_29689,N_28407);
and U31967 (N_31967,N_29912,N_29951);
and U31968 (N_31968,N_29822,N_28631);
or U31969 (N_31969,N_28817,N_29306);
or U31970 (N_31970,N_28163,N_28521);
nand U31971 (N_31971,N_28019,N_28250);
nor U31972 (N_31972,N_29682,N_27703);
nor U31973 (N_31973,N_27821,N_28810);
nor U31974 (N_31974,N_27942,N_27644);
nand U31975 (N_31975,N_29218,N_27572);
nor U31976 (N_31976,N_28462,N_29738);
and U31977 (N_31977,N_29138,N_28866);
and U31978 (N_31978,N_28415,N_27694);
or U31979 (N_31979,N_29264,N_28994);
xor U31980 (N_31980,N_28349,N_29685);
xor U31981 (N_31981,N_27888,N_29092);
xnor U31982 (N_31982,N_29880,N_27634);
xnor U31983 (N_31983,N_29815,N_27504);
or U31984 (N_31984,N_28844,N_27644);
xnor U31985 (N_31985,N_29897,N_27849);
xor U31986 (N_31986,N_28565,N_28170);
xnor U31987 (N_31987,N_28627,N_28030);
or U31988 (N_31988,N_27640,N_29579);
and U31989 (N_31989,N_29015,N_29779);
and U31990 (N_31990,N_28166,N_27709);
xor U31991 (N_31991,N_28235,N_28994);
xnor U31992 (N_31992,N_27682,N_28143);
nand U31993 (N_31993,N_27619,N_28374);
or U31994 (N_31994,N_29225,N_28134);
and U31995 (N_31995,N_27631,N_27965);
nor U31996 (N_31996,N_28682,N_28720);
nand U31997 (N_31997,N_28036,N_28795);
and U31998 (N_31998,N_29255,N_28171);
and U31999 (N_31999,N_28859,N_28378);
nand U32000 (N_32000,N_29495,N_29191);
nand U32001 (N_32001,N_28480,N_27519);
xor U32002 (N_32002,N_27511,N_28291);
and U32003 (N_32003,N_28561,N_28294);
nor U32004 (N_32004,N_28790,N_27528);
xnor U32005 (N_32005,N_28146,N_27978);
or U32006 (N_32006,N_29148,N_28999);
and U32007 (N_32007,N_29281,N_29812);
nand U32008 (N_32008,N_29849,N_29268);
xor U32009 (N_32009,N_28745,N_27700);
nand U32010 (N_32010,N_28344,N_28921);
or U32011 (N_32011,N_27928,N_28077);
and U32012 (N_32012,N_28954,N_28970);
xnor U32013 (N_32013,N_28860,N_29155);
nand U32014 (N_32014,N_28444,N_29792);
nor U32015 (N_32015,N_29461,N_29201);
nor U32016 (N_32016,N_29579,N_27512);
nand U32017 (N_32017,N_28075,N_29888);
xnor U32018 (N_32018,N_29483,N_29196);
and U32019 (N_32019,N_29255,N_28003);
nor U32020 (N_32020,N_29471,N_27834);
or U32021 (N_32021,N_27832,N_27879);
nor U32022 (N_32022,N_28677,N_29433);
and U32023 (N_32023,N_28375,N_29713);
and U32024 (N_32024,N_29738,N_29785);
or U32025 (N_32025,N_28621,N_29837);
or U32026 (N_32026,N_29265,N_27744);
xor U32027 (N_32027,N_29548,N_29433);
or U32028 (N_32028,N_27619,N_29017);
or U32029 (N_32029,N_28997,N_28995);
xor U32030 (N_32030,N_28844,N_28421);
or U32031 (N_32031,N_29905,N_29695);
nand U32032 (N_32032,N_28215,N_29200);
nand U32033 (N_32033,N_29776,N_29103);
nor U32034 (N_32034,N_29557,N_28376);
nor U32035 (N_32035,N_28757,N_28577);
nand U32036 (N_32036,N_29616,N_29345);
or U32037 (N_32037,N_29479,N_28940);
nor U32038 (N_32038,N_28194,N_29860);
nand U32039 (N_32039,N_28934,N_28591);
nor U32040 (N_32040,N_28072,N_28133);
xnor U32041 (N_32041,N_28687,N_29216);
nand U32042 (N_32042,N_29893,N_28240);
nor U32043 (N_32043,N_28507,N_29806);
and U32044 (N_32044,N_28384,N_29711);
or U32045 (N_32045,N_28473,N_28790);
and U32046 (N_32046,N_27801,N_28936);
xor U32047 (N_32047,N_29056,N_28903);
and U32048 (N_32048,N_28902,N_29938);
and U32049 (N_32049,N_29870,N_29880);
nand U32050 (N_32050,N_28468,N_28748);
xnor U32051 (N_32051,N_29595,N_27953);
nand U32052 (N_32052,N_29920,N_28975);
and U32053 (N_32053,N_28674,N_29140);
nor U32054 (N_32054,N_29625,N_29050);
nor U32055 (N_32055,N_29708,N_29564);
or U32056 (N_32056,N_28142,N_29607);
nor U32057 (N_32057,N_29476,N_28619);
xnor U32058 (N_32058,N_29840,N_29873);
and U32059 (N_32059,N_28758,N_28158);
nor U32060 (N_32060,N_28531,N_29949);
and U32061 (N_32061,N_29535,N_29874);
nor U32062 (N_32062,N_27911,N_27968);
nor U32063 (N_32063,N_28261,N_28436);
xor U32064 (N_32064,N_28192,N_29768);
or U32065 (N_32065,N_29149,N_28395);
and U32066 (N_32066,N_28778,N_29932);
nor U32067 (N_32067,N_27647,N_27683);
xnor U32068 (N_32068,N_29754,N_28729);
xor U32069 (N_32069,N_29437,N_28245);
nand U32070 (N_32070,N_28898,N_28202);
nand U32071 (N_32071,N_27940,N_29328);
or U32072 (N_32072,N_27905,N_28605);
and U32073 (N_32073,N_29296,N_29004);
or U32074 (N_32074,N_27711,N_28051);
nor U32075 (N_32075,N_28749,N_27673);
and U32076 (N_32076,N_28888,N_29166);
nor U32077 (N_32077,N_29219,N_27870);
xnor U32078 (N_32078,N_28133,N_28855);
xnor U32079 (N_32079,N_28035,N_29081);
xor U32080 (N_32080,N_29045,N_29057);
or U32081 (N_32081,N_29099,N_29782);
nand U32082 (N_32082,N_29658,N_28078);
xnor U32083 (N_32083,N_29201,N_29907);
or U32084 (N_32084,N_29428,N_29802);
and U32085 (N_32085,N_29814,N_28725);
or U32086 (N_32086,N_28335,N_28430);
nor U32087 (N_32087,N_28774,N_28733);
nand U32088 (N_32088,N_28432,N_29819);
nand U32089 (N_32089,N_29118,N_29983);
xnor U32090 (N_32090,N_29851,N_28954);
nor U32091 (N_32091,N_29644,N_28222);
and U32092 (N_32092,N_27934,N_29466);
and U32093 (N_32093,N_27995,N_28983);
nor U32094 (N_32094,N_27825,N_27795);
nor U32095 (N_32095,N_29976,N_28873);
and U32096 (N_32096,N_29985,N_29979);
nand U32097 (N_32097,N_28774,N_28849);
and U32098 (N_32098,N_28373,N_29322);
nand U32099 (N_32099,N_28254,N_28495);
nand U32100 (N_32100,N_29554,N_27578);
nand U32101 (N_32101,N_28308,N_29239);
xor U32102 (N_32102,N_29425,N_29732);
nor U32103 (N_32103,N_28047,N_28046);
nand U32104 (N_32104,N_28296,N_27878);
nand U32105 (N_32105,N_29599,N_28586);
nand U32106 (N_32106,N_28687,N_27864);
xnor U32107 (N_32107,N_27979,N_29808);
nor U32108 (N_32108,N_29863,N_27571);
nand U32109 (N_32109,N_29604,N_29724);
or U32110 (N_32110,N_28328,N_29618);
nand U32111 (N_32111,N_27650,N_29934);
nand U32112 (N_32112,N_29965,N_29198);
or U32113 (N_32113,N_28299,N_29979);
nand U32114 (N_32114,N_29282,N_28173);
nand U32115 (N_32115,N_28042,N_28057);
nor U32116 (N_32116,N_29252,N_27854);
or U32117 (N_32117,N_28803,N_27585);
nand U32118 (N_32118,N_28802,N_27915);
or U32119 (N_32119,N_29950,N_29670);
nand U32120 (N_32120,N_28131,N_28869);
and U32121 (N_32121,N_28608,N_28087);
or U32122 (N_32122,N_29506,N_29956);
nor U32123 (N_32123,N_28371,N_28281);
nor U32124 (N_32124,N_29780,N_29496);
and U32125 (N_32125,N_28582,N_28952);
nor U32126 (N_32126,N_28275,N_29760);
nand U32127 (N_32127,N_28839,N_28265);
nor U32128 (N_32128,N_28582,N_28723);
and U32129 (N_32129,N_28603,N_29184);
nor U32130 (N_32130,N_28551,N_29015);
or U32131 (N_32131,N_29048,N_29874);
nand U32132 (N_32132,N_28317,N_29480);
or U32133 (N_32133,N_29923,N_28064);
and U32134 (N_32134,N_28353,N_27908);
xor U32135 (N_32135,N_28085,N_29451);
or U32136 (N_32136,N_29064,N_28188);
and U32137 (N_32137,N_28957,N_29667);
nand U32138 (N_32138,N_28975,N_28573);
nor U32139 (N_32139,N_29132,N_29396);
nor U32140 (N_32140,N_29559,N_28162);
and U32141 (N_32141,N_29787,N_27998);
and U32142 (N_32142,N_29249,N_29899);
xor U32143 (N_32143,N_28032,N_28461);
nand U32144 (N_32144,N_27876,N_29895);
or U32145 (N_32145,N_27892,N_29702);
xor U32146 (N_32146,N_29478,N_28457);
nand U32147 (N_32147,N_27673,N_29119);
or U32148 (N_32148,N_27899,N_29866);
xnor U32149 (N_32149,N_28288,N_28988);
and U32150 (N_32150,N_28719,N_28979);
or U32151 (N_32151,N_28579,N_27880);
and U32152 (N_32152,N_28119,N_28455);
xnor U32153 (N_32153,N_29063,N_27746);
xor U32154 (N_32154,N_28507,N_28093);
or U32155 (N_32155,N_28447,N_27854);
nand U32156 (N_32156,N_29024,N_27676);
nand U32157 (N_32157,N_29011,N_28331);
xnor U32158 (N_32158,N_28476,N_28380);
nand U32159 (N_32159,N_29986,N_28070);
or U32160 (N_32160,N_28581,N_28529);
nand U32161 (N_32161,N_28775,N_29026);
nor U32162 (N_32162,N_27809,N_27638);
nor U32163 (N_32163,N_28675,N_28683);
and U32164 (N_32164,N_29277,N_29774);
or U32165 (N_32165,N_28391,N_29630);
or U32166 (N_32166,N_29955,N_27969);
nor U32167 (N_32167,N_27806,N_29735);
nand U32168 (N_32168,N_29653,N_29260);
and U32169 (N_32169,N_27753,N_29093);
or U32170 (N_32170,N_27879,N_28366);
nor U32171 (N_32171,N_29597,N_28284);
or U32172 (N_32172,N_29807,N_28079);
nand U32173 (N_32173,N_28670,N_28578);
xnor U32174 (N_32174,N_28082,N_29551);
nor U32175 (N_32175,N_29890,N_28989);
xnor U32176 (N_32176,N_28699,N_28367);
nand U32177 (N_32177,N_28008,N_29786);
or U32178 (N_32178,N_28984,N_27858);
or U32179 (N_32179,N_29464,N_29597);
and U32180 (N_32180,N_28723,N_27778);
nand U32181 (N_32181,N_27615,N_29927);
and U32182 (N_32182,N_29583,N_28887);
and U32183 (N_32183,N_28479,N_27533);
and U32184 (N_32184,N_28948,N_29943);
nor U32185 (N_32185,N_28464,N_29648);
nand U32186 (N_32186,N_29238,N_27922);
or U32187 (N_32187,N_27888,N_29527);
nor U32188 (N_32188,N_27794,N_27837);
nor U32189 (N_32189,N_27649,N_29330);
or U32190 (N_32190,N_29353,N_28622);
and U32191 (N_32191,N_28155,N_28945);
or U32192 (N_32192,N_27505,N_29822);
nor U32193 (N_32193,N_29322,N_29661);
nor U32194 (N_32194,N_29300,N_28080);
nand U32195 (N_32195,N_28948,N_28977);
or U32196 (N_32196,N_29457,N_28933);
nand U32197 (N_32197,N_27593,N_28563);
xnor U32198 (N_32198,N_27804,N_27761);
and U32199 (N_32199,N_28320,N_28549);
or U32200 (N_32200,N_28785,N_28011);
nand U32201 (N_32201,N_28375,N_28650);
xor U32202 (N_32202,N_27747,N_28081);
or U32203 (N_32203,N_28431,N_28286);
nand U32204 (N_32204,N_29697,N_29898);
nor U32205 (N_32205,N_29316,N_27936);
nand U32206 (N_32206,N_28120,N_28627);
nand U32207 (N_32207,N_27835,N_28048);
xnor U32208 (N_32208,N_29614,N_28761);
and U32209 (N_32209,N_28812,N_28708);
and U32210 (N_32210,N_29550,N_29321);
and U32211 (N_32211,N_28649,N_28426);
and U32212 (N_32212,N_29841,N_28494);
nor U32213 (N_32213,N_28140,N_27629);
and U32214 (N_32214,N_29651,N_29700);
xnor U32215 (N_32215,N_28181,N_28714);
and U32216 (N_32216,N_27772,N_28816);
xor U32217 (N_32217,N_28310,N_28128);
nand U32218 (N_32218,N_27907,N_28075);
xnor U32219 (N_32219,N_27917,N_28106);
and U32220 (N_32220,N_28368,N_28293);
or U32221 (N_32221,N_28023,N_29408);
nor U32222 (N_32222,N_28591,N_28117);
xor U32223 (N_32223,N_28847,N_28584);
and U32224 (N_32224,N_29364,N_28908);
and U32225 (N_32225,N_29002,N_29935);
nand U32226 (N_32226,N_29351,N_28152);
xor U32227 (N_32227,N_29658,N_28980);
xnor U32228 (N_32228,N_29116,N_29932);
nand U32229 (N_32229,N_27777,N_27927);
nor U32230 (N_32230,N_29334,N_29136);
xnor U32231 (N_32231,N_28596,N_27748);
nor U32232 (N_32232,N_27864,N_28965);
nor U32233 (N_32233,N_28439,N_29299);
nand U32234 (N_32234,N_29745,N_29771);
and U32235 (N_32235,N_29744,N_27641);
nor U32236 (N_32236,N_27694,N_29006);
nand U32237 (N_32237,N_28867,N_28613);
xnor U32238 (N_32238,N_29391,N_28764);
xor U32239 (N_32239,N_28998,N_28246);
xor U32240 (N_32240,N_27540,N_27982);
or U32241 (N_32241,N_29496,N_29990);
nand U32242 (N_32242,N_29062,N_27750);
nand U32243 (N_32243,N_27649,N_28215);
and U32244 (N_32244,N_27968,N_28831);
and U32245 (N_32245,N_28850,N_28629);
nor U32246 (N_32246,N_29000,N_28723);
and U32247 (N_32247,N_27921,N_28143);
or U32248 (N_32248,N_29387,N_27516);
nor U32249 (N_32249,N_29688,N_28233);
and U32250 (N_32250,N_29116,N_28571);
and U32251 (N_32251,N_27700,N_28185);
xor U32252 (N_32252,N_29417,N_28923);
or U32253 (N_32253,N_29731,N_29787);
and U32254 (N_32254,N_29983,N_29586);
nand U32255 (N_32255,N_29959,N_28027);
nand U32256 (N_32256,N_29838,N_29271);
nand U32257 (N_32257,N_29572,N_27644);
nand U32258 (N_32258,N_28901,N_29851);
and U32259 (N_32259,N_27718,N_27700);
xor U32260 (N_32260,N_27579,N_28409);
xor U32261 (N_32261,N_29207,N_27689);
xor U32262 (N_32262,N_29568,N_27763);
or U32263 (N_32263,N_28151,N_27583);
and U32264 (N_32264,N_27647,N_28675);
or U32265 (N_32265,N_28337,N_28499);
or U32266 (N_32266,N_27874,N_28638);
or U32267 (N_32267,N_29021,N_29221);
and U32268 (N_32268,N_27681,N_27796);
and U32269 (N_32269,N_29956,N_29602);
nor U32270 (N_32270,N_28439,N_28009);
and U32271 (N_32271,N_28690,N_29344);
xor U32272 (N_32272,N_28293,N_29075);
or U32273 (N_32273,N_29547,N_29026);
and U32274 (N_32274,N_28277,N_28547);
nand U32275 (N_32275,N_27798,N_27708);
and U32276 (N_32276,N_29887,N_28915);
xor U32277 (N_32277,N_29480,N_29285);
nor U32278 (N_32278,N_27919,N_29627);
or U32279 (N_32279,N_28247,N_29639);
or U32280 (N_32280,N_27705,N_29358);
and U32281 (N_32281,N_29958,N_28797);
or U32282 (N_32282,N_28189,N_29255);
or U32283 (N_32283,N_28645,N_27726);
nand U32284 (N_32284,N_28148,N_28871);
nand U32285 (N_32285,N_28758,N_29085);
xor U32286 (N_32286,N_28802,N_29566);
or U32287 (N_32287,N_29559,N_27599);
nor U32288 (N_32288,N_27921,N_27715);
nand U32289 (N_32289,N_28943,N_29391);
xnor U32290 (N_32290,N_28145,N_27817);
nor U32291 (N_32291,N_29593,N_27825);
or U32292 (N_32292,N_29361,N_29663);
or U32293 (N_32293,N_29541,N_28450);
nor U32294 (N_32294,N_27903,N_27878);
and U32295 (N_32295,N_29162,N_29732);
and U32296 (N_32296,N_29601,N_29524);
nor U32297 (N_32297,N_29613,N_29951);
nand U32298 (N_32298,N_27632,N_29611);
nand U32299 (N_32299,N_29982,N_29418);
nand U32300 (N_32300,N_28780,N_29435);
and U32301 (N_32301,N_29140,N_27776);
xnor U32302 (N_32302,N_29572,N_29948);
xor U32303 (N_32303,N_29980,N_27996);
nand U32304 (N_32304,N_28994,N_29599);
nor U32305 (N_32305,N_28652,N_28020);
xnor U32306 (N_32306,N_28749,N_28547);
nand U32307 (N_32307,N_28858,N_29940);
nand U32308 (N_32308,N_28174,N_28116);
nor U32309 (N_32309,N_28486,N_28474);
nand U32310 (N_32310,N_29336,N_27903);
and U32311 (N_32311,N_29710,N_29271);
and U32312 (N_32312,N_27820,N_28094);
nor U32313 (N_32313,N_28576,N_28833);
and U32314 (N_32314,N_28563,N_29245);
nand U32315 (N_32315,N_28827,N_29925);
and U32316 (N_32316,N_29287,N_28607);
or U32317 (N_32317,N_29638,N_28196);
xor U32318 (N_32318,N_28878,N_28425);
and U32319 (N_32319,N_27676,N_28782);
nand U32320 (N_32320,N_28951,N_28794);
xor U32321 (N_32321,N_29123,N_28566);
or U32322 (N_32322,N_28701,N_29376);
and U32323 (N_32323,N_29388,N_28079);
nand U32324 (N_32324,N_28295,N_29666);
nand U32325 (N_32325,N_28135,N_28309);
and U32326 (N_32326,N_29675,N_29636);
xor U32327 (N_32327,N_28927,N_27622);
nor U32328 (N_32328,N_28271,N_28695);
and U32329 (N_32329,N_29819,N_29509);
nand U32330 (N_32330,N_27709,N_29771);
or U32331 (N_32331,N_28257,N_27620);
nor U32332 (N_32332,N_29576,N_28901);
xor U32333 (N_32333,N_28774,N_27916);
nand U32334 (N_32334,N_28144,N_29662);
xor U32335 (N_32335,N_29162,N_28609);
and U32336 (N_32336,N_29038,N_28909);
nor U32337 (N_32337,N_28803,N_28482);
or U32338 (N_32338,N_29676,N_28383);
xor U32339 (N_32339,N_28624,N_29250);
xor U32340 (N_32340,N_28599,N_28548);
nand U32341 (N_32341,N_28262,N_28458);
or U32342 (N_32342,N_29685,N_28442);
xnor U32343 (N_32343,N_28776,N_28206);
or U32344 (N_32344,N_27520,N_27913);
and U32345 (N_32345,N_27621,N_28321);
nor U32346 (N_32346,N_28942,N_29448);
or U32347 (N_32347,N_29240,N_27710);
nor U32348 (N_32348,N_27758,N_28699);
and U32349 (N_32349,N_28694,N_28484);
nor U32350 (N_32350,N_28486,N_28058);
or U32351 (N_32351,N_29566,N_29029);
or U32352 (N_32352,N_28347,N_28646);
and U32353 (N_32353,N_29246,N_28906);
nor U32354 (N_32354,N_28531,N_27849);
nor U32355 (N_32355,N_29703,N_29565);
xnor U32356 (N_32356,N_27701,N_29517);
and U32357 (N_32357,N_29012,N_27903);
xor U32358 (N_32358,N_28519,N_29384);
nand U32359 (N_32359,N_29491,N_27816);
and U32360 (N_32360,N_28411,N_28261);
xor U32361 (N_32361,N_28479,N_29685);
xnor U32362 (N_32362,N_28157,N_29372);
xnor U32363 (N_32363,N_29490,N_29766);
nor U32364 (N_32364,N_28057,N_28451);
nor U32365 (N_32365,N_29251,N_28066);
nor U32366 (N_32366,N_28732,N_27725);
and U32367 (N_32367,N_29494,N_28847);
nor U32368 (N_32368,N_28474,N_28865);
or U32369 (N_32369,N_28550,N_29518);
and U32370 (N_32370,N_29810,N_27594);
nand U32371 (N_32371,N_27806,N_27528);
nand U32372 (N_32372,N_29865,N_28219);
or U32373 (N_32373,N_27766,N_28900);
nor U32374 (N_32374,N_29869,N_29605);
and U32375 (N_32375,N_28132,N_29792);
xnor U32376 (N_32376,N_28220,N_28889);
nand U32377 (N_32377,N_28057,N_29066);
or U32378 (N_32378,N_28477,N_28592);
and U32379 (N_32379,N_29766,N_28861);
xnor U32380 (N_32380,N_27633,N_28607);
and U32381 (N_32381,N_29323,N_29412);
xor U32382 (N_32382,N_28316,N_27966);
xnor U32383 (N_32383,N_29867,N_27633);
nor U32384 (N_32384,N_28098,N_29425);
nand U32385 (N_32385,N_28605,N_28313);
nor U32386 (N_32386,N_28824,N_28523);
nor U32387 (N_32387,N_28379,N_29162);
and U32388 (N_32388,N_27617,N_27620);
xor U32389 (N_32389,N_29511,N_27649);
and U32390 (N_32390,N_29820,N_28983);
and U32391 (N_32391,N_29980,N_27803);
and U32392 (N_32392,N_28755,N_28053);
nor U32393 (N_32393,N_28110,N_29461);
or U32394 (N_32394,N_29925,N_29834);
xor U32395 (N_32395,N_29699,N_29725);
or U32396 (N_32396,N_27832,N_29680);
and U32397 (N_32397,N_27616,N_28583);
and U32398 (N_32398,N_28389,N_27742);
nor U32399 (N_32399,N_28890,N_28270);
xor U32400 (N_32400,N_28996,N_28303);
nand U32401 (N_32401,N_27695,N_27756);
nand U32402 (N_32402,N_29220,N_28437);
and U32403 (N_32403,N_27935,N_29521);
xor U32404 (N_32404,N_28750,N_28592);
or U32405 (N_32405,N_28865,N_29823);
nor U32406 (N_32406,N_28888,N_28489);
nand U32407 (N_32407,N_28019,N_28072);
nand U32408 (N_32408,N_29882,N_27753);
nor U32409 (N_32409,N_28070,N_28089);
nand U32410 (N_32410,N_27944,N_28493);
xnor U32411 (N_32411,N_28965,N_28814);
nand U32412 (N_32412,N_29181,N_29770);
or U32413 (N_32413,N_29141,N_27668);
and U32414 (N_32414,N_29706,N_28302);
or U32415 (N_32415,N_28525,N_29412);
xnor U32416 (N_32416,N_29385,N_27521);
nand U32417 (N_32417,N_28864,N_29777);
and U32418 (N_32418,N_28929,N_28453);
nor U32419 (N_32419,N_27787,N_27890);
nand U32420 (N_32420,N_27573,N_29977);
nor U32421 (N_32421,N_29773,N_28374);
nand U32422 (N_32422,N_28304,N_29217);
nand U32423 (N_32423,N_29595,N_29612);
nor U32424 (N_32424,N_28373,N_28963);
nor U32425 (N_32425,N_28578,N_29442);
nand U32426 (N_32426,N_27839,N_28566);
or U32427 (N_32427,N_28779,N_29334);
or U32428 (N_32428,N_28794,N_28031);
nor U32429 (N_32429,N_28766,N_28308);
nand U32430 (N_32430,N_28788,N_28762);
xor U32431 (N_32431,N_28308,N_28825);
and U32432 (N_32432,N_29828,N_28981);
nand U32433 (N_32433,N_27543,N_29128);
or U32434 (N_32434,N_29808,N_28069);
nor U32435 (N_32435,N_28446,N_27901);
or U32436 (N_32436,N_28174,N_28794);
and U32437 (N_32437,N_29306,N_27613);
nand U32438 (N_32438,N_27722,N_28884);
nand U32439 (N_32439,N_29025,N_27779);
or U32440 (N_32440,N_29279,N_28245);
xor U32441 (N_32441,N_28097,N_28557);
or U32442 (N_32442,N_29974,N_28052);
xor U32443 (N_32443,N_29403,N_28953);
xor U32444 (N_32444,N_29493,N_29185);
nor U32445 (N_32445,N_28865,N_28233);
nand U32446 (N_32446,N_28067,N_27541);
and U32447 (N_32447,N_27800,N_28071);
nor U32448 (N_32448,N_28339,N_29801);
nand U32449 (N_32449,N_27962,N_29132);
nand U32450 (N_32450,N_28131,N_27504);
and U32451 (N_32451,N_29705,N_28783);
xor U32452 (N_32452,N_28486,N_27851);
and U32453 (N_32453,N_28202,N_28242);
nand U32454 (N_32454,N_28066,N_29531);
xor U32455 (N_32455,N_28114,N_28519);
xnor U32456 (N_32456,N_28369,N_27518);
xnor U32457 (N_32457,N_28626,N_27624);
or U32458 (N_32458,N_29322,N_28306);
nand U32459 (N_32459,N_28265,N_29516);
or U32460 (N_32460,N_28149,N_28560);
xnor U32461 (N_32461,N_29521,N_29111);
nand U32462 (N_32462,N_27569,N_27559);
nor U32463 (N_32463,N_28001,N_28115);
or U32464 (N_32464,N_28891,N_29988);
or U32465 (N_32465,N_28717,N_29538);
or U32466 (N_32466,N_28493,N_27682);
xor U32467 (N_32467,N_28279,N_28843);
or U32468 (N_32468,N_28566,N_28839);
nand U32469 (N_32469,N_27934,N_27562);
xor U32470 (N_32470,N_27682,N_27974);
nand U32471 (N_32471,N_29789,N_28261);
or U32472 (N_32472,N_28373,N_29740);
or U32473 (N_32473,N_28550,N_29719);
or U32474 (N_32474,N_28648,N_28170);
xor U32475 (N_32475,N_29473,N_29732);
nor U32476 (N_32476,N_29433,N_27508);
xor U32477 (N_32477,N_29868,N_28998);
xor U32478 (N_32478,N_28751,N_29325);
and U32479 (N_32479,N_29275,N_28562);
xnor U32480 (N_32480,N_29017,N_29129);
or U32481 (N_32481,N_27855,N_29236);
or U32482 (N_32482,N_28363,N_27702);
xnor U32483 (N_32483,N_27539,N_28788);
nand U32484 (N_32484,N_29490,N_28524);
nand U32485 (N_32485,N_28562,N_29355);
nand U32486 (N_32486,N_28769,N_28837);
xor U32487 (N_32487,N_29997,N_27883);
xnor U32488 (N_32488,N_28792,N_29322);
or U32489 (N_32489,N_29857,N_29746);
and U32490 (N_32490,N_29419,N_29936);
and U32491 (N_32491,N_27809,N_28735);
nor U32492 (N_32492,N_28149,N_27605);
and U32493 (N_32493,N_29320,N_29829);
xor U32494 (N_32494,N_27977,N_29968);
or U32495 (N_32495,N_27993,N_28203);
or U32496 (N_32496,N_28878,N_29795);
xnor U32497 (N_32497,N_28013,N_29270);
nand U32498 (N_32498,N_29643,N_29751);
or U32499 (N_32499,N_29696,N_28064);
nor U32500 (N_32500,N_30340,N_31752);
xor U32501 (N_32501,N_30632,N_30833);
and U32502 (N_32502,N_31872,N_30594);
nand U32503 (N_32503,N_32366,N_30970);
xnor U32504 (N_32504,N_30255,N_31085);
or U32505 (N_32505,N_31481,N_30861);
nand U32506 (N_32506,N_32069,N_30828);
xnor U32507 (N_32507,N_31762,N_31551);
nand U32508 (N_32508,N_30539,N_30895);
nor U32509 (N_32509,N_32143,N_32062);
or U32510 (N_32510,N_31044,N_30644);
nand U32511 (N_32511,N_31440,N_31069);
nand U32512 (N_32512,N_31285,N_31405);
or U32513 (N_32513,N_31870,N_31013);
and U32514 (N_32514,N_30903,N_30488);
nor U32515 (N_32515,N_32419,N_31396);
or U32516 (N_32516,N_31241,N_31091);
xnor U32517 (N_32517,N_31942,N_31247);
nor U32518 (N_32518,N_31781,N_30043);
xor U32519 (N_32519,N_30466,N_31969);
or U32520 (N_32520,N_31531,N_31049);
xor U32521 (N_32521,N_31718,N_30576);
nor U32522 (N_32522,N_30999,N_32256);
xor U32523 (N_32523,N_30480,N_30372);
nor U32524 (N_32524,N_30946,N_31798);
nand U32525 (N_32525,N_31641,N_31731);
xnor U32526 (N_32526,N_31499,N_31856);
xnor U32527 (N_32527,N_30383,N_31146);
or U32528 (N_32528,N_31910,N_32487);
xor U32529 (N_32529,N_31884,N_32036);
or U32530 (N_32530,N_31542,N_32161);
nor U32531 (N_32531,N_31136,N_30140);
nand U32532 (N_32532,N_32345,N_31796);
xnor U32533 (N_32533,N_32037,N_30408);
xnor U32534 (N_32534,N_31469,N_32023);
or U32535 (N_32535,N_32190,N_32026);
xor U32536 (N_32536,N_31135,N_30444);
or U32537 (N_32537,N_30770,N_31416);
xnor U32538 (N_32538,N_30844,N_30750);
nor U32539 (N_32539,N_31650,N_31377);
nand U32540 (N_32540,N_30399,N_32425);
or U32541 (N_32541,N_30580,N_31073);
nand U32542 (N_32542,N_30013,N_30223);
nor U32543 (N_32543,N_30469,N_30797);
and U32544 (N_32544,N_31141,N_31101);
xnor U32545 (N_32545,N_31835,N_30270);
or U32546 (N_32546,N_30416,N_32112);
or U32547 (N_32547,N_32310,N_30085);
and U32548 (N_32548,N_30356,N_31090);
xor U32549 (N_32549,N_31684,N_31735);
and U32550 (N_32550,N_31053,N_31704);
or U32551 (N_32551,N_30190,N_31140);
nand U32552 (N_32552,N_31239,N_30942);
xnor U32553 (N_32553,N_31970,N_32068);
xnor U32554 (N_32554,N_31738,N_32410);
xnor U32555 (N_32555,N_30387,N_31012);
or U32556 (N_32556,N_31240,N_31603);
xnor U32557 (N_32557,N_31654,N_30202);
or U32558 (N_32558,N_32265,N_32395);
or U32559 (N_32559,N_31382,N_31436);
xor U32560 (N_32560,N_31423,N_31930);
xor U32561 (N_32561,N_31768,N_31778);
or U32562 (N_32562,N_31895,N_31476);
nor U32563 (N_32563,N_30809,N_30003);
xnor U32564 (N_32564,N_30613,N_30597);
nand U32565 (N_32565,N_32232,N_30005);
nor U32566 (N_32566,N_31452,N_32329);
and U32567 (N_32567,N_32471,N_30868);
nand U32568 (N_32568,N_30051,N_30306);
nor U32569 (N_32569,N_31419,N_30755);
or U32570 (N_32570,N_31133,N_32268);
nand U32571 (N_32571,N_32040,N_31625);
and U32572 (N_32572,N_30441,N_31689);
nor U32573 (N_32573,N_31678,N_31034);
nand U32574 (N_32574,N_31183,N_31864);
or U32575 (N_32575,N_31501,N_30450);
nor U32576 (N_32576,N_31088,N_31984);
nor U32577 (N_32577,N_31611,N_31299);
or U32578 (N_32578,N_31609,N_30495);
xnor U32579 (N_32579,N_30272,N_31878);
and U32580 (N_32580,N_31404,N_32183);
xor U32581 (N_32581,N_31646,N_30757);
and U32582 (N_32582,N_31937,N_31275);
nand U32583 (N_32583,N_31842,N_31258);
and U32584 (N_32584,N_30351,N_30117);
and U32585 (N_32585,N_31604,N_32015);
nand U32586 (N_32586,N_32375,N_31474);
and U32587 (N_32587,N_31020,N_30607);
or U32588 (N_32588,N_30025,N_32483);
xor U32589 (N_32589,N_31791,N_30804);
xor U32590 (N_32590,N_30731,N_31394);
nor U32591 (N_32591,N_30104,N_31276);
and U32592 (N_32592,N_31026,N_31576);
nor U32593 (N_32593,N_31397,N_30534);
nand U32594 (N_32594,N_30460,N_30982);
nor U32595 (N_32595,N_30693,N_31047);
or U32596 (N_32596,N_31430,N_32218);
nand U32597 (N_32597,N_32398,N_30195);
or U32598 (N_32598,N_31690,N_31993);
xor U32599 (N_32599,N_31766,N_31729);
nand U32600 (N_32600,N_30902,N_30972);
and U32601 (N_32601,N_32133,N_31675);
nand U32602 (N_32602,N_32450,N_31225);
xnor U32603 (N_32603,N_30881,N_30978);
and U32604 (N_32604,N_30478,N_30337);
nor U32605 (N_32605,N_30121,N_31573);
nand U32606 (N_32606,N_32373,N_31407);
or U32607 (N_32607,N_31269,N_31010);
and U32608 (N_32608,N_31901,N_30887);
nand U32609 (N_32609,N_31771,N_32065);
nor U32610 (N_32610,N_30873,N_30217);
and U32611 (N_32611,N_31431,N_31896);
and U32612 (N_32612,N_32246,N_31822);
or U32613 (N_32613,N_30280,N_30886);
and U32614 (N_32614,N_31871,N_30932);
or U32615 (N_32615,N_31996,N_31277);
xnor U32616 (N_32616,N_30960,N_32052);
or U32617 (N_32617,N_31787,N_30605);
nand U32618 (N_32618,N_32423,N_30560);
nand U32619 (N_32619,N_31165,N_31504);
xnor U32620 (N_32620,N_30465,N_31888);
or U32621 (N_32621,N_31783,N_32432);
and U32622 (N_32622,N_30076,N_31446);
nand U32623 (N_32623,N_32012,N_30907);
xnor U32624 (N_32624,N_31686,N_32481);
or U32625 (N_32625,N_32048,N_32353);
nor U32626 (N_32626,N_30407,N_32418);
nor U32627 (N_32627,N_30055,N_30122);
xnor U32628 (N_32628,N_31202,N_31443);
and U32629 (N_32629,N_30850,N_30401);
or U32630 (N_32630,N_32405,N_32475);
or U32631 (N_32631,N_31972,N_30516);
nor U32632 (N_32632,N_32223,N_30393);
and U32633 (N_32633,N_30134,N_30359);
nand U32634 (N_32634,N_30634,N_30163);
nor U32635 (N_32635,N_30510,N_30133);
and U32636 (N_32636,N_30676,N_30866);
nor U32637 (N_32637,N_31544,N_31311);
or U32638 (N_32638,N_32074,N_31663);
and U32639 (N_32639,N_30691,N_31425);
nor U32640 (N_32640,N_30506,N_30323);
nor U32641 (N_32641,N_30290,N_32472);
xor U32642 (N_32642,N_31294,N_30363);
and U32643 (N_32643,N_32257,N_32426);
nor U32644 (N_32644,N_30295,N_31218);
xor U32645 (N_32645,N_31310,N_32097);
or U32646 (N_32646,N_31659,N_30740);
nor U32647 (N_32647,N_30034,N_31960);
nand U32648 (N_32648,N_30603,N_31229);
xor U32649 (N_32649,N_32184,N_31913);
nor U32650 (N_32650,N_32478,N_31074);
nor U32651 (N_32651,N_31326,N_30437);
xor U32652 (N_32652,N_30114,N_31040);
or U32653 (N_32653,N_32182,N_31224);
xnor U32654 (N_32654,N_30494,N_30264);
xor U32655 (N_32655,N_32131,N_32121);
and U32656 (N_32656,N_30662,N_32018);
or U32657 (N_32657,N_30979,N_32358);
nand U32658 (N_32658,N_31702,N_31614);
nor U32659 (N_32659,N_30412,N_30968);
nand U32660 (N_32660,N_30279,N_30775);
nand U32661 (N_32661,N_31209,N_32193);
and U32662 (N_32662,N_32394,N_31355);
and U32663 (N_32663,N_31174,N_31818);
or U32664 (N_32664,N_30829,N_30414);
xnor U32665 (N_32665,N_30105,N_32128);
nor U32666 (N_32666,N_31774,N_30966);
nor U32667 (N_32667,N_30319,N_30853);
nor U32668 (N_32668,N_32466,N_32014);
or U32669 (N_32669,N_31959,N_32046);
nand U32670 (N_32670,N_32059,N_30514);
nand U32671 (N_32671,N_30339,N_30548);
and U32672 (N_32672,N_31643,N_32239);
or U32673 (N_32673,N_30763,N_30957);
or U32674 (N_32674,N_31500,N_31869);
xor U32675 (N_32675,N_30476,N_32031);
xnor U32676 (N_32676,N_31347,N_31372);
and U32677 (N_32677,N_31914,N_31639);
xor U32678 (N_32678,N_31279,N_32399);
xnor U32679 (N_32679,N_31360,N_30878);
xnor U32680 (N_32680,N_31812,N_32490);
and U32681 (N_32681,N_31817,N_30183);
xnor U32682 (N_32682,N_32259,N_31495);
xor U32683 (N_32683,N_30382,N_31509);
nor U32684 (N_32684,N_30312,N_32420);
or U32685 (N_32685,N_31213,N_32173);
or U32686 (N_32686,N_31712,N_30536);
or U32687 (N_32687,N_31541,N_30302);
xnor U32688 (N_32688,N_31624,N_32280);
xor U32689 (N_32689,N_32007,N_31737);
nor U32690 (N_32690,N_31084,N_32449);
nor U32691 (N_32691,N_31223,N_32462);
nand U32692 (N_32692,N_32099,N_30916);
nor U32693 (N_32693,N_31666,N_32124);
and U32694 (N_32694,N_31521,N_31761);
or U32695 (N_32695,N_31645,N_30761);
and U32696 (N_32696,N_32319,N_30220);
nand U32697 (N_32697,N_31118,N_31612);
or U32698 (N_32698,N_32371,N_30404);
or U32699 (N_32699,N_32075,N_30325);
nand U32700 (N_32700,N_30839,N_30622);
and U32701 (N_32701,N_30378,N_30377);
or U32702 (N_32702,N_30214,N_32192);
or U32703 (N_32703,N_30699,N_31490);
nor U32704 (N_32704,N_30894,N_32365);
or U32705 (N_32705,N_30588,N_31580);
or U32706 (N_32706,N_31410,N_31222);
or U32707 (N_32707,N_30322,N_30764);
nor U32708 (N_32708,N_31454,N_30213);
or U32709 (N_32709,N_31743,N_31932);
xor U32710 (N_32710,N_30928,N_31707);
and U32711 (N_32711,N_30798,N_30586);
and U32712 (N_32712,N_32307,N_31600);
or U32713 (N_32713,N_32221,N_31006);
nand U32714 (N_32714,N_31099,N_30723);
or U32715 (N_32715,N_32157,N_30940);
or U32716 (N_32716,N_31777,N_32388);
nand U32717 (N_32717,N_32455,N_31456);
xnor U32718 (N_32718,N_30063,N_31636);
xnor U32719 (N_32719,N_30824,N_30008);
xor U32720 (N_32720,N_30838,N_30965);
nor U32721 (N_32721,N_31364,N_30053);
and U32722 (N_32722,N_30595,N_32339);
and U32723 (N_32723,N_31056,N_31992);
nor U32724 (N_32724,N_30896,N_30532);
nor U32725 (N_32725,N_31336,N_31522);
xnor U32726 (N_32726,N_31082,N_30637);
nor U32727 (N_32727,N_32393,N_32211);
nor U32728 (N_32728,N_31291,N_32468);
nor U32729 (N_32729,N_32202,N_31115);
nor U32730 (N_32730,N_31320,N_31994);
or U32731 (N_32731,N_30246,N_32251);
nor U32732 (N_32732,N_31890,N_31703);
and U32733 (N_32733,N_30705,N_30289);
and U32734 (N_32734,N_30297,N_32126);
nand U32735 (N_32735,N_30242,N_32095);
nand U32736 (N_32736,N_31879,N_31962);
or U32737 (N_32737,N_30386,N_30353);
nor U32738 (N_32738,N_31158,N_31716);
xnor U32739 (N_32739,N_30426,N_30483);
xnor U32740 (N_32740,N_31071,N_30474);
nor U32741 (N_32741,N_31687,N_30248);
and U32742 (N_32742,N_31676,N_31184);
nor U32743 (N_32743,N_32486,N_31851);
nor U32744 (N_32744,N_31943,N_32174);
xnor U32745 (N_32745,N_30352,N_30899);
and U32746 (N_32746,N_32364,N_30031);
or U32747 (N_32747,N_30333,N_32195);
and U32748 (N_32748,N_30354,N_31750);
nor U32749 (N_32749,N_30590,N_30796);
and U32750 (N_32750,N_30821,N_32100);
nand U32751 (N_32751,N_31935,N_31618);
and U32752 (N_32752,N_30395,N_30842);
xnor U32753 (N_32753,N_31885,N_31839);
or U32754 (N_32754,N_31862,N_31980);
nor U32755 (N_32755,N_30934,N_31867);
xnor U32756 (N_32756,N_30477,N_32269);
xnor U32757 (N_32757,N_31685,N_30923);
and U32758 (N_32758,N_31964,N_31232);
nor U32759 (N_32759,N_30834,N_31765);
nand U32760 (N_32760,N_30533,N_30253);
and U32761 (N_32761,N_30127,N_30846);
nor U32762 (N_32762,N_31036,N_31536);
nand U32763 (N_32763,N_31233,N_31242);
nand U32764 (N_32764,N_31249,N_31441);
and U32765 (N_32765,N_32130,N_31965);
and U32766 (N_32766,N_30274,N_31802);
nor U32767 (N_32767,N_32087,N_32227);
and U32768 (N_32768,N_30931,N_31097);
nor U32769 (N_32769,N_30374,N_31529);
xor U32770 (N_32770,N_32167,N_30618);
and U32771 (N_32771,N_30350,N_32109);
and U32772 (N_32772,N_31782,N_32476);
and U32773 (N_32773,N_32288,N_30102);
nand U32774 (N_32774,N_30197,N_32303);
nor U32775 (N_32775,N_30663,N_31722);
xor U32776 (N_32776,N_32281,N_32457);
xor U32777 (N_32777,N_30046,N_30449);
and U32778 (N_32778,N_31042,N_30285);
or U32779 (N_32779,N_32350,N_30727);
or U32780 (N_32780,N_31278,N_31301);
or U32781 (N_32781,N_31023,N_30915);
nand U32782 (N_32782,N_31668,N_30028);
nor U32783 (N_32783,N_31583,N_30679);
or U32784 (N_32784,N_30569,N_31078);
xnor U32785 (N_32785,N_32179,N_30068);
or U32786 (N_32786,N_30985,N_31527);
or U32787 (N_32787,N_30331,N_30816);
and U32788 (N_32788,N_32219,N_31706);
and U32789 (N_32789,N_31303,N_30511);
and U32790 (N_32790,N_32374,N_30880);
nor U32791 (N_32791,N_31831,N_31967);
and U32792 (N_32792,N_30540,N_32196);
nand U32793 (N_32793,N_32497,N_30119);
xnor U32794 (N_32794,N_30519,N_30759);
nor U32795 (N_32795,N_30059,N_31148);
xnor U32796 (N_32796,N_30448,N_32488);
or U32797 (N_32797,N_31058,N_30281);
nor U32798 (N_32798,N_32278,N_30874);
and U32799 (N_32799,N_32038,N_31161);
or U32800 (N_32800,N_31516,N_32140);
nor U32801 (N_32801,N_32261,N_31730);
nor U32802 (N_32802,N_31092,N_30097);
xnor U32803 (N_32803,N_31472,N_30888);
or U32804 (N_32804,N_31462,N_30268);
and U32805 (N_32805,N_31079,N_30981);
xor U32806 (N_32806,N_31444,N_30391);
or U32807 (N_32807,N_30461,N_31849);
and U32808 (N_32808,N_32020,N_30777);
nor U32809 (N_32809,N_31432,N_31426);
xor U32810 (N_32810,N_31715,N_30230);
xor U32811 (N_32811,N_30400,N_30701);
xnor U32812 (N_32812,N_31022,N_30115);
xor U32813 (N_32813,N_31832,N_31528);
nor U32814 (N_32814,N_30252,N_31857);
xnor U32815 (N_32815,N_31916,N_31453);
nand U32816 (N_32816,N_31840,N_32315);
nand U32817 (N_32817,N_31555,N_31900);
nor U32818 (N_32818,N_30819,N_30528);
xnor U32819 (N_32819,N_31717,N_31597);
nand U32820 (N_32820,N_30481,N_31238);
or U32821 (N_32821,N_30871,N_30309);
nor U32822 (N_32822,N_30259,N_30434);
xor U32823 (N_32823,N_30633,N_30326);
nand U32824 (N_32824,N_32258,N_30675);
or U32825 (N_32825,N_31785,N_30530);
xor U32826 (N_32826,N_31958,N_30950);
nand U32827 (N_32827,N_31596,N_31087);
nand U32828 (N_32828,N_32060,N_30825);
and U32829 (N_32829,N_31804,N_32103);
nor U32830 (N_32830,N_30423,N_30961);
nor U32831 (N_32831,N_32044,N_32215);
and U32832 (N_32832,N_30418,N_31330);
or U32833 (N_32833,N_30527,N_31934);
nand U32834 (N_32834,N_30311,N_31633);
and U32835 (N_32835,N_31581,N_30039);
xor U32836 (N_32836,N_30935,N_30219);
xnor U32837 (N_32837,N_31350,N_32204);
xor U32838 (N_32838,N_31331,N_30152);
or U32839 (N_32839,N_31054,N_32404);
nand U32840 (N_32840,N_31830,N_30815);
or U32841 (N_32841,N_32252,N_31809);
nand U32842 (N_32842,N_30566,N_32360);
or U32843 (N_32843,N_30917,N_31484);
xor U32844 (N_32844,N_32104,N_30831);
xnor U32845 (N_32845,N_30430,N_30199);
xnor U32846 (N_32846,N_31324,N_30558);
xor U32847 (N_32847,N_30145,N_30573);
and U32848 (N_32848,N_32206,N_31414);
and U32849 (N_32849,N_32108,N_32331);
xnor U32850 (N_32850,N_31800,N_32162);
or U32851 (N_32851,N_31451,N_31093);
and U32852 (N_32852,N_30172,N_30914);
or U32853 (N_32853,N_30371,N_30616);
or U32854 (N_32854,N_31898,N_32168);
or U32855 (N_32855,N_31585,N_32146);
xnor U32856 (N_32856,N_30107,N_31578);
xnor U32857 (N_32857,N_32448,N_32111);
nor U32858 (N_32858,N_31312,N_30329);
xnor U32859 (N_32859,N_30164,N_30176);
and U32860 (N_32860,N_31282,N_30572);
nand U32861 (N_32861,N_31956,N_32189);
and U32862 (N_32862,N_32032,N_31357);
xnor U32863 (N_32863,N_32186,N_30417);
or U32864 (N_32864,N_30628,N_32004);
nand U32865 (N_32865,N_30546,N_30486);
and U32866 (N_32866,N_32053,N_31941);
nand U32867 (N_32867,N_32429,N_30037);
xnor U32868 (N_32868,N_31723,N_30370);
nand U32869 (N_32869,N_30501,N_31651);
and U32870 (N_32870,N_30549,N_31671);
nor U32871 (N_32871,N_30041,N_30835);
nand U32872 (N_32872,N_31726,N_31488);
nor U32873 (N_32873,N_30865,N_32006);
or U32874 (N_32874,N_30080,N_31098);
nand U32875 (N_32875,N_31439,N_31117);
nor U32876 (N_32876,N_31848,N_32297);
nand U32877 (N_32877,N_31507,N_30784);
nor U32878 (N_32878,N_30189,N_30265);
or U32879 (N_32879,N_31400,N_30345);
and U32880 (N_32880,N_32338,N_31007);
and U32881 (N_32881,N_32271,N_32378);
and U32882 (N_32882,N_30707,N_31001);
or U32883 (N_32883,N_30084,N_30027);
nor U32884 (N_32884,N_31658,N_30807);
or U32885 (N_32885,N_30680,N_31978);
and U32886 (N_32886,N_31656,N_31710);
and U32887 (N_32887,N_30168,N_31039);
and U32888 (N_32888,N_30467,N_32066);
nand U32889 (N_32889,N_32079,N_30991);
nand U32890 (N_32890,N_32009,N_32241);
xor U32891 (N_32891,N_31100,N_31295);
xnor U32892 (N_32892,N_30656,N_31048);
and U32893 (N_32893,N_31351,N_31272);
and U32894 (N_32894,N_32230,N_31961);
nand U32895 (N_32895,N_31052,N_30535);
nand U32896 (N_32896,N_31880,N_31228);
or U32897 (N_32897,N_30012,N_32477);
and U32898 (N_32898,N_30298,N_30860);
xor U32899 (N_32899,N_31450,N_30050);
and U32900 (N_32900,N_31024,N_32160);
or U32901 (N_32901,N_30715,N_30581);
xnor U32902 (N_32902,N_30621,N_30475);
or U32903 (N_32903,N_31179,N_30889);
nor U32904 (N_32904,N_31369,N_31953);
nor U32905 (N_32905,N_32349,N_31403);
and U32906 (N_32906,N_31950,N_32090);
xor U32907 (N_32907,N_31734,N_31907);
nand U32908 (N_32908,N_31727,N_30228);
or U32909 (N_32909,N_30582,N_32050);
and U32910 (N_32910,N_30093,N_31619);
or U32911 (N_32911,N_30541,N_31065);
nand U32912 (N_32912,N_31709,N_30070);
nor U32913 (N_32913,N_31297,N_30678);
and U32914 (N_32914,N_31893,N_30987);
nor U32915 (N_32915,N_30192,N_30668);
or U32916 (N_32916,N_31801,N_30160);
xor U32917 (N_32917,N_32484,N_30882);
nand U32918 (N_32918,N_31045,N_31392);
nand U32919 (N_32919,N_30847,N_30368);
nor U32920 (N_32920,N_30704,N_31353);
nor U32921 (N_32921,N_31721,N_30989);
nand U32922 (N_32922,N_31338,N_31487);
nor U32923 (N_32923,N_30849,N_30069);
nand U32924 (N_32924,N_31828,N_31997);
nor U32925 (N_32925,N_32102,N_31083);
nand U32926 (N_32926,N_31317,N_31463);
nand U32927 (N_32927,N_30708,N_31120);
xnor U32928 (N_32928,N_31027,N_32342);
or U32929 (N_32929,N_31810,N_30938);
nor U32930 (N_32930,N_32326,N_30029);
or U32931 (N_32931,N_31672,N_31549);
nor U32932 (N_32932,N_31182,N_31323);
and U32933 (N_32933,N_31041,N_30921);
or U32934 (N_32934,N_30459,N_32286);
and U32935 (N_32935,N_31128,N_31698);
nand U32936 (N_32936,N_30032,N_30026);
nand U32937 (N_32937,N_32123,N_30876);
nor U32938 (N_32938,N_30143,N_31163);
nor U32939 (N_32939,N_30952,N_31846);
nand U32940 (N_32940,N_30648,N_31449);
nor U32941 (N_32941,N_31153,N_31003);
nor U32942 (N_32942,N_30170,N_31909);
xor U32943 (N_32943,N_30342,N_31427);
and U32944 (N_32944,N_30925,N_32422);
and U32945 (N_32945,N_31559,N_30287);
and U32946 (N_32946,N_31327,N_31915);
or U32947 (N_32947,N_31199,N_30512);
and U32948 (N_32948,N_32135,N_31471);
and U32949 (N_32949,N_30867,N_31075);
nor U32950 (N_32950,N_32073,N_30905);
and U32951 (N_32951,N_30947,N_30571);
or U32952 (N_32952,N_31605,N_32430);
nor U32953 (N_32953,N_30443,N_31928);
xor U32954 (N_32954,N_31180,N_31560);
nand U32955 (N_32955,N_31234,N_30073);
xnor U32956 (N_32956,N_30686,N_31479);
nor U32957 (N_32957,N_32470,N_31571);
nand U32958 (N_32958,N_32299,N_30507);
xnor U32959 (N_32959,N_30000,N_30254);
xor U32960 (N_32960,N_30653,N_31497);
and U32961 (N_32961,N_30619,N_30725);
or U32962 (N_32962,N_32228,N_31437);
nor U32963 (N_32963,N_31483,N_30638);
or U32964 (N_32964,N_32116,N_30305);
or U32965 (N_32965,N_31442,N_30271);
nand U32966 (N_32966,N_31626,N_31582);
and U32967 (N_32967,N_31584,N_30484);
and U32968 (N_32968,N_31577,N_31506);
xor U32969 (N_32969,N_30049,N_30801);
and U32970 (N_32970,N_31971,N_31126);
xor U32971 (N_32971,N_30071,N_30181);
xnor U32972 (N_32972,N_31070,N_32151);
xor U32973 (N_32973,N_30949,N_31307);
xor U32974 (N_32974,N_30310,N_31985);
nand U32975 (N_32975,N_31029,N_31647);
and U32976 (N_32976,N_31754,N_31906);
or U32977 (N_32977,N_32270,N_32443);
or U32978 (N_32978,N_30313,N_30706);
xor U32979 (N_32979,N_32197,N_31216);
or U32980 (N_32980,N_30373,N_30738);
nand U32981 (N_32981,N_31968,N_31923);
and U32982 (N_32982,N_30714,N_30110);
xor U32983 (N_32983,N_31477,N_31922);
nand U32984 (N_32984,N_30742,N_30225);
nor U32985 (N_32985,N_30317,N_30198);
nor U32986 (N_32986,N_32320,N_30380);
xor U32987 (N_32987,N_31459,N_31569);
xnor U32988 (N_32988,N_32367,N_31236);
nor U32989 (N_32989,N_31066,N_32141);
nor U32990 (N_32990,N_31011,N_30986);
xnor U32991 (N_32991,N_30379,N_31185);
nor U32992 (N_32992,N_31325,N_30262);
nand U32993 (N_32993,N_30455,N_31825);
nand U32994 (N_32994,N_31681,N_30939);
nand U32995 (N_32995,N_31543,N_30733);
or U32996 (N_32996,N_30496,N_31553);
xnor U32997 (N_32997,N_30741,N_32273);
or U32998 (N_32998,N_30698,N_30283);
or U32999 (N_32999,N_31017,N_31393);
and U33000 (N_33000,N_31524,N_30859);
or U33001 (N_33001,N_30002,N_30756);
nor U33002 (N_33002,N_30403,N_31535);
nor U33003 (N_33003,N_31617,N_32263);
nand U33004 (N_33004,N_30263,N_31514);
nor U33005 (N_33005,N_31464,N_32370);
nor U33006 (N_33006,N_32291,N_32117);
xor U33007 (N_33007,N_31788,N_30036);
and U33008 (N_33008,N_31669,N_30497);
and U33009 (N_33009,N_31623,N_31480);
nor U33010 (N_33010,N_30601,N_32424);
or U33011 (N_33011,N_32498,N_31019);
nor U33012 (N_33012,N_30885,N_31109);
xnor U33013 (N_33013,N_32152,N_32019);
xor U33014 (N_33014,N_31220,N_30606);
or U33015 (N_33015,N_30627,N_30789);
or U33016 (N_33016,N_32456,N_30808);
or U33017 (N_33017,N_31334,N_31122);
and U33018 (N_33018,N_30792,N_31304);
or U33019 (N_33019,N_30338,N_30453);
or U33020 (N_33020,N_32057,N_31305);
nand U33021 (N_33021,N_31503,N_31805);
or U33022 (N_33022,N_31170,N_32372);
nor U33023 (N_33023,N_31927,N_30149);
nor U33024 (N_33024,N_32137,N_30381);
nor U33025 (N_33025,N_30361,N_31362);
nand U33026 (N_33026,N_31466,N_31741);
or U33027 (N_33027,N_30433,N_31342);
or U33028 (N_33028,N_30760,N_30587);
or U33029 (N_33029,N_30623,N_31843);
nor U33030 (N_33030,N_31366,N_31564);
nor U33031 (N_33031,N_30848,N_30717);
or U33032 (N_33032,N_31986,N_32305);
and U33033 (N_33033,N_31475,N_31945);
nor U33034 (N_33034,N_31339,N_31132);
nand U33035 (N_33035,N_30139,N_32454);
and U33036 (N_33036,N_32163,N_31046);
nand U33037 (N_33037,N_31981,N_32341);
or U33038 (N_33038,N_31417,N_31660);
xnor U33039 (N_33039,N_32279,N_30951);
or U33040 (N_33040,N_31955,N_32042);
or U33041 (N_33041,N_30967,N_30650);
xor U33042 (N_33042,N_30752,N_31271);
nand U33043 (N_33043,N_31917,N_30390);
nand U33044 (N_33044,N_31770,N_30445);
or U33045 (N_33045,N_31627,N_32045);
nor U33046 (N_33046,N_31156,N_30840);
or U33047 (N_33047,N_31855,N_31751);
or U33048 (N_33048,N_30162,N_31433);
or U33049 (N_33049,N_30411,N_30826);
and U33050 (N_33050,N_31813,N_31226);
nand U33051 (N_33051,N_30300,N_30278);
or U33052 (N_33052,N_30624,N_30196);
nor U33053 (N_33053,N_32061,N_31385);
or U33054 (N_33054,N_32224,N_31705);
and U33055 (N_33055,N_30392,N_31401);
nand U33056 (N_33056,N_30232,N_30021);
or U33057 (N_33057,N_30666,N_30747);
and U33058 (N_33058,N_30427,N_30321);
nor U33059 (N_33059,N_32368,N_31205);
nor U33060 (N_33060,N_30743,N_30504);
nand U33061 (N_33061,N_31883,N_30805);
xor U33062 (N_33062,N_32234,N_30556);
nand U33063 (N_33063,N_30577,N_32205);
and U33064 (N_33064,N_30006,N_32292);
and U33065 (N_33065,N_31319,N_31590);
nand U33066 (N_33066,N_31261,N_32411);
and U33067 (N_33067,N_31060,N_30695);
xor U33068 (N_33068,N_30113,N_31395);
nor U33069 (N_33069,N_30813,N_30710);
nor U33070 (N_33070,N_31114,N_32386);
or U33071 (N_33071,N_32225,N_30276);
nor U33072 (N_33072,N_30249,N_31198);
xor U33073 (N_33073,N_31015,N_30131);
xnor U33074 (N_33074,N_31823,N_32283);
and U33075 (N_33075,N_30366,N_32262);
and U33076 (N_33076,N_30664,N_31566);
nand U33077 (N_33077,N_31283,N_30229);
and U33078 (N_33078,N_31435,N_31237);
nor U33079 (N_33079,N_30671,N_32402);
and U33080 (N_33080,N_31760,N_30958);
nor U33081 (N_33081,N_30030,N_31876);
and U33082 (N_33082,N_31892,N_30179);
nand U33083 (N_33083,N_30995,N_31207);
or U33084 (N_33084,N_31337,N_30286);
or U33085 (N_33085,N_31838,N_30221);
or U33086 (N_33086,N_30611,N_30920);
nor U33087 (N_33087,N_32433,N_30732);
xnor U33088 (N_33088,N_30016,N_30778);
nor U33089 (N_33089,N_31987,N_31063);
xor U33090 (N_33090,N_31667,N_31868);
or U33091 (N_33091,N_30201,N_31143);
or U33092 (N_33092,N_30200,N_31448);
nor U33093 (N_33093,N_30685,N_31784);
xor U33094 (N_33094,N_31557,N_32125);
nor U33095 (N_33095,N_30703,N_32028);
nor U33096 (N_33096,N_30694,N_30515);
nor U33097 (N_33097,N_30803,N_31653);
xnor U33098 (N_33098,N_30472,N_31379);
nor U33099 (N_33099,N_31328,N_31748);
nor U33100 (N_33100,N_31982,N_31266);
nand U33101 (N_33101,N_31203,N_30458);
nor U33102 (N_33102,N_31539,N_30142);
and U33103 (N_33103,N_31106,N_30419);
nand U33104 (N_33104,N_30711,N_30126);
or U33105 (N_33105,N_30659,N_30235);
or U33106 (N_33106,N_30729,N_30904);
or U33107 (N_33107,N_30617,N_30898);
and U33108 (N_33108,N_32330,N_30175);
xor U33109 (N_33109,N_31877,N_32002);
nand U33110 (N_33110,N_31235,N_32434);
nor U33111 (N_33111,N_31554,N_31378);
or U33112 (N_33112,N_31300,N_31094);
xor U33113 (N_33113,N_31176,N_31467);
xor U33114 (N_33114,N_31998,N_30737);
nand U33115 (N_33115,N_30347,N_31616);
or U33116 (N_33116,N_31391,N_30817);
nor U33117 (N_33117,N_31215,N_30665);
nor U33118 (N_33118,N_32030,N_30247);
or U33119 (N_33119,N_31370,N_30786);
nor U33120 (N_33120,N_30520,N_32198);
and U33121 (N_33121,N_31593,N_30677);
or U33122 (N_33122,N_32172,N_31990);
xnor U33123 (N_33123,N_31591,N_32359);
nor U33124 (N_33124,N_32453,N_31111);
nor U33125 (N_33125,N_31806,N_31221);
and U33126 (N_33126,N_31018,N_30781);
nand U33127 (N_33127,N_30518,N_31308);
nor U33128 (N_33128,N_32473,N_30089);
and U33129 (N_33129,N_30945,N_30349);
nand U33130 (N_33130,N_30924,N_32164);
or U33131 (N_33131,N_31976,N_31567);
nor U33132 (N_33132,N_32089,N_30498);
xnor U33133 (N_33133,N_30245,N_32134);
nor U33134 (N_33134,N_31640,N_31652);
nor U33135 (N_33135,N_30877,N_32400);
xor U33136 (N_33136,N_32445,N_30078);
nand U33137 (N_33137,N_31732,N_31505);
nand U33138 (N_33138,N_30505,N_30209);
or U33139 (N_33139,N_32311,N_30858);
and U33140 (N_33140,N_31365,N_31713);
or U33141 (N_33141,N_31677,N_30812);
nand U33142 (N_33142,N_32391,N_31096);
and U33143 (N_33143,N_31072,N_32496);
nand U33144 (N_33144,N_31649,N_32119);
xnor U33145 (N_33145,N_32442,N_32494);
or U33146 (N_33146,N_32499,N_30522);
nand U33147 (N_33147,N_30802,N_32107);
nor U33148 (N_33148,N_30344,N_30035);
or U33149 (N_33149,N_31127,N_32013);
and U33150 (N_33150,N_31465,N_30746);
nor U33151 (N_33151,N_30040,N_32158);
nand U33152 (N_33152,N_31428,N_32188);
nand U33153 (N_33153,N_31861,N_32153);
nand U33154 (N_33154,N_32324,N_31389);
or U33155 (N_33155,N_30630,N_30769);
nand U33156 (N_33156,N_32308,N_30208);
and U33157 (N_33157,N_30681,N_30207);
and U33158 (N_33158,N_30822,N_31615);
xnor U33159 (N_33159,N_32380,N_31406);
xor U33160 (N_33160,N_30579,N_31383);
xnor U33161 (N_33161,N_30503,N_30291);
and U33162 (N_33162,N_31816,N_30135);
nand U33163 (N_33163,N_31130,N_30720);
nand U33164 (N_33164,N_31995,N_31519);
nor U33165 (N_33165,N_30233,N_30185);
and U33166 (N_33166,N_32381,N_31138);
xor U33167 (N_33167,N_30918,N_31926);
nor U33168 (N_33168,N_30712,N_32495);
or U33169 (N_33169,N_30734,N_30971);
or U33170 (N_33170,N_30047,N_30702);
nand U33171 (N_33171,N_32396,N_31819);
nor U33172 (N_33172,N_31815,N_31829);
xnor U33173 (N_33173,N_30064,N_30103);
and U33174 (N_33174,N_30435,N_32145);
xor U33175 (N_33175,N_30751,N_30869);
and U33176 (N_33176,N_30062,N_31858);
nor U33177 (N_33177,N_30658,N_30394);
nor U33178 (N_33178,N_32284,N_30930);
nand U33179 (N_33179,N_32493,N_31399);
or U33180 (N_33180,N_31004,N_30672);
or U33181 (N_33181,N_30964,N_30457);
nor U33182 (N_33182,N_31445,N_30642);
nor U33183 (N_33183,N_30508,N_32155);
nor U33184 (N_33184,N_32357,N_30087);
nand U33185 (N_33185,N_30292,N_32021);
nor U33186 (N_33186,N_31173,N_30147);
nor U33187 (N_33187,N_32142,N_32409);
nor U33188 (N_33188,N_32238,N_32322);
xnor U33189 (N_33189,N_31530,N_31697);
nand U33190 (N_33190,N_31252,N_30892);
xnor U33191 (N_33191,N_31103,N_31262);
nand U33192 (N_33192,N_30988,N_32347);
xnor U33193 (N_33193,N_32054,N_30056);
or U33194 (N_33194,N_31598,N_31693);
nor U33195 (N_33195,N_30167,N_30776);
and U33196 (N_33196,N_32010,N_32222);
xnor U33197 (N_33197,N_32043,N_30529);
and U33198 (N_33198,N_30771,N_31341);
or U33199 (N_33199,N_32203,N_30206);
nand U33200 (N_33200,N_30096,N_30669);
nor U33201 (N_33201,N_32169,N_30977);
and U33202 (N_33202,N_30240,N_31939);
nand U33203 (N_33203,N_31376,N_31854);
and U33204 (N_33204,N_30863,N_31195);
or U33205 (N_33205,N_30405,N_31181);
or U33206 (N_33206,N_30688,N_31219);
nor U33207 (N_33207,N_30482,N_31525);
xor U33208 (N_33208,N_31256,N_30174);
nor U33209 (N_33209,N_31496,N_31664);
nor U33210 (N_33210,N_30155,N_30072);
nor U33211 (N_33211,N_32049,N_31187);
xor U33212 (N_33212,N_31622,N_30564);
nor U33213 (N_33213,N_32149,N_31206);
nor U33214 (N_33214,N_32011,N_30716);
nand U33215 (N_33215,N_32275,N_31638);
or U33216 (N_33216,N_32175,N_32253);
and U33217 (N_33217,N_31875,N_30446);
nand U33218 (N_33218,N_31227,N_30120);
and U33219 (N_33219,N_30910,N_30137);
xnor U33220 (N_33220,N_30335,N_30231);
xor U33221 (N_33221,N_30212,N_32084);
nand U33222 (N_33222,N_32220,N_31655);
xor U33223 (N_33223,N_30156,N_31196);
xor U33224 (N_33224,N_30525,N_32489);
or U33225 (N_33225,N_32287,N_31763);
or U33226 (N_33226,N_31924,N_30788);
or U33227 (N_33227,N_30023,N_32144);
xor U33228 (N_33228,N_32302,N_30754);
and U33229 (N_33229,N_30079,N_30625);
or U33230 (N_33230,N_30748,N_30065);
nor U33231 (N_33231,N_31005,N_32387);
xnor U33232 (N_33232,N_31243,N_30128);
and U33233 (N_33233,N_32181,N_30762);
nor U33234 (N_33234,N_30066,N_30301);
and U33235 (N_33235,N_31492,N_30724);
nand U33236 (N_33236,N_30857,N_30357);
nor U33237 (N_33237,N_31314,N_32327);
nor U33238 (N_33238,N_32458,N_32277);
and U33239 (N_33239,N_31586,N_31833);
nand U33240 (N_33240,N_31755,N_31797);
xnor U33241 (N_33241,N_31552,N_30456);
nor U33242 (N_33242,N_31670,N_30567);
nor U33243 (N_33243,N_31309,N_31248);
or U33244 (N_33244,N_31260,N_32334);
nor U33245 (N_33245,N_32041,N_30491);
or U33246 (N_33246,N_30151,N_31000);
nor U33247 (N_33247,N_32428,N_31665);
nor U33248 (N_33248,N_30856,N_30109);
xor U33249 (N_33249,N_30420,N_30111);
or U33250 (N_33250,N_31254,N_30718);
xnor U33251 (N_33251,N_30095,N_30884);
xnor U33252 (N_33252,N_30334,N_30042);
xnor U33253 (N_33253,N_32148,N_32440);
and U33254 (N_33254,N_31795,N_30389);
xor U33255 (N_33255,N_31931,N_31349);
nand U33256 (N_33256,N_30654,N_32321);
nand U33257 (N_33257,N_31188,N_31154);
or U33258 (N_33258,N_32407,N_31418);
nor U33259 (N_33259,N_31700,N_32200);
and U33260 (N_33260,N_30436,N_30210);
nand U33261 (N_33261,N_31014,N_30976);
or U33262 (N_33262,N_31966,N_31062);
xor U33263 (N_33263,N_31773,N_30883);
or U33264 (N_33264,N_32214,N_31412);
and U33265 (N_33265,N_30332,N_32248);
and U33266 (N_33266,N_30294,N_31834);
and U33267 (N_33267,N_32328,N_30171);
xor U33268 (N_33268,N_30570,N_30159);
nor U33269 (N_33269,N_31602,N_30346);
and U33270 (N_33270,N_31021,N_31786);
or U33271 (N_33271,N_31190,N_31139);
nor U33272 (N_33272,N_32033,N_32362);
nand U33273 (N_33273,N_32165,N_31200);
xor U33274 (N_33274,N_31510,N_32325);
nor U33275 (N_33275,N_32132,N_31599);
and U33276 (N_33276,N_32427,N_31438);
nor U33277 (N_33277,N_31116,N_31814);
and U33278 (N_33278,N_31189,N_32212);
nor U33279 (N_33279,N_32177,N_32035);
and U33280 (N_33280,N_31691,N_31764);
or U33281 (N_33281,N_31178,N_31523);
and U33282 (N_33282,N_32093,N_32298);
and U33283 (N_33283,N_31948,N_31398);
or U33284 (N_33284,N_31313,N_31780);
xnor U33285 (N_33285,N_31002,N_30124);
nand U33286 (N_33286,N_30355,N_30791);
or U33287 (N_33287,N_31343,N_30890);
and U33288 (N_33288,N_30470,N_32401);
xor U33289 (N_33289,N_31129,N_30471);
nand U33290 (N_33290,N_31973,N_31210);
nand U33291 (N_33291,N_32335,N_31865);
or U33292 (N_33292,N_30238,N_30973);
and U33293 (N_33293,N_31789,N_31322);
and U33294 (N_33294,N_31080,N_31201);
and U33295 (N_33295,N_30487,N_31429);
nor U33296 (N_33296,N_32114,N_30413);
and U33297 (N_33297,N_32082,N_31089);
nor U33298 (N_33298,N_32208,N_32285);
and U33299 (N_33299,N_30550,N_32136);
nand U33300 (N_33300,N_31595,N_31894);
xnor U33301 (N_33301,N_31807,N_30900);
xnor U33302 (N_33302,N_30258,N_31162);
or U33303 (N_33303,N_32187,N_32438);
and U33304 (N_33304,N_31287,N_30388);
nor U33305 (N_33305,N_31929,N_31142);
nand U33306 (N_33306,N_30341,N_32237);
nand U33307 (N_33307,N_31692,N_32436);
nor U33308 (N_33308,N_30237,N_31110);
nand U33309 (N_33309,N_32156,N_30636);
and U33310 (N_33310,N_32469,N_30800);
nand U33311 (N_33311,N_30612,N_30599);
and U33312 (N_33312,N_32343,N_30837);
or U33313 (N_33313,N_30827,N_32024);
and U33314 (N_33314,N_30236,N_32376);
nor U33315 (N_33315,N_32415,N_32382);
and U33316 (N_33316,N_31166,N_32005);
or U33317 (N_33317,N_31974,N_32055);
nor U33318 (N_33318,N_31025,N_31371);
xor U33319 (N_33319,N_30226,N_32412);
or U33320 (N_33320,N_31587,N_31212);
xnor U33321 (N_33321,N_30293,N_32003);
xor U33322 (N_33322,N_30955,N_32249);
nand U33323 (N_33323,N_31548,N_32113);
and U33324 (N_33324,N_30161,N_30667);
nor U33325 (N_33325,N_32306,N_31329);
xnor U33326 (N_33326,N_31194,N_30908);
or U33327 (N_33327,N_32389,N_31253);
and U33328 (N_33328,N_30670,N_31999);
nand U33329 (N_33329,N_31167,N_32340);
or U33330 (N_33330,N_31358,N_31102);
or U33331 (N_33331,N_31346,N_30090);
and U33332 (N_33332,N_31634,N_31979);
nor U33333 (N_33333,N_31172,N_32314);
nand U33334 (N_33334,N_31610,N_32092);
nor U33335 (N_33335,N_31860,N_31920);
xor U33336 (N_33336,N_32110,N_31486);
and U33337 (N_33337,N_31286,N_32217);
nor U33338 (N_33338,N_31674,N_32067);
xnor U33339 (N_33339,N_30944,N_30425);
nor U33340 (N_33340,N_31515,N_32385);
nand U33341 (N_33341,N_32431,N_30020);
nor U33342 (N_33342,N_31613,N_30602);
nor U33343 (N_33343,N_31635,N_31124);
nor U33344 (N_33344,N_32236,N_30852);
nor U33345 (N_33345,N_31152,N_31811);
nor U33346 (N_33346,N_32416,N_31485);
and U33347 (N_33347,N_30260,N_30620);
xnor U33348 (N_33348,N_30216,N_31575);
nor U33349 (N_33349,N_30994,N_30862);
or U33350 (N_33350,N_30033,N_32384);
nand U33351 (N_33351,N_30993,N_30830);
or U33352 (N_33352,N_31736,N_30148);
and U33353 (N_33353,N_32316,N_32264);
nor U33354 (N_33354,N_31508,N_32421);
and U33355 (N_33355,N_30969,N_30524);
nand U33356 (N_33356,N_31696,N_32344);
nand U33357 (N_33357,N_31455,N_31149);
or U33358 (N_33358,N_30136,N_32397);
or U33359 (N_33359,N_31246,N_30943);
nor U33360 (N_33360,N_32439,N_31273);
or U33361 (N_33361,N_32354,N_32247);
and U33362 (N_33362,N_31881,N_30490);
or U33363 (N_33363,N_30689,N_31380);
or U33364 (N_33364,N_32000,N_30563);
or U33365 (N_33365,N_30452,N_32016);
xor U33366 (N_33366,N_32465,N_30158);
xor U33367 (N_33367,N_30328,N_32201);
or U33368 (N_33368,N_30879,N_31108);
or U33369 (N_33369,N_30385,N_31340);
and U33370 (N_33370,N_32170,N_30574);
and U33371 (N_33371,N_32245,N_32274);
nand U33372 (N_33372,N_30990,N_31532);
xor U33373 (N_33373,N_32377,N_30187);
xor U33374 (N_33374,N_32122,N_31267);
xnor U33375 (N_33375,N_31030,N_31908);
or U33376 (N_33376,N_31280,N_30959);
nor U33377 (N_33377,N_32441,N_32226);
nor U33378 (N_33378,N_31491,N_32101);
nor U33379 (N_33379,N_30954,N_31155);
and U33380 (N_33380,N_30081,N_31408);
and U33381 (N_33381,N_30082,N_30464);
and U33382 (N_33382,N_31460,N_31104);
or U33383 (N_33383,N_30244,N_31245);
nor U33384 (N_33384,N_30537,N_31757);
and U33385 (N_33385,N_31936,N_30609);
or U33386 (N_33386,N_32120,N_31473);
xor U33387 (N_33387,N_32266,N_31147);
xor U33388 (N_33388,N_31911,N_31316);
nand U33389 (N_33389,N_30864,N_32139);
xnor U33390 (N_33390,N_31457,N_32064);
or U33391 (N_33391,N_30722,N_30773);
nand U33392 (N_33392,N_32176,N_30926);
and U33393 (N_33393,N_31518,N_30284);
xnor U33394 (N_33394,N_32029,N_30730);
and U33395 (N_33395,N_31302,N_32091);
xor U33396 (N_33396,N_31032,N_31386);
nand U33397 (N_33397,N_31513,N_30015);
and U33398 (N_33398,N_30555,N_30728);
or U33399 (N_33399,N_30424,N_32229);
nor U33400 (N_33400,N_31991,N_32294);
or U33401 (N_33401,N_31631,N_31470);
or U33402 (N_33402,N_30893,N_30551);
nor U33403 (N_33403,N_31558,N_30118);
and U33404 (N_33404,N_30001,N_31977);
and U33405 (N_33405,N_30927,N_30144);
xor U33406 (N_33406,N_30330,N_31720);
nand U33407 (N_33407,N_31946,N_31038);
and U33408 (N_33408,N_31344,N_30948);
or U33409 (N_33409,N_30845,N_30257);
nand U33410 (N_33410,N_32318,N_30188);
and U33411 (N_33411,N_30604,N_30767);
and U33412 (N_33412,N_31708,N_31565);
nand U33413 (N_33413,N_30543,N_30086);
and U33414 (N_33414,N_31606,N_31556);
or U33415 (N_33415,N_30793,N_30589);
xnor U33416 (N_33416,N_30814,N_30004);
xor U33417 (N_33417,N_31568,N_31792);
and U33418 (N_33418,N_32417,N_31356);
nand U33419 (N_33419,N_30364,N_31461);
and U33420 (N_33420,N_31051,N_30513);
and U33421 (N_33421,N_31037,N_30241);
nand U33422 (N_33422,N_32356,N_30024);
or U33423 (N_33423,N_30745,N_30017);
and U33424 (N_33424,N_31682,N_30912);
or U33425 (N_33425,N_30447,N_30521);
and U33426 (N_33426,N_32346,N_31511);
xor U33427 (N_33427,N_32180,N_32058);
and U33428 (N_33428,N_31375,N_32098);
or U33429 (N_33429,N_32317,N_30100);
xor U33430 (N_33430,N_31673,N_31899);
and U33431 (N_33431,N_31274,N_31844);
xor U33432 (N_33432,N_30234,N_31779);
or U33433 (N_33433,N_31421,N_30696);
or U33434 (N_33434,N_32289,N_32008);
xor U33435 (N_33435,N_31683,N_30299);
nand U33436 (N_33436,N_32086,N_32392);
nor U33437 (N_33437,N_30493,N_31077);
and U33438 (N_33438,N_30783,N_31028);
nand U33439 (N_33439,N_30785,N_30009);
and U33440 (N_33440,N_31157,N_31821);
nand U33441 (N_33441,N_30153,N_30044);
nor U33442 (N_33442,N_30439,N_31601);
and U33443 (N_33443,N_30592,N_30421);
or U33444 (N_33444,N_31891,N_31268);
nor U33445 (N_33445,N_30250,N_30398);
xnor U33446 (N_33446,N_31255,N_32348);
nor U33447 (N_33447,N_30014,N_30320);
nor U33448 (N_33448,N_30559,N_31373);
or U33449 (N_33449,N_32313,N_31537);
nor U33450 (N_33450,N_30011,N_30553);
nand U33451 (N_33451,N_30953,N_31434);
nor U33452 (N_33452,N_31938,N_31699);
nor U33453 (N_33453,N_30820,N_30811);
or U33454 (N_33454,N_30054,N_30075);
and U33455 (N_33455,N_31887,N_30719);
nor U33456 (N_33456,N_30489,N_30626);
or U33457 (N_33457,N_32072,N_32282);
xnor U33458 (N_33458,N_30980,N_31333);
xnor U33459 (N_33459,N_30753,N_31447);
xor U33460 (N_33460,N_31468,N_31882);
nor U33461 (N_33461,N_31756,N_31904);
xor U33462 (N_33462,N_30106,N_31321);
nand U33463 (N_33463,N_30683,N_31081);
nand U33464 (N_33464,N_30502,N_31550);
and U33465 (N_33465,N_30998,N_30454);
nor U33466 (N_33466,N_30092,N_31621);
nor U33467 (N_33467,N_31105,N_30204);
and U33468 (N_33468,N_30855,N_32240);
xnor U33469 (N_33469,N_32154,N_32267);
nand U33470 (N_33470,N_30739,N_31538);
nand U33471 (N_33471,N_30251,N_30568);
or U33472 (N_33472,N_32243,N_30674);
nand U33473 (N_33473,N_30975,N_31863);
xnor U33474 (N_33474,N_30239,N_31628);
and U33475 (N_33475,N_31306,N_31912);
nor U33476 (N_33476,N_31850,N_31131);
and U33477 (N_33477,N_31574,N_31824);
nand U33478 (N_33478,N_31502,N_31293);
and U33479 (N_33479,N_31150,N_30203);
and U33480 (N_33480,N_32406,N_32207);
nand U33481 (N_33481,N_30843,N_30099);
nand U33482 (N_33482,N_30583,N_30083);
or U33483 (N_33483,N_30600,N_31758);
nor U33484 (N_33484,N_31043,N_30429);
xor U33485 (N_33485,N_30779,N_30547);
nor U33486 (N_33486,N_32444,N_30277);
xnor U33487 (N_33487,N_31874,N_30593);
xnor U33488 (N_33488,N_30615,N_31008);
or U33489 (N_33489,N_31145,N_30610);
and U33490 (N_33490,N_31061,N_31701);
nand U33491 (N_33491,N_31740,N_30922);
nor U33492 (N_33492,N_31775,N_31837);
and U33493 (N_33493,N_32191,N_31125);
or U33494 (N_33494,N_31292,N_30673);
nor U33495 (N_33495,N_30473,N_31284);
and U33496 (N_33496,N_30983,N_30169);
or U33497 (N_33497,N_32485,N_30060);
xnor U33498 (N_33498,N_30911,N_32147);
and U33499 (N_33499,N_32210,N_31579);
or U33500 (N_33500,N_32076,N_32080);
xnor U33501 (N_33501,N_31112,N_31363);
xnor U33502 (N_33502,N_31547,N_30193);
or U33503 (N_33503,N_30937,N_32309);
xnor U33504 (N_33504,N_32435,N_30224);
nand U33505 (N_33505,N_30500,N_32301);
nand U33506 (N_33506,N_32081,N_31866);
nand U33507 (N_33507,N_32115,N_30780);
and U33508 (N_33508,N_32166,N_30608);
nand U33509 (N_33509,N_31217,N_30651);
and U33510 (N_33510,N_32300,N_31192);
nand U33511 (N_33511,N_31186,N_30348);
or U33512 (N_33512,N_30641,N_31661);
xor U33513 (N_33513,N_31742,N_31589);
or U33514 (N_33514,N_31637,N_31289);
xor U33515 (N_33515,N_31298,N_32461);
and U33516 (N_33516,N_30314,N_32333);
nor U33517 (N_33517,N_31592,N_31903);
or U33518 (N_33518,N_30261,N_30726);
nand U33519 (N_33519,N_31534,N_30222);
nand U33520 (N_33520,N_30640,N_31493);
and U33521 (N_33521,N_31517,N_31826);
nand U33522 (N_33522,N_30836,N_30744);
nor U33523 (N_33523,N_30629,N_31482);
nor U33524 (N_33524,N_31177,N_31776);
nor U33525 (N_33525,N_30038,N_31193);
or U33526 (N_33526,N_31244,N_30962);
nand U33527 (N_33527,N_30010,N_31940);
and U33528 (N_33528,N_31191,N_30647);
nand U33529 (N_33529,N_30974,N_32027);
or U33530 (N_33530,N_31629,N_30499);
or U33531 (N_33531,N_31820,N_30700);
or U33532 (N_33532,N_30963,N_31420);
nand U33533 (N_33533,N_32361,N_31031);
xor U33534 (N_33534,N_32083,N_31905);
or U33535 (N_33535,N_30897,N_31050);
or U33536 (N_33536,N_30854,N_30094);
and U33537 (N_33537,N_32078,N_31944);
and U33538 (N_33538,N_32474,N_31545);
and U33539 (N_33539,N_31680,N_30956);
nor U33540 (N_33540,N_31175,N_31359);
and U33541 (N_33541,N_30721,N_30074);
and U33542 (N_33542,N_30554,N_30327);
xor U33543 (N_33543,N_31413,N_30307);
and U33544 (N_33544,N_30178,N_31478);
and U33545 (N_33545,N_31335,N_32085);
nand U33546 (N_33546,N_31759,N_30019);
or U33547 (N_33547,N_30545,N_32071);
and U33548 (N_33548,N_30652,N_31494);
nor U33549 (N_33549,N_32106,N_30523);
and U33550 (N_33550,N_32369,N_30468);
nor U33551 (N_33551,N_32383,N_30901);
nor U33552 (N_33552,N_32094,N_31367);
xnor U33553 (N_33553,N_32480,N_31975);
or U33554 (N_33554,N_31744,N_30018);
or U33555 (N_33555,N_31171,N_30138);
xor U33556 (N_33556,N_31197,N_31057);
and U33557 (N_33557,N_30479,N_30687);
or U33558 (N_33558,N_30365,N_31949);
nand U33559 (N_33559,N_30851,N_31728);
xor U33560 (N_33560,N_30273,N_31951);
or U33561 (N_33561,N_30578,N_32118);
or U33562 (N_33562,N_31137,N_31561);
xor U33563 (N_33563,N_30316,N_30591);
or U33564 (N_33564,N_30872,N_32390);
or U33565 (N_33565,N_31409,N_30058);
xor U33566 (N_33566,N_30774,N_32403);
xnor U33567 (N_33567,N_31853,N_32056);
nand U33568 (N_33568,N_31886,N_31208);
and U33569 (N_33569,N_31009,N_30215);
nand U33570 (N_33570,N_30358,N_32355);
nor U33571 (N_33571,N_30067,N_30565);
or U33572 (N_33572,N_31231,N_30795);
or U33573 (N_33573,N_30596,N_30643);
xor U33574 (N_33574,N_32150,N_30818);
and U33575 (N_33575,N_31933,N_32491);
and U33576 (N_33576,N_31753,N_31952);
xor U33577 (N_33577,N_30735,N_30766);
nand U33578 (N_33578,N_32242,N_32244);
nor U33579 (N_33579,N_31588,N_30790);
nand U33580 (N_33580,N_31772,N_30841);
nor U33581 (N_33581,N_30269,N_31016);
nor U33582 (N_33582,N_31067,N_31873);
xnor U33583 (N_33583,N_30282,N_32171);
or U33584 (N_33584,N_30243,N_31533);
and U33585 (N_33585,N_30288,N_30141);
nor U33586 (N_33586,N_31657,N_30150);
xnor U33587 (N_33587,N_31836,N_30713);
nand U33588 (N_33588,N_32077,N_31859);
nand U33589 (N_33589,N_30146,N_30919);
nor U33590 (N_33590,N_31076,N_31288);
and U33591 (N_33591,N_32467,N_32312);
and U33592 (N_33592,N_32233,N_30166);
nor U33593 (N_33593,N_30194,N_31290);
or U33594 (N_33594,N_31368,N_30108);
nor U33595 (N_33595,N_31055,N_32492);
nor U33596 (N_33596,N_32070,N_31164);
xnor U33597 (N_33597,N_31263,N_30782);
nand U33598 (N_33598,N_31159,N_31767);
xor U33599 (N_33599,N_30631,N_31630);
and U33600 (N_33600,N_30397,N_31315);
and U33601 (N_33601,N_30266,N_32051);
nand U33602 (N_33602,N_31390,N_31270);
nor U33603 (N_33603,N_31332,N_30996);
and U33604 (N_33604,N_31725,N_31059);
xor U33605 (N_33605,N_31790,N_31747);
or U33606 (N_33606,N_30684,N_30870);
nand U33607 (N_33607,N_32235,N_32213);
nor U33608 (N_33608,N_30112,N_31845);
nand U33609 (N_33609,N_30697,N_32216);
or U33610 (N_33610,N_31724,N_30275);
or U33611 (N_33611,N_31281,N_31374);
or U33612 (N_33612,N_30130,N_30692);
nand U33613 (N_33613,N_31562,N_30690);
or U33614 (N_33614,N_31169,N_32209);
xor U33615 (N_33615,N_30343,N_31214);
nand U33616 (N_33616,N_30375,N_30182);
nand U33617 (N_33617,N_30129,N_30557);
nor U33618 (N_33618,N_32323,N_30749);
or U33619 (N_33619,N_32254,N_31632);
xor U33620 (N_33620,N_32463,N_31345);
xor U33621 (N_33621,N_32414,N_30409);
nor U33622 (N_33622,N_30992,N_31526);
nor U33623 (N_33623,N_30875,N_31841);
and U33624 (N_33624,N_32296,N_32088);
or U33625 (N_33625,N_30635,N_31745);
nand U33626 (N_33626,N_31918,N_31808);
or U33627 (N_33627,N_30442,N_30984);
and U33628 (N_33628,N_31354,N_32351);
and U33629 (N_33629,N_31086,N_32464);
nor U33630 (N_33630,N_30303,N_30318);
nand U33631 (N_33631,N_31381,N_31113);
nand U33632 (N_33632,N_30057,N_30451);
or U33633 (N_33633,N_32063,N_31989);
or U33634 (N_33634,N_32446,N_30909);
xor U33635 (N_33635,N_32047,N_30428);
xor U33636 (N_33636,N_31644,N_31134);
nand U33637 (N_33637,N_32022,N_30101);
and U33638 (N_33638,N_31988,N_30205);
xnor U33639 (N_33639,N_31746,N_31250);
and U33640 (N_33640,N_30184,N_30657);
nor U33641 (N_33641,N_30709,N_30304);
or U33642 (N_33642,N_30077,N_31411);
or U33643 (N_33643,N_30227,N_32231);
xnor U33644 (N_33644,N_32447,N_30891);
xor U33645 (N_33645,N_31498,N_31296);
nor U33646 (N_33646,N_31889,N_30186);
nand U33647 (N_33647,N_30806,N_31264);
and U33648 (N_33648,N_32460,N_32185);
nor U33649 (N_33649,N_30177,N_31620);
xnor U33650 (N_33650,N_30384,N_30267);
xor U33651 (N_33651,N_32138,N_30941);
xnor U33652 (N_33652,N_31230,N_31458);
nor U33653 (N_33653,N_30211,N_30061);
nand U33654 (N_33654,N_30218,N_30336);
nand U33655 (N_33655,N_31388,N_30832);
or U33656 (N_33656,N_30462,N_31847);
xor U33657 (N_33657,N_31594,N_30794);
and U33658 (N_33658,N_32025,N_31352);
nor U33659 (N_33659,N_30165,N_30406);
and U33660 (N_33660,N_30116,N_32352);
and U33661 (N_33661,N_30438,N_31546);
nand U33662 (N_33662,N_31642,N_30997);
and U33663 (N_33663,N_30538,N_30758);
xor U33664 (N_33664,N_32129,N_30517);
xnor U33665 (N_33665,N_30415,N_32105);
or U33666 (N_33666,N_30552,N_31107);
xnor U33667 (N_33667,N_30157,N_31035);
and U33668 (N_33668,N_31151,N_31799);
and U33669 (N_33669,N_31168,N_30823);
and U33670 (N_33670,N_30655,N_32276);
and U33671 (N_33671,N_31415,N_30765);
nand U33672 (N_33672,N_31572,N_31144);
nand U33673 (N_33673,N_30787,N_31852);
nand U33674 (N_33674,N_31204,N_31733);
nor U33675 (N_33675,N_31570,N_32479);
nand U33676 (N_33676,N_30492,N_30929);
nor U33677 (N_33677,N_30396,N_31068);
and U33678 (N_33678,N_32260,N_32096);
nor U33679 (N_33679,N_31827,N_31422);
and U33680 (N_33680,N_32363,N_30682);
xor U33681 (N_33681,N_31769,N_32001);
or U33682 (N_33682,N_32413,N_31123);
nand U33683 (N_33683,N_31402,N_31348);
or U33684 (N_33684,N_30125,N_30661);
nand U33685 (N_33685,N_31947,N_30308);
nor U33686 (N_33686,N_30542,N_31119);
nor U33687 (N_33687,N_31679,N_32437);
and U33688 (N_33688,N_31793,N_32178);
xor U33689 (N_33689,N_30526,N_31095);
and U33690 (N_33690,N_30584,N_30088);
nand U33691 (N_33691,N_30660,N_30360);
nand U33692 (N_33692,N_31711,N_31963);
nand U33693 (N_33693,N_30369,N_32290);
or U33694 (N_33694,N_31694,N_32332);
xnor U33695 (N_33695,N_32159,N_32272);
nor U33696 (N_33696,N_30132,N_31803);
and U33697 (N_33697,N_30649,N_30048);
and U33698 (N_33698,N_30173,N_31211);
xor U33699 (N_33699,N_31361,N_30639);
nand U33700 (N_33700,N_30463,N_30091);
and U33701 (N_33701,N_30052,N_32293);
or U33702 (N_33702,N_30431,N_32379);
nand U33703 (N_33703,N_32127,N_31251);
or U33704 (N_33704,N_30402,N_31540);
and U33705 (N_33705,N_30022,N_30913);
nor U33706 (N_33706,N_31954,N_30561);
or U33707 (N_33707,N_31512,N_31983);
xor U33708 (N_33708,N_30296,N_30562);
and U33709 (N_33709,N_31749,N_31719);
and U33710 (N_33710,N_31520,N_31608);
nor U33711 (N_33711,N_30936,N_31897);
or U33712 (N_33712,N_30440,N_30810);
nand U33713 (N_33713,N_30575,N_30933);
xnor U33714 (N_33714,N_30045,N_32255);
xor U33715 (N_33715,N_30362,N_31921);
nor U33716 (N_33716,N_30191,N_32295);
nand U33717 (N_33717,N_32017,N_32034);
nand U33718 (N_33718,N_30367,N_31695);
nor U33719 (N_33719,N_32459,N_31160);
and U33720 (N_33720,N_30799,N_30585);
nor U33721 (N_33721,N_31259,N_30531);
or U33722 (N_33722,N_32039,N_30123);
and U33723 (N_33723,N_31121,N_30768);
nor U33724 (N_33724,N_32482,N_31794);
and U33725 (N_33725,N_30315,N_30376);
nor U33726 (N_33726,N_30509,N_31387);
and U33727 (N_33727,N_31563,N_31902);
and U33728 (N_33728,N_32451,N_30544);
and U33729 (N_33729,N_32336,N_30154);
or U33730 (N_33730,N_30180,N_30098);
and U33731 (N_33731,N_32337,N_31265);
xor U33732 (N_33732,N_31033,N_30598);
nor U33733 (N_33733,N_30646,N_31662);
and U33734 (N_33734,N_32408,N_31424);
nand U33735 (N_33735,N_30007,N_30422);
xnor U33736 (N_33736,N_30432,N_30736);
and U33737 (N_33737,N_31925,N_31919);
nand U33738 (N_33738,N_31064,N_30324);
nand U33739 (N_33739,N_30410,N_30485);
or U33740 (N_33740,N_31714,N_30256);
nor U33741 (N_33741,N_30614,N_32250);
nand U33742 (N_33742,N_30906,N_31957);
or U33743 (N_33743,N_30772,N_32194);
and U33744 (N_33744,N_31648,N_31318);
or U33745 (N_33745,N_31739,N_31607);
or U33746 (N_33746,N_31257,N_31489);
and U33747 (N_33747,N_31688,N_31384);
or U33748 (N_33748,N_32452,N_32199);
or U33749 (N_33749,N_32304,N_30645);
xnor U33750 (N_33750,N_30362,N_31029);
or U33751 (N_33751,N_32162,N_30433);
nor U33752 (N_33752,N_31763,N_31927);
nand U33753 (N_33753,N_31634,N_30777);
nor U33754 (N_33754,N_30985,N_30022);
nor U33755 (N_33755,N_31680,N_31343);
or U33756 (N_33756,N_30728,N_31042);
nand U33757 (N_33757,N_31757,N_30849);
xnor U33758 (N_33758,N_32141,N_30099);
or U33759 (N_33759,N_31938,N_31393);
or U33760 (N_33760,N_32125,N_32242);
and U33761 (N_33761,N_32026,N_30741);
or U33762 (N_33762,N_30970,N_30745);
or U33763 (N_33763,N_30371,N_31298);
and U33764 (N_33764,N_32202,N_30578);
nand U33765 (N_33765,N_30947,N_31943);
xnor U33766 (N_33766,N_30462,N_32045);
or U33767 (N_33767,N_32185,N_32150);
nor U33768 (N_33768,N_32156,N_32326);
nand U33769 (N_33769,N_30495,N_31806);
nand U33770 (N_33770,N_30414,N_30760);
nor U33771 (N_33771,N_30012,N_31202);
and U33772 (N_33772,N_30045,N_30472);
nor U33773 (N_33773,N_31788,N_32428);
xor U33774 (N_33774,N_32032,N_32088);
and U33775 (N_33775,N_31271,N_32211);
nor U33776 (N_33776,N_31702,N_32440);
xnor U33777 (N_33777,N_32104,N_30405);
and U33778 (N_33778,N_31390,N_30190);
nor U33779 (N_33779,N_32423,N_31980);
or U33780 (N_33780,N_31003,N_30634);
nor U33781 (N_33781,N_32483,N_30854);
or U33782 (N_33782,N_30095,N_31057);
or U33783 (N_33783,N_32060,N_32045);
nor U33784 (N_33784,N_30692,N_31102);
xnor U33785 (N_33785,N_30660,N_31383);
or U33786 (N_33786,N_31360,N_31462);
or U33787 (N_33787,N_30642,N_32371);
nor U33788 (N_33788,N_30095,N_31075);
or U33789 (N_33789,N_31654,N_30975);
nand U33790 (N_33790,N_30144,N_31275);
or U33791 (N_33791,N_31864,N_31738);
nor U33792 (N_33792,N_30547,N_30007);
nand U33793 (N_33793,N_30448,N_31501);
and U33794 (N_33794,N_31941,N_32061);
nand U33795 (N_33795,N_30986,N_30708);
nand U33796 (N_33796,N_32348,N_32448);
or U33797 (N_33797,N_30246,N_30911);
xor U33798 (N_33798,N_31086,N_30015);
nand U33799 (N_33799,N_31766,N_30618);
or U33800 (N_33800,N_31440,N_30020);
or U33801 (N_33801,N_32003,N_30583);
nor U33802 (N_33802,N_32249,N_31198);
or U33803 (N_33803,N_31258,N_30049);
nand U33804 (N_33804,N_32494,N_30490);
xnor U33805 (N_33805,N_30375,N_31167);
nand U33806 (N_33806,N_32474,N_31752);
nor U33807 (N_33807,N_32119,N_31022);
or U33808 (N_33808,N_30338,N_31547);
xor U33809 (N_33809,N_30277,N_30576);
nor U33810 (N_33810,N_30853,N_31259);
nor U33811 (N_33811,N_30983,N_31545);
nand U33812 (N_33812,N_31482,N_31739);
or U33813 (N_33813,N_31778,N_31342);
and U33814 (N_33814,N_31279,N_30179);
nand U33815 (N_33815,N_31150,N_30868);
nand U33816 (N_33816,N_30790,N_31257);
nand U33817 (N_33817,N_32297,N_31116);
and U33818 (N_33818,N_30963,N_30330);
nand U33819 (N_33819,N_31874,N_32410);
nor U33820 (N_33820,N_30854,N_32460);
nor U33821 (N_33821,N_30025,N_30539);
and U33822 (N_33822,N_32222,N_30704);
or U33823 (N_33823,N_31057,N_31326);
xnor U33824 (N_33824,N_31744,N_31620);
and U33825 (N_33825,N_30485,N_30929);
xor U33826 (N_33826,N_30530,N_32392);
or U33827 (N_33827,N_32274,N_31038);
or U33828 (N_33828,N_31965,N_30234);
nor U33829 (N_33829,N_30368,N_32194);
nand U33830 (N_33830,N_30095,N_31346);
and U33831 (N_33831,N_30097,N_32289);
nand U33832 (N_33832,N_30104,N_30912);
nor U33833 (N_33833,N_30128,N_31010);
nor U33834 (N_33834,N_30361,N_30074);
or U33835 (N_33835,N_32297,N_30111);
nand U33836 (N_33836,N_31928,N_30796);
nor U33837 (N_33837,N_31490,N_30252);
or U33838 (N_33838,N_30815,N_30895);
nand U33839 (N_33839,N_32051,N_30634);
xnor U33840 (N_33840,N_31984,N_30542);
or U33841 (N_33841,N_30257,N_31261);
nor U33842 (N_33842,N_32078,N_30448);
or U33843 (N_33843,N_32107,N_30910);
and U33844 (N_33844,N_30170,N_30710);
or U33845 (N_33845,N_31891,N_31543);
xnor U33846 (N_33846,N_30403,N_30686);
or U33847 (N_33847,N_32249,N_32093);
xnor U33848 (N_33848,N_30726,N_31573);
and U33849 (N_33849,N_30992,N_30550);
and U33850 (N_33850,N_31171,N_30009);
nand U33851 (N_33851,N_31830,N_30974);
xor U33852 (N_33852,N_30715,N_31567);
nor U33853 (N_33853,N_30582,N_31804);
and U33854 (N_33854,N_31394,N_32199);
and U33855 (N_33855,N_31955,N_30947);
and U33856 (N_33856,N_31052,N_32294);
or U33857 (N_33857,N_31758,N_32298);
and U33858 (N_33858,N_31321,N_31290);
or U33859 (N_33859,N_32435,N_31996);
and U33860 (N_33860,N_31226,N_30307);
xor U33861 (N_33861,N_31910,N_30433);
xnor U33862 (N_33862,N_30212,N_30697);
or U33863 (N_33863,N_30677,N_30019);
or U33864 (N_33864,N_30547,N_32477);
nor U33865 (N_33865,N_30065,N_31087);
and U33866 (N_33866,N_30962,N_31024);
or U33867 (N_33867,N_32494,N_30297);
nor U33868 (N_33868,N_30427,N_30106);
xor U33869 (N_33869,N_31014,N_32113);
xnor U33870 (N_33870,N_32035,N_30725);
nand U33871 (N_33871,N_32136,N_32341);
or U33872 (N_33872,N_32154,N_30183);
xnor U33873 (N_33873,N_30579,N_30959);
and U33874 (N_33874,N_30856,N_32137);
nand U33875 (N_33875,N_31521,N_30930);
and U33876 (N_33876,N_32000,N_30363);
nor U33877 (N_33877,N_31888,N_31856);
and U33878 (N_33878,N_31338,N_30041);
nand U33879 (N_33879,N_30805,N_32404);
xnor U33880 (N_33880,N_31800,N_30549);
or U33881 (N_33881,N_32306,N_31481);
and U33882 (N_33882,N_30791,N_31480);
nor U33883 (N_33883,N_30625,N_32179);
xnor U33884 (N_33884,N_31067,N_32449);
and U33885 (N_33885,N_30513,N_32373);
nor U33886 (N_33886,N_30988,N_30270);
and U33887 (N_33887,N_32267,N_31814);
or U33888 (N_33888,N_31064,N_30257);
or U33889 (N_33889,N_32434,N_32155);
nor U33890 (N_33890,N_31055,N_31172);
nand U33891 (N_33891,N_30360,N_31582);
nand U33892 (N_33892,N_31980,N_30110);
xor U33893 (N_33893,N_30540,N_31170);
nand U33894 (N_33894,N_30270,N_30711);
and U33895 (N_33895,N_31737,N_32438);
nor U33896 (N_33896,N_30734,N_31391);
or U33897 (N_33897,N_31298,N_30177);
nand U33898 (N_33898,N_30622,N_31875);
and U33899 (N_33899,N_30430,N_30957);
or U33900 (N_33900,N_31126,N_31714);
and U33901 (N_33901,N_31782,N_32291);
nand U33902 (N_33902,N_30727,N_31124);
nor U33903 (N_33903,N_30731,N_32213);
nor U33904 (N_33904,N_30541,N_32118);
xnor U33905 (N_33905,N_31486,N_31573);
nand U33906 (N_33906,N_30141,N_32045);
and U33907 (N_33907,N_31047,N_31533);
nand U33908 (N_33908,N_30134,N_30067);
nor U33909 (N_33909,N_31972,N_30556);
xor U33910 (N_33910,N_31578,N_30991);
nand U33911 (N_33911,N_30655,N_32430);
xor U33912 (N_33912,N_31362,N_31668);
or U33913 (N_33913,N_32076,N_31113);
xor U33914 (N_33914,N_30729,N_30079);
or U33915 (N_33915,N_32276,N_31325);
and U33916 (N_33916,N_31968,N_30041);
or U33917 (N_33917,N_30164,N_31504);
nor U33918 (N_33918,N_30394,N_31957);
nor U33919 (N_33919,N_30963,N_31796);
or U33920 (N_33920,N_31613,N_31867);
or U33921 (N_33921,N_31858,N_32105);
nand U33922 (N_33922,N_30760,N_31540);
nand U33923 (N_33923,N_30847,N_32247);
nand U33924 (N_33924,N_30964,N_31433);
or U33925 (N_33925,N_30046,N_31791);
and U33926 (N_33926,N_30176,N_30282);
nor U33927 (N_33927,N_31693,N_30975);
nand U33928 (N_33928,N_30249,N_32078);
and U33929 (N_33929,N_31975,N_30975);
nand U33930 (N_33930,N_31289,N_31794);
nand U33931 (N_33931,N_30118,N_32133);
and U33932 (N_33932,N_30668,N_32447);
and U33933 (N_33933,N_30392,N_30218);
nand U33934 (N_33934,N_30636,N_31016);
nor U33935 (N_33935,N_30581,N_31339);
and U33936 (N_33936,N_31464,N_31364);
or U33937 (N_33937,N_31506,N_31963);
or U33938 (N_33938,N_30872,N_31690);
and U33939 (N_33939,N_31081,N_30824);
nand U33940 (N_33940,N_32404,N_30740);
or U33941 (N_33941,N_32347,N_31956);
and U33942 (N_33942,N_31504,N_32459);
xor U33943 (N_33943,N_32243,N_30404);
xnor U33944 (N_33944,N_31522,N_30813);
xor U33945 (N_33945,N_31686,N_31633);
nor U33946 (N_33946,N_30452,N_31785);
xnor U33947 (N_33947,N_30076,N_31343);
xor U33948 (N_33948,N_31971,N_30373);
or U33949 (N_33949,N_31157,N_30603);
nor U33950 (N_33950,N_30911,N_31466);
nor U33951 (N_33951,N_30972,N_31519);
xnor U33952 (N_33952,N_30516,N_30316);
xor U33953 (N_33953,N_31781,N_30586);
nor U33954 (N_33954,N_32046,N_30776);
nand U33955 (N_33955,N_30128,N_31140);
nand U33956 (N_33956,N_31316,N_30083);
nand U33957 (N_33957,N_32181,N_30644);
nand U33958 (N_33958,N_30999,N_30725);
nor U33959 (N_33959,N_30022,N_30659);
and U33960 (N_33960,N_32348,N_30906);
and U33961 (N_33961,N_30385,N_31618);
and U33962 (N_33962,N_30412,N_31490);
xnor U33963 (N_33963,N_32494,N_30537);
and U33964 (N_33964,N_31391,N_31059);
xnor U33965 (N_33965,N_30612,N_30583);
and U33966 (N_33966,N_31822,N_30197);
and U33967 (N_33967,N_31716,N_30170);
nand U33968 (N_33968,N_31842,N_32305);
nor U33969 (N_33969,N_31631,N_30949);
nor U33970 (N_33970,N_31392,N_31573);
nand U33971 (N_33971,N_31520,N_31834);
xor U33972 (N_33972,N_32083,N_30301);
and U33973 (N_33973,N_32215,N_32294);
and U33974 (N_33974,N_30986,N_31754);
nor U33975 (N_33975,N_30907,N_31448);
nor U33976 (N_33976,N_30291,N_32266);
and U33977 (N_33977,N_30029,N_31538);
or U33978 (N_33978,N_30275,N_31918);
xor U33979 (N_33979,N_31540,N_32466);
xnor U33980 (N_33980,N_32027,N_30142);
xor U33981 (N_33981,N_30897,N_30448);
or U33982 (N_33982,N_31836,N_32180);
or U33983 (N_33983,N_32009,N_30657);
or U33984 (N_33984,N_30451,N_30635);
nor U33985 (N_33985,N_31226,N_30240);
xor U33986 (N_33986,N_31329,N_31800);
nand U33987 (N_33987,N_32414,N_31449);
and U33988 (N_33988,N_32292,N_31828);
xnor U33989 (N_33989,N_30609,N_32046);
or U33990 (N_33990,N_31895,N_30557);
or U33991 (N_33991,N_30117,N_30455);
or U33992 (N_33992,N_30599,N_31725);
and U33993 (N_33993,N_31879,N_31153);
nor U33994 (N_33994,N_31869,N_30639);
nand U33995 (N_33995,N_31454,N_30120);
xor U33996 (N_33996,N_30309,N_31574);
xnor U33997 (N_33997,N_31192,N_30424);
or U33998 (N_33998,N_31089,N_32192);
or U33999 (N_33999,N_32228,N_30787);
nor U34000 (N_34000,N_32036,N_31374);
xnor U34001 (N_34001,N_31815,N_31727);
or U34002 (N_34002,N_30517,N_31508);
or U34003 (N_34003,N_32476,N_31189);
or U34004 (N_34004,N_32001,N_30056);
xnor U34005 (N_34005,N_30894,N_31756);
xor U34006 (N_34006,N_30890,N_30576);
and U34007 (N_34007,N_32409,N_30821);
nand U34008 (N_34008,N_30995,N_30919);
xor U34009 (N_34009,N_30652,N_32272);
nand U34010 (N_34010,N_30170,N_32360);
and U34011 (N_34011,N_30048,N_32488);
nand U34012 (N_34012,N_32228,N_31177);
xor U34013 (N_34013,N_30594,N_31327);
or U34014 (N_34014,N_32192,N_31110);
nand U34015 (N_34015,N_31149,N_31093);
xor U34016 (N_34016,N_32369,N_30507);
nand U34017 (N_34017,N_31740,N_31183);
xor U34018 (N_34018,N_31798,N_31989);
xnor U34019 (N_34019,N_31798,N_30680);
and U34020 (N_34020,N_30170,N_31520);
or U34021 (N_34021,N_32180,N_31564);
or U34022 (N_34022,N_31311,N_31006);
or U34023 (N_34023,N_31954,N_32087);
and U34024 (N_34024,N_30662,N_32315);
or U34025 (N_34025,N_31474,N_31814);
xnor U34026 (N_34026,N_31059,N_32455);
and U34027 (N_34027,N_31213,N_31082);
and U34028 (N_34028,N_31851,N_32368);
nand U34029 (N_34029,N_31315,N_32227);
and U34030 (N_34030,N_30957,N_31426);
and U34031 (N_34031,N_30916,N_30288);
and U34032 (N_34032,N_30138,N_31985);
nand U34033 (N_34033,N_30912,N_32134);
xor U34034 (N_34034,N_31895,N_30766);
and U34035 (N_34035,N_30850,N_32278);
or U34036 (N_34036,N_31093,N_30715);
or U34037 (N_34037,N_30587,N_30394);
nand U34038 (N_34038,N_30697,N_32160);
nor U34039 (N_34039,N_31820,N_32179);
nor U34040 (N_34040,N_32197,N_32467);
nor U34041 (N_34041,N_31159,N_31510);
xnor U34042 (N_34042,N_32098,N_30757);
or U34043 (N_34043,N_31336,N_31003);
or U34044 (N_34044,N_31338,N_31829);
nand U34045 (N_34045,N_31039,N_31466);
xor U34046 (N_34046,N_32437,N_31288);
or U34047 (N_34047,N_31653,N_31884);
nor U34048 (N_34048,N_32350,N_30557);
and U34049 (N_34049,N_30059,N_31412);
nand U34050 (N_34050,N_30550,N_31399);
xor U34051 (N_34051,N_30283,N_31970);
xor U34052 (N_34052,N_30832,N_31438);
nor U34053 (N_34053,N_30964,N_31219);
nand U34054 (N_34054,N_32137,N_30877);
or U34055 (N_34055,N_30312,N_31238);
and U34056 (N_34056,N_30644,N_31161);
nor U34057 (N_34057,N_30348,N_32161);
and U34058 (N_34058,N_32024,N_30985);
nand U34059 (N_34059,N_31225,N_31790);
nand U34060 (N_34060,N_30603,N_31649);
nor U34061 (N_34061,N_30172,N_31549);
nor U34062 (N_34062,N_30599,N_31775);
xor U34063 (N_34063,N_30672,N_32231);
and U34064 (N_34064,N_31842,N_32158);
nand U34065 (N_34065,N_30376,N_31832);
xor U34066 (N_34066,N_32301,N_30736);
or U34067 (N_34067,N_32343,N_30817);
nand U34068 (N_34068,N_31320,N_31178);
nor U34069 (N_34069,N_30316,N_32374);
xnor U34070 (N_34070,N_31738,N_31134);
nor U34071 (N_34071,N_30296,N_30062);
nand U34072 (N_34072,N_32004,N_30740);
nand U34073 (N_34073,N_32144,N_31967);
xnor U34074 (N_34074,N_30937,N_30457);
or U34075 (N_34075,N_30200,N_31993);
nor U34076 (N_34076,N_31377,N_31019);
nand U34077 (N_34077,N_31656,N_31350);
xnor U34078 (N_34078,N_30964,N_31062);
xnor U34079 (N_34079,N_32465,N_31016);
and U34080 (N_34080,N_31823,N_32457);
nand U34081 (N_34081,N_30312,N_32477);
nand U34082 (N_34082,N_32363,N_31165);
xor U34083 (N_34083,N_32213,N_31666);
nand U34084 (N_34084,N_30333,N_30342);
xnor U34085 (N_34085,N_30496,N_31057);
and U34086 (N_34086,N_30807,N_31550);
or U34087 (N_34087,N_31783,N_31403);
or U34088 (N_34088,N_31106,N_30316);
xnor U34089 (N_34089,N_30850,N_31345);
nand U34090 (N_34090,N_31532,N_30753);
and U34091 (N_34091,N_30808,N_31378);
xor U34092 (N_34092,N_32024,N_31912);
nor U34093 (N_34093,N_32252,N_30755);
and U34094 (N_34094,N_30185,N_31044);
or U34095 (N_34095,N_31251,N_31230);
or U34096 (N_34096,N_31962,N_31017);
or U34097 (N_34097,N_30946,N_31344);
nand U34098 (N_34098,N_30801,N_30055);
nand U34099 (N_34099,N_32214,N_31142);
nand U34100 (N_34100,N_30641,N_30872);
xor U34101 (N_34101,N_31949,N_30232);
and U34102 (N_34102,N_30953,N_31066);
and U34103 (N_34103,N_32494,N_30262);
xor U34104 (N_34104,N_30635,N_32055);
xnor U34105 (N_34105,N_32372,N_30559);
nor U34106 (N_34106,N_30034,N_30954);
or U34107 (N_34107,N_31030,N_30744);
nor U34108 (N_34108,N_32031,N_31975);
and U34109 (N_34109,N_32267,N_31697);
and U34110 (N_34110,N_32181,N_30541);
or U34111 (N_34111,N_31308,N_31820);
or U34112 (N_34112,N_31697,N_30306);
nand U34113 (N_34113,N_32440,N_31139);
nor U34114 (N_34114,N_30928,N_32104);
and U34115 (N_34115,N_31465,N_31601);
or U34116 (N_34116,N_31518,N_31423);
xor U34117 (N_34117,N_31873,N_31175);
or U34118 (N_34118,N_31770,N_31267);
and U34119 (N_34119,N_32047,N_30677);
and U34120 (N_34120,N_30781,N_30007);
and U34121 (N_34121,N_31566,N_32278);
nand U34122 (N_34122,N_30407,N_30252);
xnor U34123 (N_34123,N_30852,N_31219);
nor U34124 (N_34124,N_31691,N_31371);
xor U34125 (N_34125,N_30820,N_30065);
and U34126 (N_34126,N_32260,N_32028);
or U34127 (N_34127,N_30108,N_31729);
and U34128 (N_34128,N_30570,N_32326);
nor U34129 (N_34129,N_31865,N_30674);
xnor U34130 (N_34130,N_30327,N_32092);
xnor U34131 (N_34131,N_32307,N_31601);
or U34132 (N_34132,N_31606,N_32064);
and U34133 (N_34133,N_31340,N_32006);
and U34134 (N_34134,N_31579,N_30305);
nor U34135 (N_34135,N_30935,N_30800);
xnor U34136 (N_34136,N_31853,N_30704);
nor U34137 (N_34137,N_30305,N_31527);
or U34138 (N_34138,N_31672,N_30080);
and U34139 (N_34139,N_31635,N_32390);
nand U34140 (N_34140,N_30274,N_31986);
nand U34141 (N_34141,N_32296,N_31897);
or U34142 (N_34142,N_31515,N_30692);
xnor U34143 (N_34143,N_30118,N_31739);
xnor U34144 (N_34144,N_30535,N_31746);
or U34145 (N_34145,N_30493,N_31053);
and U34146 (N_34146,N_30582,N_31060);
and U34147 (N_34147,N_30133,N_30511);
nor U34148 (N_34148,N_31893,N_30809);
xor U34149 (N_34149,N_30654,N_31876);
xnor U34150 (N_34150,N_31669,N_31470);
nor U34151 (N_34151,N_31024,N_30005);
nor U34152 (N_34152,N_30665,N_31294);
nand U34153 (N_34153,N_31599,N_31175);
or U34154 (N_34154,N_30234,N_30072);
or U34155 (N_34155,N_32495,N_30425);
xor U34156 (N_34156,N_32456,N_30224);
or U34157 (N_34157,N_30692,N_30002);
xor U34158 (N_34158,N_31483,N_31926);
nand U34159 (N_34159,N_32311,N_30042);
and U34160 (N_34160,N_31599,N_30903);
nor U34161 (N_34161,N_32339,N_30124);
nor U34162 (N_34162,N_31215,N_30179);
nand U34163 (N_34163,N_30437,N_30126);
and U34164 (N_34164,N_30984,N_31353);
xor U34165 (N_34165,N_32041,N_32435);
and U34166 (N_34166,N_31776,N_31681);
nor U34167 (N_34167,N_31699,N_31780);
nand U34168 (N_34168,N_31171,N_31564);
and U34169 (N_34169,N_30580,N_31017);
nor U34170 (N_34170,N_32409,N_32262);
or U34171 (N_34171,N_31554,N_30950);
nand U34172 (N_34172,N_32494,N_31463);
nor U34173 (N_34173,N_31461,N_31961);
nand U34174 (N_34174,N_32162,N_32260);
nand U34175 (N_34175,N_31121,N_30906);
nor U34176 (N_34176,N_31498,N_31085);
nand U34177 (N_34177,N_30713,N_31149);
or U34178 (N_34178,N_32449,N_31064);
nand U34179 (N_34179,N_30386,N_30023);
or U34180 (N_34180,N_31750,N_30461);
nor U34181 (N_34181,N_31702,N_31831);
nand U34182 (N_34182,N_31672,N_31270);
nand U34183 (N_34183,N_30011,N_31892);
nor U34184 (N_34184,N_32053,N_32178);
nor U34185 (N_34185,N_30722,N_32351);
nor U34186 (N_34186,N_31292,N_32235);
xnor U34187 (N_34187,N_30193,N_31528);
and U34188 (N_34188,N_30583,N_30582);
nor U34189 (N_34189,N_32220,N_30243);
nand U34190 (N_34190,N_30235,N_31974);
nand U34191 (N_34191,N_32187,N_31132);
or U34192 (N_34192,N_30327,N_32361);
xnor U34193 (N_34193,N_31476,N_31813);
xor U34194 (N_34194,N_31513,N_32259);
or U34195 (N_34195,N_31095,N_31864);
nand U34196 (N_34196,N_30163,N_32141);
and U34197 (N_34197,N_30912,N_30824);
or U34198 (N_34198,N_31134,N_31333);
or U34199 (N_34199,N_30126,N_31436);
xnor U34200 (N_34200,N_30482,N_31969);
nand U34201 (N_34201,N_32338,N_30050);
xnor U34202 (N_34202,N_32114,N_32375);
nand U34203 (N_34203,N_31697,N_30824);
and U34204 (N_34204,N_32347,N_30845);
nor U34205 (N_34205,N_30715,N_31742);
or U34206 (N_34206,N_30719,N_30675);
nor U34207 (N_34207,N_31499,N_30871);
and U34208 (N_34208,N_30633,N_32085);
or U34209 (N_34209,N_31576,N_31429);
nand U34210 (N_34210,N_31653,N_30488);
nor U34211 (N_34211,N_30963,N_30041);
nand U34212 (N_34212,N_31632,N_31313);
or U34213 (N_34213,N_32369,N_32485);
or U34214 (N_34214,N_31833,N_30144);
xor U34215 (N_34215,N_31220,N_32452);
xnor U34216 (N_34216,N_32156,N_30094);
xnor U34217 (N_34217,N_32426,N_31283);
or U34218 (N_34218,N_31019,N_32339);
xor U34219 (N_34219,N_32070,N_30693);
nand U34220 (N_34220,N_30235,N_32228);
or U34221 (N_34221,N_31178,N_30016);
and U34222 (N_34222,N_30508,N_31388);
or U34223 (N_34223,N_32205,N_31430);
and U34224 (N_34224,N_30562,N_30973);
xnor U34225 (N_34225,N_32419,N_31557);
or U34226 (N_34226,N_30222,N_32310);
or U34227 (N_34227,N_30724,N_30076);
nand U34228 (N_34228,N_32135,N_30683);
nand U34229 (N_34229,N_30824,N_30072);
and U34230 (N_34230,N_30672,N_32118);
nor U34231 (N_34231,N_30087,N_30165);
xnor U34232 (N_34232,N_31685,N_32121);
nand U34233 (N_34233,N_30271,N_31168);
xor U34234 (N_34234,N_30409,N_30581);
nor U34235 (N_34235,N_32123,N_31864);
and U34236 (N_34236,N_30821,N_31759);
or U34237 (N_34237,N_31017,N_31943);
and U34238 (N_34238,N_31106,N_32078);
nand U34239 (N_34239,N_31157,N_30814);
nor U34240 (N_34240,N_30632,N_32107);
nor U34241 (N_34241,N_31023,N_31410);
or U34242 (N_34242,N_31081,N_31837);
or U34243 (N_34243,N_30693,N_32170);
and U34244 (N_34244,N_31297,N_31744);
and U34245 (N_34245,N_32033,N_31964);
xnor U34246 (N_34246,N_31315,N_30847);
and U34247 (N_34247,N_30291,N_30837);
and U34248 (N_34248,N_31912,N_30010);
xnor U34249 (N_34249,N_32066,N_31827);
nor U34250 (N_34250,N_31380,N_30871);
nand U34251 (N_34251,N_31027,N_30724);
nor U34252 (N_34252,N_31477,N_32030);
nand U34253 (N_34253,N_31614,N_30488);
and U34254 (N_34254,N_31641,N_30081);
nand U34255 (N_34255,N_32455,N_31672);
and U34256 (N_34256,N_32374,N_31751);
xnor U34257 (N_34257,N_32231,N_31283);
nor U34258 (N_34258,N_32308,N_30756);
or U34259 (N_34259,N_30783,N_30721);
or U34260 (N_34260,N_31890,N_30135);
and U34261 (N_34261,N_31987,N_32239);
and U34262 (N_34262,N_31822,N_31548);
nand U34263 (N_34263,N_31687,N_30334);
nor U34264 (N_34264,N_31810,N_31937);
or U34265 (N_34265,N_31604,N_31432);
and U34266 (N_34266,N_31684,N_30980);
or U34267 (N_34267,N_30833,N_31094);
and U34268 (N_34268,N_30770,N_30641);
xor U34269 (N_34269,N_30952,N_30299);
or U34270 (N_34270,N_30860,N_31096);
nand U34271 (N_34271,N_31857,N_32297);
nand U34272 (N_34272,N_30387,N_32189);
xor U34273 (N_34273,N_30250,N_31201);
and U34274 (N_34274,N_31916,N_30139);
nand U34275 (N_34275,N_31240,N_31956);
xnor U34276 (N_34276,N_30592,N_30695);
nor U34277 (N_34277,N_31827,N_31402);
or U34278 (N_34278,N_32127,N_30667);
and U34279 (N_34279,N_32125,N_30330);
xor U34280 (N_34280,N_31649,N_31545);
and U34281 (N_34281,N_30065,N_32100);
or U34282 (N_34282,N_30130,N_31467);
or U34283 (N_34283,N_30811,N_31081);
or U34284 (N_34284,N_30428,N_31728);
or U34285 (N_34285,N_31142,N_32207);
nor U34286 (N_34286,N_31456,N_31621);
nand U34287 (N_34287,N_31230,N_30023);
and U34288 (N_34288,N_32197,N_30180);
xnor U34289 (N_34289,N_31995,N_31855);
or U34290 (N_34290,N_30958,N_31483);
or U34291 (N_34291,N_32127,N_30655);
and U34292 (N_34292,N_30239,N_31623);
nand U34293 (N_34293,N_31841,N_30198);
and U34294 (N_34294,N_32250,N_32342);
nor U34295 (N_34295,N_30445,N_31894);
or U34296 (N_34296,N_31022,N_30570);
xor U34297 (N_34297,N_30894,N_31543);
or U34298 (N_34298,N_30826,N_31812);
nand U34299 (N_34299,N_30712,N_30956);
or U34300 (N_34300,N_31010,N_30724);
and U34301 (N_34301,N_32443,N_30195);
nand U34302 (N_34302,N_31191,N_30345);
nand U34303 (N_34303,N_30593,N_30299);
xor U34304 (N_34304,N_30721,N_32032);
nand U34305 (N_34305,N_30359,N_30093);
and U34306 (N_34306,N_30336,N_32269);
and U34307 (N_34307,N_31622,N_31755);
nor U34308 (N_34308,N_30498,N_31624);
xnor U34309 (N_34309,N_31740,N_30935);
and U34310 (N_34310,N_31658,N_30781);
nand U34311 (N_34311,N_30605,N_31132);
and U34312 (N_34312,N_32074,N_31442);
nor U34313 (N_34313,N_31698,N_30467);
nor U34314 (N_34314,N_31779,N_30655);
and U34315 (N_34315,N_31459,N_30878);
xnor U34316 (N_34316,N_31563,N_31377);
xnor U34317 (N_34317,N_30730,N_32226);
and U34318 (N_34318,N_31521,N_30432);
nand U34319 (N_34319,N_31776,N_31945);
and U34320 (N_34320,N_32493,N_32158);
or U34321 (N_34321,N_31032,N_30491);
xor U34322 (N_34322,N_30158,N_30517);
xnor U34323 (N_34323,N_31945,N_31355);
xnor U34324 (N_34324,N_32304,N_32336);
or U34325 (N_34325,N_31527,N_32173);
and U34326 (N_34326,N_31851,N_30254);
xor U34327 (N_34327,N_32031,N_31567);
xnor U34328 (N_34328,N_30339,N_32172);
nand U34329 (N_34329,N_30612,N_32165);
nor U34330 (N_34330,N_30182,N_31490);
nor U34331 (N_34331,N_30838,N_30503);
nor U34332 (N_34332,N_30075,N_32205);
nor U34333 (N_34333,N_30075,N_31699);
nor U34334 (N_34334,N_31784,N_31347);
or U34335 (N_34335,N_30251,N_30784);
and U34336 (N_34336,N_31051,N_30059);
nor U34337 (N_34337,N_30673,N_32054);
xor U34338 (N_34338,N_32029,N_30318);
and U34339 (N_34339,N_32052,N_31566);
nor U34340 (N_34340,N_31319,N_31439);
xor U34341 (N_34341,N_31978,N_31966);
nor U34342 (N_34342,N_30010,N_30291);
nor U34343 (N_34343,N_31666,N_31484);
nor U34344 (N_34344,N_30003,N_31835);
or U34345 (N_34345,N_30204,N_31992);
and U34346 (N_34346,N_31935,N_31296);
nand U34347 (N_34347,N_30885,N_31649);
or U34348 (N_34348,N_30797,N_31249);
or U34349 (N_34349,N_30106,N_32270);
or U34350 (N_34350,N_31625,N_31125);
or U34351 (N_34351,N_31055,N_31906);
nor U34352 (N_34352,N_31776,N_32336);
nand U34353 (N_34353,N_32044,N_31267);
nand U34354 (N_34354,N_30145,N_30227);
xnor U34355 (N_34355,N_32298,N_32152);
nand U34356 (N_34356,N_31249,N_32325);
nand U34357 (N_34357,N_32490,N_30643);
or U34358 (N_34358,N_30616,N_30292);
xor U34359 (N_34359,N_32319,N_31138);
nor U34360 (N_34360,N_30377,N_30755);
xnor U34361 (N_34361,N_31733,N_30429);
or U34362 (N_34362,N_32168,N_32110);
or U34363 (N_34363,N_31542,N_31193);
or U34364 (N_34364,N_31000,N_30277);
nor U34365 (N_34365,N_30771,N_30268);
nand U34366 (N_34366,N_30884,N_32188);
nand U34367 (N_34367,N_30166,N_32315);
nor U34368 (N_34368,N_30348,N_31703);
and U34369 (N_34369,N_30281,N_30819);
xor U34370 (N_34370,N_31128,N_30282);
xor U34371 (N_34371,N_30286,N_31788);
and U34372 (N_34372,N_30534,N_31425);
nor U34373 (N_34373,N_32087,N_31339);
xor U34374 (N_34374,N_31002,N_31110);
and U34375 (N_34375,N_31388,N_31774);
xnor U34376 (N_34376,N_30984,N_30911);
xnor U34377 (N_34377,N_31224,N_30083);
nand U34378 (N_34378,N_31752,N_31525);
or U34379 (N_34379,N_31524,N_32029);
nor U34380 (N_34380,N_30766,N_31669);
and U34381 (N_34381,N_30692,N_30524);
or U34382 (N_34382,N_31376,N_30700);
and U34383 (N_34383,N_30079,N_31280);
or U34384 (N_34384,N_31082,N_32147);
or U34385 (N_34385,N_30869,N_31957);
nand U34386 (N_34386,N_32053,N_30822);
nor U34387 (N_34387,N_32094,N_30209);
nor U34388 (N_34388,N_32481,N_31762);
or U34389 (N_34389,N_31311,N_31880);
and U34390 (N_34390,N_31402,N_31000);
xor U34391 (N_34391,N_30220,N_31877);
nor U34392 (N_34392,N_31615,N_30919);
and U34393 (N_34393,N_32272,N_30928);
nand U34394 (N_34394,N_31411,N_30274);
or U34395 (N_34395,N_32037,N_30621);
xor U34396 (N_34396,N_31529,N_31546);
or U34397 (N_34397,N_32357,N_30581);
xnor U34398 (N_34398,N_30197,N_32317);
and U34399 (N_34399,N_30595,N_30003);
xnor U34400 (N_34400,N_30783,N_30173);
and U34401 (N_34401,N_31488,N_32158);
xnor U34402 (N_34402,N_31042,N_30510);
nand U34403 (N_34403,N_31555,N_32242);
xor U34404 (N_34404,N_30064,N_31027);
nor U34405 (N_34405,N_31658,N_31435);
xor U34406 (N_34406,N_31893,N_32127);
and U34407 (N_34407,N_31551,N_30716);
nand U34408 (N_34408,N_31251,N_31305);
xnor U34409 (N_34409,N_32024,N_31491);
nor U34410 (N_34410,N_32373,N_31668);
and U34411 (N_34411,N_31425,N_32299);
nor U34412 (N_34412,N_30404,N_30836);
or U34413 (N_34413,N_31712,N_31562);
xnor U34414 (N_34414,N_30435,N_30013);
and U34415 (N_34415,N_30439,N_32054);
nand U34416 (N_34416,N_30980,N_30712);
nand U34417 (N_34417,N_30966,N_31558);
and U34418 (N_34418,N_32495,N_32171);
xor U34419 (N_34419,N_31356,N_31110);
nor U34420 (N_34420,N_30979,N_31420);
or U34421 (N_34421,N_31695,N_32059);
nand U34422 (N_34422,N_31392,N_30073);
and U34423 (N_34423,N_31384,N_32239);
xor U34424 (N_34424,N_31060,N_31672);
nand U34425 (N_34425,N_31527,N_32109);
nor U34426 (N_34426,N_32069,N_30825);
nor U34427 (N_34427,N_31896,N_30148);
and U34428 (N_34428,N_31722,N_31156);
or U34429 (N_34429,N_31195,N_31175);
xor U34430 (N_34430,N_32432,N_30661);
nor U34431 (N_34431,N_30845,N_30819);
and U34432 (N_34432,N_31954,N_30504);
xor U34433 (N_34433,N_32363,N_30676);
and U34434 (N_34434,N_30214,N_32216);
xor U34435 (N_34435,N_30705,N_31565);
or U34436 (N_34436,N_31848,N_32173);
nor U34437 (N_34437,N_31876,N_31781);
nor U34438 (N_34438,N_30210,N_31598);
or U34439 (N_34439,N_30779,N_32302);
or U34440 (N_34440,N_31641,N_31853);
nor U34441 (N_34441,N_30981,N_32315);
and U34442 (N_34442,N_30216,N_30145);
xor U34443 (N_34443,N_31203,N_31900);
or U34444 (N_34444,N_30332,N_30366);
or U34445 (N_34445,N_31658,N_30071);
or U34446 (N_34446,N_31464,N_30512);
xor U34447 (N_34447,N_32322,N_32451);
nand U34448 (N_34448,N_31179,N_30328);
and U34449 (N_34449,N_30057,N_30930);
nand U34450 (N_34450,N_31807,N_31537);
nor U34451 (N_34451,N_31376,N_30009);
xnor U34452 (N_34452,N_31196,N_32053);
or U34453 (N_34453,N_32049,N_32340);
or U34454 (N_34454,N_30309,N_30491);
or U34455 (N_34455,N_31287,N_32353);
and U34456 (N_34456,N_30070,N_31019);
xor U34457 (N_34457,N_30387,N_32321);
or U34458 (N_34458,N_31363,N_31707);
nor U34459 (N_34459,N_30268,N_30387);
nand U34460 (N_34460,N_30023,N_30927);
xnor U34461 (N_34461,N_32237,N_31436);
and U34462 (N_34462,N_31751,N_31002);
nor U34463 (N_34463,N_31910,N_31472);
nor U34464 (N_34464,N_30743,N_32072);
nor U34465 (N_34465,N_31816,N_31996);
xnor U34466 (N_34466,N_31207,N_31622);
nand U34467 (N_34467,N_30381,N_31069);
xor U34468 (N_34468,N_31738,N_30100);
nand U34469 (N_34469,N_30635,N_32259);
xnor U34470 (N_34470,N_30797,N_31434);
or U34471 (N_34471,N_32269,N_30545);
nand U34472 (N_34472,N_31948,N_31676);
xor U34473 (N_34473,N_30596,N_30095);
xor U34474 (N_34474,N_32294,N_31314);
xor U34475 (N_34475,N_31305,N_32386);
nor U34476 (N_34476,N_31583,N_31764);
nand U34477 (N_34477,N_31495,N_31153);
nor U34478 (N_34478,N_30846,N_31014);
nand U34479 (N_34479,N_30241,N_31407);
nor U34480 (N_34480,N_32057,N_31927);
and U34481 (N_34481,N_31280,N_31128);
nand U34482 (N_34482,N_30285,N_30676);
and U34483 (N_34483,N_30641,N_31733);
xor U34484 (N_34484,N_31633,N_31029);
or U34485 (N_34485,N_31253,N_30737);
nand U34486 (N_34486,N_31612,N_31185);
nand U34487 (N_34487,N_30515,N_32361);
and U34488 (N_34488,N_30829,N_31990);
nand U34489 (N_34489,N_30320,N_31305);
and U34490 (N_34490,N_31960,N_31889);
xor U34491 (N_34491,N_30961,N_30266);
nor U34492 (N_34492,N_30263,N_31602);
nor U34493 (N_34493,N_30808,N_32250);
or U34494 (N_34494,N_30395,N_30530);
and U34495 (N_34495,N_30174,N_31942);
nand U34496 (N_34496,N_31449,N_31494);
nor U34497 (N_34497,N_30095,N_32248);
or U34498 (N_34498,N_31835,N_30439);
or U34499 (N_34499,N_31950,N_30705);
and U34500 (N_34500,N_30361,N_31909);
xnor U34501 (N_34501,N_31334,N_31885);
xnor U34502 (N_34502,N_30055,N_31744);
or U34503 (N_34503,N_30347,N_31414);
nand U34504 (N_34504,N_30865,N_32070);
nor U34505 (N_34505,N_32035,N_31209);
and U34506 (N_34506,N_31235,N_32409);
and U34507 (N_34507,N_31471,N_30822);
and U34508 (N_34508,N_30701,N_32318);
and U34509 (N_34509,N_30919,N_31346);
xor U34510 (N_34510,N_32043,N_30688);
nor U34511 (N_34511,N_30195,N_31191);
nor U34512 (N_34512,N_31131,N_30256);
nand U34513 (N_34513,N_31194,N_30885);
or U34514 (N_34514,N_32380,N_31734);
nor U34515 (N_34515,N_31737,N_31128);
or U34516 (N_34516,N_32442,N_31336);
xnor U34517 (N_34517,N_30795,N_32184);
xnor U34518 (N_34518,N_32328,N_30040);
or U34519 (N_34519,N_30136,N_31593);
xnor U34520 (N_34520,N_32462,N_31975);
nand U34521 (N_34521,N_30085,N_32070);
xor U34522 (N_34522,N_30482,N_32135);
and U34523 (N_34523,N_30468,N_31203);
xnor U34524 (N_34524,N_31269,N_32116);
nor U34525 (N_34525,N_31287,N_31341);
xnor U34526 (N_34526,N_30215,N_31671);
nor U34527 (N_34527,N_31317,N_31694);
and U34528 (N_34528,N_31978,N_32257);
xor U34529 (N_34529,N_30712,N_30564);
nor U34530 (N_34530,N_31228,N_32392);
or U34531 (N_34531,N_30940,N_30095);
nand U34532 (N_34532,N_31322,N_31977);
nand U34533 (N_34533,N_30014,N_30704);
nor U34534 (N_34534,N_31325,N_31939);
xor U34535 (N_34535,N_30100,N_30727);
nor U34536 (N_34536,N_31710,N_30779);
xor U34537 (N_34537,N_30857,N_30960);
xnor U34538 (N_34538,N_32442,N_31564);
nand U34539 (N_34539,N_32143,N_30673);
and U34540 (N_34540,N_30357,N_31415);
and U34541 (N_34541,N_32041,N_31284);
and U34542 (N_34542,N_30625,N_32236);
and U34543 (N_34543,N_30516,N_30459);
nor U34544 (N_34544,N_30950,N_30041);
xnor U34545 (N_34545,N_32403,N_32301);
and U34546 (N_34546,N_30876,N_30297);
xnor U34547 (N_34547,N_32163,N_32438);
xor U34548 (N_34548,N_31201,N_30290);
nor U34549 (N_34549,N_31783,N_30494);
xnor U34550 (N_34550,N_30876,N_32140);
nand U34551 (N_34551,N_30346,N_31801);
or U34552 (N_34552,N_30401,N_30806);
nand U34553 (N_34553,N_30257,N_32039);
nor U34554 (N_34554,N_31737,N_31907);
nand U34555 (N_34555,N_30271,N_31127);
nor U34556 (N_34556,N_30655,N_31215);
xor U34557 (N_34557,N_31901,N_32408);
or U34558 (N_34558,N_32038,N_31979);
xnor U34559 (N_34559,N_31492,N_31206);
xor U34560 (N_34560,N_31288,N_30514);
xnor U34561 (N_34561,N_31997,N_30042);
nand U34562 (N_34562,N_30764,N_30539);
nor U34563 (N_34563,N_30851,N_32491);
or U34564 (N_34564,N_30971,N_30362);
nand U34565 (N_34565,N_31546,N_31544);
nand U34566 (N_34566,N_32321,N_30800);
and U34567 (N_34567,N_30506,N_32476);
nand U34568 (N_34568,N_30095,N_31778);
or U34569 (N_34569,N_30322,N_30179);
or U34570 (N_34570,N_30213,N_32178);
xor U34571 (N_34571,N_31647,N_30827);
nand U34572 (N_34572,N_30076,N_30577);
and U34573 (N_34573,N_31701,N_32073);
nor U34574 (N_34574,N_30475,N_31381);
and U34575 (N_34575,N_31989,N_31438);
and U34576 (N_34576,N_31371,N_31710);
or U34577 (N_34577,N_30609,N_32438);
or U34578 (N_34578,N_32224,N_32448);
xor U34579 (N_34579,N_32410,N_31325);
xnor U34580 (N_34580,N_31028,N_30930);
xnor U34581 (N_34581,N_31566,N_30410);
and U34582 (N_34582,N_31572,N_32360);
or U34583 (N_34583,N_31948,N_30865);
or U34584 (N_34584,N_31052,N_30419);
nand U34585 (N_34585,N_31450,N_31433);
and U34586 (N_34586,N_31647,N_31168);
and U34587 (N_34587,N_32226,N_30381);
xor U34588 (N_34588,N_31035,N_31261);
or U34589 (N_34589,N_31397,N_31400);
or U34590 (N_34590,N_32132,N_30504);
nand U34591 (N_34591,N_31662,N_32121);
xnor U34592 (N_34592,N_31269,N_30183);
or U34593 (N_34593,N_30911,N_30555);
and U34594 (N_34594,N_31875,N_30206);
nand U34595 (N_34595,N_30591,N_31046);
nor U34596 (N_34596,N_31102,N_30328);
nor U34597 (N_34597,N_30070,N_31106);
or U34598 (N_34598,N_31797,N_31127);
xor U34599 (N_34599,N_32494,N_30693);
xor U34600 (N_34600,N_32334,N_30502);
xnor U34601 (N_34601,N_31579,N_31795);
or U34602 (N_34602,N_30705,N_31590);
and U34603 (N_34603,N_30977,N_31168);
nand U34604 (N_34604,N_31384,N_32137);
xnor U34605 (N_34605,N_30234,N_31192);
or U34606 (N_34606,N_30459,N_30121);
and U34607 (N_34607,N_30039,N_31276);
or U34608 (N_34608,N_32154,N_30246);
and U34609 (N_34609,N_31650,N_31666);
or U34610 (N_34610,N_31596,N_32342);
or U34611 (N_34611,N_30998,N_30997);
nand U34612 (N_34612,N_30944,N_32435);
nor U34613 (N_34613,N_30012,N_32371);
xor U34614 (N_34614,N_30751,N_30495);
nor U34615 (N_34615,N_31432,N_30932);
nor U34616 (N_34616,N_31647,N_30145);
nor U34617 (N_34617,N_31680,N_30664);
nor U34618 (N_34618,N_32061,N_32206);
nand U34619 (N_34619,N_31739,N_31295);
xnor U34620 (N_34620,N_32268,N_30963);
and U34621 (N_34621,N_31072,N_31130);
and U34622 (N_34622,N_30565,N_30996);
xor U34623 (N_34623,N_32273,N_32009);
xnor U34624 (N_34624,N_30217,N_31568);
and U34625 (N_34625,N_32253,N_32458);
nand U34626 (N_34626,N_30217,N_30985);
and U34627 (N_34627,N_31850,N_30354);
or U34628 (N_34628,N_31768,N_31948);
and U34629 (N_34629,N_30493,N_30367);
nor U34630 (N_34630,N_31575,N_32165);
xor U34631 (N_34631,N_32334,N_31055);
or U34632 (N_34632,N_30751,N_30253);
nor U34633 (N_34633,N_32329,N_32398);
nor U34634 (N_34634,N_32100,N_30668);
nor U34635 (N_34635,N_30436,N_31640);
xor U34636 (N_34636,N_30330,N_32374);
nand U34637 (N_34637,N_30568,N_31637);
xnor U34638 (N_34638,N_30565,N_30591);
nor U34639 (N_34639,N_32170,N_31902);
nand U34640 (N_34640,N_30628,N_30723);
nor U34641 (N_34641,N_30371,N_32200);
nor U34642 (N_34642,N_30179,N_32444);
or U34643 (N_34643,N_32357,N_31346);
or U34644 (N_34644,N_32193,N_31794);
xnor U34645 (N_34645,N_31449,N_30542);
xnor U34646 (N_34646,N_30212,N_31728);
nor U34647 (N_34647,N_30376,N_31648);
xnor U34648 (N_34648,N_31592,N_30563);
nand U34649 (N_34649,N_31157,N_31554);
xor U34650 (N_34650,N_31108,N_30445);
xor U34651 (N_34651,N_31158,N_31605);
and U34652 (N_34652,N_30580,N_30239);
nand U34653 (N_34653,N_31789,N_32357);
or U34654 (N_34654,N_32035,N_31904);
nand U34655 (N_34655,N_31069,N_32484);
xor U34656 (N_34656,N_32319,N_32372);
xor U34657 (N_34657,N_31892,N_30300);
nor U34658 (N_34658,N_31057,N_30905);
nor U34659 (N_34659,N_32295,N_31555);
nor U34660 (N_34660,N_31517,N_32093);
nor U34661 (N_34661,N_30032,N_31629);
xor U34662 (N_34662,N_30017,N_31431);
nor U34663 (N_34663,N_31876,N_31958);
or U34664 (N_34664,N_31243,N_30968);
nor U34665 (N_34665,N_31797,N_30621);
nor U34666 (N_34666,N_32333,N_32234);
nand U34667 (N_34667,N_32468,N_30844);
nor U34668 (N_34668,N_30696,N_31682);
xnor U34669 (N_34669,N_30279,N_30286);
or U34670 (N_34670,N_32034,N_31081);
xor U34671 (N_34671,N_31592,N_31833);
nand U34672 (N_34672,N_31281,N_32253);
and U34673 (N_34673,N_31663,N_30708);
or U34674 (N_34674,N_32483,N_31621);
nand U34675 (N_34675,N_31562,N_30209);
nand U34676 (N_34676,N_32124,N_31916);
or U34677 (N_34677,N_31379,N_31143);
and U34678 (N_34678,N_30989,N_31694);
nor U34679 (N_34679,N_30204,N_31533);
nand U34680 (N_34680,N_30085,N_30567);
xor U34681 (N_34681,N_30844,N_30600);
and U34682 (N_34682,N_31325,N_31391);
nor U34683 (N_34683,N_32446,N_32294);
xor U34684 (N_34684,N_31671,N_31081);
xnor U34685 (N_34685,N_30974,N_32123);
xnor U34686 (N_34686,N_30768,N_31493);
or U34687 (N_34687,N_30131,N_31543);
nand U34688 (N_34688,N_31615,N_31796);
nand U34689 (N_34689,N_30772,N_31947);
and U34690 (N_34690,N_30428,N_30806);
nor U34691 (N_34691,N_32442,N_31979);
xor U34692 (N_34692,N_31241,N_32243);
xnor U34693 (N_34693,N_32029,N_30766);
and U34694 (N_34694,N_30550,N_30847);
nor U34695 (N_34695,N_31329,N_31881);
xnor U34696 (N_34696,N_31109,N_31907);
nor U34697 (N_34697,N_31724,N_31432);
nor U34698 (N_34698,N_30130,N_30341);
and U34699 (N_34699,N_30142,N_31122);
and U34700 (N_34700,N_32227,N_31135);
or U34701 (N_34701,N_31485,N_30982);
nor U34702 (N_34702,N_30907,N_31222);
or U34703 (N_34703,N_32314,N_30316);
and U34704 (N_34704,N_31288,N_30381);
xor U34705 (N_34705,N_31290,N_31888);
nor U34706 (N_34706,N_30332,N_30214);
and U34707 (N_34707,N_31633,N_30354);
xor U34708 (N_34708,N_30459,N_31835);
nand U34709 (N_34709,N_30133,N_30062);
nand U34710 (N_34710,N_31467,N_31848);
nand U34711 (N_34711,N_30824,N_32103);
nand U34712 (N_34712,N_30221,N_32191);
nor U34713 (N_34713,N_32447,N_32185);
nand U34714 (N_34714,N_32086,N_31161);
and U34715 (N_34715,N_32453,N_30262);
nand U34716 (N_34716,N_31245,N_30670);
and U34717 (N_34717,N_30284,N_32494);
and U34718 (N_34718,N_30917,N_32313);
and U34719 (N_34719,N_30192,N_32289);
nor U34720 (N_34720,N_31093,N_32450);
and U34721 (N_34721,N_30082,N_30801);
and U34722 (N_34722,N_31193,N_30015);
and U34723 (N_34723,N_32382,N_30098);
and U34724 (N_34724,N_32135,N_31186);
nor U34725 (N_34725,N_30732,N_32221);
and U34726 (N_34726,N_30050,N_30637);
xnor U34727 (N_34727,N_32157,N_30473);
xor U34728 (N_34728,N_30061,N_32380);
nand U34729 (N_34729,N_31875,N_30610);
or U34730 (N_34730,N_30941,N_30780);
or U34731 (N_34731,N_31058,N_31260);
or U34732 (N_34732,N_30798,N_30843);
and U34733 (N_34733,N_32306,N_32161);
nand U34734 (N_34734,N_30023,N_31386);
nor U34735 (N_34735,N_31187,N_31694);
or U34736 (N_34736,N_30967,N_30198);
nor U34737 (N_34737,N_31787,N_30460);
xnor U34738 (N_34738,N_31441,N_32055);
nand U34739 (N_34739,N_31952,N_30282);
and U34740 (N_34740,N_30000,N_31805);
or U34741 (N_34741,N_30250,N_31896);
or U34742 (N_34742,N_31998,N_32141);
or U34743 (N_34743,N_32311,N_31396);
or U34744 (N_34744,N_31660,N_31804);
nand U34745 (N_34745,N_30407,N_30229);
nand U34746 (N_34746,N_31636,N_30853);
and U34747 (N_34747,N_32359,N_30054);
nor U34748 (N_34748,N_32254,N_30301);
and U34749 (N_34749,N_31582,N_30176);
xnor U34750 (N_34750,N_31462,N_31124);
xor U34751 (N_34751,N_30359,N_31024);
nand U34752 (N_34752,N_30585,N_31386);
nor U34753 (N_34753,N_30359,N_31315);
nor U34754 (N_34754,N_32330,N_31360);
nand U34755 (N_34755,N_32014,N_30419);
and U34756 (N_34756,N_31339,N_31618);
nor U34757 (N_34757,N_30629,N_30512);
or U34758 (N_34758,N_31302,N_30961);
or U34759 (N_34759,N_31433,N_30556);
and U34760 (N_34760,N_30691,N_30047);
nor U34761 (N_34761,N_32177,N_31363);
or U34762 (N_34762,N_31512,N_30677);
and U34763 (N_34763,N_31497,N_31182);
nor U34764 (N_34764,N_31083,N_32294);
nand U34765 (N_34765,N_31052,N_32295);
nand U34766 (N_34766,N_32029,N_32148);
nand U34767 (N_34767,N_30530,N_31904);
and U34768 (N_34768,N_31836,N_30521);
nor U34769 (N_34769,N_32399,N_30610);
nand U34770 (N_34770,N_32082,N_31884);
or U34771 (N_34771,N_30066,N_31309);
xnor U34772 (N_34772,N_30598,N_30962);
nor U34773 (N_34773,N_31604,N_32201);
nand U34774 (N_34774,N_31241,N_31615);
nand U34775 (N_34775,N_31418,N_30153);
xor U34776 (N_34776,N_31086,N_32466);
and U34777 (N_34777,N_31193,N_30955);
or U34778 (N_34778,N_30400,N_31442);
nand U34779 (N_34779,N_31502,N_30665);
or U34780 (N_34780,N_31957,N_30442);
xnor U34781 (N_34781,N_30061,N_31511);
and U34782 (N_34782,N_30997,N_31061);
or U34783 (N_34783,N_31025,N_31338);
or U34784 (N_34784,N_31789,N_32261);
nor U34785 (N_34785,N_31045,N_31937);
nor U34786 (N_34786,N_30487,N_31674);
or U34787 (N_34787,N_30409,N_32018);
and U34788 (N_34788,N_31735,N_30312);
nand U34789 (N_34789,N_32458,N_31854);
nor U34790 (N_34790,N_30455,N_30149);
or U34791 (N_34791,N_32099,N_30867);
or U34792 (N_34792,N_30308,N_30257);
nor U34793 (N_34793,N_32210,N_31971);
nand U34794 (N_34794,N_30595,N_31902);
nand U34795 (N_34795,N_31065,N_32231);
or U34796 (N_34796,N_31178,N_30088);
and U34797 (N_34797,N_30125,N_31894);
and U34798 (N_34798,N_30511,N_32415);
nand U34799 (N_34799,N_30529,N_30612);
nor U34800 (N_34800,N_30150,N_30132);
nor U34801 (N_34801,N_30396,N_31918);
xor U34802 (N_34802,N_31039,N_30945);
nor U34803 (N_34803,N_30001,N_30705);
nand U34804 (N_34804,N_30048,N_32409);
and U34805 (N_34805,N_30650,N_31644);
or U34806 (N_34806,N_31490,N_31564);
xor U34807 (N_34807,N_31136,N_30233);
and U34808 (N_34808,N_30255,N_31483);
and U34809 (N_34809,N_30013,N_31859);
nand U34810 (N_34810,N_30034,N_31156);
xor U34811 (N_34811,N_30196,N_32152);
nand U34812 (N_34812,N_31991,N_31822);
nand U34813 (N_34813,N_31469,N_31048);
or U34814 (N_34814,N_30182,N_31951);
nor U34815 (N_34815,N_31859,N_31709);
xor U34816 (N_34816,N_32072,N_30127);
nand U34817 (N_34817,N_30627,N_30626);
nand U34818 (N_34818,N_30695,N_31735);
or U34819 (N_34819,N_30011,N_32144);
nor U34820 (N_34820,N_30094,N_30295);
nand U34821 (N_34821,N_31840,N_31149);
or U34822 (N_34822,N_30478,N_32323);
and U34823 (N_34823,N_31455,N_32011);
and U34824 (N_34824,N_31175,N_30783);
nand U34825 (N_34825,N_30842,N_32227);
nor U34826 (N_34826,N_31238,N_32058);
xor U34827 (N_34827,N_31025,N_30392);
and U34828 (N_34828,N_30038,N_31600);
xor U34829 (N_34829,N_30223,N_31407);
or U34830 (N_34830,N_31091,N_30955);
xor U34831 (N_34831,N_32290,N_32042);
or U34832 (N_34832,N_30219,N_30308);
nor U34833 (N_34833,N_31626,N_31094);
nor U34834 (N_34834,N_30440,N_30875);
nand U34835 (N_34835,N_31349,N_30020);
or U34836 (N_34836,N_31841,N_32148);
and U34837 (N_34837,N_30902,N_31878);
nand U34838 (N_34838,N_31628,N_30183);
or U34839 (N_34839,N_30126,N_31953);
xor U34840 (N_34840,N_30658,N_30933);
nand U34841 (N_34841,N_31549,N_32145);
or U34842 (N_34842,N_30538,N_31024);
nand U34843 (N_34843,N_30533,N_31112);
or U34844 (N_34844,N_30699,N_30366);
and U34845 (N_34845,N_31766,N_31540);
or U34846 (N_34846,N_30773,N_32351);
and U34847 (N_34847,N_30839,N_30798);
nor U34848 (N_34848,N_31361,N_30467);
nand U34849 (N_34849,N_30600,N_31622);
or U34850 (N_34850,N_30727,N_30774);
or U34851 (N_34851,N_30908,N_30244);
nand U34852 (N_34852,N_31796,N_30931);
nand U34853 (N_34853,N_31709,N_31564);
xnor U34854 (N_34854,N_31248,N_31836);
nand U34855 (N_34855,N_30094,N_30871);
nand U34856 (N_34856,N_31304,N_31223);
or U34857 (N_34857,N_31586,N_30203);
and U34858 (N_34858,N_31752,N_30090);
xor U34859 (N_34859,N_31232,N_31395);
nor U34860 (N_34860,N_31015,N_30983);
nor U34861 (N_34861,N_31686,N_31623);
nor U34862 (N_34862,N_32465,N_32068);
nand U34863 (N_34863,N_30842,N_31972);
nand U34864 (N_34864,N_30252,N_31711);
or U34865 (N_34865,N_31222,N_31944);
xnor U34866 (N_34866,N_31790,N_30964);
xnor U34867 (N_34867,N_30366,N_32150);
and U34868 (N_34868,N_30895,N_30053);
nand U34869 (N_34869,N_31529,N_32482);
or U34870 (N_34870,N_30651,N_31210);
or U34871 (N_34871,N_31823,N_31685);
and U34872 (N_34872,N_30445,N_31331);
nor U34873 (N_34873,N_31127,N_32499);
nor U34874 (N_34874,N_30116,N_30736);
nand U34875 (N_34875,N_30318,N_31089);
or U34876 (N_34876,N_31610,N_31675);
nor U34877 (N_34877,N_31140,N_30216);
nor U34878 (N_34878,N_32103,N_30775);
nor U34879 (N_34879,N_31076,N_31161);
and U34880 (N_34880,N_30154,N_30727);
xor U34881 (N_34881,N_32055,N_30697);
or U34882 (N_34882,N_31428,N_30439);
or U34883 (N_34883,N_30971,N_31534);
nor U34884 (N_34884,N_30239,N_30188);
and U34885 (N_34885,N_30576,N_30517);
or U34886 (N_34886,N_30711,N_31262);
or U34887 (N_34887,N_31541,N_32477);
nor U34888 (N_34888,N_32216,N_32149);
nor U34889 (N_34889,N_32090,N_31668);
or U34890 (N_34890,N_31289,N_30785);
or U34891 (N_34891,N_31426,N_32080);
and U34892 (N_34892,N_30290,N_30546);
nor U34893 (N_34893,N_32378,N_30408);
nor U34894 (N_34894,N_31663,N_30583);
xor U34895 (N_34895,N_30519,N_31453);
xnor U34896 (N_34896,N_31896,N_31095);
xnor U34897 (N_34897,N_31584,N_31744);
and U34898 (N_34898,N_30970,N_30292);
nand U34899 (N_34899,N_32381,N_31756);
and U34900 (N_34900,N_30768,N_30280);
nand U34901 (N_34901,N_30841,N_30356);
and U34902 (N_34902,N_30297,N_31145);
xnor U34903 (N_34903,N_30071,N_30303);
xor U34904 (N_34904,N_30667,N_31325);
nor U34905 (N_34905,N_32121,N_30188);
nor U34906 (N_34906,N_31029,N_30892);
xnor U34907 (N_34907,N_30427,N_32206);
or U34908 (N_34908,N_31417,N_32450);
nor U34909 (N_34909,N_31867,N_31648);
nand U34910 (N_34910,N_32239,N_30677);
or U34911 (N_34911,N_32293,N_32133);
and U34912 (N_34912,N_31434,N_30498);
nand U34913 (N_34913,N_30247,N_31394);
nor U34914 (N_34914,N_30508,N_31026);
or U34915 (N_34915,N_32028,N_31683);
nand U34916 (N_34916,N_31300,N_31210);
nand U34917 (N_34917,N_30901,N_31571);
nand U34918 (N_34918,N_31754,N_30585);
xor U34919 (N_34919,N_31134,N_31498);
nand U34920 (N_34920,N_31225,N_32425);
nand U34921 (N_34921,N_30411,N_30940);
nand U34922 (N_34922,N_30120,N_30097);
or U34923 (N_34923,N_32363,N_30607);
nor U34924 (N_34924,N_30080,N_30413);
xnor U34925 (N_34925,N_31173,N_31452);
nor U34926 (N_34926,N_30554,N_32270);
and U34927 (N_34927,N_32185,N_31875);
xor U34928 (N_34928,N_30966,N_32340);
nand U34929 (N_34929,N_30237,N_31585);
nand U34930 (N_34930,N_31596,N_30033);
xnor U34931 (N_34931,N_30005,N_32290);
xnor U34932 (N_34932,N_31383,N_30940);
and U34933 (N_34933,N_31958,N_32487);
xor U34934 (N_34934,N_31998,N_32356);
nor U34935 (N_34935,N_31100,N_30571);
xnor U34936 (N_34936,N_31321,N_31796);
nand U34937 (N_34937,N_30645,N_32451);
or U34938 (N_34938,N_30376,N_31080);
xor U34939 (N_34939,N_31692,N_32295);
or U34940 (N_34940,N_31397,N_31044);
xnor U34941 (N_34941,N_30493,N_30154);
nor U34942 (N_34942,N_31566,N_32300);
nor U34943 (N_34943,N_31264,N_30737);
and U34944 (N_34944,N_31756,N_31348);
or U34945 (N_34945,N_32352,N_32371);
and U34946 (N_34946,N_30566,N_31999);
nor U34947 (N_34947,N_32176,N_30839);
and U34948 (N_34948,N_32127,N_30447);
xnor U34949 (N_34949,N_30624,N_31316);
nor U34950 (N_34950,N_30499,N_30756);
nor U34951 (N_34951,N_32023,N_30836);
nor U34952 (N_34952,N_30625,N_30841);
nand U34953 (N_34953,N_30473,N_31407);
and U34954 (N_34954,N_30308,N_30787);
xnor U34955 (N_34955,N_31139,N_30938);
nor U34956 (N_34956,N_32292,N_32221);
xor U34957 (N_34957,N_30254,N_32463);
or U34958 (N_34958,N_31566,N_30822);
xnor U34959 (N_34959,N_30253,N_30799);
and U34960 (N_34960,N_30081,N_31864);
xor U34961 (N_34961,N_30380,N_31321);
xnor U34962 (N_34962,N_32345,N_31333);
nand U34963 (N_34963,N_31127,N_32404);
xor U34964 (N_34964,N_31581,N_32137);
and U34965 (N_34965,N_32387,N_30389);
or U34966 (N_34966,N_31686,N_31813);
nor U34967 (N_34967,N_31858,N_30713);
nand U34968 (N_34968,N_30542,N_32249);
nand U34969 (N_34969,N_31494,N_31923);
or U34970 (N_34970,N_30790,N_32273);
nor U34971 (N_34971,N_30800,N_32015);
and U34972 (N_34972,N_30385,N_30130);
nand U34973 (N_34973,N_30964,N_30592);
nor U34974 (N_34974,N_31441,N_30474);
and U34975 (N_34975,N_31505,N_31311);
xor U34976 (N_34976,N_32299,N_32290);
xor U34977 (N_34977,N_30467,N_32217);
xor U34978 (N_34978,N_30539,N_30464);
xor U34979 (N_34979,N_30974,N_31555);
nand U34980 (N_34980,N_30073,N_32233);
or U34981 (N_34981,N_30744,N_30026);
nor U34982 (N_34982,N_31848,N_30673);
and U34983 (N_34983,N_31854,N_32015);
nor U34984 (N_34984,N_31443,N_31912);
or U34985 (N_34985,N_31881,N_30574);
nand U34986 (N_34986,N_31246,N_30056);
xor U34987 (N_34987,N_32160,N_30274);
nor U34988 (N_34988,N_30579,N_30777);
nand U34989 (N_34989,N_32154,N_32091);
xnor U34990 (N_34990,N_31300,N_31280);
or U34991 (N_34991,N_30162,N_31900);
xor U34992 (N_34992,N_31840,N_30803);
xor U34993 (N_34993,N_31821,N_31175);
or U34994 (N_34994,N_32023,N_31981);
nor U34995 (N_34995,N_31294,N_30440);
nand U34996 (N_34996,N_30349,N_30363);
or U34997 (N_34997,N_31029,N_31737);
xnor U34998 (N_34998,N_30772,N_31560);
and U34999 (N_34999,N_31629,N_30797);
nand U35000 (N_35000,N_34321,N_33144);
or U35001 (N_35001,N_34871,N_33957);
xnor U35002 (N_35002,N_34434,N_32510);
nand U35003 (N_35003,N_33898,N_34925);
and U35004 (N_35004,N_34996,N_33348);
and U35005 (N_35005,N_34280,N_34405);
and U35006 (N_35006,N_34832,N_34042);
and U35007 (N_35007,N_34594,N_32578);
nor U35008 (N_35008,N_33347,N_34742);
nand U35009 (N_35009,N_33150,N_34847);
or U35010 (N_35010,N_34963,N_34284);
nand U35011 (N_35011,N_34156,N_33012);
xor U35012 (N_35012,N_34495,N_33039);
nor U35013 (N_35013,N_34320,N_33205);
and U35014 (N_35014,N_33421,N_34413);
nand U35015 (N_35015,N_33446,N_32822);
xor U35016 (N_35016,N_33302,N_33470);
xor U35017 (N_35017,N_34183,N_33016);
nand U35018 (N_35018,N_34962,N_34779);
xor U35019 (N_35019,N_33277,N_34363);
and U35020 (N_35020,N_32730,N_33418);
or U35021 (N_35021,N_34375,N_34549);
nand U35022 (N_35022,N_32585,N_34113);
or U35023 (N_35023,N_32896,N_34648);
nor U35024 (N_35024,N_34244,N_33378);
or U35025 (N_35025,N_34436,N_32518);
nor U35026 (N_35026,N_33059,N_33655);
nor U35027 (N_35027,N_34679,N_32731);
xor U35028 (N_35028,N_32936,N_33314);
nand U35029 (N_35029,N_33370,N_33000);
or U35030 (N_35030,N_34822,N_32916);
and U35031 (N_35031,N_32638,N_34262);
xor U35032 (N_35032,N_33162,N_33303);
nand U35033 (N_35033,N_32995,N_33800);
xnor U35034 (N_35034,N_32951,N_34678);
and U35035 (N_35035,N_32802,N_34386);
nor U35036 (N_35036,N_34353,N_33694);
xor U35037 (N_35037,N_34497,N_33249);
nand U35038 (N_35038,N_33168,N_33993);
and U35039 (N_35039,N_34719,N_33511);
xnor U35040 (N_35040,N_33915,N_34448);
xor U35041 (N_35041,N_32644,N_32891);
xor U35042 (N_35042,N_33074,N_33780);
nand U35043 (N_35043,N_34560,N_33923);
xnor U35044 (N_35044,N_32866,N_32875);
nor U35045 (N_35045,N_33936,N_34516);
nor U35046 (N_35046,N_34868,N_33280);
nor U35047 (N_35047,N_32751,N_34194);
and U35048 (N_35048,N_33757,N_34051);
and U35049 (N_35049,N_33424,N_33865);
xor U35050 (N_35050,N_34531,N_34544);
xor U35051 (N_35051,N_33621,N_33512);
xor U35052 (N_35052,N_34763,N_32674);
or U35053 (N_35053,N_34154,N_32668);
and U35054 (N_35054,N_34693,N_34027);
and U35055 (N_35055,N_33395,N_34293);
xor U35056 (N_35056,N_33637,N_32646);
and U35057 (N_35057,N_33760,N_33770);
nor U35058 (N_35058,N_33127,N_32877);
or U35059 (N_35059,N_34009,N_34241);
or U35060 (N_35060,N_34510,N_33774);
xor U35061 (N_35061,N_34869,N_33159);
xnor U35062 (N_35062,N_33591,N_33682);
nor U35063 (N_35063,N_33229,N_33002);
nand U35064 (N_35064,N_33636,N_34257);
xnor U35065 (N_35065,N_32840,N_34660);
xor U35066 (N_35066,N_34741,N_33350);
xor U35067 (N_35067,N_33769,N_33141);
and U35068 (N_35068,N_34374,N_34432);
nand U35069 (N_35069,N_32624,N_34961);
or U35070 (N_35070,N_33617,N_34049);
nor U35071 (N_35071,N_34715,N_34799);
and U35072 (N_35072,N_33742,N_33488);
and U35073 (N_35073,N_34317,N_34120);
nor U35074 (N_35074,N_34135,N_34443);
nand U35075 (N_35075,N_34389,N_34062);
and U35076 (N_35076,N_33029,N_33844);
nand U35077 (N_35077,N_33102,N_33836);
xnor U35078 (N_35078,N_34646,N_32832);
and U35079 (N_35079,N_33046,N_33525);
or U35080 (N_35080,N_32630,N_33459);
nor U35081 (N_35081,N_33261,N_32678);
xnor U35082 (N_35082,N_33325,N_33234);
and U35083 (N_35083,N_32736,N_32970);
and U35084 (N_35084,N_33807,N_33396);
or U35085 (N_35085,N_33641,N_34267);
nor U35086 (N_35086,N_33368,N_32548);
nand U35087 (N_35087,N_32604,N_32873);
or U35088 (N_35088,N_32829,N_33437);
or U35089 (N_35089,N_33548,N_32559);
nor U35090 (N_35090,N_34227,N_33092);
nand U35091 (N_35091,N_34199,N_34450);
xnor U35092 (N_35092,N_33916,N_33292);
and U35093 (N_35093,N_34654,N_34128);
nor U35094 (N_35094,N_32854,N_33251);
nor U35095 (N_35095,N_33560,N_34307);
or U35096 (N_35096,N_33266,N_33263);
nor U35097 (N_35097,N_33935,N_33026);
nor U35098 (N_35098,N_33887,N_32950);
or U35099 (N_35099,N_32892,N_34149);
or U35100 (N_35100,N_32582,N_34122);
nor U35101 (N_35101,N_34843,N_32557);
nor U35102 (N_35102,N_33824,N_34352);
xor U35103 (N_35103,N_33748,N_32561);
or U35104 (N_35104,N_33913,N_33164);
xnor U35105 (N_35105,N_33085,N_32969);
nor U35106 (N_35106,N_34444,N_32737);
nor U35107 (N_35107,N_33961,N_32922);
nand U35108 (N_35108,N_33593,N_33960);
xnor U35109 (N_35109,N_32629,N_34148);
and U35110 (N_35110,N_32977,N_32603);
and U35111 (N_35111,N_33466,N_34727);
or U35112 (N_35112,N_33108,N_33645);
xnor U35113 (N_35113,N_34647,N_33480);
and U35114 (N_35114,N_33499,N_34195);
nor U35115 (N_35115,N_34129,N_33040);
or U35116 (N_35116,N_34138,N_34515);
nor U35117 (N_35117,N_34109,N_33622);
nor U35118 (N_35118,N_32545,N_33216);
xor U35119 (N_35119,N_34520,N_33080);
xor U35120 (N_35120,N_33561,N_34941);
or U35121 (N_35121,N_33999,N_34038);
nand U35122 (N_35122,N_34087,N_33137);
xnor U35123 (N_35123,N_34312,N_33950);
or U35124 (N_35124,N_33296,N_34339);
or U35125 (N_35125,N_33390,N_33165);
and U35126 (N_35126,N_34596,N_34915);
nor U35127 (N_35127,N_34186,N_34787);
xor U35128 (N_35128,N_32820,N_34467);
nand U35129 (N_35129,N_32941,N_33351);
xnor U35130 (N_35130,N_33977,N_34229);
xor U35131 (N_35131,N_33096,N_32636);
or U35132 (N_35132,N_34395,N_33603);
xor U35133 (N_35133,N_33766,N_33830);
nor U35134 (N_35134,N_32806,N_34950);
and U35135 (N_35135,N_33762,N_32914);
xnor U35136 (N_35136,N_33065,N_33723);
or U35137 (N_35137,N_33627,N_34232);
nand U35138 (N_35138,N_33610,N_33199);
nor U35139 (N_35139,N_33495,N_33662);
nand U35140 (N_35140,N_34381,N_32800);
xnor U35141 (N_35141,N_33942,N_33740);
nand U35142 (N_35142,N_34850,N_32817);
nand U35143 (N_35143,N_34615,N_33030);
xor U35144 (N_35144,N_34644,N_33128);
nor U35145 (N_35145,N_34461,N_33187);
or U35146 (N_35146,N_34330,N_33650);
and U35147 (N_35147,N_32619,N_33364);
xnor U35148 (N_35148,N_34096,N_33404);
or U35149 (N_35149,N_32527,N_33743);
or U35150 (N_35150,N_33693,N_33870);
xor U35151 (N_35151,N_34757,N_32651);
and U35152 (N_35152,N_34433,N_33157);
nor U35153 (N_35153,N_33599,N_33772);
xor U35154 (N_35154,N_34652,N_33995);
or U35155 (N_35155,N_34631,N_34559);
and U35156 (N_35156,N_33947,N_34571);
and U35157 (N_35157,N_34823,N_32521);
xnor U35158 (N_35158,N_34401,N_34946);
or U35159 (N_35159,N_33872,N_34579);
nor U35160 (N_35160,N_33788,N_34604);
and U35161 (N_35161,N_32904,N_34700);
and U35162 (N_35162,N_33426,N_34171);
or U35163 (N_35163,N_33644,N_34970);
xnor U35164 (N_35164,N_34957,N_33809);
xnor U35165 (N_35165,N_32926,N_34091);
xnor U35166 (N_35166,N_33312,N_33103);
and U35167 (N_35167,N_34305,N_32750);
xnor U35168 (N_35168,N_34456,N_34713);
xnor U35169 (N_35169,N_33189,N_32958);
and U35170 (N_35170,N_32696,N_33555);
or U35171 (N_35171,N_34854,N_32520);
or U35172 (N_35172,N_33877,N_33531);
nor U35173 (N_35173,N_34285,N_34302);
and U35174 (N_35174,N_32972,N_34425);
nand U35175 (N_35175,N_33428,N_33808);
or U35176 (N_35176,N_33779,N_32990);
nor U35177 (N_35177,N_34662,N_34556);
and U35178 (N_35178,N_33532,N_32944);
nand U35179 (N_35179,N_34798,N_33005);
or U35180 (N_35180,N_33203,N_34292);
xor U35181 (N_35181,N_33543,N_33057);
nand U35182 (N_35182,N_34213,N_33295);
and U35183 (N_35183,N_33038,N_34726);
nor U35184 (N_35184,N_33520,N_32749);
or U35185 (N_35185,N_34979,N_33052);
nand U35186 (N_35186,N_33227,N_33569);
xnor U35187 (N_35187,N_32805,N_33115);
and U35188 (N_35188,N_34006,N_34377);
or U35189 (N_35189,N_32617,N_34675);
or U35190 (N_35190,N_33910,N_33828);
nand U35191 (N_35191,N_33601,N_33856);
nand U35192 (N_35192,N_33043,N_33900);
nand U35193 (N_35193,N_34037,N_33028);
nand U35194 (N_35194,N_34883,N_33465);
xor U35195 (N_35195,N_34772,N_34417);
or U35196 (N_35196,N_33385,N_33313);
nor U35197 (N_35197,N_32989,N_34641);
or U35198 (N_35198,N_33550,N_32581);
xnor U35199 (N_35199,N_34269,N_34424);
or U35200 (N_35200,N_32895,N_34756);
nor U35201 (N_35201,N_33089,N_33307);
xnor U35202 (N_35202,N_33876,N_32888);
xnor U35203 (N_35203,N_33691,N_34334);
and U35204 (N_35204,N_32858,N_33790);
nand U35205 (N_35205,N_34346,N_34001);
xor U35206 (N_35206,N_32708,N_33514);
nand U35207 (N_35207,N_33846,N_33792);
nor U35208 (N_35208,N_34501,N_32971);
and U35209 (N_35209,N_33642,N_34469);
and U35210 (N_35210,N_34905,N_33958);
or U35211 (N_35211,N_34233,N_32555);
nor U35212 (N_35212,N_34666,N_34512);
xnor U35213 (N_35213,N_32533,N_32500);
and U35214 (N_35214,N_33607,N_34688);
or U35215 (N_35215,N_34092,N_33411);
nand U35216 (N_35216,N_33355,N_33361);
or U35217 (N_35217,N_33729,N_32778);
or U35218 (N_35218,N_34259,N_33773);
nor U35219 (N_35219,N_33363,N_34766);
or U35220 (N_35220,N_33399,N_34609);
nand U35221 (N_35221,N_33899,N_34723);
xor U35222 (N_35222,N_34455,N_34539);
nor U35223 (N_35223,N_34316,N_33105);
and U35224 (N_35224,N_34837,N_32631);
xor U35225 (N_35225,N_34906,N_32899);
or U35226 (N_35226,N_34569,N_33291);
nor U35227 (N_35227,N_33112,N_32552);
nor U35228 (N_35228,N_32903,N_33657);
nand U35229 (N_35229,N_33463,N_34607);
nor U35230 (N_35230,N_34701,N_34031);
xor U35231 (N_35231,N_32852,N_34627);
nor U35232 (N_35232,N_34394,N_34537);
xor U35233 (N_35233,N_32835,N_34626);
nor U35234 (N_35234,N_33909,N_34115);
and U35235 (N_35235,N_33933,N_34892);
nand U35236 (N_35236,N_34484,N_33570);
nor U35237 (N_35237,N_33149,N_33275);
or U35238 (N_35238,N_33371,N_33563);
xnor U35239 (N_35239,N_34266,N_33737);
and U35240 (N_35240,N_34324,N_32655);
xor U35241 (N_35241,N_34606,N_33434);
or U35242 (N_35242,N_33994,N_33297);
nor U35243 (N_35243,N_34414,N_34355);
or U35244 (N_35244,N_33406,N_34474);
xor U35245 (N_35245,N_32998,N_32632);
and U35246 (N_35246,N_34791,N_34810);
xnor U35247 (N_35247,N_34802,N_34593);
xnor U35248 (N_35248,N_33687,N_34967);
and U35249 (N_35249,N_33822,N_32948);
nand U35250 (N_35250,N_33211,N_33242);
xnor U35251 (N_35251,N_33704,N_33450);
or U35252 (N_35252,N_34935,N_34612);
nor U35253 (N_35253,N_32550,N_33431);
nand U35254 (N_35254,N_33738,N_32723);
nand U35255 (N_35255,N_32567,N_33728);
nor U35256 (N_35256,N_33597,N_34958);
nor U35257 (N_35257,N_34332,N_33949);
and U35258 (N_35258,N_34438,N_32795);
and U35259 (N_35259,N_33606,N_32912);
nand U35260 (N_35260,N_34745,N_33353);
and U35261 (N_35261,N_34298,N_34240);
and U35262 (N_35262,N_33319,N_34888);
nand U35263 (N_35263,N_33321,N_34487);
or U35264 (N_35264,N_33640,N_33777);
nand U35265 (N_35265,N_34452,N_33509);
xnor U35266 (N_35266,N_33775,N_34390);
or U35267 (N_35267,N_32872,N_32687);
and U35268 (N_35268,N_33741,N_34525);
nor U35269 (N_35269,N_34093,N_33503);
nor U35270 (N_35270,N_34178,N_34538);
nor U35271 (N_35271,N_34211,N_34047);
or U35272 (N_35272,N_34327,N_34057);
and U35273 (N_35273,N_32964,N_34904);
nand U35274 (N_35274,N_34046,N_34420);
and U35275 (N_35275,N_32868,N_33415);
nor U35276 (N_35276,N_34845,N_34325);
or U35277 (N_35277,N_34916,N_33394);
and U35278 (N_35278,N_33282,N_32695);
or U35279 (N_35279,N_34658,N_33104);
nor U35280 (N_35280,N_34570,N_32766);
nor U35281 (N_35281,N_32671,N_33519);
or U35282 (N_35282,N_34349,N_32519);
and U35283 (N_35283,N_33471,N_34851);
or U35284 (N_35284,N_34121,N_33695);
nand U35285 (N_35285,N_34014,N_32662);
and U35286 (N_35286,N_33629,N_33072);
nor U35287 (N_35287,N_34749,N_34210);
or U35288 (N_35288,N_33624,N_33880);
and U35289 (N_35289,N_34770,N_34730);
nor U35290 (N_35290,N_32601,N_33546);
xor U35291 (N_35291,N_33985,N_33100);
and U35292 (N_35292,N_33575,N_34479);
or U35293 (N_35293,N_33930,N_34595);
and U35294 (N_35294,N_33449,N_34181);
nor U35295 (N_35295,N_34318,N_33182);
or U35296 (N_35296,N_34729,N_32931);
nand U35297 (N_35297,N_33990,N_33045);
nand U35298 (N_35298,N_34739,N_32901);
or U35299 (N_35299,N_34836,N_34295);
and U35300 (N_35300,N_33095,N_34776);
and U35301 (N_35301,N_34427,N_33230);
or U35302 (N_35302,N_33515,N_34496);
or U35303 (N_35303,N_33088,N_33716);
or U35304 (N_35304,N_34446,N_32774);
xnor U35305 (N_35305,N_34508,N_32517);
nand U35306 (N_35306,N_32924,N_33265);
and U35307 (N_35307,N_33849,N_33969);
nand U35308 (N_35308,N_34478,N_33857);
xnor U35309 (N_35309,N_34095,N_33153);
nor U35310 (N_35310,N_33120,N_32846);
and U35311 (N_35311,N_32568,N_34278);
nand U35312 (N_35312,N_33210,N_34864);
nor U35313 (N_35313,N_33562,N_33281);
nand U35314 (N_35314,N_32974,N_34614);
nor U35315 (N_35315,N_33568,N_33253);
or U35316 (N_35316,N_32883,N_32928);
or U35317 (N_35317,N_33823,N_34392);
nor U35318 (N_35318,N_33311,N_34174);
nor U35319 (N_35319,N_33663,N_33479);
and U35320 (N_35320,N_34918,N_33338);
nor U35321 (N_35321,N_32576,N_32610);
nor U35322 (N_35322,N_33988,N_33763);
and U35323 (N_35323,N_32734,N_34687);
xor U35324 (N_35324,N_33217,N_32560);
or U35325 (N_35325,N_33412,N_34072);
xnor U35326 (N_35326,N_33264,N_33342);
and U35327 (N_35327,N_34912,N_33707);
and U35328 (N_35328,N_33816,N_34402);
nand U35329 (N_35329,N_34069,N_34075);
nor U35330 (N_35330,N_33441,N_34873);
nand U35331 (N_35331,N_33722,N_33208);
and U35332 (N_35332,N_34786,N_34633);
and U35333 (N_35333,N_33061,N_33996);
xor U35334 (N_35334,N_32682,N_33286);
nand U35335 (N_35335,N_34026,N_34198);
and U35336 (N_35336,N_33559,N_33653);
and U35337 (N_35337,N_34754,N_32894);
nor U35338 (N_35338,N_34640,N_34220);
or U35339 (N_35339,N_34040,N_32839);
nand U35340 (N_35340,N_32616,N_33970);
or U35341 (N_35341,N_34807,N_33007);
or U35342 (N_35342,N_33982,N_33457);
or U35343 (N_35343,N_33445,N_32620);
xnor U35344 (N_35344,N_34564,N_34231);
nor U35345 (N_35345,N_34442,N_33078);
and U35346 (N_35346,N_34709,N_34929);
xor U35347 (N_35347,N_34483,N_34272);
nor U35348 (N_35348,N_33130,N_33639);
and U35349 (N_35349,N_33478,N_33146);
or U35350 (N_35350,N_32741,N_33528);
and U35351 (N_35351,N_34790,N_32673);
nand U35352 (N_35352,N_34418,N_34236);
xor U35353 (N_35353,N_34750,N_32934);
and U35354 (N_35354,N_34383,N_32718);
or U35355 (N_35355,N_32588,N_32540);
nand U35356 (N_35356,N_34590,N_34717);
xnor U35357 (N_35357,N_34264,N_32915);
nor U35358 (N_35358,N_33712,N_33320);
and U35359 (N_35359,N_33033,N_34322);
nor U35360 (N_35360,N_33798,N_32874);
nor U35361 (N_35361,N_33207,N_33925);
xor U35362 (N_35362,N_33420,N_33684);
or U35363 (N_35363,N_34553,N_34649);
nor U35364 (N_35364,N_33226,N_32975);
and U35365 (N_35365,N_34785,N_32511);
nor U35366 (N_35366,N_34792,N_32641);
and U35367 (N_35367,N_34488,N_33919);
nor U35368 (N_35368,N_33681,N_34521);
and U35369 (N_35369,N_33116,N_33576);
nor U35370 (N_35370,N_32979,N_33241);
nor U35371 (N_35371,N_33219,N_34634);
nand U35372 (N_35372,N_32523,N_34019);
and U35373 (N_35373,N_34254,N_34067);
and U35374 (N_35374,N_32698,N_33502);
nor U35375 (N_35375,N_34509,N_34992);
or U35376 (N_35376,N_32592,N_34677);
xnor U35377 (N_35377,N_33492,N_33670);
nand U35378 (N_35378,N_32591,N_33158);
or U35379 (N_35379,N_33700,N_34147);
xor U35380 (N_35380,N_32783,N_32684);
or U35381 (N_35381,N_32539,N_32833);
and U35382 (N_35382,N_33572,N_34856);
nor U35383 (N_35383,N_33076,N_33535);
nand U35384 (N_35384,N_34907,N_32670);
or U35385 (N_35385,N_34094,N_33764);
xnor U35386 (N_35386,N_34577,N_34133);
xnor U35387 (N_35387,N_34419,N_34350);
nand U35388 (N_35388,N_32532,N_33324);
xor U35389 (N_35389,N_34068,N_33091);
nor U35390 (N_35390,N_34185,N_34364);
nand U35391 (N_35391,N_34986,N_34228);
xnor U35392 (N_35392,N_33049,N_33031);
xnor U35393 (N_35393,N_33300,N_34050);
nand U35394 (N_35394,N_32823,N_34555);
and U35395 (N_35395,N_33018,N_33972);
xor U35396 (N_35396,N_34074,N_34025);
and U35397 (N_35397,N_33304,N_32770);
nand U35398 (N_35398,N_32508,N_33485);
or U35399 (N_35399,N_32953,N_33136);
xnor U35400 (N_35400,N_34784,N_33931);
and U35401 (N_35401,N_32801,N_34919);
and U35402 (N_35402,N_34956,N_33027);
nor U35403 (N_35403,N_34550,N_34933);
and U35404 (N_35404,N_33160,N_33486);
or U35405 (N_35405,N_33138,N_34993);
and U35406 (N_35406,N_33889,N_33204);
or U35407 (N_35407,N_33482,N_33813);
or U35408 (N_35408,N_34066,N_32515);
nand U35409 (N_35409,N_33021,N_34406);
or U35410 (N_35410,N_34608,N_33221);
and U35411 (N_35411,N_33125,N_34329);
or U35412 (N_35412,N_34526,N_33283);
nor U35413 (N_35413,N_34277,N_34697);
and U35414 (N_35414,N_34782,N_34765);
or U35415 (N_35415,N_33940,N_34029);
or U35416 (N_35416,N_34440,N_32705);
and U35417 (N_35417,N_33778,N_33435);
xnor U35418 (N_35418,N_33098,N_34315);
nor U35419 (N_35419,N_33333,N_33875);
and U35420 (N_35420,N_32621,N_33452);
nor U35421 (N_35421,N_33209,N_34880);
nor U35422 (N_35422,N_34561,N_34475);
xnor U35423 (N_35423,N_34968,N_32597);
xor U35424 (N_35424,N_33391,N_32573);
or U35425 (N_35425,N_34920,N_34218);
xnor U35426 (N_35426,N_34192,N_32626);
or U35427 (N_35427,N_32772,N_34161);
or U35428 (N_35428,N_34775,N_32756);
or U35429 (N_35429,N_34153,N_32850);
or U35430 (N_35430,N_33551,N_34529);
nand U35431 (N_35431,N_34557,N_33475);
nor U35432 (N_35432,N_34004,N_32654);
and U35433 (N_35433,N_34989,N_33692);
nand U35434 (N_35434,N_34473,N_33060);
nor U35435 (N_35435,N_34758,N_34441);
and U35436 (N_35436,N_33817,N_34482);
xor U35437 (N_35437,N_33014,N_33101);
nor U35438 (N_35438,N_33006,N_33821);
xor U35439 (N_35439,N_33683,N_34082);
xnor U35440 (N_35440,N_33832,N_32955);
and U35441 (N_35441,N_34347,N_33643);
and U35442 (N_35442,N_34106,N_33212);
or U35443 (N_35443,N_33058,N_34423);
nor U35444 (N_35444,N_33134,N_34548);
or U35445 (N_35445,N_34209,N_32694);
and U35446 (N_35446,N_34528,N_33791);
nand U35447 (N_35447,N_33400,N_34477);
nor U35448 (N_35448,N_34000,N_34415);
xnor U35449 (N_35449,N_34033,N_34337);
and U35450 (N_35450,N_34372,N_33267);
and U35451 (N_35451,N_34952,N_32572);
or U35452 (N_35452,N_32963,N_33938);
nor U35453 (N_35453,N_32930,N_33097);
or U35454 (N_35454,N_34629,N_34533);
and U35455 (N_35455,N_33920,N_33331);
and U35456 (N_35456,N_34672,N_34168);
nor U35457 (N_35457,N_34740,N_34387);
nor U35458 (N_35458,N_34541,N_32733);
and U35459 (N_35459,N_33504,N_32743);
and U35460 (N_35460,N_32994,N_34975);
nand U35461 (N_35461,N_33191,N_33318);
xor U35462 (N_35462,N_32815,N_33501);
nor U35463 (N_35463,N_33124,N_34724);
and U35464 (N_35464,N_33079,N_32965);
or U35465 (N_35465,N_33565,N_34796);
nand U35466 (N_35466,N_32952,N_34472);
and U35467 (N_35467,N_33863,N_33093);
nor U35468 (N_35468,N_33944,N_33652);
xnor U35469 (N_35469,N_33294,N_34485);
nor U35470 (N_35470,N_33632,N_33615);
nor U35471 (N_35471,N_34585,N_34499);
and U35472 (N_35472,N_34205,N_32623);
and U35473 (N_35473,N_34877,N_34767);
nor U35474 (N_35474,N_33335,N_32675);
or U35475 (N_35475,N_34458,N_33534);
xor U35476 (N_35476,N_33177,N_33143);
nand U35477 (N_35477,N_32633,N_34300);
nand U35478 (N_35478,N_34552,N_32849);
and U35479 (N_35479,N_33902,N_33270);
or U35480 (N_35480,N_34447,N_34587);
xor U35481 (N_35481,N_34197,N_33571);
nor U35482 (N_35482,N_32787,N_33491);
and U35483 (N_35483,N_34769,N_34494);
xnor U35484 (N_35484,N_33864,N_33186);
xor U35485 (N_35485,N_33032,N_34600);
nor U35486 (N_35486,N_33619,N_33951);
and U35487 (N_35487,N_32810,N_33952);
or U35488 (N_35488,N_34953,N_33689);
xor U35489 (N_35489,N_34777,N_34431);
and U35490 (N_35490,N_34463,N_33943);
or U35491 (N_35491,N_34221,N_32615);
and U35492 (N_35492,N_34797,N_33513);
and U35493 (N_35493,N_34833,N_34625);
nor U35494 (N_35494,N_34196,N_34621);
nand U35495 (N_35495,N_33834,N_33118);
and U35496 (N_35496,N_33440,N_33696);
nor U35497 (N_35497,N_33498,N_34809);
nand U35498 (N_35498,N_33070,N_32614);
and U35499 (N_35499,N_32506,N_34151);
nand U35500 (N_35500,N_34759,N_34780);
nand U35501 (N_35501,N_33768,N_34188);
or U35502 (N_35502,N_34959,N_34408);
xnor U35503 (N_35503,N_34720,N_33987);
and U35504 (N_35504,N_34393,N_34651);
xor U35505 (N_35505,N_34099,N_34131);
nand U35506 (N_35506,N_34744,N_34289);
or U35507 (N_35507,N_34960,N_34309);
nor U35508 (N_35508,N_34172,N_33948);
nand U35509 (N_35509,N_34492,N_33236);
xnor U35510 (N_35510,N_33148,N_32920);
nand U35511 (N_35511,N_33937,N_34603);
or U35512 (N_35512,N_33317,N_33739);
xor U35513 (N_35513,N_34323,N_33968);
and U35514 (N_35514,N_33050,N_34565);
xor U35515 (N_35515,N_34578,N_33754);
or U35516 (N_35516,N_33839,N_32602);
and U35517 (N_35517,N_34642,N_33705);
nand U35518 (N_35518,N_34985,N_33362);
nor U35519 (N_35519,N_34110,N_34704);
and U35520 (N_35520,N_33299,N_34870);
and U35521 (N_35521,N_34853,N_34200);
and U35522 (N_35522,N_33068,N_32507);
nor U35523 (N_35523,N_32870,N_33521);
nand U35524 (N_35524,N_33175,N_33954);
xnor U35525 (N_35525,N_33825,N_33003);
and U35526 (N_35526,N_34511,N_34878);
xor U35527 (N_35527,N_33557,N_32861);
nand U35528 (N_35528,N_34097,N_32625);
xor U35529 (N_35529,N_33978,N_34490);
or U35530 (N_35530,N_34846,N_33962);
and U35531 (N_35531,N_34338,N_32702);
and U35532 (N_35532,N_32685,N_33776);
nor U35533 (N_35533,N_34969,N_33380);
and U35534 (N_35534,N_33596,N_34400);
nor U35535 (N_35535,N_33556,N_33195);
xor U35536 (N_35536,N_32628,N_33429);
nand U35537 (N_35537,N_34303,N_33672);
nor U35538 (N_35538,N_34602,N_34020);
and U35539 (N_35539,N_34155,N_34685);
or U35540 (N_35540,N_34623,N_32857);
nand U35541 (N_35541,N_34982,N_32716);
nor U35542 (N_35542,N_32598,N_32844);
and U35543 (N_35543,N_32547,N_33537);
and U35544 (N_35544,N_34910,N_34706);
nand U35545 (N_35545,N_33751,N_34036);
and U35546 (N_35546,N_34812,N_33518);
or U35547 (N_35547,N_33886,N_33473);
nor U35548 (N_35548,N_34839,N_33132);
xnor U35549 (N_35549,N_34301,N_33609);
nor U35550 (N_35550,N_34283,N_33860);
and U35551 (N_35551,N_33912,N_34624);
and U35552 (N_35552,N_33494,N_32763);
xnor U35553 (N_35553,N_34369,N_33703);
and U35554 (N_35554,N_34103,N_32719);
nor U35555 (N_35555,N_34814,N_34690);
and U35556 (N_35556,N_33654,N_34725);
xor U35557 (N_35557,N_34650,N_34459);
or U35558 (N_35558,N_34551,N_33223);
or U35559 (N_35559,N_33022,N_32919);
nor U35560 (N_35560,N_33035,N_34680);
or U35561 (N_35561,N_34890,N_34670);
and U35562 (N_35562,N_34711,N_33794);
nor U35563 (N_35563,N_33544,N_34663);
or U35564 (N_35564,N_34145,N_34247);
nand U35565 (N_35565,N_32988,N_34628);
and U35566 (N_35566,N_33214,N_33287);
or U35567 (N_35567,N_33339,N_34365);
nor U35568 (N_35568,N_32725,N_32976);
or U35569 (N_35569,N_33679,N_33964);
nand U35570 (N_35570,N_33278,N_33169);
nor U35571 (N_35571,N_33747,N_32724);
xnor U35572 (N_35572,N_32594,N_32681);
nor U35573 (N_35573,N_33403,N_32530);
and U35574 (N_35574,N_32917,N_33170);
or U35575 (N_35575,N_33720,N_34336);
xnor U35576 (N_35576,N_33866,N_32762);
nor U35577 (N_35577,N_32525,N_32528);
nor U35578 (N_35578,N_32812,N_34589);
and U35579 (N_35579,N_33578,N_33932);
nand U35580 (N_35580,N_33468,N_34703);
nor U35581 (N_35581,N_34774,N_33852);
nand U35582 (N_35582,N_34238,N_33796);
xnor U35583 (N_35583,N_34189,N_33558);
nand U35584 (N_35584,N_32686,N_33590);
xor U35585 (N_35585,N_34102,N_32887);
nand U35586 (N_35586,N_34707,N_32600);
and U35587 (N_35587,N_32754,N_34219);
nand U35588 (N_35588,N_34924,N_34801);
or U35589 (N_35589,N_32947,N_34345);
or U35590 (N_35590,N_33811,N_33665);
or U35591 (N_35591,N_32786,N_33306);
nor U35592 (N_35592,N_34794,N_33927);
nand U35593 (N_35593,N_34536,N_33448);
or U35594 (N_35594,N_32885,N_34357);
nand U35595 (N_35595,N_32940,N_32622);
nor U35596 (N_35596,N_34157,N_32859);
and U35597 (N_35597,N_33117,N_33786);
nand U35598 (N_35598,N_33580,N_34524);
nand U35599 (N_35599,N_33476,N_34314);
and U35600 (N_35600,N_34972,N_34618);
nand U35601 (N_35601,N_34022,N_34088);
xor U35602 (N_35602,N_34588,N_33099);
xnor U35603 (N_35603,N_33755,N_33393);
or U35604 (N_35604,N_33896,N_32909);
and U35605 (N_35605,N_33174,N_32830);
nor U35606 (N_35606,N_32848,N_33009);
and U35607 (N_35607,N_34371,N_33373);
or U35608 (N_35608,N_32804,N_34849);
or U35609 (N_35609,N_33066,N_32522);
xor U35610 (N_35610,N_33257,N_32554);
nor U35611 (N_35611,N_34530,N_33829);
xnor U35612 (N_35612,N_32637,N_34655);
nand U35613 (N_35613,N_34965,N_34751);
or U35614 (N_35614,N_32590,N_34761);
or U35615 (N_35615,N_32529,N_34493);
nand U35616 (N_35616,N_33254,N_33733);
nand U35617 (N_35617,N_34054,N_34752);
or U35618 (N_35618,N_33472,N_34116);
nand U35619 (N_35619,N_34359,N_32808);
and U35620 (N_35620,N_33455,N_33245);
and U35621 (N_35621,N_33036,N_33481);
nor U35622 (N_35622,N_34255,N_33979);
xor U35623 (N_35623,N_33759,N_33011);
nor U35624 (N_35624,N_32889,N_32992);
nor U35625 (N_35625,N_34384,N_34464);
nand U35626 (N_35626,N_34954,N_33397);
and U35627 (N_35627,N_32732,N_32939);
nand U35628 (N_35628,N_33167,N_32929);
nand U35629 (N_35629,N_34695,N_34114);
xnor U35630 (N_35630,N_33992,N_33464);
nand U35631 (N_35631,N_33417,N_32753);
nor U35632 (N_35632,N_33422,N_34998);
and U35633 (N_35633,N_34044,N_32665);
or U35634 (N_35634,N_34665,N_32838);
nor U35635 (N_35635,N_33524,N_34344);
nand U35636 (N_35636,N_34504,N_33676);
or U35637 (N_35637,N_32982,N_34328);
xnor U35638 (N_35638,N_34333,N_33688);
and U35639 (N_35639,N_33365,N_33414);
nand U35640 (N_35640,N_34416,N_33053);
xnor U35641 (N_35641,N_32618,N_34335);
nor U35642 (N_35642,N_34983,N_34830);
xnor U35643 (N_35643,N_34505,N_32713);
nor U35644 (N_35644,N_34673,N_33714);
or U35645 (N_35645,N_33273,N_34928);
or U35646 (N_35646,N_34990,N_34908);
nor U35647 (N_35647,N_34778,N_33664);
nor U35648 (N_35648,N_34800,N_34824);
xor U35649 (N_35649,N_34018,N_34852);
nor U35650 (N_35650,N_32714,N_34828);
or U35651 (N_35651,N_34123,N_34251);
and U35652 (N_35652,N_33725,N_32788);
or U35653 (N_35653,N_34773,N_33698);
nand U35654 (N_35654,N_32634,N_33010);
and U35655 (N_35655,N_34158,N_33155);
or U35656 (N_35656,N_33781,N_33062);
nor U35657 (N_35657,N_34502,N_34712);
nand U35658 (N_35658,N_33549,N_33232);
xor U35659 (N_35659,N_33054,N_33635);
and U35660 (N_35660,N_32985,N_34584);
xor U35661 (N_35661,N_34243,N_33357);
or U35662 (N_35662,N_33129,N_33041);
and U35663 (N_35663,N_33239,N_33218);
nor U35664 (N_35664,N_33462,N_34806);
nand U35665 (N_35665,N_33734,N_33197);
xnor U35666 (N_35666,N_33496,N_33855);
nand U35667 (N_35667,N_34831,N_34126);
or U35668 (N_35668,N_33647,N_32755);
and U35669 (N_35669,N_34217,N_34944);
or U35670 (N_35670,N_33904,N_33908);
or U35671 (N_35671,N_34964,N_33814);
and U35672 (N_35672,N_32991,N_32562);
or U35673 (N_35673,N_33447,N_34005);
or U35674 (N_35674,N_32607,N_33196);
or U35675 (N_35675,N_33439,N_33787);
nand U35676 (N_35676,N_33255,N_34903);
and U35677 (N_35677,N_34947,N_34008);
xor U35678 (N_35678,N_33853,N_34003);
or U35679 (N_35679,N_32796,N_34653);
xnor U35680 (N_35680,N_32780,N_32834);
xor U35681 (N_35681,N_34112,N_33107);
or U35682 (N_35682,N_33176,N_33083);
or U35683 (N_35683,N_33522,N_32853);
or U35684 (N_35684,N_33793,N_34245);
nand U35685 (N_35685,N_32986,N_33222);
or U35686 (N_35686,N_33675,N_32807);
xnor U35687 (N_35687,N_33113,N_34523);
nor U35688 (N_35688,N_34249,N_33458);
xnor U35689 (N_35689,N_34012,N_34517);
nor U35690 (N_35690,N_34879,N_34104);
and U35691 (N_35691,N_33797,N_33585);
and U35692 (N_35692,N_33795,N_34370);
nand U35693 (N_35693,N_32967,N_32993);
or U35694 (N_35694,N_34343,N_34601);
xnor U35695 (N_35695,N_34265,N_33732);
or U35696 (N_35696,N_34304,N_32764);
nand U35697 (N_35697,N_32609,N_33469);
and U35698 (N_35698,N_33436,N_34710);
and U35699 (N_35699,N_33869,N_32649);
and U35700 (N_35700,N_33034,N_34421);
nand U35701 (N_35701,N_33553,N_33467);
xor U35702 (N_35702,N_33260,N_33454);
xnor U35703 (N_35703,N_33888,N_33804);
nor U35704 (N_35704,N_33721,N_34645);
xor U35705 (N_35705,N_32842,N_33063);
nand U35706 (N_35706,N_34900,N_33248);
nand U35707 (N_35707,N_33341,N_33516);
or U35708 (N_35708,N_33956,N_32589);
and U35709 (N_35709,N_34581,N_33044);
or U35710 (N_35710,N_34914,N_33765);
nand U35711 (N_35711,N_33114,N_33666);
nand U35712 (N_35712,N_32689,N_32549);
nor U35713 (N_35713,N_32776,N_32587);
nand U35714 (N_35714,N_34354,N_32566);
xor U35715 (N_35715,N_34881,N_34270);
nand U35716 (N_35716,N_33905,N_33837);
nor U35717 (N_35717,N_33628,N_34945);
nand U35718 (N_35718,N_32900,N_32758);
nand U35719 (N_35719,N_33966,N_32595);
or U35720 (N_35720,N_33685,N_33674);
xnor U35721 (N_35721,N_32797,N_33991);
nor U35722 (N_35722,N_34404,N_34554);
and U35723 (N_35723,N_33184,N_33945);
nor U35724 (N_35724,N_33586,N_34002);
and U35725 (N_35725,N_33037,N_32845);
xnor U35726 (N_35726,N_32680,N_33483);
nor U35727 (N_35727,N_34617,N_34605);
or U35728 (N_35728,N_34016,N_32785);
nor U35729 (N_35729,N_33785,N_33783);
or U35730 (N_35730,N_34184,N_32978);
or U35731 (N_35731,N_33749,N_33474);
nor U35732 (N_35732,N_34235,N_33181);
nor U35733 (N_35733,N_32570,N_33246);
nor U35734 (N_35734,N_34638,N_33975);
nor U35735 (N_35735,N_33015,N_33024);
nor U35736 (N_35736,N_32913,N_33432);
and U35737 (N_35737,N_33198,N_32656);
or U35738 (N_35738,N_33258,N_33604);
xnor U35739 (N_35739,N_34412,N_34207);
nor U35740 (N_35740,N_33630,N_34476);
nand U35741 (N_35741,N_32608,N_33081);
nor U35742 (N_35742,N_34190,N_34966);
or U35743 (N_35743,N_32862,N_34534);
nand U35744 (N_35744,N_33077,N_34064);
or U35745 (N_35745,N_33897,N_33349);
and U35746 (N_35746,N_34620,N_32890);
and U35747 (N_35747,N_32580,N_34518);
or U35748 (N_35748,N_33252,N_33372);
or U35749 (N_35749,N_32761,N_32918);
or U35750 (N_35750,N_32980,N_34817);
and U35751 (N_35751,N_33192,N_34737);
nor U35752 (N_35752,N_34061,N_32536);
and U35753 (N_35753,N_34882,N_33744);
nand U35754 (N_35754,N_34201,N_32884);
nor U35755 (N_35755,N_33298,N_33677);
nand U35756 (N_35756,N_33354,N_33119);
xor U35757 (N_35757,N_34694,N_33308);
nand U35758 (N_35758,N_34951,N_33656);
nand U35759 (N_35759,N_33374,N_33600);
or U35760 (N_35760,N_33847,N_34052);
nand U35761 (N_35761,N_34755,N_32667);
and U35762 (N_35762,N_34820,N_34698);
and U35763 (N_35763,N_33926,N_34111);
nand U35764 (N_35764,N_34017,N_33826);
nor U35765 (N_35765,N_33582,N_32864);
xnor U35766 (N_35766,N_34065,N_33309);
nand U35767 (N_35767,N_32663,N_34348);
nand U35768 (N_35768,N_33658,N_33710);
nor U35769 (N_35769,N_32999,N_33984);
xnor U35770 (N_35770,N_34098,N_32826);
nor U35771 (N_35771,N_32571,N_33526);
xor U35772 (N_35772,N_33868,N_34889);
and U35773 (N_35773,N_34733,N_33699);
xnor U35774 (N_35774,N_33840,N_32672);
nand U35775 (N_35775,N_34760,N_33235);
nor U35776 (N_35776,N_34942,N_32898);
nand U35777 (N_35777,N_34119,N_33151);
or U35778 (N_35778,N_32669,N_34684);
xor U35779 (N_35779,N_33017,N_34768);
nand U35780 (N_35780,N_34043,N_33974);
nor U35781 (N_35781,N_32933,N_33240);
and U35782 (N_35782,N_33955,N_32531);
nor U35783 (N_35783,N_33894,N_33638);
and U35784 (N_35784,N_33506,N_33419);
and U35785 (N_35785,N_34169,N_34180);
nor U35786 (N_35786,N_33750,N_34714);
nor U35787 (N_35787,N_34816,N_34162);
or U35788 (N_35788,N_34388,N_34150);
or U35789 (N_35789,N_33861,N_32878);
and U35790 (N_35790,N_34212,N_34842);
and U35791 (N_35791,N_34215,N_33121);
nand U35792 (N_35792,N_34470,N_34071);
nor U35793 (N_35793,N_34913,N_33989);
or U35794 (N_35794,N_33055,N_33623);
xor U35795 (N_35795,N_32911,N_34575);
or U35796 (N_35796,N_34865,N_33577);
and U35797 (N_35797,N_33375,N_34108);
xnor U35798 (N_35798,N_32775,N_33858);
nor U35799 (N_35799,N_34858,N_32541);
nor U35800 (N_35800,N_33071,N_34248);
xnor U35801 (N_35801,N_34911,N_34616);
or U35802 (N_35802,N_33959,N_34451);
or U35803 (N_35803,N_33726,N_32943);
nand U35804 (N_35804,N_34276,N_32803);
and U35805 (N_35805,N_32575,N_33611);
and U35806 (N_35806,N_32869,N_33346);
nand U35807 (N_35807,N_33384,N_33730);
nand U35808 (N_35808,N_33831,N_32757);
and U35809 (N_35809,N_34762,N_32791);
xnor U35810 (N_35810,N_32688,N_34358);
nand U35811 (N_35811,N_33369,N_33301);
or U35812 (N_35812,N_33323,N_34073);
and U35813 (N_35813,N_34909,N_34610);
nor U35814 (N_35814,N_34311,N_34866);
or U35815 (N_35815,N_32599,N_32752);
and U35816 (N_35816,N_33614,N_34367);
nand U35817 (N_35817,N_34635,N_34803);
and U35818 (N_35818,N_34743,N_33884);
nor U35819 (N_35819,N_34891,N_32740);
and U35820 (N_35820,N_32769,N_34166);
and U35821 (N_35821,N_33382,N_34974);
and U35822 (N_35822,N_33201,N_33381);
and U35823 (N_35823,N_34471,N_33388);
or U35824 (N_35824,N_33574,N_33727);
or U35825 (N_35825,N_34214,N_34558);
xnor U35826 (N_35826,N_32825,N_33051);
and U35827 (N_35827,N_32676,N_32648);
or U35828 (N_35828,N_34216,N_32968);
or U35829 (N_35829,N_34141,N_33651);
and U35830 (N_35830,N_33276,N_33326);
nand U35831 (N_35831,N_34808,N_32534);
nand U35832 (N_35832,N_33193,N_33094);
and U35833 (N_35833,N_34342,N_34274);
nor U35834 (N_35834,N_33678,N_34592);
and U35835 (N_35835,N_34056,N_34055);
xnor U35836 (N_35836,N_34795,N_32871);
and U35837 (N_35837,N_33140,N_32876);
nor U35838 (N_35838,N_34535,N_32658);
xor U35839 (N_35839,N_33202,N_34857);
xor U35840 (N_35840,N_34771,N_34860);
nand U35841 (N_35841,N_34160,N_33711);
nor U35842 (N_35842,N_33272,N_32767);
and U35843 (N_35843,N_33131,N_33903);
xnor U35844 (N_35844,N_34764,N_33859);
nor U35845 (N_35845,N_33179,N_34224);
or U35846 (N_35846,N_34310,N_33986);
or U35847 (N_35847,N_34191,N_34735);
nor U35848 (N_35848,N_32771,N_34885);
nor U35849 (N_35849,N_32728,N_33819);
xnor U35850 (N_35850,N_33456,N_33206);
and U35851 (N_35851,N_34063,N_33082);
nor U35852 (N_35852,N_33237,N_33224);
or U35853 (N_35853,N_33881,N_33172);
xnor U35854 (N_35854,N_33867,N_32809);
nor U35855 (N_35855,N_32824,N_33367);
xor U35856 (N_35856,N_33946,N_32818);
xnor U35857 (N_35857,N_33735,N_33343);
nor U35858 (N_35858,N_33998,N_34669);
and U35859 (N_35859,N_33433,N_34748);
nand U35860 (N_35860,N_33517,N_33965);
and U35861 (N_35861,N_34101,N_32860);
xor U35862 (N_35862,N_34938,N_33269);
or U35863 (N_35863,N_34164,N_33668);
or U35864 (N_35864,N_33803,N_34734);
or U35865 (N_35865,N_33171,N_32946);
nor U35866 (N_35866,N_32923,N_33883);
nor U35867 (N_35867,N_34844,N_33806);
and U35868 (N_35868,N_34746,N_33659);
nor U35869 (N_35869,N_34893,N_34622);
and U35870 (N_35870,N_33566,N_32666);
and U35871 (N_35871,N_33625,N_33510);
or U35872 (N_35872,N_34407,N_32593);
or U35873 (N_35873,N_34902,N_34855);
and U35874 (N_35874,N_33360,N_32569);
xnor U35875 (N_35875,N_33922,N_34513);
xnor U35876 (N_35876,N_34130,N_33284);
and U35877 (N_35877,N_32865,N_34481);
or U35878 (N_35878,N_34411,N_32841);
or U35879 (N_35879,N_34449,N_32938);
and U35880 (N_35880,N_32987,N_34286);
or U35881 (N_35881,N_34811,N_34611);
xor U35882 (N_35882,N_32789,N_33508);
xor U35883 (N_35883,N_34326,N_34939);
nor U35884 (N_35884,N_33753,N_32942);
and U35885 (N_35885,N_34060,N_33154);
nand U35886 (N_35886,N_34203,N_33327);
and U35887 (N_35887,N_33756,N_34202);
and U35888 (N_35888,N_33356,N_34331);
nand U35889 (N_35889,N_34991,N_32784);
nand U35890 (N_35890,N_34023,N_32935);
and U35891 (N_35891,N_34437,N_34204);
nor U35892 (N_35892,N_34643,N_33451);
xnor U35893 (N_35893,N_32773,N_34127);
or U35894 (N_35894,N_34486,N_33892);
and U35895 (N_35895,N_33019,N_32503);
and U35896 (N_35896,N_33493,N_33135);
or U35897 (N_35897,N_33086,N_34976);
and U35898 (N_35898,N_32908,N_33767);
xor U35899 (N_35899,N_33020,N_32650);
and U35900 (N_35900,N_33719,N_34894);
nand U35901 (N_35901,N_32790,N_32886);
nor U35902 (N_35902,N_32577,N_32537);
and U35903 (N_35903,N_34899,N_32579);
xor U35904 (N_35904,N_34039,N_33069);
nor U35905 (N_35905,N_33873,N_34445);
nand U35906 (N_35906,N_32516,N_34430);
or U35907 (N_35907,N_33122,N_33835);
nor U35908 (N_35908,N_33523,N_32690);
and U35909 (N_35909,N_34971,N_32906);
nor U35910 (N_35910,N_34995,N_34242);
or U35911 (N_35911,N_32504,N_33090);
or U35912 (N_35912,N_32747,N_32693);
xnor U35913 (N_35913,N_33305,N_33142);
nor U35914 (N_35914,N_34137,N_32556);
xor U35915 (N_35915,N_32701,N_34170);
nor U35916 (N_35916,N_34639,N_33939);
nand U35917 (N_35917,N_34793,N_32851);
nand U35918 (N_35918,N_34591,N_33438);
nand U35919 (N_35919,N_34230,N_33634);
nand U35920 (N_35920,N_34728,N_32726);
xnor U35921 (N_35921,N_34498,N_34380);
nor U35922 (N_35922,N_34410,N_34013);
and U35923 (N_35923,N_32831,N_34896);
nand U35924 (N_35924,N_34253,N_33161);
xor U35925 (N_35925,N_33425,N_34597);
nor U35926 (N_35926,N_34290,N_32640);
xor U35927 (N_35927,N_33680,N_33745);
xnor U35928 (N_35928,N_33409,N_34821);
xor U35929 (N_35929,N_33713,N_34948);
nand U35930 (N_35930,N_34977,N_34256);
nor U35931 (N_35931,N_34319,N_33587);
nor U35932 (N_35932,N_33190,N_34783);
or U35933 (N_35933,N_33893,N_33322);
xnor U35934 (N_35934,N_33854,N_33166);
nor U35935 (N_35935,N_34884,N_34453);
and U35936 (N_35936,N_32627,N_33731);
nand U35937 (N_35937,N_32660,N_34034);
and U35938 (N_35938,N_33156,N_33147);
xor U35939 (N_35939,N_33841,N_32927);
xnor U35940 (N_35940,N_32957,N_34261);
nor U35941 (N_35941,N_33928,N_34500);
or U35942 (N_35942,N_34268,N_34288);
xor U35943 (N_35943,N_32819,N_33746);
and U35944 (N_35944,N_32799,N_32921);
xor U35945 (N_35945,N_34084,N_33259);
and U35946 (N_35946,N_34083,N_33025);
and U35947 (N_35947,N_33133,N_33497);
nand U35948 (N_35948,N_34351,N_34275);
nor U35949 (N_35949,N_33359,N_34173);
and U35950 (N_35950,N_34362,N_33589);
nand U35951 (N_35951,N_34076,N_33183);
or U35952 (N_35952,N_34306,N_32664);
or U35953 (N_35953,N_32611,N_34582);
nand U35954 (N_35954,N_33256,N_34296);
and U35955 (N_35955,N_34514,N_34177);
nor U35956 (N_35956,N_32657,N_32792);
and U35957 (N_35957,N_33220,N_33724);
xor U35958 (N_35958,N_32546,N_32882);
nand U35959 (N_35959,N_33529,N_32813);
or U35960 (N_35960,N_32781,N_33818);
or U35961 (N_35961,N_33953,N_32722);
nand U35962 (N_35962,N_32905,N_32509);
nand U35963 (N_35963,N_33243,N_32973);
xnor U35964 (N_35964,N_33316,N_34994);
and U35965 (N_35965,N_34079,N_33633);
nand U35966 (N_35966,N_34987,N_34689);
nand U35967 (N_35967,N_34573,N_33917);
or U35968 (N_35968,N_32811,N_33225);
or U35969 (N_35969,N_32729,N_34397);
xnor U35970 (N_35970,N_32699,N_33279);
and U35971 (N_35971,N_33547,N_34932);
xor U35972 (N_35972,N_33430,N_34439);
nor U35973 (N_35973,N_32596,N_34468);
and U35974 (N_35974,N_34804,N_34045);
xor U35975 (N_35975,N_34917,N_34124);
xor U35976 (N_35976,N_34930,N_34105);
xnor U35977 (N_35977,N_34032,N_32960);
or U35978 (N_35978,N_33882,N_34699);
nand U35979 (N_35979,N_34222,N_32538);
nor U35980 (N_35980,N_33848,N_33487);
xnor U35981 (N_35981,N_33538,N_32893);
and U35982 (N_35982,N_33536,N_33626);
nand U35983 (N_35983,N_34294,N_32843);
and U35984 (N_35984,N_33595,N_32759);
nor U35985 (N_35985,N_34258,N_34692);
and U35986 (N_35986,N_33649,N_34732);
nand U35987 (N_35987,N_32794,N_33377);
and U35988 (N_35988,N_32856,N_33366);
nand U35989 (N_35989,N_32574,N_34632);
nand U35990 (N_35990,N_34815,N_33268);
nor U35991 (N_35991,N_33484,N_33843);
or U35992 (N_35992,N_33500,N_33851);
xnor U35993 (N_35993,N_34542,N_34613);
xor U35994 (N_35994,N_32712,N_34179);
xor U35995 (N_35995,N_34922,N_33976);
nor U35996 (N_35996,N_34566,N_33973);
and U35997 (N_35997,N_34273,N_34366);
or U35998 (N_35998,N_34409,N_34898);
and U35999 (N_35999,N_33612,N_32902);
xor U36000 (N_36000,N_32710,N_34619);
or U36001 (N_36001,N_32821,N_33981);
nor U36002 (N_36002,N_32715,N_33461);
xnor U36003 (N_36003,N_33250,N_34299);
nand U36004 (N_36004,N_34146,N_33701);
xor U36005 (N_36005,N_33084,N_32692);
nand U36006 (N_36006,N_32744,N_32793);
xor U36007 (N_36007,N_34165,N_32652);
nor U36008 (N_36008,N_33564,N_32816);
xor U36009 (N_36009,N_33315,N_33238);
and U36010 (N_36010,N_32945,N_34234);
nand U36011 (N_36011,N_34738,N_33332);
xor U36012 (N_36012,N_33389,N_32542);
or U36013 (N_36013,N_34193,N_33001);
or U36014 (N_36014,N_33427,N_33941);
or U36015 (N_36015,N_32661,N_34716);
nor U36016 (N_36016,N_34260,N_34382);
nor U36017 (N_36017,N_32855,N_34574);
nor U36018 (N_36018,N_33921,N_34279);
xnor U36019 (N_36019,N_33752,N_34545);
or U36020 (N_36020,N_33056,N_33194);
xor U36021 (N_36021,N_33618,N_34360);
and U36022 (N_36022,N_34667,N_33336);
xor U36023 (N_36023,N_32742,N_34926);
and U36024 (N_36024,N_33885,N_33812);
xnor U36025 (N_36025,N_34356,N_32879);
nand U36026 (N_36026,N_33328,N_34840);
xnor U36027 (N_36027,N_33906,N_32612);
nand U36028 (N_36028,N_34980,N_33608);
or U36029 (N_36029,N_34895,N_34572);
or U36030 (N_36030,N_34636,N_33231);
and U36031 (N_36031,N_34140,N_34107);
nand U36032 (N_36032,N_34090,N_34818);
nand U36033 (N_36033,N_34540,N_34167);
or U36034 (N_36034,N_33188,N_34696);
xor U36035 (N_36035,N_33274,N_34819);
or U36036 (N_36036,N_32565,N_33200);
xnor U36037 (N_36037,N_32962,N_34931);
and U36038 (N_36038,N_34206,N_33901);
and U36039 (N_36039,N_33702,N_33718);
or U36040 (N_36040,N_33289,N_33708);
nand U36041 (N_36041,N_33799,N_34175);
xnor U36042 (N_36042,N_33386,N_33352);
xor U36043 (N_36043,N_33442,N_32720);
xor U36044 (N_36044,N_33330,N_32524);
nor U36045 (N_36045,N_33573,N_32697);
or U36046 (N_36046,N_33579,N_33805);
or U36047 (N_36047,N_34263,N_33911);
nand U36048 (N_36048,N_34035,N_33443);
nand U36049 (N_36049,N_34788,N_33862);
nand U36050 (N_36050,N_33980,N_34664);
nor U36051 (N_36051,N_32782,N_33971);
nor U36052 (N_36052,N_32551,N_33379);
and U36053 (N_36053,N_33581,N_34599);
and U36054 (N_36054,N_34781,N_33244);
xnor U36055 (N_36055,N_34875,N_34630);
nor U36056 (N_36056,N_34187,N_34568);
nand U36057 (N_36057,N_34070,N_33290);
and U36058 (N_36058,N_34674,N_34250);
nor U36059 (N_36059,N_32691,N_34547);
and U36060 (N_36060,N_32925,N_33895);
and U36061 (N_36061,N_33401,N_34398);
or U36062 (N_36062,N_34118,N_34376);
or U36063 (N_36063,N_34656,N_34080);
xor U36064 (N_36064,N_34861,N_33271);
xor U36065 (N_36065,N_32505,N_33262);
and U36066 (N_36066,N_34308,N_32513);
nand U36067 (N_36067,N_34053,N_34399);
and U36068 (N_36068,N_33402,N_34867);
and U36069 (N_36069,N_33761,N_34827);
xnor U36070 (N_36070,N_32748,N_33890);
or U36071 (N_36071,N_33173,N_34159);
nand U36072 (N_36072,N_32959,N_33358);
nor U36073 (N_36073,N_33023,N_32739);
nand U36074 (N_36074,N_34058,N_34225);
or U36075 (N_36075,N_34208,N_34085);
or U36076 (N_36076,N_33845,N_33407);
and U36077 (N_36077,N_32526,N_34021);
or U36078 (N_36078,N_33444,N_34313);
nor U36079 (N_36079,N_34586,N_34462);
or U36080 (N_36080,N_34731,N_33810);
or U36081 (N_36081,N_33334,N_34246);
xnor U36082 (N_36082,N_32639,N_32981);
nor U36083 (N_36083,N_34011,N_33983);
and U36084 (N_36084,N_33879,N_34391);
nand U36085 (N_36085,N_33815,N_34691);
nor U36086 (N_36086,N_34598,N_34519);
xor U36087 (N_36087,N_34921,N_34668);
or U36088 (N_36088,N_34747,N_33598);
nand U36089 (N_36089,N_34422,N_33008);
and U36090 (N_36090,N_33075,N_33542);
nand U36091 (N_36091,N_34527,N_34223);
nand U36092 (N_36092,N_33736,N_32613);
nor U36093 (N_36093,N_34718,N_33827);
or U36094 (N_36094,N_34686,N_33228);
nand U36095 (N_36095,N_33838,N_32836);
nor U36096 (N_36096,N_32956,N_34379);
or U36097 (N_36097,N_33527,N_32727);
nor U36098 (N_36098,N_34886,N_33613);
xnor U36099 (N_36099,N_34955,N_34736);
and U36100 (N_36100,N_32867,N_33541);
nor U36101 (N_36101,N_32983,N_34134);
nand U36102 (N_36102,N_34863,N_33784);
xor U36103 (N_36103,N_32583,N_33416);
nor U36104 (N_36104,N_33967,N_34999);
nand U36105 (N_36105,N_34454,N_32765);
xor U36106 (N_36106,N_34943,N_34059);
and U36107 (N_36107,N_33871,N_33106);
xnor U36108 (N_36108,N_34671,N_33410);
nand U36109 (N_36109,N_34089,N_32647);
or U36110 (N_36110,N_33288,N_33671);
or U36111 (N_36111,N_32635,N_33540);
and U36112 (N_36112,N_33408,N_32558);
or U36113 (N_36113,N_34506,N_33109);
nand U36114 (N_36114,N_33918,N_32881);
and U36115 (N_36115,N_33067,N_33706);
nand U36116 (N_36116,N_34563,N_34271);
xor U36117 (N_36117,N_32643,N_34435);
xor U36118 (N_36118,N_33842,N_34859);
nor U36119 (N_36119,N_34041,N_34176);
or U36120 (N_36120,N_33690,N_32544);
xnor U36121 (N_36121,N_33802,N_33584);
nand U36122 (N_36122,N_33878,N_32683);
and U36123 (N_36123,N_34659,N_32837);
nand U36124 (N_36124,N_32700,N_32910);
nand U36125 (N_36125,N_34949,N_34829);
nand U36126 (N_36126,N_33907,N_34466);
nor U36127 (N_36127,N_34676,N_34583);
nand U36128 (N_36128,N_33145,N_33489);
and U36129 (N_36129,N_34874,N_32814);
nand U36130 (N_36130,N_33850,N_32584);
or U36131 (N_36131,N_34239,N_33398);
and U36132 (N_36132,N_34403,N_34872);
xor U36133 (N_36133,N_32703,N_34546);
nor U36134 (N_36134,N_33567,N_33247);
and U36135 (N_36135,N_34015,N_34152);
nand U36136 (N_36136,N_33583,N_33789);
xnor U36137 (N_36137,N_34522,N_33087);
or U36138 (N_36138,N_34708,N_32706);
nand U36139 (N_36139,N_32961,N_34981);
and U36140 (N_36140,N_32514,N_34661);
xor U36141 (N_36141,N_32535,N_33233);
and U36142 (N_36142,N_32709,N_34024);
xor U36143 (N_36143,N_32711,N_34144);
and U36144 (N_36144,N_33152,N_34182);
xor U36145 (N_36145,N_33505,N_32996);
xor U36146 (N_36146,N_34489,N_33048);
and U36147 (N_36147,N_34532,N_33477);
and U36148 (N_36148,N_34139,N_33064);
and U36149 (N_36149,N_34077,N_33533);
xor U36150 (N_36150,N_34132,N_34901);
xnor U36151 (N_36151,N_34753,N_34428);
xor U36152 (N_36152,N_32949,N_34562);
nand U36153 (N_36153,N_32966,N_32863);
nor U36154 (N_36154,N_34378,N_32563);
nand U36155 (N_36155,N_33833,N_32897);
nand U36156 (N_36156,N_34503,N_32707);
nand U36157 (N_36157,N_34341,N_32642);
or U36158 (N_36158,N_33453,N_32659);
xor U36159 (N_36159,N_32735,N_34721);
xnor U36160 (N_36160,N_34825,N_34287);
nand U36161 (N_36161,N_34385,N_34978);
xnor U36162 (N_36162,N_34834,N_33661);
or U36163 (N_36163,N_33660,N_34426);
nor U36164 (N_36164,N_34078,N_33545);
xor U36165 (N_36165,N_34086,N_32847);
nor U36166 (N_36166,N_33669,N_34480);
nor U36167 (N_36167,N_33139,N_34580);
nor U36168 (N_36168,N_34081,N_34048);
xnor U36169 (N_36169,N_33667,N_32606);
nand U36170 (N_36170,N_34340,N_34543);
or U36171 (N_36171,N_34163,N_32984);
nand U36172 (N_36172,N_33293,N_34136);
nand U36173 (N_36173,N_32745,N_33997);
and U36174 (N_36174,N_33215,N_33934);
xnor U36175 (N_36175,N_34460,N_34841);
or U36176 (N_36176,N_32827,N_33423);
nor U36177 (N_36177,N_34927,N_34997);
nand U36178 (N_36178,N_34940,N_34252);
nor U36179 (N_36179,N_33801,N_33413);
and U36180 (N_36180,N_32564,N_33620);
and U36181 (N_36181,N_33013,N_34361);
nand U36182 (N_36182,N_32721,N_34465);
nand U36183 (N_36183,N_34897,N_33929);
xnor U36184 (N_36184,N_33592,N_33178);
and U36185 (N_36185,N_32543,N_34100);
or U36186 (N_36186,N_32502,N_33686);
and U36187 (N_36187,N_32704,N_33047);
xor U36188 (N_36188,N_34835,N_34030);
and U36189 (N_36189,N_33673,N_33717);
and U36190 (N_36190,N_33631,N_32677);
and U36191 (N_36191,N_33073,N_34988);
nor U36192 (N_36192,N_34876,N_34862);
and U36193 (N_36193,N_34681,N_32937);
nor U36194 (N_36194,N_34117,N_32798);
xor U36195 (N_36195,N_33616,N_34396);
xor U36196 (N_36196,N_34683,N_34702);
and U36197 (N_36197,N_34887,N_32738);
and U36198 (N_36198,N_33460,N_34457);
nor U36199 (N_36199,N_33337,N_32997);
nor U36200 (N_36200,N_33914,N_32932);
nor U36201 (N_36201,N_33111,N_34848);
nor U36202 (N_36202,N_33552,N_32768);
nand U36203 (N_36203,N_32907,N_34722);
nor U36204 (N_36204,N_34142,N_33004);
and U36205 (N_36205,N_33891,N_33392);
or U36206 (N_36206,N_34705,N_34923);
or U36207 (N_36207,N_33405,N_34934);
or U36208 (N_36208,N_33387,N_34805);
nor U36209 (N_36209,N_33530,N_33507);
or U36210 (N_36210,N_34297,N_33126);
or U36211 (N_36211,N_34028,N_33042);
xor U36212 (N_36212,N_32605,N_33758);
xnor U36213 (N_36213,N_34507,N_34838);
nor U36214 (N_36214,N_34491,N_33345);
nand U36215 (N_36215,N_34973,N_33110);
nor U36216 (N_36216,N_33539,N_32717);
nand U36217 (N_36217,N_34657,N_32501);
and U36218 (N_36218,N_32777,N_32679);
nor U36219 (N_36219,N_33376,N_32954);
or U36220 (N_36220,N_33213,N_34429);
and U36221 (N_36221,N_34291,N_33709);
xnor U36222 (N_36222,N_33285,N_33329);
xnor U36223 (N_36223,N_32828,N_34813);
xnor U36224 (N_36224,N_34637,N_33648);
xor U36225 (N_36225,N_33874,N_33554);
nor U36226 (N_36226,N_34282,N_33340);
xor U36227 (N_36227,N_33588,N_32645);
nor U36228 (N_36228,N_34007,N_33310);
xnor U36229 (N_36229,N_33697,N_33646);
nand U36230 (N_36230,N_33715,N_32760);
xor U36231 (N_36231,N_33185,N_33820);
or U36232 (N_36232,N_34373,N_33163);
xor U36233 (N_36233,N_33344,N_32553);
nand U36234 (N_36234,N_32779,N_33602);
and U36235 (N_36235,N_33963,N_34010);
nand U36236 (N_36236,N_32586,N_33490);
nor U36237 (N_36237,N_33605,N_33924);
or U36238 (N_36238,N_32746,N_34281);
xnor U36239 (N_36239,N_34789,N_34682);
and U36240 (N_36240,N_34937,N_33123);
nor U36241 (N_36241,N_34226,N_33383);
and U36242 (N_36242,N_34125,N_34576);
or U36243 (N_36243,N_33782,N_34984);
or U36244 (N_36244,N_32512,N_33771);
xor U36245 (N_36245,N_34237,N_34936);
xnor U36246 (N_36246,N_34368,N_33594);
or U36247 (N_36247,N_33180,N_34143);
or U36248 (N_36248,N_34567,N_34826);
nor U36249 (N_36249,N_32880,N_32653);
and U36250 (N_36250,N_34539,N_34069);
and U36251 (N_36251,N_34470,N_34119);
xor U36252 (N_36252,N_33305,N_33674);
or U36253 (N_36253,N_34341,N_33888);
and U36254 (N_36254,N_34204,N_34946);
and U36255 (N_36255,N_34748,N_32817);
nor U36256 (N_36256,N_34572,N_33871);
nor U36257 (N_36257,N_34825,N_32632);
xnor U36258 (N_36258,N_34384,N_33457);
nand U36259 (N_36259,N_32723,N_32526);
nor U36260 (N_36260,N_34137,N_33912);
or U36261 (N_36261,N_32745,N_34489);
or U36262 (N_36262,N_32768,N_33867);
or U36263 (N_36263,N_34365,N_33950);
xnor U36264 (N_36264,N_34081,N_32646);
or U36265 (N_36265,N_33623,N_34374);
or U36266 (N_36266,N_34417,N_32536);
or U36267 (N_36267,N_33504,N_33784);
and U36268 (N_36268,N_32966,N_33533);
nor U36269 (N_36269,N_32800,N_34613);
and U36270 (N_36270,N_33701,N_32802);
nor U36271 (N_36271,N_33925,N_34702);
xor U36272 (N_36272,N_34145,N_34872);
and U36273 (N_36273,N_33096,N_33122);
and U36274 (N_36274,N_33462,N_34909);
nor U36275 (N_36275,N_34108,N_33054);
and U36276 (N_36276,N_34484,N_33546);
nor U36277 (N_36277,N_32689,N_32653);
or U36278 (N_36278,N_34444,N_34849);
or U36279 (N_36279,N_34833,N_32931);
nor U36280 (N_36280,N_32942,N_34481);
nor U36281 (N_36281,N_33729,N_32606);
nand U36282 (N_36282,N_33828,N_34144);
nor U36283 (N_36283,N_33728,N_34298);
nor U36284 (N_36284,N_33514,N_34930);
xor U36285 (N_36285,N_32833,N_33800);
or U36286 (N_36286,N_33336,N_33137);
or U36287 (N_36287,N_33852,N_33669);
nand U36288 (N_36288,N_34861,N_34669);
or U36289 (N_36289,N_34903,N_34135);
and U36290 (N_36290,N_33696,N_33072);
nor U36291 (N_36291,N_34162,N_34161);
nor U36292 (N_36292,N_33643,N_33383);
nor U36293 (N_36293,N_32760,N_33435);
xor U36294 (N_36294,N_33495,N_34972);
and U36295 (N_36295,N_34066,N_32975);
nand U36296 (N_36296,N_32591,N_32520);
or U36297 (N_36297,N_34142,N_34416);
xor U36298 (N_36298,N_34075,N_33581);
nor U36299 (N_36299,N_32745,N_34266);
nand U36300 (N_36300,N_33255,N_33992);
nand U36301 (N_36301,N_32785,N_33862);
xnor U36302 (N_36302,N_33980,N_33868);
or U36303 (N_36303,N_33812,N_34496);
xor U36304 (N_36304,N_33847,N_33189);
nand U36305 (N_36305,N_32854,N_33101);
nor U36306 (N_36306,N_33342,N_33440);
nand U36307 (N_36307,N_34110,N_32678);
and U36308 (N_36308,N_34946,N_32717);
xnor U36309 (N_36309,N_34642,N_32657);
and U36310 (N_36310,N_33330,N_32796);
xor U36311 (N_36311,N_34105,N_32504);
nor U36312 (N_36312,N_33242,N_34194);
xnor U36313 (N_36313,N_34563,N_34742);
xnor U36314 (N_36314,N_32561,N_34019);
or U36315 (N_36315,N_33993,N_33452);
nor U36316 (N_36316,N_34905,N_33691);
nor U36317 (N_36317,N_32911,N_34407);
and U36318 (N_36318,N_33041,N_33294);
nand U36319 (N_36319,N_33519,N_33684);
xor U36320 (N_36320,N_34389,N_34712);
nor U36321 (N_36321,N_34753,N_32597);
or U36322 (N_36322,N_34660,N_32748);
or U36323 (N_36323,N_34123,N_32950);
or U36324 (N_36324,N_32804,N_32559);
nor U36325 (N_36325,N_34927,N_34471);
or U36326 (N_36326,N_33679,N_34860);
nand U36327 (N_36327,N_33242,N_34789);
xnor U36328 (N_36328,N_34265,N_33713);
or U36329 (N_36329,N_34764,N_34114);
or U36330 (N_36330,N_34024,N_34731);
and U36331 (N_36331,N_34765,N_32734);
xor U36332 (N_36332,N_33499,N_34051);
xnor U36333 (N_36333,N_34864,N_33825);
nor U36334 (N_36334,N_34402,N_34738);
nor U36335 (N_36335,N_33494,N_34547);
nor U36336 (N_36336,N_34820,N_32563);
or U36337 (N_36337,N_34491,N_33121);
xor U36338 (N_36338,N_33086,N_33712);
nand U36339 (N_36339,N_34343,N_33700);
or U36340 (N_36340,N_34102,N_34819);
xnor U36341 (N_36341,N_32814,N_34410);
nand U36342 (N_36342,N_33669,N_34266);
nand U36343 (N_36343,N_34285,N_34339);
xor U36344 (N_36344,N_32631,N_34978);
nor U36345 (N_36345,N_33518,N_34661);
and U36346 (N_36346,N_34571,N_32618);
and U36347 (N_36347,N_34305,N_33043);
and U36348 (N_36348,N_34401,N_33014);
nand U36349 (N_36349,N_34270,N_33426);
nand U36350 (N_36350,N_34596,N_32705);
or U36351 (N_36351,N_34115,N_34022);
or U36352 (N_36352,N_34112,N_34909);
xnor U36353 (N_36353,N_34636,N_33594);
xnor U36354 (N_36354,N_34751,N_33211);
nand U36355 (N_36355,N_34299,N_34059);
nand U36356 (N_36356,N_33464,N_32937);
and U36357 (N_36357,N_34806,N_33579);
xnor U36358 (N_36358,N_32761,N_34428);
nand U36359 (N_36359,N_33621,N_33692);
and U36360 (N_36360,N_34253,N_32586);
nand U36361 (N_36361,N_34386,N_32503);
nor U36362 (N_36362,N_32654,N_33293);
nand U36363 (N_36363,N_34144,N_34471);
xnor U36364 (N_36364,N_33911,N_32608);
xor U36365 (N_36365,N_34826,N_33033);
nor U36366 (N_36366,N_33999,N_34706);
xor U36367 (N_36367,N_32593,N_34654);
nand U36368 (N_36368,N_34220,N_33699);
nor U36369 (N_36369,N_33213,N_32594);
xor U36370 (N_36370,N_34254,N_33890);
or U36371 (N_36371,N_33611,N_34890);
or U36372 (N_36372,N_33468,N_33572);
xor U36373 (N_36373,N_33006,N_34575);
nor U36374 (N_36374,N_32543,N_33218);
nor U36375 (N_36375,N_33848,N_34474);
or U36376 (N_36376,N_33041,N_34338);
nor U36377 (N_36377,N_33830,N_33418);
nor U36378 (N_36378,N_32585,N_33706);
xnor U36379 (N_36379,N_32627,N_34906);
xnor U36380 (N_36380,N_34167,N_33992);
nand U36381 (N_36381,N_34510,N_34369);
nand U36382 (N_36382,N_34176,N_33418);
nand U36383 (N_36383,N_33116,N_33121);
xor U36384 (N_36384,N_34385,N_33426);
xnor U36385 (N_36385,N_33606,N_34864);
and U36386 (N_36386,N_34422,N_34401);
xnor U36387 (N_36387,N_33767,N_34504);
and U36388 (N_36388,N_34212,N_32710);
nand U36389 (N_36389,N_34126,N_33274);
nor U36390 (N_36390,N_32993,N_33421);
and U36391 (N_36391,N_33644,N_33203);
nand U36392 (N_36392,N_32611,N_34252);
xnor U36393 (N_36393,N_32639,N_33565);
xnor U36394 (N_36394,N_32946,N_34316);
xor U36395 (N_36395,N_33723,N_33845);
nand U36396 (N_36396,N_33270,N_34081);
nor U36397 (N_36397,N_33230,N_33191);
and U36398 (N_36398,N_34373,N_33505);
nor U36399 (N_36399,N_34875,N_34122);
nand U36400 (N_36400,N_34024,N_34570);
or U36401 (N_36401,N_33029,N_34402);
nor U36402 (N_36402,N_33409,N_33312);
or U36403 (N_36403,N_34996,N_33983);
nand U36404 (N_36404,N_34096,N_32760);
nand U36405 (N_36405,N_33323,N_34196);
or U36406 (N_36406,N_34312,N_33936);
nor U36407 (N_36407,N_33991,N_32577);
or U36408 (N_36408,N_33408,N_34822);
and U36409 (N_36409,N_32641,N_33364);
or U36410 (N_36410,N_33294,N_32639);
nand U36411 (N_36411,N_34588,N_34011);
and U36412 (N_36412,N_34855,N_34444);
xor U36413 (N_36413,N_32925,N_33332);
xor U36414 (N_36414,N_33635,N_33516);
xor U36415 (N_36415,N_34320,N_33755);
or U36416 (N_36416,N_32972,N_34451);
and U36417 (N_36417,N_34619,N_34586);
xnor U36418 (N_36418,N_32754,N_34524);
or U36419 (N_36419,N_34349,N_33794);
xnor U36420 (N_36420,N_34857,N_33704);
or U36421 (N_36421,N_34705,N_33321);
xnor U36422 (N_36422,N_33590,N_34247);
or U36423 (N_36423,N_32916,N_33744);
nand U36424 (N_36424,N_32732,N_32651);
xor U36425 (N_36425,N_33454,N_34254);
xnor U36426 (N_36426,N_34625,N_33944);
nand U36427 (N_36427,N_33402,N_32512);
or U36428 (N_36428,N_32612,N_34160);
and U36429 (N_36429,N_33971,N_33633);
and U36430 (N_36430,N_34629,N_34049);
and U36431 (N_36431,N_33594,N_34730);
and U36432 (N_36432,N_34941,N_32629);
and U36433 (N_36433,N_33113,N_34135);
nor U36434 (N_36434,N_32858,N_33299);
nor U36435 (N_36435,N_34903,N_33764);
or U36436 (N_36436,N_32634,N_33759);
xnor U36437 (N_36437,N_33505,N_33643);
nand U36438 (N_36438,N_34302,N_34373);
nand U36439 (N_36439,N_33649,N_33592);
or U36440 (N_36440,N_34564,N_32797);
nand U36441 (N_36441,N_33624,N_34063);
xor U36442 (N_36442,N_32660,N_33451);
nand U36443 (N_36443,N_34553,N_32796);
or U36444 (N_36444,N_34404,N_34615);
nor U36445 (N_36445,N_34529,N_33663);
or U36446 (N_36446,N_33839,N_32608);
and U36447 (N_36447,N_33411,N_34178);
nand U36448 (N_36448,N_32793,N_33052);
nor U36449 (N_36449,N_34993,N_33667);
and U36450 (N_36450,N_32660,N_32559);
and U36451 (N_36451,N_33391,N_33922);
or U36452 (N_36452,N_34257,N_32733);
xnor U36453 (N_36453,N_34583,N_34644);
xnor U36454 (N_36454,N_33180,N_32769);
or U36455 (N_36455,N_34236,N_34686);
nand U36456 (N_36456,N_32948,N_34057);
nor U36457 (N_36457,N_34843,N_33268);
nand U36458 (N_36458,N_33986,N_34280);
nor U36459 (N_36459,N_32915,N_34558);
or U36460 (N_36460,N_33292,N_34549);
nor U36461 (N_36461,N_33433,N_33937);
nor U36462 (N_36462,N_34437,N_34378);
nand U36463 (N_36463,N_32941,N_33588);
nor U36464 (N_36464,N_33881,N_34314);
and U36465 (N_36465,N_34990,N_33876);
nand U36466 (N_36466,N_33659,N_32671);
or U36467 (N_36467,N_33189,N_32834);
xor U36468 (N_36468,N_34162,N_34406);
nor U36469 (N_36469,N_33018,N_33526);
nor U36470 (N_36470,N_34146,N_33922);
or U36471 (N_36471,N_33764,N_32674);
xnor U36472 (N_36472,N_32519,N_33016);
and U36473 (N_36473,N_32874,N_33688);
and U36474 (N_36474,N_32911,N_33010);
and U36475 (N_36475,N_33310,N_33218);
or U36476 (N_36476,N_34573,N_33294);
nand U36477 (N_36477,N_34231,N_32963);
nor U36478 (N_36478,N_33399,N_34457);
or U36479 (N_36479,N_34119,N_33308);
nor U36480 (N_36480,N_34332,N_33150);
xor U36481 (N_36481,N_33304,N_32976);
nand U36482 (N_36482,N_34679,N_32947);
and U36483 (N_36483,N_34983,N_34215);
nor U36484 (N_36484,N_34795,N_33087);
or U36485 (N_36485,N_33964,N_34908);
nand U36486 (N_36486,N_32676,N_34301);
nor U36487 (N_36487,N_33750,N_32855);
xnor U36488 (N_36488,N_34728,N_34564);
or U36489 (N_36489,N_33204,N_33741);
or U36490 (N_36490,N_34018,N_33875);
nor U36491 (N_36491,N_33325,N_34659);
xnor U36492 (N_36492,N_33291,N_34224);
nand U36493 (N_36493,N_34922,N_33598);
xor U36494 (N_36494,N_33989,N_33657);
or U36495 (N_36495,N_33485,N_33767);
xor U36496 (N_36496,N_33295,N_34519);
and U36497 (N_36497,N_34076,N_32603);
nand U36498 (N_36498,N_34230,N_32757);
and U36499 (N_36499,N_32647,N_34325);
and U36500 (N_36500,N_33330,N_33470);
nor U36501 (N_36501,N_33120,N_33357);
and U36502 (N_36502,N_32562,N_32833);
xor U36503 (N_36503,N_33156,N_33235);
or U36504 (N_36504,N_34462,N_33085);
nor U36505 (N_36505,N_33664,N_33631);
and U36506 (N_36506,N_33861,N_32905);
or U36507 (N_36507,N_34039,N_34860);
nand U36508 (N_36508,N_33314,N_33091);
xor U36509 (N_36509,N_33680,N_33883);
or U36510 (N_36510,N_33846,N_34274);
nor U36511 (N_36511,N_34500,N_34172);
or U36512 (N_36512,N_33135,N_32729);
nand U36513 (N_36513,N_33948,N_33568);
and U36514 (N_36514,N_34557,N_34569);
or U36515 (N_36515,N_34363,N_34517);
and U36516 (N_36516,N_32827,N_33916);
or U36517 (N_36517,N_33615,N_33260);
xnor U36518 (N_36518,N_33885,N_33291);
xnor U36519 (N_36519,N_34774,N_32789);
and U36520 (N_36520,N_33528,N_34122);
nor U36521 (N_36521,N_32650,N_34751);
or U36522 (N_36522,N_33292,N_33332);
or U36523 (N_36523,N_33030,N_33844);
or U36524 (N_36524,N_33052,N_34836);
nor U36525 (N_36525,N_33621,N_32928);
nor U36526 (N_36526,N_33368,N_34765);
xnor U36527 (N_36527,N_34273,N_32538);
nor U36528 (N_36528,N_33488,N_34862);
and U36529 (N_36529,N_33674,N_33215);
nor U36530 (N_36530,N_34010,N_33488);
nor U36531 (N_36531,N_34345,N_33595);
nor U36532 (N_36532,N_33263,N_34476);
and U36533 (N_36533,N_33506,N_33230);
and U36534 (N_36534,N_34537,N_34901);
nor U36535 (N_36535,N_34908,N_33776);
nor U36536 (N_36536,N_33182,N_33023);
xnor U36537 (N_36537,N_34802,N_33696);
and U36538 (N_36538,N_32965,N_34377);
or U36539 (N_36539,N_34865,N_33261);
and U36540 (N_36540,N_32928,N_34785);
nor U36541 (N_36541,N_34579,N_34521);
xor U36542 (N_36542,N_34076,N_33670);
and U36543 (N_36543,N_33133,N_32760);
nor U36544 (N_36544,N_34993,N_33454);
xor U36545 (N_36545,N_32838,N_34463);
or U36546 (N_36546,N_34969,N_33445);
and U36547 (N_36547,N_32889,N_33779);
xor U36548 (N_36548,N_33496,N_32886);
nand U36549 (N_36549,N_33804,N_34963);
nor U36550 (N_36550,N_33888,N_34499);
or U36551 (N_36551,N_33465,N_32506);
and U36552 (N_36552,N_33217,N_32542);
nor U36553 (N_36553,N_34609,N_34757);
xnor U36554 (N_36554,N_32709,N_34214);
xor U36555 (N_36555,N_33296,N_34772);
or U36556 (N_36556,N_34622,N_34051);
and U36557 (N_36557,N_33969,N_33051);
nand U36558 (N_36558,N_32520,N_34733);
nand U36559 (N_36559,N_33411,N_32574);
nor U36560 (N_36560,N_33921,N_33378);
and U36561 (N_36561,N_34532,N_34880);
xnor U36562 (N_36562,N_33785,N_33777);
xor U36563 (N_36563,N_34131,N_34434);
nor U36564 (N_36564,N_34519,N_32936);
and U36565 (N_36565,N_32993,N_34246);
nand U36566 (N_36566,N_33758,N_34363);
and U36567 (N_36567,N_32729,N_33639);
or U36568 (N_36568,N_33581,N_34803);
and U36569 (N_36569,N_34525,N_34509);
xnor U36570 (N_36570,N_32553,N_33257);
xor U36571 (N_36571,N_34534,N_34900);
or U36572 (N_36572,N_34177,N_34148);
xor U36573 (N_36573,N_33066,N_34882);
or U36574 (N_36574,N_32532,N_33528);
xnor U36575 (N_36575,N_34924,N_34524);
nor U36576 (N_36576,N_34031,N_34886);
and U36577 (N_36577,N_33708,N_33975);
nand U36578 (N_36578,N_34884,N_34945);
xor U36579 (N_36579,N_34781,N_33201);
nor U36580 (N_36580,N_34952,N_34909);
xor U36581 (N_36581,N_33437,N_34988);
nor U36582 (N_36582,N_32524,N_32674);
nand U36583 (N_36583,N_33915,N_34282);
nand U36584 (N_36584,N_34962,N_33701);
or U36585 (N_36585,N_34257,N_33512);
nand U36586 (N_36586,N_34759,N_33622);
and U36587 (N_36587,N_33007,N_33586);
xor U36588 (N_36588,N_34056,N_33905);
nand U36589 (N_36589,N_33706,N_32625);
or U36590 (N_36590,N_32543,N_34520);
and U36591 (N_36591,N_34760,N_34646);
xnor U36592 (N_36592,N_33457,N_33649);
or U36593 (N_36593,N_33605,N_33055);
nor U36594 (N_36594,N_33857,N_32753);
xor U36595 (N_36595,N_34009,N_34457);
and U36596 (N_36596,N_34219,N_34056);
and U36597 (N_36597,N_33173,N_33044);
xor U36598 (N_36598,N_32850,N_34500);
or U36599 (N_36599,N_34488,N_32510);
or U36600 (N_36600,N_33333,N_34927);
nand U36601 (N_36601,N_33262,N_33478);
nand U36602 (N_36602,N_34914,N_33712);
xor U36603 (N_36603,N_34139,N_34067);
nor U36604 (N_36604,N_34994,N_32724);
xnor U36605 (N_36605,N_34966,N_34830);
xor U36606 (N_36606,N_33427,N_33292);
or U36607 (N_36607,N_34950,N_32641);
and U36608 (N_36608,N_34339,N_34254);
nand U36609 (N_36609,N_32631,N_33732);
nor U36610 (N_36610,N_34561,N_34290);
or U36611 (N_36611,N_34053,N_33316);
nand U36612 (N_36612,N_32840,N_33822);
and U36613 (N_36613,N_33390,N_32740);
or U36614 (N_36614,N_32972,N_34686);
nor U36615 (N_36615,N_33796,N_33683);
xnor U36616 (N_36616,N_33786,N_33765);
nor U36617 (N_36617,N_34314,N_33448);
nor U36618 (N_36618,N_33946,N_32920);
xnor U36619 (N_36619,N_32987,N_33729);
nand U36620 (N_36620,N_33616,N_33423);
and U36621 (N_36621,N_32619,N_34911);
nor U36622 (N_36622,N_32852,N_32928);
or U36623 (N_36623,N_33103,N_33301);
xnor U36624 (N_36624,N_33079,N_34518);
nor U36625 (N_36625,N_34483,N_34213);
nand U36626 (N_36626,N_34783,N_33522);
or U36627 (N_36627,N_34475,N_33627);
nor U36628 (N_36628,N_33874,N_33325);
xnor U36629 (N_36629,N_32665,N_34995);
nor U36630 (N_36630,N_34034,N_32521);
nand U36631 (N_36631,N_33158,N_34051);
or U36632 (N_36632,N_34496,N_32516);
nor U36633 (N_36633,N_32595,N_33725);
nor U36634 (N_36634,N_32796,N_32960);
nand U36635 (N_36635,N_34245,N_33669);
and U36636 (N_36636,N_32701,N_33095);
nor U36637 (N_36637,N_34215,N_34432);
and U36638 (N_36638,N_34718,N_33281);
or U36639 (N_36639,N_34455,N_34661);
nand U36640 (N_36640,N_32824,N_34785);
xnor U36641 (N_36641,N_33083,N_33325);
nand U36642 (N_36642,N_32524,N_32665);
and U36643 (N_36643,N_33357,N_33894);
nor U36644 (N_36644,N_32537,N_34531);
or U36645 (N_36645,N_33434,N_33803);
xor U36646 (N_36646,N_34501,N_33140);
nor U36647 (N_36647,N_33654,N_33779);
nand U36648 (N_36648,N_33317,N_33072);
and U36649 (N_36649,N_33038,N_32770);
nand U36650 (N_36650,N_34817,N_32535);
and U36651 (N_36651,N_33203,N_34711);
nand U36652 (N_36652,N_33494,N_34321);
and U36653 (N_36653,N_33543,N_34789);
nor U36654 (N_36654,N_33440,N_33534);
xor U36655 (N_36655,N_33560,N_32737);
nand U36656 (N_36656,N_34073,N_33526);
nor U36657 (N_36657,N_34949,N_32560);
nand U36658 (N_36658,N_34653,N_34659);
xor U36659 (N_36659,N_34377,N_34235);
or U36660 (N_36660,N_32527,N_33235);
or U36661 (N_36661,N_34189,N_34216);
xnor U36662 (N_36662,N_34775,N_33982);
nor U36663 (N_36663,N_34747,N_34859);
and U36664 (N_36664,N_33007,N_34669);
nand U36665 (N_36665,N_32520,N_33422);
xnor U36666 (N_36666,N_34528,N_34243);
or U36667 (N_36667,N_32849,N_32956);
and U36668 (N_36668,N_33612,N_33480);
nor U36669 (N_36669,N_33616,N_32719);
nor U36670 (N_36670,N_34951,N_34289);
nand U36671 (N_36671,N_32685,N_34824);
nand U36672 (N_36672,N_32644,N_32890);
and U36673 (N_36673,N_34588,N_32737);
nor U36674 (N_36674,N_33130,N_34748);
or U36675 (N_36675,N_34634,N_34424);
nor U36676 (N_36676,N_34481,N_34997);
and U36677 (N_36677,N_33215,N_32944);
xor U36678 (N_36678,N_34782,N_34657);
xnor U36679 (N_36679,N_34464,N_33845);
and U36680 (N_36680,N_33847,N_34191);
or U36681 (N_36681,N_33801,N_34608);
xor U36682 (N_36682,N_33542,N_34046);
or U36683 (N_36683,N_32728,N_34267);
nand U36684 (N_36684,N_33127,N_32793);
or U36685 (N_36685,N_32770,N_33958);
and U36686 (N_36686,N_33909,N_34910);
nand U36687 (N_36687,N_34956,N_34478);
nor U36688 (N_36688,N_34545,N_33003);
and U36689 (N_36689,N_34205,N_34432);
and U36690 (N_36690,N_33938,N_33502);
xor U36691 (N_36691,N_33332,N_32530);
or U36692 (N_36692,N_34811,N_33236);
and U36693 (N_36693,N_34042,N_32664);
nand U36694 (N_36694,N_33538,N_32674);
nor U36695 (N_36695,N_34026,N_34376);
or U36696 (N_36696,N_34051,N_32659);
and U36697 (N_36697,N_33983,N_34999);
nor U36698 (N_36698,N_32746,N_33665);
and U36699 (N_36699,N_33951,N_34309);
nor U36700 (N_36700,N_34438,N_32505);
or U36701 (N_36701,N_33477,N_34191);
nand U36702 (N_36702,N_33648,N_34869);
or U36703 (N_36703,N_33422,N_34222);
and U36704 (N_36704,N_32914,N_33284);
and U36705 (N_36705,N_33865,N_32722);
nand U36706 (N_36706,N_33806,N_34446);
and U36707 (N_36707,N_32691,N_33036);
and U36708 (N_36708,N_33551,N_33871);
xnor U36709 (N_36709,N_33284,N_33016);
nor U36710 (N_36710,N_33010,N_33497);
xor U36711 (N_36711,N_33134,N_33992);
nor U36712 (N_36712,N_33022,N_34372);
and U36713 (N_36713,N_34555,N_32838);
nand U36714 (N_36714,N_34723,N_33651);
xor U36715 (N_36715,N_33199,N_32729);
or U36716 (N_36716,N_32500,N_34045);
xnor U36717 (N_36717,N_33699,N_34361);
nand U36718 (N_36718,N_33229,N_34328);
nor U36719 (N_36719,N_33085,N_34492);
nor U36720 (N_36720,N_34538,N_33945);
nand U36721 (N_36721,N_34431,N_32630);
nor U36722 (N_36722,N_34777,N_34121);
or U36723 (N_36723,N_32982,N_32604);
and U36724 (N_36724,N_34915,N_34259);
or U36725 (N_36725,N_32686,N_33346);
nand U36726 (N_36726,N_32652,N_33285);
xor U36727 (N_36727,N_34849,N_33567);
nor U36728 (N_36728,N_34229,N_34613);
xor U36729 (N_36729,N_33857,N_33287);
and U36730 (N_36730,N_33305,N_32583);
xnor U36731 (N_36731,N_33406,N_34238);
xnor U36732 (N_36732,N_33224,N_34485);
and U36733 (N_36733,N_34041,N_33956);
and U36734 (N_36734,N_32633,N_34044);
nor U36735 (N_36735,N_33963,N_33700);
or U36736 (N_36736,N_32984,N_32956);
nor U36737 (N_36737,N_34200,N_33555);
nor U36738 (N_36738,N_34111,N_33783);
or U36739 (N_36739,N_33032,N_33997);
or U36740 (N_36740,N_32565,N_33946);
nor U36741 (N_36741,N_32894,N_34324);
xor U36742 (N_36742,N_32906,N_32803);
nand U36743 (N_36743,N_34718,N_32813);
xnor U36744 (N_36744,N_33618,N_34304);
nor U36745 (N_36745,N_34012,N_32539);
or U36746 (N_36746,N_32556,N_32680);
and U36747 (N_36747,N_33978,N_33465);
nor U36748 (N_36748,N_33227,N_32984);
nand U36749 (N_36749,N_33437,N_34582);
nor U36750 (N_36750,N_34688,N_33113);
or U36751 (N_36751,N_34007,N_33421);
nor U36752 (N_36752,N_33598,N_34458);
and U36753 (N_36753,N_34403,N_34580);
nor U36754 (N_36754,N_34814,N_33834);
nand U36755 (N_36755,N_33940,N_34204);
nand U36756 (N_36756,N_33465,N_34430);
or U36757 (N_36757,N_32981,N_34768);
nor U36758 (N_36758,N_34636,N_34522);
xor U36759 (N_36759,N_33645,N_34575);
nor U36760 (N_36760,N_33244,N_33666);
or U36761 (N_36761,N_32563,N_33187);
or U36762 (N_36762,N_33051,N_34313);
nand U36763 (N_36763,N_34273,N_32787);
nand U36764 (N_36764,N_33140,N_33178);
xor U36765 (N_36765,N_34121,N_33258);
xnor U36766 (N_36766,N_32908,N_34449);
xor U36767 (N_36767,N_34354,N_33872);
nor U36768 (N_36768,N_33227,N_33660);
or U36769 (N_36769,N_33092,N_33237);
nor U36770 (N_36770,N_33675,N_34722);
xor U36771 (N_36771,N_34973,N_33158);
nor U36772 (N_36772,N_33392,N_33866);
nand U36773 (N_36773,N_34393,N_33027);
or U36774 (N_36774,N_33507,N_32880);
nand U36775 (N_36775,N_32644,N_32526);
nand U36776 (N_36776,N_34284,N_33159);
or U36777 (N_36777,N_34549,N_33620);
and U36778 (N_36778,N_33054,N_33794);
xor U36779 (N_36779,N_33844,N_34296);
and U36780 (N_36780,N_32734,N_33446);
xor U36781 (N_36781,N_32852,N_34631);
or U36782 (N_36782,N_32882,N_33578);
xnor U36783 (N_36783,N_33436,N_34809);
and U36784 (N_36784,N_34584,N_33639);
or U36785 (N_36785,N_34549,N_34048);
nand U36786 (N_36786,N_34803,N_34599);
or U36787 (N_36787,N_32820,N_34291);
nand U36788 (N_36788,N_33123,N_33247);
and U36789 (N_36789,N_33944,N_33927);
or U36790 (N_36790,N_34493,N_34843);
nor U36791 (N_36791,N_32768,N_34254);
nand U36792 (N_36792,N_33305,N_34825);
or U36793 (N_36793,N_33674,N_33990);
xnor U36794 (N_36794,N_34570,N_34537);
and U36795 (N_36795,N_33598,N_33610);
xor U36796 (N_36796,N_34006,N_34768);
nand U36797 (N_36797,N_34531,N_33119);
nor U36798 (N_36798,N_34113,N_33485);
nand U36799 (N_36799,N_33623,N_33421);
or U36800 (N_36800,N_32794,N_34320);
nand U36801 (N_36801,N_33850,N_34416);
nand U36802 (N_36802,N_33906,N_33834);
or U36803 (N_36803,N_33891,N_32852);
and U36804 (N_36804,N_34368,N_34909);
nor U36805 (N_36805,N_34261,N_33606);
xnor U36806 (N_36806,N_33123,N_34339);
xnor U36807 (N_36807,N_34632,N_34782);
nor U36808 (N_36808,N_33346,N_33465);
or U36809 (N_36809,N_32502,N_34026);
xnor U36810 (N_36810,N_32991,N_33543);
xor U36811 (N_36811,N_33317,N_33592);
nand U36812 (N_36812,N_33040,N_33909);
xnor U36813 (N_36813,N_33678,N_33939);
nand U36814 (N_36814,N_32770,N_34893);
or U36815 (N_36815,N_32587,N_34034);
xor U36816 (N_36816,N_33234,N_34934);
nor U36817 (N_36817,N_34813,N_34554);
nand U36818 (N_36818,N_33620,N_34273);
and U36819 (N_36819,N_33407,N_33025);
nor U36820 (N_36820,N_34970,N_34566);
nand U36821 (N_36821,N_32919,N_33307);
nor U36822 (N_36822,N_34739,N_34482);
or U36823 (N_36823,N_33755,N_34011);
or U36824 (N_36824,N_32813,N_34060);
and U36825 (N_36825,N_34158,N_32973);
or U36826 (N_36826,N_33593,N_32936);
or U36827 (N_36827,N_32996,N_32537);
nor U36828 (N_36828,N_34066,N_33839);
xnor U36829 (N_36829,N_34490,N_33702);
and U36830 (N_36830,N_32952,N_33819);
nor U36831 (N_36831,N_34983,N_32589);
nor U36832 (N_36832,N_32591,N_33377);
xnor U36833 (N_36833,N_34403,N_33547);
xnor U36834 (N_36834,N_34016,N_34626);
nor U36835 (N_36835,N_34328,N_33240);
nand U36836 (N_36836,N_33905,N_33265);
or U36837 (N_36837,N_32846,N_34004);
or U36838 (N_36838,N_34510,N_32645);
xnor U36839 (N_36839,N_34877,N_33503);
nor U36840 (N_36840,N_33416,N_33080);
nor U36841 (N_36841,N_32786,N_34408);
nand U36842 (N_36842,N_33366,N_33267);
or U36843 (N_36843,N_33269,N_32819);
nor U36844 (N_36844,N_34236,N_32523);
and U36845 (N_36845,N_34907,N_34653);
or U36846 (N_36846,N_32501,N_34396);
nor U36847 (N_36847,N_33597,N_33111);
or U36848 (N_36848,N_32904,N_32542);
nor U36849 (N_36849,N_34224,N_33402);
xor U36850 (N_36850,N_33629,N_34481);
and U36851 (N_36851,N_34925,N_34530);
nor U36852 (N_36852,N_32810,N_33531);
nand U36853 (N_36853,N_33339,N_33512);
or U36854 (N_36854,N_33825,N_34678);
nand U36855 (N_36855,N_34196,N_32775);
nor U36856 (N_36856,N_33383,N_32997);
xor U36857 (N_36857,N_32860,N_33872);
nand U36858 (N_36858,N_33742,N_34270);
or U36859 (N_36859,N_33434,N_34041);
nor U36860 (N_36860,N_34301,N_33250);
and U36861 (N_36861,N_34533,N_33799);
xor U36862 (N_36862,N_33718,N_34830);
xor U36863 (N_36863,N_33137,N_33689);
or U36864 (N_36864,N_33165,N_33532);
nor U36865 (N_36865,N_34100,N_33530);
or U36866 (N_36866,N_32706,N_34216);
nor U36867 (N_36867,N_34598,N_34033);
or U36868 (N_36868,N_33529,N_32922);
and U36869 (N_36869,N_33442,N_34150);
nor U36870 (N_36870,N_34866,N_32606);
and U36871 (N_36871,N_34140,N_32791);
and U36872 (N_36872,N_34970,N_33237);
and U36873 (N_36873,N_33307,N_34333);
and U36874 (N_36874,N_34490,N_34471);
or U36875 (N_36875,N_33266,N_34416);
and U36876 (N_36876,N_34286,N_33124);
or U36877 (N_36877,N_33282,N_34842);
or U36878 (N_36878,N_34430,N_33521);
or U36879 (N_36879,N_34804,N_33067);
and U36880 (N_36880,N_34427,N_34652);
xnor U36881 (N_36881,N_33326,N_34933);
and U36882 (N_36882,N_33083,N_34636);
xnor U36883 (N_36883,N_34785,N_33891);
and U36884 (N_36884,N_33719,N_32550);
nand U36885 (N_36885,N_32930,N_34454);
xnor U36886 (N_36886,N_34551,N_34984);
or U36887 (N_36887,N_33565,N_33366);
xor U36888 (N_36888,N_34089,N_33539);
xor U36889 (N_36889,N_32565,N_33253);
nor U36890 (N_36890,N_32688,N_34980);
nor U36891 (N_36891,N_34029,N_34889);
nand U36892 (N_36892,N_34253,N_32556);
or U36893 (N_36893,N_34134,N_33575);
and U36894 (N_36894,N_32762,N_33659);
nor U36895 (N_36895,N_34112,N_33529);
xor U36896 (N_36896,N_33809,N_33674);
or U36897 (N_36897,N_32545,N_32939);
xor U36898 (N_36898,N_33683,N_33562);
nor U36899 (N_36899,N_34827,N_34676);
or U36900 (N_36900,N_32705,N_33976);
nor U36901 (N_36901,N_34208,N_33159);
nor U36902 (N_36902,N_34796,N_33911);
and U36903 (N_36903,N_33067,N_33470);
nor U36904 (N_36904,N_33779,N_32502);
nand U36905 (N_36905,N_34353,N_32930);
or U36906 (N_36906,N_32870,N_34077);
xor U36907 (N_36907,N_33868,N_34104);
nor U36908 (N_36908,N_34465,N_32889);
and U36909 (N_36909,N_33140,N_33806);
nand U36910 (N_36910,N_33735,N_34432);
nand U36911 (N_36911,N_32615,N_34381);
and U36912 (N_36912,N_33140,N_33684);
xnor U36913 (N_36913,N_34839,N_33786);
nor U36914 (N_36914,N_32912,N_33354);
nand U36915 (N_36915,N_34466,N_34198);
nand U36916 (N_36916,N_33734,N_34823);
or U36917 (N_36917,N_33144,N_33199);
and U36918 (N_36918,N_33341,N_34476);
xor U36919 (N_36919,N_32706,N_33562);
nor U36920 (N_36920,N_33370,N_33450);
nand U36921 (N_36921,N_33430,N_33188);
and U36922 (N_36922,N_34190,N_33436);
xnor U36923 (N_36923,N_34536,N_33752);
xnor U36924 (N_36924,N_34629,N_33419);
and U36925 (N_36925,N_33256,N_33518);
xnor U36926 (N_36926,N_32627,N_32633);
or U36927 (N_36927,N_34057,N_33644);
and U36928 (N_36928,N_34874,N_33506);
or U36929 (N_36929,N_33079,N_33070);
nand U36930 (N_36930,N_33199,N_33476);
or U36931 (N_36931,N_32685,N_33701);
nor U36932 (N_36932,N_33817,N_33776);
nand U36933 (N_36933,N_33585,N_34482);
and U36934 (N_36934,N_34214,N_34994);
nor U36935 (N_36935,N_33732,N_33807);
nor U36936 (N_36936,N_34281,N_33476);
nor U36937 (N_36937,N_34440,N_34388);
nor U36938 (N_36938,N_33291,N_33323);
nand U36939 (N_36939,N_33878,N_33241);
xnor U36940 (N_36940,N_32728,N_33009);
nand U36941 (N_36941,N_33261,N_33554);
nand U36942 (N_36942,N_33819,N_34390);
or U36943 (N_36943,N_33692,N_32929);
nor U36944 (N_36944,N_34856,N_33305);
or U36945 (N_36945,N_34036,N_34197);
nand U36946 (N_36946,N_33649,N_32560);
xnor U36947 (N_36947,N_32569,N_32976);
nor U36948 (N_36948,N_33596,N_34628);
xor U36949 (N_36949,N_33356,N_34611);
or U36950 (N_36950,N_34471,N_34820);
nand U36951 (N_36951,N_32909,N_34433);
nor U36952 (N_36952,N_32861,N_34020);
nand U36953 (N_36953,N_33998,N_34653);
xnor U36954 (N_36954,N_33494,N_33068);
xor U36955 (N_36955,N_34480,N_34734);
nor U36956 (N_36956,N_34621,N_34455);
or U36957 (N_36957,N_33657,N_34881);
xnor U36958 (N_36958,N_34081,N_32558);
nand U36959 (N_36959,N_33340,N_34776);
nand U36960 (N_36960,N_34383,N_34269);
and U36961 (N_36961,N_34568,N_34685);
and U36962 (N_36962,N_32616,N_33775);
or U36963 (N_36963,N_32657,N_32903);
and U36964 (N_36964,N_33154,N_34252);
xor U36965 (N_36965,N_33890,N_33471);
and U36966 (N_36966,N_34521,N_34215);
or U36967 (N_36967,N_33784,N_32652);
and U36968 (N_36968,N_32844,N_34394);
and U36969 (N_36969,N_34975,N_34062);
and U36970 (N_36970,N_34991,N_33428);
or U36971 (N_36971,N_34706,N_33154);
nor U36972 (N_36972,N_32558,N_33606);
and U36973 (N_36973,N_34817,N_34269);
nand U36974 (N_36974,N_34902,N_34195);
xor U36975 (N_36975,N_33671,N_33555);
or U36976 (N_36976,N_34607,N_33426);
xor U36977 (N_36977,N_34511,N_33246);
nor U36978 (N_36978,N_33140,N_33674);
or U36979 (N_36979,N_34042,N_32638);
nand U36980 (N_36980,N_33841,N_34132);
nand U36981 (N_36981,N_34100,N_33988);
nand U36982 (N_36982,N_34129,N_34174);
xnor U36983 (N_36983,N_34707,N_34705);
nor U36984 (N_36984,N_34190,N_33655);
xor U36985 (N_36985,N_34318,N_34238);
and U36986 (N_36986,N_33432,N_32544);
or U36987 (N_36987,N_33253,N_32788);
nand U36988 (N_36988,N_34196,N_32844);
or U36989 (N_36989,N_33280,N_33993);
and U36990 (N_36990,N_34869,N_33206);
nor U36991 (N_36991,N_34835,N_34148);
nor U36992 (N_36992,N_33323,N_34171);
xnor U36993 (N_36993,N_34391,N_34467);
and U36994 (N_36994,N_34051,N_33785);
xnor U36995 (N_36995,N_34832,N_34489);
or U36996 (N_36996,N_33439,N_33901);
nand U36997 (N_36997,N_33482,N_33682);
or U36998 (N_36998,N_34060,N_33348);
or U36999 (N_36999,N_34366,N_32941);
nor U37000 (N_37000,N_33106,N_34303);
xnor U37001 (N_37001,N_33881,N_34315);
nand U37002 (N_37002,N_34202,N_33950);
or U37003 (N_37003,N_32995,N_34848);
nor U37004 (N_37004,N_33214,N_34152);
xor U37005 (N_37005,N_34191,N_33026);
nand U37006 (N_37006,N_34033,N_34068);
and U37007 (N_37007,N_32708,N_33756);
nand U37008 (N_37008,N_34289,N_32964);
or U37009 (N_37009,N_32732,N_32981);
nor U37010 (N_37010,N_33498,N_34318);
xnor U37011 (N_37011,N_33034,N_34212);
xor U37012 (N_37012,N_33200,N_34315);
nand U37013 (N_37013,N_34141,N_34037);
xor U37014 (N_37014,N_34937,N_33775);
nor U37015 (N_37015,N_34370,N_33981);
or U37016 (N_37016,N_34905,N_34593);
xnor U37017 (N_37017,N_34407,N_34205);
nor U37018 (N_37018,N_33575,N_34324);
or U37019 (N_37019,N_32710,N_33643);
nor U37020 (N_37020,N_32877,N_33329);
and U37021 (N_37021,N_34112,N_33479);
and U37022 (N_37022,N_32710,N_34950);
nor U37023 (N_37023,N_32918,N_33364);
xnor U37024 (N_37024,N_34716,N_33130);
nor U37025 (N_37025,N_33910,N_33543);
and U37026 (N_37026,N_34805,N_33313);
and U37027 (N_37027,N_34575,N_33935);
or U37028 (N_37028,N_33806,N_32951);
nor U37029 (N_37029,N_32718,N_33695);
nor U37030 (N_37030,N_33075,N_34847);
nor U37031 (N_37031,N_33001,N_33581);
xnor U37032 (N_37032,N_34209,N_34016);
or U37033 (N_37033,N_33622,N_34461);
nor U37034 (N_37034,N_34592,N_32556);
or U37035 (N_37035,N_34937,N_33337);
nor U37036 (N_37036,N_34634,N_34867);
nand U37037 (N_37037,N_34314,N_33463);
or U37038 (N_37038,N_32954,N_32766);
xor U37039 (N_37039,N_34820,N_33774);
and U37040 (N_37040,N_34929,N_33486);
nand U37041 (N_37041,N_33291,N_33398);
and U37042 (N_37042,N_32690,N_32837);
xor U37043 (N_37043,N_33701,N_32530);
nand U37044 (N_37044,N_33229,N_34070);
nor U37045 (N_37045,N_33013,N_32544);
nor U37046 (N_37046,N_34425,N_33583);
or U37047 (N_37047,N_32763,N_34983);
xnor U37048 (N_37048,N_34537,N_33789);
xnor U37049 (N_37049,N_33222,N_34237);
nor U37050 (N_37050,N_34675,N_33617);
xor U37051 (N_37051,N_33541,N_33282);
nand U37052 (N_37052,N_32664,N_34244);
or U37053 (N_37053,N_34756,N_33225);
xnor U37054 (N_37054,N_34296,N_33777);
xnor U37055 (N_37055,N_33615,N_33152);
and U37056 (N_37056,N_32663,N_33963);
nor U37057 (N_37057,N_34486,N_34707);
xnor U37058 (N_37058,N_33244,N_33706);
and U37059 (N_37059,N_34861,N_34892);
or U37060 (N_37060,N_34783,N_34809);
xor U37061 (N_37061,N_33066,N_33131);
nor U37062 (N_37062,N_33707,N_34884);
and U37063 (N_37063,N_34049,N_32690);
and U37064 (N_37064,N_34401,N_33201);
xnor U37065 (N_37065,N_34202,N_34153);
or U37066 (N_37066,N_32877,N_33780);
or U37067 (N_37067,N_32513,N_34382);
and U37068 (N_37068,N_34148,N_33191);
or U37069 (N_37069,N_33349,N_33226);
or U37070 (N_37070,N_32503,N_34957);
nor U37071 (N_37071,N_32622,N_34459);
xor U37072 (N_37072,N_32810,N_33210);
xnor U37073 (N_37073,N_33378,N_33644);
and U37074 (N_37074,N_33911,N_33342);
xnor U37075 (N_37075,N_33376,N_34080);
or U37076 (N_37076,N_34043,N_34084);
nand U37077 (N_37077,N_34638,N_34295);
nand U37078 (N_37078,N_32818,N_34747);
nand U37079 (N_37079,N_34691,N_33016);
nor U37080 (N_37080,N_34780,N_34537);
xor U37081 (N_37081,N_32583,N_32793);
and U37082 (N_37082,N_34253,N_33504);
or U37083 (N_37083,N_33512,N_34154);
xnor U37084 (N_37084,N_33939,N_34724);
xnor U37085 (N_37085,N_34726,N_33025);
nor U37086 (N_37086,N_34755,N_32720);
nor U37087 (N_37087,N_32731,N_33126);
nor U37088 (N_37088,N_34847,N_33596);
or U37089 (N_37089,N_34725,N_32938);
and U37090 (N_37090,N_33094,N_32831);
nor U37091 (N_37091,N_33399,N_33756);
nand U37092 (N_37092,N_34162,N_32632);
and U37093 (N_37093,N_33114,N_34603);
and U37094 (N_37094,N_34664,N_34477);
and U37095 (N_37095,N_33130,N_32964);
nor U37096 (N_37096,N_34295,N_34838);
and U37097 (N_37097,N_33401,N_34876);
and U37098 (N_37098,N_33618,N_34375);
nor U37099 (N_37099,N_33717,N_33342);
and U37100 (N_37100,N_34411,N_33069);
nor U37101 (N_37101,N_33321,N_34234);
or U37102 (N_37102,N_34187,N_32810);
xor U37103 (N_37103,N_32626,N_32792);
nor U37104 (N_37104,N_34649,N_33284);
nand U37105 (N_37105,N_34038,N_33947);
nand U37106 (N_37106,N_34667,N_34072);
and U37107 (N_37107,N_32566,N_34587);
nand U37108 (N_37108,N_34254,N_34497);
and U37109 (N_37109,N_33915,N_33445);
xor U37110 (N_37110,N_33818,N_34443);
or U37111 (N_37111,N_32901,N_33209);
nor U37112 (N_37112,N_33160,N_34972);
nand U37113 (N_37113,N_33992,N_34649);
nor U37114 (N_37114,N_33853,N_33914);
nand U37115 (N_37115,N_33198,N_33925);
and U37116 (N_37116,N_34169,N_34700);
xnor U37117 (N_37117,N_34671,N_34706);
nor U37118 (N_37118,N_34833,N_34218);
xnor U37119 (N_37119,N_34898,N_32707);
xor U37120 (N_37120,N_32666,N_33310);
xnor U37121 (N_37121,N_34112,N_33943);
or U37122 (N_37122,N_34158,N_34463);
xnor U37123 (N_37123,N_33124,N_33784);
or U37124 (N_37124,N_32765,N_34226);
nand U37125 (N_37125,N_33549,N_32668);
and U37126 (N_37126,N_34520,N_33968);
nor U37127 (N_37127,N_32511,N_33071);
and U37128 (N_37128,N_33420,N_33793);
nor U37129 (N_37129,N_34750,N_33132);
or U37130 (N_37130,N_34318,N_33037);
or U37131 (N_37131,N_33210,N_32842);
or U37132 (N_37132,N_33565,N_34520);
or U37133 (N_37133,N_33055,N_33249);
nand U37134 (N_37134,N_34054,N_34209);
nand U37135 (N_37135,N_33054,N_34533);
nand U37136 (N_37136,N_34845,N_34032);
nand U37137 (N_37137,N_32794,N_32909);
xor U37138 (N_37138,N_32570,N_33218);
nand U37139 (N_37139,N_33108,N_33693);
or U37140 (N_37140,N_34391,N_33739);
and U37141 (N_37141,N_34356,N_34419);
and U37142 (N_37142,N_34245,N_33082);
and U37143 (N_37143,N_34379,N_32636);
and U37144 (N_37144,N_34259,N_32784);
xnor U37145 (N_37145,N_34354,N_32889);
nand U37146 (N_37146,N_33942,N_32867);
nor U37147 (N_37147,N_33553,N_34014);
nor U37148 (N_37148,N_33102,N_33195);
or U37149 (N_37149,N_33306,N_33170);
nand U37150 (N_37150,N_33580,N_33776);
xor U37151 (N_37151,N_32877,N_34024);
xnor U37152 (N_37152,N_33440,N_34898);
or U37153 (N_37153,N_32987,N_34709);
or U37154 (N_37154,N_32852,N_32819);
or U37155 (N_37155,N_32599,N_33367);
nand U37156 (N_37156,N_33164,N_34642);
nor U37157 (N_37157,N_32873,N_33410);
nand U37158 (N_37158,N_33055,N_32586);
and U37159 (N_37159,N_34717,N_32647);
and U37160 (N_37160,N_33939,N_33494);
or U37161 (N_37161,N_34801,N_33631);
nand U37162 (N_37162,N_33750,N_32527);
or U37163 (N_37163,N_34936,N_33525);
or U37164 (N_37164,N_34600,N_34660);
xnor U37165 (N_37165,N_33985,N_34549);
xor U37166 (N_37166,N_32729,N_34818);
nand U37167 (N_37167,N_34855,N_33514);
nand U37168 (N_37168,N_32658,N_32559);
and U37169 (N_37169,N_34731,N_32847);
xnor U37170 (N_37170,N_34275,N_32721);
nor U37171 (N_37171,N_34568,N_34458);
and U37172 (N_37172,N_33318,N_33128);
or U37173 (N_37173,N_34122,N_34888);
and U37174 (N_37174,N_33588,N_33421);
nand U37175 (N_37175,N_32901,N_34555);
or U37176 (N_37176,N_32959,N_34494);
and U37177 (N_37177,N_33111,N_34995);
xor U37178 (N_37178,N_34908,N_32912);
xor U37179 (N_37179,N_34908,N_32847);
and U37180 (N_37180,N_34455,N_33511);
nand U37181 (N_37181,N_32870,N_34311);
or U37182 (N_37182,N_33858,N_34696);
nand U37183 (N_37183,N_34579,N_34892);
and U37184 (N_37184,N_34387,N_33000);
xnor U37185 (N_37185,N_34631,N_34376);
or U37186 (N_37186,N_33001,N_34797);
nand U37187 (N_37187,N_33465,N_33815);
nor U37188 (N_37188,N_32999,N_33763);
nor U37189 (N_37189,N_33539,N_34275);
nand U37190 (N_37190,N_33362,N_32700);
or U37191 (N_37191,N_34601,N_32726);
nand U37192 (N_37192,N_33896,N_33301);
and U37193 (N_37193,N_33193,N_34503);
nor U37194 (N_37194,N_33823,N_34974);
nand U37195 (N_37195,N_32621,N_33445);
or U37196 (N_37196,N_33773,N_33993);
nand U37197 (N_37197,N_32513,N_34062);
xnor U37198 (N_37198,N_34434,N_34555);
nor U37199 (N_37199,N_34867,N_33178);
nand U37200 (N_37200,N_33703,N_32621);
nand U37201 (N_37201,N_33449,N_34675);
and U37202 (N_37202,N_33570,N_32502);
xor U37203 (N_37203,N_34353,N_34394);
nand U37204 (N_37204,N_32866,N_34505);
or U37205 (N_37205,N_32502,N_32852);
xnor U37206 (N_37206,N_32972,N_32555);
or U37207 (N_37207,N_33854,N_32805);
nor U37208 (N_37208,N_32552,N_33221);
nor U37209 (N_37209,N_33505,N_34232);
xor U37210 (N_37210,N_34115,N_34089);
nor U37211 (N_37211,N_34666,N_34493);
and U37212 (N_37212,N_33367,N_32593);
xnor U37213 (N_37213,N_33230,N_33795);
xnor U37214 (N_37214,N_33053,N_34518);
nor U37215 (N_37215,N_33378,N_32654);
nor U37216 (N_37216,N_32943,N_33351);
and U37217 (N_37217,N_34279,N_33630);
and U37218 (N_37218,N_33570,N_32849);
nor U37219 (N_37219,N_34690,N_34731);
nand U37220 (N_37220,N_33761,N_33393);
nor U37221 (N_37221,N_33069,N_33714);
nor U37222 (N_37222,N_33487,N_32859);
or U37223 (N_37223,N_34052,N_33654);
nor U37224 (N_37224,N_33459,N_33169);
and U37225 (N_37225,N_34866,N_32826);
xnor U37226 (N_37226,N_34622,N_32600);
and U37227 (N_37227,N_34042,N_33886);
xnor U37228 (N_37228,N_32967,N_34427);
nand U37229 (N_37229,N_33178,N_33958);
nand U37230 (N_37230,N_34550,N_33969);
nor U37231 (N_37231,N_32585,N_34865);
nand U37232 (N_37232,N_33051,N_32585);
nand U37233 (N_37233,N_32767,N_33294);
or U37234 (N_37234,N_34945,N_33738);
and U37235 (N_37235,N_32823,N_33195);
nor U37236 (N_37236,N_34690,N_34540);
xor U37237 (N_37237,N_33508,N_33845);
or U37238 (N_37238,N_34772,N_33577);
and U37239 (N_37239,N_33551,N_34149);
xnor U37240 (N_37240,N_33095,N_32652);
and U37241 (N_37241,N_34476,N_32991);
or U37242 (N_37242,N_33869,N_34434);
xnor U37243 (N_37243,N_32525,N_34724);
xnor U37244 (N_37244,N_32677,N_33385);
nand U37245 (N_37245,N_33588,N_34447);
or U37246 (N_37246,N_33611,N_34932);
nor U37247 (N_37247,N_34277,N_33742);
xnor U37248 (N_37248,N_33097,N_32584);
xnor U37249 (N_37249,N_34944,N_33806);
nor U37250 (N_37250,N_33468,N_33700);
and U37251 (N_37251,N_32773,N_33823);
nor U37252 (N_37252,N_32666,N_34439);
or U37253 (N_37253,N_33598,N_32802);
nor U37254 (N_37254,N_33227,N_32680);
nor U37255 (N_37255,N_33796,N_34673);
and U37256 (N_37256,N_33428,N_33981);
nand U37257 (N_37257,N_32788,N_34976);
nor U37258 (N_37258,N_32743,N_33437);
or U37259 (N_37259,N_34712,N_32564);
or U37260 (N_37260,N_33788,N_33249);
or U37261 (N_37261,N_34881,N_32625);
and U37262 (N_37262,N_33181,N_33046);
xor U37263 (N_37263,N_33913,N_33687);
or U37264 (N_37264,N_32967,N_34130);
or U37265 (N_37265,N_34478,N_33484);
and U37266 (N_37266,N_32809,N_33653);
xor U37267 (N_37267,N_34200,N_34009);
xnor U37268 (N_37268,N_33983,N_33209);
nand U37269 (N_37269,N_33137,N_33339);
nor U37270 (N_37270,N_33220,N_33048);
or U37271 (N_37271,N_33953,N_33754);
or U37272 (N_37272,N_34504,N_34277);
and U37273 (N_37273,N_33755,N_33413);
nor U37274 (N_37274,N_33796,N_33087);
xnor U37275 (N_37275,N_33237,N_34874);
and U37276 (N_37276,N_33045,N_34086);
nor U37277 (N_37277,N_33823,N_34061);
or U37278 (N_37278,N_34388,N_34213);
or U37279 (N_37279,N_32702,N_34321);
or U37280 (N_37280,N_33222,N_33157);
xor U37281 (N_37281,N_34678,N_33514);
nand U37282 (N_37282,N_32572,N_33893);
or U37283 (N_37283,N_34316,N_33187);
nor U37284 (N_37284,N_34527,N_34075);
or U37285 (N_37285,N_33938,N_33014);
nand U37286 (N_37286,N_34814,N_34039);
and U37287 (N_37287,N_33780,N_34627);
or U37288 (N_37288,N_32562,N_34001);
xor U37289 (N_37289,N_33010,N_33070);
or U37290 (N_37290,N_33805,N_34662);
nor U37291 (N_37291,N_34528,N_34985);
xnor U37292 (N_37292,N_33603,N_33269);
and U37293 (N_37293,N_33429,N_34978);
nor U37294 (N_37294,N_32546,N_34667);
xor U37295 (N_37295,N_34129,N_33062);
or U37296 (N_37296,N_33980,N_33643);
nand U37297 (N_37297,N_34173,N_34693);
nor U37298 (N_37298,N_34582,N_33587);
and U37299 (N_37299,N_33460,N_34928);
nor U37300 (N_37300,N_34189,N_33022);
xnor U37301 (N_37301,N_34174,N_32977);
nor U37302 (N_37302,N_33633,N_33412);
or U37303 (N_37303,N_33792,N_34105);
xor U37304 (N_37304,N_32629,N_34647);
or U37305 (N_37305,N_34796,N_33878);
nor U37306 (N_37306,N_33431,N_34019);
xor U37307 (N_37307,N_34494,N_32891);
xnor U37308 (N_37308,N_33034,N_34545);
xnor U37309 (N_37309,N_32599,N_34797);
or U37310 (N_37310,N_34821,N_34627);
xnor U37311 (N_37311,N_33359,N_32959);
nor U37312 (N_37312,N_32756,N_33530);
and U37313 (N_37313,N_33535,N_33766);
or U37314 (N_37314,N_34379,N_34890);
xnor U37315 (N_37315,N_33119,N_33261);
or U37316 (N_37316,N_33947,N_34355);
nand U37317 (N_37317,N_32702,N_33600);
nor U37318 (N_37318,N_34624,N_33998);
nor U37319 (N_37319,N_34940,N_34562);
and U37320 (N_37320,N_34628,N_33046);
xnor U37321 (N_37321,N_33798,N_34979);
nand U37322 (N_37322,N_34086,N_34486);
nor U37323 (N_37323,N_34758,N_32802);
nand U37324 (N_37324,N_32898,N_32560);
xnor U37325 (N_37325,N_32897,N_32599);
or U37326 (N_37326,N_32794,N_32590);
nor U37327 (N_37327,N_33177,N_34561);
nand U37328 (N_37328,N_34181,N_34804);
xnor U37329 (N_37329,N_34357,N_34890);
xor U37330 (N_37330,N_33694,N_34150);
nor U37331 (N_37331,N_33305,N_32607);
xnor U37332 (N_37332,N_34118,N_34387);
xnor U37333 (N_37333,N_32871,N_32652);
or U37334 (N_37334,N_33628,N_33470);
nor U37335 (N_37335,N_33423,N_34279);
xnor U37336 (N_37336,N_32954,N_33277);
and U37337 (N_37337,N_34385,N_33424);
xnor U37338 (N_37338,N_33600,N_34837);
xor U37339 (N_37339,N_34489,N_33642);
and U37340 (N_37340,N_34901,N_32694);
or U37341 (N_37341,N_34990,N_33302);
or U37342 (N_37342,N_34872,N_33509);
nand U37343 (N_37343,N_33898,N_33622);
or U37344 (N_37344,N_34588,N_33111);
nor U37345 (N_37345,N_32670,N_32895);
nand U37346 (N_37346,N_34487,N_34426);
nand U37347 (N_37347,N_32537,N_34988);
nand U37348 (N_37348,N_32883,N_34411);
nor U37349 (N_37349,N_34484,N_33500);
nand U37350 (N_37350,N_33611,N_34110);
nor U37351 (N_37351,N_33900,N_33517);
xor U37352 (N_37352,N_33763,N_34204);
nor U37353 (N_37353,N_33290,N_34025);
and U37354 (N_37354,N_33535,N_34988);
and U37355 (N_37355,N_34683,N_34353);
or U37356 (N_37356,N_34532,N_34560);
xnor U37357 (N_37357,N_32717,N_34980);
xnor U37358 (N_37358,N_34043,N_34827);
nor U37359 (N_37359,N_33173,N_34472);
or U37360 (N_37360,N_33586,N_34237);
xor U37361 (N_37361,N_32828,N_32607);
nor U37362 (N_37362,N_32699,N_34948);
nor U37363 (N_37363,N_34277,N_33396);
nand U37364 (N_37364,N_34070,N_34292);
nor U37365 (N_37365,N_34314,N_33377);
nor U37366 (N_37366,N_33884,N_32688);
xnor U37367 (N_37367,N_34668,N_34594);
or U37368 (N_37368,N_33019,N_33862);
nand U37369 (N_37369,N_34598,N_33006);
nand U37370 (N_37370,N_33529,N_34625);
nand U37371 (N_37371,N_33503,N_34748);
xor U37372 (N_37372,N_33983,N_33958);
nor U37373 (N_37373,N_33917,N_33456);
and U37374 (N_37374,N_33990,N_34675);
nand U37375 (N_37375,N_32730,N_32728);
xnor U37376 (N_37376,N_33012,N_34462);
and U37377 (N_37377,N_33775,N_33086);
nand U37378 (N_37378,N_33663,N_34148);
or U37379 (N_37379,N_34546,N_32562);
xor U37380 (N_37380,N_32890,N_34360);
xor U37381 (N_37381,N_34102,N_32864);
xor U37382 (N_37382,N_34249,N_32742);
nand U37383 (N_37383,N_33279,N_32892);
or U37384 (N_37384,N_34803,N_32658);
or U37385 (N_37385,N_34778,N_33140);
and U37386 (N_37386,N_33261,N_34290);
or U37387 (N_37387,N_32773,N_33117);
nor U37388 (N_37388,N_33180,N_33810);
nor U37389 (N_37389,N_34905,N_34194);
and U37390 (N_37390,N_32742,N_33549);
nand U37391 (N_37391,N_33691,N_32852);
xor U37392 (N_37392,N_34592,N_34819);
nand U37393 (N_37393,N_33298,N_34698);
nand U37394 (N_37394,N_34973,N_33004);
nor U37395 (N_37395,N_32527,N_32505);
nand U37396 (N_37396,N_34329,N_33348);
xnor U37397 (N_37397,N_34979,N_33226);
nand U37398 (N_37398,N_33713,N_32543);
nor U37399 (N_37399,N_33032,N_33571);
or U37400 (N_37400,N_33811,N_33353);
nand U37401 (N_37401,N_32525,N_34688);
nor U37402 (N_37402,N_34318,N_32538);
nand U37403 (N_37403,N_33398,N_32938);
xnor U37404 (N_37404,N_34867,N_33386);
nand U37405 (N_37405,N_33293,N_32742);
and U37406 (N_37406,N_33765,N_33853);
nand U37407 (N_37407,N_32795,N_34509);
nand U37408 (N_37408,N_33218,N_34413);
and U37409 (N_37409,N_34689,N_34515);
or U37410 (N_37410,N_34137,N_34767);
nor U37411 (N_37411,N_34190,N_34941);
nand U37412 (N_37412,N_32930,N_33953);
or U37413 (N_37413,N_32693,N_33636);
nand U37414 (N_37414,N_33373,N_33741);
nand U37415 (N_37415,N_32922,N_33197);
xnor U37416 (N_37416,N_32601,N_33215);
or U37417 (N_37417,N_33039,N_34142);
and U37418 (N_37418,N_32965,N_34217);
nor U37419 (N_37419,N_34842,N_34562);
nor U37420 (N_37420,N_34690,N_34742);
xnor U37421 (N_37421,N_34984,N_34724);
xor U37422 (N_37422,N_34188,N_34859);
nand U37423 (N_37423,N_32511,N_33717);
nand U37424 (N_37424,N_33634,N_34920);
or U37425 (N_37425,N_32742,N_34114);
nor U37426 (N_37426,N_34989,N_33944);
and U37427 (N_37427,N_34679,N_33312);
and U37428 (N_37428,N_33484,N_32925);
and U37429 (N_37429,N_33631,N_32654);
or U37430 (N_37430,N_33087,N_33294);
nand U37431 (N_37431,N_34744,N_34730);
nand U37432 (N_37432,N_33655,N_34695);
or U37433 (N_37433,N_33003,N_34331);
nor U37434 (N_37434,N_32804,N_34690);
nand U37435 (N_37435,N_33345,N_33903);
xor U37436 (N_37436,N_32565,N_33558);
or U37437 (N_37437,N_32936,N_34466);
or U37438 (N_37438,N_33938,N_34810);
nor U37439 (N_37439,N_33517,N_33043);
and U37440 (N_37440,N_34294,N_32602);
and U37441 (N_37441,N_32729,N_34487);
xor U37442 (N_37442,N_33561,N_33477);
and U37443 (N_37443,N_33908,N_33416);
and U37444 (N_37444,N_33773,N_33688);
or U37445 (N_37445,N_34927,N_34063);
nor U37446 (N_37446,N_33817,N_33505);
nand U37447 (N_37447,N_33210,N_32947);
nor U37448 (N_37448,N_33490,N_34703);
or U37449 (N_37449,N_34384,N_34293);
xor U37450 (N_37450,N_32728,N_34869);
nand U37451 (N_37451,N_32883,N_33074);
nand U37452 (N_37452,N_33686,N_33831);
or U37453 (N_37453,N_32706,N_33369);
and U37454 (N_37454,N_34248,N_34152);
or U37455 (N_37455,N_33485,N_32517);
nor U37456 (N_37456,N_34925,N_33981);
and U37457 (N_37457,N_32564,N_33849);
and U37458 (N_37458,N_34869,N_33587);
and U37459 (N_37459,N_33333,N_34894);
and U37460 (N_37460,N_34398,N_32523);
nand U37461 (N_37461,N_33057,N_33539);
xor U37462 (N_37462,N_33238,N_34505);
nor U37463 (N_37463,N_33517,N_33730);
nor U37464 (N_37464,N_34637,N_33625);
nor U37465 (N_37465,N_33323,N_34527);
nor U37466 (N_37466,N_33736,N_32702);
and U37467 (N_37467,N_32813,N_32969);
nand U37468 (N_37468,N_34247,N_33756);
nand U37469 (N_37469,N_34037,N_33346);
or U37470 (N_37470,N_32881,N_33788);
xnor U37471 (N_37471,N_32800,N_32977);
and U37472 (N_37472,N_34856,N_33947);
and U37473 (N_37473,N_33417,N_33670);
nor U37474 (N_37474,N_34541,N_33778);
xor U37475 (N_37475,N_34644,N_32948);
nor U37476 (N_37476,N_34620,N_33186);
and U37477 (N_37477,N_33251,N_32927);
nor U37478 (N_37478,N_34590,N_32806);
nor U37479 (N_37479,N_34170,N_34787);
xnor U37480 (N_37480,N_34905,N_34663);
and U37481 (N_37481,N_34163,N_34671);
nor U37482 (N_37482,N_33848,N_34318);
nand U37483 (N_37483,N_34620,N_32534);
nand U37484 (N_37484,N_34818,N_34728);
xnor U37485 (N_37485,N_33962,N_34337);
and U37486 (N_37486,N_33092,N_34934);
nand U37487 (N_37487,N_33178,N_32826);
and U37488 (N_37488,N_34197,N_33122);
xor U37489 (N_37489,N_33180,N_34985);
nor U37490 (N_37490,N_34971,N_33758);
nor U37491 (N_37491,N_33388,N_33897);
nor U37492 (N_37492,N_34466,N_34430);
nor U37493 (N_37493,N_32607,N_33232);
or U37494 (N_37494,N_32968,N_34171);
or U37495 (N_37495,N_34481,N_33686);
or U37496 (N_37496,N_34963,N_33772);
or U37497 (N_37497,N_34621,N_32956);
and U37498 (N_37498,N_33366,N_32735);
or U37499 (N_37499,N_34668,N_32884);
nor U37500 (N_37500,N_35486,N_35622);
nand U37501 (N_37501,N_37153,N_35170);
xor U37502 (N_37502,N_37499,N_35482);
and U37503 (N_37503,N_36839,N_36586);
xnor U37504 (N_37504,N_35016,N_35708);
nor U37505 (N_37505,N_36663,N_36159);
and U37506 (N_37506,N_37148,N_35490);
or U37507 (N_37507,N_36906,N_35244);
nand U37508 (N_37508,N_36961,N_36414);
nand U37509 (N_37509,N_36108,N_35594);
xnor U37510 (N_37510,N_35242,N_37100);
and U37511 (N_37511,N_37365,N_37011);
nand U37512 (N_37512,N_35812,N_37237);
nor U37513 (N_37513,N_35727,N_36743);
and U37514 (N_37514,N_35414,N_36537);
or U37515 (N_37515,N_35760,N_36569);
xor U37516 (N_37516,N_35702,N_35293);
or U37517 (N_37517,N_37313,N_36628);
xnor U37518 (N_37518,N_36513,N_35000);
nand U37519 (N_37519,N_35834,N_35171);
or U37520 (N_37520,N_36449,N_36696);
or U37521 (N_37521,N_35221,N_35626);
nand U37522 (N_37522,N_36337,N_36500);
and U37523 (N_37523,N_36509,N_35849);
nand U37524 (N_37524,N_37381,N_35380);
nand U37525 (N_37525,N_37429,N_36323);
and U37526 (N_37526,N_36644,N_36905);
nand U37527 (N_37527,N_36465,N_36988);
nand U37528 (N_37528,N_35883,N_37210);
and U37529 (N_37529,N_35696,N_36223);
xor U37530 (N_37530,N_36258,N_35307);
or U37531 (N_37531,N_36396,N_37481);
or U37532 (N_37532,N_36630,N_36849);
nor U37533 (N_37533,N_35084,N_37293);
nand U37534 (N_37534,N_35701,N_36216);
or U37535 (N_37535,N_37027,N_36092);
xnor U37536 (N_37536,N_36318,N_35961);
or U37537 (N_37537,N_35771,N_36936);
nor U37538 (N_37538,N_35324,N_36479);
and U37539 (N_37539,N_36924,N_35851);
xnor U37540 (N_37540,N_36220,N_35593);
or U37541 (N_37541,N_36030,N_35091);
or U37542 (N_37542,N_35044,N_35030);
or U37543 (N_37543,N_36659,N_35524);
and U37544 (N_37544,N_35600,N_36554);
nor U37545 (N_37545,N_36055,N_35214);
and U37546 (N_37546,N_35734,N_36872);
and U37547 (N_37547,N_36836,N_36295);
and U37548 (N_37548,N_35423,N_37291);
and U37549 (N_37549,N_35781,N_35331);
xor U37550 (N_37550,N_35304,N_36789);
nand U37551 (N_37551,N_36247,N_36897);
nand U37552 (N_37552,N_35742,N_36448);
nand U37553 (N_37553,N_35080,N_37199);
nor U37554 (N_37554,N_36173,N_35390);
nor U37555 (N_37555,N_35346,N_35165);
nor U37556 (N_37556,N_36009,N_36062);
and U37557 (N_37557,N_35060,N_37345);
xnor U37558 (N_37558,N_36379,N_37456);
or U37559 (N_37559,N_37334,N_37059);
nor U37560 (N_37560,N_36380,N_35649);
and U37561 (N_37561,N_36437,N_36278);
or U37562 (N_37562,N_36947,N_36436);
xnor U37563 (N_37563,N_37179,N_37407);
xor U37564 (N_37564,N_36158,N_36395);
nor U37565 (N_37565,N_36548,N_37080);
xnor U37566 (N_37566,N_35180,N_36699);
nand U37567 (N_37567,N_37320,N_35713);
or U37568 (N_37568,N_35156,N_35752);
nand U37569 (N_37569,N_35351,N_37030);
nor U37570 (N_37570,N_36625,N_36672);
or U37571 (N_37571,N_36284,N_35506);
and U37572 (N_37572,N_35778,N_36384);
or U37573 (N_37573,N_36993,N_36647);
and U37574 (N_37574,N_36333,N_36958);
nand U37575 (N_37575,N_37187,N_36287);
xor U37576 (N_37576,N_35425,N_35500);
or U37577 (N_37577,N_36694,N_36937);
or U37578 (N_37578,N_36728,N_35595);
or U37579 (N_37579,N_36701,N_36512);
nand U37580 (N_37580,N_35412,N_37079);
nor U37581 (N_37581,N_36833,N_37105);
and U37582 (N_37582,N_36445,N_36332);
xnor U37583 (N_37583,N_37367,N_35850);
and U37584 (N_37584,N_36880,N_36022);
xor U37585 (N_37585,N_36397,N_37005);
xor U37586 (N_37586,N_35017,N_36996);
xnor U37587 (N_37587,N_36358,N_35858);
or U37588 (N_37588,N_35906,N_36079);
and U37589 (N_37589,N_36299,N_36067);
or U37590 (N_37590,N_36510,N_35587);
nand U37591 (N_37591,N_35375,N_36183);
xnor U37592 (N_37592,N_35509,N_35014);
or U37593 (N_37593,N_36048,N_36291);
nand U37594 (N_37594,N_35902,N_36099);
nor U37595 (N_37595,N_35202,N_36853);
xor U37596 (N_37596,N_35707,N_35886);
xnor U37597 (N_37597,N_36018,N_36264);
nor U37598 (N_37598,N_37496,N_35841);
nand U37599 (N_37599,N_36684,N_35190);
or U37600 (N_37600,N_35320,N_35249);
nor U37601 (N_37601,N_35297,N_36355);
nand U37602 (N_37602,N_35948,N_36931);
nor U37603 (N_37603,N_37375,N_35279);
nor U37604 (N_37604,N_35973,N_37023);
nand U37605 (N_37605,N_35415,N_36730);
or U37606 (N_37606,N_36967,N_35040);
and U37607 (N_37607,N_36913,N_35271);
nand U37608 (N_37608,N_36382,N_37034);
and U37609 (N_37609,N_35958,N_35686);
nand U37610 (N_37610,N_36852,N_36370);
nand U37611 (N_37611,N_35110,N_37378);
xor U37612 (N_37612,N_37006,N_35644);
and U37613 (N_37613,N_36590,N_36787);
or U37614 (N_37614,N_37019,N_37376);
and U37615 (N_37615,N_35144,N_37288);
or U37616 (N_37616,N_35892,N_36895);
xor U37617 (N_37617,N_35957,N_35462);
and U37618 (N_37618,N_36334,N_35381);
nand U37619 (N_37619,N_35558,N_36746);
or U37620 (N_37620,N_36733,N_36700);
nor U37621 (N_37621,N_37495,N_36960);
xor U37622 (N_37622,N_36035,N_36778);
and U37623 (N_37623,N_36838,N_35086);
nand U37624 (N_37624,N_36204,N_35181);
nor U37625 (N_37625,N_36547,N_37058);
nor U37626 (N_37626,N_36123,N_37168);
or U37627 (N_37627,N_37494,N_35083);
and U37628 (N_37628,N_35454,N_35981);
nor U37629 (N_37629,N_35130,N_36517);
xnor U37630 (N_37630,N_37130,N_36419);
nand U37631 (N_37631,N_37351,N_35693);
xor U37632 (N_37632,N_37016,N_37159);
xnor U37633 (N_37633,N_35164,N_35153);
and U37634 (N_37634,N_37125,N_36885);
or U37635 (N_37635,N_37163,N_36603);
and U37636 (N_37636,N_35545,N_35352);
and U37637 (N_37637,N_35769,N_36176);
or U37638 (N_37638,N_37324,N_37234);
and U37639 (N_37639,N_35431,N_36922);
xor U37640 (N_37640,N_37461,N_37092);
or U37641 (N_37641,N_36929,N_35237);
and U37642 (N_37642,N_37049,N_35345);
and U37643 (N_37643,N_36026,N_37477);
or U37644 (N_37644,N_36939,N_35263);
nand U37645 (N_37645,N_35737,N_36505);
xnor U37646 (N_37646,N_36503,N_36447);
or U37647 (N_37647,N_37215,N_35866);
and U37648 (N_37648,N_35444,N_35580);
or U37649 (N_37649,N_35688,N_35363);
nand U37650 (N_37650,N_36229,N_36955);
or U37651 (N_37651,N_35051,N_35995);
nor U37652 (N_37652,N_36105,N_37439);
or U37653 (N_37653,N_37004,N_35613);
xnor U37654 (N_37654,N_36984,N_36792);
nor U37655 (N_37655,N_35300,N_35126);
and U37656 (N_37656,N_35063,N_36935);
and U37657 (N_37657,N_36951,N_35275);
nor U37658 (N_37658,N_37222,N_36692);
and U37659 (N_37659,N_35777,N_37218);
xnor U37660 (N_37660,N_36296,N_36734);
xor U37661 (N_37661,N_35411,N_36294);
nand U37662 (N_37662,N_35642,N_35025);
xnor U37663 (N_37663,N_36094,N_35419);
and U37664 (N_37664,N_37454,N_36226);
xor U37665 (N_37665,N_35733,N_35168);
xnor U37666 (N_37666,N_35569,N_37194);
and U37667 (N_37667,N_35321,N_36841);
or U37668 (N_37668,N_36023,N_36591);
and U37669 (N_37669,N_35420,N_36676);
nand U37670 (N_37670,N_37175,N_36653);
and U37671 (N_37671,N_35099,N_35523);
nand U37672 (N_37672,N_35229,N_36198);
nor U37673 (N_37673,N_37075,N_37240);
xor U37674 (N_37674,N_35173,N_37250);
nand U37675 (N_37675,N_35369,N_36712);
xor U37676 (N_37676,N_37015,N_35577);
xnor U37677 (N_37677,N_35325,N_37289);
nand U37678 (N_37678,N_37248,N_36462);
nand U37679 (N_37679,N_36727,N_37347);
nor U37680 (N_37680,N_35392,N_35228);
nor U37681 (N_37681,N_35714,N_36577);
nand U37682 (N_37682,N_36398,N_37343);
or U37683 (N_37683,N_35426,N_35695);
or U37684 (N_37684,N_35955,N_35950);
and U37685 (N_37685,N_36242,N_35342);
nand U37686 (N_37686,N_35937,N_35641);
xor U37687 (N_37687,N_35521,N_35944);
nand U37688 (N_37688,N_36530,N_36902);
or U37689 (N_37689,N_36430,N_36203);
xor U37690 (N_37690,N_35532,N_35504);
xnor U37691 (N_37691,N_35788,N_35184);
or U37692 (N_37692,N_37043,N_35147);
nor U37693 (N_37693,N_35605,N_37452);
and U37694 (N_37694,N_35270,N_35929);
and U37695 (N_37695,N_37236,N_35645);
and U37696 (N_37696,N_36987,N_36522);
xnor U37697 (N_37697,N_35960,N_36240);
or U37698 (N_37698,N_36453,N_35349);
nor U37699 (N_37699,N_35028,N_36946);
or U37700 (N_37700,N_37394,N_35864);
nand U37701 (N_37701,N_36361,N_37260);
or U37702 (N_37702,N_37332,N_37106);
and U37703 (N_37703,N_37189,N_37396);
and U37704 (N_37704,N_37198,N_35374);
xor U37705 (N_37705,N_36457,N_37458);
nor U37706 (N_37706,N_36589,N_37014);
xnor U37707 (N_37707,N_37449,N_36317);
or U37708 (N_37708,N_37117,N_36248);
or U37709 (N_37709,N_37197,N_36211);
nand U37710 (N_37710,N_37388,N_35138);
or U37711 (N_37711,N_35400,N_36893);
or U37712 (N_37712,N_35719,N_36871);
nand U37713 (N_37713,N_35893,N_36281);
xnor U37714 (N_37714,N_37292,N_36777);
or U37715 (N_37715,N_37055,N_35185);
nand U37716 (N_37716,N_35759,N_36473);
and U37717 (N_37717,N_35458,N_36643);
nand U37718 (N_37718,N_35983,N_35276);
nor U37719 (N_37719,N_35724,N_35783);
nor U37720 (N_37720,N_37330,N_36146);
xnor U37721 (N_37721,N_36780,N_35544);
nor U37722 (N_37722,N_36662,N_35260);
xor U37723 (N_37723,N_35042,N_37374);
xnor U37724 (N_37724,N_35552,N_37192);
nor U37725 (N_37725,N_35456,N_36186);
xor U37726 (N_37726,N_37000,N_36388);
nor U37727 (N_37727,N_36686,N_37205);
or U37728 (N_37728,N_35898,N_35232);
nor U37729 (N_37729,N_36452,N_35939);
nor U37730 (N_37730,N_35835,N_35681);
or U37731 (N_37731,N_36869,N_36840);
nand U37732 (N_37732,N_35222,N_37102);
and U37733 (N_37733,N_37123,N_35730);
or U37734 (N_37734,N_35332,N_36666);
nor U37735 (N_37735,N_36344,N_36850);
or U37736 (N_37736,N_35679,N_35732);
or U37737 (N_37737,N_36192,N_36064);
and U37738 (N_37738,N_35932,N_36650);
xnor U37739 (N_37739,N_35637,N_36466);
nor U37740 (N_37740,N_36776,N_35988);
xor U37741 (N_37741,N_36330,N_37372);
and U37742 (N_37742,N_36506,N_35007);
and U37743 (N_37743,N_35453,N_36516);
or U37744 (N_37744,N_36335,N_36962);
or U37745 (N_37745,N_36017,N_35011);
nor U37746 (N_37746,N_37410,N_37480);
nand U37747 (N_37747,N_37277,N_37151);
xor U37748 (N_37748,N_35852,N_35853);
nand U37749 (N_37749,N_35430,N_37138);
and U37750 (N_37750,N_36868,N_36491);
xor U37751 (N_37751,N_35478,N_35823);
xor U37752 (N_37752,N_36289,N_35290);
nor U37753 (N_37753,N_36934,N_37437);
nor U37754 (N_37754,N_36280,N_36218);
nor U37755 (N_37755,N_36260,N_36718);
nor U37756 (N_37756,N_37309,N_37074);
nor U37757 (N_37757,N_35817,N_35876);
and U37758 (N_37758,N_36201,N_35818);
nor U37759 (N_37759,N_36660,N_36115);
or U37760 (N_37760,N_35703,N_36940);
and U37761 (N_37761,N_35654,N_37223);
xor U37762 (N_37762,N_35361,N_35863);
nor U37763 (N_37763,N_35251,N_35029);
nor U37764 (N_37764,N_36713,N_36570);
xor U37765 (N_37765,N_35457,N_36910);
or U37766 (N_37766,N_36781,N_35770);
or U37767 (N_37767,N_36894,N_36326);
nor U37768 (N_37768,N_36230,N_36302);
xnor U37769 (N_37769,N_35330,N_35034);
or U37770 (N_37770,N_36610,N_36339);
xor U37771 (N_37771,N_35758,N_36188);
and U37772 (N_37772,N_35924,N_37149);
or U37773 (N_37773,N_35385,N_35881);
nor U37774 (N_37774,N_36024,N_35699);
and U37775 (N_37775,N_36494,N_35623);
xor U37776 (N_37776,N_35704,N_36273);
or U37777 (N_37777,N_35306,N_37209);
nand U37778 (N_37778,N_35317,N_35940);
nor U37779 (N_37779,N_37354,N_36304);
xor U37780 (N_37780,N_36764,N_36974);
and U37781 (N_37781,N_36328,N_36954);
or U37782 (N_37782,N_35434,N_35046);
or U37783 (N_37783,N_35553,N_35090);
or U37784 (N_37784,N_36948,N_37084);
or U37785 (N_37785,N_35551,N_36131);
nor U37786 (N_37786,N_37098,N_36106);
nor U37787 (N_37787,N_36008,N_37232);
or U37788 (N_37788,N_36957,N_36862);
or U37789 (N_37789,N_36531,N_36147);
and U37790 (N_37790,N_36903,N_36275);
and U37791 (N_37791,N_37185,N_35339);
xor U37792 (N_37792,N_35808,N_37196);
and U37793 (N_37793,N_36896,N_35394);
or U37794 (N_37794,N_37263,N_35927);
nor U37795 (N_37795,N_37206,N_36674);
nor U37796 (N_37796,N_36995,N_35459);
nor U37797 (N_37797,N_35511,N_36200);
xor U37798 (N_37798,N_35735,N_37436);
and U37799 (N_37799,N_35149,N_37344);
or U37800 (N_37800,N_36907,N_37217);
xor U37801 (N_37801,N_36126,N_37107);
xnor U37802 (N_37802,N_36439,N_36593);
and U37803 (N_37803,N_35057,N_36276);
and U37804 (N_37804,N_35574,N_36341);
and U37805 (N_37805,N_37406,N_35418);
xor U37806 (N_37806,N_36464,N_37170);
or U37807 (N_37807,N_37304,N_37285);
nand U37808 (N_37808,N_37352,N_35452);
nand U37809 (N_37809,N_37216,N_37298);
or U37810 (N_37810,N_35716,N_36690);
nor U37811 (N_37811,N_36865,N_35145);
xor U37812 (N_37812,N_35987,N_36511);
xor U37813 (N_37813,N_35685,N_35048);
and U37814 (N_37814,N_35065,N_35903);
and U37815 (N_37815,N_36056,N_35360);
xnor U37816 (N_37816,N_36071,N_36357);
and U37817 (N_37817,N_36160,N_35656);
nand U37818 (N_37818,N_36536,N_35442);
or U37819 (N_37819,N_35982,N_35373);
nor U37820 (N_37820,N_35287,N_35137);
nand U37821 (N_37821,N_35053,N_35061);
xnor U37822 (N_37822,N_36648,N_35520);
and U37823 (N_37823,N_37174,N_35108);
nand U37824 (N_37824,N_35277,N_35632);
and U37825 (N_37825,N_36375,N_35526);
xor U37826 (N_37826,N_36288,N_37362);
or U37827 (N_37827,N_35246,N_35250);
xnor U37828 (N_37828,N_36976,N_37275);
and U37829 (N_37829,N_36261,N_37204);
or U37830 (N_37830,N_36167,N_36454);
nand U37831 (N_37831,N_35474,N_36773);
nand U37832 (N_37832,N_36061,N_36799);
nor U37833 (N_37833,N_35548,N_36816);
nand U37834 (N_37834,N_35041,N_36639);
and U37835 (N_37835,N_36981,N_35611);
nand U37836 (N_37836,N_35281,N_36524);
xor U37837 (N_37837,N_35743,N_36544);
or U37838 (N_37838,N_35744,N_36274);
xnor U37839 (N_37839,N_35494,N_37096);
nand U37840 (N_37840,N_36615,N_35118);
xor U37841 (N_37841,N_35436,N_36424);
nand U37842 (N_37842,N_35248,N_35806);
nor U37843 (N_37843,N_36087,N_37126);
xor U37844 (N_37844,N_36795,N_35591);
nand U37845 (N_37845,N_37225,N_36942);
xor U37846 (N_37846,N_37311,N_35493);
and U37847 (N_37847,N_35427,N_35289);
and U37848 (N_37848,N_35085,N_35407);
nor U37849 (N_37849,N_36233,N_35282);
nor U37850 (N_37850,N_36316,N_36033);
nand U37851 (N_37851,N_35070,N_35023);
or U37852 (N_37852,N_36980,N_35675);
nor U37853 (N_37853,N_36459,N_37104);
nand U37854 (N_37854,N_37093,N_35329);
and U37855 (N_37855,N_36169,N_35563);
nor U37856 (N_37856,N_36587,N_37120);
xor U37857 (N_37857,N_36352,N_35288);
xnor U37858 (N_37858,N_37331,N_37097);
or U37859 (N_37859,N_36691,N_35069);
and U37860 (N_37860,N_35174,N_37132);
and U37861 (N_37861,N_35844,N_35295);
nand U37862 (N_37862,N_36290,N_37254);
xnor U37863 (N_37863,N_36138,N_36257);
and U37864 (N_37864,N_36750,N_36673);
nand U37865 (N_37865,N_36228,N_36665);
xnor U37866 (N_37866,N_37397,N_36259);
xnor U37867 (N_37867,N_35421,N_35824);
or U37868 (N_37868,N_36710,N_36025);
nand U37869 (N_37869,N_35837,N_35203);
nor U37870 (N_37870,N_36622,N_36363);
nor U37871 (N_37871,N_35609,N_35896);
and U37872 (N_37872,N_35723,N_36911);
or U37873 (N_37873,N_36919,N_36721);
nor U37874 (N_37874,N_36137,N_36580);
and U37875 (N_37875,N_36181,N_36110);
nand U37876 (N_37876,N_36213,N_36132);
xor U37877 (N_37877,N_36786,N_36772);
xnor U37878 (N_37878,N_36251,N_35155);
xnor U37879 (N_37879,N_35314,N_35861);
xor U37880 (N_37880,N_36740,N_36508);
xnor U37881 (N_37881,N_35183,N_36645);
or U37882 (N_37882,N_35113,N_37061);
nor U37883 (N_37883,N_35334,N_35001);
or U37884 (N_37884,N_36783,N_35537);
nand U37885 (N_37885,N_36068,N_35867);
nand U37886 (N_37886,N_35634,N_35738);
nor U37887 (N_37887,N_35800,N_37425);
or U37888 (N_37888,N_36835,N_36324);
xor U37889 (N_37889,N_35140,N_37270);
and U37890 (N_37890,N_36262,N_36163);
nor U37891 (N_37891,N_37228,N_37143);
nand U37892 (N_37892,N_37101,N_36256);
or U37893 (N_37893,N_36313,N_35316);
nor U37894 (N_37894,N_36704,N_37337);
nor U37895 (N_37895,N_36152,N_35404);
and U37896 (N_37896,N_35608,N_35231);
nor U37897 (N_37897,N_37094,N_37252);
nand U37898 (N_37898,N_36250,N_35968);
nand U37899 (N_37899,N_37114,N_37068);
nand U37900 (N_37900,N_36528,N_35590);
nor U37901 (N_37901,N_36303,N_37238);
xnor U37902 (N_37902,N_35151,N_36754);
or U37903 (N_37903,N_36134,N_35488);
xor U37904 (N_37904,N_35446,N_35996);
or U37905 (N_37905,N_35116,N_36121);
and U37906 (N_37906,N_36971,N_37490);
nor U37907 (N_37907,N_37150,N_35215);
nand U37908 (N_37908,N_37326,N_35167);
nor U37909 (N_37909,N_36101,N_36706);
xor U37910 (N_37910,N_36093,N_35472);
nor U37911 (N_37911,N_37071,N_36097);
and U37912 (N_37912,N_35507,N_36107);
nor U37913 (N_37913,N_36345,N_35963);
or U37914 (N_37914,N_37111,N_37340);
xnor U37915 (N_37915,N_35751,N_37284);
xor U37916 (N_37916,N_35801,N_37133);
or U37917 (N_37917,N_35344,N_35935);
xor U37918 (N_37918,N_36966,N_36373);
xor U37919 (N_37919,N_35437,N_35554);
nor U37920 (N_37920,N_37398,N_35615);
nor U37921 (N_37921,N_35252,N_37485);
nand U37922 (N_37922,N_35158,N_36535);
nand U37923 (N_37923,N_35305,N_36843);
and U37924 (N_37924,N_35739,N_35763);
and U37925 (N_37925,N_36401,N_37491);
xnor U37926 (N_37926,N_35711,N_35663);
or U37927 (N_37927,N_35677,N_36640);
or U37928 (N_37928,N_36828,N_36405);
xnor U37929 (N_37929,N_35931,N_36817);
nor U37930 (N_37930,N_36118,N_35176);
or U37931 (N_37931,N_35211,N_36847);
and U37932 (N_37932,N_35296,N_35172);
and U37933 (N_37933,N_36185,N_36771);
nand U37934 (N_37934,N_35755,N_35031);
nor U37935 (N_37935,N_37475,N_37090);
nand U37936 (N_37936,N_36305,N_35218);
xnor U37937 (N_37937,N_36117,N_35050);
and U37938 (N_37938,N_37306,N_36595);
or U37939 (N_37939,N_35217,N_35466);
xnor U37940 (N_37940,N_35791,N_35706);
nand U37941 (N_37941,N_36949,N_35710);
nand U37942 (N_37942,N_35833,N_36238);
nor U37943 (N_37943,N_36469,N_35700);
xor U37944 (N_37944,N_35018,N_35117);
nor U37945 (N_37945,N_37411,N_35367);
and U37946 (N_37946,N_37195,N_36140);
and U37947 (N_37947,N_35241,N_35756);
nor U37948 (N_37948,N_35514,N_37087);
nand U37949 (N_37949,N_35676,N_37108);
nor U37950 (N_37950,N_36112,N_36753);
or U37951 (N_37951,N_35371,N_36438);
and U37952 (N_37952,N_36716,N_37183);
nand U37953 (N_37953,N_36613,N_35536);
or U37954 (N_37954,N_35541,N_36199);
xor U37955 (N_37955,N_36202,N_35586);
and U37956 (N_37956,N_36618,N_36421);
nand U37957 (N_37957,N_35435,N_36619);
nor U37958 (N_37958,N_35002,N_35327);
nand U37959 (N_37959,N_37042,N_36815);
xnor U37960 (N_37960,N_35135,N_35341);
xor U37961 (N_37961,N_37262,N_35607);
or U37962 (N_37962,N_35888,N_35009);
nor U37963 (N_37963,N_35784,N_35439);
nand U37964 (N_37964,N_36832,N_37416);
nand U37965 (N_37965,N_36594,N_35160);
and U37966 (N_37966,N_36766,N_36492);
and U37967 (N_37967,N_36755,N_37156);
xor U37968 (N_37968,N_35887,N_35473);
and U37969 (N_37969,N_35201,N_36471);
nor U37970 (N_37970,N_36429,N_36196);
nand U37971 (N_37971,N_36001,N_36882);
nand U37972 (N_37972,N_35697,N_36737);
and U37973 (N_37973,N_36298,N_35460);
and U37974 (N_37974,N_36717,N_35429);
nor U37975 (N_37975,N_35715,N_37053);
nand U37976 (N_37976,N_35424,N_35492);
xor U37977 (N_37977,N_35772,N_35347);
nor U37978 (N_37978,N_36308,N_37013);
and U37979 (N_37979,N_35870,N_36649);
xnor U37980 (N_37980,N_36646,N_35006);
nand U37981 (N_37981,N_35964,N_36499);
and U37982 (N_37982,N_36729,N_35827);
nor U37983 (N_37983,N_36039,N_37041);
nor U37984 (N_37984,N_37115,N_37131);
and U37985 (N_37985,N_35910,N_35628);
and U37986 (N_37986,N_37468,N_36227);
xor U37987 (N_37987,N_37167,N_36616);
nor U37988 (N_37988,N_37342,N_35633);
or U37989 (N_37989,N_35326,N_36182);
nand U37990 (N_37990,N_36926,N_35401);
nand U37991 (N_37991,N_36311,N_37088);
nand U37992 (N_37992,N_37299,N_35653);
and U37993 (N_37993,N_36521,N_37338);
nor U37994 (N_37994,N_36044,N_36945);
xor U37995 (N_37995,N_36928,N_36575);
nor U37996 (N_37996,N_35779,N_37399);
xnor U37997 (N_37997,N_35816,N_36785);
nor U37998 (N_37998,N_36496,N_37349);
nor U37999 (N_37999,N_37062,N_35912);
xnor U38000 (N_38000,N_36141,N_37065);
or U38001 (N_38001,N_36970,N_35024);
nor U38002 (N_38002,N_35949,N_35082);
nand U38003 (N_38003,N_37213,N_35479);
or U38004 (N_38004,N_35393,N_36161);
nor U38005 (N_38005,N_36051,N_35445);
and U38006 (N_38006,N_37359,N_37219);
and U38007 (N_38007,N_36043,N_36053);
nand U38008 (N_38008,N_36461,N_37370);
or U38009 (N_38009,N_36194,N_36076);
nor U38010 (N_38010,N_36190,N_35583);
nor U38011 (N_38011,N_36775,N_35647);
xor U38012 (N_38012,N_36742,N_36111);
and U38013 (N_38013,N_35915,N_37402);
or U38014 (N_38014,N_36125,N_36074);
nor U38015 (N_38015,N_36004,N_37045);
nand U38016 (N_38016,N_37369,N_35635);
or U38017 (N_38017,N_37046,N_36475);
nand U38018 (N_38018,N_35487,N_36090);
and U38019 (N_38019,N_36177,N_35163);
and U38020 (N_38020,N_35309,N_36476);
nand U38021 (N_38021,N_36760,N_35660);
or U38022 (N_38022,N_35303,N_36501);
or U38023 (N_38023,N_36830,N_36239);
nand U38024 (N_38024,N_35838,N_36002);
and U38025 (N_38025,N_36956,N_37428);
and U38026 (N_38026,N_36377,N_35977);
nor U38027 (N_38027,N_36782,N_36472);
and U38028 (N_38028,N_35498,N_37353);
nand U38029 (N_38029,N_35918,N_37028);
nor U38030 (N_38030,N_36191,N_35262);
and U38031 (N_38031,N_36652,N_37391);
or U38032 (N_38032,N_35985,N_36116);
and U38033 (N_38033,N_35829,N_37404);
xnor U38034 (N_38034,N_36480,N_36620);
xor U38035 (N_38035,N_36724,N_35104);
nor U38036 (N_38036,N_37180,N_36408);
nor U38037 (N_38037,N_36915,N_36918);
nor U38038 (N_38038,N_36671,N_36060);
and U38039 (N_38039,N_36883,N_37245);
nand U38040 (N_38040,N_36822,N_36624);
xnor U38041 (N_38041,N_35280,N_35336);
xor U38042 (N_38042,N_35767,N_35175);
or U38043 (N_38043,N_35200,N_36488);
or U38044 (N_38044,N_37157,N_37434);
nand U38045 (N_38045,N_36683,N_36858);
or U38046 (N_38046,N_35476,N_36467);
or U38047 (N_38047,N_36807,N_35391);
nor U38048 (N_38048,N_37037,N_35559);
or U38049 (N_38049,N_37155,N_37348);
and U38050 (N_38050,N_36715,N_37488);
and U38051 (N_38051,N_35683,N_36888);
nand U38052 (N_38052,N_35962,N_36381);
nand U38053 (N_38053,N_36082,N_37010);
and U38054 (N_38054,N_36189,N_36166);
and U38055 (N_38055,N_36806,N_37382);
and U38056 (N_38056,N_37498,N_36826);
or U38057 (N_38057,N_35798,N_37426);
nor U38058 (N_38058,N_36879,N_37274);
xnor U38059 (N_38059,N_36576,N_37438);
or U38060 (N_38060,N_37188,N_36600);
nor U38061 (N_38061,N_35216,N_35146);
nor U38062 (N_38062,N_37264,N_35911);
and U38063 (N_38063,N_35020,N_35366);
nand U38064 (N_38064,N_36042,N_35312);
or U38065 (N_38065,N_35067,N_36992);
and U38066 (N_38066,N_35328,N_36556);
xnor U38067 (N_38067,N_37463,N_36527);
and U38068 (N_38068,N_35847,N_35972);
xnor U38069 (N_38069,N_35133,N_36143);
nor U38070 (N_38070,N_37271,N_35247);
or U38071 (N_38071,N_37383,N_35245);
xor U38072 (N_38072,N_37323,N_35384);
and U38073 (N_38073,N_36818,N_36351);
xor U38074 (N_38074,N_35162,N_37448);
nor U38075 (N_38075,N_35026,N_37373);
nand U38076 (N_38076,N_35319,N_37276);
and U38077 (N_38077,N_35502,N_37243);
or U38078 (N_38078,N_36263,N_36978);
nand U38079 (N_38079,N_36502,N_36574);
nand U38080 (N_38080,N_35350,N_36212);
nor U38081 (N_38081,N_36006,N_37032);
nand U38082 (N_38082,N_36581,N_37303);
and U38083 (N_38083,N_35284,N_36543);
nand U38084 (N_38084,N_36312,N_36825);
xor U38085 (N_38085,N_35055,N_35785);
xnor U38086 (N_38086,N_35789,N_36168);
nor U38087 (N_38087,N_36063,N_35356);
nor U38088 (N_38088,N_36656,N_35049);
and U38089 (N_38089,N_35107,N_35516);
nand U38090 (N_38090,N_36982,N_35208);
xnor U38091 (N_38091,N_35538,N_35301);
xor U38092 (N_38092,N_36758,N_35485);
nor U38093 (N_38093,N_37443,N_36489);
nor U38094 (N_38094,N_36837,N_36820);
or U38095 (N_38095,N_35358,N_35531);
or U38096 (N_38096,N_36670,N_36638);
nor U38097 (N_38097,N_36391,N_35481);
xnor U38098 (N_38098,N_37172,N_37166);
nor U38099 (N_38099,N_36403,N_36584);
xor U38100 (N_38100,N_36286,N_37395);
and U38101 (N_38101,N_36854,N_35477);
xnor U38102 (N_38102,N_36416,N_35197);
xnor U38103 (N_38103,N_37057,N_36990);
and U38104 (N_38104,N_35189,N_36606);
nand U38105 (N_38105,N_35831,N_35993);
xnor U38106 (N_38106,N_36809,N_37012);
or U38107 (N_38107,N_37048,N_35513);
and U38108 (N_38108,N_35455,N_36386);
nand U38109 (N_38109,N_37256,N_36562);
nor U38110 (N_38110,N_36526,N_35786);
nor U38111 (N_38111,N_36784,N_36210);
nor U38112 (N_38112,N_35627,N_37118);
xor U38113 (N_38113,N_37220,N_36767);
nor U38114 (N_38114,N_35182,N_37278);
nand U38115 (N_38115,N_35921,N_36604);
nand U38116 (N_38116,N_35441,N_37158);
and U38117 (N_38117,N_35510,N_35097);
nor U38118 (N_38118,N_36425,N_35991);
xor U38119 (N_38119,N_36130,N_36222);
or U38120 (N_38120,N_35291,N_35396);
nor U38121 (N_38121,N_37401,N_36943);
nand U38122 (N_38122,N_36763,N_37400);
nor U38123 (N_38123,N_35822,N_37233);
nand U38124 (N_38124,N_35884,N_36282);
and U38125 (N_38125,N_37137,N_36005);
nor U38126 (N_38126,N_37160,N_35527);
nand U38127 (N_38127,N_36434,N_37067);
and U38128 (N_38128,N_36793,N_36070);
nand U38129 (N_38129,N_37301,N_35793);
nand U38130 (N_38130,N_37450,N_36443);
nor U38131 (N_38131,N_35451,N_36483);
nand U38132 (N_38132,N_37212,N_36205);
nor U38133 (N_38133,N_35975,N_35406);
nor U38134 (N_38134,N_35807,N_36813);
nor U38135 (N_38135,N_35631,N_35874);
and U38136 (N_38136,N_37072,N_36162);
nor U38137 (N_38137,N_35440,N_35272);
and U38138 (N_38138,N_37085,N_36393);
or U38139 (N_38139,N_37446,N_35268);
or U38140 (N_38140,N_36952,N_35383);
nand U38141 (N_38141,N_37141,N_36455);
or U38142 (N_38142,N_35525,N_35464);
nand U38143 (N_38143,N_36314,N_35413);
nand U38144 (N_38144,N_36474,N_36243);
or U38145 (N_38145,N_37462,N_35640);
xnor U38146 (N_38146,N_37145,N_35129);
xor U38147 (N_38147,N_36520,N_36555);
nor U38148 (N_38148,N_36342,N_36052);
xor U38149 (N_38149,N_35122,N_37038);
xnor U38150 (N_38150,N_36654,N_35058);
and U38151 (N_38151,N_36249,N_36667);
or U38152 (N_38152,N_36519,N_35254);
xnor U38153 (N_38153,N_35432,N_35278);
xnor U38154 (N_38154,N_37478,N_36493);
nand U38155 (N_38155,N_35499,N_36310);
xor U38156 (N_38156,N_36950,N_37135);
or U38157 (N_38157,N_35832,N_36534);
nor U38158 (N_38158,N_35604,N_36364);
nor U38159 (N_38159,N_35673,N_36482);
nor U38160 (N_38160,N_35539,N_36073);
nand U38161 (N_38161,N_36592,N_36688);
nor U38162 (N_38162,N_36679,N_37052);
nor U38163 (N_38163,N_35148,N_35934);
and U38164 (N_38164,N_35651,N_35313);
xnor U38165 (N_38165,N_36927,N_35731);
and U38166 (N_38166,N_35497,N_36794);
nor U38167 (N_38167,N_36086,N_35966);
or U38168 (N_38168,N_37258,N_37230);
xnor U38169 (N_38169,N_35682,N_37409);
and U38170 (N_38170,N_35467,N_36930);
nand U38171 (N_38171,N_35873,N_37140);
nor U38172 (N_38172,N_36422,N_37377);
and U38173 (N_38173,N_36985,N_36254);
nor U38174 (N_38174,N_36932,N_36725);
and U38175 (N_38175,N_36406,N_35566);
or U38176 (N_38176,N_36367,N_35795);
nand U38177 (N_38177,N_36568,N_35741);
or U38178 (N_38178,N_36012,N_36561);
xnor U38179 (N_38179,N_35236,N_35678);
and U38180 (N_38180,N_36407,N_35283);
xnor U38181 (N_38181,N_36523,N_36268);
nand U38182 (N_38182,N_36458,N_36349);
or U38183 (N_38183,N_37083,N_35726);
and U38184 (N_38184,N_37176,N_35100);
nand U38185 (N_38185,N_36933,N_35529);
nand U38186 (N_38186,N_36736,N_35923);
and U38187 (N_38187,N_37453,N_35687);
nor U38188 (N_38188,N_35337,N_35722);
xor U38189 (N_38189,N_36400,N_37021);
xor U38190 (N_38190,N_36253,N_35447);
xor U38191 (N_38191,N_35388,N_35266);
or U38192 (N_38192,N_36571,N_37112);
xor U38193 (N_38193,N_36450,N_37241);
xnor U38194 (N_38194,N_35124,N_36170);
nor U38195 (N_38195,N_35362,N_35826);
or U38196 (N_38196,N_37318,N_37020);
or U38197 (N_38197,N_37124,N_36959);
or U38198 (N_38198,N_37418,N_35765);
or U38199 (N_38199,N_36127,N_35954);
and U38200 (N_38200,N_35757,N_35088);
xor U38201 (N_38201,N_37226,N_35508);
and U38202 (N_38202,N_35746,N_36272);
xor U38203 (N_38203,N_36321,N_35814);
nor U38204 (N_38204,N_37116,N_35990);
or U38205 (N_38205,N_36394,N_36047);
xor U38206 (N_38206,N_35790,N_35775);
nand U38207 (N_38207,N_36972,N_36998);
nand U38208 (N_38208,N_35230,N_36080);
nor U38209 (N_38209,N_37447,N_35809);
or U38210 (N_38210,N_35668,N_35855);
and U38211 (N_38211,N_37081,N_35376);
nand U38212 (N_38212,N_36567,N_36050);
and U38213 (N_38213,N_35941,N_35959);
xor U38214 (N_38214,N_35664,N_36007);
nand U38215 (N_38215,N_36810,N_35880);
xnor U38216 (N_38216,N_36150,N_36842);
and U38217 (N_38217,N_36172,N_36735);
nand U38218 (N_38218,N_35718,N_35643);
nor U38219 (N_38219,N_35382,N_36155);
nor U38220 (N_38220,N_37024,N_35721);
xnor U38221 (N_38221,N_36297,N_37251);
xnor U38222 (N_38222,N_36149,N_36444);
and U38223 (N_38223,N_36440,N_37214);
nor U38224 (N_38224,N_35842,N_36059);
xnor U38225 (N_38225,N_35299,N_35610);
and U38226 (N_38226,N_36347,N_36368);
xnor U38227 (N_38227,N_37070,N_35377);
nand U38228 (N_38228,N_36769,N_36266);
nand U38229 (N_38229,N_36602,N_36040);
nor U38230 (N_38230,N_36237,N_37078);
or U38231 (N_38231,N_37239,N_36156);
or U38232 (N_38232,N_37484,N_35285);
or U38233 (N_38233,N_36468,N_36726);
nor U38234 (N_38234,N_36504,N_35602);
or U38235 (N_38235,N_35904,N_37040);
nand U38236 (N_38236,N_35489,N_36441);
nand U38237 (N_38237,N_37321,N_35169);
xnor U38238 (N_38238,N_35614,N_35210);
or U38239 (N_38239,N_37249,N_36546);
nand U38240 (N_38240,N_36157,N_36514);
nand U38241 (N_38241,N_35465,N_35729);
nor U38242 (N_38242,N_37033,N_36307);
or U38243 (N_38243,N_36741,N_35106);
nand U38244 (N_38244,N_36965,N_36538);
and U38245 (N_38245,N_35298,N_35976);
nand U38246 (N_38246,N_37182,N_35186);
or U38247 (N_38247,N_37122,N_36632);
nor U38248 (N_38248,N_36870,N_36019);
xnor U38249 (N_38249,N_35629,N_35143);
nand U38250 (N_38250,N_36553,N_37261);
or U38251 (N_38251,N_35019,N_36336);
and U38252 (N_38252,N_36675,N_35979);
or U38253 (N_38253,N_37029,N_36484);
or U38254 (N_38254,N_36682,N_36255);
or U38255 (N_38255,N_37315,N_37464);
and U38256 (N_38256,N_37164,N_35859);
nand U38257 (N_38257,N_36011,N_36404);
and U38258 (N_38258,N_35433,N_37273);
or U38259 (N_38259,N_36791,N_35546);
nor U38260 (N_38260,N_37327,N_36245);
nand U38261 (N_38261,N_36034,N_35517);
xnor U38262 (N_38262,N_36319,N_37190);
xnor U38263 (N_38263,N_36900,N_37471);
nand U38264 (N_38264,N_37139,N_35410);
nor U38265 (N_38265,N_37022,N_36481);
nand U38266 (N_38266,N_35035,N_36921);
nor U38267 (N_38267,N_35907,N_35582);
or U38268 (N_38268,N_35556,N_35094);
nand U38269 (N_38269,N_35557,N_35999);
and U38270 (N_38270,N_35938,N_36102);
nand U38271 (N_38271,N_37444,N_36120);
and U38272 (N_38272,N_36680,N_36540);
xnor U38273 (N_38273,N_35386,N_35845);
and U38274 (N_38274,N_35576,N_35409);
nand U38275 (N_38275,N_36891,N_36124);
nor U38276 (N_38276,N_35119,N_36578);
nor U38277 (N_38277,N_36904,N_35567);
nand U38278 (N_38278,N_37255,N_36765);
nand U38279 (N_38279,N_37227,N_36623);
xnor U38280 (N_38280,N_35836,N_36129);
nor U38281 (N_38281,N_35142,N_35547);
or U38282 (N_38282,N_36664,N_35238);
and U38283 (N_38283,N_36657,N_35102);
nor U38284 (N_38284,N_36343,N_36083);
or U38285 (N_38285,N_35909,N_37184);
and U38286 (N_38286,N_35596,N_36819);
and U38287 (N_38287,N_35840,N_35132);
or U38288 (N_38288,N_36774,N_35079);
or U38289 (N_38289,N_36707,N_37095);
and U38290 (N_38290,N_35503,N_35253);
and U38291 (N_38291,N_35308,N_35357);
and U38292 (N_38292,N_36803,N_37465);
nor U38293 (N_38293,N_35125,N_36417);
and U38294 (N_38294,N_37202,N_35905);
nor U38295 (N_38295,N_36066,N_37451);
nand U38296 (N_38296,N_36292,N_36433);
or U38297 (N_38297,N_36529,N_36607);
xor U38298 (N_38298,N_35233,N_35010);
xnor U38299 (N_38299,N_37489,N_35226);
nand U38300 (N_38300,N_36224,N_35461);
nand U38301 (N_38301,N_37076,N_35195);
nand U38302 (N_38302,N_35965,N_36693);
nand U38303 (N_38303,N_35205,N_36703);
xor U38304 (N_38304,N_36446,N_36752);
xor U38305 (N_38305,N_37486,N_36387);
or U38306 (N_38306,N_36864,N_36609);
nand U38307 (N_38307,N_35179,N_37393);
xnor U38308 (N_38308,N_37193,N_36890);
nand U38309 (N_38309,N_35389,N_35897);
or U38310 (N_38310,N_36821,N_37144);
nand U38311 (N_38311,N_35974,N_36285);
xor U38312 (N_38312,N_36359,N_35037);
xnor U38313 (N_38313,N_35639,N_36283);
or U38314 (N_38314,N_35059,N_36180);
and U38315 (N_38315,N_35914,N_36208);
xnor U38316 (N_38316,N_35560,N_35821);
or U38317 (N_38317,N_35691,N_36431);
or U38318 (N_38318,N_35370,N_35803);
xnor U38319 (N_38319,N_37246,N_36994);
nor U38320 (N_38320,N_36989,N_36426);
or U38321 (N_38321,N_36366,N_35417);
nand U38322 (N_38322,N_36812,N_35970);
and U38323 (N_38323,N_36315,N_37403);
and U38324 (N_38324,N_35745,N_35747);
xor U38325 (N_38325,N_36549,N_36678);
xnor U38326 (N_38326,N_35657,N_35178);
xnor U38327 (N_38327,N_35255,N_36757);
nand U38328 (N_38328,N_36300,N_36711);
xnor U38329 (N_38329,N_37002,N_35670);
nand U38330 (N_38330,N_35994,N_37073);
and U38331 (N_38331,N_36633,N_37302);
xnor U38332 (N_38332,N_36003,N_35782);
or U38333 (N_38333,N_35378,N_37282);
xor U38334 (N_38334,N_37044,N_35111);
nor U38335 (N_38335,N_35416,N_35690);
or U38336 (N_38336,N_37165,N_36252);
nand U38337 (N_38337,N_35512,N_36020);
nor U38338 (N_38338,N_35828,N_36748);
nand U38339 (N_38339,N_37316,N_35712);
and U38340 (N_38340,N_37476,N_35612);
xnor U38341 (N_38341,N_37483,N_37385);
nand U38342 (N_38342,N_35109,N_36507);
and U38343 (N_38343,N_35592,N_36732);
nand U38344 (N_38344,N_37493,N_36187);
nor U38345 (N_38345,N_36498,N_36234);
xor U38346 (N_38346,N_37441,N_36383);
or U38347 (N_38347,N_36542,N_36651);
xnor U38348 (N_38348,N_35398,N_36878);
or U38349 (N_38349,N_35805,N_37380);
and U38350 (N_38350,N_35530,N_35004);
and U38351 (N_38351,N_36637,N_36153);
xnor U38352 (N_38352,N_36478,N_35463);
and U38353 (N_38353,N_36797,N_36702);
xnor U38354 (N_38354,N_35533,N_36697);
or U38355 (N_38355,N_35761,N_37008);
nand U38356 (N_38356,N_36142,N_35343);
nand U38357 (N_38357,N_36325,N_36677);
and U38358 (N_38358,N_36800,N_36088);
xor U38359 (N_38359,N_35581,N_37469);
nand U38360 (N_38360,N_37363,N_35127);
and U38361 (N_38361,N_37018,N_36611);
xor U38362 (N_38362,N_37286,N_37336);
xor U38363 (N_38363,N_36058,N_35589);
or U38364 (N_38364,N_35071,N_35450);
and U38365 (N_38365,N_35638,N_36723);
nor U38366 (N_38366,N_36585,N_35549);
nor U38367 (N_38367,N_36861,N_36944);
nand U38368 (N_38368,N_37069,N_35953);
nand U38369 (N_38369,N_35997,N_35947);
nor U38370 (N_38370,N_36015,N_35986);
and U38371 (N_38371,N_36722,N_36411);
or U38372 (N_38372,N_36077,N_36969);
and U38373 (N_38373,N_35585,N_35992);
nand U38374 (N_38374,N_35936,N_35081);
and U38375 (N_38375,N_36410,N_36739);
nand U38376 (N_38376,N_36564,N_36635);
nand U38377 (N_38377,N_37329,N_35098);
nand U38378 (N_38378,N_35022,N_36719);
nand U38379 (N_38379,N_37064,N_35925);
nand U38380 (N_38380,N_37368,N_36582);
xor U38381 (N_38381,N_36376,N_37051);
nor U38382 (N_38382,N_37341,N_36756);
xnor U38383 (N_38383,N_37357,N_35408);
and U38384 (N_38384,N_35967,N_36889);
xnor U38385 (N_38385,N_35764,N_37297);
and U38386 (N_38386,N_36559,N_37272);
nand U38387 (N_38387,N_37242,N_36329);
nor U38388 (N_38388,N_35310,N_36539);
nor U38389 (N_38389,N_36165,N_36563);
xnor U38390 (N_38390,N_35799,N_36762);
nand U38391 (N_38391,N_37186,N_35839);
nand U38392 (N_38392,N_35322,N_36460);
or U38393 (N_38393,N_35820,N_36075);
or U38394 (N_38394,N_35187,N_37479);
nand U38395 (N_38395,N_36541,N_35662);
nor U38396 (N_38396,N_36197,N_37308);
and U38397 (N_38397,N_36128,N_35212);
or U38398 (N_38398,N_36845,N_35630);
nor U38399 (N_38399,N_36418,N_37154);
xor U38400 (N_38400,N_36550,N_37371);
nor U38401 (N_38401,N_35379,N_37440);
xnor U38402 (N_38402,N_36069,N_36109);
nor U38403 (N_38403,N_35919,N_35128);
nand U38404 (N_38404,N_37086,N_35039);
nand U38405 (N_38405,N_35292,N_36873);
nor U38406 (N_38406,N_35575,N_36827);
nand U38407 (N_38407,N_36144,N_37091);
nor U38408 (N_38408,N_35951,N_37201);
nor U38409 (N_38409,N_36749,N_36279);
xor U38410 (N_38410,N_36054,N_37267);
and U38411 (N_38411,N_35491,N_36293);
and U38412 (N_38412,N_37312,N_36689);
nor U38413 (N_38413,N_35815,N_36046);
or U38414 (N_38414,N_36346,N_35087);
and U38415 (N_38415,N_36588,N_37350);
nor U38416 (N_38416,N_36805,N_35860);
nand U38417 (N_38417,N_37366,N_37110);
or U38418 (N_38418,N_36389,N_36687);
or U38419 (N_38419,N_36031,N_35658);
or U38420 (N_38420,N_36860,N_35804);
or U38421 (N_38421,N_37405,N_37178);
nor U38422 (N_38422,N_36641,N_37474);
and U38423 (N_38423,N_36846,N_36867);
xor U38424 (N_38424,N_35882,N_35257);
nand U38425 (N_38425,N_35338,N_35620);
nor U38426 (N_38426,N_36557,N_36217);
nand U38427 (N_38427,N_36738,N_35223);
or U38428 (N_38428,N_35484,N_35565);
xor U38429 (N_38429,N_35054,N_36898);
xor U38430 (N_38430,N_35616,N_35121);
xor U38431 (N_38431,N_36558,N_35564);
nand U38432 (N_38432,N_35945,N_35348);
xnor U38433 (N_38433,N_37039,N_35219);
and U38434 (N_38434,N_36133,N_36309);
and U38435 (N_38435,N_35878,N_35333);
nand U38436 (N_38436,N_35015,N_36244);
nor U38437 (N_38437,N_36790,N_37433);
and U38438 (N_38438,N_36490,N_36095);
nand U38439 (N_38439,N_36597,N_35857);
xnor U38440 (N_38440,N_37417,N_37466);
or U38441 (N_38441,N_36601,N_35550);
xor U38442 (N_38442,N_35562,N_35617);
xnor U38443 (N_38443,N_37229,N_36877);
xor U38444 (N_38444,N_35674,N_36917);
xnor U38445 (N_38445,N_37244,N_37231);
and U38446 (N_38446,N_36432,N_37290);
and U38447 (N_38447,N_35621,N_36365);
nor U38448 (N_38448,N_35166,N_36271);
xnor U38449 (N_38449,N_35597,N_35908);
nor U38450 (N_38450,N_37414,N_37492);
nor U38451 (N_38451,N_36685,N_37281);
or U38452 (N_38452,N_35114,N_35933);
and U38453 (N_38453,N_37305,N_35810);
nand U38454 (N_38454,N_37472,N_35780);
and U38455 (N_38455,N_37364,N_35588);
or U38456 (N_38456,N_36209,N_37047);
nand U38457 (N_38457,N_35740,N_36207);
or U38458 (N_38458,N_37259,N_37283);
or U38459 (N_38459,N_37294,N_35198);
xor U38460 (N_38460,N_37109,N_37247);
nor U38461 (N_38461,N_36788,N_35846);
xor U38462 (N_38462,N_35998,N_35561);
and U38463 (N_38463,N_36065,N_35875);
or U38464 (N_38464,N_35397,N_35335);
nand U38465 (N_38465,N_37089,N_36886);
or U38466 (N_38466,N_37415,N_37295);
and U38467 (N_38467,N_36920,N_36306);
xor U38468 (N_38468,N_37128,N_35578);
or U38469 (N_38469,N_36338,N_35134);
xnor U38470 (N_38470,N_36953,N_35323);
or U38471 (N_38471,N_37134,N_36195);
or U38472 (N_38472,N_36041,N_35141);
and U38473 (N_38473,N_36385,N_35650);
xnor U38474 (N_38474,N_35387,N_36655);
nor U38475 (N_38475,N_35636,N_36997);
or U38476 (N_38476,N_35120,N_36372);
nor U38477 (N_38477,N_36497,N_35239);
nand U38478 (N_38478,N_35694,N_35064);
nor U38479 (N_38479,N_37467,N_35372);
or U38480 (N_38480,N_36761,N_36866);
nor U38481 (N_38481,N_37031,N_36148);
and U38482 (N_38482,N_36219,N_37322);
nor U38483 (N_38483,N_36552,N_36986);
or U38484 (N_38484,N_37099,N_35115);
or U38485 (N_38485,N_35191,N_35774);
nand U38486 (N_38486,N_35762,N_36565);
or U38487 (N_38487,N_35399,N_35573);
nand U38488 (N_38488,N_35240,N_35355);
nand U38489 (N_38489,N_37346,N_37136);
and U38490 (N_38490,N_36977,N_37268);
nand U38491 (N_38491,N_36451,N_36045);
or U38492 (N_38492,N_35862,N_37482);
or U38493 (N_38493,N_37497,N_35131);
xor U38494 (N_38494,N_36573,N_36745);
xnor U38495 (N_38495,N_37181,N_35698);
nor U38496 (N_38496,N_37408,N_36113);
nand U38497 (N_38497,N_36834,N_36744);
nand U38498 (N_38498,N_36135,N_35889);
and U38499 (N_38499,N_36089,N_35264);
xor U38500 (N_38500,N_36975,N_35469);
nor U38501 (N_38501,N_35926,N_35235);
nor U38502 (N_38502,N_37121,N_37207);
nand U38503 (N_38503,N_35220,N_35103);
and U38504 (N_38504,N_37287,N_36136);
nor U38505 (N_38505,N_35021,N_36768);
and U38506 (N_38506,N_36857,N_36399);
and U38507 (N_38507,N_36801,N_36892);
or U38508 (N_38508,N_35038,N_35225);
and U38509 (N_38509,N_35311,N_35294);
or U38510 (N_38510,N_36779,N_35978);
and U38511 (N_38511,N_36874,N_36811);
nor U38512 (N_38512,N_37487,N_36235);
or U38513 (N_38513,N_35093,N_37152);
nor U38514 (N_38514,N_36751,N_35438);
and U38515 (N_38515,N_36049,N_36265);
xnor U38516 (N_38516,N_36923,N_35665);
or U38517 (N_38517,N_36193,N_37427);
nor U38518 (N_38518,N_35402,N_35199);
or U38519 (N_38519,N_35154,N_36551);
xor U38520 (N_38520,N_37017,N_37360);
xor U38521 (N_38521,N_35483,N_35540);
xnor U38522 (N_38522,N_36078,N_37113);
nand U38523 (N_38523,N_35984,N_35952);
xnor U38524 (N_38524,N_37296,N_36215);
and U38525 (N_38525,N_36669,N_37253);
xnor U38526 (N_38526,N_35354,N_36241);
and U38527 (N_38527,N_36016,N_36000);
nor U38528 (N_38528,N_35096,N_35848);
nand U38529 (N_38529,N_37161,N_35209);
nand U38530 (N_38530,N_36442,N_35830);
nand U38531 (N_38531,N_36485,N_36798);
or U38532 (N_38532,N_37001,N_37473);
xnor U38533 (N_38533,N_36232,N_36964);
or U38534 (N_38534,N_35768,N_36331);
or U38535 (N_38535,N_36027,N_35969);
nor U38536 (N_38536,N_37077,N_36104);
nand U38537 (N_38537,N_37129,N_35101);
or U38538 (N_38538,N_35843,N_36057);
or U38539 (N_38539,N_35720,N_36010);
xnor U38540 (N_38540,N_36178,N_35725);
nand U38541 (N_38541,N_37146,N_37422);
and U38542 (N_38542,N_35942,N_36320);
or U38543 (N_38543,N_36636,N_35318);
nor U38544 (N_38544,N_35273,N_36859);
nor U38545 (N_38545,N_35928,N_35092);
nor U38546 (N_38546,N_37419,N_35073);
and U38547 (N_38547,N_37356,N_35105);
xnor U38548 (N_38548,N_35008,N_35877);
xor U38549 (N_38549,N_35519,N_35259);
nand U38550 (N_38550,N_36612,N_35709);
and U38551 (N_38551,N_35901,N_37171);
nor U38552 (N_38552,N_36029,N_35669);
and U38553 (N_38553,N_36598,N_35066);
nor U38554 (N_38554,N_35943,N_36572);
nand U38555 (N_38555,N_36392,N_36856);
or U38556 (N_38556,N_35871,N_35072);
or U38557 (N_38557,N_35032,N_35089);
nor U38558 (N_38558,N_36096,N_35584);
nand U38559 (N_38559,N_35192,N_35188);
and U38560 (N_38560,N_36925,N_36658);
nor U38561 (N_38561,N_36668,N_36705);
or U38562 (N_38562,N_37269,N_36533);
nor U38563 (N_38563,N_36695,N_35518);
nor U38564 (N_38564,N_36428,N_36681);
nor U38565 (N_38565,N_35534,N_36599);
nand U38566 (N_38566,N_36463,N_35930);
and U38567 (N_38567,N_37361,N_36327);
nand U38568 (N_38568,N_37392,N_35194);
xor U38569 (N_38569,N_37421,N_35776);
nand U38570 (N_38570,N_35265,N_35359);
xor U38571 (N_38571,N_36420,N_36139);
xor U38572 (N_38572,N_36246,N_36912);
nor U38573 (N_38573,N_35159,N_36823);
or U38574 (N_38574,N_36179,N_36084);
nor U38575 (N_38575,N_36269,N_36808);
and U38576 (N_38576,N_36525,N_35428);
and U38577 (N_38577,N_36236,N_37455);
nor U38578 (N_38578,N_35274,N_36851);
nor U38579 (N_38579,N_36999,N_35075);
or U38580 (N_38580,N_37035,N_35395);
and U38581 (N_38581,N_36909,N_35045);
or U38582 (N_38582,N_35579,N_37025);
and U38583 (N_38583,N_35571,N_37036);
and U38584 (N_38584,N_35364,N_37355);
and U38585 (N_38585,N_35543,N_36709);
and U38586 (N_38586,N_37423,N_37335);
xnor U38587 (N_38587,N_35403,N_36413);
nand U38588 (N_38588,N_35917,N_35728);
xnor U38589 (N_38589,N_35980,N_35856);
nand U38590 (N_38590,N_36532,N_35243);
nand U38591 (N_38591,N_36863,N_35448);
and U38592 (N_38592,N_35368,N_35625);
nand U38593 (N_38593,N_36037,N_36629);
nor U38594 (N_38594,N_35047,N_35754);
nand U38595 (N_38595,N_37203,N_35661);
or U38596 (N_38596,N_35797,N_37063);
nand U38597 (N_38597,N_36270,N_37300);
and U38598 (N_38598,N_35161,N_35895);
xor U38599 (N_38599,N_36021,N_37310);
nand U38600 (N_38600,N_36114,N_35825);
nand U38601 (N_38601,N_36477,N_36119);
xor U38602 (N_38602,N_37445,N_36720);
nand U38603 (N_38603,N_37200,N_35052);
xnor U38604 (N_38604,N_37054,N_35258);
and U38605 (N_38605,N_36661,N_35773);
or U38606 (N_38606,N_36214,N_36899);
or U38607 (N_38607,N_37389,N_37127);
or U38608 (N_38608,N_36908,N_36322);
nand U38609 (N_38609,N_37328,N_35033);
nand U38610 (N_38610,N_35894,N_37026);
nor U38611 (N_38611,N_36579,N_35495);
nor U38612 (N_38612,N_35568,N_36487);
and U38613 (N_38613,N_36348,N_37470);
or U38614 (N_38614,N_37339,N_37333);
or U38615 (N_38615,N_35989,N_36968);
nor U38616 (N_38616,N_37459,N_35648);
nand U38617 (N_38617,N_36032,N_36802);
xor U38618 (N_38618,N_37307,N_35150);
and U38619 (N_38619,N_35256,N_36435);
or U38620 (N_38620,N_36979,N_35542);
or U38621 (N_38621,N_36184,N_35077);
nand U38622 (N_38622,N_37325,N_35496);
nor U38623 (N_38623,N_36545,N_35480);
or U38624 (N_38624,N_37050,N_36014);
xor U38625 (N_38625,N_35036,N_37384);
xnor U38626 (N_38626,N_37314,N_35891);
and U38627 (N_38627,N_37457,N_36515);
or U38628 (N_38628,N_36103,N_36495);
nor U38629 (N_38629,N_35572,N_36804);
or U38630 (N_38630,N_35916,N_37430);
nor U38631 (N_38631,N_35555,N_36171);
xor U38632 (N_38632,N_37208,N_37386);
and U38633 (N_38633,N_35501,N_36831);
and U38634 (N_38634,N_35196,N_35717);
and U38635 (N_38635,N_36423,N_35792);
xnor U38636 (N_38636,N_36608,N_35227);
xnor U38637 (N_38637,N_36100,N_35068);
xor U38638 (N_38638,N_36151,N_36848);
xor U38639 (N_38639,N_36855,N_36634);
nand U38640 (N_38640,N_37431,N_36973);
or U38641 (N_38641,N_36098,N_36221);
or U38642 (N_38642,N_37169,N_37413);
and U38643 (N_38643,N_36824,N_35619);
and U38644 (N_38644,N_36983,N_36277);
xnor U38645 (N_38645,N_36122,N_35766);
and U38646 (N_38646,N_35750,N_37358);
nand U38647 (N_38647,N_35269,N_35449);
nand U38648 (N_38648,N_37257,N_36371);
nand U38649 (N_38649,N_36091,N_35471);
nor U38650 (N_38650,N_36081,N_36354);
nor U38651 (N_38651,N_35468,N_35193);
nand U38652 (N_38652,N_36708,N_35920);
or U38653 (N_38653,N_36154,N_35062);
and U38654 (N_38654,N_36350,N_35813);
nor U38655 (N_38655,N_37177,N_35666);
or U38656 (N_38656,N_36145,N_36456);
nor U38657 (N_38657,N_35736,N_36747);
and U38658 (N_38658,N_35123,N_35365);
xor U38659 (N_38659,N_36876,N_37435);
xnor U38660 (N_38660,N_37280,N_37211);
and U38661 (N_38661,N_36412,N_35689);
or U38662 (N_38662,N_35667,N_36614);
and U38663 (N_38663,N_37221,N_35005);
nor U38664 (N_38664,N_37319,N_35680);
or U38665 (N_38665,N_36353,N_35206);
nor U38666 (N_38666,N_36362,N_35868);
xor U38667 (N_38667,N_35422,N_37442);
nand U38668 (N_38668,N_36770,N_35659);
or U38669 (N_38669,N_37142,N_35074);
xor U38670 (N_38670,N_36267,N_36642);
or U38671 (N_38671,N_35286,N_35900);
nor U38672 (N_38672,N_35796,N_35136);
nor U38673 (N_38673,N_35177,N_37191);
xor U38674 (N_38674,N_37162,N_37279);
xnor U38675 (N_38675,N_36627,N_35794);
nor U38676 (N_38676,N_35405,N_35599);
nand U38677 (N_38677,N_35971,N_37387);
nand U38678 (N_38678,N_36390,N_36844);
nor U38679 (N_38679,N_35470,N_35315);
and U38680 (N_38680,N_37266,N_35267);
nor U38681 (N_38681,N_36875,N_35013);
and U38682 (N_38682,N_37009,N_36402);
or U38683 (N_38683,N_35570,N_35705);
and U38684 (N_38684,N_36626,N_35475);
nand U38685 (N_38685,N_36631,N_35443);
and U38686 (N_38686,N_35056,N_35624);
and U38687 (N_38687,N_36340,N_36374);
nor U38688 (N_38688,N_36914,N_35854);
nand U38689 (N_38689,N_37103,N_36963);
nand U38690 (N_38690,N_37060,N_37082);
nor U38691 (N_38691,N_36617,N_37379);
nand U38692 (N_38692,N_36621,N_36938);
nand U38693 (N_38693,N_36174,N_35535);
nor U38694 (N_38694,N_35879,N_36714);
or U38695 (N_38695,N_36360,N_35003);
or U38696 (N_38696,N_36036,N_36225);
nand U38697 (N_38697,N_35224,N_36583);
or U38698 (N_38698,N_35606,N_35618);
or U38699 (N_38699,N_36759,N_36427);
and U38700 (N_38700,N_35748,N_37460);
or U38701 (N_38701,N_36085,N_35946);
and U38702 (N_38702,N_36486,N_35027);
xor U38703 (N_38703,N_36901,N_36301);
nor U38704 (N_38704,N_36916,N_35872);
or U38705 (N_38705,N_35601,N_35956);
or U38706 (N_38706,N_35787,N_35899);
nor U38707 (N_38707,N_36175,N_36941);
and U38708 (N_38708,N_35652,N_37224);
or U38709 (N_38709,N_35207,N_35139);
nor U38710 (N_38710,N_35913,N_36829);
and U38711 (N_38711,N_36518,N_35522);
xnor U38712 (N_38712,N_36028,N_35671);
xor U38713 (N_38713,N_37390,N_36072);
nor U38714 (N_38714,N_35811,N_36605);
xnor U38715 (N_38715,N_35515,N_37412);
and U38716 (N_38716,N_35655,N_35353);
or U38717 (N_38717,N_35528,N_35885);
xor U38718 (N_38718,N_35684,N_35753);
xor U38719 (N_38719,N_36991,N_37420);
xor U38720 (N_38720,N_36596,N_35043);
xor U38721 (N_38721,N_36887,N_35598);
or U38722 (N_38722,N_35672,N_37007);
xor U38723 (N_38723,N_35204,N_35012);
or U38724 (N_38724,N_37317,N_36415);
or U38725 (N_38725,N_35505,N_36881);
nor U38726 (N_38726,N_35865,N_35603);
or U38727 (N_38727,N_36013,N_36231);
nand U38728 (N_38728,N_36566,N_37119);
and U38729 (N_38729,N_36796,N_37235);
nor U38730 (N_38730,N_36378,N_37003);
xor U38731 (N_38731,N_37147,N_35157);
nand U38732 (N_38732,N_35922,N_37424);
or U38733 (N_38733,N_36731,N_35890);
and U38734 (N_38734,N_35095,N_36369);
xor U38735 (N_38735,N_36206,N_36356);
or U38736 (N_38736,N_37265,N_36164);
or U38737 (N_38737,N_35076,N_35152);
xnor U38738 (N_38738,N_36698,N_37432);
nor U38739 (N_38739,N_36470,N_35302);
nand U38740 (N_38740,N_36038,N_36409);
xnor U38741 (N_38741,N_36560,N_35869);
and U38742 (N_38742,N_35112,N_36884);
and U38743 (N_38743,N_35749,N_35802);
and U38744 (N_38744,N_35078,N_35234);
and U38745 (N_38745,N_37056,N_37066);
nor U38746 (N_38746,N_35646,N_36814);
or U38747 (N_38747,N_35819,N_35692);
or U38748 (N_38748,N_37173,N_35340);
or U38749 (N_38749,N_35261,N_35213);
and U38750 (N_38750,N_35302,N_35318);
xnor U38751 (N_38751,N_36716,N_37305);
and U38752 (N_38752,N_36024,N_35918);
nand U38753 (N_38753,N_35178,N_37299);
and U38754 (N_38754,N_36551,N_35936);
and U38755 (N_38755,N_35056,N_36505);
nor U38756 (N_38756,N_35375,N_35088);
nand U38757 (N_38757,N_37079,N_35604);
nor U38758 (N_38758,N_35513,N_35908);
nor U38759 (N_38759,N_36872,N_35022);
and U38760 (N_38760,N_36056,N_37075);
xor U38761 (N_38761,N_36829,N_35444);
nand U38762 (N_38762,N_35056,N_36921);
xnor U38763 (N_38763,N_36319,N_36028);
and U38764 (N_38764,N_37190,N_35262);
or U38765 (N_38765,N_35005,N_37230);
or U38766 (N_38766,N_35763,N_36909);
and U38767 (N_38767,N_37231,N_35606);
or U38768 (N_38768,N_35746,N_36069);
nand U38769 (N_38769,N_35086,N_35903);
nor U38770 (N_38770,N_36820,N_37184);
and U38771 (N_38771,N_37263,N_35115);
nand U38772 (N_38772,N_37250,N_37245);
xnor U38773 (N_38773,N_36087,N_35373);
nand U38774 (N_38774,N_36501,N_35581);
nor U38775 (N_38775,N_35775,N_35628);
nor U38776 (N_38776,N_37301,N_36911);
and U38777 (N_38777,N_35212,N_35369);
nor U38778 (N_38778,N_35699,N_36375);
nand U38779 (N_38779,N_35111,N_35425);
xnor U38780 (N_38780,N_35379,N_37490);
nand U38781 (N_38781,N_37244,N_35743);
nor U38782 (N_38782,N_35589,N_35318);
or U38783 (N_38783,N_35514,N_36578);
and U38784 (N_38784,N_35540,N_36739);
xnor U38785 (N_38785,N_35165,N_36055);
and U38786 (N_38786,N_37293,N_36708);
nand U38787 (N_38787,N_37134,N_37208);
or U38788 (N_38788,N_36363,N_36732);
xnor U38789 (N_38789,N_35023,N_36045);
and U38790 (N_38790,N_35518,N_37302);
nor U38791 (N_38791,N_35346,N_35867);
xor U38792 (N_38792,N_36322,N_35716);
nor U38793 (N_38793,N_36657,N_35148);
or U38794 (N_38794,N_35441,N_37301);
and U38795 (N_38795,N_36645,N_37173);
or U38796 (N_38796,N_36634,N_35511);
xnor U38797 (N_38797,N_37317,N_37022);
nand U38798 (N_38798,N_37079,N_35370);
nor U38799 (N_38799,N_36899,N_36430);
or U38800 (N_38800,N_35657,N_36605);
xor U38801 (N_38801,N_36505,N_35591);
nor U38802 (N_38802,N_35058,N_36635);
xor U38803 (N_38803,N_36010,N_36082);
nor U38804 (N_38804,N_36096,N_37301);
nand U38805 (N_38805,N_37060,N_36462);
nand U38806 (N_38806,N_36583,N_35173);
nor U38807 (N_38807,N_35287,N_35351);
xnor U38808 (N_38808,N_36693,N_35432);
or U38809 (N_38809,N_35117,N_35990);
nand U38810 (N_38810,N_35798,N_36102);
nor U38811 (N_38811,N_36424,N_37350);
nor U38812 (N_38812,N_35235,N_36255);
xor U38813 (N_38813,N_37108,N_36005);
xor U38814 (N_38814,N_36040,N_35782);
xor U38815 (N_38815,N_37038,N_36559);
and U38816 (N_38816,N_35406,N_35792);
and U38817 (N_38817,N_35105,N_35138);
and U38818 (N_38818,N_36957,N_35107);
or U38819 (N_38819,N_36052,N_36633);
and U38820 (N_38820,N_36921,N_35127);
and U38821 (N_38821,N_36455,N_37333);
nand U38822 (N_38822,N_35453,N_35849);
and U38823 (N_38823,N_35002,N_35100);
or U38824 (N_38824,N_36803,N_36830);
nor U38825 (N_38825,N_37499,N_35918);
nand U38826 (N_38826,N_36653,N_36105);
xor U38827 (N_38827,N_37473,N_35227);
nand U38828 (N_38828,N_35635,N_35443);
or U38829 (N_38829,N_37383,N_37043);
and U38830 (N_38830,N_36313,N_37341);
or U38831 (N_38831,N_36179,N_36982);
nand U38832 (N_38832,N_36722,N_36390);
or U38833 (N_38833,N_36145,N_36362);
or U38834 (N_38834,N_36638,N_36217);
and U38835 (N_38835,N_35828,N_35765);
nand U38836 (N_38836,N_37024,N_36708);
or U38837 (N_38837,N_36243,N_36952);
xor U38838 (N_38838,N_36244,N_35301);
nor U38839 (N_38839,N_35705,N_35630);
and U38840 (N_38840,N_36567,N_37046);
and U38841 (N_38841,N_35076,N_35823);
and U38842 (N_38842,N_36874,N_37497);
nor U38843 (N_38843,N_37335,N_36250);
or U38844 (N_38844,N_36785,N_36029);
xnor U38845 (N_38845,N_35702,N_36212);
xor U38846 (N_38846,N_37414,N_37407);
xnor U38847 (N_38847,N_35040,N_35733);
and U38848 (N_38848,N_36063,N_37461);
and U38849 (N_38849,N_35350,N_36569);
or U38850 (N_38850,N_36917,N_35425);
and U38851 (N_38851,N_35470,N_37318);
or U38852 (N_38852,N_37344,N_36545);
and U38853 (N_38853,N_36161,N_35207);
or U38854 (N_38854,N_35063,N_36001);
nand U38855 (N_38855,N_36644,N_36908);
xnor U38856 (N_38856,N_36575,N_36227);
nand U38857 (N_38857,N_36791,N_36900);
nor U38858 (N_38858,N_37001,N_35270);
nor U38859 (N_38859,N_35613,N_35463);
or U38860 (N_38860,N_35517,N_36987);
nand U38861 (N_38861,N_36857,N_35494);
nor U38862 (N_38862,N_36544,N_37295);
and U38863 (N_38863,N_37344,N_36252);
or U38864 (N_38864,N_35339,N_37049);
xnor U38865 (N_38865,N_36617,N_36087);
or U38866 (N_38866,N_37318,N_35116);
nand U38867 (N_38867,N_36949,N_37484);
and U38868 (N_38868,N_36025,N_37056);
nand U38869 (N_38869,N_37282,N_36176);
xnor U38870 (N_38870,N_35853,N_35624);
and U38871 (N_38871,N_35027,N_35304);
nand U38872 (N_38872,N_35534,N_36460);
nand U38873 (N_38873,N_36114,N_35453);
or U38874 (N_38874,N_37200,N_37024);
and U38875 (N_38875,N_35004,N_36637);
xor U38876 (N_38876,N_35315,N_35511);
xnor U38877 (N_38877,N_36505,N_37013);
or U38878 (N_38878,N_37444,N_36719);
and U38879 (N_38879,N_37334,N_36132);
or U38880 (N_38880,N_36101,N_36044);
nor U38881 (N_38881,N_35948,N_36390);
or U38882 (N_38882,N_35216,N_35902);
xor U38883 (N_38883,N_37364,N_35094);
xnor U38884 (N_38884,N_35330,N_36737);
xor U38885 (N_38885,N_37146,N_35303);
or U38886 (N_38886,N_35333,N_35825);
or U38887 (N_38887,N_36495,N_35619);
nand U38888 (N_38888,N_36305,N_35874);
or U38889 (N_38889,N_35425,N_35131);
nand U38890 (N_38890,N_36981,N_36443);
nor U38891 (N_38891,N_35631,N_36679);
nand U38892 (N_38892,N_36539,N_35570);
xor U38893 (N_38893,N_36045,N_35854);
xor U38894 (N_38894,N_37147,N_35629);
xor U38895 (N_38895,N_35801,N_37251);
xnor U38896 (N_38896,N_36300,N_37358);
nand U38897 (N_38897,N_36534,N_36070);
or U38898 (N_38898,N_36648,N_37386);
nand U38899 (N_38899,N_37022,N_36466);
or U38900 (N_38900,N_37264,N_35741);
nor U38901 (N_38901,N_37473,N_36766);
and U38902 (N_38902,N_35107,N_36128);
nand U38903 (N_38903,N_36853,N_36180);
nor U38904 (N_38904,N_36433,N_36206);
nand U38905 (N_38905,N_36221,N_36920);
or U38906 (N_38906,N_35078,N_37044);
nand U38907 (N_38907,N_36468,N_37098);
nand U38908 (N_38908,N_35080,N_35584);
nand U38909 (N_38909,N_36151,N_35520);
or U38910 (N_38910,N_36310,N_35059);
nor U38911 (N_38911,N_35412,N_35926);
and U38912 (N_38912,N_35840,N_35565);
xor U38913 (N_38913,N_36766,N_37216);
or U38914 (N_38914,N_36972,N_36638);
or U38915 (N_38915,N_35650,N_37272);
or U38916 (N_38916,N_37316,N_37031);
or U38917 (N_38917,N_35099,N_36121);
and U38918 (N_38918,N_36415,N_35340);
nor U38919 (N_38919,N_37034,N_37031);
and U38920 (N_38920,N_35100,N_37281);
and U38921 (N_38921,N_35816,N_35461);
or U38922 (N_38922,N_36078,N_37473);
nand U38923 (N_38923,N_35803,N_36208);
and U38924 (N_38924,N_36702,N_36063);
xnor U38925 (N_38925,N_35094,N_35734);
xor U38926 (N_38926,N_35313,N_36199);
nand U38927 (N_38927,N_36849,N_35740);
and U38928 (N_38928,N_36898,N_37195);
and U38929 (N_38929,N_37388,N_35205);
nand U38930 (N_38930,N_35111,N_37351);
or U38931 (N_38931,N_35961,N_35986);
and U38932 (N_38932,N_36182,N_35796);
nor U38933 (N_38933,N_36028,N_36986);
nor U38934 (N_38934,N_37131,N_35246);
or U38935 (N_38935,N_35654,N_35076);
or U38936 (N_38936,N_37397,N_36382);
and U38937 (N_38937,N_36688,N_36737);
nor U38938 (N_38938,N_36899,N_35639);
and U38939 (N_38939,N_36966,N_36139);
xor U38940 (N_38940,N_36552,N_35560);
and U38941 (N_38941,N_37175,N_37003);
and U38942 (N_38942,N_36207,N_35821);
and U38943 (N_38943,N_36600,N_36657);
or U38944 (N_38944,N_35594,N_35130);
nor U38945 (N_38945,N_35678,N_36148);
xor U38946 (N_38946,N_36739,N_36280);
or U38947 (N_38947,N_35576,N_35906);
or U38948 (N_38948,N_36156,N_36852);
and U38949 (N_38949,N_37189,N_36585);
and U38950 (N_38950,N_36327,N_37283);
nor U38951 (N_38951,N_35760,N_37492);
or U38952 (N_38952,N_37465,N_35268);
and U38953 (N_38953,N_35815,N_36204);
or U38954 (N_38954,N_35346,N_36612);
nor U38955 (N_38955,N_36835,N_35543);
and U38956 (N_38956,N_36551,N_35924);
nand U38957 (N_38957,N_37165,N_35018);
nand U38958 (N_38958,N_36448,N_35808);
nand U38959 (N_38959,N_36612,N_35783);
or U38960 (N_38960,N_35827,N_35950);
and U38961 (N_38961,N_35180,N_37443);
and U38962 (N_38962,N_36857,N_36472);
nand U38963 (N_38963,N_35505,N_35687);
xnor U38964 (N_38964,N_36429,N_36499);
nand U38965 (N_38965,N_37140,N_36676);
nand U38966 (N_38966,N_35467,N_37469);
and U38967 (N_38967,N_35527,N_35358);
nor U38968 (N_38968,N_35934,N_37259);
xor U38969 (N_38969,N_35872,N_36554);
and U38970 (N_38970,N_36817,N_35076);
or U38971 (N_38971,N_35596,N_35694);
nor U38972 (N_38972,N_37112,N_36758);
xor U38973 (N_38973,N_35626,N_37060);
xnor U38974 (N_38974,N_37219,N_35937);
nor U38975 (N_38975,N_36038,N_36526);
xor U38976 (N_38976,N_37063,N_36621);
nand U38977 (N_38977,N_37135,N_37111);
or U38978 (N_38978,N_35153,N_36894);
xnor U38979 (N_38979,N_36551,N_37445);
and U38980 (N_38980,N_35932,N_37330);
nand U38981 (N_38981,N_36187,N_35164);
or U38982 (N_38982,N_35849,N_36515);
nand U38983 (N_38983,N_36807,N_35403);
and U38984 (N_38984,N_36300,N_35936);
and U38985 (N_38985,N_36807,N_37403);
and U38986 (N_38986,N_36010,N_35841);
nand U38987 (N_38987,N_36388,N_35196);
nor U38988 (N_38988,N_36270,N_35866);
nor U38989 (N_38989,N_37243,N_37301);
xor U38990 (N_38990,N_37237,N_35591);
and U38991 (N_38991,N_36374,N_37308);
nand U38992 (N_38992,N_35166,N_37313);
nor U38993 (N_38993,N_37229,N_35375);
nand U38994 (N_38994,N_37454,N_37438);
or U38995 (N_38995,N_37273,N_37408);
or U38996 (N_38996,N_35246,N_37476);
xnor U38997 (N_38997,N_36483,N_37111);
nor U38998 (N_38998,N_37307,N_36543);
nand U38999 (N_38999,N_35356,N_35831);
and U39000 (N_39000,N_36827,N_37313);
and U39001 (N_39001,N_35134,N_35101);
and U39002 (N_39002,N_35479,N_35628);
nand U39003 (N_39003,N_35784,N_37390);
nor U39004 (N_39004,N_36170,N_35699);
xor U39005 (N_39005,N_36467,N_35965);
and U39006 (N_39006,N_37161,N_35322);
or U39007 (N_39007,N_35579,N_36018);
nand U39008 (N_39008,N_35325,N_36377);
nor U39009 (N_39009,N_36989,N_36125);
nand U39010 (N_39010,N_35006,N_35440);
and U39011 (N_39011,N_37077,N_36659);
xnor U39012 (N_39012,N_35131,N_37444);
nor U39013 (N_39013,N_35618,N_37251);
or U39014 (N_39014,N_35561,N_36298);
or U39015 (N_39015,N_36727,N_35321);
xnor U39016 (N_39016,N_37333,N_35895);
nand U39017 (N_39017,N_37479,N_35973);
nor U39018 (N_39018,N_35581,N_36570);
xor U39019 (N_39019,N_35320,N_35728);
nor U39020 (N_39020,N_37418,N_36439);
nand U39021 (N_39021,N_36156,N_36155);
or U39022 (N_39022,N_35634,N_37215);
or U39023 (N_39023,N_37288,N_35014);
xnor U39024 (N_39024,N_36391,N_35513);
xnor U39025 (N_39025,N_35630,N_36251);
nor U39026 (N_39026,N_36248,N_36209);
xor U39027 (N_39027,N_36295,N_36786);
xnor U39028 (N_39028,N_36377,N_36259);
nand U39029 (N_39029,N_36988,N_36671);
and U39030 (N_39030,N_35706,N_36547);
and U39031 (N_39031,N_36555,N_35232);
and U39032 (N_39032,N_35942,N_36145);
nand U39033 (N_39033,N_37321,N_35262);
nand U39034 (N_39034,N_35477,N_36052);
nand U39035 (N_39035,N_35292,N_36927);
nand U39036 (N_39036,N_35139,N_36211);
and U39037 (N_39037,N_36074,N_37439);
or U39038 (N_39038,N_36838,N_37435);
or U39039 (N_39039,N_36888,N_35983);
nor U39040 (N_39040,N_36978,N_36821);
or U39041 (N_39041,N_35724,N_35556);
or U39042 (N_39042,N_35771,N_37066);
xnor U39043 (N_39043,N_36790,N_36051);
and U39044 (N_39044,N_36381,N_36314);
and U39045 (N_39045,N_35463,N_36817);
and U39046 (N_39046,N_35550,N_35243);
or U39047 (N_39047,N_37234,N_35257);
or U39048 (N_39048,N_35924,N_36874);
and U39049 (N_39049,N_36742,N_35623);
nand U39050 (N_39050,N_37449,N_36848);
nand U39051 (N_39051,N_37286,N_35227);
nand U39052 (N_39052,N_36229,N_36408);
xnor U39053 (N_39053,N_35542,N_36945);
xor U39054 (N_39054,N_36759,N_35039);
nand U39055 (N_39055,N_36785,N_35461);
or U39056 (N_39056,N_36181,N_36627);
and U39057 (N_39057,N_37253,N_36400);
or U39058 (N_39058,N_37450,N_35333);
nor U39059 (N_39059,N_37484,N_35700);
or U39060 (N_39060,N_37016,N_36604);
xor U39061 (N_39061,N_36558,N_35675);
xor U39062 (N_39062,N_36793,N_35164);
xnor U39063 (N_39063,N_36212,N_35816);
or U39064 (N_39064,N_36601,N_36834);
nand U39065 (N_39065,N_36975,N_36861);
and U39066 (N_39066,N_35255,N_37015);
nor U39067 (N_39067,N_36807,N_36288);
nor U39068 (N_39068,N_35919,N_35590);
nor U39069 (N_39069,N_35682,N_37008);
xnor U39070 (N_39070,N_36402,N_36661);
xnor U39071 (N_39071,N_35350,N_37312);
nand U39072 (N_39072,N_36783,N_35458);
and U39073 (N_39073,N_35725,N_35610);
or U39074 (N_39074,N_36295,N_37177);
xor U39075 (N_39075,N_37106,N_37076);
or U39076 (N_39076,N_35767,N_35107);
and U39077 (N_39077,N_35669,N_36389);
xnor U39078 (N_39078,N_36814,N_35500);
or U39079 (N_39079,N_35567,N_37375);
xnor U39080 (N_39080,N_35122,N_37062);
or U39081 (N_39081,N_36591,N_36224);
nand U39082 (N_39082,N_35375,N_37357);
and U39083 (N_39083,N_35022,N_35407);
nor U39084 (N_39084,N_35341,N_37243);
and U39085 (N_39085,N_37440,N_37118);
nor U39086 (N_39086,N_36158,N_35445);
nand U39087 (N_39087,N_35595,N_37351);
xnor U39088 (N_39088,N_35852,N_36324);
or U39089 (N_39089,N_37083,N_35978);
and U39090 (N_39090,N_37148,N_35914);
or U39091 (N_39091,N_36801,N_35705);
or U39092 (N_39092,N_36364,N_35636);
or U39093 (N_39093,N_37122,N_35938);
and U39094 (N_39094,N_35721,N_36753);
xnor U39095 (N_39095,N_35967,N_37214);
nor U39096 (N_39096,N_36341,N_36058);
nand U39097 (N_39097,N_36230,N_35237);
or U39098 (N_39098,N_36770,N_36823);
nand U39099 (N_39099,N_36631,N_35307);
and U39100 (N_39100,N_37044,N_37179);
nor U39101 (N_39101,N_35965,N_36449);
or U39102 (N_39102,N_36044,N_36303);
or U39103 (N_39103,N_36032,N_35291);
nand U39104 (N_39104,N_35872,N_36163);
nand U39105 (N_39105,N_35485,N_36254);
and U39106 (N_39106,N_36579,N_35310);
or U39107 (N_39107,N_36955,N_35948);
and U39108 (N_39108,N_35422,N_36130);
and U39109 (N_39109,N_35941,N_35531);
and U39110 (N_39110,N_36676,N_36110);
or U39111 (N_39111,N_35934,N_36880);
and U39112 (N_39112,N_36851,N_37344);
nor U39113 (N_39113,N_37010,N_35560);
or U39114 (N_39114,N_36006,N_35602);
nor U39115 (N_39115,N_36694,N_36791);
nor U39116 (N_39116,N_37273,N_36418);
or U39117 (N_39117,N_35073,N_35355);
nor U39118 (N_39118,N_37142,N_36491);
and U39119 (N_39119,N_35004,N_36293);
xor U39120 (N_39120,N_37254,N_36156);
and U39121 (N_39121,N_36124,N_36829);
nor U39122 (N_39122,N_37450,N_36541);
xor U39123 (N_39123,N_37031,N_36767);
xor U39124 (N_39124,N_35417,N_37025);
xor U39125 (N_39125,N_37288,N_35392);
nand U39126 (N_39126,N_36167,N_35700);
and U39127 (N_39127,N_36624,N_35895);
nor U39128 (N_39128,N_35373,N_36026);
nor U39129 (N_39129,N_37233,N_36062);
xnor U39130 (N_39130,N_35435,N_36595);
nor U39131 (N_39131,N_35637,N_37183);
nor U39132 (N_39132,N_36682,N_35459);
xnor U39133 (N_39133,N_35781,N_35702);
nand U39134 (N_39134,N_36791,N_37150);
and U39135 (N_39135,N_36082,N_35614);
xnor U39136 (N_39136,N_36922,N_36095);
nand U39137 (N_39137,N_35312,N_36693);
nor U39138 (N_39138,N_35910,N_36121);
and U39139 (N_39139,N_36193,N_37420);
xnor U39140 (N_39140,N_36471,N_36576);
nand U39141 (N_39141,N_35564,N_35724);
nand U39142 (N_39142,N_36998,N_35177);
nor U39143 (N_39143,N_36478,N_36733);
and U39144 (N_39144,N_36785,N_37198);
or U39145 (N_39145,N_36015,N_35771);
xnor U39146 (N_39146,N_35597,N_36957);
and U39147 (N_39147,N_36999,N_35407);
xnor U39148 (N_39148,N_37242,N_35058);
and U39149 (N_39149,N_37133,N_37340);
or U39150 (N_39150,N_37237,N_35961);
nand U39151 (N_39151,N_35296,N_36085);
nor U39152 (N_39152,N_35371,N_37257);
and U39153 (N_39153,N_35804,N_35971);
nand U39154 (N_39154,N_36104,N_36308);
nor U39155 (N_39155,N_37198,N_37212);
xor U39156 (N_39156,N_35361,N_36362);
nor U39157 (N_39157,N_35157,N_36251);
xor U39158 (N_39158,N_35392,N_35045);
or U39159 (N_39159,N_37191,N_36605);
and U39160 (N_39160,N_37059,N_35374);
xnor U39161 (N_39161,N_35730,N_35946);
and U39162 (N_39162,N_36650,N_35024);
nor U39163 (N_39163,N_37272,N_36929);
or U39164 (N_39164,N_37388,N_36825);
nand U39165 (N_39165,N_35135,N_35405);
nor U39166 (N_39166,N_36354,N_36976);
nor U39167 (N_39167,N_36344,N_35885);
and U39168 (N_39168,N_36440,N_36765);
and U39169 (N_39169,N_36920,N_35611);
nor U39170 (N_39170,N_36158,N_35240);
or U39171 (N_39171,N_36961,N_37485);
or U39172 (N_39172,N_35853,N_36765);
nor U39173 (N_39173,N_36887,N_36437);
nand U39174 (N_39174,N_35822,N_36669);
and U39175 (N_39175,N_36034,N_36235);
nor U39176 (N_39176,N_35564,N_37281);
nand U39177 (N_39177,N_35067,N_37035);
xor U39178 (N_39178,N_36800,N_35505);
xnor U39179 (N_39179,N_35339,N_36639);
nand U39180 (N_39180,N_35208,N_37325);
or U39181 (N_39181,N_36544,N_36303);
or U39182 (N_39182,N_36540,N_35217);
nor U39183 (N_39183,N_35592,N_36028);
and U39184 (N_39184,N_35557,N_35741);
xnor U39185 (N_39185,N_36892,N_35692);
or U39186 (N_39186,N_35320,N_35735);
nand U39187 (N_39187,N_37053,N_36001);
or U39188 (N_39188,N_37331,N_36269);
or U39189 (N_39189,N_37242,N_36233);
xor U39190 (N_39190,N_35993,N_35317);
nor U39191 (N_39191,N_35260,N_35564);
nor U39192 (N_39192,N_35333,N_35160);
or U39193 (N_39193,N_36601,N_35379);
or U39194 (N_39194,N_37090,N_35551);
or U39195 (N_39195,N_35800,N_36995);
and U39196 (N_39196,N_36236,N_36615);
and U39197 (N_39197,N_36418,N_36989);
nor U39198 (N_39198,N_36468,N_35335);
nand U39199 (N_39199,N_36667,N_36057);
nand U39200 (N_39200,N_35153,N_36318);
or U39201 (N_39201,N_35484,N_35143);
xor U39202 (N_39202,N_37026,N_37195);
xor U39203 (N_39203,N_37216,N_35950);
or U39204 (N_39204,N_35275,N_36884);
nor U39205 (N_39205,N_35229,N_35176);
nor U39206 (N_39206,N_35202,N_36975);
xnor U39207 (N_39207,N_35641,N_35320);
and U39208 (N_39208,N_36718,N_35344);
and U39209 (N_39209,N_36638,N_35870);
xnor U39210 (N_39210,N_36047,N_36585);
nand U39211 (N_39211,N_35106,N_35891);
nand U39212 (N_39212,N_35966,N_35004);
xnor U39213 (N_39213,N_35754,N_35099);
xor U39214 (N_39214,N_36714,N_36956);
or U39215 (N_39215,N_35943,N_36734);
xor U39216 (N_39216,N_36906,N_35706);
or U39217 (N_39217,N_36641,N_36083);
xnor U39218 (N_39218,N_35498,N_37139);
or U39219 (N_39219,N_35887,N_35283);
or U39220 (N_39220,N_36790,N_37408);
xnor U39221 (N_39221,N_37310,N_36235);
and U39222 (N_39222,N_35192,N_37411);
nor U39223 (N_39223,N_35198,N_35526);
xor U39224 (N_39224,N_35536,N_36065);
and U39225 (N_39225,N_35563,N_35777);
xnor U39226 (N_39226,N_36441,N_36010);
or U39227 (N_39227,N_36977,N_37259);
nor U39228 (N_39228,N_35425,N_36010);
and U39229 (N_39229,N_36655,N_35409);
xor U39230 (N_39230,N_36960,N_35722);
and U39231 (N_39231,N_37286,N_35911);
xnor U39232 (N_39232,N_35590,N_36359);
nor U39233 (N_39233,N_36966,N_36142);
xnor U39234 (N_39234,N_36409,N_35012);
nand U39235 (N_39235,N_37457,N_37245);
nor U39236 (N_39236,N_35047,N_36285);
or U39237 (N_39237,N_37091,N_35041);
or U39238 (N_39238,N_36976,N_37386);
xnor U39239 (N_39239,N_35237,N_36211);
or U39240 (N_39240,N_35737,N_36678);
nand U39241 (N_39241,N_35146,N_36680);
and U39242 (N_39242,N_35410,N_37258);
or U39243 (N_39243,N_35334,N_35450);
nand U39244 (N_39244,N_36016,N_35584);
or U39245 (N_39245,N_35329,N_36931);
nand U39246 (N_39246,N_35799,N_35265);
nor U39247 (N_39247,N_36720,N_35322);
or U39248 (N_39248,N_37346,N_37026);
or U39249 (N_39249,N_36725,N_35277);
nand U39250 (N_39250,N_35684,N_36659);
nor U39251 (N_39251,N_35492,N_35849);
or U39252 (N_39252,N_37337,N_36524);
and U39253 (N_39253,N_37382,N_35430);
nor U39254 (N_39254,N_36342,N_35571);
or U39255 (N_39255,N_35625,N_35199);
nand U39256 (N_39256,N_35110,N_36982);
xnor U39257 (N_39257,N_35302,N_36502);
nor U39258 (N_39258,N_36910,N_37268);
xnor U39259 (N_39259,N_37497,N_36934);
nor U39260 (N_39260,N_36893,N_35069);
nand U39261 (N_39261,N_35982,N_37356);
nor U39262 (N_39262,N_36843,N_36068);
and U39263 (N_39263,N_36453,N_35654);
nand U39264 (N_39264,N_36327,N_36195);
nand U39265 (N_39265,N_36377,N_37464);
xnor U39266 (N_39266,N_37080,N_35525);
nor U39267 (N_39267,N_36787,N_37056);
and U39268 (N_39268,N_35330,N_35594);
or U39269 (N_39269,N_35493,N_37420);
xor U39270 (N_39270,N_35367,N_35005);
or U39271 (N_39271,N_37063,N_36966);
nand U39272 (N_39272,N_37164,N_37331);
and U39273 (N_39273,N_37066,N_35908);
nor U39274 (N_39274,N_36780,N_36255);
and U39275 (N_39275,N_35351,N_36271);
xnor U39276 (N_39276,N_35673,N_35930);
nor U39277 (N_39277,N_35307,N_35506);
and U39278 (N_39278,N_35763,N_36738);
and U39279 (N_39279,N_36507,N_36464);
nand U39280 (N_39280,N_35041,N_35673);
nor U39281 (N_39281,N_35503,N_36695);
nand U39282 (N_39282,N_35072,N_36315);
or U39283 (N_39283,N_35425,N_36734);
and U39284 (N_39284,N_35098,N_35806);
and U39285 (N_39285,N_36657,N_36351);
xor U39286 (N_39286,N_37147,N_35670);
nand U39287 (N_39287,N_36627,N_37298);
or U39288 (N_39288,N_36128,N_37437);
and U39289 (N_39289,N_36400,N_37335);
and U39290 (N_39290,N_35211,N_36150);
xnor U39291 (N_39291,N_36412,N_36457);
nand U39292 (N_39292,N_35391,N_35586);
nor U39293 (N_39293,N_35984,N_35244);
or U39294 (N_39294,N_36535,N_35613);
or U39295 (N_39295,N_36353,N_37466);
or U39296 (N_39296,N_35311,N_37113);
xnor U39297 (N_39297,N_36891,N_36425);
nand U39298 (N_39298,N_35837,N_35232);
nand U39299 (N_39299,N_35286,N_36902);
nor U39300 (N_39300,N_36170,N_36264);
xor U39301 (N_39301,N_36787,N_36761);
xnor U39302 (N_39302,N_35446,N_35293);
and U39303 (N_39303,N_35966,N_35579);
xor U39304 (N_39304,N_35914,N_36774);
and U39305 (N_39305,N_37484,N_35571);
and U39306 (N_39306,N_36604,N_36752);
and U39307 (N_39307,N_37443,N_37498);
nand U39308 (N_39308,N_36372,N_36758);
and U39309 (N_39309,N_35204,N_35855);
and U39310 (N_39310,N_37412,N_35560);
and U39311 (N_39311,N_35333,N_37424);
or U39312 (N_39312,N_37115,N_36464);
or U39313 (N_39313,N_36513,N_36991);
and U39314 (N_39314,N_35287,N_36085);
nor U39315 (N_39315,N_35542,N_36891);
nor U39316 (N_39316,N_35023,N_35721);
xnor U39317 (N_39317,N_36799,N_35877);
or U39318 (N_39318,N_35914,N_35654);
nor U39319 (N_39319,N_36283,N_36068);
xnor U39320 (N_39320,N_37341,N_35604);
xnor U39321 (N_39321,N_36734,N_36042);
xor U39322 (N_39322,N_35733,N_35808);
nor U39323 (N_39323,N_36956,N_36605);
nand U39324 (N_39324,N_36584,N_36340);
nor U39325 (N_39325,N_36331,N_35207);
nand U39326 (N_39326,N_35831,N_36195);
and U39327 (N_39327,N_37223,N_37016);
nor U39328 (N_39328,N_36607,N_35195);
and U39329 (N_39329,N_35466,N_35852);
nor U39330 (N_39330,N_36565,N_36484);
xnor U39331 (N_39331,N_36838,N_37037);
nor U39332 (N_39332,N_35123,N_35601);
xnor U39333 (N_39333,N_36560,N_35639);
xnor U39334 (N_39334,N_35196,N_37218);
xnor U39335 (N_39335,N_35907,N_35621);
xor U39336 (N_39336,N_35874,N_36006);
or U39337 (N_39337,N_35375,N_36058);
and U39338 (N_39338,N_37426,N_35310);
nand U39339 (N_39339,N_35634,N_35291);
or U39340 (N_39340,N_37344,N_36988);
or U39341 (N_39341,N_36353,N_35283);
and U39342 (N_39342,N_36808,N_36498);
xnor U39343 (N_39343,N_35106,N_36655);
nand U39344 (N_39344,N_35191,N_37229);
and U39345 (N_39345,N_36002,N_36743);
or U39346 (N_39346,N_36167,N_36501);
nor U39347 (N_39347,N_36298,N_36084);
nand U39348 (N_39348,N_35583,N_35837);
or U39349 (N_39349,N_36259,N_36543);
xnor U39350 (N_39350,N_37012,N_36357);
xnor U39351 (N_39351,N_37241,N_36988);
or U39352 (N_39352,N_36628,N_35253);
nand U39353 (N_39353,N_35257,N_35931);
nor U39354 (N_39354,N_35316,N_35034);
nor U39355 (N_39355,N_36393,N_37088);
nor U39356 (N_39356,N_35516,N_35259);
nor U39357 (N_39357,N_37363,N_36146);
nand U39358 (N_39358,N_35747,N_37397);
and U39359 (N_39359,N_35149,N_35404);
or U39360 (N_39360,N_37394,N_36795);
xnor U39361 (N_39361,N_35905,N_36262);
or U39362 (N_39362,N_37293,N_36106);
nor U39363 (N_39363,N_36529,N_35353);
xor U39364 (N_39364,N_36541,N_37109);
and U39365 (N_39365,N_36147,N_35186);
nand U39366 (N_39366,N_35026,N_35650);
nand U39367 (N_39367,N_37033,N_36442);
nor U39368 (N_39368,N_36783,N_36436);
nor U39369 (N_39369,N_35243,N_35764);
xnor U39370 (N_39370,N_35475,N_36307);
nor U39371 (N_39371,N_36943,N_36646);
nand U39372 (N_39372,N_36869,N_35504);
and U39373 (N_39373,N_37265,N_37356);
nor U39374 (N_39374,N_36045,N_35518);
nand U39375 (N_39375,N_35833,N_36028);
xnor U39376 (N_39376,N_36841,N_35850);
nor U39377 (N_39377,N_37306,N_36578);
nor U39378 (N_39378,N_36648,N_36706);
xor U39379 (N_39379,N_36918,N_37140);
nand U39380 (N_39380,N_35985,N_35706);
and U39381 (N_39381,N_35449,N_35105);
nor U39382 (N_39382,N_37302,N_37315);
and U39383 (N_39383,N_36607,N_36898);
and U39384 (N_39384,N_36832,N_36098);
and U39385 (N_39385,N_37232,N_36253);
xor U39386 (N_39386,N_35677,N_37329);
or U39387 (N_39387,N_35360,N_36976);
or U39388 (N_39388,N_35585,N_35226);
or U39389 (N_39389,N_35417,N_35236);
xor U39390 (N_39390,N_36538,N_35264);
nor U39391 (N_39391,N_37497,N_35291);
or U39392 (N_39392,N_35191,N_35136);
and U39393 (N_39393,N_35953,N_37265);
or U39394 (N_39394,N_35533,N_36040);
xnor U39395 (N_39395,N_36809,N_35366);
and U39396 (N_39396,N_37057,N_35371);
and U39397 (N_39397,N_35224,N_36308);
xor U39398 (N_39398,N_35964,N_36326);
xnor U39399 (N_39399,N_36357,N_35025);
or U39400 (N_39400,N_35943,N_35754);
nand U39401 (N_39401,N_36920,N_35021);
nand U39402 (N_39402,N_35774,N_36267);
nand U39403 (N_39403,N_36668,N_35600);
nand U39404 (N_39404,N_37162,N_37172);
and U39405 (N_39405,N_36076,N_35353);
or U39406 (N_39406,N_35363,N_36048);
nand U39407 (N_39407,N_37417,N_36131);
xnor U39408 (N_39408,N_35914,N_35177);
and U39409 (N_39409,N_35909,N_37431);
and U39410 (N_39410,N_36740,N_36298);
nand U39411 (N_39411,N_37217,N_35606);
and U39412 (N_39412,N_36510,N_37300);
or U39413 (N_39413,N_35262,N_35694);
and U39414 (N_39414,N_35671,N_35676);
nor U39415 (N_39415,N_37368,N_36047);
and U39416 (N_39416,N_35249,N_35371);
nor U39417 (N_39417,N_37236,N_35253);
nand U39418 (N_39418,N_36692,N_36051);
or U39419 (N_39419,N_37411,N_37298);
and U39420 (N_39420,N_36692,N_36175);
or U39421 (N_39421,N_36654,N_37117);
or U39422 (N_39422,N_37029,N_35444);
nand U39423 (N_39423,N_35496,N_37398);
nand U39424 (N_39424,N_35634,N_36742);
and U39425 (N_39425,N_37272,N_36762);
xor U39426 (N_39426,N_35168,N_35317);
and U39427 (N_39427,N_37246,N_35949);
nand U39428 (N_39428,N_35767,N_35226);
nand U39429 (N_39429,N_36194,N_36107);
nor U39430 (N_39430,N_36452,N_36320);
nand U39431 (N_39431,N_35176,N_37387);
and U39432 (N_39432,N_35507,N_37281);
nor U39433 (N_39433,N_35795,N_36183);
or U39434 (N_39434,N_36662,N_35999);
or U39435 (N_39435,N_35602,N_37454);
xor U39436 (N_39436,N_36943,N_35373);
nor U39437 (N_39437,N_36847,N_35240);
nand U39438 (N_39438,N_36331,N_36479);
or U39439 (N_39439,N_35002,N_36382);
and U39440 (N_39440,N_35277,N_36020);
and U39441 (N_39441,N_36266,N_36295);
and U39442 (N_39442,N_35000,N_36579);
or U39443 (N_39443,N_35040,N_35355);
or U39444 (N_39444,N_36637,N_36114);
xor U39445 (N_39445,N_37060,N_37418);
or U39446 (N_39446,N_36098,N_35306);
xnor U39447 (N_39447,N_35219,N_35691);
nor U39448 (N_39448,N_36533,N_37068);
nand U39449 (N_39449,N_35076,N_35014);
nor U39450 (N_39450,N_35119,N_35632);
or U39451 (N_39451,N_37156,N_37167);
nand U39452 (N_39452,N_37419,N_37228);
nand U39453 (N_39453,N_36481,N_36089);
nor U39454 (N_39454,N_35003,N_35165);
and U39455 (N_39455,N_35104,N_36387);
nor U39456 (N_39456,N_36153,N_37452);
xnor U39457 (N_39457,N_36197,N_36805);
xnor U39458 (N_39458,N_36350,N_35266);
xor U39459 (N_39459,N_36523,N_36305);
xnor U39460 (N_39460,N_36050,N_37083);
or U39461 (N_39461,N_37391,N_35066);
nand U39462 (N_39462,N_36931,N_35445);
or U39463 (N_39463,N_36194,N_37244);
xnor U39464 (N_39464,N_35519,N_35108);
nand U39465 (N_39465,N_37444,N_36896);
and U39466 (N_39466,N_36007,N_37080);
and U39467 (N_39467,N_36629,N_37414);
xor U39468 (N_39468,N_36207,N_36357);
xnor U39469 (N_39469,N_36778,N_37356);
nor U39470 (N_39470,N_36781,N_35895);
nor U39471 (N_39471,N_36225,N_36589);
or U39472 (N_39472,N_36739,N_36487);
and U39473 (N_39473,N_35316,N_37252);
or U39474 (N_39474,N_35502,N_35685);
xor U39475 (N_39475,N_37418,N_36615);
nor U39476 (N_39476,N_35533,N_35920);
xnor U39477 (N_39477,N_35674,N_37159);
nor U39478 (N_39478,N_35860,N_36926);
or U39479 (N_39479,N_35328,N_35708);
nor U39480 (N_39480,N_37374,N_36750);
xor U39481 (N_39481,N_35169,N_35114);
nand U39482 (N_39482,N_36581,N_35653);
nand U39483 (N_39483,N_36162,N_36028);
nor U39484 (N_39484,N_35596,N_37399);
nand U39485 (N_39485,N_36766,N_35351);
xnor U39486 (N_39486,N_36672,N_36710);
nand U39487 (N_39487,N_35549,N_36145);
nand U39488 (N_39488,N_35113,N_35112);
or U39489 (N_39489,N_35208,N_36717);
or U39490 (N_39490,N_35643,N_36817);
xnor U39491 (N_39491,N_37137,N_36787);
or U39492 (N_39492,N_37163,N_36682);
xor U39493 (N_39493,N_36236,N_35709);
nand U39494 (N_39494,N_36001,N_35886);
xor U39495 (N_39495,N_36661,N_36623);
xnor U39496 (N_39496,N_35840,N_36362);
xnor U39497 (N_39497,N_36209,N_37030);
nand U39498 (N_39498,N_35418,N_37116);
nor U39499 (N_39499,N_36292,N_35897);
nor U39500 (N_39500,N_36113,N_37266);
or U39501 (N_39501,N_35068,N_35646);
xnor U39502 (N_39502,N_36291,N_36663);
or U39503 (N_39503,N_35187,N_35403);
or U39504 (N_39504,N_36231,N_36890);
nor U39505 (N_39505,N_37285,N_36146);
nor U39506 (N_39506,N_35667,N_36093);
nand U39507 (N_39507,N_36705,N_35860);
nand U39508 (N_39508,N_37152,N_35377);
and U39509 (N_39509,N_35217,N_36332);
nand U39510 (N_39510,N_36127,N_36605);
and U39511 (N_39511,N_36782,N_37367);
or U39512 (N_39512,N_37285,N_35479);
nor U39513 (N_39513,N_36848,N_35937);
nor U39514 (N_39514,N_36579,N_36392);
nor U39515 (N_39515,N_36337,N_36334);
nand U39516 (N_39516,N_36615,N_36197);
xor U39517 (N_39517,N_35840,N_36823);
and U39518 (N_39518,N_36148,N_37353);
xor U39519 (N_39519,N_37493,N_35637);
and U39520 (N_39520,N_35917,N_36597);
nor U39521 (N_39521,N_36267,N_35878);
or U39522 (N_39522,N_36383,N_36049);
xnor U39523 (N_39523,N_36497,N_36192);
nor U39524 (N_39524,N_35125,N_35311);
and U39525 (N_39525,N_36163,N_35680);
xor U39526 (N_39526,N_37399,N_36856);
xor U39527 (N_39527,N_36086,N_35939);
and U39528 (N_39528,N_37243,N_36345);
or U39529 (N_39529,N_36404,N_36356);
nor U39530 (N_39530,N_35857,N_35159);
nand U39531 (N_39531,N_37099,N_37369);
nand U39532 (N_39532,N_35929,N_35506);
and U39533 (N_39533,N_35265,N_35003);
and U39534 (N_39534,N_35741,N_36582);
xnor U39535 (N_39535,N_35136,N_35990);
nor U39536 (N_39536,N_36449,N_37093);
or U39537 (N_39537,N_35974,N_36861);
nand U39538 (N_39538,N_36411,N_36481);
nor U39539 (N_39539,N_36976,N_37300);
nor U39540 (N_39540,N_37309,N_36234);
and U39541 (N_39541,N_36104,N_37106);
nor U39542 (N_39542,N_36006,N_35627);
and U39543 (N_39543,N_35196,N_36073);
and U39544 (N_39544,N_35129,N_35491);
or U39545 (N_39545,N_35211,N_35537);
and U39546 (N_39546,N_35163,N_35724);
xnor U39547 (N_39547,N_35510,N_36191);
nor U39548 (N_39548,N_35477,N_35369);
nor U39549 (N_39549,N_35086,N_37118);
or U39550 (N_39550,N_36879,N_36331);
nor U39551 (N_39551,N_35365,N_35738);
nor U39552 (N_39552,N_37210,N_36734);
nand U39553 (N_39553,N_35466,N_35002);
nand U39554 (N_39554,N_36892,N_36009);
and U39555 (N_39555,N_35306,N_35484);
nor U39556 (N_39556,N_36002,N_37414);
or U39557 (N_39557,N_37390,N_36638);
or U39558 (N_39558,N_36480,N_36535);
and U39559 (N_39559,N_36085,N_36876);
xnor U39560 (N_39560,N_35713,N_36430);
nand U39561 (N_39561,N_35742,N_36076);
nor U39562 (N_39562,N_35578,N_36338);
or U39563 (N_39563,N_36974,N_35818);
and U39564 (N_39564,N_36505,N_37041);
nor U39565 (N_39565,N_35134,N_35881);
xor U39566 (N_39566,N_37487,N_36874);
xor U39567 (N_39567,N_36369,N_35774);
xnor U39568 (N_39568,N_35480,N_35025);
xnor U39569 (N_39569,N_36675,N_37089);
xor U39570 (N_39570,N_35686,N_36790);
and U39571 (N_39571,N_36215,N_37346);
and U39572 (N_39572,N_35787,N_36321);
or U39573 (N_39573,N_36345,N_35464);
and U39574 (N_39574,N_35327,N_35951);
nand U39575 (N_39575,N_37314,N_36102);
nor U39576 (N_39576,N_37109,N_36610);
xnor U39577 (N_39577,N_35465,N_37146);
and U39578 (N_39578,N_35310,N_35157);
xor U39579 (N_39579,N_36259,N_36126);
nor U39580 (N_39580,N_36596,N_37448);
xor U39581 (N_39581,N_36853,N_36644);
nor U39582 (N_39582,N_36466,N_36597);
nor U39583 (N_39583,N_36911,N_36395);
or U39584 (N_39584,N_37144,N_36491);
xor U39585 (N_39585,N_35474,N_35676);
and U39586 (N_39586,N_37482,N_35450);
nor U39587 (N_39587,N_36205,N_36950);
nand U39588 (N_39588,N_35326,N_37119);
nor U39589 (N_39589,N_37076,N_36736);
and U39590 (N_39590,N_36556,N_35673);
and U39591 (N_39591,N_36116,N_37249);
or U39592 (N_39592,N_35938,N_35165);
and U39593 (N_39593,N_37096,N_35828);
xor U39594 (N_39594,N_36071,N_36522);
nand U39595 (N_39595,N_36522,N_37490);
and U39596 (N_39596,N_36516,N_35527);
xnor U39597 (N_39597,N_36586,N_36742);
xor U39598 (N_39598,N_37409,N_36668);
nand U39599 (N_39599,N_37037,N_36860);
nand U39600 (N_39600,N_37241,N_35073);
xor U39601 (N_39601,N_35123,N_37329);
xnor U39602 (N_39602,N_35641,N_37368);
xor U39603 (N_39603,N_35403,N_36182);
nand U39604 (N_39604,N_36005,N_36605);
nor U39605 (N_39605,N_37485,N_36053);
and U39606 (N_39606,N_36751,N_36072);
or U39607 (N_39607,N_36352,N_35781);
nand U39608 (N_39608,N_35584,N_36068);
xor U39609 (N_39609,N_35833,N_36760);
nor U39610 (N_39610,N_36838,N_37309);
xnor U39611 (N_39611,N_35503,N_37222);
nor U39612 (N_39612,N_36439,N_37442);
nor U39613 (N_39613,N_35393,N_35112);
or U39614 (N_39614,N_36307,N_37066);
nand U39615 (N_39615,N_35069,N_36206);
nor U39616 (N_39616,N_35356,N_37441);
nand U39617 (N_39617,N_36752,N_35979);
nor U39618 (N_39618,N_35522,N_35462);
nand U39619 (N_39619,N_36059,N_36508);
nand U39620 (N_39620,N_37251,N_36552);
xnor U39621 (N_39621,N_37282,N_36676);
xnor U39622 (N_39622,N_35874,N_35792);
or U39623 (N_39623,N_37400,N_35392);
and U39624 (N_39624,N_36758,N_35080);
nand U39625 (N_39625,N_35776,N_35751);
or U39626 (N_39626,N_35138,N_36520);
xor U39627 (N_39627,N_36496,N_35707);
or U39628 (N_39628,N_35463,N_36261);
or U39629 (N_39629,N_36510,N_35156);
or U39630 (N_39630,N_37423,N_35572);
and U39631 (N_39631,N_36459,N_35405);
and U39632 (N_39632,N_36319,N_36823);
and U39633 (N_39633,N_35402,N_36175);
nor U39634 (N_39634,N_37086,N_35228);
nand U39635 (N_39635,N_36973,N_35789);
and U39636 (N_39636,N_37108,N_36955);
nor U39637 (N_39637,N_35914,N_36767);
and U39638 (N_39638,N_36154,N_35593);
xnor U39639 (N_39639,N_37322,N_37037);
xor U39640 (N_39640,N_35344,N_36570);
nand U39641 (N_39641,N_36773,N_36527);
nand U39642 (N_39642,N_35705,N_37167);
or U39643 (N_39643,N_37175,N_36126);
nor U39644 (N_39644,N_35538,N_35047);
and U39645 (N_39645,N_35848,N_37123);
and U39646 (N_39646,N_35652,N_35848);
nor U39647 (N_39647,N_36818,N_35731);
nor U39648 (N_39648,N_35228,N_35946);
xor U39649 (N_39649,N_35961,N_36172);
or U39650 (N_39650,N_35649,N_37408);
nand U39651 (N_39651,N_37464,N_35816);
or U39652 (N_39652,N_36030,N_36062);
nand U39653 (N_39653,N_37063,N_36977);
and U39654 (N_39654,N_36323,N_36968);
xnor U39655 (N_39655,N_36831,N_36139);
xnor U39656 (N_39656,N_36202,N_36504);
and U39657 (N_39657,N_35056,N_36780);
xor U39658 (N_39658,N_37444,N_36066);
nor U39659 (N_39659,N_37479,N_36568);
xnor U39660 (N_39660,N_35350,N_35969);
nor U39661 (N_39661,N_35088,N_35988);
xnor U39662 (N_39662,N_35526,N_35088);
or U39663 (N_39663,N_36151,N_36576);
nand U39664 (N_39664,N_35821,N_36935);
and U39665 (N_39665,N_37377,N_37498);
and U39666 (N_39666,N_35646,N_36711);
xor U39667 (N_39667,N_36059,N_36559);
nor U39668 (N_39668,N_35669,N_36115);
and U39669 (N_39669,N_36809,N_36354);
or U39670 (N_39670,N_36125,N_36756);
nor U39671 (N_39671,N_35846,N_36807);
and U39672 (N_39672,N_37462,N_35522);
nor U39673 (N_39673,N_35983,N_36402);
xor U39674 (N_39674,N_36857,N_37069);
nor U39675 (N_39675,N_37008,N_37462);
xor U39676 (N_39676,N_36362,N_36427);
xnor U39677 (N_39677,N_35110,N_36157);
and U39678 (N_39678,N_35756,N_35077);
nand U39679 (N_39679,N_35715,N_35425);
nor U39680 (N_39680,N_36453,N_36512);
and U39681 (N_39681,N_37483,N_36033);
xor U39682 (N_39682,N_37201,N_37428);
or U39683 (N_39683,N_37072,N_35602);
nand U39684 (N_39684,N_36107,N_36002);
xor U39685 (N_39685,N_35164,N_36483);
xnor U39686 (N_39686,N_35855,N_36193);
or U39687 (N_39687,N_35013,N_36323);
nor U39688 (N_39688,N_35268,N_35859);
or U39689 (N_39689,N_35348,N_36054);
xor U39690 (N_39690,N_37475,N_36260);
and U39691 (N_39691,N_35686,N_37259);
or U39692 (N_39692,N_37348,N_36685);
and U39693 (N_39693,N_35157,N_35596);
nand U39694 (N_39694,N_36695,N_36970);
nor U39695 (N_39695,N_36770,N_35283);
nor U39696 (N_39696,N_36344,N_35848);
nand U39697 (N_39697,N_36673,N_35531);
and U39698 (N_39698,N_35144,N_36440);
xor U39699 (N_39699,N_37306,N_37189);
or U39700 (N_39700,N_36036,N_35639);
nand U39701 (N_39701,N_36945,N_35256);
or U39702 (N_39702,N_35062,N_36284);
nand U39703 (N_39703,N_35843,N_35813);
or U39704 (N_39704,N_37042,N_35416);
or U39705 (N_39705,N_35217,N_35748);
xnor U39706 (N_39706,N_36586,N_36505);
xnor U39707 (N_39707,N_37456,N_36144);
xnor U39708 (N_39708,N_35188,N_36786);
xor U39709 (N_39709,N_35235,N_37272);
nor U39710 (N_39710,N_36780,N_37415);
and U39711 (N_39711,N_36652,N_35555);
xnor U39712 (N_39712,N_36330,N_36156);
or U39713 (N_39713,N_35734,N_36423);
nor U39714 (N_39714,N_35127,N_36393);
xor U39715 (N_39715,N_35986,N_36508);
nor U39716 (N_39716,N_35861,N_35175);
xnor U39717 (N_39717,N_35049,N_36706);
nand U39718 (N_39718,N_36414,N_36528);
nand U39719 (N_39719,N_35311,N_36258);
nand U39720 (N_39720,N_35445,N_35969);
nor U39721 (N_39721,N_36001,N_35587);
or U39722 (N_39722,N_35120,N_35840);
xnor U39723 (N_39723,N_36549,N_35593);
nor U39724 (N_39724,N_36912,N_35657);
nand U39725 (N_39725,N_36035,N_36267);
and U39726 (N_39726,N_36607,N_36293);
xor U39727 (N_39727,N_36783,N_36175);
and U39728 (N_39728,N_37349,N_36104);
xor U39729 (N_39729,N_37110,N_37164);
nor U39730 (N_39730,N_36209,N_37169);
or U39731 (N_39731,N_36319,N_35754);
xnor U39732 (N_39732,N_35301,N_36391);
nand U39733 (N_39733,N_36147,N_36304);
nor U39734 (N_39734,N_35396,N_36906);
and U39735 (N_39735,N_35136,N_36852);
and U39736 (N_39736,N_35877,N_35446);
nand U39737 (N_39737,N_36667,N_35541);
nand U39738 (N_39738,N_35041,N_36858);
nand U39739 (N_39739,N_36564,N_36558);
and U39740 (N_39740,N_37266,N_36615);
nor U39741 (N_39741,N_35634,N_35409);
and U39742 (N_39742,N_36096,N_35220);
nand U39743 (N_39743,N_36231,N_36650);
nand U39744 (N_39744,N_36667,N_37457);
nand U39745 (N_39745,N_36928,N_36243);
or U39746 (N_39746,N_37230,N_36238);
nor U39747 (N_39747,N_37130,N_35752);
nand U39748 (N_39748,N_37276,N_35685);
xnor U39749 (N_39749,N_36543,N_36069);
xor U39750 (N_39750,N_35349,N_37382);
or U39751 (N_39751,N_35773,N_36213);
nand U39752 (N_39752,N_36794,N_37037);
xnor U39753 (N_39753,N_37384,N_35958);
nor U39754 (N_39754,N_37263,N_36449);
and U39755 (N_39755,N_35759,N_36712);
xnor U39756 (N_39756,N_35884,N_36305);
nand U39757 (N_39757,N_36245,N_36141);
nand U39758 (N_39758,N_36259,N_35473);
nand U39759 (N_39759,N_35831,N_35008);
nand U39760 (N_39760,N_35867,N_35305);
or U39761 (N_39761,N_37329,N_35296);
or U39762 (N_39762,N_36508,N_35125);
xor U39763 (N_39763,N_37458,N_35571);
or U39764 (N_39764,N_35595,N_35638);
nor U39765 (N_39765,N_37309,N_37359);
nand U39766 (N_39766,N_36820,N_35398);
and U39767 (N_39767,N_35791,N_36042);
nor U39768 (N_39768,N_36008,N_35610);
nor U39769 (N_39769,N_37327,N_35500);
nand U39770 (N_39770,N_36870,N_36397);
nand U39771 (N_39771,N_35511,N_36834);
nand U39772 (N_39772,N_35581,N_36637);
nand U39773 (N_39773,N_35946,N_37090);
xor U39774 (N_39774,N_37050,N_37014);
xnor U39775 (N_39775,N_36704,N_35531);
or U39776 (N_39776,N_36454,N_36396);
xnor U39777 (N_39777,N_35898,N_35961);
nand U39778 (N_39778,N_36839,N_35363);
nand U39779 (N_39779,N_36832,N_37068);
nor U39780 (N_39780,N_35303,N_35450);
nor U39781 (N_39781,N_37475,N_37066);
nand U39782 (N_39782,N_35589,N_36720);
and U39783 (N_39783,N_35731,N_35958);
or U39784 (N_39784,N_35524,N_36262);
nand U39785 (N_39785,N_36205,N_36498);
and U39786 (N_39786,N_37296,N_36144);
xnor U39787 (N_39787,N_36164,N_36509);
or U39788 (N_39788,N_36800,N_36934);
nor U39789 (N_39789,N_35251,N_35004);
nor U39790 (N_39790,N_36887,N_36299);
and U39791 (N_39791,N_35540,N_36717);
xnor U39792 (N_39792,N_36114,N_35370);
nor U39793 (N_39793,N_36235,N_36938);
or U39794 (N_39794,N_36196,N_36244);
and U39795 (N_39795,N_37168,N_35838);
nand U39796 (N_39796,N_35562,N_35760);
nor U39797 (N_39797,N_35053,N_35249);
xor U39798 (N_39798,N_36443,N_37041);
nor U39799 (N_39799,N_37293,N_36449);
xnor U39800 (N_39800,N_35527,N_36230);
or U39801 (N_39801,N_37207,N_36906);
and U39802 (N_39802,N_36054,N_37290);
xor U39803 (N_39803,N_37314,N_36531);
nand U39804 (N_39804,N_36427,N_36336);
nand U39805 (N_39805,N_36779,N_35637);
xnor U39806 (N_39806,N_35629,N_35393);
nor U39807 (N_39807,N_37386,N_36368);
or U39808 (N_39808,N_35621,N_36671);
and U39809 (N_39809,N_37089,N_36657);
nand U39810 (N_39810,N_35009,N_35006);
or U39811 (N_39811,N_36140,N_36879);
nand U39812 (N_39812,N_35104,N_36600);
and U39813 (N_39813,N_36413,N_37493);
and U39814 (N_39814,N_35337,N_36964);
nand U39815 (N_39815,N_35947,N_35294);
nor U39816 (N_39816,N_35064,N_37043);
nand U39817 (N_39817,N_35962,N_36263);
nand U39818 (N_39818,N_36110,N_36013);
or U39819 (N_39819,N_35404,N_36715);
and U39820 (N_39820,N_36966,N_37292);
nand U39821 (N_39821,N_37320,N_37374);
xnor U39822 (N_39822,N_36809,N_35836);
xnor U39823 (N_39823,N_35978,N_35245);
or U39824 (N_39824,N_35205,N_37326);
or U39825 (N_39825,N_35559,N_35429);
xor U39826 (N_39826,N_35120,N_36233);
and U39827 (N_39827,N_36489,N_36088);
xor U39828 (N_39828,N_36147,N_35732);
nand U39829 (N_39829,N_35463,N_36745);
nand U39830 (N_39830,N_37140,N_36612);
and U39831 (N_39831,N_35386,N_35062);
and U39832 (N_39832,N_35473,N_35681);
or U39833 (N_39833,N_36071,N_37475);
nand U39834 (N_39834,N_36921,N_36308);
nand U39835 (N_39835,N_35524,N_37388);
or U39836 (N_39836,N_37189,N_36432);
and U39837 (N_39837,N_36680,N_35003);
nand U39838 (N_39838,N_36271,N_35017);
xor U39839 (N_39839,N_36436,N_36581);
xor U39840 (N_39840,N_35118,N_37191);
nand U39841 (N_39841,N_36050,N_36529);
and U39842 (N_39842,N_36349,N_37448);
nand U39843 (N_39843,N_35329,N_36641);
nand U39844 (N_39844,N_37494,N_36969);
nand U39845 (N_39845,N_35793,N_37139);
or U39846 (N_39846,N_37012,N_36458);
nand U39847 (N_39847,N_37229,N_35616);
or U39848 (N_39848,N_35461,N_35982);
or U39849 (N_39849,N_36505,N_35328);
nand U39850 (N_39850,N_37369,N_37302);
nor U39851 (N_39851,N_37332,N_37013);
nand U39852 (N_39852,N_36325,N_36002);
nand U39853 (N_39853,N_35775,N_36902);
and U39854 (N_39854,N_36920,N_35842);
nor U39855 (N_39855,N_36810,N_35509);
and U39856 (N_39856,N_35774,N_37369);
or U39857 (N_39857,N_37264,N_37390);
xor U39858 (N_39858,N_35580,N_35172);
nor U39859 (N_39859,N_35981,N_35830);
or U39860 (N_39860,N_36273,N_37262);
and U39861 (N_39861,N_35282,N_36928);
or U39862 (N_39862,N_35526,N_36526);
nand U39863 (N_39863,N_37127,N_35257);
and U39864 (N_39864,N_35803,N_36819);
and U39865 (N_39865,N_35114,N_35695);
nor U39866 (N_39866,N_36902,N_36261);
nand U39867 (N_39867,N_36429,N_35467);
or U39868 (N_39868,N_36064,N_35136);
or U39869 (N_39869,N_37314,N_36711);
or U39870 (N_39870,N_35352,N_35468);
nor U39871 (N_39871,N_35564,N_35083);
or U39872 (N_39872,N_36203,N_36071);
and U39873 (N_39873,N_35028,N_37428);
xor U39874 (N_39874,N_37090,N_37334);
nand U39875 (N_39875,N_36914,N_36324);
nor U39876 (N_39876,N_35546,N_35313);
or U39877 (N_39877,N_36132,N_35485);
or U39878 (N_39878,N_35573,N_35774);
and U39879 (N_39879,N_36701,N_36550);
xnor U39880 (N_39880,N_37076,N_35172);
or U39881 (N_39881,N_35825,N_37225);
or U39882 (N_39882,N_36784,N_36977);
nor U39883 (N_39883,N_36100,N_36969);
nor U39884 (N_39884,N_35699,N_35738);
and U39885 (N_39885,N_36622,N_35443);
nand U39886 (N_39886,N_37372,N_36264);
or U39887 (N_39887,N_36233,N_37152);
nor U39888 (N_39888,N_37081,N_36134);
xor U39889 (N_39889,N_36443,N_36347);
nor U39890 (N_39890,N_35816,N_37115);
or U39891 (N_39891,N_36929,N_37358);
xor U39892 (N_39892,N_37060,N_36684);
nand U39893 (N_39893,N_35581,N_37207);
nor U39894 (N_39894,N_36491,N_35988);
xor U39895 (N_39895,N_35039,N_36870);
nand U39896 (N_39896,N_36622,N_35291);
xor U39897 (N_39897,N_36751,N_37019);
and U39898 (N_39898,N_35111,N_36822);
xnor U39899 (N_39899,N_36988,N_35996);
nor U39900 (N_39900,N_37309,N_37173);
or U39901 (N_39901,N_37453,N_36861);
or U39902 (N_39902,N_37450,N_35710);
or U39903 (N_39903,N_36898,N_35813);
or U39904 (N_39904,N_36762,N_36361);
xnor U39905 (N_39905,N_35875,N_37056);
xnor U39906 (N_39906,N_36400,N_37446);
nand U39907 (N_39907,N_36795,N_35508);
or U39908 (N_39908,N_35386,N_36007);
nor U39909 (N_39909,N_35314,N_36391);
nand U39910 (N_39910,N_37039,N_35609);
or U39911 (N_39911,N_35402,N_35835);
xor U39912 (N_39912,N_36093,N_36294);
and U39913 (N_39913,N_36633,N_35269);
nand U39914 (N_39914,N_37084,N_36252);
nor U39915 (N_39915,N_36653,N_35617);
or U39916 (N_39916,N_35509,N_35777);
xnor U39917 (N_39917,N_36742,N_35339);
nand U39918 (N_39918,N_36235,N_36919);
and U39919 (N_39919,N_36558,N_35057);
nor U39920 (N_39920,N_36447,N_35259);
nor U39921 (N_39921,N_36536,N_36659);
xor U39922 (N_39922,N_35060,N_36609);
or U39923 (N_39923,N_35281,N_35886);
and U39924 (N_39924,N_35531,N_36273);
nand U39925 (N_39925,N_36874,N_36145);
xnor U39926 (N_39926,N_36725,N_35402);
nand U39927 (N_39927,N_36529,N_37290);
nor U39928 (N_39928,N_37173,N_37452);
xnor U39929 (N_39929,N_35645,N_36517);
and U39930 (N_39930,N_35373,N_35227);
nor U39931 (N_39931,N_36314,N_37342);
xor U39932 (N_39932,N_36213,N_36888);
xor U39933 (N_39933,N_36880,N_35425);
xnor U39934 (N_39934,N_35871,N_37293);
xnor U39935 (N_39935,N_36526,N_35777);
and U39936 (N_39936,N_37372,N_35544);
nor U39937 (N_39937,N_37299,N_35842);
or U39938 (N_39938,N_35623,N_35174);
and U39939 (N_39939,N_36329,N_36999);
nand U39940 (N_39940,N_36620,N_36013);
nand U39941 (N_39941,N_36186,N_36083);
nor U39942 (N_39942,N_35646,N_35826);
and U39943 (N_39943,N_36065,N_37080);
nand U39944 (N_39944,N_35007,N_35746);
and U39945 (N_39945,N_35008,N_35841);
nand U39946 (N_39946,N_36072,N_37413);
nor U39947 (N_39947,N_36854,N_36222);
nor U39948 (N_39948,N_35244,N_36525);
and U39949 (N_39949,N_37005,N_36298);
and U39950 (N_39950,N_37009,N_36645);
nand U39951 (N_39951,N_35961,N_36525);
nor U39952 (N_39952,N_35208,N_36665);
nand U39953 (N_39953,N_35707,N_37264);
or U39954 (N_39954,N_35869,N_37367);
and U39955 (N_39955,N_35101,N_35627);
or U39956 (N_39956,N_36097,N_35242);
nor U39957 (N_39957,N_35358,N_35054);
and U39958 (N_39958,N_36095,N_36407);
and U39959 (N_39959,N_36197,N_37458);
or U39960 (N_39960,N_36758,N_36316);
xor U39961 (N_39961,N_36364,N_35512);
nor U39962 (N_39962,N_35456,N_35127);
xnor U39963 (N_39963,N_36790,N_37068);
nand U39964 (N_39964,N_35339,N_37449);
nor U39965 (N_39965,N_37118,N_35462);
or U39966 (N_39966,N_37292,N_37443);
and U39967 (N_39967,N_36196,N_35173);
nand U39968 (N_39968,N_36310,N_36057);
or U39969 (N_39969,N_35034,N_36393);
xnor U39970 (N_39970,N_35209,N_36279);
and U39971 (N_39971,N_35572,N_36680);
and U39972 (N_39972,N_35354,N_35901);
nand U39973 (N_39973,N_36438,N_37353);
xor U39974 (N_39974,N_36882,N_36116);
and U39975 (N_39975,N_35967,N_37018);
nand U39976 (N_39976,N_37380,N_35493);
xnor U39977 (N_39977,N_37216,N_37043);
or U39978 (N_39978,N_37002,N_35302);
or U39979 (N_39979,N_36870,N_35531);
and U39980 (N_39980,N_36911,N_36344);
nor U39981 (N_39981,N_35902,N_36019);
xnor U39982 (N_39982,N_35236,N_36478);
or U39983 (N_39983,N_35505,N_36928);
and U39984 (N_39984,N_37190,N_37298);
and U39985 (N_39985,N_36358,N_36045);
nand U39986 (N_39986,N_35580,N_36533);
or U39987 (N_39987,N_37184,N_36426);
nor U39988 (N_39988,N_37433,N_37488);
or U39989 (N_39989,N_35839,N_35832);
nand U39990 (N_39990,N_36375,N_35211);
and U39991 (N_39991,N_36763,N_37256);
nor U39992 (N_39992,N_37234,N_37262);
and U39993 (N_39993,N_36039,N_35546);
nor U39994 (N_39994,N_35790,N_36993);
or U39995 (N_39995,N_37262,N_35430);
nor U39996 (N_39996,N_37093,N_35506);
nor U39997 (N_39997,N_35088,N_37130);
and U39998 (N_39998,N_36006,N_35213);
nor U39999 (N_39999,N_37025,N_35576);
xor U40000 (N_40000,N_38548,N_39160);
nand U40001 (N_40001,N_38248,N_38724);
xor U40002 (N_40002,N_39629,N_39761);
and U40003 (N_40003,N_37899,N_39607);
nor U40004 (N_40004,N_37586,N_38577);
xor U40005 (N_40005,N_37728,N_39108);
nand U40006 (N_40006,N_39102,N_38167);
xor U40007 (N_40007,N_38474,N_39058);
and U40008 (N_40008,N_39129,N_38351);
and U40009 (N_40009,N_38797,N_39801);
nand U40010 (N_40010,N_39766,N_39641);
nor U40011 (N_40011,N_38314,N_38671);
and U40012 (N_40012,N_38128,N_39551);
nor U40013 (N_40013,N_38303,N_38876);
or U40014 (N_40014,N_38052,N_38542);
xor U40015 (N_40015,N_39323,N_38963);
nor U40016 (N_40016,N_39856,N_38983);
nor U40017 (N_40017,N_39670,N_39458);
nand U40018 (N_40018,N_39914,N_37657);
and U40019 (N_40019,N_38296,N_38782);
nand U40020 (N_40020,N_37753,N_38118);
nor U40021 (N_40021,N_37833,N_38895);
and U40022 (N_40022,N_39567,N_37844);
nor U40023 (N_40023,N_38747,N_38282);
nor U40024 (N_40024,N_37952,N_39524);
xor U40025 (N_40025,N_39703,N_38780);
nand U40026 (N_40026,N_37894,N_38074);
or U40027 (N_40027,N_38423,N_38250);
xor U40028 (N_40028,N_39752,N_38631);
or U40029 (N_40029,N_38568,N_37737);
nor U40030 (N_40030,N_39133,N_38674);
and U40031 (N_40031,N_37523,N_38907);
xor U40032 (N_40032,N_37856,N_38764);
or U40033 (N_40033,N_39146,N_37722);
nand U40034 (N_40034,N_38810,N_39587);
and U40035 (N_40035,N_39943,N_39953);
or U40036 (N_40036,N_39344,N_38094);
and U40037 (N_40037,N_37669,N_38710);
or U40038 (N_40038,N_38697,N_39842);
xor U40039 (N_40039,N_38525,N_37725);
or U40040 (N_40040,N_37605,N_39969);
and U40041 (N_40041,N_38902,N_38309);
and U40042 (N_40042,N_39408,N_38765);
xor U40043 (N_40043,N_38925,N_37947);
xnor U40044 (N_40044,N_39515,N_37759);
nor U40045 (N_40045,N_39184,N_38318);
nand U40046 (N_40046,N_38905,N_38723);
xor U40047 (N_40047,N_38329,N_38239);
xnor U40048 (N_40048,N_39310,N_39814);
nand U40049 (N_40049,N_39224,N_39230);
and U40050 (N_40050,N_39002,N_38863);
nand U40051 (N_40051,N_38316,N_38550);
and U40052 (N_40052,N_39837,N_37627);
nor U40053 (N_40053,N_37865,N_39902);
nand U40054 (N_40054,N_38744,N_39859);
nand U40055 (N_40055,N_39823,N_38587);
and U40056 (N_40056,N_37784,N_37817);
or U40057 (N_40057,N_39552,N_37573);
nand U40058 (N_40058,N_39417,N_39403);
xnor U40059 (N_40059,N_39598,N_39988);
or U40060 (N_40060,N_39983,N_39213);
or U40061 (N_40061,N_38682,N_38315);
nor U40062 (N_40062,N_39589,N_37561);
and U40063 (N_40063,N_38051,N_38013);
nor U40064 (N_40064,N_39937,N_38236);
nor U40065 (N_40065,N_38801,N_38645);
or U40066 (N_40066,N_39525,N_39857);
nor U40067 (N_40067,N_37576,N_39669);
and U40068 (N_40068,N_37542,N_39092);
nand U40069 (N_40069,N_37765,N_39929);
nor U40070 (N_40070,N_39410,N_38124);
and U40071 (N_40071,N_38803,N_39152);
or U40072 (N_40072,N_39570,N_39256);
nand U40073 (N_40073,N_39155,N_38394);
or U40074 (N_40074,N_39235,N_39991);
and U40075 (N_40075,N_38770,N_38814);
nand U40076 (N_40076,N_39592,N_37895);
nand U40077 (N_40077,N_37930,N_38169);
xor U40078 (N_40078,N_38121,N_38180);
and U40079 (N_40079,N_39986,N_39557);
nand U40080 (N_40080,N_38312,N_39899);
or U40081 (N_40081,N_37734,N_39107);
xnor U40082 (N_40082,N_38229,N_37896);
and U40083 (N_40083,N_38655,N_39646);
xnor U40084 (N_40084,N_38161,N_39012);
nand U40085 (N_40085,N_39807,N_39486);
xor U40086 (N_40086,N_38428,N_37874);
nor U40087 (N_40087,N_38210,N_37937);
and U40088 (N_40088,N_39556,N_37668);
nor U40089 (N_40089,N_37604,N_37697);
xnor U40090 (N_40090,N_38806,N_37860);
or U40091 (N_40091,N_38235,N_38761);
or U40092 (N_40092,N_37956,N_37559);
nand U40093 (N_40093,N_39100,N_38625);
and U40094 (N_40094,N_39069,N_38232);
nand U40095 (N_40095,N_38756,N_37934);
or U40096 (N_40096,N_38462,N_37908);
or U40097 (N_40097,N_37763,N_38883);
and U40098 (N_40098,N_37564,N_39363);
nor U40099 (N_40099,N_38630,N_38050);
or U40100 (N_40100,N_39671,N_39478);
and U40101 (N_40101,N_37821,N_39490);
or U40102 (N_40102,N_39689,N_38352);
or U40103 (N_40103,N_39895,N_39076);
nand U40104 (N_40104,N_37507,N_37731);
xor U40105 (N_40105,N_37782,N_39581);
and U40106 (N_40106,N_38284,N_37970);
xor U40107 (N_40107,N_39151,N_37553);
and U40108 (N_40108,N_38993,N_38442);
nand U40109 (N_40109,N_37500,N_38451);
nand U40110 (N_40110,N_38837,N_39026);
nor U40111 (N_40111,N_39767,N_37904);
xor U40112 (N_40112,N_37900,N_38096);
nor U40113 (N_40113,N_38502,N_39055);
nor U40114 (N_40114,N_38258,N_37506);
and U40115 (N_40115,N_39302,N_38768);
xnor U40116 (N_40116,N_39339,N_37743);
nand U40117 (N_40117,N_38215,N_38585);
nor U40118 (N_40118,N_39804,N_38716);
nand U40119 (N_40119,N_38865,N_39800);
nand U40120 (N_40120,N_39354,N_39295);
nor U40121 (N_40121,N_39196,N_39723);
nand U40122 (N_40122,N_38365,N_39217);
xnor U40123 (N_40123,N_37603,N_39554);
nand U40124 (N_40124,N_37827,N_37946);
and U40125 (N_40125,N_38748,N_39566);
nor U40126 (N_40126,N_39187,N_38699);
or U40127 (N_40127,N_38592,N_39178);
nor U40128 (N_40128,N_39585,N_37995);
nor U40129 (N_40129,N_39872,N_38861);
nand U40130 (N_40130,N_38078,N_38030);
nand U40131 (N_40131,N_38958,N_38226);
nor U40132 (N_40132,N_39430,N_38727);
nand U40133 (N_40133,N_38054,N_38927);
or U40134 (N_40134,N_39433,N_37518);
or U40135 (N_40135,N_39584,N_39483);
nor U40136 (N_40136,N_38327,N_39582);
or U40137 (N_40137,N_37878,N_39623);
and U40138 (N_40138,N_37813,N_39046);
xor U40139 (N_40139,N_38940,N_38978);
and U40140 (N_40140,N_39432,N_37846);
and U40141 (N_40141,N_39032,N_39536);
and U40142 (N_40142,N_38920,N_38904);
and U40143 (N_40143,N_39678,N_38387);
xnor U40144 (N_40144,N_37715,N_39167);
and U40145 (N_40145,N_37872,N_39518);
nand U40146 (N_40146,N_39538,N_37544);
or U40147 (N_40147,N_39132,N_39396);
xor U40148 (N_40148,N_38741,N_37509);
xor U40149 (N_40149,N_37512,N_37723);
nand U40150 (N_40150,N_38141,N_38785);
xor U40151 (N_40151,N_39086,N_38760);
and U40152 (N_40152,N_39604,N_38243);
nand U40153 (N_40153,N_39361,N_37873);
nor U40154 (N_40154,N_39850,N_39494);
nand U40155 (N_40155,N_37704,N_39867);
or U40156 (N_40156,N_39711,N_38794);
nand U40157 (N_40157,N_39739,N_38807);
or U40158 (N_40158,N_39650,N_39870);
nand U40159 (N_40159,N_39916,N_39630);
nor U40160 (N_40160,N_39830,N_38642);
nand U40161 (N_40161,N_38117,N_37563);
or U40162 (N_40162,N_39647,N_38531);
nor U40163 (N_40163,N_38179,N_38755);
or U40164 (N_40164,N_39989,N_37767);
and U40165 (N_40165,N_38804,N_39139);
nor U40166 (N_40166,N_39891,N_39159);
xnor U40167 (N_40167,N_38076,N_39972);
nand U40168 (N_40168,N_38835,N_37768);
xor U40169 (N_40169,N_37525,N_38916);
and U40170 (N_40170,N_38516,N_37979);
nand U40171 (N_40171,N_38811,N_38650);
and U40172 (N_40172,N_37640,N_38223);
and U40173 (N_40173,N_38767,N_37510);
nor U40174 (N_40174,N_37732,N_39634);
xor U40175 (N_40175,N_39318,N_39821);
or U40176 (N_40176,N_39828,N_37965);
and U40177 (N_40177,N_37670,N_37770);
xor U40178 (N_40178,N_37959,N_39048);
nand U40179 (N_40179,N_39110,N_39239);
or U40180 (N_40180,N_39071,N_38511);
nand U40181 (N_40181,N_38687,N_37783);
xnor U40182 (N_40182,N_37879,N_39528);
nor U40183 (N_40183,N_38073,N_38844);
nand U40184 (N_40184,N_37968,N_38789);
xor U40185 (N_40185,N_38304,N_37868);
or U40186 (N_40186,N_39666,N_38523);
and U40187 (N_40187,N_39913,N_37578);
and U40188 (N_40188,N_37769,N_39450);
or U40189 (N_40189,N_39643,N_38483);
xor U40190 (N_40190,N_37819,N_38026);
or U40191 (N_40191,N_39005,N_38264);
nor U40192 (N_40192,N_39811,N_37752);
nand U40193 (N_40193,N_39887,N_38133);
and U40194 (N_40194,N_38400,N_39019);
and U40195 (N_40195,N_38341,N_37651);
nand U40196 (N_40196,N_38045,N_37633);
nand U40197 (N_40197,N_39281,N_38530);
nand U40198 (N_40198,N_37630,N_39590);
nand U40199 (N_40199,N_39888,N_39338);
xor U40200 (N_40200,N_38698,N_37793);
xnor U40201 (N_40201,N_37624,N_38553);
and U40202 (N_40202,N_38230,N_39721);
nor U40203 (N_40203,N_39818,N_38822);
nand U40204 (N_40204,N_39963,N_39639);
and U40205 (N_40205,N_37880,N_38184);
xnor U40206 (N_40206,N_38043,N_39699);
or U40207 (N_40207,N_37637,N_38111);
xnor U40208 (N_40208,N_38846,N_38153);
and U40209 (N_40209,N_37949,N_38443);
xnor U40210 (N_40210,N_37677,N_37698);
nand U40211 (N_40211,N_38166,N_39860);
nand U40212 (N_40212,N_39083,N_38473);
xnor U40213 (N_40213,N_39014,N_37811);
nand U40214 (N_40214,N_37625,N_39506);
and U40215 (N_40215,N_37683,N_39077);
nor U40216 (N_40216,N_38065,N_38424);
nor U40217 (N_40217,N_39796,N_39935);
and U40218 (N_40218,N_37859,N_39880);
xor U40219 (N_40219,N_38673,N_38055);
xor U40220 (N_40220,N_39980,N_38881);
and U40221 (N_40221,N_39246,N_38859);
nand U40222 (N_40222,N_38999,N_39288);
or U40223 (N_40223,N_39717,N_38206);
xor U40224 (N_40224,N_39145,N_39087);
nand U40225 (N_40225,N_37917,N_38418);
nand U40226 (N_40226,N_39037,N_39328);
and U40227 (N_40227,N_39770,N_39497);
xor U40228 (N_40228,N_39103,N_39233);
and U40229 (N_40229,N_38211,N_38393);
nor U40230 (N_40230,N_37925,N_38934);
and U40231 (N_40231,N_38634,N_38829);
and U40232 (N_40232,N_38189,N_39874);
xnor U40233 (N_40233,N_37528,N_37555);
or U40234 (N_40234,N_38549,N_39960);
or U40235 (N_40235,N_37809,N_38827);
nand U40236 (N_40236,N_37511,N_39783);
xor U40237 (N_40237,N_37659,N_39855);
and U40238 (N_40238,N_38856,N_38980);
nor U40239 (N_40239,N_39840,N_37781);
or U40240 (N_40240,N_38132,N_39222);
nand U40241 (N_40241,N_38265,N_38664);
nor U40242 (N_40242,N_39693,N_39117);
and U40243 (N_40243,N_38368,N_39097);
nand U40244 (N_40244,N_38746,N_38208);
or U40245 (N_40245,N_38173,N_39393);
xor U40246 (N_40246,N_37584,N_39179);
nand U40247 (N_40247,N_39386,N_39392);
and U40248 (N_40248,N_38320,N_38136);
nor U40249 (N_40249,N_38330,N_39215);
or U40250 (N_40250,N_39329,N_38696);
and U40251 (N_40251,N_39010,N_39586);
xnor U40252 (N_40252,N_39269,N_37745);
nand U40253 (N_40253,N_39404,N_38449);
and U40254 (N_40254,N_39907,N_39084);
nor U40255 (N_40255,N_38751,N_38070);
or U40256 (N_40256,N_38602,N_39695);
or U40257 (N_40257,N_37596,N_39081);
nand U40258 (N_40258,N_37923,N_39072);
nor U40259 (N_40259,N_39280,N_38938);
or U40260 (N_40260,N_37772,N_38667);
or U40261 (N_40261,N_37988,N_39161);
nor U40262 (N_40262,N_39866,N_38564);
nand U40263 (N_40263,N_38384,N_37733);
and U40264 (N_40264,N_38291,N_38757);
or U40265 (N_40265,N_39290,N_38476);
or U40266 (N_40266,N_37853,N_38385);
nor U40267 (N_40267,N_39782,N_39143);
xor U40268 (N_40268,N_39291,N_39172);
or U40269 (N_40269,N_38665,N_39777);
and U40270 (N_40270,N_39426,N_38788);
nor U40271 (N_40271,N_38053,N_38909);
nand U40272 (N_40272,N_38573,N_37685);
or U40273 (N_40273,N_38565,N_39407);
xnor U40274 (N_40274,N_38508,N_39798);
xor U40275 (N_40275,N_38851,N_38274);
nand U40276 (N_40276,N_38972,N_38008);
nor U40277 (N_40277,N_38061,N_39027);
and U40278 (N_40278,N_38112,N_38877);
nor U40279 (N_40279,N_39692,N_38843);
nor U40280 (N_40280,N_39833,N_39119);
nand U40281 (N_40281,N_38535,N_39775);
and U40282 (N_40282,N_38583,N_38499);
nand U40283 (N_40283,N_38164,N_38558);
xnor U40284 (N_40284,N_38363,N_39658);
nor U40285 (N_40285,N_39806,N_39876);
nor U40286 (N_40286,N_38255,N_38644);
or U40287 (N_40287,N_38029,N_39169);
xnor U40288 (N_40288,N_39511,N_39398);
or U40289 (N_40289,N_38155,N_37565);
or U40290 (N_40290,N_39419,N_38935);
and U40291 (N_40291,N_37619,N_39894);
or U40292 (N_40292,N_37829,N_38669);
nand U40293 (N_40293,N_38335,N_38694);
or U40294 (N_40294,N_39292,N_37903);
or U40295 (N_40295,N_38900,N_39208);
xor U40296 (N_40296,N_39690,N_39517);
nor U40297 (N_40297,N_38151,N_39476);
and U40298 (N_40298,N_37777,N_39349);
nor U40299 (N_40299,N_38556,N_38171);
nand U40300 (N_40300,N_38850,N_38256);
or U40301 (N_40301,N_39237,N_38779);
xnor U40302 (N_40302,N_38188,N_38840);
nor U40303 (N_40303,N_37588,N_37678);
or U40304 (N_40304,N_38928,N_38467);
or U40305 (N_40305,N_39025,N_38620);
and U40306 (N_40306,N_39464,N_38869);
or U40307 (N_40307,N_37701,N_39482);
nor U40308 (N_40308,N_38596,N_38639);
and U40309 (N_40309,N_39079,N_38659);
and U40310 (N_40310,N_38396,N_39682);
or U40311 (N_40311,N_39347,N_37647);
and U40312 (N_40312,N_39765,N_39687);
and U40313 (N_40313,N_38410,N_39051);
or U40314 (N_40314,N_38638,N_38679);
or U40315 (N_40315,N_38539,N_38591);
xnor U40316 (N_40316,N_39000,N_39659);
and U40317 (N_40317,N_37757,N_37626);
xnor U40318 (N_40318,N_37980,N_39204);
or U40319 (N_40319,N_38464,N_37594);
or U40320 (N_40320,N_38745,N_38098);
or U40321 (N_40321,N_39619,N_37870);
nor U40322 (N_40322,N_39321,N_37775);
nand U40323 (N_40323,N_37893,N_38600);
xor U40324 (N_40324,N_39173,N_38580);
and U40325 (N_40325,N_38060,N_39244);
nand U40326 (N_40326,N_38652,N_39945);
and U40327 (N_40327,N_38191,N_38279);
and U40328 (N_40328,N_38138,N_38971);
nor U40329 (N_40329,N_38903,N_39950);
or U40330 (N_40330,N_39406,N_39958);
or U40331 (N_40331,N_37961,N_38010);
nor U40332 (N_40332,N_38246,N_39507);
and U40333 (N_40333,N_37915,N_38005);
xor U40334 (N_40334,N_38217,N_38297);
or U40335 (N_40335,N_37803,N_39553);
or U40336 (N_40336,N_38995,N_39418);
nor U40337 (N_40337,N_38513,N_38685);
nand U40338 (N_40338,N_38914,N_37762);
and U40339 (N_40339,N_39846,N_39622);
and U40340 (N_40340,N_38609,N_38933);
xnor U40341 (N_40341,N_38581,N_38036);
and U40342 (N_40342,N_38285,N_39078);
nand U40343 (N_40343,N_38676,N_39095);
nand U40344 (N_40344,N_39547,N_37650);
xor U40345 (N_40345,N_38276,N_39477);
xor U40346 (N_40346,N_39951,N_37838);
or U40347 (N_40347,N_38287,N_39413);
or U40348 (N_40348,N_38129,N_39707);
nand U40349 (N_40349,N_39588,N_39024);
or U40350 (N_40350,N_39085,N_39401);
or U40351 (N_40351,N_37839,N_38491);
nor U40352 (N_40352,N_39467,N_39137);
or U40353 (N_40353,N_38377,N_39597);
nor U40354 (N_40354,N_39356,N_37850);
nand U40355 (N_40355,N_38527,N_39253);
xnor U40356 (N_40356,N_38786,N_38456);
and U40357 (N_40357,N_37587,N_38383);
xor U40358 (N_40358,N_39886,N_39999);
xor U40359 (N_40359,N_39740,N_38080);
nor U40360 (N_40360,N_38946,N_38186);
or U40361 (N_40361,N_39123,N_39434);
or U40362 (N_40362,N_38438,N_38796);
nor U40363 (N_40363,N_38607,N_37902);
nor U40364 (N_40364,N_39315,N_39255);
xnor U40365 (N_40365,N_38866,N_39611);
nor U40366 (N_40366,N_39308,N_38254);
xor U40367 (N_40367,N_38924,N_38706);
and U40368 (N_40368,N_38730,N_39499);
nand U40369 (N_40369,N_37661,N_37533);
or U40370 (N_40370,N_38360,N_38231);
nor U40371 (N_40371,N_39189,N_38379);
xnor U40372 (N_40372,N_37545,N_39059);
or U40373 (N_40373,N_39153,N_38367);
and U40374 (N_40374,N_39257,N_39994);
xor U40375 (N_40375,N_37711,N_37913);
nor U40376 (N_40376,N_39959,N_39883);
and U40377 (N_40377,N_38003,N_37720);
and U40378 (N_40378,N_39966,N_38889);
xor U40379 (N_40379,N_39925,N_37522);
or U40380 (N_40380,N_39109,N_38241);
nor U40381 (N_40381,N_39710,N_39150);
and U40382 (N_40382,N_39358,N_37599);
nor U40383 (N_40383,N_39089,N_39555);
or U40384 (N_40384,N_38551,N_38649);
nand U40385 (N_40385,N_37749,N_39003);
or U40386 (N_40386,N_39036,N_39734);
nand U40387 (N_40387,N_39580,N_38280);
nor U40388 (N_40388,N_38987,N_39520);
and U40389 (N_40389,N_39532,N_38197);
or U40390 (N_40390,N_38336,N_39294);
or U40391 (N_40391,N_39421,N_39331);
nor U40392 (N_40392,N_38259,N_38989);
nand U40393 (N_40393,N_38729,N_37729);
nand U40394 (N_40394,N_38345,N_39908);
or U40395 (N_40395,N_37779,N_38482);
nor U40396 (N_40396,N_38743,N_38774);
or U40397 (N_40397,N_38720,N_39794);
xor U40398 (N_40398,N_39571,N_39340);
or U40399 (N_40399,N_39140,N_39709);
xor U40400 (N_40400,N_38378,N_38375);
or U40401 (N_40401,N_37571,N_38000);
nand U40402 (N_40402,N_38959,N_39175);
nand U40403 (N_40403,N_37572,N_39183);
or U40404 (N_40404,N_38068,N_38358);
xnor U40405 (N_40405,N_37682,N_39015);
nor U40406 (N_40406,N_39044,N_37546);
nand U40407 (N_40407,N_37609,N_39971);
and U40408 (N_40408,N_38718,N_39093);
nor U40409 (N_40409,N_38064,N_39277);
or U40410 (N_40410,N_37503,N_38781);
xor U40411 (N_40411,N_39260,N_39405);
xnor U40412 (N_40412,N_39017,N_38465);
and U40413 (N_40413,N_38018,N_39768);
nor U40414 (N_40414,N_39545,N_39758);
nand U40415 (N_40415,N_38728,N_39063);
xor U40416 (N_40416,N_37556,N_38588);
xor U40417 (N_40417,N_37514,N_37841);
and U40418 (N_40418,N_37534,N_37504);
and U40419 (N_40419,N_38487,N_38269);
or U40420 (N_40420,N_37928,N_39911);
and U40421 (N_40421,N_39884,N_39023);
nand U40422 (N_40422,N_37944,N_39849);
nand U40423 (N_40423,N_39529,N_38610);
nand U40424 (N_40424,N_38249,N_37938);
xor U40425 (N_40425,N_37675,N_39445);
or U40426 (N_40426,N_39147,N_39936);
nand U40427 (N_40427,N_38648,N_38478);
and U40428 (N_40428,N_39763,N_38614);
or U40429 (N_40429,N_39459,N_39961);
nor U40430 (N_40430,N_38988,N_39090);
nand U40431 (N_40431,N_39439,N_37884);
nor U40432 (N_40432,N_37616,N_39177);
nor U40433 (N_40433,N_38198,N_38931);
and U40434 (N_40434,N_37665,N_38126);
xor U40435 (N_40435,N_38823,N_38149);
xnor U40436 (N_40436,N_39737,N_38566);
xor U40437 (N_40437,N_38102,N_38470);
or U40438 (N_40438,N_39211,N_37939);
or U40439 (N_40439,N_38216,N_37797);
or U40440 (N_40440,N_39534,N_38700);
and U40441 (N_40441,N_38095,N_37877);
and U40442 (N_40442,N_37920,N_38828);
xor U40443 (N_40443,N_38058,N_38702);
nand U40444 (N_40444,N_39377,N_39653);
xor U40445 (N_40445,N_37750,N_38137);
nor U40446 (N_40446,N_39028,N_37897);
nand U40447 (N_40447,N_39327,N_39676);
xnor U40448 (N_40448,N_39144,N_37790);
nand U40449 (N_40449,N_39033,N_39648);
or U40450 (N_40450,N_38825,N_38113);
xor U40451 (N_40451,N_39301,N_38617);
nor U40452 (N_40452,N_38471,N_39381);
xnor U40453 (N_40453,N_38268,N_38656);
and U40454 (N_40454,N_38571,N_37613);
or U40455 (N_40455,N_37606,N_38627);
nand U40456 (N_40456,N_38307,N_37551);
nor U40457 (N_40457,N_39157,N_38873);
xor U40458 (N_40458,N_37667,N_37787);
or U40459 (N_40459,N_37948,N_38956);
nand U40460 (N_40460,N_38047,N_38082);
xor U40461 (N_40461,N_38506,N_38463);
xor U40462 (N_40462,N_37910,N_39602);
and U40463 (N_40463,N_39885,N_37964);
and U40464 (N_40464,N_38611,N_38389);
nor U40465 (N_40465,N_38594,N_38019);
xnor U40466 (N_40466,N_38042,N_37941);
or U40467 (N_40467,N_37796,N_37892);
xor U40468 (N_40468,N_39496,N_38323);
nand U40469 (N_40469,N_37806,N_38975);
nand U40470 (N_40470,N_38218,N_39922);
xnor U40471 (N_40471,N_39781,N_38805);
and U40472 (N_40472,N_37644,N_39127);
nor U40473 (N_40473,N_38874,N_37807);
and U40474 (N_40474,N_39463,N_39053);
and U40475 (N_40475,N_38012,N_38401);
xor U40476 (N_40476,N_39427,N_38209);
nor U40477 (N_40477,N_38460,N_39596);
nor U40478 (N_40478,N_38172,N_37608);
nand U40479 (N_40479,N_39409,N_38622);
nand U40480 (N_40480,N_38301,N_38875);
nand U40481 (N_40481,N_39829,N_38497);
xor U40482 (N_40482,N_37997,N_39192);
nor U40483 (N_40483,N_38613,N_39871);
nor U40484 (N_40484,N_39188,N_38651);
or U40485 (N_40485,N_39389,N_39601);
nand U40486 (N_40486,N_37932,N_38635);
or U40487 (N_40487,N_39877,N_38922);
or U40488 (N_40488,N_38954,N_37852);
and U40489 (N_40489,N_37642,N_39696);
and U40490 (N_40490,N_37834,N_39190);
xor U40491 (N_40491,N_37718,N_38343);
or U40492 (N_40492,N_38714,N_37631);
and U40493 (N_40493,N_38306,N_37719);
nand U40494 (N_40494,N_38289,N_38108);
nor U40495 (N_40495,N_37971,N_38426);
xor U40496 (N_40496,N_39411,N_39722);
xor U40497 (N_40497,N_38021,N_38295);
and U40498 (N_40498,N_38599,N_39334);
or U40499 (N_40499,N_38347,N_37516);
nor U40500 (N_40500,N_39423,N_39785);
xor U40501 (N_40501,N_38890,N_39271);
and U40502 (N_40502,N_38177,N_39289);
nor U40503 (N_40503,N_39198,N_39742);
nand U40504 (N_40504,N_37526,N_39106);
or U40505 (N_40505,N_38769,N_39614);
or U40506 (N_40506,N_39539,N_39706);
xor U40507 (N_40507,N_38708,N_38257);
nand U40508 (N_40508,N_38022,N_39034);
and U40509 (N_40509,N_38662,N_39638);
and U40510 (N_40510,N_38455,N_38390);
or U40511 (N_40511,N_37891,N_38116);
nand U40512 (N_40512,N_39337,N_38842);
or U40513 (N_40513,N_38386,N_39284);
or U40514 (N_40514,N_39508,N_38948);
xor U40515 (N_40515,N_39893,N_38813);
or U40516 (N_40516,N_38572,N_39826);
xor U40517 (N_40517,N_38193,N_39612);
nand U40518 (N_40518,N_39131,N_38270);
nand U40519 (N_40519,N_39724,N_39569);
nand U40520 (N_40520,N_39975,N_38808);
nor U40521 (N_40521,N_39632,N_38071);
nor U40522 (N_40522,N_37687,N_38143);
nand U40523 (N_40523,N_38783,N_38641);
xor U40524 (N_40524,N_37854,N_39812);
nor U40525 (N_40525,N_39957,N_38691);
or U40526 (N_40526,N_37581,N_39454);
or U40527 (N_40527,N_37808,N_38083);
and U40528 (N_40528,N_39248,N_39784);
and U40529 (N_40529,N_38417,N_39435);
nor U40530 (N_40530,N_38452,N_39514);
or U40531 (N_40531,N_38448,N_38404);
or U40532 (N_40532,N_38382,N_39955);
nand U40533 (N_40533,N_39573,N_38009);
nand U40534 (N_40534,N_37875,N_39346);
xnor U40535 (N_40535,N_37695,N_37935);
nor U40536 (N_40536,N_38242,N_39174);
xor U40537 (N_40537,N_39018,N_38409);
nand U40538 (N_40538,N_38292,N_38308);
xnor U40539 (N_40539,N_38795,N_38546);
xor U40540 (N_40540,N_38195,N_38445);
nand U40541 (N_40541,N_37774,N_39191);
nor U40542 (N_40542,N_38115,N_38559);
nand U40543 (N_40543,N_39898,N_39485);
nand U40544 (N_40544,N_37812,N_39942);
nand U40545 (N_40545,N_39306,N_39940);
nor U40546 (N_40546,N_39049,N_38252);
xnor U40547 (N_40547,N_38359,N_37802);
nand U40548 (N_40548,N_39762,N_38266);
nand U40549 (N_40549,N_38949,N_38561);
xnor U40550 (N_40550,N_39162,N_38500);
and U40551 (N_40551,N_37820,N_37869);
and U40552 (N_40552,N_38758,N_39073);
or U40553 (N_40553,N_38271,N_37635);
nand U40554 (N_40554,N_38072,N_37689);
nor U40555 (N_40555,N_37638,N_38518);
nor U40556 (N_40556,N_38833,N_38888);
or U40557 (N_40557,N_39652,N_38666);
and U40558 (N_40558,N_38589,N_38845);
nand U40559 (N_40559,N_37748,N_38926);
xor U40560 (N_40560,N_37990,N_38552);
or U40561 (N_40561,N_39273,N_38974);
xor U40562 (N_40562,N_39941,N_39373);
xor U40563 (N_40563,N_38737,N_39789);
nor U40564 (N_40564,N_37996,N_38961);
nor U40565 (N_40565,N_39440,N_37562);
and U40566 (N_40566,N_39992,N_38369);
xor U40567 (N_40567,N_39757,N_38668);
or U40568 (N_40568,N_38294,N_38120);
nor U40569 (N_40569,N_38985,N_39399);
xor U40570 (N_40570,N_39933,N_37933);
and U40571 (N_40571,N_38187,N_39954);
and U40572 (N_40572,N_38753,N_38221);
or U40573 (N_40573,N_38704,N_37520);
nor U40574 (N_40574,N_39105,N_38317);
and U40575 (N_40575,N_39088,N_38468);
xnor U40576 (N_40576,N_37529,N_38885);
nor U40577 (N_40577,N_38640,N_39663);
nand U40578 (N_40578,N_38380,N_38355);
nand U40579 (N_40579,N_37842,N_38604);
and U40580 (N_40580,N_39926,N_39543);
nand U40581 (N_40581,N_39265,N_39825);
and U40582 (N_40582,N_38407,N_38233);
or U40583 (N_40583,N_39997,N_39564);
nand U40584 (N_40584,N_39965,N_39351);
and U40585 (N_40585,N_38624,N_38520);
xnor U40586 (N_40586,N_39640,N_38929);
or U40587 (N_40587,N_38033,N_38688);
xnor U40588 (N_40588,N_38575,N_37680);
nor U40589 (N_40589,N_39832,N_37824);
xor U40590 (N_40590,N_37740,N_38181);
nor U40591 (N_40591,N_38134,N_37674);
or U40592 (N_40592,N_38953,N_38089);
nand U40593 (N_40593,N_39822,N_37862);
xor U40594 (N_40594,N_39008,N_38984);
nor U40595 (N_40595,N_38251,N_37771);
xnor U40596 (N_40596,N_38776,N_39621);
nor U40597 (N_40597,N_37831,N_38273);
or U40598 (N_40598,N_38964,N_38841);
nor U40599 (N_40599,N_39387,N_37577);
xnor U40600 (N_40600,N_39625,N_38402);
nand U40601 (N_40601,N_39094,N_38338);
or U40602 (N_40602,N_38263,N_39939);
nor U40603 (N_40603,N_37539,N_39229);
xor U40604 (N_40604,N_38541,N_38192);
or U40605 (N_40605,N_38154,N_38411);
nand U40606 (N_40606,N_37672,N_39062);
nor U40607 (N_40607,N_37825,N_38201);
or U40608 (N_40608,N_38534,N_38416);
xor U40609 (N_40609,N_39091,N_39182);
xnor U40610 (N_40610,N_38576,N_39158);
xor U40611 (N_40611,N_39384,N_38821);
nor U40612 (N_40612,N_38415,N_38701);
and U40613 (N_40613,N_38826,N_39357);
xnor U40614 (N_40614,N_37958,N_39715);
nor U40615 (N_40615,N_37521,N_39156);
or U40616 (N_40616,N_38447,N_38420);
or U40617 (N_40617,N_37798,N_37681);
and U40618 (N_40618,N_37830,N_39043);
xnor U40619 (N_40619,N_37658,N_38777);
xnor U40620 (N_40620,N_38340,N_39274);
or U40621 (N_40621,N_38434,N_37712);
xnor U40622 (N_40622,N_39863,N_38678);
xor U40623 (N_40623,N_38880,N_39165);
nor U40624 (N_40624,N_39769,N_38945);
xor U40625 (N_40625,N_38537,N_39719);
nand U40626 (N_40626,N_38125,N_39572);
and U40627 (N_40627,N_37866,N_39541);
xnor U40628 (N_40628,N_38152,N_38749);
or U40629 (N_40629,N_38286,N_39952);
and U40630 (N_40630,N_38818,N_39600);
xnor U40631 (N_40631,N_38654,N_37795);
nand U40632 (N_40632,N_39824,N_39755);
or U40633 (N_40633,N_39512,N_38658);
nor U40634 (N_40634,N_39293,N_39270);
and U40635 (N_40635,N_37876,N_39258);
and U40636 (N_40636,N_38996,N_38574);
xor U40637 (N_40637,N_39462,N_37814);
nor U40638 (N_40638,N_38897,N_39847);
and U40639 (N_40639,N_38979,N_38101);
xor U40640 (N_40640,N_39704,N_39491);
nor U40641 (N_40641,N_38224,N_38006);
or U40642 (N_40642,N_38220,N_38435);
nor U40643 (N_40643,N_38707,N_39793);
xor U40644 (N_40644,N_39168,N_38834);
and U40645 (N_40645,N_39021,N_38034);
nand U40646 (N_40646,N_38114,N_39115);
nand U40647 (N_40647,N_39488,N_39243);
or U40648 (N_40648,N_38762,N_37989);
and U40649 (N_40649,N_39903,N_38371);
nand U40650 (N_40650,N_39054,N_39052);
or U40651 (N_40651,N_37531,N_39714);
xnor U40652 (N_40652,N_39948,N_38519);
or U40653 (N_40653,N_38908,N_37554);
nand U40654 (N_40654,N_39546,N_38163);
nor U40655 (N_40655,N_39057,N_39299);
nand U40656 (N_40656,N_38353,N_38578);
nor U40657 (N_40657,N_37991,N_39428);
and U40658 (N_40658,N_37690,N_39200);
nor U40659 (N_40659,N_39390,N_39918);
nor U40660 (N_40660,N_38947,N_39668);
or U40661 (N_40661,N_38991,N_37984);
nor U40662 (N_40662,N_38792,N_39684);
nor U40663 (N_40663,N_39031,N_39838);
and U40664 (N_40664,N_37909,N_39045);
nand U40665 (N_40665,N_39111,N_38864);
and U40666 (N_40666,N_39424,N_39447);
nor U40667 (N_40667,N_39901,N_37943);
and U40668 (N_40668,N_39449,N_38469);
nand U40669 (N_40669,N_39041,N_38529);
nand U40670 (N_40670,N_37972,N_37721);
or U40671 (N_40671,N_38496,N_38941);
nand U40672 (N_40672,N_37632,N_39324);
and U40673 (N_40673,N_37560,N_38579);
and U40674 (N_40674,N_38349,N_37810);
xnor U40675 (N_40675,N_39786,N_37593);
nand U40676 (N_40676,N_37579,N_38182);
and U40677 (N_40677,N_37598,N_37566);
or U40678 (N_40678,N_39309,N_37582);
or U40679 (N_40679,N_39697,N_39510);
xor U40680 (N_40680,N_38509,N_39070);
or U40681 (N_40681,N_37963,N_39774);
or U40682 (N_40682,N_38998,N_38326);
xnor U40683 (N_40683,N_39627,N_39320);
nor U40684 (N_40684,N_38398,N_38538);
and U40685 (N_40685,N_39996,N_38075);
and U40686 (N_40686,N_39773,N_39171);
xor U40687 (N_40687,N_39210,N_38512);
or U40688 (N_40688,N_39559,N_38293);
or U40689 (N_40689,N_38791,N_37634);
and U40690 (N_40690,N_39415,N_38812);
nand U40691 (N_40691,N_39262,N_39688);
nand U40692 (N_40692,N_39912,N_38918);
or U40693 (N_40693,N_38809,N_39836);
xor U40694 (N_40694,N_39104,N_37864);
nor U40695 (N_40695,N_38868,N_37709);
or U40696 (N_40696,N_39082,N_38362);
nor U40697 (N_40697,N_38479,N_37648);
xnor U40698 (N_40698,N_39383,N_37998);
or U40699 (N_40699,N_38772,N_37548);
xnor U40700 (N_40700,N_37921,N_39312);
nor U40701 (N_40701,N_38107,N_37622);
nand U40702 (N_40702,N_39820,N_39125);
xnor U40703 (N_40703,N_37601,N_39397);
or U40704 (N_40704,N_39148,N_39206);
nand U40705 (N_40705,N_39560,N_39674);
xor U40706 (N_40706,N_39974,N_39114);
and U40707 (N_40707,N_39446,N_37501);
nor U40708 (N_40708,N_39353,N_39928);
xor U40709 (N_40709,N_39562,N_38399);
and U40710 (N_40710,N_37886,N_37716);
and U40711 (N_40711,N_39287,N_39927);
or U40712 (N_40712,N_39743,N_39416);
nor U40713 (N_40713,N_37639,N_39713);
nand U40714 (N_40714,N_38740,N_39465);
and U40715 (N_40715,N_39875,N_39685);
and U40716 (N_40716,N_39261,N_38099);
and U40717 (N_40717,N_39799,N_37726);
nor U40718 (N_40718,N_39780,N_39466);
and U40719 (N_40719,N_38454,N_38917);
nand U40720 (N_40720,N_37773,N_39635);
and U40721 (N_40721,N_39307,N_38689);
xnor U40722 (N_40722,N_39591,N_38647);
nor U40723 (N_40723,N_39068,N_39050);
nor U40724 (N_40724,N_38077,N_38742);
nand U40725 (N_40725,N_38930,N_38160);
and U40726 (N_40726,N_39577,N_37791);
nand U40727 (N_40727,N_39128,N_38441);
nand U40728 (N_40728,N_39726,N_38049);
and U40729 (N_40729,N_39201,N_39220);
and U40730 (N_40730,N_38450,N_38608);
or U40731 (N_40731,N_39788,N_37652);
or U40732 (N_40732,N_37758,N_37666);
nor U40733 (N_40733,N_38750,N_39851);
nand U40734 (N_40734,N_37867,N_38046);
nand U40735 (N_40735,N_38272,N_37730);
nor U40736 (N_40736,N_39352,N_38838);
nand U40737 (N_40737,N_37558,N_38563);
and U40738 (N_40738,N_37914,N_39660);
nand U40739 (N_40739,N_38175,N_39915);
or U40740 (N_40740,N_39135,N_38703);
nor U40741 (N_40741,N_39495,N_38752);
nand U40742 (N_40742,N_37957,N_39296);
or U40743 (N_40743,N_37643,N_38225);
and U40744 (N_40744,N_38488,N_38555);
nor U40745 (N_40745,N_37889,N_38898);
nand U40746 (N_40746,N_37614,N_39608);
nor U40747 (N_40747,N_38227,N_38731);
nor U40748 (N_40748,N_38247,N_39376);
nor U40749 (N_40749,N_39437,N_38016);
nand U40750 (N_40750,N_39325,N_38732);
xnor U40751 (N_40751,N_38200,N_38521);
nor U40752 (N_40752,N_39134,N_38693);
and U40753 (N_40753,N_38194,N_39892);
and U40754 (N_40754,N_38901,N_38376);
and U40755 (N_40755,N_39332,N_39480);
and U40756 (N_40756,N_38148,N_37585);
and U40757 (N_40757,N_38734,N_37960);
nor U40758 (N_40758,N_38093,N_39620);
and U40759 (N_40759,N_39195,N_37699);
nor U40760 (N_40760,N_37540,N_39964);
or U40761 (N_40761,N_38867,N_38886);
nor U40762 (N_40762,N_38754,N_38997);
nand U40763 (N_40763,N_39575,N_39456);
or U40764 (N_40764,N_38505,N_38739);
nand U40765 (N_40765,N_37705,N_37926);
and U40766 (N_40766,N_38122,N_37918);
or U40767 (N_40767,N_38331,N_38636);
and U40768 (N_40768,N_38853,N_39748);
nor U40769 (N_40769,N_37794,N_39400);
nand U40770 (N_40770,N_39574,N_39197);
and U40771 (N_40771,N_39234,N_37663);
nand U40772 (N_40772,N_39568,N_39987);
and U40773 (N_40773,N_39720,N_39815);
nor U40774 (N_40774,N_39618,N_38800);
xnor U40775 (N_40775,N_39637,N_38854);
nand U40776 (N_40776,N_39412,N_39730);
or U40777 (N_40777,N_39792,N_38203);
nand U40778 (N_40778,N_39205,N_39848);
xnor U40779 (N_40779,N_38207,N_37617);
nor U40780 (N_40780,N_39380,N_39313);
nand U40781 (N_40781,N_37848,N_39683);
and U40782 (N_40782,N_38477,N_39022);
nor U40783 (N_40783,N_38643,N_37591);
nand U40784 (N_40784,N_38283,N_38784);
or U40785 (N_40785,N_37756,N_38490);
xnor U40786 (N_40786,N_39651,N_39728);
nor U40787 (N_40787,N_39662,N_39225);
xnor U40788 (N_40788,N_39531,N_38976);
nand U40789 (N_40789,N_39917,N_37535);
or U40790 (N_40790,N_37741,N_39747);
or U40791 (N_40791,N_38213,N_37645);
and U40792 (N_40792,N_39113,N_37919);
xor U40793 (N_40793,N_38878,N_37655);
or U40794 (N_40794,N_37708,N_39579);
nor U40795 (N_40795,N_39667,N_39921);
and U40796 (N_40796,N_38965,N_37927);
nand U40797 (N_40797,N_37955,N_38891);
xnor U40798 (N_40798,N_38830,N_37881);
nor U40799 (N_40799,N_38457,N_38267);
nor U40800 (N_40800,N_38504,N_38446);
and U40801 (N_40801,N_39194,N_37818);
or U40802 (N_40802,N_39616,N_37656);
xor U40803 (N_40803,N_39075,N_39231);
nor U40804 (N_40804,N_37929,N_38238);
and U40805 (N_40805,N_38489,N_38858);
nor U40806 (N_40806,N_37822,N_37536);
xor U40807 (N_40807,N_38484,N_39549);
or U40808 (N_40808,N_37676,N_38119);
nand U40809 (N_40809,N_39968,N_37799);
nand U40810 (N_40810,N_39909,N_38960);
or U40811 (N_40811,N_38593,N_37696);
and U40812 (N_40812,N_39605,N_37727);
or U40813 (N_40813,N_38709,N_39594);
nor U40814 (N_40814,N_38582,N_38726);
or U40815 (N_40815,N_39443,N_38884);
or U40816 (N_40816,N_38144,N_39138);
nand U40817 (N_40817,N_37924,N_39448);
nand U40818 (N_40818,N_39042,N_37912);
nor U40819 (N_40819,N_37832,N_38260);
or U40820 (N_40820,N_38882,N_39655);
nor U40821 (N_40821,N_37863,N_38025);
and U40822 (N_40822,N_38715,N_37849);
nand U40823 (N_40823,N_39493,N_37836);
nand U40824 (N_40824,N_39956,N_39263);
nor U40825 (N_40825,N_39947,N_37583);
nor U40826 (N_40826,N_38472,N_38942);
nor U40827 (N_40827,N_39333,N_38816);
xor U40828 (N_40828,N_38894,N_39121);
and U40829 (N_40829,N_38969,N_38951);
or U40830 (N_40830,N_38632,N_38526);
nand U40831 (N_40831,N_39944,N_37538);
nand U40832 (N_40832,N_38855,N_38421);
and U40833 (N_40833,N_39249,N_39548);
and U40834 (N_40834,N_39267,N_38039);
and U40835 (N_40835,N_39735,N_39489);
and U40836 (N_40836,N_38494,N_39932);
and U40837 (N_40837,N_39778,N_37974);
and U40838 (N_40838,N_39523,N_38439);
nor U40839 (N_40839,N_38437,N_39672);
nand U40840 (N_40840,N_39475,N_38717);
xor U40841 (N_40841,N_38560,N_39881);
nand U40842 (N_40842,N_37845,N_39897);
and U40843 (N_40843,N_37703,N_37788);
and U40844 (N_40844,N_38766,N_37700);
xor U40845 (N_40845,N_38820,N_38319);
xor U40846 (N_40846,N_38104,N_39420);
xor U40847 (N_40847,N_38852,N_37597);
nor U40848 (N_40848,N_39372,N_37575);
nand U40849 (N_40849,N_38196,N_39595);
and U40850 (N_40850,N_38228,N_39065);
or U40851 (N_40851,N_39732,N_39371);
nor U40852 (N_40852,N_37761,N_37592);
nor U40853 (N_40853,N_38562,N_39878);
or U40854 (N_40854,N_39232,N_38950);
or U40855 (N_40855,N_38615,N_38584);
or U40856 (N_40856,N_39976,N_37888);
nor U40857 (N_40857,N_38381,N_39216);
xor U40858 (N_40858,N_38943,N_38899);
xnor U40859 (N_40859,N_38857,N_39006);
and U40860 (N_40860,N_37589,N_37786);
and U40861 (N_40861,N_37567,N_38150);
nand U40862 (N_40862,N_37710,N_39455);
and U40863 (N_40863,N_39680,N_38536);
xnor U40864 (N_40864,N_39348,N_38162);
xor U40865 (N_40865,N_37549,N_39985);
or U40866 (N_40866,N_38084,N_37541);
nand U40867 (N_40867,N_39995,N_39492);
nand U40868 (N_40868,N_39136,N_38603);
nor U40869 (N_40869,N_37898,N_38939);
nand U40870 (N_40870,N_38059,N_37954);
nor U40871 (N_40871,N_39852,N_38966);
xor U40872 (N_40872,N_38533,N_39609);
xnor U40873 (N_40873,N_39831,N_39862);
and U40874 (N_40874,N_39429,N_39444);
nor U40875 (N_40875,N_39864,N_39727);
and U40876 (N_40876,N_37754,N_38165);
or U40877 (N_40877,N_39973,N_37901);
nand U40878 (N_40878,N_37611,N_39516);
nor U40879 (N_40879,N_38277,N_38431);
xor U40880 (N_40880,N_39934,N_39064);
xnor U40881 (N_40881,N_37532,N_38344);
nand U40882 (N_40882,N_39981,N_38567);
nand U40883 (N_40883,N_39481,N_37664);
xor U40884 (N_40884,N_38031,N_38787);
nand U40885 (N_40885,N_39750,N_37981);
nor U40886 (N_40886,N_38007,N_38515);
and U40887 (N_40887,N_39099,N_39414);
xnor U40888 (N_40888,N_37612,N_38994);
nand U40889 (N_40889,N_38313,N_37950);
nand U40890 (N_40890,N_39460,N_38763);
or U40891 (N_40891,N_39001,N_37580);
or U40892 (N_40892,N_38024,N_37621);
or U40893 (N_40893,N_38973,N_38066);
or U40894 (N_40894,N_39664,N_38507);
nor U40895 (N_40895,N_39473,N_38370);
and U40896 (N_40896,N_39038,N_39236);
xor U40897 (N_40897,N_38621,N_38305);
and U40898 (N_40898,N_38253,N_38722);
nand U40899 (N_40899,N_38035,N_37887);
nor U40900 (N_40900,N_37693,N_39819);
and U40901 (N_40901,N_37969,N_38332);
or U40902 (N_40902,N_39606,N_39238);
or U40903 (N_40903,N_39369,N_39362);
and U40904 (N_40904,N_39441,N_38015);
and U40905 (N_40905,N_39438,N_39753);
xnor U40906 (N_40906,N_39754,N_39470);
or U40907 (N_40907,N_38879,N_39242);
xnor U40908 (N_40908,N_38595,N_38480);
nor U40909 (N_40909,N_37684,N_37840);
nand U40910 (N_40910,N_39181,N_39827);
or U40911 (N_40911,N_39154,N_37978);
nand U40912 (N_40912,N_38159,N_38105);
nor U40913 (N_40913,N_38214,N_38919);
nand U40914 (N_40914,N_38372,N_39268);
nand U40915 (N_40915,N_38261,N_39779);
nand U40916 (N_40916,N_39350,N_37976);
or U40917 (N_40917,N_38183,N_38028);
xnor U40918 (N_40918,N_39080,N_38146);
and U40919 (N_40919,N_39869,N_39661);
or U40920 (N_40920,N_39163,N_38130);
nand U40921 (N_40921,N_38913,N_38660);
and U40922 (N_40922,N_38815,N_37543);
and U40923 (N_40923,N_39422,N_37828);
and U40924 (N_40924,N_39472,N_39803);
nor U40925 (N_40925,N_37861,N_38738);
nand U40926 (N_40926,N_39040,N_38131);
or U40927 (N_40927,N_38514,N_39451);
or U40928 (N_40928,N_37982,N_38799);
or U40929 (N_40929,N_39865,N_37744);
and U40930 (N_40930,N_37987,N_38346);
or U40931 (N_40931,N_39868,N_38366);
or U40932 (N_40932,N_39378,N_37953);
xnor U40933 (N_40933,N_38278,N_39379);
nand U40934 (N_40934,N_39771,N_38453);
and U40935 (N_40935,N_37911,N_39285);
and U40936 (N_40936,N_37962,N_37847);
or U40937 (N_40937,N_37568,N_39978);
nor U40938 (N_40938,N_39061,N_37519);
xnor U40939 (N_40939,N_38778,N_38350);
nand U40940 (N_40940,N_38736,N_38977);
xor U40941 (N_40941,N_39202,N_39617);
nor U40942 (N_40942,N_39385,N_39311);
xor U40943 (N_40943,N_37517,N_38037);
xor U40944 (N_40944,N_37671,N_37524);
xor U40945 (N_40945,N_38337,N_39141);
nor U40946 (N_40946,N_38027,N_37975);
or U40947 (N_40947,N_38466,N_39367);
or U40948 (N_40948,N_38923,N_37764);
and U40949 (N_40949,N_37590,N_38412);
xnor U40950 (N_40950,N_38554,N_39644);
nor U40951 (N_40951,N_38690,N_39341);
and U40952 (N_40952,N_38142,N_37985);
and U40953 (N_40953,N_39599,N_38001);
and U40954 (N_40954,N_39170,N_38110);
nor U40955 (N_40955,N_39214,N_37755);
and U40956 (N_40956,N_38719,N_39283);
xor U40957 (N_40957,N_38436,N_39558);
xor U40958 (N_40958,N_37906,N_39853);
nand U40959 (N_40959,N_39802,N_38802);
and U40960 (N_40960,N_39657,N_39905);
and U40961 (N_40961,N_39809,N_38906);
nand U40962 (N_40962,N_38616,N_39185);
nand U40963 (N_40963,N_38790,N_39264);
or U40964 (N_40964,N_38085,N_39919);
nor U40965 (N_40965,N_39776,N_38798);
and U40966 (N_40966,N_37835,N_38981);
and U40967 (N_40967,N_39839,N_38824);
or U40968 (N_40968,N_38836,N_38493);
xnor U40969 (N_40969,N_38677,N_39645);
and U40970 (N_40970,N_39904,N_39527);
xor U40971 (N_40971,N_37694,N_38176);
nor U40972 (N_40972,N_37785,N_38092);
and U40973 (N_40973,N_38081,N_39176);
and U40974 (N_40974,N_38601,N_39615);
nor U40975 (N_40975,N_38713,N_37505);
and U40976 (N_40976,N_39395,N_37738);
or U40977 (N_40977,N_37607,N_39011);
nor U40978 (N_40978,N_39364,N_39718);
nand U40979 (N_40979,N_37574,N_38896);
and U40980 (N_40980,N_38091,N_38299);
xor U40981 (N_40981,N_38819,N_38680);
nor U40982 (N_40982,N_38373,N_39442);
nor U40983 (N_40983,N_39513,N_39118);
or U40984 (N_40984,N_38444,N_39759);
nand U40985 (N_40985,N_39649,N_39039);
nand U40986 (N_40986,N_38915,N_39984);
or U40987 (N_40987,N_37973,N_39382);
nand U40988 (N_40988,N_38090,N_39879);
xnor U40989 (N_40989,N_38174,N_39537);
nand U40990 (N_40990,N_39474,N_39240);
and U40991 (N_40991,N_37792,N_38461);
nor U40992 (N_40992,N_38944,N_37736);
and U40993 (N_40993,N_39858,N_38429);
nor U40994 (N_40994,N_38532,N_39550);
nand U40995 (N_40995,N_39744,N_37931);
xor U40996 (N_40996,N_39368,N_38887);
xnor U40997 (N_40997,N_38721,N_38681);
and U40998 (N_40998,N_38413,N_39509);
and U40999 (N_40999,N_38205,N_39326);
or U41000 (N_41000,N_39336,N_39760);
xnor U41001 (N_41001,N_39841,N_39199);
nor U41002 (N_41002,N_39861,N_39526);
or U41003 (N_41003,N_38670,N_39751);
xor U41004 (N_41004,N_39479,N_39375);
nor U41005 (N_41005,N_39388,N_39681);
nand U41006 (N_41006,N_38495,N_38322);
and U41007 (N_41007,N_39316,N_39808);
nand U41008 (N_41008,N_38910,N_39613);
nand U41009 (N_41009,N_37885,N_39209);
and U41010 (N_41010,N_39164,N_38921);
and U41011 (N_41011,N_38324,N_38893);
or U41012 (N_41012,N_38023,N_38079);
and U41013 (N_41013,N_39533,N_37855);
nand U41014 (N_41014,N_39817,N_37776);
or U41015 (N_41015,N_39772,N_38485);
nor U41016 (N_41016,N_39193,N_38832);
and U41017 (N_41017,N_39503,N_37951);
nand U41018 (N_41018,N_38486,N_37780);
nand U41019 (N_41019,N_38653,N_39522);
or U41020 (N_41020,N_37826,N_39245);
nor U41021 (N_41021,N_39938,N_37602);
nand U41022 (N_41022,N_39716,N_39035);
nor U41023 (N_41023,N_38598,N_37649);
and U41024 (N_41024,N_38178,N_37570);
xor U41025 (N_41025,N_38540,N_39686);
xor U41026 (N_41026,N_38618,N_38771);
or U41027 (N_41027,N_37702,N_38127);
and U41028 (N_41028,N_37513,N_37550);
and U41029 (N_41029,N_39979,N_38067);
nand U41030 (N_41030,N_39923,N_37883);
and U41031 (N_41031,N_39746,N_39542);
and U41032 (N_41032,N_39247,N_39484);
nor U41033 (N_41033,N_37942,N_37994);
and U41034 (N_41034,N_39228,N_37751);
and U41035 (N_41035,N_38321,N_37618);
nor U41036 (N_41036,N_38962,N_38543);
and U41037 (N_41037,N_39431,N_39227);
nand U41038 (N_41038,N_39565,N_38501);
or U41039 (N_41039,N_38199,N_37805);
nor U41040 (N_41040,N_39665,N_39790);
or U41041 (N_41041,N_39067,N_39126);
nand U41042 (N_41042,N_38202,N_38310);
and U41043 (N_41043,N_38952,N_38892);
nand U41044 (N_41044,N_39345,N_38528);
nand U41045 (N_41045,N_38190,N_39251);
xor U41046 (N_41046,N_39845,N_38237);
nand U41047 (N_41047,N_39949,N_39370);
xnor U41048 (N_41048,N_37823,N_38395);
nor U41049 (N_41049,N_39004,N_37907);
xor U41050 (N_41050,N_38775,N_39203);
xor U41051 (N_41051,N_38204,N_39020);
or U41052 (N_41052,N_38522,N_38711);
nor U41053 (N_41053,N_39226,N_39835);
xnor U41054 (N_41054,N_37936,N_38057);
nor U41055 (N_41055,N_38356,N_37502);
nor U41056 (N_41056,N_39101,N_38735);
nand U41057 (N_41057,N_38361,N_38062);
nor U41058 (N_41058,N_39583,N_38406);
or U41059 (N_41059,N_38569,N_38968);
nand U41060 (N_41060,N_39130,N_37992);
nand U41061 (N_41061,N_39967,N_39124);
or U41062 (N_41062,N_37688,N_37746);
nand U41063 (N_41063,N_39745,N_39990);
and U41064 (N_41064,N_39593,N_39029);
nand U41065 (N_41065,N_39461,N_39679);
or U41066 (N_41066,N_38427,N_38302);
or U41067 (N_41067,N_39563,N_39452);
or U41068 (N_41068,N_38992,N_39365);
and U41069 (N_41069,N_39656,N_38860);
nor U41070 (N_41070,N_38219,N_38325);
or U41071 (N_41071,N_38440,N_38871);
or U41072 (N_41072,N_38262,N_37620);
or U41073 (N_41073,N_39394,N_37800);
and U41074 (N_41074,N_39166,N_39576);
nor U41075 (N_41075,N_38684,N_39610);
nand U41076 (N_41076,N_37857,N_39425);
and U41077 (N_41077,N_39254,N_39355);
xnor U41078 (N_41078,N_39504,N_38106);
xor U41079 (N_41079,N_39343,N_38623);
nand U41080 (N_41080,N_38425,N_39700);
nor U41081 (N_41081,N_38063,N_38657);
nand U41082 (N_41082,N_38357,N_37569);
xor U41083 (N_41083,N_37760,N_37653);
and U41084 (N_41084,N_38432,N_39813);
and U41085 (N_41085,N_39970,N_39795);
nand U41086 (N_41086,N_39675,N_39007);
xnor U41087 (N_41087,N_38069,N_39900);
xor U41088 (N_41088,N_38705,N_39906);
xnor U41089 (N_41089,N_39098,N_38123);
and U41090 (N_41090,N_39998,N_39319);
and U41091 (N_41091,N_39030,N_39276);
xor U41092 (N_41092,N_39931,N_38103);
xnor U41093 (N_41093,N_38032,N_37986);
or U41094 (N_41094,N_38619,N_39142);
nand U41095 (N_41095,N_39843,N_39009);
or U41096 (N_41096,N_38288,N_39741);
and U41097 (N_41097,N_39402,N_38597);
and U41098 (N_41098,N_39736,N_39854);
nor U41099 (N_41099,N_39920,N_39890);
nand U41100 (N_41100,N_39212,N_38109);
and U41101 (N_41101,N_37537,N_38403);
nor U41102 (N_41102,N_39149,N_38388);
nand U41103 (N_41103,N_39603,N_37691);
nor U41104 (N_41104,N_39122,N_38135);
and U41105 (N_41105,N_39816,N_38156);
and U41106 (N_41106,N_38245,N_37858);
and U41107 (N_41107,N_38339,N_38817);
nor U41108 (N_41108,N_38222,N_38663);
nor U41109 (N_41109,N_38870,N_39066);
and U41110 (N_41110,N_38524,N_38333);
and U41111 (N_41111,N_37967,N_39756);
and U41112 (N_41112,N_38170,N_38088);
and U41113 (N_41113,N_39300,N_39303);
or U41114 (N_41114,N_38695,N_37724);
nand U41115 (N_41115,N_39791,N_39374);
nor U41116 (N_41116,N_39930,N_38475);
nand U41117 (N_41117,N_39278,N_38281);
nand U41118 (N_41118,N_38545,N_39180);
and U41119 (N_41119,N_38848,N_39074);
or U41120 (N_41120,N_39335,N_39305);
or U41121 (N_41121,N_38041,N_38038);
nor U41122 (N_41122,N_39521,N_37692);
and U41123 (N_41123,N_38517,N_37707);
or U41124 (N_41124,N_39578,N_39342);
nand U41125 (N_41125,N_39501,N_37940);
or U41126 (N_41126,N_38002,N_38967);
or U41127 (N_41127,N_38298,N_38831);
nor U41128 (N_41128,N_38017,N_39738);
xnor U41129 (N_41129,N_37557,N_38328);
or U41130 (N_41130,N_39505,N_38646);
nand U41131 (N_41131,N_38586,N_39112);
and U41132 (N_41132,N_39628,N_38014);
and U41133 (N_41133,N_38422,N_37679);
xnor U41134 (N_41134,N_39834,N_38955);
nor U41135 (N_41135,N_37654,N_37646);
nor U41136 (N_41136,N_37983,N_39844);
nand U41137 (N_41137,N_39223,N_38364);
or U41138 (N_41138,N_38712,N_38004);
xor U41139 (N_41139,N_39540,N_37527);
xor U41140 (N_41140,N_39272,N_39882);
xor U41141 (N_41141,N_39502,N_38862);
and U41142 (N_41142,N_39787,N_39705);
or U41143 (N_41143,N_37660,N_38793);
or U41144 (N_41144,N_38957,N_38481);
nand U41145 (N_41145,N_39708,N_38839);
xor U41146 (N_41146,N_38408,N_38492);
or U41147 (N_41147,N_38145,N_38590);
nand U41148 (N_41148,N_38725,N_37515);
or U41149 (N_41149,N_39013,N_39360);
or U41150 (N_41150,N_39279,N_37530);
and U41151 (N_41151,N_38932,N_39391);
xnor U41152 (N_41152,N_39218,N_39297);
nor U41153 (N_41153,N_38459,N_38937);
xnor U41154 (N_41154,N_39749,N_38147);
xor U41155 (N_41155,N_38570,N_38936);
nor U41156 (N_41156,N_38414,N_38234);
xor U41157 (N_41157,N_39712,N_38290);
or U41158 (N_41158,N_39654,N_38733);
or U41159 (N_41159,N_38275,N_38311);
xnor U41160 (N_41160,N_37837,N_38849);
xnor U41161 (N_41161,N_38510,N_37686);
nand U41162 (N_41162,N_38672,N_37739);
nand U41163 (N_41163,N_39056,N_39436);
nor U41164 (N_41164,N_38168,N_39797);
nand U41165 (N_41165,N_38086,N_37610);
or U41166 (N_41166,N_38157,N_38354);
or U41167 (N_41167,N_38661,N_38629);
xor U41168 (N_41168,N_37890,N_38397);
or U41169 (N_41169,N_39633,N_37508);
and U41170 (N_41170,N_37977,N_37636);
or U41171 (N_41171,N_38606,N_39487);
nor U41172 (N_41172,N_38628,N_39221);
or U41173 (N_41173,N_37714,N_39810);
and U41174 (N_41174,N_39673,N_38097);
nor U41175 (N_41175,N_38100,N_38139);
or U41176 (N_41176,N_37778,N_37871);
and U41177 (N_41177,N_37816,N_38430);
xor U41178 (N_41178,N_38637,N_38686);
or U41179 (N_41179,N_38334,N_37742);
nor U41180 (N_41180,N_37641,N_38044);
nor U41181 (N_41181,N_39282,N_39366);
xor U41182 (N_41182,N_39453,N_38986);
nor U41183 (N_41183,N_39469,N_39698);
nor U41184 (N_41184,N_38020,N_38040);
or U41185 (N_41185,N_38185,N_39116);
and U41186 (N_41186,N_39498,N_38374);
and U41187 (N_41187,N_39471,N_38872);
xor U41188 (N_41188,N_37623,N_39642);
xnor U41189 (N_41189,N_38773,N_39266);
nor U41190 (N_41190,N_39286,N_37717);
and U41191 (N_41191,N_39544,N_37628);
nand U41192 (N_41192,N_39910,N_39314);
or U41193 (N_41193,N_37882,N_39060);
nand U41194 (N_41194,N_37966,N_38140);
nand U41195 (N_41195,N_38675,N_38503);
and U41196 (N_41196,N_39694,N_38544);
nand U41197 (N_41197,N_39701,N_37993);
xnor U41198 (N_41198,N_38633,N_37615);
nor U41199 (N_41199,N_39702,N_39873);
and U41200 (N_41200,N_39946,N_37547);
and U41201 (N_41201,N_39241,N_37851);
or U41202 (N_41202,N_39977,N_37673);
and U41203 (N_41203,N_38405,N_39993);
xor U41204 (N_41204,N_39457,N_38911);
nand U41205 (N_41205,N_39677,N_38348);
and U41206 (N_41206,N_38605,N_37789);
nand U41207 (N_41207,N_39016,N_37662);
or U41208 (N_41208,N_39924,N_39317);
nor U41209 (N_41209,N_39252,N_38087);
xnor U41210 (N_41210,N_39982,N_39207);
nor U41211 (N_41211,N_39304,N_39250);
xnor U41212 (N_41212,N_39275,N_39047);
and U41213 (N_41213,N_39219,N_37600);
xor U41214 (N_41214,N_39468,N_37922);
nand U41215 (N_41215,N_38547,N_38683);
nor U41216 (N_41216,N_39731,N_37804);
nand U41217 (N_41217,N_37801,N_38300);
nand U41218 (N_41218,N_38692,N_38626);
xor U41219 (N_41219,N_38212,N_38759);
nor U41220 (N_41220,N_38048,N_38240);
xor U41221 (N_41221,N_37706,N_39725);
or U41222 (N_41222,N_37843,N_39896);
nor U41223 (N_41223,N_38612,N_39298);
nor U41224 (N_41224,N_38912,N_37905);
or U41225 (N_41225,N_38433,N_39764);
nor U41226 (N_41226,N_38392,N_39500);
xor U41227 (N_41227,N_39561,N_39631);
nand U41228 (N_41228,N_38498,N_39636);
nand U41229 (N_41229,N_37713,N_38056);
or U41230 (N_41230,N_39624,N_38557);
nand U41231 (N_41231,N_38244,N_37766);
or U41232 (N_41232,N_39626,N_39322);
nand U41233 (N_41233,N_37945,N_39259);
nand U41234 (N_41234,N_37595,N_37552);
and U41235 (N_41235,N_39096,N_39359);
nand U41236 (N_41236,N_38847,N_38342);
or U41237 (N_41237,N_37735,N_39330);
nand U41238 (N_41238,N_39186,N_39691);
nor U41239 (N_41239,N_39535,N_38970);
nand U41240 (N_41240,N_39962,N_38990);
xnor U41241 (N_41241,N_37815,N_39805);
nor U41242 (N_41242,N_37999,N_38419);
nand U41243 (N_41243,N_38458,N_38011);
or U41244 (N_41244,N_38158,N_39889);
or U41245 (N_41245,N_38391,N_39519);
xor U41246 (N_41246,N_37916,N_38982);
and U41247 (N_41247,N_39120,N_39729);
or U41248 (N_41248,N_39530,N_37747);
and U41249 (N_41249,N_37629,N_39733);
nor U41250 (N_41250,N_39877,N_38305);
and U41251 (N_41251,N_38288,N_39729);
nand U41252 (N_41252,N_38176,N_39760);
nand U41253 (N_41253,N_39544,N_38588);
nand U41254 (N_41254,N_39288,N_38658);
nand U41255 (N_41255,N_39009,N_39611);
or U41256 (N_41256,N_38809,N_39318);
and U41257 (N_41257,N_37727,N_39530);
nand U41258 (N_41258,N_38487,N_39714);
or U41259 (N_41259,N_39595,N_38406);
and U41260 (N_41260,N_39531,N_38188);
or U41261 (N_41261,N_38462,N_39174);
and U41262 (N_41262,N_39467,N_38872);
nand U41263 (N_41263,N_39639,N_38592);
nand U41264 (N_41264,N_39174,N_37788);
xor U41265 (N_41265,N_39392,N_39183);
or U41266 (N_41266,N_38167,N_37616);
xor U41267 (N_41267,N_37799,N_39234);
or U41268 (N_41268,N_38283,N_38649);
xnor U41269 (N_41269,N_38740,N_38618);
or U41270 (N_41270,N_39817,N_38154);
nand U41271 (N_41271,N_37649,N_37923);
and U41272 (N_41272,N_37522,N_39778);
or U41273 (N_41273,N_38051,N_39115);
or U41274 (N_41274,N_38409,N_38935);
or U41275 (N_41275,N_37894,N_39099);
and U41276 (N_41276,N_39377,N_39262);
nand U41277 (N_41277,N_39804,N_38053);
xor U41278 (N_41278,N_37719,N_38850);
or U41279 (N_41279,N_37899,N_38521);
and U41280 (N_41280,N_37739,N_38026);
xnor U41281 (N_41281,N_38231,N_39610);
nand U41282 (N_41282,N_39196,N_39852);
xor U41283 (N_41283,N_39302,N_38816);
nand U41284 (N_41284,N_38792,N_37615);
and U41285 (N_41285,N_39802,N_39250);
xor U41286 (N_41286,N_38711,N_39638);
nor U41287 (N_41287,N_38414,N_38506);
or U41288 (N_41288,N_39974,N_39036);
nand U41289 (N_41289,N_38502,N_37618);
xnor U41290 (N_41290,N_38016,N_38254);
nand U41291 (N_41291,N_38096,N_38038);
nand U41292 (N_41292,N_37725,N_37680);
nand U41293 (N_41293,N_39020,N_38234);
or U41294 (N_41294,N_37900,N_39645);
xor U41295 (N_41295,N_37502,N_38374);
nor U41296 (N_41296,N_38366,N_38771);
or U41297 (N_41297,N_38293,N_39642);
and U41298 (N_41298,N_39259,N_38184);
or U41299 (N_41299,N_38076,N_37639);
and U41300 (N_41300,N_39364,N_39132);
and U41301 (N_41301,N_39698,N_37938);
and U41302 (N_41302,N_39572,N_39131);
or U41303 (N_41303,N_38678,N_39035);
xnor U41304 (N_41304,N_39578,N_38248);
or U41305 (N_41305,N_38134,N_39286);
or U41306 (N_41306,N_38608,N_39808);
xor U41307 (N_41307,N_37582,N_39982);
xnor U41308 (N_41308,N_39188,N_39442);
nor U41309 (N_41309,N_38777,N_37804);
or U41310 (N_41310,N_37526,N_37808);
xnor U41311 (N_41311,N_37747,N_38711);
xnor U41312 (N_41312,N_38697,N_39088);
xor U41313 (N_41313,N_39089,N_39331);
xor U41314 (N_41314,N_38043,N_38090);
nand U41315 (N_41315,N_39959,N_38574);
xor U41316 (N_41316,N_39027,N_38550);
or U41317 (N_41317,N_38603,N_38174);
nor U41318 (N_41318,N_39816,N_37551);
or U41319 (N_41319,N_38996,N_38224);
xnor U41320 (N_41320,N_39594,N_39225);
and U41321 (N_41321,N_38433,N_38676);
or U41322 (N_41322,N_38800,N_37738);
and U41323 (N_41323,N_37730,N_39714);
and U41324 (N_41324,N_39840,N_39417);
or U41325 (N_41325,N_37615,N_38593);
and U41326 (N_41326,N_39064,N_39398);
nor U41327 (N_41327,N_37733,N_39749);
and U41328 (N_41328,N_39008,N_38530);
nand U41329 (N_41329,N_39587,N_39894);
xnor U41330 (N_41330,N_38963,N_39533);
or U41331 (N_41331,N_39196,N_39823);
or U41332 (N_41332,N_37736,N_38752);
xor U41333 (N_41333,N_38936,N_38619);
xor U41334 (N_41334,N_37539,N_38630);
or U41335 (N_41335,N_39675,N_38472);
nand U41336 (N_41336,N_38057,N_38605);
and U41337 (N_41337,N_38251,N_39347);
and U41338 (N_41338,N_38263,N_38811);
xnor U41339 (N_41339,N_39474,N_37603);
xor U41340 (N_41340,N_39229,N_38461);
or U41341 (N_41341,N_37884,N_38085);
and U41342 (N_41342,N_39941,N_39755);
or U41343 (N_41343,N_38602,N_39599);
nor U41344 (N_41344,N_38192,N_37969);
and U41345 (N_41345,N_37737,N_38088);
or U41346 (N_41346,N_38191,N_37954);
nand U41347 (N_41347,N_38805,N_39998);
nand U41348 (N_41348,N_39498,N_39447);
nor U41349 (N_41349,N_37954,N_37698);
and U41350 (N_41350,N_39518,N_39966);
xor U41351 (N_41351,N_38117,N_39550);
or U41352 (N_41352,N_39411,N_37759);
and U41353 (N_41353,N_38648,N_37658);
or U41354 (N_41354,N_38278,N_37669);
nand U41355 (N_41355,N_39577,N_38645);
or U41356 (N_41356,N_39849,N_39002);
xnor U41357 (N_41357,N_38229,N_39455);
and U41358 (N_41358,N_39316,N_37845);
nand U41359 (N_41359,N_38306,N_39709);
xor U41360 (N_41360,N_38438,N_39341);
nand U41361 (N_41361,N_37906,N_38685);
nor U41362 (N_41362,N_38332,N_39712);
or U41363 (N_41363,N_39954,N_38075);
nand U41364 (N_41364,N_37886,N_39874);
nand U41365 (N_41365,N_39717,N_38427);
nand U41366 (N_41366,N_38918,N_39760);
xnor U41367 (N_41367,N_39139,N_39177);
nand U41368 (N_41368,N_38820,N_39574);
nor U41369 (N_41369,N_39139,N_38103);
nand U41370 (N_41370,N_39282,N_38060);
and U41371 (N_41371,N_38944,N_38217);
nor U41372 (N_41372,N_37912,N_39845);
and U41373 (N_41373,N_39014,N_37683);
xor U41374 (N_41374,N_38825,N_37623);
nand U41375 (N_41375,N_39896,N_39589);
nand U41376 (N_41376,N_39618,N_39370);
nor U41377 (N_41377,N_38365,N_38313);
nand U41378 (N_41378,N_37675,N_38984);
nor U41379 (N_41379,N_38171,N_38552);
and U41380 (N_41380,N_38964,N_38656);
or U41381 (N_41381,N_39490,N_39017);
nand U41382 (N_41382,N_38504,N_38168);
xnor U41383 (N_41383,N_38567,N_38620);
or U41384 (N_41384,N_37926,N_39601);
xor U41385 (N_41385,N_38717,N_39302);
or U41386 (N_41386,N_39917,N_37587);
or U41387 (N_41387,N_39329,N_37681);
and U41388 (N_41388,N_39981,N_39477);
or U41389 (N_41389,N_37842,N_39499);
xnor U41390 (N_41390,N_37711,N_39477);
xor U41391 (N_41391,N_39680,N_37914);
nor U41392 (N_41392,N_37694,N_38325);
or U41393 (N_41393,N_39863,N_39198);
nor U41394 (N_41394,N_39463,N_39414);
xnor U41395 (N_41395,N_37884,N_39500);
nor U41396 (N_41396,N_39509,N_38350);
xnor U41397 (N_41397,N_39792,N_39883);
xnor U41398 (N_41398,N_39639,N_39810);
xor U41399 (N_41399,N_38036,N_38629);
nand U41400 (N_41400,N_38610,N_39832);
or U41401 (N_41401,N_39078,N_39079);
and U41402 (N_41402,N_38893,N_38126);
nor U41403 (N_41403,N_37522,N_39393);
nand U41404 (N_41404,N_37754,N_38081);
nand U41405 (N_41405,N_39133,N_38198);
nand U41406 (N_41406,N_39455,N_38010);
nor U41407 (N_41407,N_38182,N_38505);
nor U41408 (N_41408,N_38713,N_39788);
nor U41409 (N_41409,N_39523,N_39986);
and U41410 (N_41410,N_39496,N_39614);
nand U41411 (N_41411,N_38944,N_39444);
nand U41412 (N_41412,N_37722,N_37584);
nand U41413 (N_41413,N_39192,N_39215);
nor U41414 (N_41414,N_38355,N_38350);
nand U41415 (N_41415,N_39252,N_37867);
and U41416 (N_41416,N_39173,N_39002);
nand U41417 (N_41417,N_38814,N_39013);
nand U41418 (N_41418,N_38186,N_39898);
and U41419 (N_41419,N_39728,N_38128);
xor U41420 (N_41420,N_38505,N_38349);
nand U41421 (N_41421,N_39689,N_39000);
xnor U41422 (N_41422,N_39171,N_39904);
or U41423 (N_41423,N_38445,N_37516);
and U41424 (N_41424,N_37939,N_39591);
or U41425 (N_41425,N_38496,N_38497);
and U41426 (N_41426,N_37719,N_39882);
and U41427 (N_41427,N_39133,N_37651);
nor U41428 (N_41428,N_39834,N_38723);
nand U41429 (N_41429,N_38262,N_37744);
xnor U41430 (N_41430,N_38762,N_39148);
or U41431 (N_41431,N_39447,N_38940);
or U41432 (N_41432,N_39670,N_38692);
nor U41433 (N_41433,N_37520,N_38676);
xnor U41434 (N_41434,N_38586,N_37975);
nor U41435 (N_41435,N_37695,N_38410);
or U41436 (N_41436,N_39880,N_38263);
nand U41437 (N_41437,N_39371,N_38266);
and U41438 (N_41438,N_39616,N_39477);
or U41439 (N_41439,N_37542,N_39184);
nor U41440 (N_41440,N_39235,N_38734);
xnor U41441 (N_41441,N_38133,N_39782);
xnor U41442 (N_41442,N_39441,N_37681);
or U41443 (N_41443,N_39001,N_38576);
or U41444 (N_41444,N_37548,N_38644);
nand U41445 (N_41445,N_38338,N_39867);
xnor U41446 (N_41446,N_38628,N_39820);
xor U41447 (N_41447,N_39573,N_37778);
xnor U41448 (N_41448,N_38246,N_39614);
nor U41449 (N_41449,N_39012,N_38592);
and U41450 (N_41450,N_37771,N_37748);
nor U41451 (N_41451,N_38300,N_38831);
xor U41452 (N_41452,N_38213,N_39487);
xor U41453 (N_41453,N_37686,N_38913);
xor U41454 (N_41454,N_39337,N_37837);
or U41455 (N_41455,N_38460,N_37560);
nor U41456 (N_41456,N_39205,N_39361);
xor U41457 (N_41457,N_39595,N_38420);
xnor U41458 (N_41458,N_38602,N_38073);
and U41459 (N_41459,N_38091,N_38431);
and U41460 (N_41460,N_38863,N_37656);
and U41461 (N_41461,N_39216,N_38394);
xnor U41462 (N_41462,N_38198,N_39604);
or U41463 (N_41463,N_39857,N_37592);
xnor U41464 (N_41464,N_38463,N_39042);
and U41465 (N_41465,N_39680,N_38296);
or U41466 (N_41466,N_38165,N_37736);
or U41467 (N_41467,N_37795,N_38759);
or U41468 (N_41468,N_39167,N_38710);
xor U41469 (N_41469,N_38612,N_38217);
or U41470 (N_41470,N_37785,N_38503);
nand U41471 (N_41471,N_39791,N_38927);
or U41472 (N_41472,N_37773,N_38629);
or U41473 (N_41473,N_38395,N_38451);
xor U41474 (N_41474,N_38163,N_37968);
and U41475 (N_41475,N_38273,N_38086);
and U41476 (N_41476,N_38698,N_38237);
xor U41477 (N_41477,N_38475,N_39971);
nor U41478 (N_41478,N_39555,N_39339);
xor U41479 (N_41479,N_39915,N_37527);
xnor U41480 (N_41480,N_38903,N_39055);
or U41481 (N_41481,N_37585,N_38591);
xnor U41482 (N_41482,N_39753,N_38241);
xnor U41483 (N_41483,N_38081,N_38182);
nor U41484 (N_41484,N_37666,N_38612);
or U41485 (N_41485,N_39944,N_39783);
xor U41486 (N_41486,N_38170,N_38151);
nand U41487 (N_41487,N_38883,N_39972);
nand U41488 (N_41488,N_38300,N_38096);
and U41489 (N_41489,N_39096,N_39854);
nor U41490 (N_41490,N_38062,N_38891);
and U41491 (N_41491,N_38009,N_39843);
nand U41492 (N_41492,N_38701,N_39342);
or U41493 (N_41493,N_38421,N_39583);
nor U41494 (N_41494,N_39247,N_38196);
or U41495 (N_41495,N_38203,N_38259);
and U41496 (N_41496,N_38469,N_38657);
xor U41497 (N_41497,N_37658,N_39623);
nand U41498 (N_41498,N_38463,N_38500);
or U41499 (N_41499,N_39258,N_39268);
and U41500 (N_41500,N_39336,N_39235);
xnor U41501 (N_41501,N_38493,N_39112);
nand U41502 (N_41502,N_38090,N_39790);
or U41503 (N_41503,N_39530,N_38621);
nor U41504 (N_41504,N_38140,N_38355);
and U41505 (N_41505,N_38015,N_39888);
or U41506 (N_41506,N_38532,N_38918);
xnor U41507 (N_41507,N_39996,N_38227);
and U41508 (N_41508,N_38512,N_38649);
nand U41509 (N_41509,N_39252,N_38391);
nand U41510 (N_41510,N_37689,N_38973);
or U41511 (N_41511,N_39105,N_39586);
or U41512 (N_41512,N_39621,N_38210);
xor U41513 (N_41513,N_37540,N_39186);
nand U41514 (N_41514,N_39193,N_39736);
xnor U41515 (N_41515,N_39686,N_39866);
nand U41516 (N_41516,N_39572,N_38759);
and U41517 (N_41517,N_38237,N_39505);
nor U41518 (N_41518,N_38117,N_39764);
and U41519 (N_41519,N_37883,N_37562);
and U41520 (N_41520,N_38289,N_38541);
and U41521 (N_41521,N_38956,N_37976);
or U41522 (N_41522,N_37818,N_38566);
xnor U41523 (N_41523,N_39919,N_39588);
nand U41524 (N_41524,N_39664,N_37525);
nand U41525 (N_41525,N_39888,N_38460);
or U41526 (N_41526,N_39225,N_39575);
and U41527 (N_41527,N_38171,N_39410);
nand U41528 (N_41528,N_37746,N_38643);
xor U41529 (N_41529,N_39960,N_39711);
or U41530 (N_41530,N_39550,N_38469);
xor U41531 (N_41531,N_37829,N_39048);
nand U41532 (N_41532,N_38107,N_39950);
and U41533 (N_41533,N_37708,N_38555);
nand U41534 (N_41534,N_38458,N_38695);
and U41535 (N_41535,N_37609,N_37800);
and U41536 (N_41536,N_38155,N_39052);
xnor U41537 (N_41537,N_38015,N_39362);
nand U41538 (N_41538,N_37903,N_39749);
nor U41539 (N_41539,N_39505,N_38432);
nor U41540 (N_41540,N_38601,N_38546);
xnor U41541 (N_41541,N_38381,N_39062);
nor U41542 (N_41542,N_39996,N_37657);
or U41543 (N_41543,N_38492,N_38028);
xnor U41544 (N_41544,N_38943,N_39367);
and U41545 (N_41545,N_38675,N_37656);
or U41546 (N_41546,N_38095,N_38304);
nand U41547 (N_41547,N_39473,N_39210);
xnor U41548 (N_41548,N_37963,N_39836);
nor U41549 (N_41549,N_39932,N_38677);
nand U41550 (N_41550,N_38833,N_39216);
and U41551 (N_41551,N_38757,N_38242);
nand U41552 (N_41552,N_39541,N_38673);
or U41553 (N_41553,N_39113,N_37960);
or U41554 (N_41554,N_39738,N_38635);
nor U41555 (N_41555,N_37695,N_39776);
xor U41556 (N_41556,N_37919,N_38707);
xor U41557 (N_41557,N_39373,N_38903);
and U41558 (N_41558,N_37938,N_38854);
nand U41559 (N_41559,N_38409,N_39347);
nand U41560 (N_41560,N_37710,N_39036);
nand U41561 (N_41561,N_39688,N_38108);
and U41562 (N_41562,N_38148,N_39686);
and U41563 (N_41563,N_38622,N_38996);
nor U41564 (N_41564,N_37878,N_37973);
nor U41565 (N_41565,N_39444,N_38866);
nand U41566 (N_41566,N_38212,N_38877);
nand U41567 (N_41567,N_37913,N_39061);
nand U41568 (N_41568,N_37589,N_37510);
or U41569 (N_41569,N_37938,N_39678);
nand U41570 (N_41570,N_38745,N_38700);
nor U41571 (N_41571,N_38825,N_39825);
xor U41572 (N_41572,N_38727,N_37899);
nor U41573 (N_41573,N_38027,N_39198);
xor U41574 (N_41574,N_39436,N_38970);
nand U41575 (N_41575,N_38761,N_38012);
or U41576 (N_41576,N_38148,N_39137);
or U41577 (N_41577,N_38798,N_39172);
or U41578 (N_41578,N_38315,N_39780);
nor U41579 (N_41579,N_38214,N_39738);
nor U41580 (N_41580,N_39319,N_37587);
nand U41581 (N_41581,N_37515,N_39593);
and U41582 (N_41582,N_38250,N_39895);
nor U41583 (N_41583,N_39035,N_38061);
and U41584 (N_41584,N_37759,N_37866);
xnor U41585 (N_41585,N_37923,N_38569);
nand U41586 (N_41586,N_37901,N_39434);
nor U41587 (N_41587,N_38949,N_38146);
or U41588 (N_41588,N_38612,N_39372);
xnor U41589 (N_41589,N_39331,N_39448);
or U41590 (N_41590,N_37507,N_39383);
nor U41591 (N_41591,N_37907,N_38435);
xnor U41592 (N_41592,N_38191,N_37698);
nand U41593 (N_41593,N_38176,N_38822);
xnor U41594 (N_41594,N_39252,N_37721);
and U41595 (N_41595,N_39430,N_39693);
nor U41596 (N_41596,N_37845,N_38715);
and U41597 (N_41597,N_38583,N_37543);
xor U41598 (N_41598,N_39952,N_38762);
nor U41599 (N_41599,N_37951,N_39775);
nor U41600 (N_41600,N_39596,N_39287);
and U41601 (N_41601,N_39539,N_39096);
nand U41602 (N_41602,N_39618,N_38596);
and U41603 (N_41603,N_38963,N_39083);
nor U41604 (N_41604,N_39640,N_38527);
nor U41605 (N_41605,N_37566,N_38998);
or U41606 (N_41606,N_38393,N_37604);
or U41607 (N_41607,N_38992,N_38050);
or U41608 (N_41608,N_39419,N_38920);
nand U41609 (N_41609,N_39346,N_39743);
nor U41610 (N_41610,N_37550,N_39979);
nor U41611 (N_41611,N_38264,N_39258);
and U41612 (N_41612,N_38612,N_37583);
or U41613 (N_41613,N_39565,N_37917);
nor U41614 (N_41614,N_37869,N_39724);
and U41615 (N_41615,N_37710,N_38341);
nand U41616 (N_41616,N_39012,N_39177);
nor U41617 (N_41617,N_39751,N_39701);
and U41618 (N_41618,N_39584,N_37966);
nor U41619 (N_41619,N_38020,N_39823);
or U41620 (N_41620,N_38758,N_38097);
nand U41621 (N_41621,N_39264,N_39660);
or U41622 (N_41622,N_39136,N_38664);
and U41623 (N_41623,N_39782,N_37793);
nor U41624 (N_41624,N_39635,N_38243);
and U41625 (N_41625,N_39585,N_38401);
or U41626 (N_41626,N_38864,N_38358);
xnor U41627 (N_41627,N_39362,N_39788);
or U41628 (N_41628,N_38915,N_38053);
or U41629 (N_41629,N_37907,N_38852);
or U41630 (N_41630,N_37547,N_39925);
or U41631 (N_41631,N_38890,N_39673);
xor U41632 (N_41632,N_38966,N_38982);
nor U41633 (N_41633,N_38078,N_39379);
xor U41634 (N_41634,N_39556,N_39498);
and U41635 (N_41635,N_38460,N_38833);
and U41636 (N_41636,N_39959,N_37759);
nand U41637 (N_41637,N_38218,N_37857);
nand U41638 (N_41638,N_39007,N_39685);
nor U41639 (N_41639,N_38920,N_39504);
xor U41640 (N_41640,N_39830,N_39189);
xnor U41641 (N_41641,N_39197,N_38570);
nand U41642 (N_41642,N_37896,N_39776);
and U41643 (N_41643,N_39691,N_37521);
nand U41644 (N_41644,N_38883,N_37737);
nand U41645 (N_41645,N_38559,N_39421);
or U41646 (N_41646,N_39171,N_38192);
nand U41647 (N_41647,N_38548,N_38830);
and U41648 (N_41648,N_37574,N_38764);
or U41649 (N_41649,N_37577,N_39466);
or U41650 (N_41650,N_37853,N_38482);
nor U41651 (N_41651,N_38734,N_38095);
xnor U41652 (N_41652,N_38507,N_39133);
xor U41653 (N_41653,N_38599,N_39728);
nand U41654 (N_41654,N_38711,N_39941);
and U41655 (N_41655,N_39682,N_38248);
nand U41656 (N_41656,N_38750,N_38816);
nand U41657 (N_41657,N_37778,N_39948);
nand U41658 (N_41658,N_39419,N_38291);
or U41659 (N_41659,N_39131,N_39184);
nor U41660 (N_41660,N_38772,N_38393);
xor U41661 (N_41661,N_38355,N_37627);
or U41662 (N_41662,N_38052,N_37688);
xnor U41663 (N_41663,N_38902,N_39506);
xnor U41664 (N_41664,N_39153,N_39661);
nor U41665 (N_41665,N_39847,N_37673);
xor U41666 (N_41666,N_39316,N_38043);
or U41667 (N_41667,N_37670,N_39920);
nor U41668 (N_41668,N_37953,N_38385);
or U41669 (N_41669,N_38926,N_39571);
xnor U41670 (N_41670,N_38915,N_38009);
nor U41671 (N_41671,N_37662,N_39753);
xor U41672 (N_41672,N_39705,N_37753);
xnor U41673 (N_41673,N_39304,N_38502);
and U41674 (N_41674,N_38484,N_39252);
nand U41675 (N_41675,N_38640,N_39149);
or U41676 (N_41676,N_38020,N_39190);
and U41677 (N_41677,N_38661,N_39734);
or U41678 (N_41678,N_38366,N_39898);
nor U41679 (N_41679,N_39835,N_38453);
nand U41680 (N_41680,N_38765,N_38788);
or U41681 (N_41681,N_39126,N_39598);
nand U41682 (N_41682,N_39717,N_38089);
xor U41683 (N_41683,N_38402,N_37978);
nor U41684 (N_41684,N_39222,N_39254);
nand U41685 (N_41685,N_38942,N_38180);
and U41686 (N_41686,N_38481,N_37603);
nand U41687 (N_41687,N_38418,N_38585);
or U41688 (N_41688,N_37570,N_38363);
or U41689 (N_41689,N_39942,N_39972);
or U41690 (N_41690,N_39722,N_38881);
nand U41691 (N_41691,N_38397,N_38040);
nor U41692 (N_41692,N_37772,N_39313);
nor U41693 (N_41693,N_38808,N_38604);
nor U41694 (N_41694,N_39783,N_38391);
nor U41695 (N_41695,N_39548,N_38978);
xnor U41696 (N_41696,N_37770,N_39841);
nor U41697 (N_41697,N_39587,N_38246);
and U41698 (N_41698,N_39610,N_38670);
nand U41699 (N_41699,N_37601,N_37747);
nor U41700 (N_41700,N_38994,N_38856);
nand U41701 (N_41701,N_39372,N_37605);
xnor U41702 (N_41702,N_39283,N_37503);
xnor U41703 (N_41703,N_38532,N_39970);
xor U41704 (N_41704,N_39805,N_37536);
nor U41705 (N_41705,N_38704,N_38239);
xnor U41706 (N_41706,N_39279,N_39384);
xnor U41707 (N_41707,N_39100,N_38285);
xor U41708 (N_41708,N_39297,N_37846);
or U41709 (N_41709,N_38100,N_38182);
or U41710 (N_41710,N_38561,N_38110);
nand U41711 (N_41711,N_38371,N_38596);
or U41712 (N_41712,N_37913,N_37625);
or U41713 (N_41713,N_39871,N_39214);
and U41714 (N_41714,N_37570,N_38618);
nor U41715 (N_41715,N_37745,N_39188);
xor U41716 (N_41716,N_37851,N_39302);
and U41717 (N_41717,N_38832,N_38571);
nand U41718 (N_41718,N_39575,N_37856);
or U41719 (N_41719,N_39820,N_39457);
nor U41720 (N_41720,N_37568,N_37735);
and U41721 (N_41721,N_38569,N_38374);
or U41722 (N_41722,N_39496,N_37627);
or U41723 (N_41723,N_39975,N_39212);
nor U41724 (N_41724,N_38270,N_38761);
and U41725 (N_41725,N_38633,N_38428);
and U41726 (N_41726,N_39691,N_38437);
xor U41727 (N_41727,N_37954,N_37897);
xor U41728 (N_41728,N_38808,N_38338);
nand U41729 (N_41729,N_38972,N_37546);
xor U41730 (N_41730,N_39290,N_38510);
or U41731 (N_41731,N_39015,N_39223);
xor U41732 (N_41732,N_38243,N_37518);
xnor U41733 (N_41733,N_37562,N_39284);
nand U41734 (N_41734,N_38892,N_38105);
or U41735 (N_41735,N_39877,N_37687);
or U41736 (N_41736,N_39262,N_37804);
nor U41737 (N_41737,N_38417,N_39900);
nor U41738 (N_41738,N_39890,N_39989);
or U41739 (N_41739,N_38769,N_38064);
xnor U41740 (N_41740,N_38078,N_37707);
or U41741 (N_41741,N_38933,N_37519);
xor U41742 (N_41742,N_39656,N_38718);
nand U41743 (N_41743,N_39530,N_39963);
nor U41744 (N_41744,N_37895,N_37833);
and U41745 (N_41745,N_37858,N_39562);
nand U41746 (N_41746,N_37931,N_38074);
nor U41747 (N_41747,N_39407,N_37627);
or U41748 (N_41748,N_39930,N_39413);
xor U41749 (N_41749,N_39110,N_38443);
xor U41750 (N_41750,N_38410,N_39862);
and U41751 (N_41751,N_39256,N_39613);
or U41752 (N_41752,N_38058,N_37590);
nand U41753 (N_41753,N_39459,N_38838);
nand U41754 (N_41754,N_39442,N_38972);
nand U41755 (N_41755,N_38727,N_39091);
nand U41756 (N_41756,N_38665,N_39999);
nor U41757 (N_41757,N_37774,N_38572);
or U41758 (N_41758,N_38002,N_38193);
or U41759 (N_41759,N_38163,N_38176);
nor U41760 (N_41760,N_39946,N_39580);
nor U41761 (N_41761,N_39715,N_39003);
nand U41762 (N_41762,N_38550,N_39516);
or U41763 (N_41763,N_38260,N_38913);
or U41764 (N_41764,N_38873,N_39863);
and U41765 (N_41765,N_38902,N_39623);
nand U41766 (N_41766,N_38534,N_38544);
or U41767 (N_41767,N_37814,N_39445);
nor U41768 (N_41768,N_38739,N_38140);
xnor U41769 (N_41769,N_39310,N_38086);
nand U41770 (N_41770,N_38142,N_38613);
nand U41771 (N_41771,N_38499,N_38851);
nand U41772 (N_41772,N_39996,N_39350);
nor U41773 (N_41773,N_39260,N_39384);
nand U41774 (N_41774,N_39483,N_38867);
and U41775 (N_41775,N_38727,N_38237);
nor U41776 (N_41776,N_38028,N_39261);
nor U41777 (N_41777,N_38679,N_39776);
nor U41778 (N_41778,N_39835,N_37571);
and U41779 (N_41779,N_38678,N_39546);
xor U41780 (N_41780,N_38453,N_38015);
nand U41781 (N_41781,N_38415,N_37911);
and U41782 (N_41782,N_37838,N_39170);
and U41783 (N_41783,N_39889,N_39059);
nand U41784 (N_41784,N_37723,N_37566);
or U41785 (N_41785,N_37669,N_37867);
xnor U41786 (N_41786,N_38899,N_38312);
nand U41787 (N_41787,N_38773,N_39072);
xor U41788 (N_41788,N_37701,N_37601);
xor U41789 (N_41789,N_38825,N_37639);
nand U41790 (N_41790,N_37739,N_38152);
xnor U41791 (N_41791,N_37957,N_38629);
and U41792 (N_41792,N_39539,N_38638);
nand U41793 (N_41793,N_39191,N_38143);
and U41794 (N_41794,N_38882,N_39262);
or U41795 (N_41795,N_38238,N_37579);
nand U41796 (N_41796,N_37952,N_39256);
nand U41797 (N_41797,N_38921,N_38863);
and U41798 (N_41798,N_39188,N_39909);
xor U41799 (N_41799,N_38218,N_37831);
and U41800 (N_41800,N_38891,N_38436);
or U41801 (N_41801,N_39616,N_39324);
xnor U41802 (N_41802,N_37894,N_39029);
or U41803 (N_41803,N_38780,N_37741);
and U41804 (N_41804,N_38101,N_39757);
nand U41805 (N_41805,N_38026,N_37822);
or U41806 (N_41806,N_39079,N_39827);
and U41807 (N_41807,N_37859,N_38096);
nand U41808 (N_41808,N_39859,N_37735);
or U41809 (N_41809,N_39806,N_39263);
xnor U41810 (N_41810,N_39136,N_38768);
and U41811 (N_41811,N_39252,N_39588);
xor U41812 (N_41812,N_38555,N_39638);
xor U41813 (N_41813,N_39176,N_38156);
nor U41814 (N_41814,N_37641,N_38052);
or U41815 (N_41815,N_39789,N_37643);
xor U41816 (N_41816,N_37943,N_38808);
nor U41817 (N_41817,N_37624,N_39032);
and U41818 (N_41818,N_39228,N_38001);
nand U41819 (N_41819,N_39893,N_39214);
nand U41820 (N_41820,N_39936,N_38486);
or U41821 (N_41821,N_39977,N_38536);
and U41822 (N_41822,N_38058,N_38325);
nor U41823 (N_41823,N_37585,N_39000);
or U41824 (N_41824,N_39160,N_38495);
nand U41825 (N_41825,N_39016,N_39332);
xnor U41826 (N_41826,N_39133,N_38079);
nor U41827 (N_41827,N_38577,N_38757);
nand U41828 (N_41828,N_39283,N_37860);
xnor U41829 (N_41829,N_37888,N_39152);
nor U41830 (N_41830,N_38897,N_37829);
xnor U41831 (N_41831,N_38038,N_38592);
or U41832 (N_41832,N_37640,N_38443);
nor U41833 (N_41833,N_39438,N_38797);
xor U41834 (N_41834,N_38394,N_39979);
or U41835 (N_41835,N_39611,N_39100);
or U41836 (N_41836,N_39889,N_39102);
and U41837 (N_41837,N_37928,N_37907);
and U41838 (N_41838,N_38677,N_39153);
or U41839 (N_41839,N_38878,N_39014);
nand U41840 (N_41840,N_38452,N_37924);
or U41841 (N_41841,N_38473,N_39257);
and U41842 (N_41842,N_39741,N_37505);
nand U41843 (N_41843,N_38409,N_39523);
nor U41844 (N_41844,N_39165,N_38783);
nor U41845 (N_41845,N_37953,N_39289);
xor U41846 (N_41846,N_39294,N_38246);
and U41847 (N_41847,N_39685,N_39719);
nor U41848 (N_41848,N_37964,N_39023);
nand U41849 (N_41849,N_39631,N_38259);
nor U41850 (N_41850,N_39778,N_37832);
nor U41851 (N_41851,N_38075,N_38798);
or U41852 (N_41852,N_38932,N_37722);
and U41853 (N_41853,N_38109,N_38832);
xnor U41854 (N_41854,N_39683,N_37633);
nand U41855 (N_41855,N_38481,N_39426);
xnor U41856 (N_41856,N_39903,N_37723);
nand U41857 (N_41857,N_37769,N_39307);
or U41858 (N_41858,N_39050,N_37533);
xor U41859 (N_41859,N_38666,N_39351);
or U41860 (N_41860,N_38512,N_37511);
or U41861 (N_41861,N_38891,N_38195);
or U41862 (N_41862,N_38158,N_38215);
xnor U41863 (N_41863,N_39838,N_39273);
or U41864 (N_41864,N_38925,N_37920);
or U41865 (N_41865,N_38740,N_38260);
or U41866 (N_41866,N_38453,N_39254);
and U41867 (N_41867,N_38038,N_38810);
nor U41868 (N_41868,N_37887,N_37572);
nand U41869 (N_41869,N_38726,N_37648);
nor U41870 (N_41870,N_38039,N_39574);
and U41871 (N_41871,N_38303,N_39524);
or U41872 (N_41872,N_38736,N_39269);
xor U41873 (N_41873,N_39282,N_39864);
or U41874 (N_41874,N_39431,N_38017);
nand U41875 (N_41875,N_39524,N_37689);
and U41876 (N_41876,N_38425,N_37930);
and U41877 (N_41877,N_38929,N_38750);
nand U41878 (N_41878,N_38442,N_38859);
or U41879 (N_41879,N_38224,N_38030);
nor U41880 (N_41880,N_39073,N_39825);
or U41881 (N_41881,N_38441,N_38268);
nor U41882 (N_41882,N_37928,N_38310);
and U41883 (N_41883,N_38000,N_37947);
nand U41884 (N_41884,N_39063,N_39110);
nor U41885 (N_41885,N_38121,N_37849);
xnor U41886 (N_41886,N_39410,N_38516);
and U41887 (N_41887,N_39224,N_39660);
xor U41888 (N_41888,N_38845,N_38003);
nand U41889 (N_41889,N_38425,N_38563);
or U41890 (N_41890,N_39169,N_38845);
nor U41891 (N_41891,N_38427,N_39763);
nor U41892 (N_41892,N_39713,N_38107);
nand U41893 (N_41893,N_38678,N_38233);
xnor U41894 (N_41894,N_37727,N_37666);
or U41895 (N_41895,N_39359,N_39324);
xnor U41896 (N_41896,N_39116,N_38103);
or U41897 (N_41897,N_38146,N_37649);
nor U41898 (N_41898,N_38282,N_39557);
and U41899 (N_41899,N_37613,N_39884);
or U41900 (N_41900,N_38330,N_37715);
xor U41901 (N_41901,N_38063,N_39924);
nand U41902 (N_41902,N_39257,N_39951);
nand U41903 (N_41903,N_39450,N_38557);
nor U41904 (N_41904,N_38410,N_38747);
or U41905 (N_41905,N_38827,N_37882);
and U41906 (N_41906,N_37749,N_39797);
nand U41907 (N_41907,N_38146,N_39546);
and U41908 (N_41908,N_39558,N_39830);
or U41909 (N_41909,N_37715,N_37806);
nor U41910 (N_41910,N_37519,N_38505);
or U41911 (N_41911,N_39268,N_39884);
and U41912 (N_41912,N_38152,N_39184);
or U41913 (N_41913,N_37728,N_38089);
or U41914 (N_41914,N_39418,N_38719);
nand U41915 (N_41915,N_39953,N_39483);
nor U41916 (N_41916,N_39059,N_38906);
nand U41917 (N_41917,N_37844,N_38281);
and U41918 (N_41918,N_38010,N_38446);
nor U41919 (N_41919,N_38037,N_39291);
and U41920 (N_41920,N_39410,N_38150);
and U41921 (N_41921,N_39013,N_38991);
nand U41922 (N_41922,N_38119,N_37953);
or U41923 (N_41923,N_39067,N_39402);
nor U41924 (N_41924,N_39455,N_38536);
or U41925 (N_41925,N_39140,N_38697);
nor U41926 (N_41926,N_37925,N_38106);
and U41927 (N_41927,N_39942,N_38618);
and U41928 (N_41928,N_38328,N_37767);
nand U41929 (N_41929,N_37720,N_39760);
and U41930 (N_41930,N_39205,N_37533);
nor U41931 (N_41931,N_39014,N_38401);
or U41932 (N_41932,N_37926,N_39316);
and U41933 (N_41933,N_37550,N_39275);
nor U41934 (N_41934,N_39383,N_38855);
or U41935 (N_41935,N_38143,N_38493);
xor U41936 (N_41936,N_39899,N_39090);
nand U41937 (N_41937,N_38695,N_39111);
and U41938 (N_41938,N_38291,N_38383);
nor U41939 (N_41939,N_39868,N_39213);
nor U41940 (N_41940,N_38458,N_38196);
nor U41941 (N_41941,N_38084,N_38445);
or U41942 (N_41942,N_38213,N_37656);
or U41943 (N_41943,N_38038,N_37858);
xnor U41944 (N_41944,N_37577,N_39694);
nand U41945 (N_41945,N_38003,N_39836);
and U41946 (N_41946,N_38800,N_39845);
nand U41947 (N_41947,N_39318,N_39788);
xor U41948 (N_41948,N_39745,N_39071);
xor U41949 (N_41949,N_37841,N_39775);
xor U41950 (N_41950,N_38332,N_38612);
xor U41951 (N_41951,N_39806,N_39941);
or U41952 (N_41952,N_37880,N_39263);
or U41953 (N_41953,N_39846,N_39775);
xnor U41954 (N_41954,N_38527,N_38966);
xnor U41955 (N_41955,N_38384,N_39708);
xnor U41956 (N_41956,N_37520,N_39278);
or U41957 (N_41957,N_38997,N_39185);
and U41958 (N_41958,N_38471,N_38912);
nor U41959 (N_41959,N_37867,N_38783);
xor U41960 (N_41960,N_38466,N_37947);
xnor U41961 (N_41961,N_38891,N_38795);
nor U41962 (N_41962,N_39836,N_39319);
and U41963 (N_41963,N_38169,N_39061);
nor U41964 (N_41964,N_37572,N_37527);
nor U41965 (N_41965,N_38612,N_39638);
nor U41966 (N_41966,N_37657,N_39148);
or U41967 (N_41967,N_38224,N_38175);
and U41968 (N_41968,N_38326,N_37843);
xor U41969 (N_41969,N_38283,N_38935);
xnor U41970 (N_41970,N_37679,N_39388);
or U41971 (N_41971,N_37812,N_39548);
or U41972 (N_41972,N_39276,N_38016);
nand U41973 (N_41973,N_39201,N_39666);
or U41974 (N_41974,N_38080,N_38007);
nor U41975 (N_41975,N_37522,N_38346);
or U41976 (N_41976,N_37691,N_39767);
or U41977 (N_41977,N_37882,N_39016);
nor U41978 (N_41978,N_39932,N_39971);
or U41979 (N_41979,N_38945,N_39415);
xnor U41980 (N_41980,N_38906,N_39981);
nor U41981 (N_41981,N_39272,N_39420);
and U41982 (N_41982,N_39351,N_37547);
or U41983 (N_41983,N_39657,N_39885);
or U41984 (N_41984,N_37770,N_37655);
or U41985 (N_41985,N_39838,N_37633);
xor U41986 (N_41986,N_39222,N_37932);
or U41987 (N_41987,N_38525,N_38356);
nand U41988 (N_41988,N_38810,N_38041);
nand U41989 (N_41989,N_39017,N_39533);
and U41990 (N_41990,N_38652,N_38128);
and U41991 (N_41991,N_38726,N_38619);
and U41992 (N_41992,N_38170,N_37802);
nor U41993 (N_41993,N_38846,N_39645);
and U41994 (N_41994,N_38923,N_39445);
and U41995 (N_41995,N_39018,N_38533);
xnor U41996 (N_41996,N_39020,N_39984);
xnor U41997 (N_41997,N_37546,N_38091);
nor U41998 (N_41998,N_38405,N_39178);
nand U41999 (N_41999,N_38598,N_39046);
xor U42000 (N_42000,N_39286,N_39434);
xor U42001 (N_42001,N_37961,N_38549);
xor U42002 (N_42002,N_39764,N_39616);
xor U42003 (N_42003,N_39593,N_39443);
and U42004 (N_42004,N_39300,N_39736);
and U42005 (N_42005,N_38892,N_37693);
nor U42006 (N_42006,N_39456,N_37654);
nor U42007 (N_42007,N_38518,N_39352);
or U42008 (N_42008,N_38690,N_39457);
and U42009 (N_42009,N_37753,N_38139);
xor U42010 (N_42010,N_37526,N_39994);
and U42011 (N_42011,N_39459,N_39231);
xor U42012 (N_42012,N_39804,N_39405);
nand U42013 (N_42013,N_39515,N_37842);
nor U42014 (N_42014,N_38532,N_38820);
nor U42015 (N_42015,N_39641,N_39596);
nor U42016 (N_42016,N_39909,N_37538);
xor U42017 (N_42017,N_37945,N_38251);
nor U42018 (N_42018,N_39174,N_39619);
nand U42019 (N_42019,N_39111,N_38289);
or U42020 (N_42020,N_38137,N_38668);
or U42021 (N_42021,N_38941,N_38739);
xnor U42022 (N_42022,N_38130,N_38833);
and U42023 (N_42023,N_39095,N_39319);
xnor U42024 (N_42024,N_38429,N_38740);
or U42025 (N_42025,N_38663,N_38676);
nand U42026 (N_42026,N_38617,N_37573);
and U42027 (N_42027,N_39779,N_39241);
xnor U42028 (N_42028,N_38560,N_39231);
and U42029 (N_42029,N_38848,N_39331);
nor U42030 (N_42030,N_37575,N_38382);
or U42031 (N_42031,N_38372,N_38281);
xor U42032 (N_42032,N_38320,N_37622);
and U42033 (N_42033,N_37701,N_39917);
nand U42034 (N_42034,N_38780,N_39499);
nor U42035 (N_42035,N_37677,N_38938);
nor U42036 (N_42036,N_38151,N_38652);
nand U42037 (N_42037,N_38305,N_39068);
nand U42038 (N_42038,N_38448,N_37508);
nand U42039 (N_42039,N_37996,N_38678);
nor U42040 (N_42040,N_38085,N_37940);
xor U42041 (N_42041,N_38451,N_37836);
nand U42042 (N_42042,N_39158,N_38517);
nor U42043 (N_42043,N_39329,N_39560);
nor U42044 (N_42044,N_38220,N_39121);
and U42045 (N_42045,N_39382,N_38421);
or U42046 (N_42046,N_39343,N_39524);
or U42047 (N_42047,N_39128,N_38376);
xnor U42048 (N_42048,N_38194,N_38358);
or U42049 (N_42049,N_39387,N_39274);
xor U42050 (N_42050,N_39364,N_39214);
and U42051 (N_42051,N_38828,N_37946);
nand U42052 (N_42052,N_38271,N_37865);
nor U42053 (N_42053,N_39094,N_38349);
nand U42054 (N_42054,N_38504,N_39120);
nor U42055 (N_42055,N_37866,N_39733);
xor U42056 (N_42056,N_39630,N_37649);
xor U42057 (N_42057,N_39005,N_37639);
xor U42058 (N_42058,N_39805,N_38097);
nand U42059 (N_42059,N_39059,N_37757);
nor U42060 (N_42060,N_38493,N_39128);
or U42061 (N_42061,N_37778,N_38127);
and U42062 (N_42062,N_39440,N_39086);
nand U42063 (N_42063,N_38133,N_39110);
nand U42064 (N_42064,N_38696,N_38336);
and U42065 (N_42065,N_38529,N_39819);
nor U42066 (N_42066,N_37539,N_38404);
or U42067 (N_42067,N_38342,N_38636);
nor U42068 (N_42068,N_39031,N_37880);
or U42069 (N_42069,N_39090,N_38624);
nand U42070 (N_42070,N_38757,N_38487);
and U42071 (N_42071,N_39316,N_39677);
and U42072 (N_42072,N_39209,N_37787);
or U42073 (N_42073,N_39201,N_38503);
and U42074 (N_42074,N_39783,N_37885);
nor U42075 (N_42075,N_39654,N_39204);
nand U42076 (N_42076,N_38320,N_39913);
or U42077 (N_42077,N_38608,N_37899);
nand U42078 (N_42078,N_39730,N_39939);
and U42079 (N_42079,N_38500,N_38977);
and U42080 (N_42080,N_39334,N_39995);
nor U42081 (N_42081,N_38193,N_39866);
nand U42082 (N_42082,N_39480,N_38164);
xor U42083 (N_42083,N_38880,N_39380);
and U42084 (N_42084,N_37771,N_39448);
or U42085 (N_42085,N_39498,N_39476);
xor U42086 (N_42086,N_39891,N_38008);
xnor U42087 (N_42087,N_39666,N_37915);
xnor U42088 (N_42088,N_39731,N_39729);
and U42089 (N_42089,N_38784,N_37588);
or U42090 (N_42090,N_37633,N_38871);
nor U42091 (N_42091,N_39443,N_37988);
xnor U42092 (N_42092,N_37667,N_39150);
xnor U42093 (N_42093,N_39306,N_38849);
and U42094 (N_42094,N_39261,N_39594);
and U42095 (N_42095,N_37919,N_38182);
nor U42096 (N_42096,N_39394,N_39416);
nor U42097 (N_42097,N_39412,N_38435);
and U42098 (N_42098,N_39023,N_39955);
and U42099 (N_42099,N_37791,N_38481);
nand U42100 (N_42100,N_37773,N_39614);
xnor U42101 (N_42101,N_39066,N_38940);
nand U42102 (N_42102,N_37798,N_38814);
nor U42103 (N_42103,N_39098,N_39115);
or U42104 (N_42104,N_39388,N_38537);
nor U42105 (N_42105,N_39450,N_37585);
and U42106 (N_42106,N_39777,N_39710);
and U42107 (N_42107,N_38210,N_39331);
nor U42108 (N_42108,N_38732,N_38855);
xnor U42109 (N_42109,N_38223,N_39282);
or U42110 (N_42110,N_38459,N_39827);
xnor U42111 (N_42111,N_38421,N_39772);
xnor U42112 (N_42112,N_38445,N_39007);
or U42113 (N_42113,N_37767,N_39401);
xor U42114 (N_42114,N_39140,N_38700);
nor U42115 (N_42115,N_39825,N_39662);
or U42116 (N_42116,N_38214,N_37740);
and U42117 (N_42117,N_38397,N_38369);
and U42118 (N_42118,N_38548,N_39385);
nand U42119 (N_42119,N_38629,N_38780);
or U42120 (N_42120,N_38399,N_39618);
or U42121 (N_42121,N_38376,N_38178);
xor U42122 (N_42122,N_39523,N_38293);
nand U42123 (N_42123,N_39317,N_39191);
xnor U42124 (N_42124,N_39223,N_37809);
or U42125 (N_42125,N_39406,N_39574);
and U42126 (N_42126,N_38938,N_37715);
nand U42127 (N_42127,N_37567,N_39966);
xor U42128 (N_42128,N_38315,N_39136);
and U42129 (N_42129,N_39723,N_39314);
or U42130 (N_42130,N_38602,N_39228);
nand U42131 (N_42131,N_39037,N_37885);
and U42132 (N_42132,N_37505,N_37610);
xnor U42133 (N_42133,N_39136,N_38782);
or U42134 (N_42134,N_39717,N_38588);
xor U42135 (N_42135,N_39335,N_39561);
nor U42136 (N_42136,N_37567,N_39688);
nand U42137 (N_42137,N_39168,N_37860);
nor U42138 (N_42138,N_38656,N_39326);
and U42139 (N_42139,N_38795,N_39952);
nor U42140 (N_42140,N_38166,N_38538);
or U42141 (N_42141,N_39556,N_39838);
and U42142 (N_42142,N_39715,N_38063);
and U42143 (N_42143,N_39672,N_39245);
xnor U42144 (N_42144,N_37937,N_39113);
and U42145 (N_42145,N_39065,N_39941);
or U42146 (N_42146,N_38255,N_38196);
and U42147 (N_42147,N_38858,N_37813);
and U42148 (N_42148,N_37557,N_38597);
or U42149 (N_42149,N_38790,N_39017);
nand U42150 (N_42150,N_39645,N_37807);
and U42151 (N_42151,N_38659,N_37824);
xnor U42152 (N_42152,N_38345,N_39313);
nor U42153 (N_42153,N_38881,N_38570);
nand U42154 (N_42154,N_37956,N_39632);
and U42155 (N_42155,N_38647,N_37602);
or U42156 (N_42156,N_39606,N_39097);
or U42157 (N_42157,N_38229,N_39167);
xnor U42158 (N_42158,N_37827,N_39087);
xnor U42159 (N_42159,N_38852,N_37758);
nand U42160 (N_42160,N_38532,N_39607);
or U42161 (N_42161,N_38055,N_38987);
nor U42162 (N_42162,N_38930,N_37825);
nand U42163 (N_42163,N_37974,N_39356);
or U42164 (N_42164,N_38141,N_39915);
or U42165 (N_42165,N_38942,N_38005);
xor U42166 (N_42166,N_39092,N_39500);
or U42167 (N_42167,N_39908,N_38643);
nand U42168 (N_42168,N_39926,N_39507);
nor U42169 (N_42169,N_38422,N_37987);
nor U42170 (N_42170,N_37841,N_38795);
xnor U42171 (N_42171,N_37671,N_38680);
and U42172 (N_42172,N_37798,N_39271);
nand U42173 (N_42173,N_39718,N_37983);
nand U42174 (N_42174,N_39272,N_39818);
and U42175 (N_42175,N_39742,N_38997);
and U42176 (N_42176,N_38831,N_38126);
or U42177 (N_42177,N_37682,N_38493);
or U42178 (N_42178,N_39839,N_39436);
nor U42179 (N_42179,N_39165,N_39490);
xnor U42180 (N_42180,N_39060,N_37888);
nor U42181 (N_42181,N_38563,N_39149);
or U42182 (N_42182,N_39717,N_38510);
nor U42183 (N_42183,N_38342,N_37552);
and U42184 (N_42184,N_38610,N_37634);
nand U42185 (N_42185,N_37920,N_39380);
nand U42186 (N_42186,N_39650,N_38080);
or U42187 (N_42187,N_37784,N_39216);
nand U42188 (N_42188,N_38184,N_37903);
or U42189 (N_42189,N_37930,N_38368);
nor U42190 (N_42190,N_38807,N_39114);
or U42191 (N_42191,N_38716,N_37926);
nand U42192 (N_42192,N_39707,N_38813);
and U42193 (N_42193,N_39843,N_39628);
nor U42194 (N_42194,N_39205,N_37730);
nor U42195 (N_42195,N_38882,N_38257);
xnor U42196 (N_42196,N_39210,N_38798);
nand U42197 (N_42197,N_37585,N_37976);
nor U42198 (N_42198,N_39743,N_38686);
xnor U42199 (N_42199,N_39785,N_38238);
nor U42200 (N_42200,N_38645,N_39820);
nand U42201 (N_42201,N_37636,N_39611);
nand U42202 (N_42202,N_39992,N_39494);
or U42203 (N_42203,N_37815,N_39243);
xnor U42204 (N_42204,N_37638,N_39728);
xnor U42205 (N_42205,N_39456,N_37728);
and U42206 (N_42206,N_38768,N_38562);
and U42207 (N_42207,N_38585,N_37815);
nor U42208 (N_42208,N_39097,N_39350);
xnor U42209 (N_42209,N_38004,N_37921);
or U42210 (N_42210,N_38512,N_39571);
and U42211 (N_42211,N_39899,N_38423);
xnor U42212 (N_42212,N_39238,N_39492);
or U42213 (N_42213,N_37729,N_39192);
or U42214 (N_42214,N_39120,N_39448);
nand U42215 (N_42215,N_39558,N_39413);
nor U42216 (N_42216,N_37940,N_38492);
xnor U42217 (N_42217,N_38079,N_39657);
or U42218 (N_42218,N_39592,N_39565);
xnor U42219 (N_42219,N_39433,N_39945);
nor U42220 (N_42220,N_38207,N_38211);
or U42221 (N_42221,N_37921,N_39511);
nand U42222 (N_42222,N_37822,N_39259);
nand U42223 (N_42223,N_38881,N_38710);
nand U42224 (N_42224,N_39894,N_37544);
xnor U42225 (N_42225,N_37537,N_38004);
nand U42226 (N_42226,N_38547,N_39324);
and U42227 (N_42227,N_39200,N_38438);
nand U42228 (N_42228,N_38103,N_37835);
nand U42229 (N_42229,N_38098,N_38692);
and U42230 (N_42230,N_37639,N_38650);
nand U42231 (N_42231,N_38972,N_37823);
and U42232 (N_42232,N_39623,N_38058);
nand U42233 (N_42233,N_39212,N_38086);
nand U42234 (N_42234,N_38222,N_39883);
xnor U42235 (N_42235,N_38461,N_38141);
or U42236 (N_42236,N_37938,N_39738);
and U42237 (N_42237,N_39131,N_38518);
nor U42238 (N_42238,N_39422,N_38327);
xor U42239 (N_42239,N_37520,N_38823);
and U42240 (N_42240,N_38673,N_38722);
xor U42241 (N_42241,N_39014,N_38389);
and U42242 (N_42242,N_39475,N_38370);
nor U42243 (N_42243,N_39250,N_39536);
and U42244 (N_42244,N_38590,N_37604);
nor U42245 (N_42245,N_38340,N_38071);
and U42246 (N_42246,N_38545,N_38631);
nor U42247 (N_42247,N_38976,N_38146);
xor U42248 (N_42248,N_39142,N_37755);
xor U42249 (N_42249,N_38741,N_37726);
or U42250 (N_42250,N_38776,N_39275);
xnor U42251 (N_42251,N_37767,N_37603);
and U42252 (N_42252,N_37680,N_38975);
and U42253 (N_42253,N_39066,N_37655);
nor U42254 (N_42254,N_37704,N_39623);
xor U42255 (N_42255,N_39473,N_38249);
xnor U42256 (N_42256,N_37877,N_39392);
nand U42257 (N_42257,N_38468,N_39690);
or U42258 (N_42258,N_38396,N_39623);
and U42259 (N_42259,N_38372,N_39287);
xnor U42260 (N_42260,N_39972,N_39537);
xnor U42261 (N_42261,N_37671,N_38900);
nor U42262 (N_42262,N_39093,N_39536);
nand U42263 (N_42263,N_39081,N_39474);
xor U42264 (N_42264,N_39505,N_38394);
xor U42265 (N_42265,N_37964,N_38586);
and U42266 (N_42266,N_39809,N_38340);
nand U42267 (N_42267,N_38445,N_39825);
or U42268 (N_42268,N_39869,N_39687);
xnor U42269 (N_42269,N_39891,N_37659);
nor U42270 (N_42270,N_38730,N_38482);
nor U42271 (N_42271,N_38709,N_39333);
or U42272 (N_42272,N_39869,N_38593);
xor U42273 (N_42273,N_37678,N_38909);
xnor U42274 (N_42274,N_38756,N_37711);
nor U42275 (N_42275,N_39912,N_38087);
xnor U42276 (N_42276,N_38146,N_38460);
nor U42277 (N_42277,N_39043,N_38590);
nand U42278 (N_42278,N_38881,N_38684);
or U42279 (N_42279,N_39122,N_39311);
xor U42280 (N_42280,N_38356,N_37907);
or U42281 (N_42281,N_39473,N_38106);
or U42282 (N_42282,N_39618,N_37546);
nor U42283 (N_42283,N_38789,N_38998);
or U42284 (N_42284,N_38197,N_38360);
or U42285 (N_42285,N_39312,N_39191);
and U42286 (N_42286,N_38617,N_39117);
nand U42287 (N_42287,N_38961,N_38867);
or U42288 (N_42288,N_37765,N_38503);
or U42289 (N_42289,N_39190,N_37675);
nor U42290 (N_42290,N_38726,N_39758);
and U42291 (N_42291,N_39531,N_38308);
or U42292 (N_42292,N_37663,N_39578);
nand U42293 (N_42293,N_39896,N_38687);
or U42294 (N_42294,N_38965,N_39542);
and U42295 (N_42295,N_39886,N_37877);
and U42296 (N_42296,N_39727,N_39468);
and U42297 (N_42297,N_39954,N_38813);
nor U42298 (N_42298,N_37913,N_39908);
and U42299 (N_42299,N_38860,N_38419);
or U42300 (N_42300,N_38139,N_37997);
and U42301 (N_42301,N_39986,N_39559);
nand U42302 (N_42302,N_38937,N_37642);
and U42303 (N_42303,N_37950,N_39559);
or U42304 (N_42304,N_38410,N_38033);
xnor U42305 (N_42305,N_38527,N_38559);
xor U42306 (N_42306,N_37900,N_39525);
xnor U42307 (N_42307,N_38942,N_39964);
and U42308 (N_42308,N_38359,N_39276);
nand U42309 (N_42309,N_39391,N_38620);
or U42310 (N_42310,N_39606,N_38286);
and U42311 (N_42311,N_38412,N_39368);
nand U42312 (N_42312,N_38704,N_38050);
nor U42313 (N_42313,N_39577,N_39377);
or U42314 (N_42314,N_39968,N_37740);
nor U42315 (N_42315,N_39489,N_39268);
or U42316 (N_42316,N_37670,N_38849);
nand U42317 (N_42317,N_37921,N_37654);
or U42318 (N_42318,N_38675,N_37977);
nand U42319 (N_42319,N_37614,N_39903);
nand U42320 (N_42320,N_39607,N_38279);
and U42321 (N_42321,N_38637,N_39135);
nor U42322 (N_42322,N_39270,N_38963);
nand U42323 (N_42323,N_38228,N_39047);
xor U42324 (N_42324,N_38904,N_39043);
nand U42325 (N_42325,N_37783,N_38979);
and U42326 (N_42326,N_38402,N_38155);
nor U42327 (N_42327,N_38054,N_38682);
or U42328 (N_42328,N_39901,N_39143);
xnor U42329 (N_42329,N_37738,N_37802);
or U42330 (N_42330,N_38474,N_39090);
or U42331 (N_42331,N_39340,N_39876);
xor U42332 (N_42332,N_39973,N_38628);
or U42333 (N_42333,N_39361,N_38077);
nor U42334 (N_42334,N_38646,N_38754);
nand U42335 (N_42335,N_38086,N_39659);
nand U42336 (N_42336,N_39269,N_39440);
or U42337 (N_42337,N_37681,N_39590);
xor U42338 (N_42338,N_38529,N_39158);
and U42339 (N_42339,N_39905,N_39889);
or U42340 (N_42340,N_38198,N_38358);
xor U42341 (N_42341,N_39071,N_38180);
xor U42342 (N_42342,N_38254,N_38114);
nand U42343 (N_42343,N_39259,N_39543);
nor U42344 (N_42344,N_39564,N_37535);
nand U42345 (N_42345,N_38329,N_38076);
or U42346 (N_42346,N_39138,N_38068);
nor U42347 (N_42347,N_39426,N_37841);
nand U42348 (N_42348,N_38641,N_39925);
nand U42349 (N_42349,N_37752,N_39274);
or U42350 (N_42350,N_38110,N_39013);
and U42351 (N_42351,N_38805,N_38331);
and U42352 (N_42352,N_38410,N_39715);
nor U42353 (N_42353,N_37776,N_38651);
or U42354 (N_42354,N_37587,N_38961);
nor U42355 (N_42355,N_37818,N_38096);
and U42356 (N_42356,N_37713,N_37623);
xor U42357 (N_42357,N_39871,N_38571);
and U42358 (N_42358,N_39249,N_38505);
and U42359 (N_42359,N_39147,N_38436);
and U42360 (N_42360,N_39594,N_38308);
xnor U42361 (N_42361,N_38487,N_39399);
and U42362 (N_42362,N_38093,N_39391);
nor U42363 (N_42363,N_38573,N_38765);
nand U42364 (N_42364,N_38408,N_39480);
and U42365 (N_42365,N_37943,N_38980);
or U42366 (N_42366,N_38461,N_37720);
nand U42367 (N_42367,N_39232,N_38486);
and U42368 (N_42368,N_37719,N_38138);
and U42369 (N_42369,N_39050,N_37723);
xnor U42370 (N_42370,N_38481,N_39285);
and U42371 (N_42371,N_37972,N_38107);
nand U42372 (N_42372,N_38536,N_39231);
nand U42373 (N_42373,N_39642,N_38641);
nand U42374 (N_42374,N_37625,N_38263);
and U42375 (N_42375,N_38915,N_39944);
or U42376 (N_42376,N_39248,N_39889);
nor U42377 (N_42377,N_39281,N_38183);
nor U42378 (N_42378,N_39735,N_37703);
or U42379 (N_42379,N_37503,N_38374);
nand U42380 (N_42380,N_38615,N_38238);
and U42381 (N_42381,N_39827,N_39647);
nor U42382 (N_42382,N_37800,N_38462);
and U42383 (N_42383,N_39348,N_39251);
nand U42384 (N_42384,N_37976,N_38104);
nand U42385 (N_42385,N_39265,N_39590);
nand U42386 (N_42386,N_38287,N_39814);
nand U42387 (N_42387,N_38476,N_39788);
xor U42388 (N_42388,N_38701,N_39099);
nand U42389 (N_42389,N_39739,N_39101);
and U42390 (N_42390,N_39983,N_39304);
nand U42391 (N_42391,N_38738,N_39528);
and U42392 (N_42392,N_38059,N_39623);
nor U42393 (N_42393,N_39442,N_39937);
nand U42394 (N_42394,N_38158,N_37828);
xnor U42395 (N_42395,N_38006,N_37776);
nand U42396 (N_42396,N_39212,N_38608);
xnor U42397 (N_42397,N_39959,N_38162);
xor U42398 (N_42398,N_39056,N_38842);
xor U42399 (N_42399,N_39933,N_38586);
or U42400 (N_42400,N_39398,N_38752);
nor U42401 (N_42401,N_38035,N_37769);
xor U42402 (N_42402,N_38947,N_39107);
or U42403 (N_42403,N_39533,N_38637);
and U42404 (N_42404,N_39918,N_37551);
nor U42405 (N_42405,N_39230,N_39456);
or U42406 (N_42406,N_37786,N_38750);
and U42407 (N_42407,N_37594,N_38786);
xnor U42408 (N_42408,N_39941,N_38066);
nand U42409 (N_42409,N_39964,N_38572);
nand U42410 (N_42410,N_39796,N_38451);
nand U42411 (N_42411,N_39245,N_39369);
xor U42412 (N_42412,N_39221,N_39666);
and U42413 (N_42413,N_38296,N_39997);
and U42414 (N_42414,N_37944,N_39083);
xnor U42415 (N_42415,N_37946,N_39995);
nand U42416 (N_42416,N_39009,N_37702);
nor U42417 (N_42417,N_39416,N_39277);
and U42418 (N_42418,N_37913,N_37517);
or U42419 (N_42419,N_39110,N_38343);
xor U42420 (N_42420,N_38312,N_38726);
nor U42421 (N_42421,N_38268,N_39593);
nand U42422 (N_42422,N_39123,N_38367);
and U42423 (N_42423,N_39716,N_37651);
xor U42424 (N_42424,N_39990,N_39784);
nand U42425 (N_42425,N_38342,N_38470);
and U42426 (N_42426,N_38650,N_37886);
nor U42427 (N_42427,N_38690,N_38513);
nand U42428 (N_42428,N_39953,N_38680);
and U42429 (N_42429,N_39217,N_38176);
nor U42430 (N_42430,N_38114,N_37981);
and U42431 (N_42431,N_38052,N_37762);
and U42432 (N_42432,N_38728,N_39257);
or U42433 (N_42433,N_39299,N_39928);
nor U42434 (N_42434,N_38921,N_39818);
nor U42435 (N_42435,N_37700,N_39877);
nand U42436 (N_42436,N_38828,N_39617);
xor U42437 (N_42437,N_37541,N_39190);
and U42438 (N_42438,N_39495,N_38168);
nand U42439 (N_42439,N_38562,N_39292);
xnor U42440 (N_42440,N_38095,N_37748);
or U42441 (N_42441,N_38295,N_39291);
nand U42442 (N_42442,N_39697,N_38718);
xor U42443 (N_42443,N_39634,N_37943);
xor U42444 (N_42444,N_39563,N_38762);
or U42445 (N_42445,N_38011,N_38818);
xnor U42446 (N_42446,N_39475,N_38084);
or U42447 (N_42447,N_39158,N_38909);
xor U42448 (N_42448,N_39187,N_39310);
or U42449 (N_42449,N_37545,N_38976);
xnor U42450 (N_42450,N_39505,N_37638);
nand U42451 (N_42451,N_38828,N_38881);
nand U42452 (N_42452,N_38520,N_38159);
or U42453 (N_42453,N_38802,N_38217);
xnor U42454 (N_42454,N_37983,N_38173);
nor U42455 (N_42455,N_38558,N_38027);
nor U42456 (N_42456,N_39915,N_38470);
xnor U42457 (N_42457,N_39550,N_39816);
or U42458 (N_42458,N_39757,N_39289);
or U42459 (N_42459,N_37982,N_38138);
xnor U42460 (N_42460,N_39796,N_38235);
nor U42461 (N_42461,N_38284,N_38521);
xor U42462 (N_42462,N_38193,N_39893);
or U42463 (N_42463,N_39685,N_38778);
or U42464 (N_42464,N_37678,N_38890);
nand U42465 (N_42465,N_37517,N_37682);
or U42466 (N_42466,N_38119,N_38884);
nor U42467 (N_42467,N_39282,N_38115);
nor U42468 (N_42468,N_39244,N_38711);
xnor U42469 (N_42469,N_37504,N_38549);
nor U42470 (N_42470,N_38693,N_38555);
nor U42471 (N_42471,N_38024,N_39074);
or U42472 (N_42472,N_39743,N_38615);
or U42473 (N_42473,N_38902,N_39118);
or U42474 (N_42474,N_38172,N_37604);
nand U42475 (N_42475,N_39134,N_38615);
nand U42476 (N_42476,N_39306,N_39209);
or U42477 (N_42477,N_38355,N_38217);
or U42478 (N_42478,N_37896,N_39312);
xor U42479 (N_42479,N_39385,N_38325);
nand U42480 (N_42480,N_38141,N_39860);
nor U42481 (N_42481,N_38983,N_39902);
and U42482 (N_42482,N_37743,N_39216);
xor U42483 (N_42483,N_38604,N_38583);
and U42484 (N_42484,N_39106,N_37662);
xnor U42485 (N_42485,N_38039,N_39068);
xnor U42486 (N_42486,N_37718,N_38765);
xnor U42487 (N_42487,N_37633,N_38668);
xor U42488 (N_42488,N_38887,N_39100);
and U42489 (N_42489,N_39639,N_38200);
nor U42490 (N_42490,N_37695,N_38270);
nand U42491 (N_42491,N_39639,N_38453);
nor U42492 (N_42492,N_37637,N_38561);
nand U42493 (N_42493,N_39295,N_38293);
and U42494 (N_42494,N_39152,N_38902);
nor U42495 (N_42495,N_37619,N_38956);
xor U42496 (N_42496,N_38461,N_38745);
or U42497 (N_42497,N_39901,N_39059);
nor U42498 (N_42498,N_38335,N_37994);
xor U42499 (N_42499,N_37823,N_39696);
nor U42500 (N_42500,N_41444,N_40029);
or U42501 (N_42501,N_42006,N_41804);
nand U42502 (N_42502,N_41726,N_41348);
xnor U42503 (N_42503,N_40562,N_40806);
or U42504 (N_42504,N_42384,N_41617);
nor U42505 (N_42505,N_42194,N_40566);
xor U42506 (N_42506,N_40018,N_40924);
and U42507 (N_42507,N_41578,N_42029);
nand U42508 (N_42508,N_40438,N_40898);
nor U42509 (N_42509,N_41093,N_41687);
nor U42510 (N_42510,N_42411,N_40249);
nand U42511 (N_42511,N_40041,N_41473);
nor U42512 (N_42512,N_41279,N_40916);
nand U42513 (N_42513,N_40414,N_41339);
and U42514 (N_42514,N_40514,N_41012);
or U42515 (N_42515,N_40919,N_40221);
or U42516 (N_42516,N_42340,N_41776);
nor U42517 (N_42517,N_42028,N_42446);
nor U42518 (N_42518,N_41501,N_40167);
nor U42519 (N_42519,N_40084,N_40853);
or U42520 (N_42520,N_40446,N_41358);
and U42521 (N_42521,N_41320,N_42138);
xnor U42522 (N_42522,N_41963,N_40386);
nand U42523 (N_42523,N_40954,N_41820);
and U42524 (N_42524,N_41765,N_41952);
xnor U42525 (N_42525,N_41427,N_40907);
or U42526 (N_42526,N_41483,N_40235);
xnor U42527 (N_42527,N_41833,N_41714);
nor U42528 (N_42528,N_42232,N_42053);
nor U42529 (N_42529,N_40594,N_40330);
nand U42530 (N_42530,N_40184,N_41899);
xnor U42531 (N_42531,N_40461,N_41156);
xnor U42532 (N_42532,N_40054,N_40050);
nor U42533 (N_42533,N_41318,N_41336);
or U42534 (N_42534,N_40344,N_41353);
nand U42535 (N_42535,N_40533,N_42247);
and U42536 (N_42536,N_40978,N_41625);
xnor U42537 (N_42537,N_42346,N_42464);
nand U42538 (N_42538,N_40708,N_40311);
nor U42539 (N_42539,N_42011,N_40232);
xnor U42540 (N_42540,N_40653,N_42465);
or U42541 (N_42541,N_40309,N_42491);
nor U42542 (N_42542,N_41744,N_41423);
or U42543 (N_42543,N_42067,N_40930);
xor U42544 (N_42544,N_41017,N_41253);
and U42545 (N_42545,N_40355,N_40038);
xor U42546 (N_42546,N_40039,N_42259);
nand U42547 (N_42547,N_41360,N_41314);
and U42548 (N_42548,N_41165,N_41872);
or U42549 (N_42549,N_40314,N_41231);
xnor U42550 (N_42550,N_42368,N_40748);
xor U42551 (N_42551,N_41095,N_42208);
nor U42552 (N_42552,N_41521,N_40664);
nor U42553 (N_42553,N_41303,N_40228);
nand U42554 (N_42554,N_41556,N_41595);
or U42555 (N_42555,N_42495,N_41527);
nor U42556 (N_42556,N_41582,N_41228);
and U42557 (N_42557,N_41875,N_41920);
xnor U42558 (N_42558,N_41539,N_42226);
or U42559 (N_42559,N_40250,N_42198);
and U42560 (N_42560,N_41665,N_40417);
and U42561 (N_42561,N_42039,N_41881);
and U42562 (N_42562,N_41964,N_40460);
nand U42563 (N_42563,N_41727,N_40540);
or U42564 (N_42564,N_40683,N_40493);
nor U42565 (N_42565,N_40879,N_40335);
nor U42566 (N_42566,N_42016,N_42468);
and U42567 (N_42567,N_41688,N_40921);
nor U42568 (N_42568,N_41293,N_41417);
or U42569 (N_42569,N_42275,N_40037);
nand U42570 (N_42570,N_42493,N_41045);
and U42571 (N_42571,N_41456,N_40139);
xnor U42572 (N_42572,N_40152,N_41808);
xor U42573 (N_42573,N_41131,N_40476);
and U42574 (N_42574,N_41201,N_41056);
and U42575 (N_42575,N_41402,N_41119);
nand U42576 (N_42576,N_41710,N_42474);
nand U42577 (N_42577,N_42216,N_42266);
nor U42578 (N_42578,N_42037,N_42410);
or U42579 (N_42579,N_42321,N_40056);
nand U42580 (N_42580,N_40302,N_42445);
xor U42581 (N_42581,N_41407,N_41758);
nand U42582 (N_42582,N_42412,N_40313);
and U42583 (N_42583,N_42088,N_41421);
nor U42584 (N_42584,N_41633,N_42407);
nand U42585 (N_42585,N_41437,N_42063);
or U42586 (N_42586,N_40797,N_42119);
and U42587 (N_42587,N_42424,N_40340);
nor U42588 (N_42588,N_40768,N_40948);
nor U42589 (N_42589,N_41666,N_42314);
or U42590 (N_42590,N_40905,N_41190);
nor U42591 (N_42591,N_40080,N_41500);
nand U42592 (N_42592,N_41817,N_42252);
and U42593 (N_42593,N_41123,N_42034);
or U42594 (N_42594,N_40960,N_40821);
nand U42595 (N_42595,N_40837,N_41340);
nor U42596 (N_42596,N_40223,N_41486);
nor U42597 (N_42597,N_40471,N_42455);
and U42598 (N_42598,N_40856,N_41815);
nor U42599 (N_42599,N_40716,N_40440);
xor U42600 (N_42600,N_41342,N_42284);
xnor U42601 (N_42601,N_42221,N_42361);
nand U42602 (N_42602,N_41007,N_41570);
or U42603 (N_42603,N_40858,N_40765);
xnor U42604 (N_42604,N_41040,N_41106);
nand U42605 (N_42605,N_41674,N_41929);
nand U42606 (N_42606,N_41529,N_40349);
and U42607 (N_42607,N_42038,N_40226);
or U42608 (N_42608,N_40961,N_42349);
nand U42609 (N_42609,N_41614,N_41142);
nor U42610 (N_42610,N_41632,N_42112);
xor U42611 (N_42611,N_41153,N_42440);
and U42612 (N_42612,N_41592,N_41036);
xnor U42613 (N_42613,N_40261,N_41404);
nand U42614 (N_42614,N_41781,N_40096);
and U42615 (N_42615,N_40774,N_42106);
nor U42616 (N_42616,N_42470,N_40178);
nand U42617 (N_42617,N_41917,N_40789);
xor U42618 (N_42618,N_40124,N_42336);
nor U42619 (N_42619,N_40483,N_40169);
nand U42620 (N_42620,N_42432,N_41946);
nor U42621 (N_42621,N_41626,N_41606);
or U42622 (N_42622,N_41124,N_40390);
nor U42623 (N_42623,N_42073,N_41168);
nand U42624 (N_42624,N_41835,N_40798);
or U42625 (N_42625,N_41728,N_42402);
nand U42626 (N_42626,N_41267,N_41459);
and U42627 (N_42627,N_41021,N_42327);
or U42628 (N_42628,N_40450,N_41465);
nor U42629 (N_42629,N_42125,N_40537);
or U42630 (N_42630,N_40265,N_40260);
nand U42631 (N_42631,N_42100,N_41514);
or U42632 (N_42632,N_41120,N_40772);
or U42633 (N_42633,N_41874,N_41957);
nand U42634 (N_42634,N_40757,N_42234);
xor U42635 (N_42635,N_41322,N_40962);
nor U42636 (N_42636,N_40865,N_42295);
nand U42637 (N_42637,N_41611,N_42204);
nor U42638 (N_42638,N_42017,N_42451);
xnor U42639 (N_42639,N_41082,N_41209);
xnor U42640 (N_42640,N_40183,N_41182);
xor U42641 (N_42641,N_40827,N_40936);
and U42642 (N_42642,N_41931,N_40076);
and U42643 (N_42643,N_41939,N_41559);
and U42644 (N_42644,N_41673,N_41535);
and U42645 (N_42645,N_40667,N_40530);
and U42646 (N_42646,N_41542,N_42105);
or U42647 (N_42647,N_40549,N_41911);
nand U42648 (N_42648,N_40792,N_42127);
nand U42649 (N_42649,N_40573,N_42307);
xnor U42650 (N_42650,N_41363,N_40326);
xnor U42651 (N_42651,N_41419,N_42399);
nand U42652 (N_42652,N_41669,N_40724);
nand U42653 (N_42653,N_41934,N_40477);
nand U42654 (N_42654,N_40803,N_41885);
and U42655 (N_42655,N_41230,N_40244);
nor U42656 (N_42656,N_41395,N_41802);
nand U42657 (N_42657,N_41172,N_42463);
nor U42658 (N_42658,N_40788,N_40331);
nor U42659 (N_42659,N_41111,N_41510);
xor U42660 (N_42660,N_41430,N_40648);
and U42661 (N_42661,N_40563,N_41850);
nand U42662 (N_42662,N_41830,N_42081);
or U42663 (N_42663,N_40132,N_41059);
or U42664 (N_42664,N_41143,N_40603);
and U42665 (N_42665,N_42027,N_41273);
nor U42666 (N_42666,N_41656,N_41265);
nor U42667 (N_42667,N_42183,N_40310);
nand U42668 (N_42668,N_40997,N_40551);
and U42669 (N_42669,N_40149,N_42049);
nor U42670 (N_42670,N_42182,N_40306);
and U42671 (N_42671,N_41431,N_40052);
or U42672 (N_42672,N_41378,N_41426);
nor U42673 (N_42673,N_41927,N_41855);
xnor U42674 (N_42674,N_42084,N_41063);
nor U42675 (N_42675,N_42083,N_42090);
or U42676 (N_42676,N_40177,N_40951);
or U42677 (N_42677,N_40763,N_41335);
or U42678 (N_42678,N_40336,N_41118);
nand U42679 (N_42679,N_41742,N_41275);
xor U42680 (N_42680,N_41264,N_40318);
nand U42681 (N_42681,N_40148,N_40475);
nand U42682 (N_42682,N_41174,N_40108);
nand U42683 (N_42683,N_41411,N_42184);
or U42684 (N_42684,N_42209,N_41296);
xnor U42685 (N_42685,N_40248,N_42370);
or U42686 (N_42686,N_41568,N_42270);
nor U42687 (N_42687,N_42235,N_41104);
and U42688 (N_42688,N_42020,N_40732);
nor U42689 (N_42689,N_41821,N_40363);
nor U42690 (N_42690,N_42010,N_40393);
nand U42691 (N_42691,N_40628,N_41607);
and U42692 (N_42692,N_41079,N_41720);
xor U42693 (N_42693,N_41986,N_41774);
nor U42694 (N_42694,N_41098,N_41311);
or U42695 (N_42695,N_41893,N_42434);
and U42696 (N_42696,N_41943,N_41278);
nor U42697 (N_42697,N_41838,N_40238);
and U42698 (N_42698,N_40125,N_41246);
nand U42699 (N_42699,N_41281,N_41824);
or U42700 (N_42700,N_41133,N_40230);
xor U42701 (N_42701,N_40854,N_41724);
or U42702 (N_42702,N_42363,N_40728);
and U42703 (N_42703,N_42256,N_41947);
xor U42704 (N_42704,N_41132,N_42196);
nand U42705 (N_42705,N_41244,N_41889);
xnor U42706 (N_42706,N_40947,N_41725);
xor U42707 (N_42707,N_42394,N_41088);
or U42708 (N_42708,N_41642,N_41506);
xor U42709 (N_42709,N_42276,N_41756);
xnor U42710 (N_42710,N_42002,N_42312);
nor U42711 (N_42711,N_42228,N_42348);
xor U42712 (N_42712,N_42462,N_41741);
nor U42713 (N_42713,N_41643,N_42378);
xor U42714 (N_42714,N_42079,N_40672);
nor U42715 (N_42715,N_40432,N_40053);
nor U42716 (N_42716,N_41574,N_42390);
xnor U42717 (N_42717,N_40480,N_41519);
xor U42718 (N_42718,N_40329,N_42335);
nor U42719 (N_42719,N_40985,N_41385);
and U42720 (N_42720,N_41645,N_42126);
nor U42721 (N_42721,N_40299,N_41676);
xnor U42722 (N_42722,N_40459,N_40861);
or U42723 (N_42723,N_42377,N_41247);
and U42724 (N_42724,N_40602,N_41452);
xor U42725 (N_42725,N_41967,N_40946);
xor U42726 (N_42726,N_41200,N_42397);
and U42727 (N_42727,N_42143,N_40101);
nor U42728 (N_42728,N_41677,N_40590);
nor U42729 (N_42729,N_40333,N_40506);
xor U42730 (N_42730,N_41461,N_41609);
or U42731 (N_42731,N_40544,N_41579);
or U42732 (N_42732,N_40419,N_42164);
nand U42733 (N_42733,N_41409,N_41705);
xnor U42734 (N_42734,N_40599,N_40776);
or U42735 (N_42735,N_40753,N_42122);
nand U42736 (N_42736,N_42166,N_42117);
nand U42737 (N_42737,N_40731,N_40676);
and U42738 (N_42738,N_42482,N_41738);
xor U42739 (N_42739,N_40661,N_40980);
or U42740 (N_42740,N_41865,N_40192);
nand U42741 (N_42741,N_42167,N_40146);
and U42742 (N_42742,N_41167,N_40147);
and U42743 (N_42743,N_40744,N_42129);
nand U42744 (N_42744,N_41186,N_42219);
nand U42745 (N_42745,N_40224,N_41584);
nor U42746 (N_42746,N_41152,N_42007);
xnor U42747 (N_42747,N_42302,N_40212);
and U42748 (N_42748,N_41962,N_40927);
nor U42749 (N_42749,N_40567,N_42444);
xnor U42750 (N_42750,N_40103,N_42294);
or U42751 (N_42751,N_40973,N_41715);
and U42752 (N_42752,N_41467,N_42174);
nand U42753 (N_42753,N_40649,N_40348);
nand U42754 (N_42754,N_42169,N_41690);
and U42755 (N_42755,N_41729,N_42347);
and U42756 (N_42756,N_40441,N_41619);
or U42757 (N_42757,N_41896,N_41085);
xor U42758 (N_42758,N_40814,N_40523);
xor U42759 (N_42759,N_40819,N_41572);
and U42760 (N_42760,N_41475,N_40091);
or U42761 (N_42761,N_40379,N_40781);
xnor U42762 (N_42762,N_41793,N_40892);
and U42763 (N_42763,N_40357,N_40399);
nand U42764 (N_42764,N_41050,N_40654);
or U42765 (N_42765,N_41347,N_41890);
and U42766 (N_42766,N_40082,N_40397);
or U42767 (N_42767,N_41832,N_40580);
or U42768 (N_42768,N_42113,N_42099);
nor U42769 (N_42769,N_41206,N_41463);
nand U42770 (N_42770,N_40154,N_41258);
xnor U42771 (N_42771,N_41637,N_40527);
xnor U42772 (N_42772,N_41863,N_41357);
and U42773 (N_42773,N_41003,N_41408);
nand U42774 (N_42774,N_40209,N_42050);
and U42775 (N_42775,N_41438,N_42210);
or U42776 (N_42776,N_41531,N_41700);
xnor U42777 (N_42777,N_40293,N_41026);
and U42778 (N_42778,N_41775,N_41768);
and U42779 (N_42779,N_41594,N_41518);
nor U42780 (N_42780,N_42065,N_40011);
xor U42781 (N_42781,N_41051,N_40779);
nand U42782 (N_42782,N_40904,N_40449);
nor U42783 (N_42783,N_41921,N_40682);
xnor U42784 (N_42784,N_42150,N_42396);
and U42785 (N_42785,N_40714,N_40877);
or U42786 (N_42786,N_41827,N_40982);
or U42787 (N_42787,N_42323,N_42452);
xor U42788 (N_42788,N_40785,N_40750);
xor U42789 (N_42789,N_40118,N_42236);
xnor U42790 (N_42790,N_40616,N_42393);
xnor U42791 (N_42791,N_40504,N_42439);
xor U42792 (N_42792,N_41540,N_40833);
xor U42793 (N_42793,N_41383,N_40994);
and U42794 (N_42794,N_41976,N_40914);
nand U42795 (N_42795,N_42499,N_40706);
or U42796 (N_42796,N_40470,N_41065);
nor U42797 (N_42797,N_41573,N_42492);
nor U42798 (N_42798,N_42200,N_42203);
nand U42799 (N_42799,N_40862,N_41101);
nand U42800 (N_42800,N_42004,N_40083);
nand U42801 (N_42801,N_42304,N_41207);
and U42802 (N_42802,N_40105,N_41703);
nor U42803 (N_42803,N_40134,N_42199);
nor U42804 (N_42804,N_41166,N_40660);
or U42805 (N_42805,N_41499,N_41307);
nand U42806 (N_42806,N_40911,N_40025);
and U42807 (N_42807,N_41956,N_41325);
and U42808 (N_42808,N_41718,N_41203);
nor U42809 (N_42809,N_41707,N_42391);
and U42810 (N_42810,N_42218,N_41750);
nand U42811 (N_42811,N_40687,N_42369);
or U42812 (N_42812,N_40621,N_41600);
nor U42813 (N_42813,N_40231,N_40722);
nand U42814 (N_42814,N_40220,N_42450);
nand U42815 (N_42815,N_40155,N_41842);
or U42816 (N_42816,N_41041,N_40233);
xnor U42817 (N_42817,N_42395,N_40063);
xor U42818 (N_42818,N_40909,N_41128);
nand U42819 (N_42819,N_40635,N_40456);
xnor U42820 (N_42820,N_42147,N_40636);
xor U42821 (N_42821,N_42414,N_41942);
and U42822 (N_42822,N_42461,N_42477);
and U42823 (N_42823,N_41678,N_41317);
xor U42824 (N_42824,N_42457,N_40085);
or U42825 (N_42825,N_40113,N_41077);
and U42826 (N_42826,N_40388,N_40161);
nand U42827 (N_42827,N_41066,N_41269);
nand U42828 (N_42828,N_40607,N_41599);
nor U42829 (N_42829,N_41616,N_40019);
or U42830 (N_42830,N_42193,N_40920);
or U42831 (N_42831,N_42280,N_40141);
nand U42832 (N_42832,N_40888,N_40342);
or U42833 (N_42833,N_40702,N_40109);
xnor U42834 (N_42834,N_40887,N_42315);
nor U42835 (N_42835,N_40696,N_40135);
nand U42836 (N_42836,N_42253,N_40385);
and U42837 (N_42837,N_42262,N_42139);
nand U42838 (N_42838,N_41796,N_42466);
or U42839 (N_42839,N_42403,N_40572);
nand U42840 (N_42840,N_40592,N_41277);
or U42841 (N_42841,N_41990,N_41525);
nor U42842 (N_42842,N_42287,N_40780);
or U42843 (N_42843,N_41966,N_40705);
xnor U42844 (N_42844,N_41401,N_40035);
or U42845 (N_42845,N_41257,N_42405);
nor U42846 (N_42846,N_41495,N_41447);
nor U42847 (N_42847,N_40402,N_42429);
or U42848 (N_42848,N_41301,N_42163);
xnor U42849 (N_42849,N_40413,N_40274);
nor U42850 (N_42850,N_40875,N_40401);
or U42851 (N_42851,N_40087,N_40384);
nor U42852 (N_42852,N_41555,N_40110);
nand U42853 (N_42853,N_40014,N_41091);
and U42854 (N_42854,N_42350,N_40194);
and U42855 (N_42855,N_40832,N_41912);
nand U42856 (N_42856,N_40938,N_41014);
nor U42857 (N_42857,N_40458,N_40639);
or U42858 (N_42858,N_40000,N_40346);
or U42859 (N_42859,N_41816,N_41323);
nor U42860 (N_42860,N_40894,N_41693);
or U42861 (N_42861,N_41538,N_41588);
or U42862 (N_42862,N_40902,N_41073);
xor U42863 (N_42863,N_41226,N_41978);
or U42864 (N_42864,N_41552,N_42014);
and U42865 (N_42865,N_41762,N_42267);
nor U42866 (N_42866,N_42291,N_41918);
or U42867 (N_42867,N_40009,N_41659);
or U42868 (N_42868,N_41205,N_40584);
nand U42869 (N_42869,N_40433,N_40764);
nor U42870 (N_42870,N_41234,N_40574);
or U42871 (N_42871,N_40322,N_40350);
nor U42872 (N_42872,N_42033,N_41685);
or U42873 (N_42873,N_41694,N_41869);
xnor U42874 (N_42874,N_42435,N_40766);
nor U42875 (N_42875,N_40984,N_41736);
and U42876 (N_42876,N_40822,N_42175);
and U42877 (N_42877,N_40734,N_41405);
nand U42878 (N_42878,N_41851,N_40266);
nor U42879 (N_42879,N_40496,N_41458);
and U42880 (N_42880,N_41806,N_42292);
and U42881 (N_42881,N_41446,N_41297);
and U42882 (N_42882,N_42289,N_41549);
and U42883 (N_42883,N_42286,N_40880);
nor U42884 (N_42884,N_41284,N_42121);
nand U42885 (N_42885,N_40452,N_40756);
nor U42886 (N_42886,N_41581,N_42191);
nor U42887 (N_42887,N_42171,N_42015);
nor U42888 (N_42888,N_40626,N_42398);
and U42889 (N_42889,N_41936,N_40860);
nand U42890 (N_42890,N_41882,N_41748);
and U42891 (N_42891,N_41382,N_40680);
nor U42892 (N_42892,N_41433,N_41670);
and U42893 (N_42893,N_40615,N_40102);
nor U42894 (N_42894,N_41585,N_42064);
nor U42895 (N_42895,N_41196,N_40881);
nand U42896 (N_42896,N_40501,N_41454);
xnor U42897 (N_42897,N_41328,N_40424);
nor U42898 (N_42898,N_41177,N_42264);
nand U42899 (N_42899,N_41248,N_41298);
and U42900 (N_42900,N_40842,N_41413);
and U42901 (N_42901,N_42421,N_41173);
and U42902 (N_42902,N_42258,N_41286);
nor U42903 (N_42903,N_41792,N_40193);
and U42904 (N_42904,N_42485,N_41951);
xnor U42905 (N_42905,N_41508,N_41941);
nor U42906 (N_42906,N_41711,N_41873);
and U42907 (N_42907,N_40629,N_40488);
nand U42908 (N_42908,N_41880,N_41398);
and U42909 (N_42909,N_40442,N_42447);
and U42910 (N_42910,N_42104,N_40730);
and U42911 (N_42911,N_42288,N_40694);
nand U42912 (N_42912,N_40871,N_41735);
nor U42913 (N_42913,N_41960,N_41862);
or U42914 (N_42914,N_42358,N_41811);
xnor U42915 (N_42915,N_40679,N_41983);
or U42916 (N_42916,N_42072,N_40640);
xor U42917 (N_42917,N_41497,N_41300);
nand U42918 (N_42918,N_42145,N_40737);
nand U42919 (N_42919,N_41341,N_41108);
or U42920 (N_42920,N_40367,N_41054);
xnor U42921 (N_42921,N_41753,N_40754);
and U42922 (N_42922,N_41192,N_40246);
and U42923 (N_42923,N_41959,N_41105);
xnor U42924 (N_42924,N_41795,N_41590);
or U42925 (N_42925,N_42030,N_40013);
and U42926 (N_42926,N_40651,N_40435);
nor U42927 (N_42927,N_41148,N_40777);
and U42928 (N_42928,N_40499,N_41681);
nor U42929 (N_42929,N_42488,N_42459);
nand U42930 (N_42930,N_42362,N_40280);
and U42931 (N_42931,N_41137,N_42144);
nor U42932 (N_42932,N_41373,N_42195);
or U42933 (N_42933,N_41680,N_40188);
and U42934 (N_42934,N_41330,N_42415);
or U42935 (N_42935,N_41530,N_40351);
nand U42936 (N_42936,N_42352,N_41557);
or U42937 (N_42937,N_40074,N_41919);
and U42938 (N_42938,N_41615,N_42243);
nand U42939 (N_42939,N_42159,N_42331);
and U42940 (N_42940,N_41502,N_41777);
xor U42941 (N_42941,N_41602,N_41212);
or U42942 (N_42942,N_40300,N_40334);
xnor U42943 (N_42943,N_40116,N_40404);
nor U42944 (N_42944,N_41866,N_41164);
xor U42945 (N_42945,N_40075,N_42176);
or U42946 (N_42946,N_41217,N_40568);
nor U42947 (N_42947,N_41432,N_41895);
xnor U42948 (N_42948,N_40620,N_40817);
nand U42949 (N_42949,N_40752,N_41958);
nand U42950 (N_42950,N_40498,N_41136);
nand U42951 (N_42951,N_40186,N_40173);
or U42952 (N_42952,N_40931,N_42009);
nand U42953 (N_42953,N_40126,N_40278);
nor U42954 (N_42954,N_41224,N_40673);
xnor U42955 (N_42955,N_40298,N_40992);
and U42956 (N_42956,N_42300,N_41886);
nand U42957 (N_42957,N_41580,N_40067);
xnor U42958 (N_42958,N_41695,N_40794);
nand U42959 (N_42959,N_40923,N_41587);
nor U42960 (N_42960,N_42242,N_40319);
nand U42961 (N_42961,N_42035,N_40117);
nor U42962 (N_42962,N_41980,N_41251);
xnor U42963 (N_42963,N_41825,N_40988);
and U42964 (N_42964,N_40203,N_40870);
or U42965 (N_42965,N_40699,N_41276);
and U42966 (N_42966,N_42116,N_41075);
and U42967 (N_42967,N_41179,N_41770);
nand U42968 (N_42968,N_42071,N_42324);
nor U42969 (N_42969,N_40006,N_42371);
nand U42970 (N_42970,N_42325,N_42436);
xor U42971 (N_42971,N_41110,N_40421);
and U42972 (N_42972,N_40910,N_42168);
or U42973 (N_42973,N_41757,N_41836);
nor U42974 (N_42974,N_41996,N_40239);
nand U42975 (N_42975,N_42149,N_40229);
nor U42976 (N_42976,N_42305,N_40205);
xor U42977 (N_42977,N_40542,N_41139);
or U42978 (N_42978,N_40127,N_42416);
or U42979 (N_42979,N_40935,N_41147);
nand U42980 (N_42980,N_40507,N_40423);
nand U42981 (N_42981,N_40729,N_40809);
nand U42982 (N_42982,N_41924,N_42472);
or U42983 (N_42983,N_42093,N_41352);
or U42984 (N_42984,N_40825,N_40849);
xor U42985 (N_42985,N_40739,N_41564);
nor U42986 (N_42986,N_41517,N_42301);
nand U42987 (N_42987,N_42332,N_40159);
xor U42988 (N_42988,N_41789,N_40267);
or U42989 (N_42989,N_41553,N_41708);
nand U42990 (N_42990,N_40328,N_42443);
nand U42991 (N_42991,N_40150,N_41998);
or U42992 (N_42992,N_41161,N_40622);
nand U42993 (N_42993,N_42045,N_41365);
nand U42994 (N_42994,N_40122,N_40608);
nor U42995 (N_42995,N_40610,N_40200);
or U42996 (N_42996,N_41810,N_41788);
nand U42997 (N_42997,N_42047,N_42473);
nand U42998 (N_42998,N_40878,N_40465);
nand U42999 (N_42999,N_41127,N_41117);
xnor U43000 (N_43000,N_42356,N_42026);
nor U43001 (N_43001,N_40347,N_41638);
or U43002 (N_43002,N_41879,N_42357);
nor U43003 (N_43003,N_41261,N_41070);
or U43004 (N_43004,N_41387,N_41989);
or U43005 (N_43005,N_42478,N_40307);
and U43006 (N_43006,N_40003,N_41049);
nand U43007 (N_43007,N_42320,N_41222);
or U43008 (N_43008,N_41785,N_41664);
and U43009 (N_43009,N_41283,N_41441);
nor U43010 (N_43010,N_41018,N_40570);
nand U43011 (N_43011,N_40895,N_40040);
nand U43012 (N_43012,N_40813,N_41513);
xnor U43013 (N_43013,N_41979,N_40364);
xnor U43014 (N_43014,N_40451,N_40426);
nor U43015 (N_43015,N_41002,N_40297);
xnor U43016 (N_43016,N_42409,N_40271);
and U43017 (N_43017,N_40093,N_40073);
nand U43018 (N_43018,N_40048,N_42186);
nor U43019 (N_43019,N_40944,N_41369);
or U43020 (N_43020,N_41107,N_42068);
and U43021 (N_43021,N_40755,N_40681);
xnor U43022 (N_43022,N_42261,N_41791);
and U43023 (N_43023,N_40826,N_40133);
nand U43024 (N_43024,N_40295,N_41183);
xnor U43025 (N_43025,N_42215,N_41653);
and U43026 (N_43026,N_41618,N_40374);
nand U43027 (N_43027,N_41255,N_42018);
nor U43028 (N_43028,N_42433,N_41443);
and U43029 (N_43029,N_41543,N_42469);
nor U43030 (N_43030,N_41894,N_41930);
and U43031 (N_43031,N_42343,N_41932);
or U43032 (N_43032,N_40976,N_42322);
nand U43033 (N_43033,N_40520,N_42230);
nor U43034 (N_43034,N_42279,N_40535);
and U43035 (N_43035,N_41968,N_40955);
or U43036 (N_43036,N_42339,N_41861);
xnor U43037 (N_43037,N_42202,N_41309);
nand U43038 (N_43038,N_40671,N_41146);
nand U43039 (N_43039,N_40528,N_41324);
xnor U43040 (N_43040,N_41523,N_40829);
or U43041 (N_43041,N_41747,N_41194);
and U43042 (N_43042,N_40596,N_42086);
and U43043 (N_43043,N_41099,N_40835);
and U43044 (N_43044,N_40064,N_40987);
xnor U43045 (N_43045,N_41982,N_41610);
xor U43046 (N_43046,N_40691,N_41266);
and U43047 (N_43047,N_40698,N_40160);
nand U43048 (N_43048,N_41884,N_41233);
or U43049 (N_43049,N_42254,N_41494);
nand U43050 (N_43050,N_40587,N_40720);
nor U43051 (N_43051,N_40359,N_40381);
xnor U43052 (N_43052,N_40721,N_42227);
or U43053 (N_43053,N_42299,N_40263);
nor U43054 (N_43054,N_40352,N_40700);
xor U43055 (N_43055,N_40872,N_40508);
nor U43056 (N_43056,N_41274,N_41566);
nand U43057 (N_43057,N_40536,N_40556);
and U43058 (N_43058,N_40304,N_41445);
and U43059 (N_43059,N_41987,N_41280);
or U43060 (N_43060,N_42298,N_41565);
xor U43061 (N_43061,N_41096,N_40142);
and U43062 (N_43062,N_40941,N_40585);
xor U43063 (N_43063,N_40198,N_41151);
xor U43064 (N_43064,N_40028,N_40791);
nand U43065 (N_43065,N_40595,N_41381);
and U43066 (N_43066,N_40020,N_42238);
or U43067 (N_43067,N_42330,N_40023);
or U43068 (N_43068,N_42096,N_40343);
or U43069 (N_43069,N_41702,N_41532);
nor U43070 (N_43070,N_42179,N_42054);
nor U43071 (N_43071,N_40005,N_41425);
nand U43072 (N_43072,N_40180,N_41299);
nor U43073 (N_43073,N_40863,N_41622);
or U43074 (N_43074,N_40068,N_41295);
xor U43075 (N_43075,N_42479,N_41229);
or U43076 (N_43076,N_40467,N_41292);
xor U43077 (N_43077,N_41709,N_40655);
and U43078 (N_43078,N_41086,N_41472);
and U43079 (N_43079,N_40623,N_41754);
and U43080 (N_43080,N_40338,N_40358);
or U43081 (N_43081,N_41460,N_40004);
or U43082 (N_43082,N_41985,N_40360);
xnor U43083 (N_43083,N_40016,N_42313);
xnor U43084 (N_43084,N_41094,N_40517);
or U43085 (N_43085,N_42036,N_41149);
xnor U43086 (N_43086,N_40007,N_40718);
and U43087 (N_43087,N_42360,N_40939);
or U43088 (N_43088,N_42153,N_41406);
xnor U43089 (N_43089,N_40253,N_41024);
and U43090 (N_43090,N_41944,N_40824);
or U43091 (N_43091,N_41355,N_42353);
nor U43092 (N_43092,N_41883,N_40922);
nor U43093 (N_43093,N_40519,N_41620);
nand U43094 (N_43094,N_40487,N_40908);
and U43095 (N_43095,N_40883,N_41033);
or U43096 (N_43096,N_41926,N_42044);
xnor U43097 (N_43097,N_40104,N_41623);
nand U43098 (N_43098,N_40554,N_40378);
nor U43099 (N_43099,N_40571,N_42087);
and U43100 (N_43100,N_40784,N_40787);
xnor U43101 (N_43101,N_40474,N_40320);
xor U43102 (N_43102,N_42115,N_41420);
nand U43103 (N_43103,N_41981,N_40709);
nor U43104 (N_43104,N_42097,N_41717);
xnor U43105 (N_43105,N_40092,N_40024);
and U43106 (N_43106,N_41558,N_40816);
xor U43107 (N_43107,N_40071,N_40371);
or U43108 (N_43108,N_40240,N_40131);
nand U43109 (N_43109,N_41937,N_42379);
or U43110 (N_43110,N_42374,N_40315);
xnor U43111 (N_43111,N_40650,N_41682);
xnor U43112 (N_43112,N_40502,N_42310);
nor U43113 (N_43113,N_42245,N_41635);
and U43114 (N_43114,N_40407,N_40268);
xnor U43115 (N_43115,N_40889,N_41701);
nand U43116 (N_43116,N_42205,N_40066);
and U43117 (N_43117,N_41121,N_41503);
nand U43118 (N_43118,N_41034,N_40601);
nand U43119 (N_43119,N_40218,N_41822);
nand U43120 (N_43120,N_42181,N_40538);
xor U43121 (N_43121,N_40675,N_40415);
nand U43122 (N_43122,N_42487,N_41170);
and U43123 (N_43123,N_41215,N_40369);
or U43124 (N_43124,N_40400,N_41515);
xnor U43125 (N_43125,N_41903,N_42022);
nor U43126 (N_43126,N_40942,N_40468);
nand U43127 (N_43127,N_41282,N_41953);
or U43128 (N_43128,N_40055,N_41739);
nand U43129 (N_43129,N_41800,N_40531);
nor U43130 (N_43130,N_40264,N_40505);
nand U43131 (N_43131,N_40632,N_40525);
nand U43132 (N_43132,N_41629,N_41593);
xor U43133 (N_43133,N_42160,N_42388);
nand U43134 (N_43134,N_40582,N_42005);
and U43135 (N_43135,N_40581,N_41256);
nand U43136 (N_43136,N_40996,N_42052);
nand U43137 (N_43137,N_42185,N_41468);
or U43138 (N_43138,N_40543,N_40513);
or U43139 (N_43139,N_41740,N_42490);
and U43140 (N_43140,N_42486,N_42158);
xnor U43141 (N_43141,N_42311,N_40642);
xor U43142 (N_43142,N_40839,N_42082);
and U43143 (N_43143,N_40715,N_40859);
nand U43144 (N_43144,N_42366,N_40738);
and U43145 (N_43145,N_40245,N_41436);
nor U43146 (N_43146,N_42013,N_40588);
nor U43147 (N_43147,N_41745,N_41178);
or U43148 (N_43148,N_41773,N_41723);
or U43149 (N_43149,N_40900,N_40560);
nand U43150 (N_43150,N_41954,N_40222);
xor U43151 (N_43151,N_40725,N_41772);
nor U43152 (N_43152,N_40106,N_40312);
nand U43153 (N_43153,N_41654,N_42272);
or U43154 (N_43154,N_40929,N_41991);
xnor U43155 (N_43155,N_41871,N_42293);
and U43156 (N_43156,N_41332,N_40002);
nand U43157 (N_43157,N_42003,N_40325);
nor U43158 (N_43158,N_40641,N_40665);
nand U43159 (N_43159,N_41380,N_41853);
or U43160 (N_43160,N_42173,N_40550);
nor U43161 (N_43161,N_42091,N_40899);
or U43162 (N_43162,N_40368,N_41846);
nor U43163 (N_43163,N_40285,N_41828);
or U43164 (N_43164,N_42103,N_40795);
xor U43165 (N_43165,N_40678,N_42372);
nor U43166 (N_43166,N_41520,N_42448);
nand U43167 (N_43167,N_42380,N_41219);
xnor U43168 (N_43168,N_41933,N_41922);
or U43169 (N_43169,N_40276,N_41092);
xnor U43170 (N_43170,N_40617,N_40604);
nor U43171 (N_43171,N_40123,N_41589);
xnor U43172 (N_43172,N_40674,N_42076);
and U43173 (N_43173,N_42207,N_41906);
or U43174 (N_43174,N_40042,N_40296);
xnor U43175 (N_43175,N_40612,N_40012);
nand U43176 (N_43176,N_40812,N_40197);
and U43177 (N_43177,N_41076,N_42430);
xnor U43178 (N_43178,N_41025,N_41449);
nor U43179 (N_43179,N_40855,N_41412);
nand U43180 (N_43180,N_40989,N_40383);
nor U43181 (N_43181,N_41892,N_40624);
xnor U43182 (N_43182,N_40234,N_42094);
nor U43183 (N_43183,N_40707,N_40983);
nand U43184 (N_43184,N_40445,N_40796);
and U43185 (N_43185,N_41852,N_41392);
nor U43186 (N_43186,N_41057,N_41371);
and U43187 (N_43187,N_40521,N_41344);
nand U43188 (N_43188,N_40852,N_40583);
nor U43189 (N_43189,N_41887,N_41254);
nand U43190 (N_43190,N_42146,N_41291);
xor U43191 (N_43191,N_42265,N_41062);
or U43192 (N_43192,N_40974,N_40723);
nor U43193 (N_43193,N_42229,N_41512);
xor U43194 (N_43194,N_40500,N_40166);
xnor U43195 (N_43195,N_40434,N_40256);
or U43196 (N_43196,N_41290,N_42032);
nand U43197 (N_43197,N_42180,N_40395);
xnor U43198 (N_43198,N_40657,N_40840);
and U43199 (N_43199,N_42211,N_40416);
nand U43200 (N_43200,N_42417,N_40077);
nor U43201 (N_43201,N_40771,N_41157);
and U43202 (N_43202,N_40986,N_41268);
or U43203 (N_43203,N_41994,N_42189);
xor U43204 (N_43204,N_42308,N_40422);
nand U43205 (N_43205,N_41948,N_41083);
xor U43206 (N_43206,N_42237,N_42225);
xnor U43207 (N_43207,N_40630,N_40156);
xor U43208 (N_43208,N_40060,N_41771);
or U43209 (N_43209,N_42136,N_40569);
and U43210 (N_43210,N_40666,N_41679);
nor U43211 (N_43211,N_41089,N_42297);
nand U43212 (N_43212,N_40686,N_41271);
nand U43213 (N_43213,N_41158,N_40008);
xor U43214 (N_43214,N_42019,N_40743);
xor U43215 (N_43215,N_40546,N_41193);
and U43216 (N_43216,N_40703,N_42107);
or U43217 (N_43217,N_40712,N_40217);
or U43218 (N_43218,N_40130,N_41238);
and U43219 (N_43219,N_40637,N_40409);
nor U43220 (N_43220,N_41250,N_40614);
nand U43221 (N_43221,N_42213,N_41812);
and U43222 (N_43222,N_41915,N_42244);
xor U43223 (N_43223,N_41969,N_40945);
and U43224 (N_43224,N_40157,N_40999);
xnor U43225 (N_43225,N_40685,N_41305);
or U43226 (N_43226,N_40726,N_40219);
and U43227 (N_43227,N_42128,N_40032);
or U43228 (N_43228,N_40270,N_42161);
xor U43229 (N_43229,N_41176,N_40586);
xor U43230 (N_43230,N_42001,N_41048);
nor U43231 (N_43231,N_41109,N_41011);
nor U43232 (N_43232,N_40492,N_41346);
or U43233 (N_43233,N_41498,N_41496);
nor U43234 (N_43234,N_40933,N_42427);
nand U43235 (N_43235,N_40204,N_40589);
nor U43236 (N_43236,N_41651,N_41097);
or U43237 (N_43237,N_41187,N_40557);
nand U43238 (N_43238,N_41029,N_41090);
and U43239 (N_43239,N_40489,N_41016);
or U43240 (N_43240,N_41663,N_41337);
nand U43241 (N_43241,N_40481,N_40370);
and U43242 (N_43242,N_41184,N_42040);
and U43243 (N_43243,N_41545,N_42101);
nor U43244 (N_43244,N_40807,N_41047);
and U43245 (N_43245,N_40548,N_40375);
and U43246 (N_43246,N_41597,N_40289);
or U43247 (N_43247,N_40886,N_42376);
and U43248 (N_43248,N_40713,N_40515);
nor U43249 (N_43249,N_40633,N_40281);
nand U43250 (N_43250,N_41841,N_40398);
and U43251 (N_43251,N_42385,N_41422);
and U43252 (N_43252,N_41798,N_41285);
or U43253 (N_43253,N_41042,N_41801);
nor U43254 (N_43254,N_41252,N_40775);
or U43255 (N_43255,N_41220,N_40801);
or U43256 (N_43256,N_41591,N_40128);
and U43257 (N_43257,N_41790,N_42095);
and U43258 (N_43258,N_41973,N_42201);
nand U43259 (N_43259,N_40211,N_41410);
nor U43260 (N_43260,N_41858,N_40059);
nand U43261 (N_43261,N_42337,N_41416);
and U43262 (N_43262,N_41243,N_42042);
and U43263 (N_43263,N_41150,N_41831);
or U43264 (N_43264,N_41972,N_42418);
nor U43265 (N_43265,N_40332,N_41845);
nor U43266 (N_43266,N_41794,N_42406);
xor U43267 (N_43267,N_42061,N_40482);
nand U43268 (N_43268,N_40843,N_41389);
nand U43269 (N_43269,N_40030,N_40669);
or U43270 (N_43270,N_40275,N_42217);
nor U43271 (N_43271,N_41999,N_40998);
and U43272 (N_43272,N_41778,N_41550);
nor U43273 (N_43273,N_40176,N_40991);
nand U43274 (N_43274,N_40373,N_40890);
and U43275 (N_43275,N_40828,N_40926);
xor U43276 (N_43276,N_41214,N_41140);
or U43277 (N_43277,N_40663,N_40112);
nand U43278 (N_43278,N_40026,N_40165);
or U43279 (N_43279,N_41627,N_41560);
or U43280 (N_43280,N_41902,N_41160);
nand U43281 (N_43281,N_40677,N_41649);
xor U43282 (N_43282,N_41464,N_41006);
nor U43283 (N_43283,N_42471,N_42268);
nand U43284 (N_43284,N_41154,N_41805);
xor U43285 (N_43285,N_40565,N_41658);
xnor U43286 (N_43286,N_40526,N_40915);
nor U43287 (N_43287,N_41974,N_41797);
xor U43288 (N_43288,N_40214,N_42120);
xor U43289 (N_43289,N_40269,N_41908);
nor U43290 (N_43290,N_41396,N_40429);
nor U43291 (N_43291,N_41236,N_42441);
or U43292 (N_43292,N_40283,N_42387);
nand U43293 (N_43293,N_41784,N_41672);
and U43294 (N_43294,N_42354,N_42497);
nor U43295 (N_43295,N_42051,N_40897);
nor U43296 (N_43296,N_40943,N_42329);
xnor U43297 (N_43297,N_40403,N_40216);
nand U43298 (N_43298,N_41477,N_40354);
and U43299 (N_43299,N_42041,N_41060);
or U43300 (N_43300,N_41189,N_41370);
and U43301 (N_43301,N_40179,N_41843);
or U43302 (N_43302,N_41971,N_42344);
nor U43303 (N_43303,N_40022,N_42074);
nand U43304 (N_43304,N_40286,N_40746);
or U43305 (N_43305,N_40172,N_40247);
xnor U43306 (N_43306,N_42059,N_41533);
and U43307 (N_43307,N_40695,N_40979);
xnor U43308 (N_43308,N_41442,N_42318);
nor U43309 (N_43309,N_40191,N_41660);
xnor U43310 (N_43310,N_41769,N_40258);
xor U43311 (N_43311,N_40408,N_42130);
nand U43312 (N_43312,N_42137,N_41904);
or U43313 (N_43313,N_40027,N_41586);
and U43314 (N_43314,N_41913,N_42333);
or U43315 (N_43315,N_41262,N_42077);
nor U43316 (N_43316,N_41509,N_42000);
or U43317 (N_43317,N_41115,N_42282);
xnor U43318 (N_43318,N_41304,N_41849);
nand U43319 (N_43319,N_42108,N_41746);
xnor U43320 (N_43320,N_40958,N_40279);
xnor U43321 (N_43321,N_40252,N_42151);
nand U43322 (N_43322,N_40428,N_40045);
and U43323 (N_43323,N_41528,N_40044);
nor U43324 (N_43324,N_42110,N_41302);
xnor U43325 (N_43325,N_42098,N_40021);
nand U43326 (N_43326,N_41046,N_42023);
nand U43327 (N_43327,N_40462,N_40062);
nand U43328 (N_43328,N_41481,N_41429);
nand U43329 (N_43329,N_41241,N_40043);
and U43330 (N_43330,N_41379,N_40195);
or U43331 (N_43331,N_40206,N_41898);
nor U43332 (N_43332,N_41448,N_42426);
nand U43333 (N_43333,N_42365,N_41975);
nand U43334 (N_43334,N_41984,N_40511);
or U43335 (N_43335,N_41466,N_40928);
and U43336 (N_43336,N_41197,N_40874);
and U43337 (N_43337,N_40394,N_42404);
and U43338 (N_43338,N_40145,N_41199);
nand U43339 (N_43339,N_41245,N_42132);
and U43340 (N_43340,N_40376,N_41009);
and U43341 (N_43341,N_40479,N_42241);
or U43342 (N_43342,N_40959,N_41326);
nor U43343 (N_43343,N_42142,N_42135);
and U43344 (N_43344,N_41541,N_41755);
xnor U43345 (N_43345,N_40949,N_40372);
nand U43346 (N_43346,N_41598,N_42057);
or U43347 (N_43347,N_40036,N_41038);
and U43348 (N_43348,N_40163,N_41761);
nand U43349 (N_43349,N_41878,N_40662);
or U43350 (N_43350,N_40284,N_40741);
xor U43351 (N_43351,N_41035,N_40425);
nand U43352 (N_43352,N_41240,N_42214);
nor U43353 (N_43353,N_42141,N_40917);
and U43354 (N_43354,N_41544,N_42248);
nand U43355 (N_43355,N_41450,N_40081);
xnor U43356 (N_43356,N_40541,N_42157);
xnor U43357 (N_43357,N_41662,N_41916);
and U43358 (N_43358,N_41516,N_40701);
nor U43359 (N_43359,N_40406,N_40387);
or U43360 (N_43360,N_40818,N_40613);
and U43361 (N_43361,N_41561,N_42222);
nand U43362 (N_43362,N_41813,N_40740);
nand U43363 (N_43363,N_41575,N_42480);
nand U43364 (N_43364,N_40575,N_40181);
nor U43365 (N_43365,N_40802,N_41321);
xor U43366 (N_43366,N_41782,N_41630);
or U43367 (N_43367,N_40447,N_42281);
nor U43368 (N_43368,N_41043,N_41191);
nand U43369 (N_43369,N_40095,N_41113);
or U43370 (N_43370,N_42425,N_41657);
xnor U43371 (N_43371,N_42048,N_40208);
and U43372 (N_43372,N_41759,N_40345);
xnor U43373 (N_43373,N_40138,N_42392);
xor U43374 (N_43374,N_42131,N_41876);
nand U43375 (N_43375,N_41393,N_41327);
nor U43376 (N_43376,N_40906,N_40638);
nand U43377 (N_43377,N_40201,N_41204);
nor U43378 (N_43378,N_42489,N_40993);
and U43379 (N_43379,N_40199,N_40820);
or U43380 (N_43380,N_41032,N_41474);
and U43381 (N_43381,N_42481,N_40047);
xnor U43382 (N_43382,N_40516,N_40735);
nand U43383 (N_43383,N_41760,N_41650);
xor U43384 (N_43384,N_41646,N_41135);
nor U43385 (N_43385,N_41631,N_41039);
or U43386 (N_43386,N_42269,N_41722);
nor U43387 (N_43387,N_40086,N_41534);
and U43388 (N_43388,N_40576,N_40704);
and U43389 (N_43389,N_41013,N_41030);
and U43390 (N_43390,N_40494,N_41155);
nor U43391 (N_43391,N_41488,N_41418);
or U43392 (N_43392,N_40136,N_40305);
nand U43393 (N_43393,N_40846,N_40439);
xor U43394 (N_43394,N_40760,N_41001);
and U43395 (N_43395,N_40841,N_42188);
nor U43396 (N_43396,N_40965,N_42382);
and U43397 (N_43397,N_40237,N_40937);
nand U43398 (N_43398,N_41213,N_41628);
and U43399 (N_43399,N_41955,N_40972);
nand U43400 (N_43400,N_40301,N_41624);
and U43401 (N_43401,N_40975,N_41208);
nand U43402 (N_43402,N_40097,N_40079);
xnor U43403 (N_43403,N_41505,N_41272);
and U43404 (N_43404,N_42290,N_41900);
nand U43405 (N_43405,N_40545,N_40090);
nor U43406 (N_43406,N_41536,N_40981);
xnor U43407 (N_43407,N_42475,N_41546);
nand U43408 (N_43408,N_40805,N_40869);
and U43409 (N_43409,N_42069,N_42496);
xor U43410 (N_43410,N_41100,N_41713);
nand U43411 (N_43411,N_41310,N_41130);
nor U43412 (N_43412,N_41004,N_40799);
xnor U43413 (N_43413,N_41671,N_41997);
and U43414 (N_43414,N_41786,N_40606);
and U43415 (N_43415,N_40324,N_42386);
and U43416 (N_43416,N_41315,N_41260);
and U43417 (N_43417,N_41485,N_42060);
and U43418 (N_43418,N_42367,N_41188);
xor U43419 (N_43419,N_41834,N_40436);
and U43420 (N_43420,N_41455,N_41857);
nand U43421 (N_43421,N_40288,N_41367);
xor U43422 (N_43422,N_41377,N_41044);
nor U43423 (N_43423,N_41374,N_41289);
nand U43424 (N_43424,N_40693,N_41384);
xor U43425 (N_43425,N_42177,N_41605);
nor U43426 (N_43426,N_42341,N_40867);
nor U43427 (N_43427,N_41202,N_40495);
or U43428 (N_43428,N_40457,N_40327);
nand U43429 (N_43429,N_40684,N_41891);
and U43430 (N_43430,N_41333,N_40168);
and U43431 (N_43431,N_42148,N_40913);
and U43432 (N_43432,N_41394,N_40362);
and U43433 (N_43433,N_41116,N_40761);
xnor U43434 (N_43434,N_41376,N_40392);
and U43435 (N_43435,N_42190,N_40643);
or U43436 (N_43436,N_40225,N_40001);
and U43437 (N_43437,N_40552,N_42021);
xor U43438 (N_43438,N_40033,N_41507);
nand U43439 (N_43439,N_40782,N_40262);
xor U43440 (N_43440,N_40838,N_41814);
or U43441 (N_43441,N_41020,N_41639);
nand U43442 (N_43442,N_41779,N_41270);
and U43443 (N_43443,N_40210,N_40524);
nor U43444 (N_43444,N_40472,N_42442);
or U43445 (N_43445,N_42456,N_42123);
or U43446 (N_43446,N_41415,N_41319);
nand U43447 (N_43447,N_40031,N_41400);
or U43448 (N_43448,N_42419,N_41308);
or U43449 (N_43449,N_41242,N_40361);
xnor U43450 (N_43450,N_42152,N_40609);
and U43451 (N_43451,N_41000,N_41856);
and U43452 (N_43452,N_41860,N_41749);
xor U43453 (N_43453,N_40140,N_40463);
or U43454 (N_43454,N_40411,N_42255);
or U43455 (N_43455,N_41081,N_40129);
and U43456 (N_43456,N_40811,N_41259);
nor U43457 (N_43457,N_42056,N_40611);
nor U43458 (N_43458,N_42118,N_40605);
or U43459 (N_43459,N_40273,N_42375);
xor U43460 (N_43460,N_41287,N_41524);
nand U43461 (N_43461,N_41185,N_40243);
nand U43462 (N_43462,N_41451,N_40970);
or U43463 (N_43463,N_41848,N_41037);
xor U43464 (N_43464,N_41522,N_41719);
xor U43465 (N_43465,N_41648,N_41935);
xor U43466 (N_43466,N_41368,N_40619);
and U43467 (N_43467,N_41144,N_41571);
xor U43468 (N_43468,N_40884,N_40189);
and U43469 (N_43469,N_41159,N_41055);
nor U43470 (N_43470,N_41877,N_41223);
xor U43471 (N_43471,N_41019,N_41476);
nand U43472 (N_43472,N_41171,N_41995);
xor U43473 (N_43473,N_40317,N_41766);
xor U43474 (N_43474,N_40598,N_40850);
nand U43475 (N_43475,N_40215,N_40341);
or U43476 (N_43476,N_42381,N_41484);
or U43477 (N_43477,N_40688,N_42401);
xor U43478 (N_43478,N_40366,N_40547);
and U43479 (N_43479,N_41819,N_41612);
or U43480 (N_43480,N_40971,N_41537);
nor U43481 (N_43481,N_41084,N_41583);
nor U43482 (N_43482,N_41103,N_40323);
nor U43483 (N_43483,N_40017,N_42296);
nor U43484 (N_43484,N_42285,N_40762);
nand U43485 (N_43485,N_41490,N_41087);
and U43486 (N_43486,N_40600,N_42273);
or U43487 (N_43487,N_41608,N_41453);
and U43488 (N_43488,N_42062,N_41763);
xor U43489 (N_43489,N_41864,N_41064);
and U43490 (N_43490,N_41993,N_42154);
and U43491 (N_43491,N_40207,N_41356);
or U43492 (N_43492,N_42240,N_40990);
or U43493 (N_43493,N_41479,N_40448);
nor U43494 (N_43494,N_40316,N_41232);
and U43495 (N_43495,N_42155,N_42345);
nor U43496 (N_43496,N_40272,N_41235);
nor U43497 (N_43497,N_41823,N_40444);
nand U43498 (N_43498,N_41644,N_41362);
xor U43499 (N_43499,N_40597,N_40430);
nor U43500 (N_43500,N_42389,N_41022);
and U43501 (N_43501,N_41198,N_41391);
nand U43502 (N_43502,N_40844,N_42085);
xnor U43503 (N_43503,N_41078,N_41636);
or U43504 (N_43504,N_41847,N_40631);
xor U43505 (N_43505,N_41799,N_41675);
or U43506 (N_43506,N_40454,N_41061);
xor U43507 (N_43507,N_42055,N_40485);
nand U43508 (N_43508,N_40503,N_42025);
or U43509 (N_43509,N_42467,N_42206);
xor U43510 (N_43510,N_42431,N_42075);
nand U43511 (N_43511,N_41162,N_41028);
xnor U43512 (N_43512,N_40934,N_40830);
xor U43513 (N_43513,N_40957,N_41641);
xnor U43514 (N_43514,N_40532,N_41712);
xor U43515 (N_43515,N_41175,N_42260);
or U43516 (N_43516,N_40089,N_40078);
nand U43517 (N_43517,N_41706,N_41027);
and U43518 (N_43518,N_41596,N_42460);
and U43519 (N_43519,N_42239,N_40618);
xor U43520 (N_43520,N_40711,N_41910);
and U43521 (N_43521,N_40255,N_41928);
xor U43522 (N_43522,N_40196,N_41780);
nand U43523 (N_43523,N_41005,N_40963);
or U43524 (N_43524,N_42383,N_41210);
nor U43525 (N_43525,N_42428,N_42043);
nor U43526 (N_43526,N_42165,N_41751);
or U43527 (N_43527,N_41634,N_42342);
nand U43528 (N_43528,N_40736,N_40710);
xnor U43529 (N_43529,N_40034,N_41901);
and U43530 (N_43530,N_41704,N_42080);
nand U43531 (N_43531,N_40783,N_41491);
nand U43532 (N_43532,N_42422,N_42408);
nand U43533 (N_43533,N_40903,N_41689);
xor U43534 (N_43534,N_41181,N_40719);
nor U43535 (N_43535,N_41316,N_42271);
or U43536 (N_43536,N_41699,N_40733);
xor U43537 (N_43537,N_40057,N_42058);
nor U43538 (N_43538,N_41737,N_41667);
nor U43539 (N_43539,N_41721,N_40953);
nor U43540 (N_43540,N_41372,N_41734);
nand U43541 (N_43541,N_40410,N_41216);
or U43542 (N_43542,N_41783,N_41940);
nand U43543 (N_43543,N_40758,N_40486);
nor U43544 (N_43544,N_40478,N_42303);
nand U43545 (N_43545,N_41603,N_41548);
xnor U43546 (N_43546,N_41640,N_42046);
xor U43547 (N_43547,N_40115,N_40469);
xor U43548 (N_43548,N_42172,N_40769);
xor U43549 (N_43549,N_41074,N_41837);
or U43550 (N_43550,N_42277,N_42224);
nand U43551 (N_43551,N_41126,N_42092);
or U43552 (N_43552,N_40114,N_42140);
nand U43553 (N_43553,N_40810,N_40473);
xnor U43554 (N_43554,N_40497,N_41428);
nor U43555 (N_43555,N_40964,N_40656);
xor U43556 (N_43556,N_40847,N_41359);
nor U43557 (N_43557,N_41696,N_42102);
nand U43558 (N_43558,N_42212,N_40453);
or U43559 (N_43559,N_40455,N_41141);
nand U43560 (N_43560,N_40171,N_41211);
nand U43561 (N_43561,N_41482,N_40773);
xnor U43562 (N_43562,N_40559,N_41399);
and U43563 (N_43563,N_41731,N_41691);
or U43564 (N_43564,N_41897,N_41195);
nor U43565 (N_43565,N_40094,N_40793);
or U43566 (N_43566,N_40634,N_40727);
nor U43567 (N_43567,N_41803,N_40510);
or U43568 (N_43568,N_40891,N_42257);
xor U43569 (N_43569,N_41249,N_40065);
nor U43570 (N_43570,N_41752,N_40437);
xor U43571 (N_43571,N_41125,N_41052);
and U43572 (N_43572,N_40896,N_40162);
and U43573 (N_43573,N_40625,N_40144);
or U43574 (N_43574,N_40558,N_41180);
xnor U43575 (N_43575,N_42114,N_42364);
or U43576 (N_43576,N_41551,N_41692);
or U43577 (N_43577,N_40786,N_40287);
and U43578 (N_43578,N_41970,N_41457);
and U43579 (N_43579,N_41511,N_40553);
xor U43580 (N_43580,N_41263,N_41068);
nor U43581 (N_43581,N_40061,N_40236);
or U43582 (N_43582,N_40882,N_40966);
xnor U43583 (N_43583,N_41733,N_40290);
nand U43584 (N_43584,N_42197,N_41567);
and U43585 (N_43585,N_42223,N_42338);
and U43586 (N_43586,N_42454,N_41493);
xor U43587 (N_43587,N_41435,N_41015);
nand U43588 (N_43588,N_40187,N_41716);
or U43589 (N_43589,N_40058,N_40932);
nand U43590 (N_43590,N_42066,N_42249);
or U43591 (N_43591,N_41237,N_40627);
xor U43592 (N_43592,N_41988,N_40645);
or U43593 (N_43593,N_40834,N_40534);
or U43594 (N_43594,N_42355,N_41569);
and U43595 (N_43595,N_42070,N_40491);
nor U43596 (N_43596,N_40591,N_41977);
nand U43597 (N_43597,N_40647,N_42246);
nand U43598 (N_43598,N_40742,N_42317);
nand U43599 (N_43599,N_41909,N_41386);
xor U43600 (N_43600,N_41489,N_40509);
nand U43601 (N_43601,N_42031,N_40956);
nor U43602 (N_43602,N_41683,N_41102);
nor U43603 (N_43603,N_42170,N_40518);
nand U43604 (N_43604,N_40893,N_42484);
or U43605 (N_43605,N_40070,N_40912);
nor U43606 (N_43606,N_41023,N_42359);
or U43607 (N_43607,N_40174,N_42156);
nor U43608 (N_43608,N_40120,N_40512);
nor U43609 (N_43609,N_40015,N_40670);
or U43610 (N_43610,N_40490,N_40143);
nand U43611 (N_43611,N_40182,N_41354);
nand U43612 (N_43612,N_41122,N_42024);
nand U43613 (N_43613,N_40876,N_40770);
nand U43614 (N_43614,N_40697,N_41375);
nor U43615 (N_43615,N_42437,N_41686);
nor U43616 (N_43616,N_41388,N_41577);
nor U43617 (N_43617,N_41547,N_41965);
nor U43618 (N_43618,N_42178,N_40227);
or U43619 (N_43619,N_40464,N_40241);
nor U43620 (N_43620,N_42328,N_41859);
or U43621 (N_43621,N_42162,N_41312);
nand U43622 (N_43622,N_41697,N_40668);
nor U43623 (N_43623,N_41129,N_41008);
and U43624 (N_43624,N_40337,N_40391);
and U43625 (N_43625,N_40242,N_42089);
and U43626 (N_43626,N_40555,N_41563);
or U43627 (N_43627,N_40405,N_40658);
xor U43628 (N_43628,N_41390,N_40356);
nor U43629 (N_43629,N_40069,N_41364);
nand U43630 (N_43630,N_41840,N_41112);
and U43631 (N_43631,N_42453,N_41655);
xnor U43632 (N_43632,N_41471,N_42220);
and U43633 (N_43633,N_42187,N_40484);
nand U43634 (N_43634,N_40749,N_40099);
and U43635 (N_43635,N_41067,N_41661);
nor U43636 (N_43636,N_41787,N_40564);
nor U43637 (N_43637,N_42449,N_40857);
and U43638 (N_43638,N_40845,N_40901);
xor U43639 (N_43639,N_41071,N_42423);
nand U43640 (N_43640,N_41440,N_42413);
and U43641 (N_43641,N_40759,N_40522);
xnor U43642 (N_43642,N_41504,N_42012);
nor U43643 (N_43643,N_41907,N_41945);
and U43644 (N_43644,N_41492,N_41163);
or U43645 (N_43645,N_40690,N_40321);
nand U43646 (N_43646,N_41554,N_41684);
xnor U43647 (N_43647,N_41950,N_41888);
and U43648 (N_43648,N_40291,N_42319);
or U43649 (N_43649,N_41424,N_40151);
xor U43650 (N_43650,N_40804,N_41366);
nand U43651 (N_43651,N_41288,N_40644);
or U43652 (N_43652,N_41218,N_42494);
nand U43653 (N_43653,N_41134,N_40380);
and U43654 (N_43654,N_41345,N_41462);
nor U43655 (N_43655,N_41526,N_42274);
and U43656 (N_43656,N_40010,N_42250);
nand U43657 (N_43657,N_41576,N_42420);
nor U43658 (N_43658,N_41867,N_40111);
and U43659 (N_43659,N_41343,N_40046);
nand U43660 (N_43660,N_40800,N_41294);
or U43661 (N_43661,N_41403,N_41730);
nor U43662 (N_43662,N_40751,N_40185);
or U43663 (N_43663,N_41138,N_41306);
nor U43664 (N_43664,N_41923,N_41905);
nor U43665 (N_43665,N_42373,N_40339);
nor U43666 (N_43666,N_40808,N_42008);
nand U43667 (N_43667,N_42231,N_41169);
nand U43668 (N_43668,N_41221,N_41349);
nand U43669 (N_43669,N_41053,N_40277);
nand U43670 (N_43670,N_41072,N_41938);
or U43671 (N_43671,N_41031,N_41329);
and U43672 (N_43672,N_40396,N_40170);
nand U43673 (N_43673,N_41949,N_40175);
and U43674 (N_43674,N_40578,N_41487);
or U43675 (N_43675,N_41478,N_40088);
xnor U43676 (N_43676,N_41809,N_41338);
nand U43677 (N_43677,N_42078,N_40969);
or U43678 (N_43678,N_41562,N_40747);
nand U43679 (N_43679,N_41732,N_40652);
xor U43680 (N_43680,N_42283,N_42483);
xnor U43681 (N_43681,N_41397,N_40292);
nor U43682 (N_43682,N_40815,N_40646);
and U43683 (N_43683,N_41414,N_40308);
nor U43684 (N_43684,N_40353,N_40885);
nand U43685 (N_43685,N_40382,N_40918);
nor U43686 (N_43686,N_42111,N_40251);
nor U43687 (N_43687,N_40051,N_40049);
nor U43688 (N_43688,N_41227,N_42316);
nand U43689 (N_43689,N_41647,N_41925);
and U43690 (N_43690,N_40977,N_40443);
xnor U43691 (N_43691,N_40389,N_41961);
nor U43692 (N_43692,N_41145,N_40593);
or U43693 (N_43693,N_42351,N_41069);
nor U43694 (N_43694,N_42133,N_40873);
and U43695 (N_43695,N_41844,N_41604);
or U43696 (N_43696,N_41439,N_41058);
xnor U43697 (N_43697,N_40213,N_40282);
nand U43698 (N_43698,N_40431,N_42233);
nand U43699 (N_43699,N_40745,N_40100);
nor U43700 (N_43700,N_40119,N_40967);
xnor U43701 (N_43701,N_41764,N_40831);
or U43702 (N_43702,N_41839,N_40158);
xnor U43703 (N_43703,N_40098,N_42458);
nor U43704 (N_43704,N_41621,N_41469);
nand U43705 (N_43705,N_41868,N_40257);
nand U43706 (N_43706,N_42192,N_40420);
nor U43707 (N_43707,N_41225,N_41351);
nor U43708 (N_43708,N_40579,N_42334);
nor U43709 (N_43709,N_42476,N_40790);
xnor U43710 (N_43710,N_40851,N_40950);
nand U43711 (N_43711,N_41434,N_41080);
xnor U43712 (N_43712,N_40940,N_41767);
nor U43713 (N_43713,N_40864,N_41668);
nor U43714 (N_43714,N_40072,N_42278);
nor U43715 (N_43715,N_41480,N_40836);
nor U43716 (N_43716,N_40365,N_42438);
xor U43717 (N_43717,N_40539,N_41829);
nor U43718 (N_43718,N_41818,N_40925);
xnor U43719 (N_43719,N_40995,N_42124);
or U43720 (N_43720,N_42498,N_41652);
and U43721 (N_43721,N_40377,N_40107);
xnor U43722 (N_43722,N_40952,N_40848);
and U43723 (N_43723,N_40968,N_40767);
xnor U43724 (N_43724,N_41350,N_42309);
nor U43725 (N_43725,N_41807,N_40418);
or U43726 (N_43726,N_40778,N_41331);
or U43727 (N_43727,N_41239,N_40466);
and U43728 (N_43728,N_42109,N_41114);
nor U43729 (N_43729,N_41826,N_41914);
nand U43730 (N_43730,N_40561,N_40689);
xor U43731 (N_43731,N_40412,N_42306);
nand U43732 (N_43732,N_41313,N_41470);
nor U43733 (N_43733,N_42263,N_41992);
xnor U43734 (N_43734,N_41854,N_40153);
or U43735 (N_43735,N_40164,N_42400);
nor U43736 (N_43736,N_40866,N_40202);
nor U43737 (N_43737,N_40717,N_40692);
xnor U43738 (N_43738,N_41870,N_42251);
and U43739 (N_43739,N_40294,N_40303);
xor U43740 (N_43740,N_40137,N_40427);
and U43741 (N_43741,N_41698,N_41601);
and U43742 (N_43742,N_42134,N_41334);
nor U43743 (N_43743,N_40577,N_40529);
nand U43744 (N_43744,N_42326,N_41613);
nand U43745 (N_43745,N_41361,N_40121);
or U43746 (N_43746,N_41743,N_40259);
or U43747 (N_43747,N_40823,N_40254);
and U43748 (N_43748,N_40190,N_40659);
nand U43749 (N_43749,N_40868,N_41010);
nor U43750 (N_43750,N_41262,N_40201);
nor U43751 (N_43751,N_40093,N_41215);
xnor U43752 (N_43752,N_40741,N_42222);
nand U43753 (N_43753,N_40888,N_42099);
xor U43754 (N_43754,N_40202,N_42295);
and U43755 (N_43755,N_41269,N_41289);
xor U43756 (N_43756,N_41901,N_40239);
nand U43757 (N_43757,N_42160,N_42193);
nor U43758 (N_43758,N_40446,N_40544);
nor U43759 (N_43759,N_40197,N_41688);
xor U43760 (N_43760,N_40476,N_42073);
nor U43761 (N_43761,N_40687,N_41701);
xnor U43762 (N_43762,N_42331,N_41433);
and U43763 (N_43763,N_41062,N_41206);
and U43764 (N_43764,N_41684,N_40784);
nand U43765 (N_43765,N_41890,N_41512);
xnor U43766 (N_43766,N_41256,N_41701);
nand U43767 (N_43767,N_41454,N_40756);
nor U43768 (N_43768,N_40367,N_40248);
and U43769 (N_43769,N_40939,N_41520);
nand U43770 (N_43770,N_42189,N_41401);
nor U43771 (N_43771,N_40741,N_41780);
xnor U43772 (N_43772,N_41343,N_41112);
xnor U43773 (N_43773,N_40144,N_42495);
or U43774 (N_43774,N_41980,N_40140);
xor U43775 (N_43775,N_40612,N_41311);
xnor U43776 (N_43776,N_41127,N_40865);
or U43777 (N_43777,N_41425,N_40341);
nor U43778 (N_43778,N_41324,N_41835);
or U43779 (N_43779,N_42220,N_42387);
or U43780 (N_43780,N_40589,N_40257);
nor U43781 (N_43781,N_40088,N_41420);
or U43782 (N_43782,N_40072,N_41996);
or U43783 (N_43783,N_42468,N_42078);
and U43784 (N_43784,N_40953,N_41799);
or U43785 (N_43785,N_41544,N_42224);
nand U43786 (N_43786,N_41943,N_41967);
nand U43787 (N_43787,N_40751,N_41910);
nor U43788 (N_43788,N_40627,N_41333);
or U43789 (N_43789,N_40865,N_42239);
or U43790 (N_43790,N_41352,N_41001);
nor U43791 (N_43791,N_40309,N_40811);
and U43792 (N_43792,N_42317,N_41353);
and U43793 (N_43793,N_41498,N_41695);
nor U43794 (N_43794,N_42316,N_42208);
nor U43795 (N_43795,N_41368,N_42107);
nor U43796 (N_43796,N_41994,N_40399);
or U43797 (N_43797,N_40520,N_40960);
or U43798 (N_43798,N_40908,N_41706);
and U43799 (N_43799,N_41281,N_40624);
xor U43800 (N_43800,N_42495,N_40635);
and U43801 (N_43801,N_40385,N_42103);
or U43802 (N_43802,N_40361,N_42388);
xnor U43803 (N_43803,N_41957,N_42375);
nand U43804 (N_43804,N_40340,N_41455);
xnor U43805 (N_43805,N_40234,N_41467);
or U43806 (N_43806,N_40815,N_40903);
and U43807 (N_43807,N_41941,N_42347);
nand U43808 (N_43808,N_42238,N_40739);
and U43809 (N_43809,N_41118,N_40262);
and U43810 (N_43810,N_40262,N_40709);
nand U43811 (N_43811,N_42051,N_40408);
and U43812 (N_43812,N_40570,N_41719);
and U43813 (N_43813,N_41213,N_41632);
xor U43814 (N_43814,N_41324,N_42329);
xnor U43815 (N_43815,N_40152,N_41638);
nand U43816 (N_43816,N_40273,N_42058);
and U43817 (N_43817,N_41871,N_40637);
nand U43818 (N_43818,N_41131,N_40502);
or U43819 (N_43819,N_42022,N_42425);
or U43820 (N_43820,N_40198,N_40070);
nor U43821 (N_43821,N_40468,N_40166);
or U43822 (N_43822,N_41338,N_41396);
and U43823 (N_43823,N_41437,N_40428);
nand U43824 (N_43824,N_40186,N_40906);
and U43825 (N_43825,N_40646,N_42425);
or U43826 (N_43826,N_42294,N_40177);
nor U43827 (N_43827,N_40241,N_40056);
and U43828 (N_43828,N_41709,N_41505);
and U43829 (N_43829,N_40768,N_40226);
nand U43830 (N_43830,N_41375,N_41542);
xnor U43831 (N_43831,N_41807,N_40423);
and U43832 (N_43832,N_41213,N_41167);
or U43833 (N_43833,N_41490,N_40045);
or U43834 (N_43834,N_41954,N_41544);
nand U43835 (N_43835,N_41568,N_40516);
xor U43836 (N_43836,N_41604,N_40085);
xnor U43837 (N_43837,N_41125,N_40591);
nor U43838 (N_43838,N_40079,N_42379);
nor U43839 (N_43839,N_40998,N_41020);
or U43840 (N_43840,N_42157,N_40942);
or U43841 (N_43841,N_42400,N_40964);
nand U43842 (N_43842,N_40195,N_41388);
nand U43843 (N_43843,N_40332,N_40676);
and U43844 (N_43844,N_41169,N_41223);
nor U43845 (N_43845,N_41625,N_41117);
or U43846 (N_43846,N_40251,N_41872);
xor U43847 (N_43847,N_42243,N_40908);
xnor U43848 (N_43848,N_40163,N_41684);
nor U43849 (N_43849,N_40095,N_41149);
xor U43850 (N_43850,N_40328,N_40728);
or U43851 (N_43851,N_42475,N_41422);
and U43852 (N_43852,N_40407,N_41512);
or U43853 (N_43853,N_42213,N_40429);
nand U43854 (N_43854,N_40154,N_40107);
nand U43855 (N_43855,N_40073,N_41967);
or U43856 (N_43856,N_40312,N_40452);
and U43857 (N_43857,N_40461,N_40883);
nand U43858 (N_43858,N_40321,N_41547);
nor U43859 (N_43859,N_40485,N_41167);
nor U43860 (N_43860,N_40262,N_42139);
nor U43861 (N_43861,N_41330,N_40949);
nor U43862 (N_43862,N_42030,N_41367);
or U43863 (N_43863,N_41871,N_41039);
xor U43864 (N_43864,N_41058,N_41837);
xnor U43865 (N_43865,N_40905,N_40307);
xor U43866 (N_43866,N_42041,N_41159);
xnor U43867 (N_43867,N_42253,N_42095);
nand U43868 (N_43868,N_42317,N_41097);
and U43869 (N_43869,N_41862,N_40486);
or U43870 (N_43870,N_40994,N_40753);
and U43871 (N_43871,N_40621,N_40884);
and U43872 (N_43872,N_40485,N_41572);
or U43873 (N_43873,N_40121,N_40085);
xnor U43874 (N_43874,N_40619,N_42384);
and U43875 (N_43875,N_40689,N_40679);
and U43876 (N_43876,N_41586,N_41004);
or U43877 (N_43877,N_40678,N_40064);
xnor U43878 (N_43878,N_40708,N_41931);
xor U43879 (N_43879,N_42460,N_41657);
or U43880 (N_43880,N_40074,N_40075);
or U43881 (N_43881,N_40775,N_40636);
nand U43882 (N_43882,N_40879,N_40870);
and U43883 (N_43883,N_42485,N_41889);
xnor U43884 (N_43884,N_40362,N_41233);
nor U43885 (N_43885,N_40643,N_41542);
nor U43886 (N_43886,N_42032,N_41077);
and U43887 (N_43887,N_41195,N_41109);
and U43888 (N_43888,N_40091,N_40185);
nand U43889 (N_43889,N_42037,N_40999);
nand U43890 (N_43890,N_40897,N_40715);
xor U43891 (N_43891,N_40508,N_41032);
nor U43892 (N_43892,N_41254,N_41665);
nor U43893 (N_43893,N_40249,N_42318);
nand U43894 (N_43894,N_40402,N_42142);
or U43895 (N_43895,N_41406,N_41292);
nor U43896 (N_43896,N_41507,N_42020);
xor U43897 (N_43897,N_41161,N_41382);
nor U43898 (N_43898,N_40966,N_40220);
nand U43899 (N_43899,N_40691,N_40891);
nand U43900 (N_43900,N_41278,N_40806);
xnor U43901 (N_43901,N_41187,N_41389);
nor U43902 (N_43902,N_42469,N_41308);
nand U43903 (N_43903,N_40490,N_42289);
xor U43904 (N_43904,N_40009,N_42254);
or U43905 (N_43905,N_40477,N_41113);
xnor U43906 (N_43906,N_40780,N_42284);
nand U43907 (N_43907,N_42414,N_40058);
nor U43908 (N_43908,N_41653,N_40597);
xnor U43909 (N_43909,N_40094,N_40171);
or U43910 (N_43910,N_42206,N_40430);
nor U43911 (N_43911,N_40081,N_40710);
nand U43912 (N_43912,N_41799,N_41126);
nand U43913 (N_43913,N_42310,N_40018);
nor U43914 (N_43914,N_41795,N_41275);
nor U43915 (N_43915,N_40757,N_42241);
nor U43916 (N_43916,N_42247,N_40774);
xnor U43917 (N_43917,N_41959,N_42332);
nor U43918 (N_43918,N_40245,N_40406);
nor U43919 (N_43919,N_40046,N_42381);
nor U43920 (N_43920,N_41011,N_40435);
or U43921 (N_43921,N_41378,N_40460);
and U43922 (N_43922,N_40060,N_40580);
and U43923 (N_43923,N_41150,N_40071);
xor U43924 (N_43924,N_40240,N_42416);
xor U43925 (N_43925,N_41483,N_41120);
and U43926 (N_43926,N_40163,N_40855);
nand U43927 (N_43927,N_42133,N_42143);
or U43928 (N_43928,N_41846,N_40097);
nor U43929 (N_43929,N_41265,N_40689);
or U43930 (N_43930,N_41689,N_41698);
nand U43931 (N_43931,N_42009,N_41843);
xnor U43932 (N_43932,N_41486,N_40835);
nand U43933 (N_43933,N_40768,N_41068);
xnor U43934 (N_43934,N_41620,N_40397);
nand U43935 (N_43935,N_42359,N_41911);
xnor U43936 (N_43936,N_41991,N_40505);
and U43937 (N_43937,N_41279,N_41769);
and U43938 (N_43938,N_41673,N_41405);
nand U43939 (N_43939,N_41589,N_42326);
nor U43940 (N_43940,N_40744,N_40479);
xor U43941 (N_43941,N_41776,N_42007);
nand U43942 (N_43942,N_42147,N_42018);
nor U43943 (N_43943,N_41651,N_41957);
xor U43944 (N_43944,N_41684,N_41577);
nand U43945 (N_43945,N_40751,N_40461);
xor U43946 (N_43946,N_41191,N_40894);
nand U43947 (N_43947,N_42286,N_42260);
nand U43948 (N_43948,N_41038,N_41348);
or U43949 (N_43949,N_41086,N_40955);
and U43950 (N_43950,N_40410,N_40529);
nor U43951 (N_43951,N_40298,N_42363);
nor U43952 (N_43952,N_40031,N_42225);
nor U43953 (N_43953,N_41217,N_42340);
xor U43954 (N_43954,N_40764,N_40781);
or U43955 (N_43955,N_40585,N_41027);
nor U43956 (N_43956,N_40657,N_40709);
nand U43957 (N_43957,N_41353,N_41139);
or U43958 (N_43958,N_42260,N_40512);
xnor U43959 (N_43959,N_41559,N_40031);
nor U43960 (N_43960,N_40728,N_40619);
xor U43961 (N_43961,N_42081,N_41361);
nor U43962 (N_43962,N_40083,N_41064);
xor U43963 (N_43963,N_41459,N_40958);
or U43964 (N_43964,N_40297,N_41937);
nand U43965 (N_43965,N_40461,N_41162);
or U43966 (N_43966,N_41028,N_42003);
and U43967 (N_43967,N_42004,N_40258);
xnor U43968 (N_43968,N_41995,N_40195);
or U43969 (N_43969,N_41061,N_40678);
nor U43970 (N_43970,N_40439,N_42426);
nor U43971 (N_43971,N_41680,N_41774);
and U43972 (N_43972,N_41141,N_41064);
nand U43973 (N_43973,N_40491,N_41269);
or U43974 (N_43974,N_40955,N_40185);
or U43975 (N_43975,N_42009,N_40399);
nand U43976 (N_43976,N_40139,N_41371);
nor U43977 (N_43977,N_41235,N_41194);
xor U43978 (N_43978,N_41912,N_42315);
xor U43979 (N_43979,N_40803,N_41377);
and U43980 (N_43980,N_42086,N_40877);
xnor U43981 (N_43981,N_42219,N_42064);
and U43982 (N_43982,N_41087,N_41963);
nor U43983 (N_43983,N_41520,N_41539);
and U43984 (N_43984,N_41995,N_41258);
and U43985 (N_43985,N_41679,N_42255);
or U43986 (N_43986,N_40865,N_40258);
xor U43987 (N_43987,N_41919,N_42379);
or U43988 (N_43988,N_41827,N_42118);
nand U43989 (N_43989,N_40737,N_41836);
or U43990 (N_43990,N_41265,N_42128);
or U43991 (N_43991,N_40928,N_41844);
xnor U43992 (N_43992,N_40323,N_41180);
or U43993 (N_43993,N_40875,N_41370);
xor U43994 (N_43994,N_42002,N_40156);
and U43995 (N_43995,N_41206,N_40807);
xnor U43996 (N_43996,N_42326,N_40732);
and U43997 (N_43997,N_42204,N_40199);
nor U43998 (N_43998,N_40837,N_40482);
nor U43999 (N_43999,N_40021,N_42437);
nand U44000 (N_44000,N_40827,N_42139);
or U44001 (N_44001,N_42126,N_41496);
nand U44002 (N_44002,N_42487,N_41673);
and U44003 (N_44003,N_40789,N_41422);
nor U44004 (N_44004,N_40597,N_40501);
or U44005 (N_44005,N_42381,N_41741);
or U44006 (N_44006,N_41247,N_40472);
nor U44007 (N_44007,N_40902,N_40347);
or U44008 (N_44008,N_42142,N_41188);
xnor U44009 (N_44009,N_41977,N_40735);
nor U44010 (N_44010,N_42271,N_40336);
nand U44011 (N_44011,N_40511,N_41408);
xor U44012 (N_44012,N_41385,N_41262);
nand U44013 (N_44013,N_40557,N_41208);
and U44014 (N_44014,N_41231,N_41055);
or U44015 (N_44015,N_42259,N_42280);
and U44016 (N_44016,N_41280,N_40245);
nor U44017 (N_44017,N_41560,N_42040);
xor U44018 (N_44018,N_42201,N_40342);
and U44019 (N_44019,N_40611,N_41624);
nand U44020 (N_44020,N_40148,N_41092);
nor U44021 (N_44021,N_42018,N_41164);
nor U44022 (N_44022,N_41482,N_40352);
or U44023 (N_44023,N_42106,N_41275);
nor U44024 (N_44024,N_42310,N_40784);
or U44025 (N_44025,N_41110,N_42223);
or U44026 (N_44026,N_41203,N_40856);
nor U44027 (N_44027,N_40983,N_41892);
nand U44028 (N_44028,N_41429,N_42250);
and U44029 (N_44029,N_41832,N_40576);
nand U44030 (N_44030,N_41064,N_41532);
nor U44031 (N_44031,N_40269,N_40108);
nor U44032 (N_44032,N_41998,N_40223);
nand U44033 (N_44033,N_42022,N_40543);
and U44034 (N_44034,N_40002,N_41447);
or U44035 (N_44035,N_40324,N_41061);
or U44036 (N_44036,N_40741,N_41186);
and U44037 (N_44037,N_42256,N_42046);
xor U44038 (N_44038,N_41507,N_41134);
nand U44039 (N_44039,N_41104,N_40428);
or U44040 (N_44040,N_42481,N_42223);
nand U44041 (N_44041,N_40562,N_42436);
nand U44042 (N_44042,N_41069,N_41685);
and U44043 (N_44043,N_40124,N_41989);
nor U44044 (N_44044,N_40647,N_41119);
nand U44045 (N_44045,N_40707,N_40523);
nand U44046 (N_44046,N_40054,N_41389);
nand U44047 (N_44047,N_40691,N_41390);
xor U44048 (N_44048,N_41469,N_42119);
nand U44049 (N_44049,N_40724,N_40081);
nand U44050 (N_44050,N_40114,N_41663);
nand U44051 (N_44051,N_40362,N_41336);
or U44052 (N_44052,N_41691,N_41572);
nand U44053 (N_44053,N_40058,N_41882);
and U44054 (N_44054,N_41456,N_40531);
nand U44055 (N_44055,N_40457,N_41752);
and U44056 (N_44056,N_40936,N_40515);
nand U44057 (N_44057,N_41821,N_42175);
and U44058 (N_44058,N_41193,N_41523);
and U44059 (N_44059,N_41297,N_41916);
or U44060 (N_44060,N_40338,N_42475);
and U44061 (N_44061,N_40715,N_40431);
or U44062 (N_44062,N_41767,N_40244);
or U44063 (N_44063,N_40197,N_41573);
or U44064 (N_44064,N_42179,N_41501);
nor U44065 (N_44065,N_42089,N_40910);
or U44066 (N_44066,N_41088,N_42007);
or U44067 (N_44067,N_41346,N_42343);
and U44068 (N_44068,N_42145,N_41010);
and U44069 (N_44069,N_42114,N_41965);
or U44070 (N_44070,N_41184,N_41153);
nand U44071 (N_44071,N_41467,N_42353);
nand U44072 (N_44072,N_42002,N_41159);
nor U44073 (N_44073,N_40195,N_40530);
and U44074 (N_44074,N_40344,N_40728);
xnor U44075 (N_44075,N_40132,N_41440);
and U44076 (N_44076,N_41441,N_40394);
xnor U44077 (N_44077,N_41745,N_40271);
xnor U44078 (N_44078,N_41164,N_40738);
xor U44079 (N_44079,N_42475,N_41405);
and U44080 (N_44080,N_40552,N_40134);
or U44081 (N_44081,N_42105,N_41170);
nor U44082 (N_44082,N_42206,N_41624);
or U44083 (N_44083,N_40505,N_40873);
or U44084 (N_44084,N_42445,N_40640);
nand U44085 (N_44085,N_42230,N_41643);
and U44086 (N_44086,N_40428,N_42124);
or U44087 (N_44087,N_42376,N_40476);
nor U44088 (N_44088,N_40601,N_41832);
xor U44089 (N_44089,N_41297,N_40394);
or U44090 (N_44090,N_42172,N_41904);
xnor U44091 (N_44091,N_40844,N_41281);
nand U44092 (N_44092,N_40307,N_42257);
xnor U44093 (N_44093,N_40124,N_41544);
nor U44094 (N_44094,N_41283,N_42003);
nor U44095 (N_44095,N_41206,N_40036);
or U44096 (N_44096,N_41267,N_40877);
xor U44097 (N_44097,N_41215,N_41495);
nor U44098 (N_44098,N_40738,N_41884);
or U44099 (N_44099,N_40734,N_40040);
xnor U44100 (N_44100,N_42467,N_40312);
or U44101 (N_44101,N_41865,N_41863);
and U44102 (N_44102,N_40115,N_41454);
xnor U44103 (N_44103,N_42052,N_40937);
nor U44104 (N_44104,N_41843,N_40715);
nor U44105 (N_44105,N_41951,N_42348);
nor U44106 (N_44106,N_41515,N_40195);
nand U44107 (N_44107,N_41332,N_41982);
xor U44108 (N_44108,N_41139,N_40582);
nand U44109 (N_44109,N_41129,N_42395);
and U44110 (N_44110,N_42017,N_40419);
nor U44111 (N_44111,N_42191,N_42230);
xor U44112 (N_44112,N_40625,N_42245);
xnor U44113 (N_44113,N_40891,N_41759);
xnor U44114 (N_44114,N_41087,N_40124);
nand U44115 (N_44115,N_40383,N_41554);
nor U44116 (N_44116,N_40905,N_41679);
nor U44117 (N_44117,N_41740,N_40272);
xnor U44118 (N_44118,N_41257,N_41538);
or U44119 (N_44119,N_41596,N_40968);
nor U44120 (N_44120,N_42346,N_42270);
and U44121 (N_44121,N_40704,N_40327);
xor U44122 (N_44122,N_42133,N_41232);
and U44123 (N_44123,N_41880,N_41080);
and U44124 (N_44124,N_40738,N_40353);
nand U44125 (N_44125,N_41961,N_40486);
xor U44126 (N_44126,N_42156,N_42370);
xor U44127 (N_44127,N_40498,N_42277);
xnor U44128 (N_44128,N_40901,N_41348);
nor U44129 (N_44129,N_40992,N_41633);
and U44130 (N_44130,N_42095,N_41538);
xor U44131 (N_44131,N_42451,N_40516);
or U44132 (N_44132,N_41052,N_41609);
nand U44133 (N_44133,N_40354,N_41613);
and U44134 (N_44134,N_40041,N_41535);
nand U44135 (N_44135,N_40546,N_41548);
nor U44136 (N_44136,N_40302,N_42418);
and U44137 (N_44137,N_41399,N_41078);
nand U44138 (N_44138,N_41505,N_41339);
nor U44139 (N_44139,N_40943,N_41985);
nand U44140 (N_44140,N_41936,N_42023);
and U44141 (N_44141,N_42254,N_41356);
or U44142 (N_44142,N_42233,N_40804);
or U44143 (N_44143,N_41909,N_42266);
or U44144 (N_44144,N_40210,N_42231);
nor U44145 (N_44145,N_40547,N_42419);
nor U44146 (N_44146,N_40327,N_40381);
and U44147 (N_44147,N_40162,N_42343);
nand U44148 (N_44148,N_40425,N_40467);
nand U44149 (N_44149,N_40283,N_42052);
nor U44150 (N_44150,N_41520,N_40912);
and U44151 (N_44151,N_41368,N_41489);
xor U44152 (N_44152,N_41107,N_40367);
xor U44153 (N_44153,N_40308,N_40206);
and U44154 (N_44154,N_41841,N_42255);
or U44155 (N_44155,N_41803,N_42108);
xnor U44156 (N_44156,N_41843,N_41769);
or U44157 (N_44157,N_41772,N_40372);
nor U44158 (N_44158,N_40984,N_41364);
and U44159 (N_44159,N_42169,N_41576);
nand U44160 (N_44160,N_41677,N_41571);
and U44161 (N_44161,N_40435,N_41082);
nand U44162 (N_44162,N_41688,N_41642);
or U44163 (N_44163,N_41136,N_42147);
and U44164 (N_44164,N_42134,N_40614);
and U44165 (N_44165,N_42206,N_42481);
or U44166 (N_44166,N_42115,N_41812);
xnor U44167 (N_44167,N_41152,N_40065);
nor U44168 (N_44168,N_41726,N_41127);
nor U44169 (N_44169,N_40193,N_42172);
xnor U44170 (N_44170,N_40196,N_42389);
nand U44171 (N_44171,N_41820,N_41447);
xor U44172 (N_44172,N_41929,N_41320);
and U44173 (N_44173,N_41643,N_40980);
xnor U44174 (N_44174,N_42496,N_41535);
nor U44175 (N_44175,N_40011,N_41617);
nor U44176 (N_44176,N_41516,N_40131);
and U44177 (N_44177,N_40020,N_42248);
and U44178 (N_44178,N_40689,N_41519);
nand U44179 (N_44179,N_40315,N_40324);
xor U44180 (N_44180,N_40069,N_40435);
and U44181 (N_44181,N_41946,N_40732);
and U44182 (N_44182,N_40634,N_42309);
and U44183 (N_44183,N_41318,N_40893);
nor U44184 (N_44184,N_41004,N_42143);
or U44185 (N_44185,N_42441,N_41578);
or U44186 (N_44186,N_41861,N_42413);
nor U44187 (N_44187,N_40862,N_42239);
nor U44188 (N_44188,N_40266,N_40780);
nand U44189 (N_44189,N_40658,N_42433);
or U44190 (N_44190,N_41567,N_41575);
nand U44191 (N_44191,N_40031,N_40696);
nor U44192 (N_44192,N_40496,N_40309);
nor U44193 (N_44193,N_42293,N_42101);
or U44194 (N_44194,N_41850,N_40145);
nor U44195 (N_44195,N_40231,N_41010);
and U44196 (N_44196,N_40608,N_40079);
or U44197 (N_44197,N_40018,N_42380);
or U44198 (N_44198,N_41578,N_40756);
xor U44199 (N_44199,N_40841,N_41125);
or U44200 (N_44200,N_40908,N_40844);
xor U44201 (N_44201,N_40660,N_42402);
nand U44202 (N_44202,N_40537,N_41806);
nand U44203 (N_44203,N_42211,N_40303);
nor U44204 (N_44204,N_41838,N_42109);
and U44205 (N_44205,N_41281,N_42147);
or U44206 (N_44206,N_42199,N_40271);
nand U44207 (N_44207,N_41431,N_41514);
nand U44208 (N_44208,N_41310,N_42058);
xor U44209 (N_44209,N_40119,N_40242);
xor U44210 (N_44210,N_40779,N_42114);
or U44211 (N_44211,N_40871,N_41355);
xor U44212 (N_44212,N_42151,N_40307);
or U44213 (N_44213,N_42235,N_41571);
xnor U44214 (N_44214,N_40610,N_40853);
nand U44215 (N_44215,N_40343,N_40528);
and U44216 (N_44216,N_40637,N_40489);
or U44217 (N_44217,N_41982,N_40327);
nor U44218 (N_44218,N_41553,N_41228);
and U44219 (N_44219,N_40378,N_41694);
xnor U44220 (N_44220,N_42278,N_40576);
xnor U44221 (N_44221,N_41415,N_42331);
xor U44222 (N_44222,N_42285,N_40778);
xnor U44223 (N_44223,N_41529,N_42304);
xor U44224 (N_44224,N_40955,N_41721);
and U44225 (N_44225,N_41250,N_40627);
nand U44226 (N_44226,N_41571,N_40741);
nand U44227 (N_44227,N_40358,N_41548);
or U44228 (N_44228,N_40370,N_42022);
nand U44229 (N_44229,N_40709,N_40617);
nand U44230 (N_44230,N_40768,N_42399);
xnor U44231 (N_44231,N_41283,N_40954);
nor U44232 (N_44232,N_41860,N_41885);
nand U44233 (N_44233,N_40479,N_42004);
and U44234 (N_44234,N_41314,N_41777);
and U44235 (N_44235,N_42319,N_40977);
nand U44236 (N_44236,N_40533,N_41528);
and U44237 (N_44237,N_40666,N_41149);
nand U44238 (N_44238,N_40677,N_41949);
xnor U44239 (N_44239,N_40055,N_41408);
and U44240 (N_44240,N_42039,N_40020);
nor U44241 (N_44241,N_41541,N_41750);
nand U44242 (N_44242,N_40874,N_41298);
and U44243 (N_44243,N_41663,N_40326);
and U44244 (N_44244,N_41137,N_41897);
or U44245 (N_44245,N_41970,N_40337);
nor U44246 (N_44246,N_41540,N_40580);
and U44247 (N_44247,N_40995,N_40323);
or U44248 (N_44248,N_42284,N_40596);
and U44249 (N_44249,N_40907,N_42488);
and U44250 (N_44250,N_41500,N_41243);
nand U44251 (N_44251,N_42423,N_41036);
or U44252 (N_44252,N_41169,N_41316);
nand U44253 (N_44253,N_42102,N_42408);
nor U44254 (N_44254,N_41132,N_41497);
xnor U44255 (N_44255,N_41041,N_40459);
or U44256 (N_44256,N_41923,N_40189);
xnor U44257 (N_44257,N_40314,N_42022);
nand U44258 (N_44258,N_40527,N_41778);
xnor U44259 (N_44259,N_41791,N_40526);
or U44260 (N_44260,N_41573,N_41609);
xor U44261 (N_44261,N_40033,N_40520);
nor U44262 (N_44262,N_41892,N_40931);
nor U44263 (N_44263,N_42335,N_40687);
or U44264 (N_44264,N_41861,N_41787);
and U44265 (N_44265,N_42093,N_42186);
xor U44266 (N_44266,N_41543,N_40564);
and U44267 (N_44267,N_40660,N_41722);
xnor U44268 (N_44268,N_42100,N_41021);
or U44269 (N_44269,N_41504,N_42110);
or U44270 (N_44270,N_42219,N_41358);
and U44271 (N_44271,N_41477,N_41571);
xnor U44272 (N_44272,N_42306,N_42369);
nand U44273 (N_44273,N_40087,N_41370);
nor U44274 (N_44274,N_41924,N_41720);
xor U44275 (N_44275,N_42352,N_41267);
nand U44276 (N_44276,N_40026,N_41672);
nor U44277 (N_44277,N_41186,N_40252);
and U44278 (N_44278,N_40161,N_40536);
and U44279 (N_44279,N_41348,N_40880);
nand U44280 (N_44280,N_41998,N_40957);
and U44281 (N_44281,N_42334,N_42419);
nor U44282 (N_44282,N_41388,N_41949);
or U44283 (N_44283,N_41086,N_42139);
nand U44284 (N_44284,N_40696,N_40889);
or U44285 (N_44285,N_40684,N_40005);
or U44286 (N_44286,N_41124,N_40704);
or U44287 (N_44287,N_41332,N_40094);
xnor U44288 (N_44288,N_40217,N_41236);
and U44289 (N_44289,N_41288,N_41448);
or U44290 (N_44290,N_41034,N_40995);
or U44291 (N_44291,N_40471,N_40612);
or U44292 (N_44292,N_40336,N_42191);
or U44293 (N_44293,N_40800,N_41621);
nand U44294 (N_44294,N_41730,N_40101);
nand U44295 (N_44295,N_40770,N_41610);
or U44296 (N_44296,N_41591,N_41647);
nor U44297 (N_44297,N_40580,N_42397);
nor U44298 (N_44298,N_40076,N_40146);
nor U44299 (N_44299,N_42444,N_40864);
nor U44300 (N_44300,N_42427,N_40249);
nand U44301 (N_44301,N_41261,N_40168);
and U44302 (N_44302,N_42067,N_42156);
or U44303 (N_44303,N_42378,N_40523);
xor U44304 (N_44304,N_42284,N_40505);
nor U44305 (N_44305,N_42235,N_42131);
nor U44306 (N_44306,N_40839,N_40503);
xor U44307 (N_44307,N_40860,N_41634);
xnor U44308 (N_44308,N_41154,N_40960);
xnor U44309 (N_44309,N_42089,N_40678);
or U44310 (N_44310,N_42334,N_41603);
nor U44311 (N_44311,N_41969,N_40575);
nor U44312 (N_44312,N_40122,N_42285);
and U44313 (N_44313,N_41155,N_42193);
xor U44314 (N_44314,N_41030,N_41143);
or U44315 (N_44315,N_41474,N_41481);
nand U44316 (N_44316,N_42343,N_40047);
xnor U44317 (N_44317,N_41179,N_40054);
or U44318 (N_44318,N_40629,N_40063);
and U44319 (N_44319,N_40554,N_42012);
nand U44320 (N_44320,N_42241,N_41825);
or U44321 (N_44321,N_40668,N_42258);
nand U44322 (N_44322,N_41228,N_41873);
or U44323 (N_44323,N_41384,N_41550);
nand U44324 (N_44324,N_40314,N_40419);
xor U44325 (N_44325,N_41204,N_42230);
nor U44326 (N_44326,N_41800,N_41959);
xor U44327 (N_44327,N_41138,N_42292);
nor U44328 (N_44328,N_41439,N_41459);
or U44329 (N_44329,N_40089,N_41092);
nor U44330 (N_44330,N_40518,N_41238);
nand U44331 (N_44331,N_41858,N_41082);
or U44332 (N_44332,N_41797,N_40553);
xor U44333 (N_44333,N_41685,N_41591);
and U44334 (N_44334,N_41485,N_40516);
or U44335 (N_44335,N_40327,N_42084);
and U44336 (N_44336,N_42037,N_40255);
nand U44337 (N_44337,N_42069,N_40127);
nor U44338 (N_44338,N_40800,N_41632);
xnor U44339 (N_44339,N_42466,N_42054);
nand U44340 (N_44340,N_41509,N_41781);
or U44341 (N_44341,N_40195,N_41721);
nand U44342 (N_44342,N_40318,N_40121);
nor U44343 (N_44343,N_40211,N_41649);
or U44344 (N_44344,N_40886,N_40170);
or U44345 (N_44345,N_40527,N_41051);
nor U44346 (N_44346,N_40437,N_42063);
nand U44347 (N_44347,N_41423,N_40545);
and U44348 (N_44348,N_42282,N_40096);
nor U44349 (N_44349,N_41255,N_41818);
nor U44350 (N_44350,N_40981,N_40851);
xor U44351 (N_44351,N_41115,N_40275);
or U44352 (N_44352,N_42140,N_41201);
nand U44353 (N_44353,N_40401,N_42075);
xor U44354 (N_44354,N_40153,N_41021);
nor U44355 (N_44355,N_42337,N_41398);
and U44356 (N_44356,N_41637,N_42371);
nand U44357 (N_44357,N_40567,N_40248);
or U44358 (N_44358,N_41678,N_40288);
xor U44359 (N_44359,N_40818,N_40312);
nand U44360 (N_44360,N_42147,N_40752);
and U44361 (N_44361,N_41531,N_41003);
nand U44362 (N_44362,N_41950,N_40468);
nor U44363 (N_44363,N_42424,N_40761);
xnor U44364 (N_44364,N_40249,N_40203);
nand U44365 (N_44365,N_40748,N_42414);
or U44366 (N_44366,N_41081,N_40087);
and U44367 (N_44367,N_40195,N_40565);
and U44368 (N_44368,N_41220,N_40530);
and U44369 (N_44369,N_40355,N_40017);
xnor U44370 (N_44370,N_40090,N_42435);
nor U44371 (N_44371,N_41214,N_42445);
and U44372 (N_44372,N_41334,N_40701);
nor U44373 (N_44373,N_40117,N_40378);
nor U44374 (N_44374,N_41076,N_40192);
nor U44375 (N_44375,N_40485,N_40533);
or U44376 (N_44376,N_40175,N_40307);
and U44377 (N_44377,N_41067,N_42364);
nand U44378 (N_44378,N_42136,N_40457);
and U44379 (N_44379,N_41863,N_40554);
nand U44380 (N_44380,N_40310,N_41867);
or U44381 (N_44381,N_40858,N_41976);
xnor U44382 (N_44382,N_41754,N_40082);
or U44383 (N_44383,N_42325,N_41395);
or U44384 (N_44384,N_40834,N_41713);
and U44385 (N_44385,N_40365,N_41967);
nor U44386 (N_44386,N_41316,N_40773);
and U44387 (N_44387,N_40426,N_42360);
or U44388 (N_44388,N_40607,N_40152);
nand U44389 (N_44389,N_40946,N_42012);
and U44390 (N_44390,N_41218,N_42469);
nand U44391 (N_44391,N_42389,N_40023);
and U44392 (N_44392,N_42017,N_40079);
nand U44393 (N_44393,N_40806,N_41277);
xor U44394 (N_44394,N_40498,N_40628);
nor U44395 (N_44395,N_40917,N_41207);
or U44396 (N_44396,N_41231,N_40916);
nor U44397 (N_44397,N_41158,N_42173);
nor U44398 (N_44398,N_40441,N_40343);
nand U44399 (N_44399,N_40407,N_40346);
nand U44400 (N_44400,N_40706,N_41657);
xor U44401 (N_44401,N_41682,N_40242);
nor U44402 (N_44402,N_41959,N_40189);
xnor U44403 (N_44403,N_40727,N_40097);
and U44404 (N_44404,N_40913,N_41432);
xnor U44405 (N_44405,N_40605,N_40420);
nor U44406 (N_44406,N_41639,N_41392);
or U44407 (N_44407,N_41442,N_42450);
and U44408 (N_44408,N_40234,N_41234);
and U44409 (N_44409,N_42145,N_42023);
nand U44410 (N_44410,N_40251,N_40800);
or U44411 (N_44411,N_41351,N_41402);
and U44412 (N_44412,N_41276,N_40074);
nand U44413 (N_44413,N_40241,N_40812);
xnor U44414 (N_44414,N_40784,N_42293);
and U44415 (N_44415,N_40597,N_41078);
or U44416 (N_44416,N_41573,N_42471);
nand U44417 (N_44417,N_42062,N_40590);
nor U44418 (N_44418,N_41720,N_40822);
nand U44419 (N_44419,N_42439,N_41725);
xor U44420 (N_44420,N_40143,N_41030);
nor U44421 (N_44421,N_41110,N_40865);
xor U44422 (N_44422,N_41249,N_40103);
nor U44423 (N_44423,N_41054,N_41370);
xnor U44424 (N_44424,N_42307,N_41691);
nor U44425 (N_44425,N_42312,N_41844);
and U44426 (N_44426,N_41239,N_40179);
or U44427 (N_44427,N_40313,N_40104);
or U44428 (N_44428,N_40946,N_41617);
and U44429 (N_44429,N_40161,N_40814);
nor U44430 (N_44430,N_41469,N_40720);
and U44431 (N_44431,N_40964,N_41371);
nand U44432 (N_44432,N_41281,N_40409);
nand U44433 (N_44433,N_41956,N_42084);
xor U44434 (N_44434,N_41992,N_40675);
or U44435 (N_44435,N_40929,N_40051);
nor U44436 (N_44436,N_42175,N_40716);
nand U44437 (N_44437,N_40821,N_40502);
nor U44438 (N_44438,N_40186,N_40494);
nand U44439 (N_44439,N_41846,N_40125);
xnor U44440 (N_44440,N_41142,N_41767);
xor U44441 (N_44441,N_40703,N_42127);
xnor U44442 (N_44442,N_40185,N_41120);
xor U44443 (N_44443,N_40885,N_42255);
nor U44444 (N_44444,N_42260,N_41444);
nor U44445 (N_44445,N_41236,N_41461);
and U44446 (N_44446,N_40792,N_42423);
and U44447 (N_44447,N_40271,N_41916);
or U44448 (N_44448,N_40492,N_41662);
nor U44449 (N_44449,N_40209,N_42192);
or U44450 (N_44450,N_40703,N_41917);
or U44451 (N_44451,N_40583,N_42482);
and U44452 (N_44452,N_41166,N_40555);
nand U44453 (N_44453,N_42015,N_41530);
nor U44454 (N_44454,N_41031,N_40629);
and U44455 (N_44455,N_42305,N_41533);
nand U44456 (N_44456,N_42331,N_41799);
nor U44457 (N_44457,N_40183,N_40725);
or U44458 (N_44458,N_40612,N_42384);
and U44459 (N_44459,N_40085,N_40969);
and U44460 (N_44460,N_42079,N_41903);
nand U44461 (N_44461,N_40809,N_40274);
or U44462 (N_44462,N_41415,N_41946);
or U44463 (N_44463,N_41096,N_42209);
and U44464 (N_44464,N_42221,N_40404);
and U44465 (N_44465,N_41395,N_41711);
or U44466 (N_44466,N_41062,N_40107);
and U44467 (N_44467,N_40061,N_41428);
nor U44468 (N_44468,N_40857,N_41089);
xor U44469 (N_44469,N_40637,N_41177);
nand U44470 (N_44470,N_41312,N_42496);
and U44471 (N_44471,N_41960,N_42300);
and U44472 (N_44472,N_40336,N_41245);
and U44473 (N_44473,N_41717,N_41706);
nand U44474 (N_44474,N_42389,N_40263);
xnor U44475 (N_44475,N_40372,N_41938);
xnor U44476 (N_44476,N_41531,N_40133);
or U44477 (N_44477,N_42193,N_40604);
and U44478 (N_44478,N_40747,N_42191);
or U44479 (N_44479,N_42326,N_40382);
nor U44480 (N_44480,N_42168,N_42255);
nand U44481 (N_44481,N_42387,N_42206);
nor U44482 (N_44482,N_40659,N_40073);
or U44483 (N_44483,N_41448,N_41166);
or U44484 (N_44484,N_40578,N_41710);
nor U44485 (N_44485,N_41722,N_41855);
xnor U44486 (N_44486,N_40805,N_42455);
nor U44487 (N_44487,N_42060,N_40918);
xor U44488 (N_44488,N_40276,N_40364);
nor U44489 (N_44489,N_41497,N_41764);
xor U44490 (N_44490,N_41401,N_41822);
or U44491 (N_44491,N_42204,N_41996);
and U44492 (N_44492,N_40470,N_42347);
nand U44493 (N_44493,N_40010,N_40150);
and U44494 (N_44494,N_41890,N_41502);
xor U44495 (N_44495,N_41802,N_41989);
and U44496 (N_44496,N_41321,N_41259);
nor U44497 (N_44497,N_40681,N_41787);
nand U44498 (N_44498,N_42103,N_41921);
nand U44499 (N_44499,N_40885,N_42254);
nor U44500 (N_44500,N_40403,N_40214);
or U44501 (N_44501,N_40946,N_41023);
nand U44502 (N_44502,N_40777,N_41264);
or U44503 (N_44503,N_40933,N_42161);
and U44504 (N_44504,N_40509,N_42454);
nor U44505 (N_44505,N_40551,N_42161);
xnor U44506 (N_44506,N_42024,N_42195);
nor U44507 (N_44507,N_42007,N_40491);
nor U44508 (N_44508,N_41757,N_40266);
and U44509 (N_44509,N_42204,N_41797);
xor U44510 (N_44510,N_40691,N_42033);
or U44511 (N_44511,N_40473,N_40460);
or U44512 (N_44512,N_40182,N_40073);
nand U44513 (N_44513,N_40086,N_40176);
or U44514 (N_44514,N_42242,N_41655);
xnor U44515 (N_44515,N_42483,N_42191);
xnor U44516 (N_44516,N_41951,N_41854);
xnor U44517 (N_44517,N_41870,N_42449);
nor U44518 (N_44518,N_41792,N_40689);
nor U44519 (N_44519,N_41054,N_40847);
and U44520 (N_44520,N_41368,N_41477);
nor U44521 (N_44521,N_41558,N_40452);
or U44522 (N_44522,N_41391,N_42065);
or U44523 (N_44523,N_41468,N_40690);
xnor U44524 (N_44524,N_41424,N_40764);
nor U44525 (N_44525,N_40227,N_42078);
nor U44526 (N_44526,N_42460,N_40645);
xnor U44527 (N_44527,N_40406,N_41118);
nor U44528 (N_44528,N_41037,N_41563);
xor U44529 (N_44529,N_40505,N_40807);
xnor U44530 (N_44530,N_42422,N_42366);
nor U44531 (N_44531,N_41785,N_41026);
nor U44532 (N_44532,N_40891,N_41161);
or U44533 (N_44533,N_41869,N_41892);
nor U44534 (N_44534,N_42084,N_41149);
nor U44535 (N_44535,N_40827,N_40696);
xnor U44536 (N_44536,N_40412,N_41937);
xor U44537 (N_44537,N_40032,N_41453);
and U44538 (N_44538,N_41229,N_40658);
and U44539 (N_44539,N_40986,N_40053);
nand U44540 (N_44540,N_41224,N_40384);
nor U44541 (N_44541,N_41650,N_41793);
nand U44542 (N_44542,N_40147,N_42307);
nand U44543 (N_44543,N_41253,N_42432);
xor U44544 (N_44544,N_41417,N_42042);
or U44545 (N_44545,N_41655,N_41872);
xor U44546 (N_44546,N_40417,N_40298);
or U44547 (N_44547,N_41106,N_42414);
or U44548 (N_44548,N_41106,N_41211);
nand U44549 (N_44549,N_42322,N_42495);
xor U44550 (N_44550,N_40080,N_40135);
xnor U44551 (N_44551,N_40152,N_40081);
xor U44552 (N_44552,N_41774,N_42485);
nor U44553 (N_44553,N_41303,N_40555);
nand U44554 (N_44554,N_40270,N_42120);
nor U44555 (N_44555,N_41681,N_42196);
and U44556 (N_44556,N_42144,N_42413);
nor U44557 (N_44557,N_40115,N_40481);
and U44558 (N_44558,N_42434,N_40979);
nand U44559 (N_44559,N_40716,N_42116);
nand U44560 (N_44560,N_41988,N_40982);
or U44561 (N_44561,N_41001,N_41672);
nand U44562 (N_44562,N_41629,N_41783);
and U44563 (N_44563,N_42285,N_40889);
or U44564 (N_44564,N_41820,N_40520);
or U44565 (N_44565,N_40142,N_42489);
nor U44566 (N_44566,N_41029,N_41387);
or U44567 (N_44567,N_42166,N_42278);
and U44568 (N_44568,N_41493,N_40042);
and U44569 (N_44569,N_42005,N_41361);
and U44570 (N_44570,N_40497,N_41392);
and U44571 (N_44571,N_41486,N_40723);
nand U44572 (N_44572,N_41944,N_42098);
nor U44573 (N_44573,N_40443,N_40840);
xnor U44574 (N_44574,N_40716,N_41105);
or U44575 (N_44575,N_42078,N_40112);
and U44576 (N_44576,N_42121,N_42192);
nor U44577 (N_44577,N_41744,N_41727);
and U44578 (N_44578,N_40372,N_42056);
xor U44579 (N_44579,N_41074,N_40114);
and U44580 (N_44580,N_41096,N_41697);
nand U44581 (N_44581,N_41235,N_41915);
xor U44582 (N_44582,N_40804,N_40188);
nor U44583 (N_44583,N_41058,N_42166);
or U44584 (N_44584,N_42479,N_40722);
and U44585 (N_44585,N_41381,N_40446);
or U44586 (N_44586,N_40751,N_40125);
xor U44587 (N_44587,N_41510,N_42400);
and U44588 (N_44588,N_41809,N_40411);
nand U44589 (N_44589,N_41798,N_41599);
nor U44590 (N_44590,N_41007,N_42178);
xnor U44591 (N_44591,N_41480,N_41229);
or U44592 (N_44592,N_41009,N_41019);
or U44593 (N_44593,N_41390,N_40314);
xnor U44594 (N_44594,N_40429,N_40799);
nor U44595 (N_44595,N_41089,N_42004);
xnor U44596 (N_44596,N_40235,N_41486);
xnor U44597 (N_44597,N_40333,N_41151);
nor U44598 (N_44598,N_42090,N_42410);
or U44599 (N_44599,N_41488,N_41642);
xnor U44600 (N_44600,N_40874,N_40457);
nand U44601 (N_44601,N_42286,N_40854);
and U44602 (N_44602,N_41492,N_41305);
or U44603 (N_44603,N_40163,N_41454);
nor U44604 (N_44604,N_40547,N_40851);
xor U44605 (N_44605,N_40388,N_42359);
nor U44606 (N_44606,N_41708,N_41606);
nor U44607 (N_44607,N_40325,N_41303);
nor U44608 (N_44608,N_40642,N_40263);
nor U44609 (N_44609,N_40893,N_42450);
xnor U44610 (N_44610,N_42320,N_41729);
nand U44611 (N_44611,N_41505,N_42236);
and U44612 (N_44612,N_41556,N_40943);
nand U44613 (N_44613,N_40941,N_42483);
xnor U44614 (N_44614,N_42007,N_42391);
nor U44615 (N_44615,N_42400,N_41549);
nand U44616 (N_44616,N_41415,N_41900);
xor U44617 (N_44617,N_40780,N_41495);
or U44618 (N_44618,N_42336,N_41670);
nand U44619 (N_44619,N_41115,N_40776);
nor U44620 (N_44620,N_40560,N_40786);
xnor U44621 (N_44621,N_40722,N_40501);
nor U44622 (N_44622,N_40270,N_40674);
nand U44623 (N_44623,N_42130,N_42051);
or U44624 (N_44624,N_40312,N_42328);
xor U44625 (N_44625,N_41879,N_40968);
nor U44626 (N_44626,N_40086,N_40600);
nand U44627 (N_44627,N_40993,N_42164);
nand U44628 (N_44628,N_41814,N_42380);
nand U44629 (N_44629,N_40461,N_42082);
or U44630 (N_44630,N_41695,N_40637);
or U44631 (N_44631,N_41203,N_40174);
and U44632 (N_44632,N_40775,N_41175);
and U44633 (N_44633,N_41959,N_40965);
nand U44634 (N_44634,N_40675,N_41683);
nand U44635 (N_44635,N_40380,N_40305);
and U44636 (N_44636,N_40800,N_42414);
and U44637 (N_44637,N_41879,N_41660);
xnor U44638 (N_44638,N_41866,N_40839);
xor U44639 (N_44639,N_42047,N_41373);
or U44640 (N_44640,N_41443,N_41862);
and U44641 (N_44641,N_40915,N_41857);
xnor U44642 (N_44642,N_42415,N_41794);
and U44643 (N_44643,N_40552,N_41212);
and U44644 (N_44644,N_42392,N_42068);
xnor U44645 (N_44645,N_41490,N_40085);
xnor U44646 (N_44646,N_40478,N_41854);
nand U44647 (N_44647,N_40355,N_42472);
nand U44648 (N_44648,N_40343,N_40825);
or U44649 (N_44649,N_40589,N_41939);
or U44650 (N_44650,N_40017,N_42048);
xnor U44651 (N_44651,N_41813,N_41622);
nand U44652 (N_44652,N_40854,N_41038);
and U44653 (N_44653,N_41835,N_40666);
nand U44654 (N_44654,N_40691,N_41585);
nor U44655 (N_44655,N_40787,N_41088);
nand U44656 (N_44656,N_40570,N_42423);
xnor U44657 (N_44657,N_41808,N_41369);
nand U44658 (N_44658,N_41210,N_40237);
and U44659 (N_44659,N_41644,N_40008);
and U44660 (N_44660,N_41099,N_41425);
and U44661 (N_44661,N_41094,N_42263);
nand U44662 (N_44662,N_40470,N_41829);
nor U44663 (N_44663,N_40558,N_41253);
nand U44664 (N_44664,N_40644,N_41673);
xnor U44665 (N_44665,N_40881,N_42003);
and U44666 (N_44666,N_40786,N_41406);
and U44667 (N_44667,N_42100,N_40364);
nor U44668 (N_44668,N_40292,N_42371);
and U44669 (N_44669,N_40226,N_41937);
nand U44670 (N_44670,N_41481,N_40757);
or U44671 (N_44671,N_42374,N_41229);
or U44672 (N_44672,N_40438,N_42270);
nor U44673 (N_44673,N_42305,N_42457);
nand U44674 (N_44674,N_41266,N_41375);
or U44675 (N_44675,N_40000,N_41419);
xnor U44676 (N_44676,N_41764,N_41975);
xor U44677 (N_44677,N_40479,N_41015);
or U44678 (N_44678,N_41444,N_42322);
nor U44679 (N_44679,N_42297,N_40293);
and U44680 (N_44680,N_41545,N_40153);
xnor U44681 (N_44681,N_40800,N_40057);
and U44682 (N_44682,N_42176,N_42497);
nand U44683 (N_44683,N_42081,N_40953);
and U44684 (N_44684,N_42341,N_41391);
or U44685 (N_44685,N_40328,N_41296);
nand U44686 (N_44686,N_41855,N_41371);
nand U44687 (N_44687,N_41544,N_41285);
and U44688 (N_44688,N_40801,N_40181);
nor U44689 (N_44689,N_42427,N_42277);
nor U44690 (N_44690,N_40748,N_40755);
nand U44691 (N_44691,N_41495,N_41507);
and U44692 (N_44692,N_41705,N_41298);
or U44693 (N_44693,N_40217,N_40672);
nor U44694 (N_44694,N_40051,N_40585);
or U44695 (N_44695,N_41250,N_40377);
nor U44696 (N_44696,N_40912,N_41834);
or U44697 (N_44697,N_41668,N_42056);
and U44698 (N_44698,N_40488,N_42182);
xnor U44699 (N_44699,N_42155,N_40788);
or U44700 (N_44700,N_41834,N_40930);
or U44701 (N_44701,N_40286,N_42013);
xor U44702 (N_44702,N_40691,N_41568);
or U44703 (N_44703,N_40620,N_41097);
nand U44704 (N_44704,N_40802,N_41756);
nand U44705 (N_44705,N_41232,N_40250);
or U44706 (N_44706,N_41795,N_40188);
xor U44707 (N_44707,N_41893,N_41599);
nor U44708 (N_44708,N_41039,N_41889);
nor U44709 (N_44709,N_41123,N_40625);
and U44710 (N_44710,N_41132,N_41334);
nand U44711 (N_44711,N_40487,N_40932);
nand U44712 (N_44712,N_40359,N_40527);
nand U44713 (N_44713,N_40714,N_41063);
and U44714 (N_44714,N_42036,N_40827);
or U44715 (N_44715,N_41034,N_40925);
nand U44716 (N_44716,N_42400,N_42318);
or U44717 (N_44717,N_40642,N_41040);
xor U44718 (N_44718,N_40634,N_42342);
nand U44719 (N_44719,N_40464,N_40446);
nor U44720 (N_44720,N_40195,N_41799);
xnor U44721 (N_44721,N_41027,N_40704);
nor U44722 (N_44722,N_40821,N_40900);
nor U44723 (N_44723,N_40934,N_40048);
xor U44724 (N_44724,N_40200,N_40497);
and U44725 (N_44725,N_41112,N_40119);
or U44726 (N_44726,N_41524,N_41354);
nor U44727 (N_44727,N_40388,N_41097);
nand U44728 (N_44728,N_40476,N_42219);
nand U44729 (N_44729,N_40827,N_41667);
xor U44730 (N_44730,N_40359,N_40202);
xor U44731 (N_44731,N_41111,N_41745);
xnor U44732 (N_44732,N_40399,N_40864);
xnor U44733 (N_44733,N_42056,N_42349);
nand U44734 (N_44734,N_40370,N_42333);
or U44735 (N_44735,N_41454,N_40475);
and U44736 (N_44736,N_42290,N_41248);
nand U44737 (N_44737,N_41502,N_41802);
nor U44738 (N_44738,N_41492,N_42018);
or U44739 (N_44739,N_41020,N_40017);
nor U44740 (N_44740,N_41862,N_41138);
or U44741 (N_44741,N_41634,N_40051);
nand U44742 (N_44742,N_40675,N_42157);
and U44743 (N_44743,N_40118,N_41591);
xnor U44744 (N_44744,N_41590,N_41532);
xnor U44745 (N_44745,N_42301,N_42398);
nand U44746 (N_44746,N_40312,N_40577);
xnor U44747 (N_44747,N_40228,N_41121);
and U44748 (N_44748,N_40078,N_42236);
nand U44749 (N_44749,N_41907,N_42408);
or U44750 (N_44750,N_41531,N_41750);
or U44751 (N_44751,N_41243,N_41850);
nor U44752 (N_44752,N_40400,N_40375);
nand U44753 (N_44753,N_41370,N_40387);
nand U44754 (N_44754,N_40133,N_42049);
nand U44755 (N_44755,N_41640,N_42262);
or U44756 (N_44756,N_40740,N_40134);
or U44757 (N_44757,N_41561,N_42463);
nand U44758 (N_44758,N_41790,N_41847);
nand U44759 (N_44759,N_41321,N_41867);
and U44760 (N_44760,N_40358,N_40680);
and U44761 (N_44761,N_41258,N_42314);
nand U44762 (N_44762,N_41685,N_41868);
nor U44763 (N_44763,N_40128,N_42168);
nor U44764 (N_44764,N_41543,N_40397);
xnor U44765 (N_44765,N_40440,N_41386);
nand U44766 (N_44766,N_40210,N_41677);
nand U44767 (N_44767,N_40869,N_41839);
or U44768 (N_44768,N_42237,N_41698);
or U44769 (N_44769,N_42434,N_42338);
xor U44770 (N_44770,N_42235,N_41432);
nor U44771 (N_44771,N_41731,N_41426);
or U44772 (N_44772,N_40689,N_41464);
and U44773 (N_44773,N_40659,N_41519);
xor U44774 (N_44774,N_42065,N_41977);
nor U44775 (N_44775,N_42452,N_40567);
and U44776 (N_44776,N_40043,N_40445);
nand U44777 (N_44777,N_40162,N_41852);
nand U44778 (N_44778,N_42273,N_41637);
or U44779 (N_44779,N_41350,N_40679);
or U44780 (N_44780,N_42473,N_41590);
xnor U44781 (N_44781,N_41154,N_42258);
xnor U44782 (N_44782,N_41699,N_41979);
and U44783 (N_44783,N_41029,N_41422);
xor U44784 (N_44784,N_41167,N_41381);
xor U44785 (N_44785,N_41022,N_41741);
and U44786 (N_44786,N_41227,N_41559);
xnor U44787 (N_44787,N_42400,N_40083);
and U44788 (N_44788,N_41836,N_41353);
or U44789 (N_44789,N_41558,N_40435);
and U44790 (N_44790,N_41998,N_42356);
xor U44791 (N_44791,N_41016,N_40061);
and U44792 (N_44792,N_41367,N_42027);
nand U44793 (N_44793,N_41669,N_40491);
or U44794 (N_44794,N_41802,N_40959);
nor U44795 (N_44795,N_40256,N_40492);
nor U44796 (N_44796,N_42269,N_41237);
and U44797 (N_44797,N_41055,N_40151);
nand U44798 (N_44798,N_40935,N_40656);
and U44799 (N_44799,N_40818,N_41231);
and U44800 (N_44800,N_40431,N_42405);
nand U44801 (N_44801,N_41413,N_41847);
or U44802 (N_44802,N_40042,N_42257);
xor U44803 (N_44803,N_41458,N_41943);
nand U44804 (N_44804,N_41102,N_41608);
nor U44805 (N_44805,N_42160,N_40408);
or U44806 (N_44806,N_40550,N_40886);
xor U44807 (N_44807,N_42111,N_40916);
or U44808 (N_44808,N_42435,N_40158);
or U44809 (N_44809,N_41247,N_42418);
nand U44810 (N_44810,N_40638,N_40253);
and U44811 (N_44811,N_40826,N_41040);
and U44812 (N_44812,N_42001,N_42342);
and U44813 (N_44813,N_41718,N_41183);
nor U44814 (N_44814,N_41526,N_40854);
and U44815 (N_44815,N_40202,N_41107);
or U44816 (N_44816,N_42481,N_40094);
xnor U44817 (N_44817,N_42302,N_40708);
and U44818 (N_44818,N_41338,N_41961);
xor U44819 (N_44819,N_41335,N_42311);
xnor U44820 (N_44820,N_41046,N_41745);
nor U44821 (N_44821,N_41652,N_42416);
nand U44822 (N_44822,N_42254,N_41286);
xnor U44823 (N_44823,N_41086,N_40831);
nor U44824 (N_44824,N_40098,N_40963);
xor U44825 (N_44825,N_42399,N_40259);
xor U44826 (N_44826,N_41117,N_41050);
or U44827 (N_44827,N_40302,N_41165);
nor U44828 (N_44828,N_42340,N_40886);
nor U44829 (N_44829,N_40347,N_40901);
nor U44830 (N_44830,N_41557,N_40859);
nand U44831 (N_44831,N_40181,N_41357);
nand U44832 (N_44832,N_40940,N_42057);
nor U44833 (N_44833,N_40069,N_40087);
and U44834 (N_44834,N_41652,N_41928);
xnor U44835 (N_44835,N_42058,N_42040);
and U44836 (N_44836,N_40899,N_41060);
or U44837 (N_44837,N_41834,N_42485);
xnor U44838 (N_44838,N_40207,N_41447);
and U44839 (N_44839,N_40684,N_40992);
xnor U44840 (N_44840,N_40836,N_41647);
or U44841 (N_44841,N_41560,N_41889);
and U44842 (N_44842,N_40308,N_42311);
and U44843 (N_44843,N_40236,N_41184);
nand U44844 (N_44844,N_41317,N_42497);
nand U44845 (N_44845,N_40431,N_40934);
and U44846 (N_44846,N_41260,N_42218);
or U44847 (N_44847,N_42062,N_41193);
xor U44848 (N_44848,N_40813,N_40126);
xnor U44849 (N_44849,N_41336,N_42415);
nor U44850 (N_44850,N_40089,N_41729);
nor U44851 (N_44851,N_41309,N_40184);
nand U44852 (N_44852,N_41515,N_42116);
nor U44853 (N_44853,N_42247,N_41803);
nand U44854 (N_44854,N_40370,N_41682);
xor U44855 (N_44855,N_42057,N_40648);
xnor U44856 (N_44856,N_42493,N_41274);
nand U44857 (N_44857,N_42262,N_40028);
nand U44858 (N_44858,N_41887,N_41767);
xor U44859 (N_44859,N_40100,N_41177);
nand U44860 (N_44860,N_41240,N_41872);
or U44861 (N_44861,N_40888,N_40946);
and U44862 (N_44862,N_41034,N_40093);
nor U44863 (N_44863,N_41950,N_42238);
nor U44864 (N_44864,N_41054,N_40551);
and U44865 (N_44865,N_41695,N_41871);
nor U44866 (N_44866,N_41863,N_40728);
and U44867 (N_44867,N_40024,N_40686);
or U44868 (N_44868,N_41914,N_40823);
and U44869 (N_44869,N_41429,N_42167);
nor U44870 (N_44870,N_41269,N_41353);
and U44871 (N_44871,N_40151,N_40623);
nand U44872 (N_44872,N_40129,N_40757);
or U44873 (N_44873,N_41533,N_40244);
and U44874 (N_44874,N_40336,N_41004);
nand U44875 (N_44875,N_40974,N_40965);
nand U44876 (N_44876,N_40655,N_41312);
and U44877 (N_44877,N_40976,N_41463);
and U44878 (N_44878,N_40200,N_40417);
nand U44879 (N_44879,N_41618,N_40404);
and U44880 (N_44880,N_41034,N_41549);
nand U44881 (N_44881,N_41251,N_41388);
or U44882 (N_44882,N_40140,N_41431);
nand U44883 (N_44883,N_42082,N_41254);
nand U44884 (N_44884,N_42259,N_41597);
nor U44885 (N_44885,N_42220,N_42339);
and U44886 (N_44886,N_40173,N_41364);
xnor U44887 (N_44887,N_40814,N_40408);
or U44888 (N_44888,N_41744,N_40857);
nor U44889 (N_44889,N_42091,N_40192);
or U44890 (N_44890,N_41896,N_40971);
xnor U44891 (N_44891,N_40189,N_40557);
or U44892 (N_44892,N_40015,N_41457);
or U44893 (N_44893,N_41021,N_40602);
and U44894 (N_44894,N_40753,N_41075);
nand U44895 (N_44895,N_40814,N_41932);
and U44896 (N_44896,N_41646,N_41069);
or U44897 (N_44897,N_42102,N_41462);
nor U44898 (N_44898,N_41275,N_41129);
nor U44899 (N_44899,N_41237,N_40586);
or U44900 (N_44900,N_42420,N_40089);
and U44901 (N_44901,N_40462,N_42262);
nor U44902 (N_44902,N_41076,N_40148);
or U44903 (N_44903,N_41458,N_40944);
and U44904 (N_44904,N_41669,N_41730);
nor U44905 (N_44905,N_40756,N_42074);
xnor U44906 (N_44906,N_41819,N_41785);
nand U44907 (N_44907,N_40127,N_40581);
and U44908 (N_44908,N_40667,N_41691);
xnor U44909 (N_44909,N_41153,N_41951);
xor U44910 (N_44910,N_40388,N_41626);
nand U44911 (N_44911,N_41247,N_40766);
xnor U44912 (N_44912,N_40516,N_41516);
and U44913 (N_44913,N_40009,N_40353);
nor U44914 (N_44914,N_41189,N_41632);
xor U44915 (N_44915,N_40548,N_41416);
or U44916 (N_44916,N_41499,N_41456);
and U44917 (N_44917,N_41989,N_40276);
and U44918 (N_44918,N_42238,N_42227);
and U44919 (N_44919,N_41249,N_41906);
nor U44920 (N_44920,N_40007,N_41364);
nand U44921 (N_44921,N_41835,N_41692);
and U44922 (N_44922,N_41200,N_41070);
and U44923 (N_44923,N_40618,N_42464);
nor U44924 (N_44924,N_42375,N_41844);
or U44925 (N_44925,N_42134,N_41744);
nor U44926 (N_44926,N_41560,N_41325);
nand U44927 (N_44927,N_40660,N_40792);
nor U44928 (N_44928,N_41501,N_41675);
nand U44929 (N_44929,N_40130,N_42392);
xor U44930 (N_44930,N_40237,N_41242);
nor U44931 (N_44931,N_40135,N_41784);
and U44932 (N_44932,N_41706,N_40635);
nor U44933 (N_44933,N_41729,N_41981);
xor U44934 (N_44934,N_41462,N_42260);
or U44935 (N_44935,N_42450,N_40157);
or U44936 (N_44936,N_41980,N_40707);
or U44937 (N_44937,N_41578,N_40454);
nand U44938 (N_44938,N_41786,N_40758);
nor U44939 (N_44939,N_41187,N_40071);
or U44940 (N_44940,N_41152,N_42477);
nor U44941 (N_44941,N_40579,N_40062);
or U44942 (N_44942,N_40568,N_40230);
or U44943 (N_44943,N_42181,N_42323);
nor U44944 (N_44944,N_41098,N_41475);
or U44945 (N_44945,N_41999,N_41545);
xor U44946 (N_44946,N_40901,N_42206);
and U44947 (N_44947,N_40461,N_40627);
nand U44948 (N_44948,N_40333,N_40206);
xor U44949 (N_44949,N_41536,N_42134);
or U44950 (N_44950,N_41815,N_40191);
nor U44951 (N_44951,N_40341,N_41578);
or U44952 (N_44952,N_41217,N_41426);
and U44953 (N_44953,N_42431,N_42199);
nor U44954 (N_44954,N_41381,N_40943);
nor U44955 (N_44955,N_41602,N_41713);
nor U44956 (N_44956,N_41983,N_40202);
nor U44957 (N_44957,N_40684,N_42163);
nor U44958 (N_44958,N_40057,N_40920);
or U44959 (N_44959,N_40468,N_40091);
or U44960 (N_44960,N_41236,N_40342);
nor U44961 (N_44961,N_40060,N_41135);
xnor U44962 (N_44962,N_41053,N_42484);
xnor U44963 (N_44963,N_41975,N_41139);
nand U44964 (N_44964,N_40142,N_41025);
xnor U44965 (N_44965,N_40154,N_41380);
and U44966 (N_44966,N_41458,N_42316);
and U44967 (N_44967,N_40458,N_40883);
and U44968 (N_44968,N_40998,N_40944);
xor U44969 (N_44969,N_42348,N_42384);
nor U44970 (N_44970,N_42461,N_41090);
nor U44971 (N_44971,N_41118,N_40023);
nand U44972 (N_44972,N_41530,N_41961);
nor U44973 (N_44973,N_42263,N_40383);
nand U44974 (N_44974,N_41554,N_40968);
and U44975 (N_44975,N_40332,N_41264);
nand U44976 (N_44976,N_42291,N_42279);
nor U44977 (N_44977,N_41011,N_40773);
nand U44978 (N_44978,N_40446,N_40793);
nor U44979 (N_44979,N_40708,N_41211);
nand U44980 (N_44980,N_42471,N_40690);
xor U44981 (N_44981,N_41041,N_41899);
or U44982 (N_44982,N_42042,N_41766);
and U44983 (N_44983,N_40305,N_40845);
nand U44984 (N_44984,N_40429,N_40009);
and U44985 (N_44985,N_40093,N_41009);
xnor U44986 (N_44986,N_41111,N_41223);
and U44987 (N_44987,N_42305,N_40414);
xnor U44988 (N_44988,N_41160,N_42232);
nand U44989 (N_44989,N_40405,N_40484);
or U44990 (N_44990,N_41832,N_40403);
and U44991 (N_44991,N_41966,N_40126);
xnor U44992 (N_44992,N_40812,N_40500);
or U44993 (N_44993,N_40518,N_42480);
or U44994 (N_44994,N_40546,N_40610);
or U44995 (N_44995,N_41696,N_41112);
and U44996 (N_44996,N_40655,N_41199);
and U44997 (N_44997,N_40963,N_40601);
xor U44998 (N_44998,N_40279,N_41571);
nor U44999 (N_44999,N_40203,N_41203);
nand U45000 (N_45000,N_43793,N_44925);
and U45001 (N_45001,N_44632,N_44056);
xnor U45002 (N_45002,N_43986,N_43437);
nand U45003 (N_45003,N_44391,N_42758);
nand U45004 (N_45004,N_44902,N_43252);
nand U45005 (N_45005,N_42577,N_42948);
nand U45006 (N_45006,N_43739,N_43085);
nor U45007 (N_45007,N_42616,N_44170);
and U45008 (N_45008,N_43471,N_44659);
or U45009 (N_45009,N_43358,N_43025);
nand U45010 (N_45010,N_43428,N_44145);
or U45011 (N_45011,N_44096,N_44641);
nand U45012 (N_45012,N_42505,N_43960);
nand U45013 (N_45013,N_42870,N_44859);
xor U45014 (N_45014,N_43074,N_43187);
xnor U45015 (N_45015,N_43152,N_42843);
nor U45016 (N_45016,N_43936,N_43422);
nor U45017 (N_45017,N_43202,N_42744);
xnor U45018 (N_45018,N_44916,N_43811);
nand U45019 (N_45019,N_43657,N_43041);
nor U45020 (N_45020,N_43978,N_44546);
nor U45021 (N_45021,N_43545,N_43588);
xnor U45022 (N_45022,N_44515,N_44009);
nor U45023 (N_45023,N_44273,N_43870);
and U45024 (N_45024,N_43365,N_43043);
and U45025 (N_45025,N_43660,N_43629);
nor U45026 (N_45026,N_44032,N_43408);
xor U45027 (N_45027,N_43664,N_44441);
or U45028 (N_45028,N_43779,N_44123);
or U45029 (N_45029,N_43282,N_44443);
or U45030 (N_45030,N_42919,N_43393);
or U45031 (N_45031,N_43760,N_44351);
or U45032 (N_45032,N_42699,N_42680);
nand U45033 (N_45033,N_44678,N_42994);
xnor U45034 (N_45034,N_44476,N_43906);
nor U45035 (N_45035,N_44864,N_43119);
nor U45036 (N_45036,N_44030,N_43593);
or U45037 (N_45037,N_43353,N_44679);
nor U45038 (N_45038,N_43255,N_44188);
nand U45039 (N_45039,N_44375,N_43451);
and U45040 (N_45040,N_43191,N_43797);
nor U45041 (N_45041,N_42689,N_44027);
xnor U45042 (N_45042,N_43964,N_42816);
or U45043 (N_45043,N_43620,N_43171);
xnor U45044 (N_45044,N_43090,N_42541);
xor U45045 (N_45045,N_44656,N_44344);
nand U45046 (N_45046,N_43951,N_43616);
nor U45047 (N_45047,N_44455,N_42667);
and U45048 (N_45048,N_44177,N_43704);
xnor U45049 (N_45049,N_42598,N_43646);
or U45050 (N_45050,N_43814,N_44790);
nor U45051 (N_45051,N_44020,N_42895);
nand U45052 (N_45052,N_43264,N_43359);
or U45053 (N_45053,N_43362,N_43210);
nor U45054 (N_45054,N_44231,N_43265);
xor U45055 (N_45055,N_43898,N_42836);
and U45056 (N_45056,N_44459,N_43653);
nand U45057 (N_45057,N_42669,N_44286);
nand U45058 (N_45058,N_43744,N_43416);
nor U45059 (N_45059,N_44920,N_43027);
xnor U45060 (N_45060,N_43614,N_42537);
xor U45061 (N_45061,N_44555,N_42884);
and U45062 (N_45062,N_42708,N_44708);
nand U45063 (N_45063,N_44624,N_43999);
or U45064 (N_45064,N_44384,N_44274);
xnor U45065 (N_45065,N_44658,N_44756);
and U45066 (N_45066,N_44205,N_43435);
and U45067 (N_45067,N_43730,N_43195);
nor U45068 (N_45068,N_43968,N_44400);
nor U45069 (N_45069,N_44069,N_43763);
nor U45070 (N_45070,N_44106,N_43488);
nor U45071 (N_45071,N_43812,N_44892);
xnor U45072 (N_45072,N_43497,N_44345);
and U45073 (N_45073,N_44878,N_43843);
xnor U45074 (N_45074,N_44843,N_43256);
and U45075 (N_45075,N_44971,N_43231);
nor U45076 (N_45076,N_43444,N_43126);
xor U45077 (N_45077,N_44138,N_43272);
nand U45078 (N_45078,N_43762,N_43950);
and U45079 (N_45079,N_43879,N_42853);
nand U45080 (N_45080,N_43032,N_44114);
or U45081 (N_45081,N_44374,N_43016);
nand U45082 (N_45082,N_42612,N_44178);
xor U45083 (N_45083,N_43240,N_42978);
nor U45084 (N_45084,N_43735,N_43316);
nor U45085 (N_45085,N_43778,N_43295);
xor U45086 (N_45086,N_42812,N_44084);
and U45087 (N_45087,N_43273,N_43184);
or U45088 (N_45088,N_44002,N_43791);
xnor U45089 (N_45089,N_44222,N_42620);
nor U45090 (N_45090,N_44074,N_44760);
and U45091 (N_45091,N_44480,N_44039);
xor U45092 (N_45092,N_44379,N_44129);
nand U45093 (N_45093,N_44538,N_42881);
xnor U45094 (N_45094,N_43097,N_44111);
and U45095 (N_45095,N_44457,N_43692);
nor U45096 (N_45096,N_43003,N_43686);
xor U45097 (N_45097,N_44922,N_43133);
nand U45098 (N_45098,N_43918,N_42794);
nor U45099 (N_45099,N_43156,N_42628);
and U45100 (N_45100,N_44058,N_44744);
or U45101 (N_45101,N_44073,N_44752);
nor U45102 (N_45102,N_43606,N_43092);
or U45103 (N_45103,N_44448,N_42961);
or U45104 (N_45104,N_44303,N_42963);
and U45105 (N_45105,N_42516,N_43373);
nor U45106 (N_45106,N_44442,N_42518);
xnor U45107 (N_45107,N_44022,N_42769);
nand U45108 (N_45108,N_43630,N_44917);
and U45109 (N_45109,N_42522,N_44826);
or U45110 (N_45110,N_44957,N_42642);
nand U45111 (N_45111,N_44028,N_43239);
nor U45112 (N_45112,N_44890,N_44246);
or U45113 (N_45113,N_43904,N_44288);
or U45114 (N_45114,N_44095,N_44031);
nand U45115 (N_45115,N_44169,N_42572);
nand U45116 (N_45116,N_43648,N_42707);
nand U45117 (N_45117,N_44425,N_44268);
xor U45118 (N_45118,N_43542,N_43350);
nand U45119 (N_45119,N_44521,N_42539);
or U45120 (N_45120,N_44429,N_44665);
xor U45121 (N_45121,N_43182,N_44849);
nand U45122 (N_45122,N_43116,N_43123);
and U45123 (N_45123,N_44600,N_44766);
and U45124 (N_45124,N_42914,N_43626);
nand U45125 (N_45125,N_43607,N_43439);
xnor U45126 (N_45126,N_44065,N_42797);
or U45127 (N_45127,N_44547,N_42981);
or U45128 (N_45128,N_44907,N_43530);
nor U45129 (N_45129,N_43698,N_43882);
nor U45130 (N_45130,N_43540,N_44577);
and U45131 (N_45131,N_43312,N_44939);
and U45132 (N_45132,N_44329,N_43414);
nand U45133 (N_45133,N_44385,N_42524);
and U45134 (N_45134,N_42549,N_42988);
or U45135 (N_45135,N_42776,N_43214);
nand U45136 (N_45136,N_44104,N_43624);
or U45137 (N_45137,N_43771,N_44157);
nor U45138 (N_45138,N_43302,N_44275);
nor U45139 (N_45139,N_44047,N_43063);
nand U45140 (N_45140,N_42866,N_43463);
xnor U45141 (N_45141,N_44970,N_42998);
and U45142 (N_45142,N_42946,N_44565);
xor U45143 (N_45143,N_44540,N_44248);
and U45144 (N_45144,N_44699,N_43993);
nor U45145 (N_45145,N_42555,N_44097);
nor U45146 (N_45146,N_43315,N_44530);
xor U45147 (N_45147,N_43637,N_42611);
and U45148 (N_45148,N_44034,N_43243);
and U45149 (N_45149,N_44534,N_44083);
xnor U45150 (N_45150,N_44652,N_43233);
xor U45151 (N_45151,N_42888,N_43891);
xnor U45152 (N_45152,N_44276,N_43010);
and U45153 (N_45153,N_43389,N_43874);
nor U45154 (N_45154,N_43671,N_43107);
nand U45155 (N_45155,N_42973,N_43656);
and U45156 (N_45156,N_43561,N_44412);
or U45157 (N_45157,N_44545,N_44748);
and U45158 (N_45158,N_42875,N_44932);
and U45159 (N_45159,N_42532,N_43384);
and U45160 (N_45160,N_44691,N_44527);
and U45161 (N_45161,N_42921,N_44943);
and U45162 (N_45162,N_44332,N_43563);
nand U45163 (N_45163,N_44202,N_43232);
and U45164 (N_45164,N_43207,N_43553);
or U45165 (N_45165,N_43838,N_44848);
xnor U45166 (N_45166,N_42661,N_44264);
or U45167 (N_45167,N_43203,N_44861);
xnor U45168 (N_45168,N_44837,N_44173);
nor U45169 (N_45169,N_43851,N_44586);
and U45170 (N_45170,N_42641,N_42785);
xor U45171 (N_45171,N_43305,N_43649);
nand U45172 (N_45172,N_43903,N_43609);
nand U45173 (N_45173,N_42559,N_44589);
nor U45174 (N_45174,N_44883,N_44858);
and U45175 (N_45175,N_43959,N_42602);
nand U45176 (N_45176,N_44422,N_43114);
nor U45177 (N_45177,N_42824,N_44258);
xor U45178 (N_45178,N_43871,N_44376);
and U45179 (N_45179,N_44635,N_42639);
or U45180 (N_45180,N_42664,N_43176);
nand U45181 (N_45181,N_43714,N_43672);
nor U45182 (N_45182,N_43192,N_43493);
and U45183 (N_45183,N_43592,N_42712);
nand U45184 (N_45184,N_44423,N_42735);
nor U45185 (N_45185,N_43780,N_42803);
or U45186 (N_45186,N_43111,N_42711);
or U45187 (N_45187,N_42892,N_44751);
nor U45188 (N_45188,N_44259,N_43445);
and U45189 (N_45189,N_43004,N_43582);
and U45190 (N_45190,N_43804,N_44529);
xor U45191 (N_45191,N_44816,N_43237);
or U45192 (N_45192,N_44912,N_42774);
nor U45193 (N_45193,N_44539,N_43644);
or U45194 (N_45194,N_44889,N_43336);
xor U45195 (N_45195,N_42659,N_43100);
nor U45196 (N_45196,N_43805,N_44532);
nand U45197 (N_45197,N_43250,N_42815);
or U45198 (N_45198,N_44704,N_44280);
and U45199 (N_45199,N_42966,N_43225);
and U45200 (N_45200,N_43854,N_43684);
nand U45201 (N_45201,N_42819,N_43896);
nand U45202 (N_45202,N_43121,N_44479);
nand U45203 (N_45203,N_43566,N_43211);
or U45204 (N_45204,N_42779,N_44979);
or U45205 (N_45205,N_44301,N_44147);
nor U45206 (N_45206,N_42916,N_44763);
nand U45207 (N_45207,N_43244,N_44502);
or U45208 (N_45208,N_43460,N_42975);
nor U45209 (N_45209,N_43223,N_42786);
or U45210 (N_45210,N_43454,N_42567);
or U45211 (N_45211,N_43828,N_42780);
and U45212 (N_45212,N_44955,N_44120);
xor U45213 (N_45213,N_44124,N_42937);
and U45214 (N_45214,N_43535,N_44648);
or U45215 (N_45215,N_42514,N_43911);
or U45216 (N_45216,N_43356,N_44285);
and U45217 (N_45217,N_42727,N_44117);
nand U45218 (N_45218,N_42640,N_43743);
xor U45219 (N_45219,N_43247,N_43775);
xnor U45220 (N_45220,N_44582,N_44518);
or U45221 (N_45221,N_44828,N_44794);
or U45222 (N_45222,N_42992,N_42701);
xnor U45223 (N_45223,N_44194,N_42872);
xnor U45224 (N_45224,N_44645,N_44218);
and U45225 (N_45225,N_43505,N_42950);
nor U45226 (N_45226,N_42847,N_43822);
and U45227 (N_45227,N_44987,N_44456);
or U45228 (N_45228,N_44492,N_44711);
nor U45229 (N_45229,N_44371,N_43324);
and U45230 (N_45230,N_42897,N_43995);
xor U45231 (N_45231,N_43064,N_44976);
xor U45232 (N_45232,N_44126,N_44324);
and U45233 (N_45233,N_44315,N_44821);
and U45234 (N_45234,N_44198,N_43757);
nor U45235 (N_45235,N_44392,N_44703);
nor U45236 (N_45236,N_44846,N_44353);
nor U45237 (N_45237,N_43136,N_43059);
or U45238 (N_45238,N_43981,N_44526);
xor U45239 (N_45239,N_44747,N_43519);
nor U45240 (N_45240,N_44463,N_44511);
or U45241 (N_45241,N_42957,N_44651);
nand U45242 (N_45242,N_43155,N_43477);
or U45243 (N_45243,N_43550,N_43270);
xor U45244 (N_45244,N_43023,N_43321);
nand U45245 (N_45245,N_42827,N_44898);
xor U45246 (N_45246,N_43722,N_44099);
or U45247 (N_45247,N_42704,N_44272);
and U45248 (N_45248,N_43317,N_43222);
nand U45249 (N_45249,N_43619,N_42583);
and U45250 (N_45250,N_44396,N_43426);
nand U45251 (N_45251,N_44077,N_43813);
xor U45252 (N_45252,N_44797,N_44533);
nand U45253 (N_45253,N_42840,N_44764);
and U45254 (N_45254,N_44601,N_44851);
nand U45255 (N_45255,N_42976,N_44026);
xnor U45256 (N_45256,N_44989,N_42662);
or U45257 (N_45257,N_43260,N_42943);
xnor U45258 (N_45258,N_44444,N_43788);
nor U45259 (N_45259,N_43937,N_44298);
nor U45260 (N_45260,N_44626,N_43570);
and U45261 (N_45261,N_44486,N_44113);
or U45262 (N_45262,N_44642,N_43430);
nor U45263 (N_45263,N_44695,N_43469);
and U45264 (N_45264,N_42793,N_44404);
or U45265 (N_45265,N_43967,N_42817);
or U45266 (N_45266,N_42959,N_44478);
nand U45267 (N_45267,N_43200,N_42630);
nand U45268 (N_45268,N_42784,N_44112);
nor U45269 (N_45269,N_44269,N_44171);
nor U45270 (N_45270,N_43703,N_43761);
nor U45271 (N_45271,N_42542,N_44841);
nor U45272 (N_45272,N_44241,N_43532);
or U45273 (N_45273,N_44220,N_44776);
nor U45274 (N_45274,N_42918,N_43663);
and U45275 (N_45275,N_43832,N_43835);
xor U45276 (N_45276,N_43948,N_43777);
nand U45277 (N_45277,N_44525,N_44265);
nor U45278 (N_45278,N_42682,N_43035);
and U45279 (N_45279,N_43511,N_43015);
nand U45280 (N_45280,N_43411,N_42771);
or U45281 (N_45281,N_44578,N_43333);
nor U45282 (N_45282,N_44927,N_43522);
nor U45283 (N_45283,N_43372,N_42883);
nor U45284 (N_45284,N_44901,N_43647);
xnor U45285 (N_45285,N_42958,N_43303);
and U45286 (N_45286,N_42698,N_42731);
nor U45287 (N_45287,N_42566,N_44991);
or U45288 (N_45288,N_43106,N_42599);
nand U45289 (N_45289,N_44687,N_43881);
and U45290 (N_45290,N_44806,N_44936);
xnor U45291 (N_45291,N_43000,N_44029);
nand U45292 (N_45292,N_44913,N_43249);
xor U45293 (N_45293,N_42710,N_43745);
or U45294 (N_45294,N_42681,N_44594);
xnor U45295 (N_45295,N_44591,N_44514);
or U45296 (N_45296,N_43508,N_42561);
and U45297 (N_45297,N_43162,N_44471);
and U45298 (N_45298,N_44762,N_43533);
xor U45299 (N_45299,N_43334,N_42908);
xnor U45300 (N_45300,N_43500,N_43976);
nor U45301 (N_45301,N_43473,N_44155);
nor U45302 (N_45302,N_43067,N_43168);
and U45303 (N_45303,N_44214,N_43135);
xnor U45304 (N_45304,N_42984,N_44551);
nor U45305 (N_45305,N_42925,N_43556);
xnor U45306 (N_45306,N_44331,N_44688);
and U45307 (N_45307,N_43529,N_44761);
nand U45308 (N_45308,N_42552,N_43160);
or U45309 (N_45309,N_43687,N_44399);
nor U45310 (N_45310,N_44380,N_43901);
and U45311 (N_45311,N_42747,N_42782);
nand U45312 (N_45312,N_42829,N_43631);
nor U45313 (N_45313,N_44713,N_43710);
or U45314 (N_45314,N_44357,N_43031);
nor U45315 (N_45315,N_43355,N_44232);
and U45316 (N_45316,N_42761,N_44325);
nand U45317 (N_45317,N_43044,N_43905);
nand U45318 (N_45318,N_44720,N_42750);
nor U45319 (N_45319,N_43919,N_43515);
nand U45320 (N_45320,N_43782,N_44312);
or U45321 (N_45321,N_44394,N_44512);
nand U45322 (N_45322,N_43691,N_43888);
xor U45323 (N_45323,N_42923,N_43461);
or U45324 (N_45324,N_44543,N_43309);
xnor U45325 (N_45325,N_43039,N_43892);
nor U45326 (N_45326,N_43839,N_43907);
nor U45327 (N_45327,N_44309,N_44070);
nor U45328 (N_45328,N_44661,N_43122);
and U45329 (N_45329,N_44895,N_44307);
nor U45330 (N_45330,N_42852,N_43065);
and U45331 (N_45331,N_44544,N_44239);
nor U45332 (N_45332,N_43855,N_44715);
xor U45333 (N_45333,N_44054,N_43789);
xnor U45334 (N_45334,N_42801,N_44805);
nand U45335 (N_45335,N_43679,N_44649);
nand U45336 (N_45336,N_43987,N_43404);
and U45337 (N_45337,N_44388,N_44834);
xnor U45338 (N_45338,N_44207,N_44853);
nor U45339 (N_45339,N_44603,N_43577);
xor U45340 (N_45340,N_44235,N_44838);
or U45341 (N_45341,N_44507,N_42841);
nor U45342 (N_45342,N_44793,N_43052);
or U45343 (N_45343,N_43610,N_43875);
xnor U45344 (N_45344,N_42685,N_43559);
nor U45345 (N_45345,N_44537,N_42700);
xnor U45346 (N_45346,N_44407,N_44311);
nor U45347 (N_45347,N_44305,N_43965);
or U45348 (N_45348,N_43348,N_44436);
nand U45349 (N_45349,N_44677,N_44081);
or U45350 (N_45350,N_44004,N_43224);
xnor U45351 (N_45351,N_43028,N_44224);
nand U45352 (N_45352,N_43397,N_42676);
nand U45353 (N_45353,N_43661,N_44115);
nand U45354 (N_45354,N_42609,N_43456);
nor U45355 (N_45355,N_43680,N_43857);
or U45356 (N_45356,N_44203,N_44299);
nand U45357 (N_45357,N_43277,N_42636);
and U45358 (N_45358,N_43737,N_43758);
xor U45359 (N_45359,N_44076,N_43747);
nand U45360 (N_45360,N_42833,N_43276);
nor U45361 (N_45361,N_43831,N_44277);
xor U45362 (N_45362,N_43652,N_44005);
xnor U45363 (N_45363,N_43169,N_44962);
nor U45364 (N_45364,N_42544,N_43419);
and U45365 (N_45365,N_42519,N_44663);
nand U45366 (N_45366,N_42938,N_42821);
and U45367 (N_45367,N_43339,N_43138);
nand U45368 (N_45368,N_43022,N_44686);
xor U45369 (N_45369,N_44839,N_44014);
or U45370 (N_45370,N_43318,N_44701);
or U45371 (N_45371,N_43885,N_44079);
and U45372 (N_45372,N_44814,N_42693);
and U45373 (N_45373,N_44672,N_42755);
and U45374 (N_45374,N_43371,N_43297);
or U45375 (N_45375,N_43311,N_43554);
nand U45376 (N_45376,N_44599,N_44063);
and U45377 (N_45377,N_44675,N_44567);
nor U45378 (N_45378,N_43058,N_43980);
and U45379 (N_45379,N_43740,N_43306);
nor U45380 (N_45380,N_44775,N_44339);
nand U45381 (N_45381,N_44639,N_43257);
and U45382 (N_45382,N_44043,N_42606);
nand U45383 (N_45383,N_44745,N_44180);
nand U45384 (N_45384,N_44061,N_44416);
and U45385 (N_45385,N_44431,N_44446);
xnor U45386 (N_45386,N_44795,N_44778);
or U45387 (N_45387,N_43894,N_43693);
nor U45388 (N_45388,N_43830,N_44897);
nand U45389 (N_45389,N_44796,N_43412);
and U45390 (N_45390,N_44850,N_44882);
xnor U45391 (N_45391,N_43575,N_44614);
xor U45392 (N_45392,N_44865,N_44560);
or U45393 (N_45393,N_42979,N_44266);
nor U45394 (N_45394,N_43287,N_44042);
xor U45395 (N_45395,N_43081,N_44025);
nor U45396 (N_45396,N_44372,N_43886);
xnor U45397 (N_45397,N_44938,N_44033);
and U45398 (N_45398,N_44296,N_42718);
xnor U45399 (N_45399,N_43021,N_44992);
and U45400 (N_45400,N_43925,N_43957);
nor U45401 (N_45401,N_44464,N_43095);
nor U45402 (N_45402,N_43018,N_42533);
and U45403 (N_45403,N_43314,N_43727);
and U45404 (N_45404,N_44243,N_44852);
or U45405 (N_45405,N_44041,N_43229);
xor U45406 (N_45406,N_44712,N_43382);
or U45407 (N_45407,N_44562,N_44334);
nand U45408 (N_45408,N_43280,N_44908);
nand U45409 (N_45409,N_42590,N_44994);
nand U45410 (N_45410,N_43406,N_43185);
nor U45411 (N_45411,N_43816,N_42789);
nor U45412 (N_45412,N_44293,N_43803);
nor U45413 (N_45413,N_43285,N_44613);
or U45414 (N_45414,N_42634,N_43345);
nor U45415 (N_45415,N_42967,N_44923);
or U45416 (N_45416,N_44630,N_44705);
nand U45417 (N_45417,N_44689,N_44596);
and U45418 (N_45418,N_43707,N_44135);
or U45419 (N_45419,N_43528,N_43518);
and U45420 (N_45420,N_44341,N_44000);
and U45421 (N_45421,N_43524,N_44162);
or U45422 (N_45422,N_42756,N_44668);
or U45423 (N_45423,N_44819,N_42858);
xor U45424 (N_45424,N_43271,N_43069);
and U45425 (N_45425,N_44732,N_44267);
or U45426 (N_45426,N_44072,N_42798);
xor U45427 (N_45427,N_42969,N_42861);
xor U45428 (N_45428,N_42721,N_44433);
nor U45429 (N_45429,N_43618,N_44295);
nor U45430 (N_45430,N_42878,N_44584);
or U45431 (N_45431,N_43890,N_44383);
nand U45432 (N_45432,N_44845,N_42882);
or U45433 (N_45433,N_43713,N_44142);
nor U45434 (N_45434,N_44506,N_43066);
or U45435 (N_45435,N_43860,N_42722);
nor U45436 (N_45436,N_42927,N_42603);
nand U45437 (N_45437,N_44765,N_43926);
nor U45438 (N_45438,N_44330,N_44451);
xnor U45439 (N_45439,N_42535,N_43313);
xor U45440 (N_45440,N_44389,N_43694);
and U45441 (N_45441,N_44190,N_43706);
nor U45442 (N_45442,N_44657,N_43546);
xnor U45443 (N_45443,N_44185,N_44234);
nor U45444 (N_45444,N_44781,N_44996);
or U45445 (N_45445,N_43551,N_44051);
or U45446 (N_45446,N_44817,N_43215);
or U45447 (N_45447,N_43129,N_43982);
or U45448 (N_45448,N_42986,N_43234);
nand U45449 (N_45449,N_44815,N_43024);
or U45450 (N_45450,N_44420,N_43970);
xor U45451 (N_45451,N_44980,N_43387);
xor U45452 (N_45452,N_44857,N_44948);
nor U45453 (N_45453,N_42930,N_42551);
xnor U45454 (N_45454,N_44487,N_43494);
or U45455 (N_45455,N_42509,N_44873);
nor U45456 (N_45456,N_44333,N_44319);
nor U45457 (N_45457,N_43578,N_42538);
xnor U45458 (N_45458,N_42907,N_42868);
and U45459 (N_45459,N_44365,N_44755);
xor U45460 (N_45460,N_44974,N_42666);
nor U45461 (N_45461,N_44036,N_43405);
xor U45462 (N_45462,N_44110,N_44617);
and U45463 (N_45463,N_42586,N_42980);
nor U45464 (N_45464,N_42935,N_44789);
or U45465 (N_45465,N_44006,N_44870);
or U45466 (N_45466,N_42525,N_42691);
or U45467 (N_45467,N_44349,N_42831);
or U45468 (N_45468,N_44888,N_42517);
nand U45469 (N_45469,N_43776,N_44592);
nor U45470 (N_45470,N_44090,N_42740);
nand U45471 (N_45471,N_43292,N_43596);
and U45472 (N_45472,N_42876,N_44316);
xnor U45473 (N_45473,N_43433,N_44066);
and U45474 (N_45474,N_43047,N_42686);
and U45475 (N_45475,N_43091,N_44403);
nor U45476 (N_45476,N_43038,N_42901);
xor U45477 (N_45477,N_44482,N_43172);
or U45478 (N_45478,N_42738,N_44647);
or U45479 (N_45479,N_44395,N_42902);
or U45480 (N_45480,N_42631,N_44210);
or U45481 (N_45481,N_44508,N_44832);
nor U45482 (N_45482,N_43434,N_42655);
and U45483 (N_45483,N_42594,N_43873);
and U45484 (N_45484,N_43075,N_43351);
or U45485 (N_45485,N_43584,N_44313);
and U45486 (N_45486,N_42607,N_42762);
nor U45487 (N_45487,N_44426,N_43583);
and U45488 (N_45488,N_44767,N_43966);
nand U45489 (N_45489,N_43984,N_44103);
nand U45490 (N_45490,N_43258,N_44835);
nand U45491 (N_45491,N_44430,N_44156);
xor U45492 (N_45492,N_43983,N_43503);
and U45493 (N_45493,N_43729,N_44602);
nand U45494 (N_45494,N_43054,N_43726);
nand U45495 (N_45495,N_42777,N_42729);
or U45496 (N_45496,N_43806,N_42936);
or U45497 (N_45497,N_44595,N_44472);
and U45498 (N_45498,N_42857,N_42719);
xor U45499 (N_45499,N_44256,N_43792);
nor U45500 (N_45500,N_44460,N_44985);
xnor U45501 (N_45501,N_42818,N_43383);
and U45502 (N_45502,N_44133,N_44719);
or U45503 (N_45503,N_43701,N_43774);
nor U45504 (N_45504,N_44012,N_42972);
xor U45505 (N_45505,N_43591,N_44068);
and U45506 (N_45506,N_42800,N_44721);
or U45507 (N_45507,N_42880,N_43322);
xnor U45508 (N_45508,N_42851,N_43717);
nand U45509 (N_45509,N_44571,N_43643);
nand U45510 (N_45510,N_42996,N_42960);
xnor U45511 (N_45511,N_44271,N_43681);
nand U45512 (N_45512,N_43094,N_43056);
nor U45513 (N_45513,N_42624,N_42893);
and U45514 (N_45514,N_44187,N_42933);
nand U45515 (N_45515,N_44150,N_44951);
or U45516 (N_45516,N_44304,N_43601);
or U45517 (N_45517,N_43300,N_43893);
or U45518 (N_45518,N_44952,N_44958);
and U45519 (N_45519,N_43495,N_43576);
or U45520 (N_45520,N_43140,N_44320);
nor U45521 (N_45521,N_43246,N_44473);
nand U45522 (N_45522,N_43952,N_44812);
or U45523 (N_45523,N_42879,N_44481);
nand U45524 (N_45524,N_44730,N_43979);
and U45525 (N_45525,N_44326,N_42945);
xnor U45526 (N_45526,N_43379,N_43083);
xnor U45527 (N_45527,N_43953,N_43360);
nand U45528 (N_45528,N_42743,N_42617);
and U45529 (N_45529,N_43725,N_44310);
or U45530 (N_45530,N_43924,N_43453);
or U45531 (N_45531,N_43286,N_43705);
or U45532 (N_45532,N_44556,N_42500);
nor U45533 (N_45533,N_44450,N_42723);
or U45534 (N_45534,N_43971,N_43923);
nor U45535 (N_45535,N_44250,N_43877);
nand U45536 (N_45536,N_42553,N_43150);
xor U45537 (N_45537,N_42904,N_43988);
and U45538 (N_45538,N_43539,N_44179);
nand U45539 (N_45539,N_42545,N_44887);
and U45540 (N_45540,N_42728,N_43179);
and U45541 (N_45541,N_44726,N_43174);
xor U45542 (N_45542,N_44219,N_42865);
xnor U45543 (N_45543,N_44080,N_44386);
nand U45544 (N_45544,N_42576,N_44741);
and U45545 (N_45545,N_44753,N_43520);
and U45546 (N_45546,N_44340,N_43513);
and U45547 (N_45547,N_43392,N_44465);
nand U45548 (N_45548,N_44398,N_42554);
xor U45549 (N_45549,N_44503,N_42956);
nand U45550 (N_45550,N_44397,N_43666);
and U45551 (N_45551,N_44109,N_42949);
or U45552 (N_45552,N_43868,N_43659);
and U45553 (N_45553,N_44306,N_43254);
and U45554 (N_45554,N_43883,N_43654);
nor U45555 (N_45555,N_43565,N_44107);
and U45556 (N_45556,N_44377,N_44282);
and U45557 (N_45557,N_43751,N_43386);
nor U45558 (N_45558,N_44101,N_43946);
and U45559 (N_45559,N_44044,N_44942);
or U45560 (N_45560,N_43555,N_44566);
or U45561 (N_45561,N_43534,N_43325);
or U45562 (N_45562,N_43400,N_44322);
or U45563 (N_45563,N_44736,N_42810);
xnor U45564 (N_45564,N_44694,N_42739);
nand U45565 (N_45565,N_43450,N_42725);
nor U45566 (N_45566,N_44559,N_44364);
or U45567 (N_45567,N_44754,N_44255);
nor U45568 (N_45568,N_43772,N_43368);
nand U45569 (N_45569,N_44308,N_44035);
nand U45570 (N_45570,N_42890,N_44801);
or U45571 (N_45571,N_42652,N_42767);
nor U45572 (N_45572,N_44724,N_44137);
xor U45573 (N_45573,N_43947,N_43370);
or U45574 (N_45574,N_43079,N_42846);
and U45575 (N_45575,N_43489,N_44549);
or U45576 (N_45576,N_43259,N_43756);
nor U45577 (N_45577,N_42531,N_43177);
nor U45578 (N_45578,N_43819,N_44833);
nor U45579 (N_45579,N_43766,N_44682);
nor U45580 (N_45580,N_43699,N_44427);
and U45581 (N_45581,N_44609,N_44019);
and U45582 (N_45582,N_44884,N_43912);
nor U45583 (N_45583,N_43352,N_44130);
nor U45584 (N_45584,N_43829,N_43103);
nand U45585 (N_45585,N_43390,N_44419);
nand U45586 (N_45586,N_43800,N_43181);
or U45587 (N_45587,N_44021,N_43139);
or U45588 (N_45588,N_43677,N_44750);
xnor U45589 (N_45589,N_43622,N_43850);
or U45590 (N_45590,N_43998,N_42896);
and U45591 (N_45591,N_42802,N_44159);
nor U45592 (N_45592,N_43046,N_44911);
or U45593 (N_45593,N_42683,N_42604);
nand U45594 (N_45594,N_44439,N_44606);
and U45595 (N_45595,N_42790,N_44615);
nand U45596 (N_45596,N_42570,N_43842);
and U45597 (N_45597,N_44292,N_43034);
nand U45598 (N_45598,N_44281,N_44863);
and U45599 (N_45599,N_42696,N_44924);
or U45600 (N_45600,N_42871,N_43266);
nand U45601 (N_45601,N_42665,N_43279);
xnor U45602 (N_45602,N_42720,N_44102);
nand U45603 (N_45603,N_42928,N_44523);
and U45604 (N_45604,N_44953,N_44909);
nand U45605 (N_45605,N_43670,N_42588);
nor U45606 (N_45606,N_42990,N_43608);
and U45607 (N_45607,N_43189,N_43204);
or U45608 (N_45608,N_42621,N_44999);
nor U45609 (N_45609,N_44553,N_43146);
and U45610 (N_45610,N_43164,N_42768);
nor U45611 (N_45611,N_42637,N_43338);
nor U45612 (N_45612,N_44249,N_43221);
nor U45613 (N_45613,N_43955,N_43547);
or U45614 (N_45614,N_43665,N_44743);
or U45615 (N_45615,N_43770,N_44671);
xor U45616 (N_45616,N_44915,N_43319);
or U45617 (N_45617,N_43486,N_42703);
nor U45618 (N_45618,N_43323,N_42845);
nor U45619 (N_45619,N_42670,N_44401);
nand U45620 (N_45620,N_44964,N_42911);
nor U45621 (N_45621,N_44588,N_42856);
and U45622 (N_45622,N_44166,N_44496);
and U45623 (N_45623,N_43198,N_43628);
nor U45624 (N_45624,N_44604,N_44574);
and U45625 (N_45625,N_44702,N_42520);
and U45626 (N_45626,N_44226,N_44900);
nor U45627 (N_45627,N_44780,N_42842);
nor U45628 (N_45628,N_43824,N_44640);
and U45629 (N_45629,N_44573,N_44154);
and U45630 (N_45630,N_43634,N_43053);
nand U45631 (N_45631,N_44370,N_43235);
nand U45632 (N_45632,N_44856,N_44877);
and U45633 (N_45633,N_43787,N_44929);
and U45634 (N_45634,N_43969,N_44206);
or U45635 (N_45635,N_43543,N_42807);
nand U45636 (N_45636,N_42867,N_44728);
nand U45637 (N_45637,N_43481,N_44204);
or U45638 (N_45638,N_44820,N_43746);
nor U45639 (N_45639,N_44557,N_44983);
nor U45640 (N_45640,N_44666,N_43381);
and U45641 (N_45641,N_44469,N_43357);
or U45642 (N_45642,N_43569,N_44733);
and U45643 (N_45643,N_44491,N_42991);
or U45644 (N_45644,N_44055,N_44519);
or U45645 (N_45645,N_43636,N_44568);
nand U45646 (N_45646,N_43029,N_43178);
and U45647 (N_45647,N_43742,N_44337);
and U45648 (N_45648,N_44082,N_44140);
xnor U45649 (N_45649,N_43219,N_43394);
or U45650 (N_45650,N_44408,N_44361);
xnor U45651 (N_45651,N_42556,N_44217);
xor U45652 (N_45652,N_43042,N_44823);
or U45653 (N_45653,N_42674,N_42563);
xnor U45654 (N_45654,N_42571,N_42814);
or U45655 (N_45655,N_44017,N_43668);
nand U45656 (N_45656,N_44684,N_43175);
or U45657 (N_45657,N_44449,N_44373);
or U45658 (N_45658,N_44903,N_42909);
nor U45659 (N_45659,N_43754,N_43402);
and U45660 (N_45660,N_44535,N_42605);
or U45661 (N_45661,N_43476,N_42885);
xnor U45662 (N_45662,N_44866,N_44984);
nor U45663 (N_45663,N_43504,N_42905);
and U45664 (N_45664,N_44787,N_44064);
xor U45665 (N_45665,N_43030,N_43199);
xnor U45666 (N_45666,N_44946,N_42783);
nor U45667 (N_45667,N_44608,N_44742);
nand U45668 (N_45668,N_44490,N_42585);
nor U45669 (N_45669,N_43127,N_44788);
and U45670 (N_45670,N_42862,N_42903);
nor U45671 (N_45671,N_43994,N_43712);
and U45672 (N_45672,N_43278,N_43410);
or U45673 (N_45673,N_42732,N_43440);
nor U45674 (N_45674,N_44520,N_44139);
or U45675 (N_45675,N_42593,N_43396);
nor U45676 (N_45676,N_44875,N_43452);
or U45677 (N_45677,N_44896,N_42792);
nand U45678 (N_45678,N_44972,N_43424);
or U45679 (N_45679,N_43688,N_42715);
or U45680 (N_45680,N_42929,N_44966);
nand U45681 (N_45681,N_44045,N_42799);
nand U45682 (N_45682,N_43752,N_42684);
and U45683 (N_45683,N_42965,N_43604);
or U45684 (N_45684,N_44696,N_44784);
or U45685 (N_45685,N_43602,N_44100);
and U45686 (N_45686,N_43996,N_44252);
nor U45687 (N_45687,N_44417,N_44215);
xor U45688 (N_45688,N_43026,N_44718);
nor U45689 (N_45689,N_44590,N_44466);
or U45690 (N_45690,N_42863,N_42565);
or U45691 (N_45691,N_43263,N_42688);
nand U45692 (N_45692,N_42997,N_43864);
or U45693 (N_45693,N_44894,N_42705);
and U45694 (N_45694,N_44092,N_44247);
xnor U45695 (N_45695,N_44947,N_42772);
xor U45696 (N_45696,N_42504,N_44242);
xor U45697 (N_45697,N_43093,N_44011);
or U45698 (N_45698,N_43837,N_43033);
and U45699 (N_45699,N_43682,N_43310);
or U45700 (N_45700,N_43773,N_44452);
nor U45701 (N_45701,N_44868,N_43344);
xor U45702 (N_45702,N_44636,N_43275);
and U45703 (N_45703,N_43597,N_44148);
or U45704 (N_45704,N_44125,N_43073);
xnor U45705 (N_45705,N_44184,N_42501);
nand U45706 (N_45706,N_44993,N_42734);
xor U45707 (N_45707,N_42717,N_44230);
nor U45708 (N_45708,N_42569,N_44824);
or U45709 (N_45709,N_43599,N_43962);
xor U45710 (N_45710,N_44144,N_43961);
xor U45711 (N_45711,N_43538,N_43009);
and U45712 (N_45712,N_43230,N_43929);
nor U45713 (N_45713,N_44141,N_43149);
or U45714 (N_45714,N_44616,N_43425);
xnor U45715 (N_45715,N_44522,N_43809);
and U45716 (N_45716,N_43429,N_44517);
or U45717 (N_45717,N_42526,N_43415);
xor U45718 (N_45718,N_43696,N_44263);
nand U45719 (N_45719,N_43459,N_42742);
xnor U45720 (N_45720,N_44347,N_43834);
nand U45721 (N_45721,N_43134,N_43342);
nor U45722 (N_45722,N_43940,N_44493);
and U45723 (N_45723,N_44623,N_44654);
and U45724 (N_45724,N_42982,N_43226);
or U45725 (N_45725,N_42737,N_44680);
nor U45726 (N_45726,N_43567,N_43443);
nor U45727 (N_45727,N_44693,N_43786);
and U45728 (N_45728,N_43523,N_44289);
or U45729 (N_45729,N_44803,N_42820);
nor U45730 (N_45730,N_44418,N_44638);
xnor U45731 (N_45731,N_44619,N_43190);
and U45732 (N_45732,N_44918,N_44674);
xor U45733 (N_45733,N_44118,N_43188);
nor U45734 (N_45734,N_43755,N_44108);
xor U45735 (N_45735,N_42778,N_42912);
xor U45736 (N_45736,N_44071,N_42557);
nand U45737 (N_45737,N_44160,N_44437);
nand U45738 (N_45738,N_43335,N_42511);
nor U45739 (N_45739,N_44181,N_43484);
nor U45740 (N_45740,N_43859,N_43491);
or U45741 (N_45741,N_42974,N_43061);
and U45742 (N_45742,N_44318,N_43331);
xnor U45743 (N_45743,N_44737,N_42839);
or U45744 (N_45744,N_43212,N_44228);
nor U45745 (N_45745,N_44881,N_42964);
or U45746 (N_45746,N_43939,N_43076);
and U45747 (N_45747,N_42889,N_43045);
xnor U45748 (N_45748,N_42543,N_43262);
nor U45749 (N_45749,N_43750,N_43253);
xor U45750 (N_45750,N_44510,N_44294);
nor U45751 (N_45751,N_44008,N_44046);
xor U45752 (N_45752,N_43914,N_44683);
nor U45753 (N_45753,N_43236,N_43487);
nand U45754 (N_45754,N_43084,N_42618);
xnor U45755 (N_45755,N_44810,N_44921);
nor U45756 (N_45756,N_42579,N_43464);
nand U45757 (N_45757,N_44700,N_44057);
or U45758 (N_45758,N_43909,N_44367);
nand U45759 (N_45759,N_43974,N_42528);
and U45760 (N_45760,N_44931,N_43872);
nand U45761 (N_45761,N_42832,N_44505);
and U45762 (N_45762,N_43521,N_43008);
and U45763 (N_45763,N_42977,N_43417);
xor U45764 (N_45764,N_42764,N_42550);
nor U45765 (N_45765,N_44227,N_44569);
nor U45766 (N_45766,N_44284,N_42697);
xnor U45767 (N_45767,N_44628,N_44963);
xnor U45768 (N_45768,N_43180,N_44692);
or U45769 (N_45769,N_44414,N_43632);
nand U45770 (N_45770,N_43820,N_44738);
nor U45771 (N_45771,N_43147,N_44003);
nand U45772 (N_45772,N_43366,N_42917);
and U45773 (N_45773,N_44685,N_43594);
nor U45774 (N_45774,N_43474,N_43808);
or U45775 (N_45775,N_44769,N_44977);
or U45776 (N_45776,N_44960,N_43818);
nor U45777 (N_45777,N_43669,N_44352);
and U45778 (N_45778,N_44670,N_43132);
xnor U45779 (N_45779,N_42692,N_43077);
or U45780 (N_45780,N_44211,N_43124);
nand U45781 (N_45781,N_44279,N_44893);
nand U45782 (N_45782,N_42534,N_44673);
and U45783 (N_45783,N_43196,N_44186);
or U45784 (N_45784,N_44474,N_43101);
and U45785 (N_45785,N_43991,N_43897);
nand U45786 (N_45786,N_43759,N_44174);
nor U45787 (N_45787,N_42530,N_42788);
xor U45788 (N_45788,N_42813,N_43612);
nor U45789 (N_45789,N_43088,N_42540);
xnor U45790 (N_45790,N_42582,N_43328);
or U45791 (N_45791,N_43611,N_42626);
xnor U45792 (N_45792,N_44886,N_43407);
nor U45793 (N_45793,N_43213,N_42654);
or U45794 (N_45794,N_44676,N_43466);
and U45795 (N_45795,N_44461,N_44062);
nor U45796 (N_45796,N_42894,N_44827);
or U45797 (N_45797,N_44664,N_42968);
and U45798 (N_45798,N_44244,N_44906);
and U45799 (N_45799,N_42805,N_44758);
and U45800 (N_45800,N_44727,N_43005);
nand U45801 (N_45801,N_43662,N_43399);
and U45802 (N_45802,N_44010,N_44151);
nor U45803 (N_45803,N_42999,N_44904);
or U45804 (N_45804,N_43082,N_42724);
xnor U45805 (N_45805,N_43769,N_44260);
and U45806 (N_45806,N_43507,N_43364);
nand U45807 (N_45807,N_43595,N_44809);
and U45808 (N_45808,N_42615,N_42503);
xnor U45809 (N_45809,N_44576,N_43401);
or U45810 (N_45810,N_42864,N_42906);
or U45811 (N_45811,N_43143,N_42536);
or U45812 (N_45812,N_44818,N_44610);
xor U45813 (N_45813,N_43927,N_43330);
nor U45814 (N_45814,N_43154,N_43954);
and U45815 (N_45815,N_44193,N_44798);
xnor U45816 (N_45816,N_44413,N_43183);
nor U45817 (N_45817,N_43479,N_44934);
and U45818 (N_45818,N_43600,N_44581);
nand U45819 (N_45819,N_42922,N_44216);
and U45820 (N_45820,N_44175,N_43801);
nor U45821 (N_45821,N_43749,N_42597);
and U45822 (N_45822,N_43633,N_43764);
and U45823 (N_45823,N_43050,N_42873);
and U45824 (N_45824,N_43337,N_43012);
and U45825 (N_45825,N_43942,N_44094);
nand U45826 (N_45826,N_43549,N_42660);
xnor U45827 (N_45827,N_43472,N_43462);
nor U45828 (N_45828,N_44360,N_44462);
or U45829 (N_45829,N_43468,N_43449);
nand U45830 (N_45830,N_44053,N_42826);
xnor U45831 (N_45831,N_43349,N_44722);
or U45832 (N_45832,N_44967,N_43810);
nand U45833 (N_45833,N_42759,N_43332);
nor U45834 (N_45834,N_42855,N_43783);
and U45835 (N_45835,N_44988,N_44368);
nor U45836 (N_45836,N_42989,N_42926);
nor U45837 (N_45837,N_42589,N_43586);
nor U45838 (N_45838,N_43733,N_43625);
nor U45839 (N_45839,N_43571,N_44660);
nand U45840 (N_45840,N_44078,N_43833);
nand U45841 (N_45841,N_44200,N_42508);
xor U45842 (N_45842,N_43732,N_44593);
nor U45843 (N_45843,N_43689,N_44131);
or U45844 (N_45844,N_43963,N_44049);
and U45845 (N_45845,N_42952,N_44965);
and U45846 (N_45846,N_44143,N_42581);
and U45847 (N_45847,N_44885,N_43186);
nand U45848 (N_45848,N_42521,N_43078);
or U45849 (N_45849,N_43941,N_42601);
xnor U45850 (N_45850,N_42770,N_43037);
xor U45851 (N_45851,N_44278,N_44830);
nor U45852 (N_45852,N_42900,N_43574);
nand U45853 (N_45853,N_43673,N_42995);
xor U45854 (N_45854,N_43301,N_44773);
nand U45855 (N_45855,N_44489,N_44434);
or U45856 (N_45856,N_44997,N_42653);
nor U45857 (N_45857,N_42679,N_43836);
nor U45858 (N_45858,N_44409,N_42787);
xnor U45859 (N_45859,N_42614,N_44024);
and U45860 (N_45860,N_44725,N_43869);
and U45861 (N_45861,N_42877,N_44093);
and U45862 (N_45862,N_44323,N_42656);
or U45863 (N_45863,N_43900,N_42924);
and U45864 (N_45864,N_44808,N_43506);
and U45865 (N_45865,N_44050,N_43989);
or U45866 (N_45866,N_43548,N_44829);
nand U45867 (N_45867,N_44621,N_44023);
and U45868 (N_45868,N_42834,N_44541);
or U45869 (N_45869,N_43856,N_43720);
nor U45870 (N_45870,N_43598,N_43099);
or U45871 (N_45871,N_42837,N_44650);
or U45872 (N_45872,N_43290,N_43227);
and U45873 (N_45873,N_42749,N_43541);
or U45874 (N_45874,N_43931,N_42746);
nand U45875 (N_45875,N_42811,N_44158);
nand U45876 (N_45876,N_44643,N_44350);
nand U45877 (N_45877,N_43852,N_44802);
or U45878 (N_45878,N_44105,N_43655);
nor U45879 (N_45879,N_43639,N_43579);
nor U45880 (N_45880,N_43436,N_43294);
and U45881 (N_45881,N_43552,N_44734);
xnor U45882 (N_45882,N_43765,N_44428);
nor U45883 (N_45883,N_43956,N_43062);
nand U45884 (N_45884,N_43723,N_44362);
xor U45885 (N_45885,N_44563,N_43205);
nand U45886 (N_45886,N_43395,N_44238);
and U45887 (N_45887,N_44620,N_42643);
or U45888 (N_45888,N_43340,N_44928);
nor U45889 (N_45889,N_44653,N_44424);
nand U45890 (N_45890,N_43849,N_44136);
nor U45891 (N_45891,N_43560,N_44587);
nand U45892 (N_45892,N_44862,N_43721);
and U45893 (N_45893,N_44229,N_43446);
or U45894 (N_45894,N_42548,N_42507);
and U45895 (N_45895,N_44192,N_44941);
xor U45896 (N_45896,N_44453,N_43617);
nor U45897 (N_45897,N_43884,N_43623);
nand U45898 (N_45898,N_43442,N_42622);
nand U45899 (N_45899,N_44213,N_42745);
xor U45900 (N_45900,N_44655,N_43973);
or U45901 (N_45901,N_43327,N_42899);
or U45902 (N_45902,N_43935,N_44872);
xnor U45903 (N_45903,N_42733,N_42592);
and U45904 (N_45904,N_42702,N_42954);
xor U45905 (N_45905,N_43848,N_42632);
and U45906 (N_45906,N_43418,N_44087);
xor U45907 (N_45907,N_43346,N_42753);
nor U45908 (N_45908,N_43572,N_43251);
xor U45909 (N_45909,N_43120,N_44637);
or U45910 (N_45910,N_44607,N_42694);
nand U45911 (N_45911,N_43977,N_43173);
nand U45912 (N_45912,N_44378,N_44800);
nand U45913 (N_45913,N_44940,N_42663);
nor U45914 (N_45914,N_43403,N_42736);
and U45915 (N_45915,N_42940,N_44844);
xor U45916 (N_45916,N_44122,N_44366);
xor U45917 (N_45917,N_43421,N_44633);
and U45918 (N_45918,N_43784,N_44134);
or U45919 (N_45919,N_43369,N_43447);
nor U45920 (N_45920,N_42651,N_43475);
xnor U45921 (N_45921,N_44302,N_44225);
or U45922 (N_45922,N_42647,N_43715);
nand U45923 (N_45923,N_43562,N_43589);
nand U45924 (N_45924,N_42523,N_42587);
nand U45925 (N_45925,N_42580,N_43153);
or U45926 (N_45926,N_44874,N_42687);
and U45927 (N_45927,N_43220,N_43580);
and U45928 (N_45928,N_43413,N_43499);
nor U45929 (N_45929,N_42849,N_42910);
and U45930 (N_45930,N_44164,N_43304);
and U45931 (N_45931,N_44314,N_43863);
xor U45932 (N_45932,N_43568,N_44804);
nand U45933 (N_45933,N_43496,N_43438);
xor U45934 (N_45934,N_42574,N_43281);
or U45935 (N_45935,N_43526,N_43458);
xnor U45936 (N_45936,N_44342,N_43242);
nor U45937 (N_45937,N_43197,N_44435);
or U45938 (N_45938,N_43678,N_44625);
nor U45939 (N_45939,N_43071,N_44914);
nand U45940 (N_45940,N_43934,N_42510);
or U45941 (N_45941,N_43531,N_42835);
and U45942 (N_45942,N_43910,N_43667);
nand U45943 (N_45943,N_44196,N_43525);
nand U45944 (N_45944,N_44950,N_43354);
or U45945 (N_45945,N_42648,N_43341);
or U45946 (N_45946,N_44089,N_44735);
and U45947 (N_45947,N_44411,N_44432);
and U45948 (N_45948,N_42823,N_44116);
nor U45949 (N_45949,N_43853,N_43683);
and U45950 (N_45950,N_44622,N_43209);
or U45951 (N_45951,N_43070,N_43840);
nand U45952 (N_45952,N_43768,N_44132);
and U45953 (N_45953,N_43296,N_42560);
or U45954 (N_45954,N_42649,N_44287);
or U45955 (N_45955,N_43347,N_42709);
and U45956 (N_45956,N_42859,N_43821);
nand U45957 (N_45957,N_44669,N_44233);
xnor U45958 (N_45958,N_42627,N_43916);
xor U45959 (N_45959,N_44254,N_42941);
nand U45960 (N_45960,N_43700,N_43990);
nor U45961 (N_45961,N_43501,N_42766);
and U45962 (N_45962,N_43642,N_44237);
nand U45963 (N_45963,N_44961,N_43573);
xor U45964 (N_45964,N_43080,N_44612);
nand U45965 (N_45965,N_42944,N_44910);
xnor U45966 (N_45966,N_44328,N_43564);
nor U45967 (N_45967,N_43245,N_44860);
nand U45968 (N_45968,N_44440,N_43641);
and U45969 (N_45969,N_43409,N_42754);
and U45970 (N_45970,N_43465,N_44037);
xor U45971 (N_45971,N_44811,N_44899);
nor U45972 (N_45972,N_44709,N_42714);
xnor U45973 (N_45973,N_44998,N_44475);
nor U45974 (N_45974,N_44297,N_43615);
and U45975 (N_45975,N_43299,N_44001);
nand U45976 (N_45976,N_44016,N_44945);
and U45977 (N_45977,N_44840,N_44498);
or U45978 (N_45978,N_43510,N_42808);
xnor U45979 (N_45979,N_43498,N_43378);
and U45980 (N_45980,N_43007,N_44343);
xnor U45981 (N_45981,N_43517,N_44716);
or U45982 (N_45982,N_44189,N_43796);
nor U45983 (N_45983,N_44085,N_43587);
nor U45984 (N_45984,N_44415,N_44869);
nor U45985 (N_45985,N_44494,N_44513);
xnor U45986 (N_45986,N_42646,N_44067);
nand U45987 (N_45987,N_44554,N_43376);
and U45988 (N_45988,N_43118,N_43006);
xor U45989 (N_45989,N_44410,N_42886);
nand U45990 (N_45990,N_43590,N_43388);
and U45991 (N_45991,N_44572,N_44393);
xnor U45992 (N_45992,N_44146,N_43603);
and U45993 (N_45993,N_43794,N_44497);
nor U45994 (N_45994,N_42645,N_44631);
and U45995 (N_45995,N_44245,N_43057);
xnor U45996 (N_45996,N_44707,N_44597);
nor U45997 (N_45997,N_42506,N_43899);
nand U45998 (N_45998,N_44667,N_42650);
and U45999 (N_45999,N_43753,N_43374);
nor U46000 (N_46000,N_43343,N_43895);
nor U46001 (N_46001,N_44978,N_44052);
nor U46002 (N_46002,N_44059,N_43908);
xnor U46003 (N_46003,N_43527,N_43002);
or U46004 (N_46004,N_44167,N_43104);
xor U46005 (N_46005,N_44710,N_42677);
and U46006 (N_46006,N_44060,N_43915);
xor U46007 (N_46007,N_44791,N_44969);
xor U46008 (N_46008,N_43267,N_43795);
nand U46009 (N_46009,N_43738,N_44926);
nand U46010 (N_46010,N_42795,N_44561);
nand U46011 (N_46011,N_43040,N_44197);
and U46012 (N_46012,N_42751,N_44458);
and U46013 (N_46013,N_42741,N_43105);
and U46014 (N_46014,N_43117,N_44813);
nand U46015 (N_46015,N_43014,N_43512);
and U46016 (N_46016,N_44973,N_42690);
xnor U46017 (N_46017,N_44445,N_43001);
xnor U46018 (N_46018,N_44421,N_43887);
nor U46019 (N_46019,N_44598,N_42854);
and U46020 (N_46020,N_43847,N_42985);
or U46021 (N_46021,N_44954,N_42828);
or U46022 (N_46022,N_44583,N_44782);
nor U46023 (N_46023,N_44467,N_44986);
and U46024 (N_46024,N_43902,N_42830);
nand U46025 (N_46025,N_44038,N_44807);
xnor U46026 (N_46026,N_42760,N_44495);
and U46027 (N_46027,N_43020,N_44774);
and U46028 (N_46028,N_44359,N_44831);
nand U46029 (N_46029,N_43398,N_43928);
xnor U46030 (N_46030,N_44346,N_42781);
xnor U46031 (N_46031,N_44356,N_44959);
and U46032 (N_46032,N_44088,N_43823);
xnor U46033 (N_46033,N_43544,N_43702);
and U46034 (N_46034,N_43718,N_44291);
and U46035 (N_46035,N_42527,N_43917);
nor U46036 (N_46036,N_44585,N_42564);
xnor U46037 (N_46037,N_44119,N_44317);
and U46038 (N_46038,N_43238,N_42512);
xnor U46039 (N_46039,N_44933,N_43455);
and U46040 (N_46040,N_43478,N_44690);
and U46041 (N_46041,N_43827,N_44799);
or U46042 (N_46042,N_42993,N_43375);
and U46043 (N_46043,N_44363,N_43972);
or U46044 (N_46044,N_43218,N_44867);
nand U46045 (N_46045,N_44580,N_44777);
xnor U46046 (N_46046,N_44176,N_43109);
or U46047 (N_46047,N_42822,N_42730);
nor U46048 (N_46048,N_42825,N_44740);
or U46049 (N_46049,N_43151,N_43798);
xor U46050 (N_46050,N_44662,N_44739);
nor U46051 (N_46051,N_44575,N_43086);
or U46052 (N_46052,N_44221,N_43308);
nand U46053 (N_46053,N_43716,N_43128);
xor U46054 (N_46054,N_44015,N_43741);
nor U46055 (N_46055,N_43536,N_44406);
and U46056 (N_46056,N_43144,N_43651);
nand U46057 (N_46057,N_44018,N_44438);
nor U46058 (N_46058,N_44558,N_44516);
xor U46059 (N_46059,N_44152,N_44091);
nand U46060 (N_46060,N_42657,N_43361);
xnor U46061 (N_46061,N_42775,N_44153);
or U46062 (N_46062,N_44552,N_44251);
xnor U46063 (N_46063,N_42844,N_44706);
xnor U46064 (N_46064,N_44390,N_43690);
or U46065 (N_46065,N_42971,N_42573);
xnor U46066 (N_46066,N_44855,N_43125);
nand U46067 (N_46067,N_43817,N_43248);
xnor U46068 (N_46068,N_42623,N_43537);
nor U46069 (N_46069,N_43288,N_42600);
or U46070 (N_46070,N_43930,N_44746);
xor U46071 (N_46071,N_44354,N_44772);
nor U46072 (N_46072,N_44618,N_43638);
nand U46073 (N_46073,N_44355,N_42962);
nand U46074 (N_46074,N_42638,N_42672);
and U46075 (N_46075,N_44854,N_43785);
nand U46076 (N_46076,N_43866,N_43709);
or U46077 (N_46077,N_43293,N_44201);
nor U46078 (N_46078,N_42529,N_43431);
and U46079 (N_46079,N_43997,N_43585);
xnor U46080 (N_46080,N_44876,N_43685);
nand U46081 (N_46081,N_43767,N_44040);
and U46082 (N_46082,N_44335,N_42546);
xnor U46083 (N_46083,N_42970,N_44358);
and U46084 (N_46084,N_44891,N_44485);
nor U46085 (N_46085,N_42673,N_44321);
xor U46086 (N_46086,N_43055,N_43470);
xnor U46087 (N_46087,N_43060,N_43790);
and U46088 (N_46088,N_44161,N_44262);
nor U46089 (N_46089,N_43613,N_43096);
xor U46090 (N_46090,N_43627,N_42763);
nand U46091 (N_46091,N_43921,N_42635);
nor U46092 (N_46092,N_43675,N_42934);
nor U46093 (N_46093,N_44369,N_43320);
nor U46094 (N_46094,N_43441,N_43329);
or U46095 (N_46095,N_42848,N_44405);
or U46096 (N_46096,N_43363,N_44770);
or U46097 (N_46097,N_44975,N_44937);
or U46098 (N_46098,N_42595,N_44300);
xnor U46099 (N_46099,N_44382,N_44253);
or U46100 (N_46100,N_44714,N_44785);
nand U46101 (N_46101,N_44381,N_43289);
nor U46102 (N_46102,N_44731,N_43734);
nand U46103 (N_46103,N_43581,N_42596);
nor U46104 (N_46104,N_42983,N_43228);
nor U46105 (N_46105,N_43131,N_43161);
xnor U46106 (N_46106,N_44086,N_44128);
xor U46107 (N_46107,N_42955,N_44212);
nor U46108 (N_46108,N_44550,N_43201);
or U46109 (N_46109,N_43516,N_44483);
nor U46110 (N_46110,N_43098,N_43112);
and U46111 (N_46111,N_43049,N_44542);
nand U46112 (N_46112,N_43170,N_44500);
or U46113 (N_46113,N_42591,N_42502);
nand U46114 (N_46114,N_44182,N_44477);
nor U46115 (N_46115,N_43815,N_43876);
or U46116 (N_46116,N_44075,N_43208);
nand U46117 (N_46117,N_43291,N_43194);
nor U46118 (N_46118,N_43841,N_44504);
nand U46119 (N_46119,N_44749,N_44919);
nor U46120 (N_46120,N_43975,N_44771);
nor U46121 (N_46121,N_44570,N_43298);
nor U46122 (N_46122,N_44121,N_43943);
or U46123 (N_46123,N_43922,N_44956);
and U46124 (N_46124,N_44484,N_43867);
xor U46125 (N_46125,N_43158,N_43845);
or U46126 (N_46126,N_44387,N_43167);
and U46127 (N_46127,N_42891,N_43113);
xor U46128 (N_46128,N_44447,N_42898);
nand U46129 (N_46129,N_42568,N_44007);
or U46130 (N_46130,N_44717,N_44270);
nand U46131 (N_46131,N_42931,N_42806);
nand U46132 (N_46132,N_42675,N_43110);
xor U46133 (N_46133,N_44564,N_43932);
and U46134 (N_46134,N_43724,N_42547);
and U46135 (N_46135,N_43557,N_44013);
nand U46136 (N_46136,N_43142,N_43674);
nor U46137 (N_46137,N_43206,N_42915);
and U46138 (N_46138,N_44195,N_44488);
nand U46139 (N_46139,N_43377,N_42850);
and U46140 (N_46140,N_42951,N_42578);
xor U46141 (N_46141,N_43502,N_44208);
nand U46142 (N_46142,N_44779,N_43108);
xor U46143 (N_46143,N_43483,N_42575);
or U46144 (N_46144,N_44338,N_42838);
and U46145 (N_46145,N_44880,N_42765);
or U46146 (N_46146,N_43858,N_43089);
and U46147 (N_46147,N_42706,N_44822);
or U46148 (N_46148,N_42584,N_43640);
nor U46149 (N_46149,N_42809,N_44847);
xnor U46150 (N_46150,N_43621,N_43825);
nor U46151 (N_46151,N_43423,N_44524);
or U46152 (N_46152,N_44470,N_44995);
xor U46153 (N_46153,N_44990,N_43826);
nor U46154 (N_46154,N_43427,N_43985);
and U46155 (N_46155,N_42804,N_43558);
and U46156 (N_46156,N_43865,N_44348);
nor U46157 (N_46157,N_44786,N_42713);
nand U46158 (N_46158,N_43048,N_43645);
and U46159 (N_46159,N_43992,N_43261);
or U46160 (N_46160,N_43514,N_43492);
and U46161 (N_46161,N_44634,N_44165);
nor U46162 (N_46162,N_44697,N_42913);
or U46163 (N_46163,N_42942,N_44240);
nor U46164 (N_46164,N_44944,N_42796);
nor U46165 (N_46165,N_44982,N_44127);
and U46166 (N_46166,N_42748,N_44172);
xor U46167 (N_46167,N_44199,N_42869);
nand U46168 (N_46168,N_43945,N_42860);
nand U46169 (N_46169,N_43861,N_44871);
or U46170 (N_46170,N_42619,N_44681);
xor U46171 (N_46171,N_44548,N_43448);
nand U46172 (N_46172,N_42610,N_43051);
nor U46173 (N_46173,N_43509,N_43949);
nor U46174 (N_46174,N_43695,N_43268);
xor U46175 (N_46175,N_43141,N_43087);
xor U46176 (N_46176,N_44290,N_43938);
and U46177 (N_46177,N_42633,N_43920);
and U46178 (N_46178,N_44605,N_43862);
nor U46179 (N_46179,N_44768,N_44336);
xnor U46180 (N_46180,N_43420,N_43944);
nand U46181 (N_46181,N_44611,N_42562);
nand U46182 (N_46182,N_43802,N_42987);
or U46183 (N_46183,N_44257,N_42515);
nor U46184 (N_46184,N_43036,N_44930);
nand U46185 (N_46185,N_44402,N_42920);
xnor U46186 (N_46186,N_43846,N_44842);
or U46187 (N_46187,N_43385,N_44283);
xnor U46188 (N_46188,N_44163,N_43432);
xnor U46189 (N_46189,N_43728,N_43157);
nand U46190 (N_46190,N_44191,N_43658);
xor U46191 (N_46191,N_42773,N_43391);
nor U46192 (N_46192,N_44261,N_42947);
or U46193 (N_46193,N_42726,N_43159);
or U46194 (N_46194,N_43605,N_44236);
xnor U46195 (N_46195,N_42608,N_44646);
nand U46196 (N_46196,N_44723,N_43072);
nor U46197 (N_46197,N_43165,N_43889);
xor U46198 (N_46198,N_43781,N_43676);
nor U46199 (N_46199,N_43708,N_44968);
nor U46200 (N_46200,N_42644,N_43490);
and U46201 (N_46201,N_44981,N_43482);
nand U46202 (N_46202,N_43807,N_44825);
nand U46203 (N_46203,N_43284,N_43457);
or U46204 (N_46204,N_43148,N_42678);
and U46205 (N_46205,N_42887,N_42953);
and U46206 (N_46206,N_43115,N_44468);
and U46207 (N_46207,N_43731,N_44757);
xor U46208 (N_46208,N_43068,N_44536);
and U46209 (N_46209,N_43697,N_44499);
and U46210 (N_46210,N_42558,N_43307);
and U46211 (N_46211,N_44759,N_43166);
xor U46212 (N_46212,N_43102,N_42671);
xor U46213 (N_46213,N_44098,N_44531);
nand U46214 (N_46214,N_43137,N_44501);
nor U46215 (N_46215,N_42932,N_44454);
xnor U46216 (N_46216,N_42874,N_42513);
and U46217 (N_46217,N_43933,N_42625);
and U46218 (N_46218,N_43467,N_44048);
nor U46219 (N_46219,N_42939,N_44792);
nand U46220 (N_46220,N_43878,N_43913);
nand U46221 (N_46221,N_43241,N_44935);
and U46222 (N_46222,N_43748,N_43269);
and U46223 (N_46223,N_43193,N_43736);
xor U46224 (N_46224,N_42791,N_44528);
nor U46225 (N_46225,N_43011,N_42752);
nor U46226 (N_46226,N_42629,N_43019);
and U46227 (N_46227,N_43216,N_44223);
or U46228 (N_46228,N_44644,N_44836);
xnor U46229 (N_46229,N_43880,N_43145);
xnor U46230 (N_46230,N_43635,N_42658);
or U46231 (N_46231,N_44627,N_43367);
nor U46232 (N_46232,N_43799,N_44698);
xnor U46233 (N_46233,N_44729,N_43844);
and U46234 (N_46234,N_44149,N_44327);
or U46235 (N_46235,N_44783,N_43017);
xnor U46236 (N_46236,N_42668,N_43217);
or U46237 (N_46237,N_43711,N_43283);
and U46238 (N_46238,N_43013,N_43274);
and U46239 (N_46239,N_44509,N_42613);
xnor U46240 (N_46240,N_44183,N_44579);
and U46241 (N_46241,N_43719,N_44905);
xor U46242 (N_46242,N_43480,N_42757);
or U46243 (N_46243,N_43380,N_43485);
or U46244 (N_46244,N_44879,N_44209);
or U46245 (N_46245,N_44949,N_44168);
and U46246 (N_46246,N_43130,N_42695);
nand U46247 (N_46247,N_43326,N_43163);
nand U46248 (N_46248,N_42716,N_43958);
and U46249 (N_46249,N_43650,N_44629);
nand U46250 (N_46250,N_44514,N_43229);
nor U46251 (N_46251,N_43373,N_42900);
nand U46252 (N_46252,N_44747,N_43861);
or U46253 (N_46253,N_42760,N_42949);
or U46254 (N_46254,N_44436,N_42833);
and U46255 (N_46255,N_44831,N_44113);
and U46256 (N_46256,N_44766,N_43658);
and U46257 (N_46257,N_42669,N_44142);
nand U46258 (N_46258,N_44514,N_42723);
xnor U46259 (N_46259,N_42656,N_43210);
xnor U46260 (N_46260,N_42645,N_44197);
xor U46261 (N_46261,N_44201,N_44547);
nor U46262 (N_46262,N_43102,N_44200);
or U46263 (N_46263,N_43215,N_44170);
or U46264 (N_46264,N_43570,N_44838);
or U46265 (N_46265,N_44214,N_43051);
xnor U46266 (N_46266,N_42904,N_43493);
xnor U46267 (N_46267,N_43282,N_44874);
xor U46268 (N_46268,N_42872,N_44356);
and U46269 (N_46269,N_42916,N_44181);
xnor U46270 (N_46270,N_43511,N_44305);
nor U46271 (N_46271,N_42659,N_44329);
xor U46272 (N_46272,N_44382,N_43371);
xnor U46273 (N_46273,N_43870,N_42600);
nand U46274 (N_46274,N_43070,N_42804);
or U46275 (N_46275,N_43569,N_44171);
and U46276 (N_46276,N_42921,N_44879);
nand U46277 (N_46277,N_44973,N_42976);
xor U46278 (N_46278,N_44409,N_43193);
nor U46279 (N_46279,N_44372,N_44338);
xnor U46280 (N_46280,N_43967,N_42914);
or U46281 (N_46281,N_43685,N_42734);
and U46282 (N_46282,N_44484,N_44981);
nand U46283 (N_46283,N_43010,N_44405);
nor U46284 (N_46284,N_44337,N_43851);
nor U46285 (N_46285,N_43583,N_44509);
nor U46286 (N_46286,N_42672,N_44280);
nand U46287 (N_46287,N_44772,N_44095);
nor U46288 (N_46288,N_44388,N_43877);
and U46289 (N_46289,N_42625,N_42753);
xnor U46290 (N_46290,N_44432,N_43502);
and U46291 (N_46291,N_44744,N_42958);
xnor U46292 (N_46292,N_44713,N_44729);
xor U46293 (N_46293,N_44095,N_42814);
or U46294 (N_46294,N_42859,N_44504);
nand U46295 (N_46295,N_43979,N_44349);
xnor U46296 (N_46296,N_44568,N_43956);
xor U46297 (N_46297,N_44274,N_43503);
nand U46298 (N_46298,N_42555,N_44611);
nor U46299 (N_46299,N_42780,N_44541);
xnor U46300 (N_46300,N_43524,N_44035);
nor U46301 (N_46301,N_44654,N_44673);
or U46302 (N_46302,N_43614,N_43761);
and U46303 (N_46303,N_44004,N_44520);
nor U46304 (N_46304,N_44925,N_43758);
nor U46305 (N_46305,N_44779,N_44419);
nor U46306 (N_46306,N_44493,N_44964);
and U46307 (N_46307,N_44472,N_43003);
nand U46308 (N_46308,N_43351,N_43583);
nor U46309 (N_46309,N_43795,N_44118);
or U46310 (N_46310,N_44741,N_43325);
xnor U46311 (N_46311,N_43478,N_44960);
and U46312 (N_46312,N_44548,N_44100);
xnor U46313 (N_46313,N_42553,N_42719);
nor U46314 (N_46314,N_43378,N_44684);
and U46315 (N_46315,N_43419,N_43784);
and U46316 (N_46316,N_43734,N_44698);
nand U46317 (N_46317,N_43204,N_42697);
xor U46318 (N_46318,N_44258,N_42778);
nor U46319 (N_46319,N_44025,N_44200);
or U46320 (N_46320,N_43874,N_43127);
or U46321 (N_46321,N_43009,N_43602);
nor U46322 (N_46322,N_44984,N_44746);
or U46323 (N_46323,N_43021,N_42869);
and U46324 (N_46324,N_43081,N_42917);
or U46325 (N_46325,N_44267,N_44628);
nor U46326 (N_46326,N_44418,N_43752);
nand U46327 (N_46327,N_44054,N_43743);
or U46328 (N_46328,N_42680,N_42930);
nand U46329 (N_46329,N_44372,N_43703);
and U46330 (N_46330,N_44249,N_43257);
and U46331 (N_46331,N_42895,N_42751);
xor U46332 (N_46332,N_44703,N_43041);
and U46333 (N_46333,N_44354,N_44272);
and U46334 (N_46334,N_43466,N_43841);
nand U46335 (N_46335,N_44590,N_43887);
xor U46336 (N_46336,N_43416,N_43597);
nand U46337 (N_46337,N_42890,N_43834);
xnor U46338 (N_46338,N_44003,N_43021);
xor U46339 (N_46339,N_44589,N_44997);
and U46340 (N_46340,N_43610,N_43614);
xnor U46341 (N_46341,N_43388,N_42752);
nand U46342 (N_46342,N_42941,N_42550);
or U46343 (N_46343,N_43427,N_44861);
or U46344 (N_46344,N_42967,N_43387);
nand U46345 (N_46345,N_42696,N_44585);
nand U46346 (N_46346,N_44406,N_44340);
nand U46347 (N_46347,N_42681,N_42856);
or U46348 (N_46348,N_43268,N_44054);
xnor U46349 (N_46349,N_43758,N_43258);
or U46350 (N_46350,N_44036,N_43872);
and U46351 (N_46351,N_42869,N_44095);
nand U46352 (N_46352,N_43004,N_44772);
nand U46353 (N_46353,N_44239,N_42785);
xor U46354 (N_46354,N_43982,N_43962);
nand U46355 (N_46355,N_42565,N_43093);
and U46356 (N_46356,N_43643,N_43371);
xnor U46357 (N_46357,N_43455,N_43506);
nor U46358 (N_46358,N_44208,N_42663);
nand U46359 (N_46359,N_44010,N_42837);
xnor U46360 (N_46360,N_44985,N_44770);
xor U46361 (N_46361,N_42925,N_44656);
nand U46362 (N_46362,N_44799,N_43124);
or U46363 (N_46363,N_43561,N_44880);
or U46364 (N_46364,N_43288,N_44203);
nor U46365 (N_46365,N_43515,N_44146);
and U46366 (N_46366,N_44788,N_43496);
or U46367 (N_46367,N_43295,N_43450);
and U46368 (N_46368,N_44453,N_44909);
nor U46369 (N_46369,N_43268,N_43816);
xnor U46370 (N_46370,N_43717,N_42945);
and U46371 (N_46371,N_43972,N_43261);
and U46372 (N_46372,N_43643,N_43149);
nand U46373 (N_46373,N_42616,N_42907);
or U46374 (N_46374,N_43939,N_43262);
nand U46375 (N_46375,N_44078,N_43792);
nand U46376 (N_46376,N_43212,N_44359);
or U46377 (N_46377,N_44746,N_42913);
nor U46378 (N_46378,N_43458,N_42632);
xnor U46379 (N_46379,N_44962,N_44415);
nor U46380 (N_46380,N_43817,N_43143);
and U46381 (N_46381,N_44976,N_44100);
and U46382 (N_46382,N_44082,N_44144);
nor U46383 (N_46383,N_44635,N_44098);
and U46384 (N_46384,N_44323,N_42879);
xnor U46385 (N_46385,N_43298,N_44291);
or U46386 (N_46386,N_43128,N_43149);
xnor U46387 (N_46387,N_44245,N_44910);
nor U46388 (N_46388,N_42711,N_44943);
nand U46389 (N_46389,N_42945,N_43416);
or U46390 (N_46390,N_44272,N_42748);
nand U46391 (N_46391,N_43898,N_43670);
nand U46392 (N_46392,N_43297,N_42766);
and U46393 (N_46393,N_44633,N_43298);
and U46394 (N_46394,N_42757,N_44725);
nor U46395 (N_46395,N_43108,N_44206);
and U46396 (N_46396,N_44606,N_43060);
nand U46397 (N_46397,N_44605,N_43606);
or U46398 (N_46398,N_42768,N_44054);
or U46399 (N_46399,N_44755,N_44642);
nand U46400 (N_46400,N_43521,N_43173);
nor U46401 (N_46401,N_43494,N_44837);
or U46402 (N_46402,N_44152,N_42842);
nor U46403 (N_46403,N_44574,N_43086);
nor U46404 (N_46404,N_43997,N_43671);
and U46405 (N_46405,N_44265,N_44412);
nor U46406 (N_46406,N_43290,N_42540);
or U46407 (N_46407,N_44277,N_42917);
nor U46408 (N_46408,N_44015,N_43017);
or U46409 (N_46409,N_42760,N_44072);
and U46410 (N_46410,N_43760,N_43172);
and U46411 (N_46411,N_44916,N_44363);
nand U46412 (N_46412,N_42613,N_44272);
or U46413 (N_46413,N_44641,N_44683);
nor U46414 (N_46414,N_44673,N_42512);
and U46415 (N_46415,N_43748,N_42639);
nand U46416 (N_46416,N_44586,N_42693);
and U46417 (N_46417,N_43155,N_44164);
nand U46418 (N_46418,N_44148,N_42745);
nor U46419 (N_46419,N_44282,N_43745);
nor U46420 (N_46420,N_42967,N_44081);
nand U46421 (N_46421,N_43973,N_44817);
and U46422 (N_46422,N_44372,N_43897);
nand U46423 (N_46423,N_44524,N_43055);
and U46424 (N_46424,N_42616,N_43602);
xor U46425 (N_46425,N_43633,N_44529);
and U46426 (N_46426,N_43339,N_44119);
or U46427 (N_46427,N_43598,N_44649);
nor U46428 (N_46428,N_43844,N_43358);
and U46429 (N_46429,N_43965,N_44116);
or U46430 (N_46430,N_42663,N_43240);
xor U46431 (N_46431,N_44627,N_44670);
and U46432 (N_46432,N_43185,N_44686);
nand U46433 (N_46433,N_44377,N_43609);
xor U46434 (N_46434,N_44726,N_43771);
and U46435 (N_46435,N_42581,N_44298);
or U46436 (N_46436,N_43554,N_44251);
xnor U46437 (N_46437,N_42950,N_44014);
or U46438 (N_46438,N_44585,N_44529);
nor U46439 (N_46439,N_43321,N_44414);
xor U46440 (N_46440,N_43471,N_44473);
nor U46441 (N_46441,N_43467,N_43660);
nor U46442 (N_46442,N_44341,N_43590);
or U46443 (N_46443,N_43048,N_44280);
xnor U46444 (N_46444,N_44966,N_43226);
or U46445 (N_46445,N_42769,N_43743);
nand U46446 (N_46446,N_43729,N_42585);
nand U46447 (N_46447,N_44743,N_44864);
or U46448 (N_46448,N_44101,N_44545);
nand U46449 (N_46449,N_42917,N_43943);
or U46450 (N_46450,N_43406,N_42648);
nand U46451 (N_46451,N_43326,N_43432);
nand U46452 (N_46452,N_44612,N_43456);
xor U46453 (N_46453,N_44056,N_43407);
or U46454 (N_46454,N_42922,N_44975);
and U46455 (N_46455,N_42761,N_43862);
nand U46456 (N_46456,N_44563,N_43231);
and U46457 (N_46457,N_42645,N_44005);
nor U46458 (N_46458,N_43055,N_44166);
nand U46459 (N_46459,N_42824,N_43880);
or U46460 (N_46460,N_42599,N_43041);
nor U46461 (N_46461,N_43210,N_43171);
or U46462 (N_46462,N_44843,N_44136);
and U46463 (N_46463,N_43023,N_44437);
xor U46464 (N_46464,N_44957,N_43259);
and U46465 (N_46465,N_43654,N_44737);
xor U46466 (N_46466,N_44922,N_43822);
and U46467 (N_46467,N_44048,N_43101);
and U46468 (N_46468,N_44728,N_43560);
or U46469 (N_46469,N_43844,N_44122);
nor U46470 (N_46470,N_44739,N_43059);
xnor U46471 (N_46471,N_42792,N_44018);
or U46472 (N_46472,N_43750,N_43528);
nand U46473 (N_46473,N_44804,N_43208);
nand U46474 (N_46474,N_44422,N_43529);
and U46475 (N_46475,N_43901,N_44327);
xor U46476 (N_46476,N_44410,N_44885);
nand U46477 (N_46477,N_44595,N_44866);
nand U46478 (N_46478,N_44409,N_42771);
or U46479 (N_46479,N_42512,N_42693);
or U46480 (N_46480,N_42636,N_43027);
or U46481 (N_46481,N_44549,N_44813);
or U46482 (N_46482,N_44310,N_44588);
nor U46483 (N_46483,N_42675,N_44159);
and U46484 (N_46484,N_43566,N_43321);
or U46485 (N_46485,N_44492,N_44152);
nand U46486 (N_46486,N_44626,N_43424);
xnor U46487 (N_46487,N_43429,N_42534);
or U46488 (N_46488,N_43250,N_42777);
xor U46489 (N_46489,N_43675,N_44596);
or U46490 (N_46490,N_44680,N_42743);
nand U46491 (N_46491,N_43126,N_44560);
or U46492 (N_46492,N_44708,N_44262);
nand U46493 (N_46493,N_44435,N_43541);
xnor U46494 (N_46494,N_44419,N_43761);
nor U46495 (N_46495,N_43233,N_43690);
nor U46496 (N_46496,N_44324,N_44913);
xnor U46497 (N_46497,N_43510,N_44918);
nand U46498 (N_46498,N_43746,N_43710);
xnor U46499 (N_46499,N_43863,N_43710);
or U46500 (N_46500,N_44496,N_43453);
nand U46501 (N_46501,N_44828,N_43832);
nor U46502 (N_46502,N_44144,N_44719);
xnor U46503 (N_46503,N_44650,N_42814);
nor U46504 (N_46504,N_43621,N_43550);
nand U46505 (N_46505,N_44444,N_43097);
xnor U46506 (N_46506,N_44924,N_43364);
xnor U46507 (N_46507,N_44053,N_43294);
and U46508 (N_46508,N_43813,N_42655);
and U46509 (N_46509,N_43795,N_44602);
or U46510 (N_46510,N_42910,N_43010);
xor U46511 (N_46511,N_43746,N_43080);
xnor U46512 (N_46512,N_44196,N_43753);
and U46513 (N_46513,N_44849,N_44905);
and U46514 (N_46514,N_43839,N_43352);
xor U46515 (N_46515,N_42893,N_42519);
or U46516 (N_46516,N_42524,N_43045);
nand U46517 (N_46517,N_44801,N_43606);
and U46518 (N_46518,N_42962,N_44611);
and U46519 (N_46519,N_44050,N_43357);
xor U46520 (N_46520,N_42621,N_42636);
xnor U46521 (N_46521,N_44863,N_43554);
and U46522 (N_46522,N_43531,N_44501);
xor U46523 (N_46523,N_44084,N_43885);
nor U46524 (N_46524,N_43300,N_44491);
and U46525 (N_46525,N_42635,N_42994);
xnor U46526 (N_46526,N_43183,N_43263);
or U46527 (N_46527,N_44058,N_44797);
nor U46528 (N_46528,N_43126,N_44841);
and U46529 (N_46529,N_44381,N_44858);
or U46530 (N_46530,N_42814,N_44720);
or U46531 (N_46531,N_43631,N_42786);
or U46532 (N_46532,N_43151,N_44808);
nor U46533 (N_46533,N_43050,N_44520);
and U46534 (N_46534,N_43641,N_42915);
and U46535 (N_46535,N_42794,N_44817);
xnor U46536 (N_46536,N_44597,N_42509);
nor U46537 (N_46537,N_44316,N_43091);
nand U46538 (N_46538,N_44339,N_44047);
and U46539 (N_46539,N_44761,N_42722);
xnor U46540 (N_46540,N_43345,N_43269);
xnor U46541 (N_46541,N_44584,N_42676);
nand U46542 (N_46542,N_44179,N_42601);
and U46543 (N_46543,N_42971,N_44923);
or U46544 (N_46544,N_42755,N_44103);
nor U46545 (N_46545,N_43390,N_43167);
nand U46546 (N_46546,N_42623,N_44013);
xnor U46547 (N_46547,N_43514,N_43923);
xor U46548 (N_46548,N_44041,N_43562);
nor U46549 (N_46549,N_44820,N_44243);
and U46550 (N_46550,N_43211,N_42544);
and U46551 (N_46551,N_43301,N_43741);
nor U46552 (N_46552,N_44308,N_42994);
xnor U46553 (N_46553,N_44611,N_43145);
or U46554 (N_46554,N_43791,N_43228);
nor U46555 (N_46555,N_43618,N_42815);
nand U46556 (N_46556,N_43682,N_44565);
nor U46557 (N_46557,N_43363,N_43915);
xor U46558 (N_46558,N_44711,N_44775);
nor U46559 (N_46559,N_44430,N_42500);
and U46560 (N_46560,N_43621,N_43334);
xor U46561 (N_46561,N_42639,N_43223);
nand U46562 (N_46562,N_43040,N_43516);
and U46563 (N_46563,N_43559,N_44038);
or U46564 (N_46564,N_44666,N_44482);
and U46565 (N_46565,N_43200,N_44531);
or U46566 (N_46566,N_44428,N_44062);
nor U46567 (N_46567,N_43198,N_43819);
xor U46568 (N_46568,N_43555,N_44031);
and U46569 (N_46569,N_44004,N_42997);
and U46570 (N_46570,N_44254,N_42750);
nor U46571 (N_46571,N_44014,N_44827);
nand U46572 (N_46572,N_43448,N_43397);
nor U46573 (N_46573,N_44644,N_42788);
or U46574 (N_46574,N_43239,N_42896);
xor U46575 (N_46575,N_43549,N_42602);
and U46576 (N_46576,N_42628,N_43974);
nor U46577 (N_46577,N_43306,N_43341);
and U46578 (N_46578,N_44541,N_44062);
or U46579 (N_46579,N_44440,N_44822);
nand U46580 (N_46580,N_44204,N_43318);
nor U46581 (N_46581,N_42837,N_44474);
nand U46582 (N_46582,N_44494,N_43533);
and U46583 (N_46583,N_44505,N_43987);
or U46584 (N_46584,N_43126,N_43152);
nor U46585 (N_46585,N_43516,N_43122);
xor U46586 (N_46586,N_44694,N_42895);
nor U46587 (N_46587,N_43096,N_44739);
nor U46588 (N_46588,N_44533,N_44220);
or U46589 (N_46589,N_44080,N_42812);
nand U46590 (N_46590,N_44815,N_43682);
and U46591 (N_46591,N_44182,N_44816);
xnor U46592 (N_46592,N_44784,N_42823);
or U46593 (N_46593,N_44796,N_44168);
xor U46594 (N_46594,N_42878,N_43529);
nor U46595 (N_46595,N_43546,N_44661);
nand U46596 (N_46596,N_42949,N_43678);
or U46597 (N_46597,N_42616,N_43820);
nand U46598 (N_46598,N_44070,N_42822);
nor U46599 (N_46599,N_43093,N_43095);
or U46600 (N_46600,N_43584,N_43443);
nand U46601 (N_46601,N_44905,N_43255);
nand U46602 (N_46602,N_42606,N_43038);
nor U46603 (N_46603,N_43432,N_43903);
xnor U46604 (N_46604,N_44659,N_42662);
nand U46605 (N_46605,N_42519,N_44637);
nor U46606 (N_46606,N_42651,N_44533);
nor U46607 (N_46607,N_43024,N_43383);
nor U46608 (N_46608,N_42522,N_44382);
nor U46609 (N_46609,N_44288,N_43633);
and U46610 (N_46610,N_42995,N_44606);
nand U46611 (N_46611,N_42665,N_42712);
and U46612 (N_46612,N_43217,N_44743);
and U46613 (N_46613,N_44807,N_42810);
or U46614 (N_46614,N_42670,N_43431);
xor U46615 (N_46615,N_44322,N_43660);
xnor U46616 (N_46616,N_42508,N_44799);
nor U46617 (N_46617,N_43383,N_44972);
and U46618 (N_46618,N_42889,N_42520);
nand U46619 (N_46619,N_44539,N_43179);
nand U46620 (N_46620,N_43433,N_43767);
nand U46621 (N_46621,N_43590,N_43533);
nand U46622 (N_46622,N_42865,N_42738);
xor U46623 (N_46623,N_44148,N_43857);
or U46624 (N_46624,N_44924,N_42622);
and U46625 (N_46625,N_44597,N_43745);
xor U46626 (N_46626,N_43541,N_43595);
nor U46627 (N_46627,N_44295,N_44977);
and U46628 (N_46628,N_44715,N_43240);
or U46629 (N_46629,N_44316,N_44566);
nand U46630 (N_46630,N_43382,N_44313);
nand U46631 (N_46631,N_44868,N_44764);
or U46632 (N_46632,N_43343,N_43845);
xnor U46633 (N_46633,N_43242,N_43012);
or U46634 (N_46634,N_43659,N_43888);
nand U46635 (N_46635,N_42518,N_44318);
nand U46636 (N_46636,N_43064,N_43937);
or U46637 (N_46637,N_43850,N_42894);
nand U46638 (N_46638,N_43563,N_44169);
and U46639 (N_46639,N_43320,N_42835);
or U46640 (N_46640,N_44930,N_44269);
nand U46641 (N_46641,N_43121,N_43281);
nand U46642 (N_46642,N_42756,N_44258);
and U46643 (N_46643,N_44148,N_43932);
nor U46644 (N_46644,N_43802,N_44565);
xnor U46645 (N_46645,N_44537,N_42591);
nor U46646 (N_46646,N_43033,N_44017);
and U46647 (N_46647,N_44571,N_44088);
xnor U46648 (N_46648,N_44867,N_44862);
xnor U46649 (N_46649,N_43953,N_43267);
xnor U46650 (N_46650,N_43624,N_43519);
nor U46651 (N_46651,N_44643,N_44338);
xor U46652 (N_46652,N_42729,N_43445);
nand U46653 (N_46653,N_44945,N_43233);
and U46654 (N_46654,N_44101,N_44754);
xnor U46655 (N_46655,N_44339,N_44648);
xor U46656 (N_46656,N_44170,N_44968);
nor U46657 (N_46657,N_44685,N_44675);
and U46658 (N_46658,N_43740,N_42799);
nor U46659 (N_46659,N_43401,N_44661);
xor U46660 (N_46660,N_44428,N_44212);
or U46661 (N_46661,N_43061,N_42892);
or U46662 (N_46662,N_42538,N_43587);
xor U46663 (N_46663,N_43185,N_44029);
xnor U46664 (N_46664,N_43883,N_42691);
nor U46665 (N_46665,N_44488,N_43913);
nand U46666 (N_46666,N_43631,N_43561);
and U46667 (N_46667,N_43824,N_43739);
and U46668 (N_46668,N_44155,N_43374);
xnor U46669 (N_46669,N_44401,N_43773);
xnor U46670 (N_46670,N_44304,N_42639);
xnor U46671 (N_46671,N_42527,N_43629);
nand U46672 (N_46672,N_43281,N_44688);
or U46673 (N_46673,N_42971,N_42697);
xnor U46674 (N_46674,N_44831,N_42969);
nor U46675 (N_46675,N_43369,N_43496);
and U46676 (N_46676,N_44472,N_43259);
or U46677 (N_46677,N_44279,N_42842);
xnor U46678 (N_46678,N_43732,N_44943);
and U46679 (N_46679,N_43431,N_44226);
nand U46680 (N_46680,N_43119,N_43175);
nor U46681 (N_46681,N_43391,N_42642);
xnor U46682 (N_46682,N_43851,N_43232);
nand U46683 (N_46683,N_44541,N_42971);
and U46684 (N_46684,N_44708,N_44450);
nor U46685 (N_46685,N_42646,N_43980);
or U46686 (N_46686,N_43410,N_44730);
or U46687 (N_46687,N_42852,N_44362);
and U46688 (N_46688,N_44419,N_44224);
nor U46689 (N_46689,N_42639,N_43903);
xnor U46690 (N_46690,N_43029,N_42908);
and U46691 (N_46691,N_44136,N_43486);
or U46692 (N_46692,N_43416,N_43995);
or U46693 (N_46693,N_44075,N_44047);
and U46694 (N_46694,N_44496,N_43973);
nor U46695 (N_46695,N_44436,N_44554);
and U46696 (N_46696,N_44058,N_43955);
nor U46697 (N_46697,N_44494,N_42539);
xnor U46698 (N_46698,N_43491,N_43792);
xnor U46699 (N_46699,N_43934,N_44936);
nand U46700 (N_46700,N_43138,N_43373);
xor U46701 (N_46701,N_44703,N_43577);
nand U46702 (N_46702,N_44428,N_44807);
or U46703 (N_46703,N_44003,N_44020);
nand U46704 (N_46704,N_43191,N_42802);
or U46705 (N_46705,N_43006,N_43839);
and U46706 (N_46706,N_43306,N_43143);
and U46707 (N_46707,N_44049,N_44713);
nand U46708 (N_46708,N_44293,N_44522);
or U46709 (N_46709,N_43501,N_42969);
nor U46710 (N_46710,N_43777,N_44815);
or U46711 (N_46711,N_42635,N_43496);
or U46712 (N_46712,N_44491,N_43087);
nand U46713 (N_46713,N_43036,N_44695);
nand U46714 (N_46714,N_42820,N_42635);
xor U46715 (N_46715,N_43501,N_42981);
and U46716 (N_46716,N_43660,N_44444);
or U46717 (N_46717,N_44263,N_44344);
nor U46718 (N_46718,N_43279,N_43505);
nand U46719 (N_46719,N_43453,N_43137);
xnor U46720 (N_46720,N_42785,N_43327);
and U46721 (N_46721,N_43911,N_44849);
or U46722 (N_46722,N_42560,N_43488);
xnor U46723 (N_46723,N_44274,N_42684);
nand U46724 (N_46724,N_43699,N_44847);
and U46725 (N_46725,N_44930,N_43674);
and U46726 (N_46726,N_44296,N_44039);
xnor U46727 (N_46727,N_43037,N_44375);
or U46728 (N_46728,N_44802,N_43807);
xnor U46729 (N_46729,N_43744,N_43224);
or U46730 (N_46730,N_43141,N_44178);
nor U46731 (N_46731,N_43095,N_43868);
xor U46732 (N_46732,N_44926,N_44839);
nand U46733 (N_46733,N_43322,N_44247);
and U46734 (N_46734,N_44227,N_43619);
nor U46735 (N_46735,N_43094,N_44011);
xnor U46736 (N_46736,N_44685,N_43963);
nand U46737 (N_46737,N_43482,N_43563);
or U46738 (N_46738,N_44790,N_43528);
nor U46739 (N_46739,N_43171,N_44704);
and U46740 (N_46740,N_43164,N_42521);
nand U46741 (N_46741,N_43607,N_44896);
nand U46742 (N_46742,N_44228,N_44878);
nand U46743 (N_46743,N_42583,N_44691);
nor U46744 (N_46744,N_43611,N_44958);
and U46745 (N_46745,N_43720,N_43833);
nor U46746 (N_46746,N_43078,N_43067);
and U46747 (N_46747,N_42924,N_44405);
nand U46748 (N_46748,N_43102,N_43932);
and U46749 (N_46749,N_43260,N_42564);
nand U46750 (N_46750,N_44590,N_43272);
xor U46751 (N_46751,N_43923,N_42550);
or U46752 (N_46752,N_43455,N_44662);
xnor U46753 (N_46753,N_44802,N_44724);
nand U46754 (N_46754,N_44634,N_43777);
xor U46755 (N_46755,N_44629,N_44354);
nand U46756 (N_46756,N_43038,N_43391);
xnor U46757 (N_46757,N_44109,N_43518);
xnor U46758 (N_46758,N_44718,N_44930);
nand U46759 (N_46759,N_43895,N_44317);
or U46760 (N_46760,N_44916,N_44036);
nor U46761 (N_46761,N_43542,N_42953);
or U46762 (N_46762,N_44180,N_42592);
and U46763 (N_46763,N_42668,N_43294);
nor U46764 (N_46764,N_44550,N_44581);
and U46765 (N_46765,N_44224,N_44241);
nand U46766 (N_46766,N_42894,N_43728);
nor U46767 (N_46767,N_42533,N_42786);
xor U46768 (N_46768,N_43562,N_42512);
nor U46769 (N_46769,N_42775,N_43433);
or U46770 (N_46770,N_42586,N_42858);
nor U46771 (N_46771,N_44552,N_44077);
or U46772 (N_46772,N_42591,N_43771);
nand U46773 (N_46773,N_44609,N_42653);
or U46774 (N_46774,N_44044,N_42812);
xor U46775 (N_46775,N_44778,N_44874);
nand U46776 (N_46776,N_43221,N_42656);
xnor U46777 (N_46777,N_42903,N_44005);
or U46778 (N_46778,N_43673,N_44872);
xnor U46779 (N_46779,N_44171,N_44126);
nor U46780 (N_46780,N_43721,N_42762);
or U46781 (N_46781,N_43252,N_43837);
or U46782 (N_46782,N_42559,N_44488);
nor U46783 (N_46783,N_42991,N_43009);
or U46784 (N_46784,N_43841,N_42930);
nand U46785 (N_46785,N_43814,N_42928);
nand U46786 (N_46786,N_42554,N_43404);
nor U46787 (N_46787,N_44226,N_42776);
nand U46788 (N_46788,N_44414,N_43509);
nor U46789 (N_46789,N_44911,N_44999);
and U46790 (N_46790,N_44829,N_43270);
and U46791 (N_46791,N_44004,N_42614);
and U46792 (N_46792,N_43164,N_43959);
and U46793 (N_46793,N_44650,N_44052);
nand U46794 (N_46794,N_42898,N_44285);
or U46795 (N_46795,N_44728,N_43441);
and U46796 (N_46796,N_43561,N_43770);
nand U46797 (N_46797,N_42526,N_44837);
xnor U46798 (N_46798,N_43227,N_43305);
nor U46799 (N_46799,N_42649,N_44272);
nor U46800 (N_46800,N_43214,N_44814);
nor U46801 (N_46801,N_42516,N_43198);
nand U46802 (N_46802,N_44434,N_44759);
and U46803 (N_46803,N_44626,N_42909);
or U46804 (N_46804,N_44393,N_43596);
xnor U46805 (N_46805,N_44007,N_42504);
or U46806 (N_46806,N_44182,N_44582);
or U46807 (N_46807,N_42770,N_44924);
or U46808 (N_46808,N_44157,N_43922);
xnor U46809 (N_46809,N_43159,N_44459);
and U46810 (N_46810,N_44348,N_43728);
nor U46811 (N_46811,N_44290,N_44679);
xnor U46812 (N_46812,N_42902,N_44066);
nand U46813 (N_46813,N_44108,N_44407);
and U46814 (N_46814,N_44049,N_42534);
xnor U46815 (N_46815,N_44297,N_43238);
xor U46816 (N_46816,N_44776,N_43487);
xor U46817 (N_46817,N_44317,N_43306);
xor U46818 (N_46818,N_44238,N_43605);
and U46819 (N_46819,N_44017,N_44125);
nor U46820 (N_46820,N_44693,N_44973);
xor U46821 (N_46821,N_43342,N_44718);
xnor U46822 (N_46822,N_44728,N_44287);
nand U46823 (N_46823,N_42793,N_44335);
xor U46824 (N_46824,N_42580,N_43065);
and U46825 (N_46825,N_44779,N_43527);
and U46826 (N_46826,N_43889,N_44365);
or U46827 (N_46827,N_42782,N_43210);
xor U46828 (N_46828,N_42807,N_43328);
xor U46829 (N_46829,N_44064,N_43370);
and U46830 (N_46830,N_44216,N_43122);
nor U46831 (N_46831,N_42702,N_44027);
nor U46832 (N_46832,N_44208,N_43126);
and U46833 (N_46833,N_44468,N_42969);
nand U46834 (N_46834,N_44542,N_44771);
nand U46835 (N_46835,N_43034,N_43085);
or U46836 (N_46836,N_43017,N_42870);
and U46837 (N_46837,N_43079,N_44075);
nor U46838 (N_46838,N_42520,N_44234);
xnor U46839 (N_46839,N_44158,N_42752);
or U46840 (N_46840,N_43650,N_43154);
nand U46841 (N_46841,N_43522,N_43797);
and U46842 (N_46842,N_43322,N_43734);
and U46843 (N_46843,N_44497,N_44098);
and U46844 (N_46844,N_42691,N_42917);
xor U46845 (N_46845,N_42740,N_42708);
nor U46846 (N_46846,N_43472,N_44443);
or U46847 (N_46847,N_43369,N_43870);
xnor U46848 (N_46848,N_43754,N_42573);
xnor U46849 (N_46849,N_43457,N_44642);
and U46850 (N_46850,N_43163,N_44078);
xor U46851 (N_46851,N_43044,N_43063);
and U46852 (N_46852,N_44596,N_43846);
nor U46853 (N_46853,N_43119,N_42974);
nand U46854 (N_46854,N_44438,N_43098);
nor U46855 (N_46855,N_43576,N_43663);
or U46856 (N_46856,N_42985,N_44881);
nand U46857 (N_46857,N_42611,N_43122);
nand U46858 (N_46858,N_43558,N_42757);
nand U46859 (N_46859,N_43751,N_44838);
and U46860 (N_46860,N_44005,N_43977);
nor U46861 (N_46861,N_44322,N_43549);
xnor U46862 (N_46862,N_42600,N_43180);
nand U46863 (N_46863,N_43685,N_44140);
or U46864 (N_46864,N_42782,N_43104);
xor U46865 (N_46865,N_42565,N_43427);
or U46866 (N_46866,N_42912,N_44401);
xnor U46867 (N_46867,N_42795,N_42576);
xnor U46868 (N_46868,N_44165,N_42627);
nand U46869 (N_46869,N_42942,N_44885);
nor U46870 (N_46870,N_43090,N_42877);
and U46871 (N_46871,N_43258,N_44049);
nand U46872 (N_46872,N_43566,N_43389);
and U46873 (N_46873,N_44854,N_43376);
xor U46874 (N_46874,N_43213,N_43203);
nor U46875 (N_46875,N_42990,N_44359);
xor U46876 (N_46876,N_43494,N_43306);
xor U46877 (N_46877,N_43746,N_44598);
nor U46878 (N_46878,N_43323,N_43018);
and U46879 (N_46879,N_44293,N_42984);
nor U46880 (N_46880,N_44377,N_43000);
nand U46881 (N_46881,N_43563,N_42534);
nor U46882 (N_46882,N_43751,N_43331);
xnor U46883 (N_46883,N_44722,N_44142);
and U46884 (N_46884,N_42696,N_42686);
xor U46885 (N_46885,N_43344,N_43187);
nand U46886 (N_46886,N_44889,N_43822);
or U46887 (N_46887,N_43664,N_44507);
or U46888 (N_46888,N_43779,N_42975);
and U46889 (N_46889,N_43270,N_43108);
and U46890 (N_46890,N_44533,N_44176);
xnor U46891 (N_46891,N_44894,N_44795);
xor U46892 (N_46892,N_43835,N_44193);
or U46893 (N_46893,N_44386,N_44574);
nand U46894 (N_46894,N_42605,N_43458);
nor U46895 (N_46895,N_44829,N_44114);
nand U46896 (N_46896,N_44835,N_43360);
or U46897 (N_46897,N_43376,N_44011);
nor U46898 (N_46898,N_43597,N_43619);
xor U46899 (N_46899,N_44735,N_43967);
or U46900 (N_46900,N_44022,N_43887);
xor U46901 (N_46901,N_42846,N_44726);
nand U46902 (N_46902,N_43141,N_44733);
or U46903 (N_46903,N_43837,N_43116);
and U46904 (N_46904,N_44774,N_44718);
xor U46905 (N_46905,N_43640,N_42594);
and U46906 (N_46906,N_42840,N_44769);
nand U46907 (N_46907,N_44258,N_43380);
or U46908 (N_46908,N_42738,N_43351);
nor U46909 (N_46909,N_43919,N_43606);
nand U46910 (N_46910,N_44530,N_44093);
or U46911 (N_46911,N_44472,N_44205);
nor U46912 (N_46912,N_42991,N_43656);
nand U46913 (N_46913,N_43981,N_43604);
xor U46914 (N_46914,N_43134,N_44799);
nand U46915 (N_46915,N_43327,N_42734);
nor U46916 (N_46916,N_42837,N_43638);
or U46917 (N_46917,N_43779,N_43864);
nor U46918 (N_46918,N_44865,N_43353);
nand U46919 (N_46919,N_44829,N_42953);
nor U46920 (N_46920,N_43053,N_44253);
or U46921 (N_46921,N_42817,N_42684);
and U46922 (N_46922,N_43702,N_43644);
xnor U46923 (N_46923,N_44508,N_44758);
or U46924 (N_46924,N_44145,N_43930);
nand U46925 (N_46925,N_44285,N_44853);
nand U46926 (N_46926,N_42947,N_43257);
and U46927 (N_46927,N_44854,N_42618);
nand U46928 (N_46928,N_42765,N_44266);
or U46929 (N_46929,N_43907,N_44309);
nor U46930 (N_46930,N_43604,N_42929);
and U46931 (N_46931,N_43630,N_42622);
nand U46932 (N_46932,N_44795,N_42834);
nor U46933 (N_46933,N_44663,N_42537);
or U46934 (N_46934,N_44612,N_44097);
nand U46935 (N_46935,N_43225,N_44261);
xnor U46936 (N_46936,N_43904,N_44755);
nand U46937 (N_46937,N_44895,N_42639);
xnor U46938 (N_46938,N_44574,N_42782);
nand U46939 (N_46939,N_43234,N_42712);
xor U46940 (N_46940,N_43677,N_44782);
and U46941 (N_46941,N_44551,N_43003);
or U46942 (N_46942,N_44348,N_44401);
or U46943 (N_46943,N_42872,N_43311);
xnor U46944 (N_46944,N_42759,N_43012);
and U46945 (N_46945,N_43227,N_43910);
or U46946 (N_46946,N_42594,N_44548);
or U46947 (N_46947,N_42528,N_44599);
nand U46948 (N_46948,N_44962,N_42552);
or U46949 (N_46949,N_44348,N_43221);
nand U46950 (N_46950,N_42911,N_44968);
or U46951 (N_46951,N_43228,N_42725);
and U46952 (N_46952,N_43184,N_43044);
nor U46953 (N_46953,N_44085,N_43974);
xor U46954 (N_46954,N_43618,N_43772);
nand U46955 (N_46955,N_44662,N_43043);
xor U46956 (N_46956,N_43525,N_44588);
nand U46957 (N_46957,N_43809,N_43638);
or U46958 (N_46958,N_44855,N_44516);
and U46959 (N_46959,N_42829,N_44138);
and U46960 (N_46960,N_43070,N_43015);
or U46961 (N_46961,N_44089,N_42544);
or U46962 (N_46962,N_43418,N_44942);
nand U46963 (N_46963,N_42683,N_43208);
and U46964 (N_46964,N_43975,N_44529);
xnor U46965 (N_46965,N_42609,N_43745);
or U46966 (N_46966,N_44614,N_43344);
and U46967 (N_46967,N_44191,N_44182);
and U46968 (N_46968,N_42680,N_43837);
nand U46969 (N_46969,N_44080,N_43854);
nor U46970 (N_46970,N_44703,N_43403);
nand U46971 (N_46971,N_43549,N_43245);
and U46972 (N_46972,N_42730,N_42503);
xor U46973 (N_46973,N_42879,N_44785);
and U46974 (N_46974,N_42766,N_42658);
and U46975 (N_46975,N_43539,N_43804);
and U46976 (N_46976,N_44429,N_43820);
xor U46977 (N_46977,N_42991,N_44776);
nand U46978 (N_46978,N_42966,N_44322);
or U46979 (N_46979,N_44564,N_43920);
nor U46980 (N_46980,N_43315,N_43892);
or U46981 (N_46981,N_44315,N_42954);
and U46982 (N_46982,N_42766,N_44849);
or U46983 (N_46983,N_43623,N_44888);
xor U46984 (N_46984,N_44096,N_44607);
and U46985 (N_46985,N_44563,N_43448);
and U46986 (N_46986,N_42606,N_42777);
xnor U46987 (N_46987,N_43110,N_42506);
nand U46988 (N_46988,N_43313,N_44189);
nand U46989 (N_46989,N_44547,N_44410);
and U46990 (N_46990,N_44888,N_43467);
or U46991 (N_46991,N_43633,N_42618);
xor U46992 (N_46992,N_43798,N_44297);
nand U46993 (N_46993,N_43015,N_43538);
and U46994 (N_46994,N_43114,N_42972);
nor U46995 (N_46995,N_42720,N_42615);
xnor U46996 (N_46996,N_44983,N_43199);
xnor U46997 (N_46997,N_43803,N_44636);
xnor U46998 (N_46998,N_44867,N_44654);
nor U46999 (N_46999,N_42520,N_43763);
nand U47000 (N_47000,N_42971,N_42985);
xor U47001 (N_47001,N_44609,N_44607);
nand U47002 (N_47002,N_44980,N_42969);
nor U47003 (N_47003,N_43379,N_44628);
or U47004 (N_47004,N_43129,N_42851);
nand U47005 (N_47005,N_42554,N_43349);
nand U47006 (N_47006,N_44937,N_44706);
or U47007 (N_47007,N_43818,N_42721);
or U47008 (N_47008,N_42729,N_42689);
nand U47009 (N_47009,N_42590,N_44399);
or U47010 (N_47010,N_43263,N_44397);
and U47011 (N_47011,N_43043,N_44267);
nor U47012 (N_47012,N_42953,N_44544);
nand U47013 (N_47013,N_44049,N_44761);
and U47014 (N_47014,N_44633,N_43377);
nand U47015 (N_47015,N_43844,N_43853);
nand U47016 (N_47016,N_44213,N_43817);
or U47017 (N_47017,N_44176,N_44883);
nand U47018 (N_47018,N_44088,N_44395);
nor U47019 (N_47019,N_43553,N_43440);
or U47020 (N_47020,N_44304,N_44037);
and U47021 (N_47021,N_43555,N_44738);
nand U47022 (N_47022,N_43134,N_42771);
nand U47023 (N_47023,N_44266,N_43801);
or U47024 (N_47024,N_42758,N_43468);
xnor U47025 (N_47025,N_44565,N_44195);
and U47026 (N_47026,N_44916,N_44370);
nor U47027 (N_47027,N_44749,N_44893);
or U47028 (N_47028,N_44246,N_44610);
or U47029 (N_47029,N_43608,N_44554);
and U47030 (N_47030,N_43147,N_43700);
nor U47031 (N_47031,N_44028,N_43782);
or U47032 (N_47032,N_43489,N_43584);
nor U47033 (N_47033,N_43359,N_44624);
nand U47034 (N_47034,N_44186,N_43478);
or U47035 (N_47035,N_42523,N_43956);
nand U47036 (N_47036,N_44530,N_42985);
xor U47037 (N_47037,N_44544,N_42741);
nor U47038 (N_47038,N_43105,N_43121);
nor U47039 (N_47039,N_43965,N_44454);
and U47040 (N_47040,N_44549,N_44177);
xnor U47041 (N_47041,N_44580,N_43964);
nand U47042 (N_47042,N_44673,N_43159);
xnor U47043 (N_47043,N_43558,N_43435);
nand U47044 (N_47044,N_44892,N_42573);
nand U47045 (N_47045,N_43709,N_43162);
and U47046 (N_47046,N_42717,N_44925);
and U47047 (N_47047,N_43146,N_44724);
nand U47048 (N_47048,N_42931,N_43637);
nor U47049 (N_47049,N_44188,N_42585);
nand U47050 (N_47050,N_43782,N_43008);
xor U47051 (N_47051,N_43737,N_43860);
nor U47052 (N_47052,N_43754,N_42927);
xor U47053 (N_47053,N_42757,N_42545);
and U47054 (N_47054,N_43454,N_43992);
xor U47055 (N_47055,N_44834,N_44542);
or U47056 (N_47056,N_43364,N_42535);
and U47057 (N_47057,N_44009,N_43509);
and U47058 (N_47058,N_44414,N_43245);
nand U47059 (N_47059,N_43993,N_43990);
or U47060 (N_47060,N_44866,N_44742);
nand U47061 (N_47061,N_42881,N_43622);
and U47062 (N_47062,N_43656,N_44703);
and U47063 (N_47063,N_44779,N_43786);
or U47064 (N_47064,N_43360,N_43293);
nand U47065 (N_47065,N_44315,N_44850);
nand U47066 (N_47066,N_42626,N_42592);
xor U47067 (N_47067,N_42692,N_44020);
or U47068 (N_47068,N_42564,N_44894);
xor U47069 (N_47069,N_43632,N_43935);
or U47070 (N_47070,N_42856,N_43161);
nand U47071 (N_47071,N_44133,N_42985);
or U47072 (N_47072,N_42895,N_43706);
xor U47073 (N_47073,N_43604,N_43967);
and U47074 (N_47074,N_43382,N_42672);
nand U47075 (N_47075,N_43447,N_44534);
xnor U47076 (N_47076,N_44693,N_43651);
xor U47077 (N_47077,N_43354,N_44128);
and U47078 (N_47078,N_42753,N_42516);
nor U47079 (N_47079,N_44230,N_44244);
nor U47080 (N_47080,N_44249,N_44285);
and U47081 (N_47081,N_42785,N_44047);
or U47082 (N_47082,N_42858,N_44527);
and U47083 (N_47083,N_44264,N_43071);
or U47084 (N_47084,N_43815,N_44652);
xnor U47085 (N_47085,N_43762,N_43860);
xor U47086 (N_47086,N_42778,N_43513);
nand U47087 (N_47087,N_44173,N_44148);
nor U47088 (N_47088,N_42882,N_43086);
xor U47089 (N_47089,N_43197,N_44992);
xor U47090 (N_47090,N_44908,N_42974);
and U47091 (N_47091,N_43829,N_43329);
nor U47092 (N_47092,N_43514,N_42589);
or U47093 (N_47093,N_42785,N_43591);
nand U47094 (N_47094,N_44959,N_43863);
nand U47095 (N_47095,N_44734,N_43884);
or U47096 (N_47096,N_43455,N_44738);
and U47097 (N_47097,N_43864,N_44959);
or U47098 (N_47098,N_43172,N_43092);
or U47099 (N_47099,N_44413,N_44532);
nor U47100 (N_47100,N_44437,N_44489);
nand U47101 (N_47101,N_43018,N_44974);
and U47102 (N_47102,N_43666,N_44174);
or U47103 (N_47103,N_42810,N_43211);
nand U47104 (N_47104,N_43153,N_44328);
nand U47105 (N_47105,N_44372,N_43429);
and U47106 (N_47106,N_42796,N_44415);
and U47107 (N_47107,N_44000,N_42831);
nor U47108 (N_47108,N_43166,N_42869);
and U47109 (N_47109,N_42614,N_42629);
nand U47110 (N_47110,N_43789,N_44556);
or U47111 (N_47111,N_44833,N_42533);
nor U47112 (N_47112,N_42994,N_42937);
xor U47113 (N_47113,N_44666,N_44416);
and U47114 (N_47114,N_42864,N_44534);
nand U47115 (N_47115,N_44631,N_42704);
nand U47116 (N_47116,N_43975,N_42643);
nand U47117 (N_47117,N_44979,N_43985);
nand U47118 (N_47118,N_43198,N_43555);
and U47119 (N_47119,N_43305,N_43187);
xnor U47120 (N_47120,N_43198,N_44999);
or U47121 (N_47121,N_44155,N_44873);
and U47122 (N_47122,N_43236,N_44750);
or U47123 (N_47123,N_43557,N_43603);
nand U47124 (N_47124,N_44843,N_43321);
nor U47125 (N_47125,N_44611,N_44463);
nand U47126 (N_47126,N_42940,N_43511);
and U47127 (N_47127,N_42863,N_44966);
or U47128 (N_47128,N_43760,N_43843);
nor U47129 (N_47129,N_42860,N_43273);
nand U47130 (N_47130,N_44538,N_42603);
nand U47131 (N_47131,N_43206,N_44118);
nand U47132 (N_47132,N_43939,N_43030);
nor U47133 (N_47133,N_44672,N_44346);
nor U47134 (N_47134,N_44481,N_44436);
or U47135 (N_47135,N_44512,N_44046);
or U47136 (N_47136,N_43872,N_44316);
xnor U47137 (N_47137,N_44500,N_43896);
and U47138 (N_47138,N_43579,N_43998);
or U47139 (N_47139,N_43442,N_43913);
nor U47140 (N_47140,N_44376,N_44462);
or U47141 (N_47141,N_43021,N_44564);
xnor U47142 (N_47142,N_44521,N_43362);
or U47143 (N_47143,N_42528,N_44499);
and U47144 (N_47144,N_44594,N_42743);
nor U47145 (N_47145,N_44241,N_44306);
nand U47146 (N_47146,N_44337,N_44721);
and U47147 (N_47147,N_42891,N_43663);
nand U47148 (N_47148,N_42501,N_44548);
or U47149 (N_47149,N_44867,N_44320);
nand U47150 (N_47150,N_42870,N_44806);
or U47151 (N_47151,N_43997,N_43991);
or U47152 (N_47152,N_44916,N_44711);
nand U47153 (N_47153,N_43752,N_43614);
xnor U47154 (N_47154,N_43992,N_43855);
or U47155 (N_47155,N_42863,N_43735);
nor U47156 (N_47156,N_44292,N_43558);
nor U47157 (N_47157,N_44200,N_44901);
nand U47158 (N_47158,N_44873,N_43705);
nand U47159 (N_47159,N_42909,N_44493);
xnor U47160 (N_47160,N_44040,N_43235);
or U47161 (N_47161,N_44158,N_42767);
nand U47162 (N_47162,N_42588,N_43551);
or U47163 (N_47163,N_44032,N_43332);
nor U47164 (N_47164,N_42594,N_43984);
nand U47165 (N_47165,N_44244,N_43202);
or U47166 (N_47166,N_43610,N_43010);
nand U47167 (N_47167,N_43251,N_43525);
nand U47168 (N_47168,N_42543,N_42759);
xor U47169 (N_47169,N_43355,N_44524);
or U47170 (N_47170,N_44627,N_44643);
nor U47171 (N_47171,N_43853,N_43306);
nor U47172 (N_47172,N_43537,N_44587);
or U47173 (N_47173,N_43792,N_42552);
nand U47174 (N_47174,N_44263,N_44821);
or U47175 (N_47175,N_43574,N_43240);
or U47176 (N_47176,N_44291,N_43752);
nand U47177 (N_47177,N_43998,N_44010);
nor U47178 (N_47178,N_43201,N_44895);
nor U47179 (N_47179,N_43794,N_43072);
or U47180 (N_47180,N_43627,N_43273);
nor U47181 (N_47181,N_44572,N_44999);
or U47182 (N_47182,N_44596,N_43452);
or U47183 (N_47183,N_43621,N_42535);
and U47184 (N_47184,N_43693,N_42763);
nand U47185 (N_47185,N_43860,N_42651);
nor U47186 (N_47186,N_43874,N_44398);
nand U47187 (N_47187,N_43337,N_42922);
nor U47188 (N_47188,N_44989,N_42537);
and U47189 (N_47189,N_43881,N_44925);
nor U47190 (N_47190,N_44266,N_43148);
and U47191 (N_47191,N_44858,N_43464);
nand U47192 (N_47192,N_44745,N_43403);
xor U47193 (N_47193,N_42807,N_43234);
and U47194 (N_47194,N_43477,N_42569);
xnor U47195 (N_47195,N_43128,N_44085);
and U47196 (N_47196,N_44844,N_43205);
nor U47197 (N_47197,N_44735,N_43651);
and U47198 (N_47198,N_44256,N_43860);
nor U47199 (N_47199,N_43775,N_44598);
or U47200 (N_47200,N_44884,N_43391);
and U47201 (N_47201,N_44784,N_44703);
nand U47202 (N_47202,N_43370,N_44410);
or U47203 (N_47203,N_44242,N_43667);
nand U47204 (N_47204,N_43872,N_44236);
and U47205 (N_47205,N_42787,N_44534);
nand U47206 (N_47206,N_43794,N_43043);
nand U47207 (N_47207,N_43153,N_43065);
and U47208 (N_47208,N_44255,N_43644);
or U47209 (N_47209,N_42697,N_43487);
and U47210 (N_47210,N_43111,N_43434);
nand U47211 (N_47211,N_43010,N_44919);
xor U47212 (N_47212,N_42630,N_43063);
nand U47213 (N_47213,N_44888,N_43531);
or U47214 (N_47214,N_43562,N_44696);
or U47215 (N_47215,N_44362,N_42990);
nand U47216 (N_47216,N_43266,N_44023);
nand U47217 (N_47217,N_43325,N_44654);
nand U47218 (N_47218,N_43487,N_43971);
or U47219 (N_47219,N_43908,N_44820);
and U47220 (N_47220,N_43048,N_43481);
xor U47221 (N_47221,N_42748,N_43032);
or U47222 (N_47222,N_43231,N_43532);
nand U47223 (N_47223,N_44336,N_43046);
and U47224 (N_47224,N_44130,N_43054);
and U47225 (N_47225,N_43705,N_44520);
or U47226 (N_47226,N_43291,N_43787);
or U47227 (N_47227,N_44667,N_44128);
nand U47228 (N_47228,N_44468,N_43562);
xnor U47229 (N_47229,N_43451,N_42564);
nand U47230 (N_47230,N_42728,N_44270);
or U47231 (N_47231,N_43519,N_44170);
or U47232 (N_47232,N_44198,N_43282);
and U47233 (N_47233,N_44724,N_44818);
nor U47234 (N_47234,N_42760,N_44062);
nand U47235 (N_47235,N_44068,N_42952);
nor U47236 (N_47236,N_44489,N_44648);
and U47237 (N_47237,N_43840,N_43125);
or U47238 (N_47238,N_43054,N_43971);
nand U47239 (N_47239,N_43775,N_43191);
and U47240 (N_47240,N_44458,N_44380);
and U47241 (N_47241,N_43706,N_43363);
nor U47242 (N_47242,N_43518,N_44743);
and U47243 (N_47243,N_42872,N_44534);
and U47244 (N_47244,N_42587,N_43479);
nor U47245 (N_47245,N_42555,N_44883);
nand U47246 (N_47246,N_44514,N_43150);
and U47247 (N_47247,N_44842,N_44539);
or U47248 (N_47248,N_42970,N_44506);
nand U47249 (N_47249,N_44039,N_43221);
xor U47250 (N_47250,N_42612,N_44323);
or U47251 (N_47251,N_43997,N_43929);
nand U47252 (N_47252,N_44512,N_44978);
nor U47253 (N_47253,N_44239,N_43146);
and U47254 (N_47254,N_43300,N_44918);
or U47255 (N_47255,N_44097,N_42845);
and U47256 (N_47256,N_44227,N_43893);
nor U47257 (N_47257,N_42704,N_43010);
and U47258 (N_47258,N_43479,N_43514);
nor U47259 (N_47259,N_44589,N_44756);
or U47260 (N_47260,N_44146,N_42608);
nand U47261 (N_47261,N_42669,N_44961);
or U47262 (N_47262,N_44364,N_44833);
nand U47263 (N_47263,N_44866,N_44939);
and U47264 (N_47264,N_43174,N_42931);
and U47265 (N_47265,N_43845,N_42770);
xnor U47266 (N_47266,N_43243,N_43658);
and U47267 (N_47267,N_42529,N_43400);
nor U47268 (N_47268,N_42592,N_43950);
nand U47269 (N_47269,N_43696,N_42882);
and U47270 (N_47270,N_43562,N_42974);
nand U47271 (N_47271,N_43567,N_43508);
xnor U47272 (N_47272,N_44529,N_44237);
xnor U47273 (N_47273,N_44023,N_43691);
and U47274 (N_47274,N_44316,N_44178);
or U47275 (N_47275,N_43864,N_43922);
xnor U47276 (N_47276,N_42599,N_43435);
or U47277 (N_47277,N_44245,N_43379);
nor U47278 (N_47278,N_42896,N_44756);
nand U47279 (N_47279,N_42503,N_42606);
and U47280 (N_47280,N_44954,N_43135);
xnor U47281 (N_47281,N_44369,N_42876);
xnor U47282 (N_47282,N_44277,N_43653);
or U47283 (N_47283,N_43190,N_44281);
and U47284 (N_47284,N_44100,N_44628);
and U47285 (N_47285,N_43613,N_43475);
xor U47286 (N_47286,N_42935,N_42678);
xor U47287 (N_47287,N_43369,N_44458);
or U47288 (N_47288,N_43413,N_44117);
xnor U47289 (N_47289,N_42747,N_42966);
nor U47290 (N_47290,N_44443,N_44946);
nor U47291 (N_47291,N_43534,N_43130);
xnor U47292 (N_47292,N_44563,N_44861);
and U47293 (N_47293,N_43655,N_43333);
xnor U47294 (N_47294,N_43670,N_44585);
xnor U47295 (N_47295,N_43366,N_43660);
or U47296 (N_47296,N_44449,N_43253);
nor U47297 (N_47297,N_44285,N_42849);
xnor U47298 (N_47298,N_42760,N_44377);
nand U47299 (N_47299,N_44120,N_43339);
or U47300 (N_47300,N_44953,N_42596);
or U47301 (N_47301,N_44861,N_42918);
nand U47302 (N_47302,N_43841,N_44129);
or U47303 (N_47303,N_43380,N_42562);
nor U47304 (N_47304,N_44707,N_43992);
xor U47305 (N_47305,N_44132,N_43604);
nand U47306 (N_47306,N_44889,N_42625);
nor U47307 (N_47307,N_42732,N_43139);
nand U47308 (N_47308,N_44867,N_42932);
xnor U47309 (N_47309,N_42703,N_43888);
nor U47310 (N_47310,N_43109,N_44997);
nand U47311 (N_47311,N_44712,N_43045);
or U47312 (N_47312,N_42683,N_43325);
nor U47313 (N_47313,N_42574,N_43352);
nor U47314 (N_47314,N_42618,N_44464);
nor U47315 (N_47315,N_44245,N_44956);
nand U47316 (N_47316,N_44623,N_43322);
nor U47317 (N_47317,N_42651,N_44772);
or U47318 (N_47318,N_44285,N_43096);
or U47319 (N_47319,N_44909,N_43841);
or U47320 (N_47320,N_44033,N_43791);
xnor U47321 (N_47321,N_43994,N_44364);
xor U47322 (N_47322,N_44909,N_42653);
or U47323 (N_47323,N_43737,N_43888);
xor U47324 (N_47324,N_43166,N_44512);
nor U47325 (N_47325,N_42513,N_43843);
xor U47326 (N_47326,N_44535,N_43358);
nor U47327 (N_47327,N_43468,N_44379);
nor U47328 (N_47328,N_44898,N_43832);
nor U47329 (N_47329,N_44154,N_43356);
and U47330 (N_47330,N_42791,N_43217);
or U47331 (N_47331,N_42701,N_44974);
or U47332 (N_47332,N_44874,N_44863);
nand U47333 (N_47333,N_44544,N_42955);
and U47334 (N_47334,N_44465,N_44657);
nand U47335 (N_47335,N_43003,N_43704);
nand U47336 (N_47336,N_43643,N_43688);
and U47337 (N_47337,N_44300,N_43750);
and U47338 (N_47338,N_43791,N_42943);
and U47339 (N_47339,N_43473,N_44067);
xnor U47340 (N_47340,N_44937,N_44481);
xnor U47341 (N_47341,N_44529,N_43262);
nor U47342 (N_47342,N_42678,N_42515);
nand U47343 (N_47343,N_43851,N_43287);
nor U47344 (N_47344,N_42692,N_43939);
xor U47345 (N_47345,N_43905,N_42704);
nor U47346 (N_47346,N_44373,N_44657);
xnor U47347 (N_47347,N_43344,N_42593);
xor U47348 (N_47348,N_43924,N_43575);
or U47349 (N_47349,N_44758,N_43420);
or U47350 (N_47350,N_44080,N_43292);
nand U47351 (N_47351,N_42885,N_43507);
nand U47352 (N_47352,N_42970,N_44112);
nor U47353 (N_47353,N_44393,N_44215);
nand U47354 (N_47354,N_44041,N_44617);
xnor U47355 (N_47355,N_44680,N_44815);
xnor U47356 (N_47356,N_43657,N_44980);
or U47357 (N_47357,N_43912,N_43152);
nand U47358 (N_47358,N_44712,N_44180);
and U47359 (N_47359,N_43501,N_44277);
nand U47360 (N_47360,N_44864,N_44811);
and U47361 (N_47361,N_42684,N_44958);
nand U47362 (N_47362,N_42913,N_43727);
xor U47363 (N_47363,N_43002,N_43878);
and U47364 (N_47364,N_42898,N_44631);
or U47365 (N_47365,N_43208,N_42596);
and U47366 (N_47366,N_44706,N_42660);
or U47367 (N_47367,N_43731,N_43390);
and U47368 (N_47368,N_43239,N_42970);
xor U47369 (N_47369,N_43866,N_43707);
nand U47370 (N_47370,N_43509,N_44037);
nor U47371 (N_47371,N_44892,N_43937);
nor U47372 (N_47372,N_43742,N_42606);
or U47373 (N_47373,N_43833,N_44966);
nand U47374 (N_47374,N_44540,N_42843);
nor U47375 (N_47375,N_44746,N_44415);
nor U47376 (N_47376,N_44839,N_43900);
or U47377 (N_47377,N_43740,N_43063);
or U47378 (N_47378,N_42853,N_44581);
and U47379 (N_47379,N_43801,N_43467);
nor U47380 (N_47380,N_43212,N_43236);
and U47381 (N_47381,N_44150,N_43652);
or U47382 (N_47382,N_44450,N_44381);
nand U47383 (N_47383,N_43611,N_44905);
nor U47384 (N_47384,N_44526,N_44008);
and U47385 (N_47385,N_42509,N_42770);
nand U47386 (N_47386,N_43490,N_43672);
or U47387 (N_47387,N_44423,N_44100);
nand U47388 (N_47388,N_43369,N_44959);
nor U47389 (N_47389,N_43032,N_43203);
or U47390 (N_47390,N_44378,N_44912);
and U47391 (N_47391,N_42825,N_43908);
and U47392 (N_47392,N_43552,N_42720);
or U47393 (N_47393,N_44124,N_43233);
nand U47394 (N_47394,N_43115,N_44640);
or U47395 (N_47395,N_44151,N_43882);
xnor U47396 (N_47396,N_44417,N_44931);
or U47397 (N_47397,N_43960,N_43320);
and U47398 (N_47398,N_43150,N_42958);
nor U47399 (N_47399,N_44353,N_43055);
nor U47400 (N_47400,N_44629,N_44634);
and U47401 (N_47401,N_44237,N_43125);
or U47402 (N_47402,N_43159,N_43528);
or U47403 (N_47403,N_44186,N_44437);
nand U47404 (N_47404,N_44725,N_43458);
nand U47405 (N_47405,N_44724,N_44610);
xnor U47406 (N_47406,N_42503,N_43420);
nand U47407 (N_47407,N_43137,N_44064);
or U47408 (N_47408,N_44119,N_43175);
or U47409 (N_47409,N_44774,N_44953);
and U47410 (N_47410,N_44385,N_42882);
and U47411 (N_47411,N_43102,N_44492);
xor U47412 (N_47412,N_43535,N_42560);
nor U47413 (N_47413,N_44418,N_44509);
and U47414 (N_47414,N_44994,N_42891);
nand U47415 (N_47415,N_42660,N_43169);
xnor U47416 (N_47416,N_44175,N_42673);
nand U47417 (N_47417,N_43964,N_43526);
xor U47418 (N_47418,N_42910,N_44536);
or U47419 (N_47419,N_42870,N_43893);
and U47420 (N_47420,N_44816,N_44823);
nor U47421 (N_47421,N_44343,N_43966);
nor U47422 (N_47422,N_44801,N_44771);
xor U47423 (N_47423,N_44799,N_44917);
nor U47424 (N_47424,N_44648,N_43134);
and U47425 (N_47425,N_43060,N_43258);
xnor U47426 (N_47426,N_43068,N_43658);
nor U47427 (N_47427,N_42716,N_44368);
and U47428 (N_47428,N_44974,N_43737);
or U47429 (N_47429,N_44847,N_44775);
and U47430 (N_47430,N_43110,N_44061);
nand U47431 (N_47431,N_44863,N_42826);
or U47432 (N_47432,N_43878,N_44343);
or U47433 (N_47433,N_44412,N_44674);
xor U47434 (N_47434,N_43025,N_43073);
or U47435 (N_47435,N_42889,N_44562);
or U47436 (N_47436,N_43357,N_44289);
or U47437 (N_47437,N_44524,N_44708);
or U47438 (N_47438,N_44955,N_44556);
or U47439 (N_47439,N_44021,N_43849);
nand U47440 (N_47440,N_42721,N_43314);
xnor U47441 (N_47441,N_43825,N_44092);
xnor U47442 (N_47442,N_42521,N_44511);
nor U47443 (N_47443,N_44430,N_43137);
xor U47444 (N_47444,N_44447,N_44288);
nor U47445 (N_47445,N_43647,N_44099);
or U47446 (N_47446,N_44462,N_43258);
or U47447 (N_47447,N_43695,N_44330);
or U47448 (N_47448,N_43189,N_43188);
and U47449 (N_47449,N_42500,N_43787);
xnor U47450 (N_47450,N_43135,N_44169);
or U47451 (N_47451,N_44644,N_44139);
xor U47452 (N_47452,N_43519,N_44659);
nor U47453 (N_47453,N_43842,N_43665);
and U47454 (N_47454,N_42851,N_42674);
or U47455 (N_47455,N_43990,N_43817);
nand U47456 (N_47456,N_43856,N_44575);
or U47457 (N_47457,N_43069,N_42549);
nand U47458 (N_47458,N_43349,N_43465);
nor U47459 (N_47459,N_43770,N_44307);
and U47460 (N_47460,N_43894,N_44407);
nand U47461 (N_47461,N_44502,N_44334);
nand U47462 (N_47462,N_44595,N_44424);
or U47463 (N_47463,N_44074,N_44267);
nor U47464 (N_47464,N_44081,N_44574);
xnor U47465 (N_47465,N_43846,N_44495);
xnor U47466 (N_47466,N_42780,N_43966);
xnor U47467 (N_47467,N_42680,N_43076);
or U47468 (N_47468,N_44712,N_42914);
nand U47469 (N_47469,N_43769,N_43521);
or U47470 (N_47470,N_44458,N_44753);
nand U47471 (N_47471,N_44646,N_43592);
xnor U47472 (N_47472,N_44857,N_43164);
or U47473 (N_47473,N_42839,N_42646);
nor U47474 (N_47474,N_43711,N_43540);
nor U47475 (N_47475,N_42884,N_42952);
xnor U47476 (N_47476,N_43066,N_42736);
xor U47477 (N_47477,N_43612,N_42692);
and U47478 (N_47478,N_44691,N_43116);
nor U47479 (N_47479,N_42664,N_44537);
xnor U47480 (N_47480,N_44954,N_44155);
or U47481 (N_47481,N_43216,N_42718);
or U47482 (N_47482,N_44375,N_44772);
nor U47483 (N_47483,N_43039,N_43695);
nand U47484 (N_47484,N_42551,N_42728);
xnor U47485 (N_47485,N_44589,N_43482);
nand U47486 (N_47486,N_43085,N_43434);
nand U47487 (N_47487,N_44003,N_43228);
nor U47488 (N_47488,N_43582,N_43660);
and U47489 (N_47489,N_42964,N_43242);
or U47490 (N_47490,N_43386,N_44123);
and U47491 (N_47491,N_42974,N_44569);
xor U47492 (N_47492,N_42979,N_43962);
xor U47493 (N_47493,N_42639,N_43206);
and U47494 (N_47494,N_43389,N_43070);
xnor U47495 (N_47495,N_44046,N_42741);
nand U47496 (N_47496,N_42867,N_42892);
and U47497 (N_47497,N_42731,N_43471);
or U47498 (N_47498,N_42880,N_43656);
nand U47499 (N_47499,N_44564,N_44854);
xnor U47500 (N_47500,N_47041,N_46355);
or U47501 (N_47501,N_46099,N_45657);
and U47502 (N_47502,N_46799,N_45852);
or U47503 (N_47503,N_47478,N_46402);
nand U47504 (N_47504,N_45286,N_46165);
or U47505 (N_47505,N_46352,N_45388);
nand U47506 (N_47506,N_46228,N_45382);
and U47507 (N_47507,N_46568,N_47479);
nor U47508 (N_47508,N_45512,N_46337);
or U47509 (N_47509,N_45648,N_45617);
nand U47510 (N_47510,N_46199,N_45797);
nor U47511 (N_47511,N_46862,N_47317);
nand U47512 (N_47512,N_45924,N_45149);
nand U47513 (N_47513,N_46774,N_46012);
xor U47514 (N_47514,N_46676,N_47440);
nand U47515 (N_47515,N_45975,N_45554);
xor U47516 (N_47516,N_46324,N_46223);
or U47517 (N_47517,N_45997,N_45386);
nand U47518 (N_47518,N_46122,N_46481);
nor U47519 (N_47519,N_46020,N_46921);
nor U47520 (N_47520,N_45171,N_46156);
xnor U47521 (N_47521,N_46196,N_45047);
nor U47522 (N_47522,N_45285,N_46398);
xor U47523 (N_47523,N_47212,N_45435);
or U47524 (N_47524,N_45375,N_46823);
nor U47525 (N_47525,N_46654,N_46954);
xor U47526 (N_47526,N_47249,N_46691);
and U47527 (N_47527,N_46150,N_45760);
nand U47528 (N_47528,N_47059,N_45489);
nand U47529 (N_47529,N_45390,N_46760);
xor U47530 (N_47530,N_47449,N_46282);
nor U47531 (N_47531,N_46773,N_45459);
xnor U47532 (N_47532,N_45707,N_46916);
nor U47533 (N_47533,N_46567,N_45332);
xnor U47534 (N_47534,N_47241,N_45800);
or U47535 (N_47535,N_45372,N_45102);
nor U47536 (N_47536,N_45619,N_45984);
or U47537 (N_47537,N_45548,N_47339);
nor U47538 (N_47538,N_46872,N_45625);
or U47539 (N_47539,N_46838,N_47211);
nor U47540 (N_47540,N_45170,N_45727);
nor U47541 (N_47541,N_45376,N_45414);
nor U47542 (N_47542,N_46254,N_45497);
xor U47543 (N_47543,N_45508,N_47204);
nor U47544 (N_47544,N_47409,N_47065);
and U47545 (N_47545,N_45348,N_45563);
xor U47546 (N_47546,N_45603,N_45338);
nor U47547 (N_47547,N_45865,N_45598);
or U47548 (N_47548,N_45493,N_47288);
xnor U47549 (N_47549,N_45889,N_46794);
or U47550 (N_47550,N_45343,N_47218);
nand U47551 (N_47551,N_47124,N_45484);
or U47552 (N_47552,N_46325,N_46335);
or U47553 (N_47553,N_47246,N_45736);
xnor U47554 (N_47554,N_46029,N_47025);
or U47555 (N_47555,N_46261,N_45274);
nand U47556 (N_47556,N_46217,N_45881);
nand U47557 (N_47557,N_46442,N_46317);
or U47558 (N_47558,N_46665,N_45642);
xor U47559 (N_47559,N_45296,N_45798);
xor U47560 (N_47560,N_45306,N_47399);
nor U47561 (N_47561,N_45206,N_46790);
nor U47562 (N_47562,N_46775,N_46582);
nor U47563 (N_47563,N_47370,N_47395);
nor U47564 (N_47564,N_46108,N_45037);
nor U47565 (N_47565,N_46057,N_46844);
xnor U47566 (N_47566,N_45662,N_47032);
or U47567 (N_47567,N_46070,N_46024);
nor U47568 (N_47568,N_47360,N_47049);
and U47569 (N_47569,N_46763,N_45048);
nor U47570 (N_47570,N_45240,N_45530);
nand U47571 (N_47571,N_46717,N_46801);
nor U47572 (N_47572,N_46544,N_45947);
nand U47573 (N_47573,N_45265,N_45911);
and U47574 (N_47574,N_46967,N_46171);
and U47575 (N_47575,N_47203,N_46450);
xnor U47576 (N_47576,N_45153,N_46569);
and U47577 (N_47577,N_46472,N_47183);
nor U47578 (N_47578,N_47263,N_45453);
or U47579 (N_47579,N_45537,N_46501);
nand U47580 (N_47580,N_46634,N_46572);
or U47581 (N_47581,N_45117,N_45620);
and U47582 (N_47582,N_47092,N_46283);
nand U47583 (N_47583,N_46419,N_47105);
xnor U47584 (N_47584,N_47293,N_46269);
nand U47585 (N_47585,N_46725,N_45927);
or U47586 (N_47586,N_46966,N_45813);
or U47587 (N_47587,N_46265,N_47470);
nor U47588 (N_47588,N_46396,N_45495);
and U47589 (N_47589,N_46868,N_47029);
nor U47590 (N_47590,N_45886,N_46574);
xnor U47591 (N_47591,N_45829,N_46158);
nor U47592 (N_47592,N_45143,N_47345);
nand U47593 (N_47593,N_45570,N_45860);
xnor U47594 (N_47594,N_46278,N_47134);
nor U47595 (N_47595,N_45267,N_46362);
nand U47596 (N_47596,N_46015,N_46004);
nand U47597 (N_47597,N_45576,N_47337);
nor U47598 (N_47598,N_45328,N_47496);
nor U47599 (N_47599,N_47385,N_45590);
nand U47600 (N_47600,N_46575,N_46128);
or U47601 (N_47601,N_46837,N_47490);
or U47602 (N_47602,N_47300,N_47443);
or U47603 (N_47603,N_45472,N_46959);
nor U47604 (N_47604,N_45297,N_45091);
and U47605 (N_47605,N_45588,N_46898);
xor U47606 (N_47606,N_46886,N_46458);
nor U47607 (N_47607,N_45669,N_46348);
or U47608 (N_47608,N_46590,N_47018);
and U47609 (N_47609,N_46144,N_45200);
or U47610 (N_47610,N_47027,N_46752);
nand U47611 (N_47611,N_47486,N_47022);
nor U47612 (N_47612,N_45364,N_46615);
and U47613 (N_47613,N_46891,N_45611);
nor U47614 (N_47614,N_45049,N_46573);
and U47615 (N_47615,N_47031,N_47289);
nor U47616 (N_47616,N_45515,N_45458);
nor U47617 (N_47617,N_47464,N_45849);
nand U47618 (N_47618,N_45845,N_45202);
xor U47619 (N_47619,N_45953,N_45340);
nand U47620 (N_47620,N_45945,N_47233);
nand U47621 (N_47621,N_45215,N_46422);
nor U47622 (N_47622,N_46816,N_45269);
nor U47623 (N_47623,N_46599,N_45966);
nor U47624 (N_47624,N_45719,N_46761);
xnor U47625 (N_47625,N_46277,N_46330);
and U47626 (N_47626,N_45197,N_47149);
nand U47627 (N_47627,N_46424,N_45226);
nor U47628 (N_47628,N_45794,N_46197);
nor U47629 (N_47629,N_47026,N_45418);
xor U47630 (N_47630,N_45094,N_45958);
and U47631 (N_47631,N_46849,N_46043);
or U47632 (N_47632,N_45228,N_45580);
xor U47633 (N_47633,N_45347,N_45161);
xor U47634 (N_47634,N_47209,N_47167);
xnor U47635 (N_47635,N_45146,N_47111);
and U47636 (N_47636,N_46174,N_46386);
nor U47637 (N_47637,N_47202,N_46133);
or U47638 (N_47638,N_46680,N_46280);
nor U47639 (N_47639,N_45535,N_46409);
nand U47640 (N_47640,N_46384,N_46475);
xor U47641 (N_47641,N_47445,N_45893);
and U47642 (N_47642,N_46484,N_47356);
nand U47643 (N_47643,N_47348,N_45956);
nand U47644 (N_47644,N_46098,N_45632);
and U47645 (N_47645,N_47043,N_46477);
xor U47646 (N_47646,N_45618,N_45943);
nand U47647 (N_47647,N_45686,N_45661);
nand U47648 (N_47648,N_46579,N_46668);
xnor U47649 (N_47649,N_47067,N_45636);
and U47650 (N_47650,N_46366,N_45071);
xnor U47651 (N_47651,N_45747,N_45990);
nor U47652 (N_47652,N_47116,N_45791);
nor U47653 (N_47653,N_46955,N_46183);
or U47654 (N_47654,N_45008,N_46909);
xor U47655 (N_47655,N_46048,N_47215);
xnor U47656 (N_47656,N_46192,N_45859);
or U47657 (N_47657,N_46440,N_45068);
xnor U47658 (N_47658,N_45216,N_47351);
nand U47659 (N_47659,N_45635,N_45142);
nor U47660 (N_47660,N_47103,N_45804);
and U47661 (N_47661,N_47201,N_46910);
and U47662 (N_47662,N_45962,N_45052);
nor U47663 (N_47663,N_45607,N_45626);
and U47664 (N_47664,N_45908,N_46787);
or U47665 (N_47665,N_47007,N_45688);
xor U47666 (N_47666,N_45383,N_47061);
or U47667 (N_47667,N_46163,N_47028);
or U47668 (N_47668,N_45868,N_47467);
and U47669 (N_47669,N_47117,N_46646);
nor U47670 (N_47670,N_45126,N_47423);
or U47671 (N_47671,N_46427,N_45028);
and U47672 (N_47672,N_47210,N_46081);
or U47673 (N_47673,N_46190,N_46353);
xor U47674 (N_47674,N_45043,N_47431);
xnor U47675 (N_47675,N_47138,N_46310);
nor U47676 (N_47676,N_45536,N_46834);
xnor U47677 (N_47677,N_45787,N_45345);
and U47678 (N_47678,N_46167,N_47035);
nor U47679 (N_47679,N_47133,N_45124);
or U47680 (N_47680,N_47427,N_45120);
xor U47681 (N_47681,N_46902,N_47268);
nand U47682 (N_47682,N_47331,N_45898);
or U47683 (N_47683,N_46227,N_47097);
or U47684 (N_47684,N_45644,N_45315);
nor U47685 (N_47685,N_46919,N_45641);
nand U47686 (N_47686,N_45704,N_45780);
or U47687 (N_47687,N_46857,N_46006);
nor U47688 (N_47688,N_47161,N_46389);
nand U47689 (N_47689,N_46947,N_45211);
nor U47690 (N_47690,N_47400,N_45457);
xnor U47691 (N_47691,N_45569,N_45987);
xor U47692 (N_47692,N_45327,N_45505);
xor U47693 (N_47693,N_46956,N_47272);
nor U47694 (N_47694,N_46843,N_46072);
nand U47695 (N_47695,N_45768,N_45322);
xor U47696 (N_47696,N_46251,N_46581);
nor U47697 (N_47697,N_46711,N_45394);
xnor U47698 (N_47698,N_46965,N_47039);
nand U47699 (N_47699,N_45991,N_45424);
and U47700 (N_47700,N_45498,N_45708);
nand U47701 (N_47701,N_46306,N_46023);
nand U47702 (N_47702,N_46333,N_47159);
nand U47703 (N_47703,N_45770,N_45125);
or U47704 (N_47704,N_47315,N_47240);
and U47705 (N_47705,N_45317,N_47160);
and U47706 (N_47706,N_45182,N_47324);
xor U47707 (N_47707,N_45359,N_46627);
and U47708 (N_47708,N_46981,N_47376);
nand U47709 (N_47709,N_46840,N_45925);
and U47710 (N_47710,N_45754,N_47066);
and U47711 (N_47711,N_45235,N_46038);
nand U47712 (N_47712,N_47454,N_46874);
xnor U47713 (N_47713,N_46314,N_45932);
nor U47714 (N_47714,N_46155,N_45951);
and U47715 (N_47715,N_45089,N_46187);
xnor U47716 (N_47716,N_45693,N_45410);
nor U47717 (N_47717,N_46082,N_46548);
or U47718 (N_47718,N_45788,N_45176);
xnor U47719 (N_47719,N_45887,N_46974);
or U47720 (N_47720,N_45069,N_47005);
and U47721 (N_47721,N_46364,N_46796);
xnor U47722 (N_47722,N_46944,N_46999);
nand U47723 (N_47723,N_46776,N_45050);
xor U47724 (N_47724,N_45273,N_46851);
or U47725 (N_47725,N_47270,N_46385);
or U47726 (N_47726,N_45078,N_45259);
and U47727 (N_47727,N_45963,N_45428);
and U47728 (N_47728,N_45731,N_46757);
or U47729 (N_47729,N_45287,N_46336);
and U47730 (N_47730,N_45012,N_47274);
and U47731 (N_47731,N_46215,N_47081);
xnor U47732 (N_47732,N_46554,N_45702);
nand U47733 (N_47733,N_47230,N_45423);
and U47734 (N_47734,N_46119,N_45298);
or U47735 (N_47735,N_46011,N_45503);
nand U47736 (N_47736,N_46139,N_45398);
and U47737 (N_47737,N_46970,N_46556);
nor U47738 (N_47738,N_47308,N_47190);
and U47739 (N_47739,N_45746,N_45716);
nand U47740 (N_47740,N_46800,N_45807);
nand U47741 (N_47741,N_46264,N_46617);
or U47742 (N_47742,N_47350,N_45450);
and U47743 (N_47743,N_46123,N_46658);
nand U47744 (N_47744,N_47238,N_45329);
xor U47745 (N_47745,N_45729,N_45201);
and U47746 (N_47746,N_46541,N_45204);
xnor U47747 (N_47747,N_46211,N_46958);
xor U47748 (N_47748,N_46037,N_46244);
xor U47749 (N_47749,N_46263,N_46625);
and U47750 (N_47750,N_45264,N_46421);
and U47751 (N_47751,N_46381,N_46455);
and U47752 (N_47752,N_45682,N_46670);
nor U47753 (N_47753,N_45998,N_45035);
or U47754 (N_47754,N_46830,N_46542);
or U47755 (N_47755,N_45272,N_45853);
nor U47756 (N_47756,N_45342,N_47329);
nor U47757 (N_47757,N_46168,N_45681);
and U47758 (N_47758,N_46297,N_45465);
nand U47759 (N_47759,N_45792,N_46019);
or U47760 (N_47760,N_45511,N_45725);
xnor U47761 (N_47761,N_47387,N_46273);
nor U47762 (N_47762,N_45628,N_45335);
or U47763 (N_47763,N_46061,N_46041);
nand U47764 (N_47764,N_45742,N_47327);
nor U47765 (N_47765,N_46587,N_45130);
xor U47766 (N_47766,N_45610,N_45647);
or U47767 (N_47767,N_45544,N_47229);
or U47768 (N_47768,N_46311,N_45930);
and U47769 (N_47769,N_46430,N_45584);
or U47770 (N_47770,N_45821,N_47070);
xnor U47771 (N_47771,N_46594,N_46588);
or U47772 (N_47772,N_46049,N_45882);
xor U47773 (N_47773,N_46439,N_47282);
nand U47774 (N_47774,N_47355,N_45637);
nor U47775 (N_47775,N_46447,N_47176);
nor U47776 (N_47776,N_47307,N_45769);
nand U47777 (N_47777,N_46560,N_45468);
nor U47778 (N_47778,N_46201,N_47413);
nor U47779 (N_47779,N_45038,N_46734);
or U47780 (N_47780,N_46968,N_47453);
nand U47781 (N_47781,N_47334,N_47362);
xor U47782 (N_47782,N_46678,N_45026);
or U47783 (N_47783,N_46855,N_46116);
or U47784 (N_47784,N_46690,N_46570);
nor U47785 (N_47785,N_47325,N_46929);
xor U47786 (N_47786,N_45802,N_45982);
or U47787 (N_47787,N_45353,N_46847);
nor U47788 (N_47788,N_45336,N_47353);
and U47789 (N_47789,N_46495,N_46731);
or U47790 (N_47790,N_46810,N_47471);
nor U47791 (N_47791,N_46022,N_46259);
or U47792 (N_47792,N_45596,N_46606);
nand U47793 (N_47793,N_46688,N_47011);
and U47794 (N_47794,N_46404,N_45278);
or U47795 (N_47795,N_47237,N_45004);
xor U47796 (N_47796,N_45163,N_47402);
or U47797 (N_47797,N_46933,N_47141);
nand U47798 (N_47798,N_47302,N_46071);
nand U47799 (N_47799,N_46681,N_46002);
or U47800 (N_47800,N_45021,N_45018);
xnor U47801 (N_47801,N_45502,N_46808);
and U47802 (N_47802,N_46613,N_47472);
nor U47803 (N_47803,N_45977,N_45973);
xnor U47804 (N_47804,N_45462,N_45413);
nand U47805 (N_47805,N_45407,N_46492);
and U47806 (N_47806,N_46789,N_47436);
nand U47807 (N_47807,N_46528,N_46418);
and U47808 (N_47808,N_45397,N_46453);
xor U47809 (N_47809,N_46976,N_45695);
and U47810 (N_47810,N_45121,N_46347);
xnor U47811 (N_47811,N_46846,N_46637);
xnor U47812 (N_47812,N_46946,N_46812);
or U47813 (N_47813,N_45250,N_45587);
or U47814 (N_47814,N_47231,N_47421);
nor U47815 (N_47815,N_47119,N_46301);
nand U47816 (N_47816,N_46060,N_47450);
or U47817 (N_47817,N_45473,N_45876);
nor U47818 (N_47818,N_46879,N_45475);
nand U47819 (N_47819,N_46591,N_46644);
nor U47820 (N_47820,N_46236,N_46302);
nor U47821 (N_47821,N_47122,N_46675);
or U47822 (N_47822,N_45949,N_47216);
nor U47823 (N_47823,N_45942,N_45151);
xor U47824 (N_47824,N_46531,N_47038);
and U47825 (N_47825,N_45295,N_46601);
xor U47826 (N_47826,N_45756,N_47250);
xor U47827 (N_47827,N_47247,N_45492);
or U47828 (N_47828,N_45152,N_45350);
or U47829 (N_47829,N_47239,N_45850);
nand U47830 (N_47830,N_45717,N_45673);
nor U47831 (N_47831,N_46985,N_46126);
nor U47832 (N_47832,N_46861,N_46718);
xor U47833 (N_47833,N_47180,N_46166);
nand U47834 (N_47834,N_45878,N_47298);
or U47835 (N_47835,N_47390,N_45401);
and U47836 (N_47836,N_46189,N_45679);
nand U47837 (N_47837,N_45811,N_45959);
nor U47838 (N_47838,N_46137,N_45749);
and U47839 (N_47839,N_46674,N_47137);
xnor U47840 (N_47840,N_45801,N_45779);
nor U47841 (N_47841,N_45365,N_47046);
or U47842 (N_47842,N_45758,N_45324);
nor U47843 (N_47843,N_46488,N_45744);
nor U47844 (N_47844,N_45903,N_45281);
nand U47845 (N_47845,N_46883,N_45373);
nand U47846 (N_47846,N_46343,N_47087);
or U47847 (N_47847,N_45039,N_46331);
xnor U47848 (N_47848,N_47392,N_46899);
xor U47849 (N_47849,N_45155,N_46360);
nor U47850 (N_47850,N_46287,N_46719);
xor U47851 (N_47851,N_46964,N_45592);
and U47852 (N_47852,N_45545,N_46512);
xnor U47853 (N_47853,N_45141,N_46181);
xnor U47854 (N_47854,N_46509,N_46724);
xnor U47855 (N_47855,N_45782,N_46177);
nand U47856 (N_47856,N_46040,N_46247);
and U47857 (N_47857,N_45507,N_47276);
and U47858 (N_47858,N_45456,N_46989);
nor U47859 (N_47859,N_47352,N_45477);
and U47860 (N_47860,N_45169,N_46520);
nand U47861 (N_47861,N_45223,N_46322);
or U47862 (N_47862,N_46927,N_47148);
or U47863 (N_47863,N_47044,N_46334);
nand U47864 (N_47864,N_47379,N_46432);
and U47865 (N_47865,N_45586,N_46864);
nand U47866 (N_47866,N_45292,N_45349);
nor U47867 (N_47867,N_46505,N_45422);
nand U47868 (N_47868,N_45869,N_47121);
and U47869 (N_47869,N_47401,N_46094);
xnor U47870 (N_47870,N_47438,N_46180);
nand U47871 (N_47871,N_45086,N_45344);
and U47872 (N_47872,N_46235,N_46349);
nor U47873 (N_47873,N_47197,N_46521);
xor U47874 (N_47874,N_46961,N_45271);
or U47875 (N_47875,N_46704,N_47320);
and U47876 (N_47876,N_46755,N_46697);
nand U47877 (N_47877,N_45217,N_46257);
and U47878 (N_47878,N_47085,N_45391);
nand U47879 (N_47879,N_46397,N_46824);
nor U47880 (N_47880,N_46924,N_45241);
or U47881 (N_47881,N_45525,N_46772);
nor U47882 (N_47882,N_45723,N_46661);
nand U47883 (N_47883,N_46622,N_45188);
and U47884 (N_47884,N_46417,N_47226);
and U47885 (N_47885,N_45985,N_46701);
or U47886 (N_47886,N_45366,N_45168);
nand U47887 (N_47887,N_46683,N_46434);
nand U47888 (N_47888,N_46125,N_47013);
nor U47889 (N_47889,N_47264,N_45989);
nand U47890 (N_47890,N_45416,N_46727);
or U47891 (N_47891,N_47484,N_46293);
or U47892 (N_47892,N_45931,N_47393);
or U47893 (N_47893,N_45894,N_46523);
or U47894 (N_47894,N_47182,N_45016);
and U47895 (N_47895,N_45670,N_46739);
or U47896 (N_47896,N_46062,N_46001);
and U47897 (N_47897,N_47223,N_45581);
nand U47898 (N_47898,N_46825,N_45741);
and U47899 (N_47899,N_46925,N_46785);
nand U47900 (N_47900,N_47483,N_46890);
and U47901 (N_47901,N_45463,N_46744);
nand U47902 (N_47902,N_45195,N_45015);
nand U47903 (N_47903,N_45178,N_47030);
nand U47904 (N_47904,N_46221,N_46344);
nand U47905 (N_47905,N_46239,N_46149);
nor U47906 (N_47906,N_47075,N_46241);
and U47907 (N_47907,N_46841,N_45560);
nand U47908 (N_47908,N_45730,N_45109);
nor U47909 (N_47909,N_45726,N_47297);
nor U47910 (N_47910,N_45995,N_45466);
or U47911 (N_47911,N_46246,N_45805);
nor U47912 (N_47912,N_46547,N_46372);
and U47913 (N_47913,N_46873,N_45950);
nor U47914 (N_47914,N_47143,N_46741);
and U47915 (N_47915,N_47369,N_45743);
nand U47916 (N_47916,N_45356,N_46249);
xnor U47917 (N_47917,N_47474,N_45270);
nand U47918 (N_47918,N_45764,N_47146);
and U47919 (N_47919,N_45290,N_46905);
or U47920 (N_47920,N_47073,N_47466);
and U47921 (N_47921,N_45253,N_46949);
nand U47922 (N_47922,N_46435,N_45752);
nor U47923 (N_47923,N_45119,N_47155);
xor U47924 (N_47924,N_45482,N_45843);
and U47925 (N_47925,N_45280,N_46391);
xor U47926 (N_47926,N_45072,N_45885);
and U47927 (N_47927,N_46142,N_45645);
or U47928 (N_47928,N_46405,N_46498);
xnor U47929 (N_47929,N_45833,N_47433);
or U47930 (N_47930,N_46457,N_46903);
nor U47931 (N_47931,N_45935,N_47126);
nand U47932 (N_47932,N_45460,N_46563);
nor U47933 (N_47933,N_45313,N_46111);
or U47934 (N_47934,N_47213,N_47336);
and U47935 (N_47935,N_47068,N_46401);
or U47936 (N_47936,N_45377,N_45183);
and U47937 (N_47937,N_47430,N_46876);
nand U47938 (N_47938,N_47330,N_45160);
nor U47939 (N_47939,N_45096,N_46839);
nor U47940 (N_47940,N_45937,N_46783);
and U47941 (N_47941,N_45604,N_45131);
xnor U47942 (N_47942,N_45426,N_46220);
xnor U47943 (N_47943,N_46535,N_47008);
nor U47944 (N_47944,N_46565,N_46686);
xor U47945 (N_47945,N_45065,N_46500);
nand U47946 (N_47946,N_45858,N_46533);
and U47947 (N_47947,N_45999,N_47191);
xnor U47948 (N_47948,N_45221,N_46877);
or U47949 (N_47949,N_46917,N_46382);
xnor U47950 (N_47950,N_47359,N_46508);
or U47951 (N_47951,N_45370,N_45158);
nand U47952 (N_47952,N_47136,N_45961);
and U47953 (N_47953,N_46708,N_46957);
xnor U47954 (N_47954,N_45572,N_46673);
or U47955 (N_47955,N_46437,N_46807);
nor U47956 (N_47956,N_46003,N_45583);
nor U47957 (N_47957,N_46340,N_45638);
and U47958 (N_47958,N_46095,N_45384);
and U47959 (N_47959,N_46551,N_45711);
and U47960 (N_47960,N_46511,N_46940);
and U47961 (N_47961,N_46585,N_45835);
xnor U47962 (N_47962,N_47397,N_45058);
nand U47963 (N_47963,N_46892,N_45055);
or U47964 (N_47964,N_46345,N_46159);
xor U47965 (N_47965,N_47139,N_45134);
nor U47966 (N_47966,N_45556,N_46605);
nand U47967 (N_47967,N_46988,N_46756);
nor U47968 (N_47968,N_46318,N_45738);
or U47969 (N_47969,N_46005,N_47132);
or U47970 (N_47970,N_46894,N_45709);
nor U47971 (N_47971,N_45874,N_47113);
or U47972 (N_47972,N_46354,N_45765);
nor U47973 (N_47973,N_46815,N_46666);
or U47974 (N_47974,N_47072,N_46134);
or U47975 (N_47975,N_45652,N_47418);
nor U47976 (N_47976,N_45732,N_45863);
nor U47977 (N_47977,N_45566,N_45913);
nor U47978 (N_47978,N_46593,N_47076);
nor U47979 (N_47979,N_46113,N_46743);
and U47980 (N_47980,N_45230,N_46914);
and U47981 (N_47981,N_46135,N_45486);
nor U47982 (N_47982,N_46932,N_46758);
or U47983 (N_47983,N_45334,N_45060);
and U47984 (N_47984,N_46702,N_46543);
and U47985 (N_47985,N_45775,N_47269);
nand U47986 (N_47986,N_47234,N_47396);
nor U47987 (N_47987,N_46842,N_46503);
xnor U47988 (N_47988,N_46130,N_45630);
nor U47989 (N_47989,N_47295,N_45421);
nor U47990 (N_47990,N_45087,N_46173);
nor U47991 (N_47991,N_46030,N_47489);
and U47992 (N_47992,N_45692,N_46915);
and U47993 (N_47993,N_46305,N_45888);
or U47994 (N_47994,N_46896,N_47086);
nor U47995 (N_47995,N_45815,N_46614);
and U47996 (N_47996,N_46558,N_46426);
xor U47997 (N_47997,N_45243,N_45614);
or U47998 (N_47998,N_45276,N_45753);
nand U47999 (N_47999,N_47104,N_45419);
nand U48000 (N_48000,N_46233,N_46466);
nor U48001 (N_48001,N_46782,N_45248);
and U48002 (N_48002,N_46361,N_46482);
nor U48003 (N_48003,N_46991,N_45229);
xnor U48004 (N_48004,N_46191,N_46468);
or U48005 (N_48005,N_47322,N_47294);
and U48006 (N_48006,N_47045,N_45088);
nor U48007 (N_48007,N_45331,N_45803);
nand U48008 (N_48008,N_45936,N_46065);
xnor U48009 (N_48009,N_45452,N_45755);
xnor U48010 (N_48010,N_46200,N_45062);
and U48011 (N_48011,N_46996,N_47034);
and U48012 (N_48012,N_45902,N_47195);
or U48013 (N_48013,N_47286,N_46035);
xnor U48014 (N_48014,N_45806,N_46827);
nor U48015 (N_48015,N_45319,N_46703);
or U48016 (N_48016,N_46388,N_45013);
nor U48017 (N_48017,N_45745,N_45621);
and U48018 (N_48018,N_45257,N_46561);
xor U48019 (N_48019,N_45371,N_47316);
or U48020 (N_48020,N_45192,N_45042);
and U48021 (N_48021,N_46860,N_46088);
and U48022 (N_48022,N_45436,N_46987);
xor U48023 (N_48023,N_45380,N_45897);
and U48024 (N_48024,N_45409,N_45411);
nand U48025 (N_48025,N_45517,N_45699);
or U48026 (N_48026,N_45011,N_46545);
or U48027 (N_48027,N_46657,N_45655);
or U48028 (N_48028,N_45114,N_46831);
xor U48029 (N_48029,N_45020,N_47388);
xnor U48030 (N_48030,N_45057,N_45653);
xnor U48031 (N_48031,N_47499,N_46008);
or U48032 (N_48032,N_45282,N_46600);
or U48033 (N_48033,N_45672,N_45871);
xor U48034 (N_48034,N_47287,N_45862);
and U48035 (N_48035,N_46713,N_45831);
and U48036 (N_48036,N_45595,N_45713);
and U48037 (N_48037,N_47426,N_47262);
nand U48038 (N_48038,N_45772,N_46695);
nor U48039 (N_48039,N_46051,N_46176);
or U48040 (N_48040,N_46736,N_47372);
nand U48041 (N_48041,N_45451,N_46298);
nand U48042 (N_48042,N_46243,N_45097);
and U48043 (N_48043,N_47123,N_47382);
or U48044 (N_48044,N_45654,N_46102);
and U48045 (N_48045,N_45565,N_46138);
nor U48046 (N_48046,N_46083,N_46747);
xor U48047 (N_48047,N_46328,N_45663);
xor U48048 (N_48048,N_46225,N_46323);
nor U48049 (N_48049,N_45320,N_46630);
nor U48050 (N_48050,N_47358,N_46380);
nand U48051 (N_48051,N_45928,N_46234);
nor U48052 (N_48052,N_45550,N_45667);
and U48053 (N_48053,N_47221,N_45499);
or U48054 (N_48054,N_46408,N_46266);
nor U48055 (N_48055,N_45866,N_47410);
and U48056 (N_48056,N_47089,N_46332);
nand U48057 (N_48057,N_47292,N_46608);
nor U48058 (N_48058,N_45916,N_45737);
nor U48059 (N_48059,N_45983,N_46609);
nor U48060 (N_48060,N_45106,N_45774);
and U48061 (N_48061,N_46555,N_47112);
xor U48062 (N_48062,N_46031,N_45019);
xor U48063 (N_48063,N_45193,N_46365);
or U48064 (N_48064,N_47492,N_47235);
xor U48065 (N_48065,N_46032,N_46705);
xnor U48066 (N_48066,N_47169,N_45133);
xnor U48067 (N_48067,N_46090,N_47064);
xor U48068 (N_48068,N_47020,N_47452);
and U48069 (N_48069,N_47260,N_46875);
nor U48070 (N_48070,N_45955,N_46084);
nor U48071 (N_48071,N_47477,N_47328);
xor U48072 (N_48072,N_46639,N_46820);
nor U48073 (N_48073,N_46050,N_45222);
nor U48074 (N_48074,N_45759,N_45198);
nand U48075 (N_48075,N_46268,N_47405);
or U48076 (N_48076,N_45481,N_47151);
nor U48077 (N_48077,N_45233,N_45568);
nor U48078 (N_48078,N_47056,N_46920);
nand U48079 (N_48079,N_46312,N_47108);
nor U48080 (N_48080,N_46393,N_46017);
nand U48081 (N_48081,N_45249,N_47357);
or U48082 (N_48082,N_45938,N_45701);
nor U48083 (N_48083,N_45464,N_46486);
or U48084 (N_48084,N_46854,N_45857);
or U48085 (N_48085,N_45793,N_45415);
nand U48086 (N_48086,N_46693,N_45355);
and U48087 (N_48087,N_45325,N_45631);
and U48088 (N_48088,N_46937,N_46647);
or U48089 (N_48089,N_47448,N_46490);
xnor U48090 (N_48090,N_46742,N_45639);
xnor U48091 (N_48091,N_46656,N_46660);
nand U48092 (N_48092,N_46245,N_45101);
nor U48093 (N_48093,N_47217,N_45809);
and U48094 (N_48094,N_46814,N_46240);
xor U48095 (N_48095,N_46745,N_46294);
nor U48096 (N_48096,N_47480,N_46671);
nor U48097 (N_48097,N_45822,N_45819);
and U48098 (N_48098,N_47098,N_45678);
or U48099 (N_48099,N_45056,N_45976);
or U48100 (N_48100,N_46633,N_45491);
xnor U48101 (N_48101,N_46315,N_46616);
nor U48102 (N_48102,N_45310,N_46788);
nor U48103 (N_48103,N_45242,N_46699);
xor U48104 (N_48104,N_47366,N_45140);
xnor U48105 (N_48105,N_47023,N_45551);
and U48106 (N_48106,N_46689,N_46506);
nand U48107 (N_48107,N_46804,N_47265);
nor U48108 (N_48108,N_46923,N_47420);
nor U48109 (N_48109,N_46018,N_45720);
xnor U48110 (N_48110,N_45157,N_46597);
xor U48111 (N_48111,N_47091,N_46852);
nor U48112 (N_48112,N_46677,N_45734);
nor U48113 (N_48113,N_46291,N_47174);
xor U48114 (N_48114,N_46087,N_45939);
xor U48115 (N_48115,N_45470,N_47083);
xnor U48116 (N_48116,N_46286,N_46527);
nand U48117 (N_48117,N_47140,N_45258);
nand U48118 (N_48118,N_45519,N_46053);
nor U48119 (N_48119,N_45640,N_45099);
or U48120 (N_48120,N_47373,N_45909);
or U48121 (N_48121,N_46603,N_46073);
nand U48122 (N_48122,N_45196,N_46464);
xnor U48123 (N_48123,N_46728,N_46452);
and U48124 (N_48124,N_46068,N_47162);
or U48125 (N_48125,N_45132,N_45165);
nand U48126 (N_48126,N_45361,N_46832);
or U48127 (N_48127,N_46904,N_46195);
and U48128 (N_48128,N_46682,N_46663);
or U48129 (N_48129,N_45174,N_46882);
xor U48130 (N_48130,N_46536,N_45789);
nand U48131 (N_48131,N_45778,N_45559);
or U48132 (N_48132,N_45289,N_45425);
or U48133 (N_48133,N_46411,N_47411);
nand U48134 (N_48134,N_46226,N_45115);
xnor U48135 (N_48135,N_45461,N_46953);
nor U48136 (N_48136,N_46667,N_45437);
nor U48137 (N_48137,N_45156,N_45172);
nand U48138 (N_48138,N_45761,N_45552);
xnor U48139 (N_48139,N_45389,N_46132);
xnor U48140 (N_48140,N_46653,N_46580);
and U48141 (N_48141,N_46733,N_45031);
or U48142 (N_48142,N_46395,N_45527);
xnor U48143 (N_48143,N_45912,N_46218);
or U48144 (N_48144,N_46491,N_45767);
and U48145 (N_48145,N_45705,N_47279);
nor U48146 (N_48146,N_45040,N_45085);
and U48147 (N_48147,N_46934,N_46753);
or U48148 (N_48148,N_46515,N_46433);
and U48149 (N_48149,N_46759,N_46651);
xnor U48150 (N_48150,N_47173,N_46777);
or U48151 (N_48151,N_46679,N_45352);
nor U48152 (N_48152,N_46918,N_45358);
xnor U48153 (N_48153,N_45417,N_45922);
and U48154 (N_48154,N_45478,N_47347);
and U48155 (N_48155,N_46078,N_46339);
or U48156 (N_48156,N_45981,N_47090);
nand U48157 (N_48157,N_45602,N_45312);
nand U48158 (N_48158,N_45080,N_46692);
nand U48159 (N_48159,N_45538,N_47458);
and U48160 (N_48160,N_45284,N_46648);
and U48161 (N_48161,N_46394,N_45624);
xor U48162 (N_48162,N_46640,N_47129);
nor U48163 (N_48163,N_46441,N_46209);
and U48164 (N_48164,N_46369,N_45010);
or U48165 (N_48165,N_45714,N_46935);
nor U48166 (N_48166,N_46213,N_47380);
nand U48167 (N_48167,N_46712,N_45333);
nand U48168 (N_48168,N_46009,N_46162);
xor U48169 (N_48169,N_47318,N_47178);
or U48170 (N_48170,N_46771,N_46836);
nor U48171 (N_48171,N_45643,N_46750);
and U48172 (N_48172,N_46604,N_46390);
nand U48173 (N_48173,N_46865,N_46186);
or U48174 (N_48174,N_47062,N_45799);
nor U48175 (N_48175,N_47290,N_45079);
or U48176 (N_48176,N_45175,N_46252);
nand U48177 (N_48177,N_47446,N_47326);
or U48178 (N_48178,N_45051,N_46112);
nor U48179 (N_48179,N_45855,N_46454);
xor U48180 (N_48180,N_46576,N_46906);
nor U48181 (N_48181,N_46473,N_45546);
xor U48182 (N_48182,N_46510,N_47063);
xor U48183 (N_48183,N_45275,N_46120);
nor U48184 (N_48184,N_46281,N_46097);
and U48185 (N_48185,N_45408,N_46636);
nor U48186 (N_48186,N_46885,N_47319);
nor U48187 (N_48187,N_45919,N_46350);
xor U48188 (N_48188,N_45480,N_46080);
and U48189 (N_48189,N_45190,N_46307);
and U48190 (N_48190,N_45712,N_45986);
nand U48191 (N_48191,N_46858,N_45664);
nor U48192 (N_48192,N_46564,N_47375);
nand U48193 (N_48193,N_45254,N_47100);
or U48194 (N_48194,N_46407,N_46013);
or U48195 (N_48195,N_47441,N_45444);
xor U48196 (N_48196,N_45646,N_45135);
and U48197 (N_48197,N_46198,N_46769);
and U48198 (N_48198,N_45771,N_47252);
nor U48199 (N_48199,N_45210,N_47004);
nor U48200 (N_48200,N_45571,N_47152);
xor U48201 (N_48201,N_45514,N_46373);
and U48202 (N_48202,N_46694,N_45762);
and U48203 (N_48203,N_46881,N_47243);
xnor U48204 (N_48204,N_46058,N_46975);
or U48205 (N_48205,N_46295,N_45186);
nand U48206 (N_48206,N_45660,N_45914);
xor U48207 (N_48207,N_46485,N_46595);
or U48208 (N_48208,N_45128,N_46532);
nand U48209 (N_48209,N_45447,N_45689);
xor U48210 (N_48210,N_46516,N_45735);
and U48211 (N_48211,N_45609,N_46971);
xor U48212 (N_48212,N_46562,N_46982);
nor U48213 (N_48213,N_47001,N_47128);
nand U48214 (N_48214,N_45212,N_47042);
nand U48215 (N_48215,N_46143,N_45077);
or U48216 (N_48216,N_45879,N_46412);
or U48217 (N_48217,N_46726,N_46036);
or U48218 (N_48218,N_45659,N_45154);
or U48219 (N_48219,N_46992,N_46951);
nor U48220 (N_48220,N_45402,N_46577);
nor U48221 (N_48221,N_45523,N_45541);
nand U48222 (N_48222,N_46027,N_46546);
xor U48223 (N_48223,N_45834,N_46641);
and U48224 (N_48224,N_45111,N_46272);
nor U48225 (N_48225,N_46583,N_45786);
or U48226 (N_48226,N_45066,N_45524);
or U48227 (N_48227,N_45307,N_45449);
and U48228 (N_48228,N_45420,N_45203);
nand U48229 (N_48229,N_46208,N_46368);
or U48230 (N_48230,N_46121,N_46007);
xnor U48231 (N_48231,N_45668,N_46300);
and U48232 (N_48232,N_45367,N_45083);
or U48233 (N_48233,N_45053,N_45854);
nor U48234 (N_48234,N_46379,N_47214);
xor U48235 (N_48235,N_47147,N_47109);
nand U48236 (N_48236,N_47135,N_47493);
nand U48237 (N_48237,N_45608,N_45177);
nand U48238 (N_48238,N_46487,N_45368);
or U48239 (N_48239,N_45110,N_45529);
nor U48240 (N_48240,N_46055,N_45090);
xor U48241 (N_48241,N_45247,N_47368);
or U48242 (N_48242,N_47102,N_45899);
xnor U48243 (N_48243,N_46645,N_47096);
nor U48244 (N_48244,N_45509,N_46715);
nand U48245 (N_48245,N_46066,N_45393);
nor U48246 (N_48246,N_45400,N_47094);
nor U48247 (N_48247,N_45820,N_46596);
or U48248 (N_48248,N_47407,N_45875);
or U48249 (N_48249,N_46729,N_47482);
or U48250 (N_48250,N_46880,N_46911);
nor U48251 (N_48251,N_45033,N_46141);
nor U48252 (N_48252,N_45326,N_45757);
nor U48253 (N_48253,N_46662,N_46629);
and U48254 (N_48254,N_46000,N_45440);
xor U48255 (N_48255,N_45081,N_46631);
and U48256 (N_48256,N_45234,N_46416);
and U48257 (N_48257,N_47057,N_45148);
nand U48258 (N_48258,N_46443,N_46930);
nand U48259 (N_48259,N_45836,N_45856);
nor U48260 (N_48260,N_47451,N_46290);
or U48261 (N_48261,N_46067,N_45808);
nor U48262 (N_48262,N_45360,N_45615);
and U48263 (N_48263,N_46476,N_46994);
or U48264 (N_48264,N_46255,N_45238);
or U48265 (N_48265,N_45847,N_46045);
xnor U48266 (N_48266,N_45543,N_46939);
xnor U48267 (N_48267,N_45225,N_46737);
nand U48268 (N_48268,N_45122,N_46338);
nor U48269 (N_48269,N_47428,N_46232);
nor U48270 (N_48270,N_45300,N_46478);
nor U48271 (N_48271,N_47172,N_45261);
and U48272 (N_48272,N_47079,N_46878);
and U48273 (N_48273,N_46519,N_45840);
nor U48274 (N_48274,N_47257,N_46172);
nand U48275 (N_48275,N_45599,N_45763);
nand U48276 (N_48276,N_46552,N_47391);
nor U48277 (N_48277,N_45205,N_45184);
xor U48278 (N_48278,N_47200,N_45837);
and U48279 (N_48279,N_45064,N_46431);
or U48280 (N_48280,N_46231,N_45980);
xor U48281 (N_48281,N_46998,N_46969);
or U48282 (N_48282,N_45944,N_46962);
nand U48283 (N_48283,N_46931,N_47363);
nand U48284 (N_48284,N_45246,N_47283);
and U48285 (N_48285,N_45880,N_47404);
nand U48286 (N_48286,N_45266,N_46471);
nor U48287 (N_48287,N_45773,N_45490);
and U48288 (N_48288,N_46320,N_45314);
nand U48289 (N_48289,N_46124,N_45108);
xnor U48290 (N_48290,N_46428,N_45777);
or U48291 (N_48291,N_47434,N_46502);
or U48292 (N_48292,N_45994,N_46351);
xor U48293 (N_48293,N_47082,N_45910);
nand U48294 (N_48294,N_45542,N_46664);
nor U48295 (N_48295,N_46106,N_45232);
or U48296 (N_48296,N_47186,N_46963);
and U48297 (N_48297,N_46222,N_45316);
or U48298 (N_48298,N_45810,N_46069);
nor U48299 (N_48299,N_46374,N_46375);
and U48300 (N_48300,N_47171,N_45024);
or U48301 (N_48301,N_45137,N_46376);
or U48302 (N_48302,N_46722,N_45185);
nand U48303 (N_48303,N_45005,N_46463);
xnor U48304 (N_48304,N_46612,N_46105);
nor U48305 (N_48305,N_46474,N_45231);
nor U48306 (N_48306,N_47341,N_47253);
and U48307 (N_48307,N_45113,N_45748);
or U48308 (N_48308,N_45917,N_46672);
nand U48309 (N_48309,N_46046,N_45301);
and U48310 (N_48310,N_47439,N_46136);
nor U48311 (N_48311,N_47419,N_45159);
nor U48312 (N_48312,N_46203,N_45500);
nand U48313 (N_48313,N_46042,N_45164);
nor U48314 (N_48314,N_45522,N_46148);
xnor U48315 (N_48315,N_46383,N_47099);
xor U48316 (N_48316,N_46732,N_45677);
xor U48317 (N_48317,N_47187,N_47313);
and U48318 (N_48318,N_45518,N_47468);
nand U48319 (N_48319,N_47256,N_45891);
or U48320 (N_48320,N_45351,N_47469);
xnor U48321 (N_48321,N_47144,N_46079);
and U48322 (N_48322,N_46714,N_45941);
xnor U48323 (N_48323,N_47301,N_47154);
or U48324 (N_48324,N_47175,N_45650);
or U48325 (N_48325,N_46377,N_45220);
or U48326 (N_48326,N_46188,N_47101);
nor U48327 (N_48327,N_47227,N_47425);
nor U48328 (N_48328,N_46410,N_46805);
xor U48329 (N_48329,N_46085,N_46973);
xor U48330 (N_48330,N_46256,N_45093);
or U48331 (N_48331,N_45283,N_47060);
xnor U48332 (N_48332,N_46624,N_47006);
nand U48333 (N_48333,N_46219,N_46449);
and U48334 (N_48334,N_46033,N_46751);
and U48335 (N_48335,N_47157,N_45558);
xnor U48336 (N_48336,N_45208,N_46900);
nor U48337 (N_48337,N_45357,N_47192);
nor U48338 (N_48338,N_45236,N_45612);
nor U48339 (N_48339,N_46901,N_45277);
and U48340 (N_48340,N_47497,N_47389);
nor U48341 (N_48341,N_45023,N_46161);
xnor U48342 (N_48342,N_46738,N_47456);
nand U48343 (N_48343,N_46465,N_47305);
and U48344 (N_48344,N_47002,N_45387);
or U48345 (N_48345,N_46887,N_47338);
or U48346 (N_48346,N_45433,N_45784);
and U48347 (N_48347,N_46399,N_46496);
nand U48348 (N_48348,N_47444,N_46540);
xor U48349 (N_48349,N_45098,N_46179);
or U48350 (N_48350,N_45627,N_46993);
xor U48351 (N_48351,N_46592,N_45303);
nor U48352 (N_48352,N_45967,N_45070);
nor U48353 (N_48353,N_45790,N_47078);
xor U48354 (N_48354,N_45526,N_46248);
nor U48355 (N_48355,N_47142,N_45873);
nor U48356 (N_48356,N_46619,N_45504);
and U48357 (N_48357,N_45513,N_46980);
nand U48358 (N_48358,N_46623,N_46821);
nor U48359 (N_48359,N_45751,N_47403);
and U48360 (N_48360,N_45684,N_45562);
xor U48361 (N_48361,N_46943,N_47349);
nor U48362 (N_48362,N_46762,N_46778);
nand U48363 (N_48363,N_46260,N_45323);
or U48364 (N_48364,N_45706,N_47364);
or U48365 (N_48365,N_45830,N_46826);
nor U48366 (N_48366,N_46518,N_45207);
xor U48367 (N_48367,N_45227,N_47285);
nand U48368 (N_48368,N_47168,N_46154);
or U48369 (N_48369,N_46363,N_45045);
xnor U48370 (N_48370,N_47054,N_45818);
nor U48371 (N_48371,N_47118,N_45474);
nand U48372 (N_48372,N_47024,N_46869);
or U48373 (N_48373,N_45658,N_45851);
nor U48374 (N_48374,N_45308,N_45006);
and U48375 (N_48375,N_47258,N_45698);
nor U48376 (N_48376,N_45063,N_47437);
nand U48377 (N_48377,N_45406,N_45405);
xor U48378 (N_48378,N_46414,N_47259);
and U48379 (N_48379,N_46169,N_46093);
nor U48380 (N_48380,N_46092,N_46309);
or U48381 (N_48381,N_46716,N_46928);
nand U48382 (N_48382,N_45992,N_46438);
xnor U48383 (N_48383,N_45895,N_47381);
nor U48384 (N_48384,N_46822,N_46793);
nand U48385 (N_48385,N_46052,N_45861);
or U48386 (N_48386,N_47051,N_45034);
nand U48387 (N_48387,N_45346,N_46258);
and U48388 (N_48388,N_45483,N_45262);
or U48389 (N_48389,N_46765,N_47340);
nor U48390 (N_48390,N_47010,N_46803);
nand U48391 (N_48391,N_46406,N_47333);
nand U48392 (N_48392,N_47000,N_47219);
nor U48393 (N_48393,N_45575,N_46607);
nand U48394 (N_48394,N_47303,N_45469);
and U48395 (N_48395,N_46359,N_45446);
xnor U48396 (N_48396,N_45739,N_45674);
or U48397 (N_48397,N_46436,N_45445);
or U48398 (N_48398,N_45442,N_46781);
or U48399 (N_48399,N_46091,N_46448);
and U48400 (N_48400,N_46444,N_45721);
nand U48401 (N_48401,N_46296,N_46371);
xor U48402 (N_48402,N_45675,N_47130);
nor U48403 (N_48403,N_47120,N_45683);
nand U48404 (N_48404,N_46710,N_45318);
xor U48405 (N_48405,N_45901,N_45988);
or U48406 (N_48406,N_45485,N_45591);
nand U48407 (N_48407,N_47457,N_46709);
or U48408 (N_48408,N_45785,N_45567);
xnor U48409 (N_48409,N_45260,N_45691);
nor U48410 (N_48410,N_45904,N_46856);
nand U48411 (N_48411,N_47424,N_45180);
or U48412 (N_48412,N_47384,N_45251);
or U48413 (N_48413,N_45455,N_45915);
xor U48414 (N_48414,N_45244,N_46936);
and U48415 (N_48415,N_45487,N_45392);
xor U48416 (N_48416,N_46289,N_46870);
nor U48417 (N_48417,N_45703,N_46204);
xnor U48418 (N_48418,N_46655,N_45696);
xor U48419 (N_48419,N_46888,N_47415);
nor U48420 (N_48420,N_45321,N_47198);
nor U48421 (N_48421,N_46889,N_47071);
or U48422 (N_48422,N_45531,N_46586);
nand U48423 (N_48423,N_46160,N_46735);
and U48424 (N_48424,N_45561,N_47460);
xor U48425 (N_48425,N_47069,N_46770);
nor U48426 (N_48426,N_46984,N_45404);
xor U48427 (N_48427,N_45964,N_46025);
xor U48428 (N_48428,N_46507,N_46754);
nor U48429 (N_48429,N_47261,N_46871);
xnor U48430 (N_48430,N_45395,N_45001);
nand U48431 (N_48431,N_46990,N_47016);
and U48432 (N_48432,N_47194,N_45279);
and U48433 (N_48433,N_45864,N_46271);
or U48434 (N_48434,N_46779,N_45827);
xnor U48435 (N_48435,N_46370,N_46326);
nor U48436 (N_48436,N_47074,N_46461);
nor U48437 (N_48437,N_46074,N_45676);
nand U48438 (N_48438,N_46420,N_47414);
nand U48439 (N_48439,N_46446,N_45585);
xnor U48440 (N_48440,N_45194,N_45844);
nor U48441 (N_48441,N_45553,N_47255);
nand U48442 (N_48442,N_47416,N_45337);
or U48443 (N_48443,N_45796,N_45199);
nor U48444 (N_48444,N_45189,N_45957);
xor U48445 (N_48445,N_46652,N_47244);
nor U48446 (N_48446,N_47196,N_46479);
nor U48447 (N_48447,N_45311,N_45883);
and U48448 (N_48448,N_46445,N_47378);
nor U48449 (N_48449,N_45291,N_46866);
and U48450 (N_48450,N_47367,N_45539);
and U48451 (N_48451,N_46210,N_46504);
or U48452 (N_48452,N_47224,N_46850);
and U48453 (N_48453,N_45354,N_47205);
nand U48454 (N_48454,N_45733,N_46423);
nand U48455 (N_48455,N_46182,N_45671);
nand U48456 (N_48456,N_46140,N_45237);
and U48457 (N_48457,N_45996,N_45501);
xnor U48458 (N_48458,N_46740,N_45656);
or U48459 (N_48459,N_45061,N_47199);
nand U48460 (N_48460,N_46649,N_47225);
or U48461 (N_48461,N_46611,N_47475);
and U48462 (N_48462,N_47222,N_46525);
or U48463 (N_48463,N_46034,N_46685);
xnor U48464 (N_48464,N_46926,N_46288);
or U48465 (N_48465,N_47040,N_46206);
xnor U48466 (N_48466,N_46895,N_46459);
nor U48467 (N_48467,N_45954,N_46153);
nand U48468 (N_48468,N_46809,N_46467);
xnor U48469 (N_48469,N_47476,N_45929);
xor U48470 (N_48470,N_45823,N_45722);
nor U48471 (N_48471,N_47145,N_46983);
nand U48472 (N_48472,N_47332,N_46316);
or U48473 (N_48473,N_47447,N_45496);
nand U48474 (N_48474,N_47052,N_47267);
or U48475 (N_48475,N_46986,N_46589);
or U48476 (N_48476,N_45214,N_46321);
or U48477 (N_48477,N_47106,N_45412);
xor U48478 (N_48478,N_47036,N_47465);
nor U48479 (N_48479,N_45027,N_46114);
and U48480 (N_48480,N_46127,N_45213);
or U48481 (N_48481,N_46303,N_45838);
nor U48482 (N_48482,N_47012,N_46522);
nor U48483 (N_48483,N_46400,N_45870);
or U48484 (N_48484,N_45969,N_45032);
and U48485 (N_48485,N_45379,N_46107);
nand U48486 (N_48486,N_46811,N_45593);
and U48487 (N_48487,N_45685,N_46549);
or U48488 (N_48488,N_46039,N_47114);
and U48489 (N_48489,N_46096,N_46584);
or U48490 (N_48490,N_45030,N_47275);
xnor U48491 (N_48491,N_45103,N_47254);
xnor U48492 (N_48492,N_46669,N_45623);
nand U48493 (N_48493,N_45816,N_46659);
nand U48494 (N_48494,N_46853,N_47184);
nor U48495 (N_48495,N_45680,N_46274);
or U48496 (N_48496,N_45781,N_46537);
or U48497 (N_48497,N_45127,N_45434);
xor U48498 (N_48498,N_46797,N_47053);
nor U48499 (N_48499,N_45092,N_47179);
xor U48500 (N_48500,N_47080,N_46950);
nand U48501 (N_48501,N_46942,N_47310);
and U48502 (N_48502,N_46063,N_46185);
or U48503 (N_48503,N_45826,N_45573);
or U48504 (N_48504,N_46214,N_45105);
and U48505 (N_48505,N_47245,N_45118);
nand U48506 (N_48506,N_46460,N_46539);
and U48507 (N_48507,N_46979,N_45448);
and U48508 (N_48508,N_45339,N_46978);
or U48509 (N_48509,N_45993,N_46913);
or U48510 (N_48510,N_46292,N_46275);
nand U48511 (N_48511,N_47487,N_46304);
xnor U48512 (N_48512,N_46908,N_47273);
nand U48513 (N_48513,N_46456,N_45634);
xor U48514 (N_48514,N_47055,N_47193);
nor U48515 (N_48515,N_45817,N_46819);
nand U48516 (N_48516,N_47377,N_46429);
nand U48517 (N_48517,N_45946,N_46285);
nand U48518 (N_48518,N_46329,N_45697);
or U48519 (N_48519,N_45044,N_47181);
nand U48520 (N_48520,N_46696,N_46075);
xnor U48521 (N_48521,N_45084,N_46977);
or U48522 (N_48522,N_45832,N_46635);
nor U48523 (N_48523,N_46483,N_46907);
nand U48524 (N_48524,N_47021,N_47309);
xor U48525 (N_48525,N_47473,N_47084);
or U48526 (N_48526,N_47494,N_45467);
xor U48527 (N_48527,N_46514,N_45173);
and U48528 (N_48528,N_46212,N_45107);
nand U48529 (N_48529,N_47156,N_47163);
nand U48530 (N_48530,N_46538,N_46828);
xor U48531 (N_48531,N_46721,N_45629);
nand U48532 (N_48532,N_45952,N_45740);
or U48533 (N_48533,N_45100,N_47047);
and U48534 (N_48534,N_46578,N_46730);
or U48535 (N_48535,N_45933,N_47342);
xor U48536 (N_48536,N_46764,N_46392);
nand U48537 (N_48537,N_45441,N_47048);
and U48538 (N_48538,N_47277,N_45877);
nand U48539 (N_48539,N_45009,N_46064);
xnor U48540 (N_48540,N_46118,N_46184);
and U48541 (N_48541,N_46131,N_46557);
or U48542 (N_48542,N_46270,N_46566);
or U48543 (N_48543,N_45166,N_45574);
xor U48544 (N_48544,N_45921,N_45687);
xor U48545 (N_48545,N_47077,N_45890);
nand U48546 (N_48546,N_45218,N_47278);
nor U48547 (N_48547,N_47343,N_47150);
nand U48548 (N_48548,N_46086,N_46117);
nor U48549 (N_48549,N_47455,N_45454);
xnor U48550 (N_48550,N_47394,N_47429);
nor U48551 (N_48551,N_46047,N_46706);
nand U48552 (N_48552,N_47017,N_46178);
or U48553 (N_48553,N_45601,N_45403);
or U48554 (N_48554,N_45906,N_45439);
xor U48555 (N_48555,N_45528,N_47166);
nor U48556 (N_48556,N_46104,N_47271);
nand U48557 (N_48557,N_45007,N_45940);
nor U48558 (N_48558,N_45649,N_46829);
nand U48559 (N_48559,N_47284,N_47014);
and U48560 (N_48560,N_45181,N_45187);
or U48561 (N_48561,N_45074,N_47374);
nand U48562 (N_48562,N_46780,N_45665);
nand U48563 (N_48563,N_45129,N_45718);
nand U48564 (N_48564,N_46299,N_46250);
nand U48565 (N_48565,N_47188,N_45167);
nor U48566 (N_48566,N_46207,N_45666);
xnor U48567 (N_48567,N_46530,N_46026);
xnor U48568 (N_48568,N_45960,N_45600);
and U48569 (N_48569,N_46626,N_45907);
and U48570 (N_48570,N_47354,N_45252);
or U48571 (N_48571,N_45073,N_46995);
and U48572 (N_48572,N_46216,N_46193);
nand U48573 (N_48573,N_45540,N_47033);
nor U48574 (N_48574,N_45268,N_47462);
or U48575 (N_48575,N_45112,N_46101);
nor U48576 (N_48576,N_47019,N_45597);
and U48577 (N_48577,N_46610,N_46859);
nor U48578 (N_48578,N_46598,N_45082);
nand U48579 (N_48579,N_45255,N_46356);
nor U48580 (N_48580,N_47232,N_46945);
and U48581 (N_48581,N_45399,N_45594);
nand U48582 (N_48582,N_45896,N_46746);
or U48583 (N_48583,N_45432,N_45972);
nand U48584 (N_48584,N_45814,N_45812);
or U48585 (N_48585,N_47009,N_46115);
nor U48586 (N_48586,N_45605,N_45059);
and U48587 (N_48587,N_47459,N_45245);
nor U48588 (N_48588,N_45123,N_46016);
xor U48589 (N_48589,N_47398,N_47314);
nor U48590 (N_48590,N_46147,N_46014);
and U48591 (N_48591,N_47299,N_46021);
or U48592 (N_48592,N_45577,N_45516);
nor U48593 (N_48593,N_45839,N_46469);
and U48594 (N_48594,N_45872,N_46175);
nand U48595 (N_48595,N_45589,N_47220);
xnor U48596 (N_48596,N_45476,N_46684);
or U48597 (N_48597,N_46089,N_47280);
nor U48598 (N_48598,N_46267,N_47386);
nor U48599 (N_48599,N_45965,N_46893);
xnor U48600 (N_48600,N_47461,N_46077);
nor U48601 (N_48601,N_46941,N_47110);
nand U48602 (N_48602,N_47371,N_45138);
nand U48603 (N_48603,N_45104,N_45029);
nand U48604 (N_48604,N_46059,N_46863);
nand U48605 (N_48605,N_47095,N_45934);
nor U48606 (N_48606,N_46493,N_45054);
and U48607 (N_48607,N_46813,N_45330);
and U48608 (N_48608,N_45842,N_45948);
nor U48609 (N_48609,N_46054,N_45533);
xnor U48610 (N_48610,N_45606,N_46357);
nor U48611 (N_48611,N_46109,N_45616);
and U48612 (N_48612,N_47003,N_46795);
nand U48613 (N_48613,N_45022,N_46571);
nand U48614 (N_48614,N_45613,N_46526);
nand U48615 (N_48615,N_47266,N_46346);
nor U48616 (N_48616,N_45920,N_47498);
and U48617 (N_48617,N_46922,N_45690);
or U48618 (N_48618,N_46798,N_45095);
and U48619 (N_48619,N_45488,N_45968);
xor U48620 (N_48620,N_46620,N_45014);
nor U48621 (N_48621,N_46387,N_46524);
or U48622 (N_48622,N_46833,N_46748);
nor U48623 (N_48623,N_46602,N_45427);
or U48624 (N_48624,N_47323,N_45521);
xor U48625 (N_48625,N_46707,N_45363);
and U48626 (N_48626,N_47131,N_47281);
or U48627 (N_48627,N_45905,N_47365);
nor U48628 (N_48628,N_46687,N_46319);
nor U48629 (N_48629,N_46242,N_45036);
or U48630 (N_48630,N_46997,N_46768);
xor U48631 (N_48631,N_46470,N_46358);
nor U48632 (N_48632,N_45003,N_45825);
nand U48633 (N_48633,N_47242,N_46262);
nor U48634 (N_48634,N_47344,N_45136);
or U48635 (N_48635,N_46237,N_46308);
and U48636 (N_48636,N_45557,N_45002);
and U48637 (N_48637,N_47115,N_46786);
or U48638 (N_48638,N_46378,N_46253);
nor U48639 (N_48639,N_46489,N_46517);
and U48640 (N_48640,N_45362,N_47412);
xor U48641 (N_48641,N_46791,N_47207);
xor U48642 (N_48642,N_45884,N_46462);
nor U48643 (N_48643,N_45900,N_46628);
and U48644 (N_48644,N_45776,N_46621);
nand U48645 (N_48645,N_47432,N_45239);
nand U48646 (N_48646,N_45017,N_45046);
nand U48647 (N_48647,N_46529,N_47463);
or U48648 (N_48648,N_46279,N_45381);
nor U48649 (N_48649,N_46164,N_45710);
nor U48650 (N_48650,N_45067,N_47125);
and U48651 (N_48651,N_46802,N_46723);
xor U48652 (N_48652,N_46952,N_45534);
nand U48653 (N_48653,N_45892,N_45506);
xnor U48654 (N_48654,N_46110,N_46367);
nand U48655 (N_48655,N_47442,N_45622);
xor U48656 (N_48656,N_47491,N_45633);
or U48657 (N_48657,N_45750,N_45494);
or U48658 (N_48658,N_46151,N_47177);
nand U48659 (N_48659,N_45162,N_47296);
or U48660 (N_48660,N_45139,N_46948);
xnor U48661 (N_48661,N_46413,N_45076);
nor U48662 (N_48662,N_45848,N_46553);
or U48663 (N_48663,N_47208,N_46497);
xnor U48664 (N_48664,N_46835,N_45191);
nor U48665 (N_48665,N_46229,N_46848);
or U48666 (N_48666,N_45549,N_46642);
nor U48667 (N_48667,N_47189,N_47346);
or U48668 (N_48668,N_47107,N_46720);
nor U48669 (N_48669,N_45396,N_45179);
nand U48670 (N_48670,N_47417,N_46749);
xnor U48671 (N_48671,N_46972,N_45075);
or U48672 (N_48672,N_45302,N_46044);
and U48673 (N_48673,N_47408,N_47248);
nand U48674 (N_48674,N_47170,N_46806);
xnor U48675 (N_48675,N_47321,N_47361);
and U48676 (N_48676,N_46766,N_46152);
or U48677 (N_48677,N_45564,N_45369);
nand U48678 (N_48678,N_45431,N_45299);
and U48679 (N_48679,N_46767,N_45578);
or U48680 (N_48680,N_46313,N_45000);
nand U48681 (N_48681,N_47291,N_47312);
xnor U48682 (N_48682,N_46205,N_45116);
xor U48683 (N_48683,N_45841,N_47485);
and U48684 (N_48684,N_45304,N_46513);
nor U48685 (N_48685,N_45294,N_46643);
xor U48686 (N_48686,N_47488,N_46817);
nor U48687 (N_48687,N_46618,N_46103);
and U48688 (N_48688,N_45374,N_46480);
xor U48689 (N_48689,N_45700,N_45479);
nand U48690 (N_48690,N_46145,N_45438);
or U48691 (N_48691,N_46550,N_45783);
nor U48692 (N_48692,N_46451,N_45979);
or U48693 (N_48693,N_46700,N_46170);
nand U48694 (N_48694,N_46230,N_46897);
or U48695 (N_48695,N_47165,N_45219);
xor U48696 (N_48696,N_46698,N_45974);
and U48697 (N_48697,N_45923,N_46276);
nand U48698 (N_48698,N_46499,N_47383);
or U48699 (N_48699,N_46010,N_46194);
or U48700 (N_48700,N_47185,N_45224);
nor U48701 (N_48701,N_46534,N_47495);
nand U48702 (N_48702,N_46960,N_45547);
xnor U48703 (N_48703,N_47058,N_46818);
nand U48704 (N_48704,N_47304,N_45579);
xnor U48705 (N_48705,N_45443,N_46559);
nand U48706 (N_48706,N_45970,N_45918);
or U48707 (N_48707,N_47206,N_46284);
and U48708 (N_48708,N_46202,N_47158);
and U48709 (N_48709,N_45471,N_46327);
nor U48710 (N_48710,N_45430,N_47422);
or U48711 (N_48711,N_46912,N_47251);
xor U48712 (N_48712,N_46632,N_46238);
xnor U48713 (N_48713,N_45651,N_45263);
or U48714 (N_48714,N_46224,N_46157);
nand U48715 (N_48715,N_46638,N_45288);
or U48716 (N_48716,N_45147,N_46028);
nand U48717 (N_48717,N_47088,N_47127);
xor U48718 (N_48718,N_47435,N_47093);
and U48719 (N_48719,N_45385,N_47153);
nand U48720 (N_48720,N_47228,N_46341);
or U48721 (N_48721,N_45145,N_45724);
nor U48722 (N_48722,N_45532,N_45824);
or U48723 (N_48723,N_46415,N_45694);
nor U48724 (N_48724,N_45309,N_45867);
nand U48725 (N_48725,N_45144,N_46784);
nand U48726 (N_48726,N_45150,N_47050);
nor U48727 (N_48727,N_46146,N_46056);
or U48728 (N_48728,N_45341,N_46938);
nor U48729 (N_48729,N_47481,N_45209);
nor U48730 (N_48730,N_46792,N_45795);
xnor U48731 (N_48731,N_47164,N_47037);
and U48732 (N_48732,N_46100,N_45926);
xor U48733 (N_48733,N_46403,N_46650);
nor U48734 (N_48734,N_45293,N_45041);
nand U48735 (N_48735,N_46342,N_46425);
and U48736 (N_48736,N_46884,N_47311);
nor U48737 (N_48737,N_45378,N_47306);
or U48738 (N_48738,N_47015,N_45555);
or U48739 (N_48739,N_46845,N_46129);
and U48740 (N_48740,N_45429,N_45828);
or U48741 (N_48741,N_45305,N_45256);
nor U48742 (N_48742,N_45766,N_45582);
nand U48743 (N_48743,N_45025,N_45978);
or U48744 (N_48744,N_45971,N_45510);
nor U48745 (N_48745,N_47236,N_47406);
nor U48746 (N_48746,N_46867,N_46076);
and U48747 (N_48747,N_45846,N_45728);
or U48748 (N_48748,N_45520,N_46494);
or U48749 (N_48749,N_47335,N_45715);
xor U48750 (N_48750,N_45800,N_45877);
nor U48751 (N_48751,N_45057,N_47178);
nor U48752 (N_48752,N_45153,N_45727);
nand U48753 (N_48753,N_46312,N_45349);
nand U48754 (N_48754,N_47193,N_45352);
and U48755 (N_48755,N_45691,N_45409);
nand U48756 (N_48756,N_45235,N_46506);
xnor U48757 (N_48757,N_46427,N_45610);
nand U48758 (N_48758,N_47207,N_45851);
xor U48759 (N_48759,N_46172,N_45198);
xnor U48760 (N_48760,N_46641,N_46042);
nor U48761 (N_48761,N_47461,N_46453);
nor U48762 (N_48762,N_45350,N_46678);
or U48763 (N_48763,N_45582,N_45825);
nand U48764 (N_48764,N_46807,N_46623);
nor U48765 (N_48765,N_45102,N_47200);
or U48766 (N_48766,N_47022,N_45541);
xnor U48767 (N_48767,N_46794,N_45446);
nor U48768 (N_48768,N_46603,N_47362);
xor U48769 (N_48769,N_46956,N_45261);
and U48770 (N_48770,N_45916,N_46652);
and U48771 (N_48771,N_45380,N_46411);
xnor U48772 (N_48772,N_45544,N_46159);
nand U48773 (N_48773,N_46788,N_47247);
or U48774 (N_48774,N_46782,N_45728);
nor U48775 (N_48775,N_47357,N_45723);
nor U48776 (N_48776,N_45539,N_46126);
nand U48777 (N_48777,N_45296,N_45450);
xor U48778 (N_48778,N_46153,N_46719);
and U48779 (N_48779,N_47171,N_45788);
and U48780 (N_48780,N_45065,N_46475);
nand U48781 (N_48781,N_45175,N_45097);
nor U48782 (N_48782,N_46836,N_47283);
nor U48783 (N_48783,N_47336,N_46189);
xnor U48784 (N_48784,N_45350,N_45821);
nand U48785 (N_48785,N_45003,N_45495);
or U48786 (N_48786,N_47396,N_46735);
nand U48787 (N_48787,N_46973,N_46762);
nand U48788 (N_48788,N_45878,N_46260);
or U48789 (N_48789,N_45978,N_45226);
or U48790 (N_48790,N_45866,N_47063);
or U48791 (N_48791,N_46906,N_46334);
nand U48792 (N_48792,N_46750,N_47499);
xor U48793 (N_48793,N_45291,N_47168);
nand U48794 (N_48794,N_46695,N_46326);
or U48795 (N_48795,N_45852,N_45594);
and U48796 (N_48796,N_46022,N_45592);
xor U48797 (N_48797,N_45177,N_45088);
nand U48798 (N_48798,N_46948,N_46618);
or U48799 (N_48799,N_46314,N_46421);
xor U48800 (N_48800,N_45992,N_46614);
and U48801 (N_48801,N_45805,N_45245);
nand U48802 (N_48802,N_46425,N_45683);
xor U48803 (N_48803,N_47451,N_46631);
nor U48804 (N_48804,N_45910,N_46557);
or U48805 (N_48805,N_46014,N_46030);
nand U48806 (N_48806,N_47008,N_45715);
and U48807 (N_48807,N_47081,N_46907);
or U48808 (N_48808,N_45533,N_47109);
nor U48809 (N_48809,N_47427,N_47240);
nor U48810 (N_48810,N_45544,N_46699);
xnor U48811 (N_48811,N_45297,N_45290);
nand U48812 (N_48812,N_46473,N_47103);
xnor U48813 (N_48813,N_46656,N_46799);
xor U48814 (N_48814,N_45658,N_45979);
nor U48815 (N_48815,N_47200,N_47283);
xor U48816 (N_48816,N_47115,N_46406);
nor U48817 (N_48817,N_45417,N_46423);
nor U48818 (N_48818,N_46031,N_45657);
or U48819 (N_48819,N_45340,N_46977);
xnor U48820 (N_48820,N_46581,N_46048);
nand U48821 (N_48821,N_47026,N_46825);
nand U48822 (N_48822,N_46211,N_45719);
nand U48823 (N_48823,N_45231,N_46955);
nor U48824 (N_48824,N_45733,N_46443);
or U48825 (N_48825,N_47490,N_46116);
nand U48826 (N_48826,N_45706,N_47256);
nor U48827 (N_48827,N_45406,N_46495);
xnor U48828 (N_48828,N_46633,N_47018);
or U48829 (N_48829,N_47448,N_46335);
and U48830 (N_48830,N_45721,N_46042);
or U48831 (N_48831,N_45298,N_45186);
and U48832 (N_48832,N_46562,N_46192);
nand U48833 (N_48833,N_46874,N_45516);
and U48834 (N_48834,N_47123,N_46573);
nand U48835 (N_48835,N_47094,N_47072);
and U48836 (N_48836,N_46950,N_46681);
nand U48837 (N_48837,N_45667,N_45987);
nor U48838 (N_48838,N_47100,N_47453);
nand U48839 (N_48839,N_46591,N_47100);
xnor U48840 (N_48840,N_45978,N_46843);
nand U48841 (N_48841,N_45370,N_46931);
xnor U48842 (N_48842,N_46713,N_46440);
nand U48843 (N_48843,N_46925,N_47401);
nor U48844 (N_48844,N_47430,N_46888);
or U48845 (N_48845,N_46907,N_46279);
xor U48846 (N_48846,N_45853,N_47344);
nand U48847 (N_48847,N_46001,N_47453);
or U48848 (N_48848,N_46630,N_47077);
or U48849 (N_48849,N_46152,N_46904);
nand U48850 (N_48850,N_47020,N_46555);
nor U48851 (N_48851,N_45998,N_46513);
xnor U48852 (N_48852,N_45671,N_47481);
or U48853 (N_48853,N_47335,N_45989);
xor U48854 (N_48854,N_46096,N_47291);
nor U48855 (N_48855,N_45230,N_46863);
nand U48856 (N_48856,N_46615,N_47326);
xnor U48857 (N_48857,N_45964,N_45211);
xor U48858 (N_48858,N_45724,N_45844);
and U48859 (N_48859,N_45611,N_45248);
or U48860 (N_48860,N_46079,N_47159);
or U48861 (N_48861,N_46132,N_47302);
nor U48862 (N_48862,N_47381,N_46036);
xnor U48863 (N_48863,N_47023,N_45133);
nor U48864 (N_48864,N_46758,N_45277);
nand U48865 (N_48865,N_46837,N_46695);
xor U48866 (N_48866,N_47232,N_45133);
and U48867 (N_48867,N_46064,N_45324);
nand U48868 (N_48868,N_46953,N_47232);
and U48869 (N_48869,N_46840,N_45856);
nand U48870 (N_48870,N_47124,N_45600);
xor U48871 (N_48871,N_46874,N_46466);
nor U48872 (N_48872,N_47235,N_46980);
nor U48873 (N_48873,N_45454,N_47161);
nor U48874 (N_48874,N_47457,N_46023);
or U48875 (N_48875,N_45136,N_46410);
xnor U48876 (N_48876,N_46315,N_45526);
nand U48877 (N_48877,N_47391,N_47196);
xnor U48878 (N_48878,N_45740,N_45598);
or U48879 (N_48879,N_46350,N_46646);
nor U48880 (N_48880,N_45064,N_47081);
xor U48881 (N_48881,N_46702,N_45193);
and U48882 (N_48882,N_45327,N_46813);
xor U48883 (N_48883,N_46493,N_46426);
nand U48884 (N_48884,N_45229,N_47188);
or U48885 (N_48885,N_45920,N_47368);
and U48886 (N_48886,N_47178,N_45137);
xor U48887 (N_48887,N_46593,N_45876);
xor U48888 (N_48888,N_46499,N_46635);
and U48889 (N_48889,N_46339,N_47341);
nand U48890 (N_48890,N_47150,N_46380);
nand U48891 (N_48891,N_45684,N_46741);
nand U48892 (N_48892,N_46824,N_46959);
nor U48893 (N_48893,N_47174,N_47262);
nor U48894 (N_48894,N_45675,N_47068);
nand U48895 (N_48895,N_45314,N_45102);
nand U48896 (N_48896,N_45222,N_46986);
nand U48897 (N_48897,N_45924,N_46994);
and U48898 (N_48898,N_45432,N_45656);
xnor U48899 (N_48899,N_46267,N_46165);
or U48900 (N_48900,N_46003,N_46254);
or U48901 (N_48901,N_46817,N_47100);
nor U48902 (N_48902,N_47499,N_45900);
xor U48903 (N_48903,N_45758,N_45055);
xor U48904 (N_48904,N_46854,N_45099);
nand U48905 (N_48905,N_45941,N_46909);
or U48906 (N_48906,N_47363,N_45004);
or U48907 (N_48907,N_45152,N_46049);
nand U48908 (N_48908,N_46494,N_46931);
xor U48909 (N_48909,N_45401,N_45017);
xor U48910 (N_48910,N_47174,N_45357);
or U48911 (N_48911,N_46708,N_45449);
or U48912 (N_48912,N_45616,N_46761);
xnor U48913 (N_48913,N_45078,N_46330);
nand U48914 (N_48914,N_45158,N_47472);
and U48915 (N_48915,N_45886,N_46235);
nor U48916 (N_48916,N_46428,N_47417);
xnor U48917 (N_48917,N_45989,N_46130);
nor U48918 (N_48918,N_45820,N_47188);
or U48919 (N_48919,N_46922,N_46189);
and U48920 (N_48920,N_47155,N_46673);
nand U48921 (N_48921,N_45290,N_47330);
nand U48922 (N_48922,N_46223,N_45254);
nand U48923 (N_48923,N_47136,N_46846);
or U48924 (N_48924,N_45524,N_46169);
nor U48925 (N_48925,N_45212,N_46761);
nor U48926 (N_48926,N_46698,N_46552);
nor U48927 (N_48927,N_46049,N_45225);
and U48928 (N_48928,N_45591,N_47221);
nand U48929 (N_48929,N_45368,N_46532);
nor U48930 (N_48930,N_45831,N_45476);
xnor U48931 (N_48931,N_45309,N_46173);
xnor U48932 (N_48932,N_45700,N_47456);
nand U48933 (N_48933,N_45354,N_46835);
nor U48934 (N_48934,N_45213,N_45797);
and U48935 (N_48935,N_47406,N_46455);
nor U48936 (N_48936,N_46745,N_45174);
nand U48937 (N_48937,N_45873,N_47145);
and U48938 (N_48938,N_46419,N_46082);
or U48939 (N_48939,N_46629,N_46323);
or U48940 (N_48940,N_46044,N_47450);
nand U48941 (N_48941,N_45850,N_46195);
nor U48942 (N_48942,N_45743,N_46129);
and U48943 (N_48943,N_46867,N_46381);
and U48944 (N_48944,N_47137,N_45251);
and U48945 (N_48945,N_45117,N_46531);
nand U48946 (N_48946,N_45370,N_45254);
or U48947 (N_48947,N_45090,N_46499);
xor U48948 (N_48948,N_45104,N_45341);
nand U48949 (N_48949,N_46775,N_45168);
or U48950 (N_48950,N_46644,N_46991);
and U48951 (N_48951,N_45301,N_45607);
xor U48952 (N_48952,N_45922,N_46279);
or U48953 (N_48953,N_45529,N_45273);
or U48954 (N_48954,N_45458,N_46698);
nor U48955 (N_48955,N_45094,N_45135);
nand U48956 (N_48956,N_46790,N_46205);
xor U48957 (N_48957,N_47344,N_45909);
nand U48958 (N_48958,N_45450,N_46078);
or U48959 (N_48959,N_46021,N_46239);
xor U48960 (N_48960,N_46334,N_45465);
and U48961 (N_48961,N_45121,N_46493);
nor U48962 (N_48962,N_47436,N_45502);
and U48963 (N_48963,N_46445,N_45695);
nand U48964 (N_48964,N_47068,N_46910);
nand U48965 (N_48965,N_46548,N_46866);
nand U48966 (N_48966,N_47331,N_45624);
nor U48967 (N_48967,N_45192,N_45748);
xnor U48968 (N_48968,N_45918,N_46252);
xor U48969 (N_48969,N_46406,N_46047);
nor U48970 (N_48970,N_47024,N_45414);
or U48971 (N_48971,N_46721,N_45814);
nand U48972 (N_48972,N_45453,N_47170);
or U48973 (N_48973,N_46307,N_45071);
nand U48974 (N_48974,N_45531,N_46087);
or U48975 (N_48975,N_45303,N_46342);
and U48976 (N_48976,N_47280,N_45719);
nor U48977 (N_48977,N_45409,N_46417);
or U48978 (N_48978,N_45571,N_45038);
or U48979 (N_48979,N_46909,N_46396);
nor U48980 (N_48980,N_45610,N_46076);
and U48981 (N_48981,N_46096,N_45344);
or U48982 (N_48982,N_45483,N_47440);
nand U48983 (N_48983,N_46165,N_45951);
xor U48984 (N_48984,N_45412,N_47313);
or U48985 (N_48985,N_46445,N_46304);
xor U48986 (N_48986,N_45560,N_46052);
nand U48987 (N_48987,N_45087,N_47023);
or U48988 (N_48988,N_46363,N_46994);
and U48989 (N_48989,N_46855,N_46183);
and U48990 (N_48990,N_47000,N_45695);
nand U48991 (N_48991,N_45721,N_46794);
or U48992 (N_48992,N_46942,N_45083);
or U48993 (N_48993,N_46455,N_45465);
or U48994 (N_48994,N_46977,N_46512);
xor U48995 (N_48995,N_46778,N_45545);
nand U48996 (N_48996,N_45303,N_45987);
xnor U48997 (N_48997,N_46652,N_47050);
nand U48998 (N_48998,N_46885,N_45848);
or U48999 (N_48999,N_45467,N_47029);
nor U49000 (N_49000,N_46867,N_45564);
xor U49001 (N_49001,N_46989,N_45940);
nor U49002 (N_49002,N_47293,N_45733);
xor U49003 (N_49003,N_45024,N_45436);
and U49004 (N_49004,N_47140,N_46710);
or U49005 (N_49005,N_45434,N_45419);
and U49006 (N_49006,N_45899,N_45616);
or U49007 (N_49007,N_46784,N_45297);
and U49008 (N_49008,N_45273,N_46400);
and U49009 (N_49009,N_47257,N_47102);
nand U49010 (N_49010,N_47054,N_45700);
nand U49011 (N_49011,N_47219,N_47044);
nor U49012 (N_49012,N_47185,N_47229);
or U49013 (N_49013,N_45104,N_45747);
nor U49014 (N_49014,N_46405,N_46598);
xor U49015 (N_49015,N_47140,N_46945);
and U49016 (N_49016,N_45742,N_47158);
nor U49017 (N_49017,N_47136,N_47063);
nor U49018 (N_49018,N_45436,N_45247);
and U49019 (N_49019,N_46901,N_45283);
or U49020 (N_49020,N_45946,N_47163);
and U49021 (N_49021,N_45327,N_45908);
and U49022 (N_49022,N_47380,N_46502);
nand U49023 (N_49023,N_46687,N_47045);
and U49024 (N_49024,N_45908,N_45310);
nand U49025 (N_49025,N_45105,N_45849);
nand U49026 (N_49026,N_45587,N_45212);
nor U49027 (N_49027,N_45261,N_47102);
nor U49028 (N_49028,N_45011,N_46623);
and U49029 (N_49029,N_47495,N_45586);
nand U49030 (N_49030,N_45130,N_46491);
or U49031 (N_49031,N_47479,N_46295);
nand U49032 (N_49032,N_45430,N_46216);
or U49033 (N_49033,N_46472,N_46304);
and U49034 (N_49034,N_45305,N_45987);
or U49035 (N_49035,N_45588,N_45697);
nor U49036 (N_49036,N_46213,N_45637);
xor U49037 (N_49037,N_45776,N_45330);
nor U49038 (N_49038,N_45984,N_45614);
nand U49039 (N_49039,N_47202,N_46266);
or U49040 (N_49040,N_46269,N_46331);
nor U49041 (N_49041,N_46146,N_46140);
nor U49042 (N_49042,N_47178,N_45298);
nor U49043 (N_49043,N_45771,N_47195);
xnor U49044 (N_49044,N_45659,N_45613);
xor U49045 (N_49045,N_45167,N_46658);
nor U49046 (N_49046,N_47464,N_47237);
nand U49047 (N_49047,N_46038,N_46568);
or U49048 (N_49048,N_47181,N_46416);
nor U49049 (N_49049,N_47380,N_47425);
or U49050 (N_49050,N_45592,N_45711);
nor U49051 (N_49051,N_45818,N_45543);
and U49052 (N_49052,N_45363,N_45438);
nor U49053 (N_49053,N_45636,N_45894);
or U49054 (N_49054,N_46464,N_46517);
xor U49055 (N_49055,N_47202,N_45239);
nand U49056 (N_49056,N_47398,N_45113);
or U49057 (N_49057,N_45393,N_45463);
nor U49058 (N_49058,N_45373,N_45517);
and U49059 (N_49059,N_46792,N_45292);
and U49060 (N_49060,N_47028,N_46148);
or U49061 (N_49061,N_46727,N_46868);
nand U49062 (N_49062,N_46262,N_46830);
nand U49063 (N_49063,N_46197,N_46263);
or U49064 (N_49064,N_46132,N_45371);
and U49065 (N_49065,N_46545,N_46854);
nand U49066 (N_49066,N_47026,N_46773);
and U49067 (N_49067,N_45316,N_46567);
nand U49068 (N_49068,N_45602,N_45738);
nor U49069 (N_49069,N_45770,N_47186);
or U49070 (N_49070,N_46539,N_45650);
or U49071 (N_49071,N_46273,N_46151);
xor U49072 (N_49072,N_45123,N_45659);
xnor U49073 (N_49073,N_45836,N_45347);
nand U49074 (N_49074,N_47206,N_46377);
xor U49075 (N_49075,N_46132,N_46506);
and U49076 (N_49076,N_46896,N_46406);
or U49077 (N_49077,N_46514,N_46292);
nor U49078 (N_49078,N_47250,N_46428);
nand U49079 (N_49079,N_47441,N_46229);
and U49080 (N_49080,N_47024,N_47133);
and U49081 (N_49081,N_46002,N_45248);
nand U49082 (N_49082,N_47003,N_46265);
or U49083 (N_49083,N_46300,N_46032);
xor U49084 (N_49084,N_45223,N_46701);
nand U49085 (N_49085,N_45984,N_47480);
nor U49086 (N_49086,N_46307,N_46163);
or U49087 (N_49087,N_45990,N_47407);
nand U49088 (N_49088,N_46166,N_47412);
nand U49089 (N_49089,N_47104,N_45070);
xnor U49090 (N_49090,N_46185,N_47262);
or U49091 (N_49091,N_46662,N_47409);
nand U49092 (N_49092,N_45221,N_47225);
nand U49093 (N_49093,N_47229,N_46494);
and U49094 (N_49094,N_47312,N_45291);
nand U49095 (N_49095,N_45533,N_45116);
xnor U49096 (N_49096,N_46975,N_45220);
nor U49097 (N_49097,N_45558,N_47028);
and U49098 (N_49098,N_46071,N_45072);
nor U49099 (N_49099,N_45246,N_46339);
nand U49100 (N_49100,N_45916,N_45179);
and U49101 (N_49101,N_45912,N_46806);
nand U49102 (N_49102,N_46791,N_46797);
xor U49103 (N_49103,N_45714,N_45732);
and U49104 (N_49104,N_46801,N_47390);
nand U49105 (N_49105,N_45899,N_46916);
nor U49106 (N_49106,N_45834,N_45331);
and U49107 (N_49107,N_45229,N_45868);
xnor U49108 (N_49108,N_45712,N_45305);
and U49109 (N_49109,N_46165,N_46289);
xnor U49110 (N_49110,N_45849,N_45156);
or U49111 (N_49111,N_45534,N_45161);
xnor U49112 (N_49112,N_46979,N_45926);
nor U49113 (N_49113,N_46409,N_45411);
nor U49114 (N_49114,N_45970,N_45657);
xnor U49115 (N_49115,N_47474,N_46136);
and U49116 (N_49116,N_45043,N_45680);
and U49117 (N_49117,N_45626,N_45923);
xnor U49118 (N_49118,N_46046,N_45405);
nand U49119 (N_49119,N_47489,N_46923);
or U49120 (N_49120,N_45387,N_46939);
and U49121 (N_49121,N_46418,N_46660);
nand U49122 (N_49122,N_47141,N_45532);
and U49123 (N_49123,N_46964,N_45815);
nand U49124 (N_49124,N_45061,N_46676);
nor U49125 (N_49125,N_46291,N_46961);
nand U49126 (N_49126,N_45879,N_47135);
xnor U49127 (N_49127,N_46375,N_47001);
or U49128 (N_49128,N_46972,N_46192);
xor U49129 (N_49129,N_46147,N_45463);
and U49130 (N_49130,N_45823,N_45998);
nand U49131 (N_49131,N_46216,N_45140);
xor U49132 (N_49132,N_47164,N_46080);
xnor U49133 (N_49133,N_45716,N_46384);
nor U49134 (N_49134,N_45184,N_46562);
or U49135 (N_49135,N_47067,N_47172);
or U49136 (N_49136,N_45121,N_45830);
or U49137 (N_49137,N_45813,N_47369);
nand U49138 (N_49138,N_47335,N_45964);
and U49139 (N_49139,N_45121,N_47474);
nor U49140 (N_49140,N_46565,N_45736);
nor U49141 (N_49141,N_46795,N_45428);
and U49142 (N_49142,N_46424,N_45876);
xnor U49143 (N_49143,N_45729,N_45022);
nand U49144 (N_49144,N_45175,N_45421);
and U49145 (N_49145,N_45879,N_45678);
nor U49146 (N_49146,N_47179,N_46746);
nor U49147 (N_49147,N_46624,N_45682);
nor U49148 (N_49148,N_45473,N_45025);
xor U49149 (N_49149,N_47426,N_46057);
xnor U49150 (N_49150,N_46035,N_46568);
nor U49151 (N_49151,N_45476,N_47346);
nand U49152 (N_49152,N_46767,N_45059);
nand U49153 (N_49153,N_46154,N_45714);
nor U49154 (N_49154,N_45857,N_46209);
nand U49155 (N_49155,N_45289,N_46016);
nor U49156 (N_49156,N_46744,N_45694);
nor U49157 (N_49157,N_46266,N_46053);
nor U49158 (N_49158,N_45493,N_46576);
nor U49159 (N_49159,N_46969,N_45711);
xnor U49160 (N_49160,N_46740,N_45818);
nor U49161 (N_49161,N_47104,N_46109);
and U49162 (N_49162,N_45673,N_46730);
xnor U49163 (N_49163,N_47129,N_45591);
or U49164 (N_49164,N_47021,N_47335);
xnor U49165 (N_49165,N_46505,N_45906);
or U49166 (N_49166,N_46489,N_47443);
or U49167 (N_49167,N_45343,N_46310);
xor U49168 (N_49168,N_45363,N_45292);
nand U49169 (N_49169,N_46665,N_47051);
and U49170 (N_49170,N_46104,N_46346);
and U49171 (N_49171,N_45355,N_46162);
or U49172 (N_49172,N_46888,N_46831);
or U49173 (N_49173,N_46919,N_45809);
nor U49174 (N_49174,N_47368,N_46460);
nor U49175 (N_49175,N_45643,N_46837);
and U49176 (N_49176,N_45635,N_46325);
and U49177 (N_49177,N_45528,N_47221);
nor U49178 (N_49178,N_47005,N_45903);
nand U49179 (N_49179,N_47428,N_45794);
and U49180 (N_49180,N_45150,N_45568);
nand U49181 (N_49181,N_45047,N_46590);
and U49182 (N_49182,N_46195,N_46124);
nand U49183 (N_49183,N_46756,N_46802);
nand U49184 (N_49184,N_46652,N_45233);
nand U49185 (N_49185,N_46238,N_46319);
or U49186 (N_49186,N_46391,N_47197);
and U49187 (N_49187,N_45302,N_47126);
nor U49188 (N_49188,N_45039,N_46768);
nor U49189 (N_49189,N_47343,N_45402);
or U49190 (N_49190,N_47201,N_47177);
or U49191 (N_49191,N_47333,N_46783);
nand U49192 (N_49192,N_46710,N_45853);
nor U49193 (N_49193,N_45553,N_45772);
xor U49194 (N_49194,N_47264,N_46251);
nand U49195 (N_49195,N_47002,N_45993);
nand U49196 (N_49196,N_45053,N_45706);
and U49197 (N_49197,N_46274,N_45797);
and U49198 (N_49198,N_46772,N_45118);
nor U49199 (N_49199,N_45132,N_45239);
and U49200 (N_49200,N_46397,N_45039);
nor U49201 (N_49201,N_46003,N_47332);
nand U49202 (N_49202,N_47049,N_45508);
nor U49203 (N_49203,N_45090,N_45128);
xor U49204 (N_49204,N_46814,N_45639);
nand U49205 (N_49205,N_46009,N_46712);
nor U49206 (N_49206,N_46847,N_45370);
nor U49207 (N_49207,N_45970,N_45913);
or U49208 (N_49208,N_46407,N_46783);
xor U49209 (N_49209,N_47404,N_45373);
xor U49210 (N_49210,N_45283,N_46428);
nand U49211 (N_49211,N_45748,N_46937);
and U49212 (N_49212,N_46961,N_47428);
nor U49213 (N_49213,N_46009,N_47435);
or U49214 (N_49214,N_45110,N_45737);
nand U49215 (N_49215,N_46233,N_46053);
or U49216 (N_49216,N_46605,N_46050);
nor U49217 (N_49217,N_45006,N_46099);
or U49218 (N_49218,N_45841,N_46788);
or U49219 (N_49219,N_45506,N_46066);
xnor U49220 (N_49220,N_47411,N_46019);
or U49221 (N_49221,N_45096,N_46107);
nor U49222 (N_49222,N_45391,N_46643);
or U49223 (N_49223,N_45517,N_45575);
nor U49224 (N_49224,N_45550,N_46744);
nor U49225 (N_49225,N_45098,N_46362);
nand U49226 (N_49226,N_45498,N_45222);
xor U49227 (N_49227,N_46890,N_45643);
nand U49228 (N_49228,N_45063,N_45675);
nand U49229 (N_49229,N_46127,N_46549);
or U49230 (N_49230,N_46621,N_46085);
nand U49231 (N_49231,N_45118,N_46258);
nor U49232 (N_49232,N_45462,N_46005);
nor U49233 (N_49233,N_46285,N_45633);
and U49234 (N_49234,N_47431,N_45022);
xor U49235 (N_49235,N_46007,N_46048);
and U49236 (N_49236,N_47238,N_45097);
xor U49237 (N_49237,N_47119,N_46417);
xor U49238 (N_49238,N_45945,N_46680);
and U49239 (N_49239,N_47211,N_47104);
xor U49240 (N_49240,N_45037,N_47298);
nor U49241 (N_49241,N_45723,N_46817);
xor U49242 (N_49242,N_47457,N_46129);
or U49243 (N_49243,N_45627,N_45607);
and U49244 (N_49244,N_45364,N_47442);
xor U49245 (N_49245,N_45796,N_45996);
nor U49246 (N_49246,N_46076,N_46749);
xor U49247 (N_49247,N_47145,N_45206);
nor U49248 (N_49248,N_45151,N_45998);
nand U49249 (N_49249,N_45356,N_46378);
and U49250 (N_49250,N_46190,N_47139);
and U49251 (N_49251,N_45710,N_46510);
and U49252 (N_49252,N_46763,N_45970);
and U49253 (N_49253,N_45306,N_45116);
nor U49254 (N_49254,N_46697,N_47007);
xnor U49255 (N_49255,N_47337,N_47306);
nor U49256 (N_49256,N_47150,N_47152);
and U49257 (N_49257,N_45768,N_47079);
nor U49258 (N_49258,N_46529,N_47450);
and U49259 (N_49259,N_46429,N_47384);
nor U49260 (N_49260,N_45590,N_45262);
nand U49261 (N_49261,N_45416,N_47376);
nor U49262 (N_49262,N_45829,N_46328);
xor U49263 (N_49263,N_45484,N_46925);
nand U49264 (N_49264,N_46811,N_46243);
nand U49265 (N_49265,N_45203,N_46093);
nand U49266 (N_49266,N_45306,N_47188);
nand U49267 (N_49267,N_46778,N_47363);
xnor U49268 (N_49268,N_45545,N_47217);
nand U49269 (N_49269,N_47499,N_45325);
and U49270 (N_49270,N_47026,N_47109);
xor U49271 (N_49271,N_45855,N_46037);
xor U49272 (N_49272,N_47198,N_46907);
xnor U49273 (N_49273,N_46262,N_45717);
nor U49274 (N_49274,N_46538,N_45727);
xor U49275 (N_49275,N_47089,N_47498);
nand U49276 (N_49276,N_46053,N_47021);
or U49277 (N_49277,N_45350,N_46841);
nor U49278 (N_49278,N_45598,N_46732);
nor U49279 (N_49279,N_47080,N_46682);
nand U49280 (N_49280,N_45352,N_45519);
and U49281 (N_49281,N_45268,N_47221);
or U49282 (N_49282,N_46601,N_46833);
or U49283 (N_49283,N_45182,N_45437);
or U49284 (N_49284,N_47438,N_45880);
nor U49285 (N_49285,N_46444,N_45211);
or U49286 (N_49286,N_47080,N_47383);
and U49287 (N_49287,N_47087,N_45325);
and U49288 (N_49288,N_45422,N_47342);
nor U49289 (N_49289,N_45373,N_45638);
and U49290 (N_49290,N_45261,N_47032);
xnor U49291 (N_49291,N_47260,N_46789);
xnor U49292 (N_49292,N_47240,N_45338);
nor U49293 (N_49293,N_46960,N_45132);
or U49294 (N_49294,N_45766,N_45288);
nor U49295 (N_49295,N_45719,N_46130);
and U49296 (N_49296,N_46271,N_46167);
xnor U49297 (N_49297,N_46225,N_47389);
nand U49298 (N_49298,N_47259,N_46664);
nor U49299 (N_49299,N_46724,N_46278);
and U49300 (N_49300,N_45954,N_45650);
or U49301 (N_49301,N_46085,N_47212);
and U49302 (N_49302,N_45154,N_46807);
nor U49303 (N_49303,N_45889,N_45788);
or U49304 (N_49304,N_45631,N_46323);
nand U49305 (N_49305,N_45765,N_47054);
and U49306 (N_49306,N_45757,N_46786);
nand U49307 (N_49307,N_46141,N_45638);
or U49308 (N_49308,N_46906,N_45572);
nor U49309 (N_49309,N_46356,N_46863);
xnor U49310 (N_49310,N_46430,N_47221);
nand U49311 (N_49311,N_46382,N_45086);
and U49312 (N_49312,N_46046,N_46894);
or U49313 (N_49313,N_45767,N_45355);
and U49314 (N_49314,N_45728,N_45178);
and U49315 (N_49315,N_45199,N_45571);
nand U49316 (N_49316,N_47410,N_45268);
xor U49317 (N_49317,N_45050,N_47249);
nor U49318 (N_49318,N_46889,N_46048);
nor U49319 (N_49319,N_46004,N_45385);
nand U49320 (N_49320,N_47338,N_45926);
or U49321 (N_49321,N_45858,N_47327);
nor U49322 (N_49322,N_46055,N_46018);
or U49323 (N_49323,N_46132,N_46570);
nand U49324 (N_49324,N_46367,N_45131);
or U49325 (N_49325,N_47070,N_45729);
xor U49326 (N_49326,N_46079,N_46535);
nor U49327 (N_49327,N_47022,N_45483);
and U49328 (N_49328,N_46219,N_45911);
nand U49329 (N_49329,N_45681,N_46823);
and U49330 (N_49330,N_45728,N_45883);
xnor U49331 (N_49331,N_47126,N_45504);
nand U49332 (N_49332,N_47234,N_47063);
and U49333 (N_49333,N_46642,N_46285);
xnor U49334 (N_49334,N_45178,N_46916);
nor U49335 (N_49335,N_45810,N_45716);
nand U49336 (N_49336,N_45807,N_45510);
and U49337 (N_49337,N_45742,N_47414);
xor U49338 (N_49338,N_45091,N_45479);
nand U49339 (N_49339,N_47408,N_45479);
nor U49340 (N_49340,N_45252,N_46794);
and U49341 (N_49341,N_45002,N_45497);
and U49342 (N_49342,N_45533,N_46875);
xnor U49343 (N_49343,N_47112,N_46646);
xor U49344 (N_49344,N_45167,N_45454);
xor U49345 (N_49345,N_45943,N_45980);
and U49346 (N_49346,N_47088,N_47023);
nor U49347 (N_49347,N_46587,N_47429);
xnor U49348 (N_49348,N_45433,N_47297);
nor U49349 (N_49349,N_46862,N_46519);
nor U49350 (N_49350,N_47174,N_45074);
and U49351 (N_49351,N_47468,N_47282);
nor U49352 (N_49352,N_46466,N_46588);
nand U49353 (N_49353,N_46640,N_46417);
xnor U49354 (N_49354,N_47078,N_45631);
and U49355 (N_49355,N_45319,N_46821);
and U49356 (N_49356,N_47418,N_45185);
nand U49357 (N_49357,N_46857,N_47395);
nor U49358 (N_49358,N_47068,N_45701);
nand U49359 (N_49359,N_46175,N_45828);
nand U49360 (N_49360,N_46194,N_46061);
nand U49361 (N_49361,N_45125,N_45249);
nand U49362 (N_49362,N_45283,N_45589);
xnor U49363 (N_49363,N_46777,N_45960);
or U49364 (N_49364,N_46060,N_45420);
nand U49365 (N_49365,N_46802,N_45288);
nor U49366 (N_49366,N_45988,N_47456);
nand U49367 (N_49367,N_46739,N_45094);
xnor U49368 (N_49368,N_47482,N_46259);
nor U49369 (N_49369,N_46725,N_45663);
nor U49370 (N_49370,N_45227,N_47393);
and U49371 (N_49371,N_47461,N_45404);
nor U49372 (N_49372,N_46179,N_46210);
or U49373 (N_49373,N_46078,N_45542);
nand U49374 (N_49374,N_46703,N_46763);
nor U49375 (N_49375,N_45749,N_45436);
xnor U49376 (N_49376,N_45765,N_47150);
and U49377 (N_49377,N_45002,N_46655);
nor U49378 (N_49378,N_45187,N_46359);
nand U49379 (N_49379,N_47216,N_45351);
nand U49380 (N_49380,N_46077,N_45166);
or U49381 (N_49381,N_45246,N_47059);
and U49382 (N_49382,N_45890,N_47389);
xnor U49383 (N_49383,N_46143,N_46499);
nor U49384 (N_49384,N_46141,N_47353);
nor U49385 (N_49385,N_45988,N_47122);
and U49386 (N_49386,N_46104,N_46327);
xnor U49387 (N_49387,N_45852,N_45360);
nand U49388 (N_49388,N_46686,N_46493);
or U49389 (N_49389,N_45428,N_47186);
or U49390 (N_49390,N_47063,N_46844);
nand U49391 (N_49391,N_45021,N_45565);
nand U49392 (N_49392,N_46091,N_46198);
xor U49393 (N_49393,N_46773,N_45811);
nor U49394 (N_49394,N_46630,N_46500);
nor U49395 (N_49395,N_46056,N_46489);
nand U49396 (N_49396,N_45271,N_45244);
or U49397 (N_49397,N_46320,N_47292);
and U49398 (N_49398,N_45033,N_47096);
and U49399 (N_49399,N_46486,N_45171);
and U49400 (N_49400,N_46116,N_46490);
and U49401 (N_49401,N_46003,N_45327);
nor U49402 (N_49402,N_46323,N_46998);
xnor U49403 (N_49403,N_46996,N_46701);
nand U49404 (N_49404,N_47411,N_45820);
nand U49405 (N_49405,N_46031,N_46941);
or U49406 (N_49406,N_47360,N_46097);
nand U49407 (N_49407,N_46831,N_46455);
nand U49408 (N_49408,N_46070,N_45998);
nor U49409 (N_49409,N_46536,N_47187);
and U49410 (N_49410,N_45098,N_46586);
nand U49411 (N_49411,N_47110,N_45952);
nor U49412 (N_49412,N_46787,N_47323);
nand U49413 (N_49413,N_45436,N_46366);
nor U49414 (N_49414,N_46874,N_45792);
and U49415 (N_49415,N_47001,N_46746);
nand U49416 (N_49416,N_45762,N_46937);
nand U49417 (N_49417,N_45407,N_46725);
xnor U49418 (N_49418,N_47010,N_45599);
xor U49419 (N_49419,N_46075,N_47400);
nand U49420 (N_49420,N_45597,N_45463);
and U49421 (N_49421,N_46502,N_45300);
nand U49422 (N_49422,N_45676,N_47068);
xnor U49423 (N_49423,N_46900,N_46170);
nor U49424 (N_49424,N_45107,N_46426);
and U49425 (N_49425,N_47444,N_46445);
nand U49426 (N_49426,N_47395,N_47325);
nand U49427 (N_49427,N_45775,N_46886);
nand U49428 (N_49428,N_45149,N_46268);
or U49429 (N_49429,N_45068,N_45846);
nand U49430 (N_49430,N_46461,N_45705);
and U49431 (N_49431,N_46514,N_45065);
or U49432 (N_49432,N_45190,N_45096);
xor U49433 (N_49433,N_45747,N_45670);
nand U49434 (N_49434,N_45295,N_45567);
nor U49435 (N_49435,N_46530,N_45104);
nor U49436 (N_49436,N_45029,N_45538);
nor U49437 (N_49437,N_45875,N_45625);
nand U49438 (N_49438,N_45520,N_46572);
or U49439 (N_49439,N_46697,N_45010);
nand U49440 (N_49440,N_46599,N_45599);
xnor U49441 (N_49441,N_46792,N_46528);
or U49442 (N_49442,N_46783,N_46052);
xor U49443 (N_49443,N_45797,N_47057);
nor U49444 (N_49444,N_45092,N_46437);
nor U49445 (N_49445,N_45452,N_45231);
and U49446 (N_49446,N_45020,N_46298);
nand U49447 (N_49447,N_47134,N_45802);
xnor U49448 (N_49448,N_45722,N_46378);
or U49449 (N_49449,N_46720,N_46520);
xor U49450 (N_49450,N_46742,N_46053);
xor U49451 (N_49451,N_47216,N_47478);
xor U49452 (N_49452,N_46516,N_45121);
nor U49453 (N_49453,N_46917,N_45830);
nand U49454 (N_49454,N_46118,N_45389);
and U49455 (N_49455,N_45391,N_46083);
and U49456 (N_49456,N_46196,N_45869);
and U49457 (N_49457,N_45966,N_46817);
nand U49458 (N_49458,N_46028,N_46735);
nand U49459 (N_49459,N_45701,N_47019);
or U49460 (N_49460,N_46131,N_46463);
or U49461 (N_49461,N_47312,N_46023);
xor U49462 (N_49462,N_45685,N_46482);
or U49463 (N_49463,N_47179,N_46030);
nor U49464 (N_49464,N_45769,N_46333);
xnor U49465 (N_49465,N_45945,N_46997);
and U49466 (N_49466,N_45149,N_46826);
and U49467 (N_49467,N_45519,N_45730);
and U49468 (N_49468,N_46620,N_47404);
nand U49469 (N_49469,N_45091,N_47283);
xor U49470 (N_49470,N_45127,N_46035);
and U49471 (N_49471,N_45550,N_45812);
nor U49472 (N_49472,N_47367,N_45820);
or U49473 (N_49473,N_46628,N_45066);
nor U49474 (N_49474,N_45423,N_45795);
nand U49475 (N_49475,N_45808,N_45189);
and U49476 (N_49476,N_46247,N_46325);
xnor U49477 (N_49477,N_46943,N_45437);
xor U49478 (N_49478,N_46848,N_45065);
nand U49479 (N_49479,N_46129,N_46631);
and U49480 (N_49480,N_46537,N_45679);
xnor U49481 (N_49481,N_45128,N_46650);
xor U49482 (N_49482,N_45284,N_45497);
nand U49483 (N_49483,N_47303,N_47032);
and U49484 (N_49484,N_45920,N_45819);
nand U49485 (N_49485,N_46314,N_46131);
or U49486 (N_49486,N_47156,N_45683);
or U49487 (N_49487,N_45818,N_46683);
and U49488 (N_49488,N_45913,N_47266);
or U49489 (N_49489,N_45798,N_46929);
nor U49490 (N_49490,N_45198,N_46049);
nor U49491 (N_49491,N_47105,N_45218);
nor U49492 (N_49492,N_45040,N_45436);
nand U49493 (N_49493,N_45614,N_45172);
nor U49494 (N_49494,N_45195,N_45847);
or U49495 (N_49495,N_45021,N_46722);
xnor U49496 (N_49496,N_45094,N_45502);
nor U49497 (N_49497,N_45287,N_47278);
nand U49498 (N_49498,N_45498,N_46097);
xor U49499 (N_49499,N_46984,N_46451);
nand U49500 (N_49500,N_45419,N_45360);
and U49501 (N_49501,N_47054,N_47236);
and U49502 (N_49502,N_45410,N_45850);
or U49503 (N_49503,N_45562,N_46561);
nor U49504 (N_49504,N_46713,N_46821);
xnor U49505 (N_49505,N_47105,N_45828);
xor U49506 (N_49506,N_47256,N_46105);
or U49507 (N_49507,N_45456,N_45647);
xnor U49508 (N_49508,N_46751,N_46838);
xor U49509 (N_49509,N_46231,N_47122);
and U49510 (N_49510,N_46779,N_45443);
xnor U49511 (N_49511,N_46379,N_46108);
nand U49512 (N_49512,N_45713,N_45611);
xor U49513 (N_49513,N_45561,N_47235);
xnor U49514 (N_49514,N_46036,N_45214);
nand U49515 (N_49515,N_45414,N_46482);
nor U49516 (N_49516,N_45782,N_46525);
or U49517 (N_49517,N_47135,N_47342);
xor U49518 (N_49518,N_46432,N_46215);
and U49519 (N_49519,N_45694,N_45122);
nand U49520 (N_49520,N_45452,N_45751);
nor U49521 (N_49521,N_46214,N_45235);
and U49522 (N_49522,N_46518,N_47343);
or U49523 (N_49523,N_46689,N_46257);
nand U49524 (N_49524,N_45599,N_47175);
nor U49525 (N_49525,N_46737,N_46380);
and U49526 (N_49526,N_45972,N_45153);
or U49527 (N_49527,N_45625,N_46611);
xor U49528 (N_49528,N_47011,N_46998);
nand U49529 (N_49529,N_47402,N_45472);
and U49530 (N_49530,N_46718,N_46334);
xnor U49531 (N_49531,N_47249,N_46464);
nor U49532 (N_49532,N_45753,N_45052);
or U49533 (N_49533,N_47116,N_45280);
and U49534 (N_49534,N_46587,N_47289);
xnor U49535 (N_49535,N_46088,N_47391);
or U49536 (N_49536,N_45799,N_45759);
xnor U49537 (N_49537,N_45159,N_47190);
xor U49538 (N_49538,N_46527,N_45154);
or U49539 (N_49539,N_46480,N_46467);
nor U49540 (N_49540,N_45322,N_46069);
nor U49541 (N_49541,N_46471,N_45655);
or U49542 (N_49542,N_45491,N_45656);
nor U49543 (N_49543,N_46693,N_45274);
and U49544 (N_49544,N_46186,N_46424);
or U49545 (N_49545,N_45809,N_47148);
or U49546 (N_49546,N_46574,N_45003);
nor U49547 (N_49547,N_46440,N_45104);
nor U49548 (N_49548,N_46281,N_47147);
nand U49549 (N_49549,N_47185,N_46528);
nor U49550 (N_49550,N_45449,N_46982);
nand U49551 (N_49551,N_46052,N_46056);
xor U49552 (N_49552,N_46248,N_45204);
nor U49553 (N_49553,N_46669,N_45219);
nor U49554 (N_49554,N_45857,N_46856);
nor U49555 (N_49555,N_46380,N_46042);
nor U49556 (N_49556,N_45736,N_45315);
and U49557 (N_49557,N_46854,N_46587);
nand U49558 (N_49558,N_47207,N_47138);
or U49559 (N_49559,N_45574,N_45208);
xor U49560 (N_49560,N_46007,N_45875);
and U49561 (N_49561,N_45613,N_46008);
xnor U49562 (N_49562,N_46748,N_47132);
or U49563 (N_49563,N_46858,N_45780);
or U49564 (N_49564,N_46843,N_47052);
nand U49565 (N_49565,N_45213,N_45175);
or U49566 (N_49566,N_47176,N_45774);
xor U49567 (N_49567,N_45968,N_45622);
or U49568 (N_49568,N_47480,N_46426);
xor U49569 (N_49569,N_45764,N_45338);
nand U49570 (N_49570,N_46738,N_46963);
nand U49571 (N_49571,N_46748,N_47040);
xnor U49572 (N_49572,N_46898,N_47212);
nor U49573 (N_49573,N_45046,N_47002);
or U49574 (N_49574,N_46222,N_46754);
nand U49575 (N_49575,N_45718,N_47026);
and U49576 (N_49576,N_45069,N_45624);
nor U49577 (N_49577,N_47441,N_46445);
xnor U49578 (N_49578,N_46301,N_45717);
or U49579 (N_49579,N_45811,N_45079);
or U49580 (N_49580,N_45470,N_46117);
and U49581 (N_49581,N_46187,N_46314);
or U49582 (N_49582,N_46194,N_46940);
or U49583 (N_49583,N_47307,N_47460);
nand U49584 (N_49584,N_45239,N_45989);
or U49585 (N_49585,N_46022,N_47345);
and U49586 (N_49586,N_47332,N_47269);
nand U49587 (N_49587,N_46497,N_46909);
and U49588 (N_49588,N_47328,N_46275);
nand U49589 (N_49589,N_45227,N_45534);
and U49590 (N_49590,N_46128,N_46808);
or U49591 (N_49591,N_47485,N_46935);
nor U49592 (N_49592,N_46497,N_45021);
and U49593 (N_49593,N_46568,N_46001);
and U49594 (N_49594,N_46903,N_46670);
xnor U49595 (N_49595,N_47150,N_45001);
xor U49596 (N_49596,N_46240,N_45764);
or U49597 (N_49597,N_47266,N_46455);
or U49598 (N_49598,N_46205,N_45395);
or U49599 (N_49599,N_45883,N_45473);
xnor U49600 (N_49600,N_45356,N_47258);
xor U49601 (N_49601,N_45183,N_47327);
or U49602 (N_49602,N_47266,N_47306);
and U49603 (N_49603,N_46161,N_46989);
or U49604 (N_49604,N_46883,N_46016);
or U49605 (N_49605,N_45499,N_45015);
nand U49606 (N_49606,N_46785,N_46500);
xnor U49607 (N_49607,N_47253,N_45831);
nor U49608 (N_49608,N_46701,N_47316);
or U49609 (N_49609,N_45348,N_46625);
or U49610 (N_49610,N_46724,N_47029);
nor U49611 (N_49611,N_46603,N_45345);
and U49612 (N_49612,N_45035,N_45812);
nand U49613 (N_49613,N_46033,N_47301);
and U49614 (N_49614,N_47224,N_45477);
nand U49615 (N_49615,N_45952,N_45672);
nand U49616 (N_49616,N_47170,N_46171);
nor U49617 (N_49617,N_45469,N_46771);
xnor U49618 (N_49618,N_46378,N_47023);
nor U49619 (N_49619,N_45745,N_45487);
or U49620 (N_49620,N_47179,N_45144);
or U49621 (N_49621,N_47311,N_45723);
or U49622 (N_49622,N_47136,N_47108);
or U49623 (N_49623,N_45979,N_46127);
or U49624 (N_49624,N_45158,N_47204);
and U49625 (N_49625,N_46495,N_45594);
xnor U49626 (N_49626,N_46095,N_46233);
and U49627 (N_49627,N_47485,N_46819);
or U49628 (N_49628,N_46950,N_45501);
nand U49629 (N_49629,N_47326,N_46491);
nor U49630 (N_49630,N_46615,N_46705);
xnor U49631 (N_49631,N_45041,N_45746);
xor U49632 (N_49632,N_45515,N_45516);
and U49633 (N_49633,N_45969,N_46496);
and U49634 (N_49634,N_45222,N_47244);
or U49635 (N_49635,N_46709,N_45310);
xnor U49636 (N_49636,N_45867,N_45853);
nor U49637 (N_49637,N_45052,N_46124);
xnor U49638 (N_49638,N_46325,N_46101);
xnor U49639 (N_49639,N_45971,N_45238);
xnor U49640 (N_49640,N_45590,N_47458);
nand U49641 (N_49641,N_46671,N_47316);
or U49642 (N_49642,N_47142,N_45321);
xor U49643 (N_49643,N_47217,N_46589);
nand U49644 (N_49644,N_45629,N_45782);
nand U49645 (N_49645,N_46673,N_46954);
nor U49646 (N_49646,N_46673,N_45186);
and U49647 (N_49647,N_46296,N_46968);
nand U49648 (N_49648,N_47314,N_45730);
nand U49649 (N_49649,N_46623,N_46526);
nand U49650 (N_49650,N_47131,N_46690);
or U49651 (N_49651,N_46037,N_46164);
xor U49652 (N_49652,N_45623,N_46214);
nand U49653 (N_49653,N_45967,N_47187);
and U49654 (N_49654,N_47341,N_45006);
nor U49655 (N_49655,N_45400,N_45628);
and U49656 (N_49656,N_45774,N_46469);
nor U49657 (N_49657,N_47308,N_46312);
or U49658 (N_49658,N_45562,N_47398);
nor U49659 (N_49659,N_47178,N_45076);
nand U49660 (N_49660,N_45916,N_46447);
nand U49661 (N_49661,N_46472,N_47412);
and U49662 (N_49662,N_46377,N_45498);
xnor U49663 (N_49663,N_45399,N_47421);
or U49664 (N_49664,N_47488,N_45590);
or U49665 (N_49665,N_46817,N_45126);
or U49666 (N_49666,N_46314,N_46148);
nor U49667 (N_49667,N_47225,N_47157);
nand U49668 (N_49668,N_45673,N_46591);
nand U49669 (N_49669,N_45955,N_45746);
nand U49670 (N_49670,N_45925,N_47293);
or U49671 (N_49671,N_46148,N_47110);
nand U49672 (N_49672,N_45154,N_47192);
xor U49673 (N_49673,N_45468,N_46326);
nor U49674 (N_49674,N_45743,N_46683);
nor U49675 (N_49675,N_46698,N_45020);
or U49676 (N_49676,N_46312,N_46299);
and U49677 (N_49677,N_45975,N_45278);
nand U49678 (N_49678,N_46933,N_46042);
and U49679 (N_49679,N_45393,N_47053);
nor U49680 (N_49680,N_47479,N_45095);
or U49681 (N_49681,N_46761,N_45731);
xor U49682 (N_49682,N_45806,N_47268);
and U49683 (N_49683,N_45721,N_45058);
nand U49684 (N_49684,N_46418,N_46732);
nand U49685 (N_49685,N_45570,N_45613);
or U49686 (N_49686,N_45211,N_46327);
nand U49687 (N_49687,N_46802,N_45276);
or U49688 (N_49688,N_45463,N_45090);
or U49689 (N_49689,N_45812,N_45064);
nand U49690 (N_49690,N_46783,N_47306);
xnor U49691 (N_49691,N_47140,N_46901);
nand U49692 (N_49692,N_46992,N_47205);
or U49693 (N_49693,N_46315,N_47252);
nand U49694 (N_49694,N_45124,N_46242);
xor U49695 (N_49695,N_45117,N_46585);
nand U49696 (N_49696,N_45433,N_45108);
nor U49697 (N_49697,N_47058,N_45443);
nand U49698 (N_49698,N_45174,N_45870);
nand U49699 (N_49699,N_46680,N_46787);
xnor U49700 (N_49700,N_45439,N_45315);
or U49701 (N_49701,N_46924,N_46909);
and U49702 (N_49702,N_45108,N_47031);
xor U49703 (N_49703,N_45677,N_45216);
and U49704 (N_49704,N_45809,N_45525);
and U49705 (N_49705,N_46010,N_45725);
xnor U49706 (N_49706,N_46670,N_45832);
xor U49707 (N_49707,N_45987,N_46492);
or U49708 (N_49708,N_45723,N_45113);
xnor U49709 (N_49709,N_46010,N_47205);
xnor U49710 (N_49710,N_45141,N_45165);
and U49711 (N_49711,N_47229,N_45018);
xor U49712 (N_49712,N_45065,N_47472);
xnor U49713 (N_49713,N_47379,N_46377);
xnor U49714 (N_49714,N_47099,N_46871);
nand U49715 (N_49715,N_46467,N_45088);
and U49716 (N_49716,N_47402,N_45849);
nand U49717 (N_49717,N_47016,N_46771);
and U49718 (N_49718,N_45972,N_45956);
nor U49719 (N_49719,N_46453,N_46351);
nor U49720 (N_49720,N_45554,N_45479);
or U49721 (N_49721,N_46552,N_45460);
or U49722 (N_49722,N_45395,N_45293);
or U49723 (N_49723,N_46221,N_47071);
nand U49724 (N_49724,N_45356,N_45274);
and U49725 (N_49725,N_46743,N_45898);
or U49726 (N_49726,N_47072,N_47024);
nor U49727 (N_49727,N_47421,N_46753);
and U49728 (N_49728,N_46953,N_45475);
nand U49729 (N_49729,N_45044,N_46362);
and U49730 (N_49730,N_45073,N_45339);
and U49731 (N_49731,N_45590,N_46335);
and U49732 (N_49732,N_46387,N_46832);
nor U49733 (N_49733,N_46821,N_47350);
or U49734 (N_49734,N_46301,N_46267);
and U49735 (N_49735,N_46554,N_46601);
or U49736 (N_49736,N_46759,N_47004);
nor U49737 (N_49737,N_45675,N_46836);
and U49738 (N_49738,N_46996,N_46370);
nand U49739 (N_49739,N_47359,N_46985);
nand U49740 (N_49740,N_45037,N_46977);
and U49741 (N_49741,N_45346,N_46078);
xor U49742 (N_49742,N_46564,N_46617);
and U49743 (N_49743,N_45495,N_45339);
nand U49744 (N_49744,N_47115,N_45919);
xnor U49745 (N_49745,N_46473,N_45255);
and U49746 (N_49746,N_45755,N_45471);
xnor U49747 (N_49747,N_45458,N_45671);
xor U49748 (N_49748,N_45094,N_45655);
or U49749 (N_49749,N_45258,N_45483);
nand U49750 (N_49750,N_47307,N_46959);
or U49751 (N_49751,N_45554,N_45419);
xor U49752 (N_49752,N_45720,N_47406);
nand U49753 (N_49753,N_46137,N_46543);
nor U49754 (N_49754,N_47098,N_46489);
and U49755 (N_49755,N_47073,N_45531);
and U49756 (N_49756,N_45302,N_46126);
xor U49757 (N_49757,N_46015,N_46393);
nand U49758 (N_49758,N_46497,N_45705);
nor U49759 (N_49759,N_46654,N_45101);
nand U49760 (N_49760,N_45308,N_46829);
nand U49761 (N_49761,N_45320,N_46663);
or U49762 (N_49762,N_47476,N_45574);
nand U49763 (N_49763,N_45851,N_45807);
or U49764 (N_49764,N_46129,N_45384);
xor U49765 (N_49765,N_45869,N_46699);
and U49766 (N_49766,N_47336,N_46309);
and U49767 (N_49767,N_46951,N_45430);
and U49768 (N_49768,N_45418,N_45945);
or U49769 (N_49769,N_45785,N_45004);
xnor U49770 (N_49770,N_46461,N_46830);
and U49771 (N_49771,N_46037,N_45373);
nor U49772 (N_49772,N_46197,N_45124);
or U49773 (N_49773,N_45071,N_45085);
and U49774 (N_49774,N_45219,N_45141);
nand U49775 (N_49775,N_45281,N_47143);
nor U49776 (N_49776,N_47208,N_46444);
and U49777 (N_49777,N_47010,N_46777);
nand U49778 (N_49778,N_45108,N_45475);
nand U49779 (N_49779,N_45026,N_46596);
and U49780 (N_49780,N_46899,N_46892);
and U49781 (N_49781,N_47006,N_47069);
xor U49782 (N_49782,N_45172,N_47087);
nor U49783 (N_49783,N_45418,N_46159);
and U49784 (N_49784,N_47160,N_47228);
xor U49785 (N_49785,N_46328,N_45170);
nor U49786 (N_49786,N_45067,N_46295);
or U49787 (N_49787,N_46528,N_45566);
nor U49788 (N_49788,N_45971,N_46042);
and U49789 (N_49789,N_45727,N_47351);
or U49790 (N_49790,N_46781,N_45046);
nor U49791 (N_49791,N_45830,N_45006);
or U49792 (N_49792,N_46163,N_46949);
nand U49793 (N_49793,N_46915,N_46472);
or U49794 (N_49794,N_46907,N_47433);
nor U49795 (N_49795,N_47193,N_46919);
and U49796 (N_49796,N_46630,N_45180);
or U49797 (N_49797,N_46517,N_46046);
or U49798 (N_49798,N_45256,N_46161);
and U49799 (N_49799,N_45453,N_46866);
xnor U49800 (N_49800,N_45250,N_46578);
and U49801 (N_49801,N_46358,N_46418);
nand U49802 (N_49802,N_45530,N_45193);
xor U49803 (N_49803,N_46261,N_45187);
nand U49804 (N_49804,N_47189,N_45366);
and U49805 (N_49805,N_46015,N_46276);
nand U49806 (N_49806,N_46023,N_45140);
or U49807 (N_49807,N_45896,N_47086);
nor U49808 (N_49808,N_46802,N_47330);
nand U49809 (N_49809,N_45375,N_45946);
nand U49810 (N_49810,N_46789,N_46319);
xnor U49811 (N_49811,N_47429,N_46816);
and U49812 (N_49812,N_46981,N_45005);
nand U49813 (N_49813,N_46385,N_47177);
and U49814 (N_49814,N_45367,N_45010);
and U49815 (N_49815,N_45952,N_46063);
nor U49816 (N_49816,N_47459,N_45198);
and U49817 (N_49817,N_46638,N_46358);
and U49818 (N_49818,N_45840,N_45355);
nand U49819 (N_49819,N_45300,N_46313);
and U49820 (N_49820,N_46067,N_47406);
and U49821 (N_49821,N_45355,N_46247);
and U49822 (N_49822,N_47007,N_45046);
nor U49823 (N_49823,N_46417,N_47088);
nor U49824 (N_49824,N_45717,N_46151);
or U49825 (N_49825,N_45977,N_46649);
nor U49826 (N_49826,N_45529,N_46094);
and U49827 (N_49827,N_45758,N_47374);
xor U49828 (N_49828,N_45154,N_46384);
nand U49829 (N_49829,N_46042,N_47063);
xor U49830 (N_49830,N_47276,N_45215);
and U49831 (N_49831,N_45551,N_45422);
and U49832 (N_49832,N_45885,N_45356);
xor U49833 (N_49833,N_45445,N_45446);
and U49834 (N_49834,N_46636,N_46484);
or U49835 (N_49835,N_46998,N_47457);
or U49836 (N_49836,N_46671,N_45436);
and U49837 (N_49837,N_46262,N_46973);
and U49838 (N_49838,N_47416,N_46846);
and U49839 (N_49839,N_46769,N_45808);
xnor U49840 (N_49840,N_47167,N_46202);
or U49841 (N_49841,N_45901,N_47499);
nand U49842 (N_49842,N_46716,N_46114);
or U49843 (N_49843,N_46193,N_45989);
nand U49844 (N_49844,N_46987,N_46268);
and U49845 (N_49845,N_45508,N_45230);
nor U49846 (N_49846,N_46014,N_47167);
and U49847 (N_49847,N_45164,N_45001);
and U49848 (N_49848,N_47390,N_45195);
or U49849 (N_49849,N_46620,N_46924);
nor U49850 (N_49850,N_45349,N_46239);
xnor U49851 (N_49851,N_46844,N_46881);
and U49852 (N_49852,N_46659,N_47062);
nand U49853 (N_49853,N_45598,N_46367);
xnor U49854 (N_49854,N_45284,N_45701);
nor U49855 (N_49855,N_46975,N_46583);
xor U49856 (N_49856,N_45534,N_45345);
or U49857 (N_49857,N_46748,N_45700);
xnor U49858 (N_49858,N_45286,N_46795);
xor U49859 (N_49859,N_46189,N_45084);
and U49860 (N_49860,N_45066,N_45678);
or U49861 (N_49861,N_45241,N_46901);
and U49862 (N_49862,N_45250,N_45636);
nand U49863 (N_49863,N_46190,N_46168);
and U49864 (N_49864,N_46995,N_45566);
and U49865 (N_49865,N_46869,N_45994);
xor U49866 (N_49866,N_45353,N_45340);
and U49867 (N_49867,N_45623,N_46388);
nand U49868 (N_49868,N_46746,N_46732);
xnor U49869 (N_49869,N_45809,N_45674);
or U49870 (N_49870,N_45637,N_46148);
or U49871 (N_49871,N_45573,N_46263);
or U49872 (N_49872,N_45815,N_47170);
nand U49873 (N_49873,N_45748,N_45716);
or U49874 (N_49874,N_45525,N_47004);
or U49875 (N_49875,N_45613,N_45567);
and U49876 (N_49876,N_46772,N_47164);
nor U49877 (N_49877,N_47114,N_46134);
or U49878 (N_49878,N_47496,N_47209);
xnor U49879 (N_49879,N_47349,N_46292);
nand U49880 (N_49880,N_46089,N_46263);
nand U49881 (N_49881,N_46835,N_46571);
nor U49882 (N_49882,N_47478,N_45520);
or U49883 (N_49883,N_45908,N_45222);
xor U49884 (N_49884,N_47302,N_45711);
or U49885 (N_49885,N_46213,N_46401);
or U49886 (N_49886,N_46614,N_45043);
and U49887 (N_49887,N_47199,N_45205);
nand U49888 (N_49888,N_45055,N_45933);
and U49889 (N_49889,N_46169,N_46215);
nor U49890 (N_49890,N_46500,N_45828);
or U49891 (N_49891,N_45775,N_46813);
nor U49892 (N_49892,N_45700,N_46249);
and U49893 (N_49893,N_45779,N_46314);
nand U49894 (N_49894,N_46397,N_45252);
nand U49895 (N_49895,N_47322,N_47345);
nand U49896 (N_49896,N_46185,N_46747);
or U49897 (N_49897,N_47219,N_46984);
and U49898 (N_49898,N_47125,N_46546);
nand U49899 (N_49899,N_47372,N_47177);
or U49900 (N_49900,N_45260,N_45995);
nand U49901 (N_49901,N_45813,N_46412);
and U49902 (N_49902,N_47402,N_45742);
nand U49903 (N_49903,N_46217,N_45665);
xor U49904 (N_49904,N_46144,N_46998);
xnor U49905 (N_49905,N_45895,N_46118);
nand U49906 (N_49906,N_46867,N_45616);
and U49907 (N_49907,N_45306,N_46115);
and U49908 (N_49908,N_45592,N_45867);
nor U49909 (N_49909,N_46010,N_45484);
or U49910 (N_49910,N_45107,N_45117);
nand U49911 (N_49911,N_47377,N_47485);
nor U49912 (N_49912,N_46784,N_47460);
or U49913 (N_49913,N_47430,N_47472);
and U49914 (N_49914,N_47419,N_45560);
nand U49915 (N_49915,N_47006,N_47132);
and U49916 (N_49916,N_47488,N_47374);
nand U49917 (N_49917,N_46619,N_45457);
or U49918 (N_49918,N_46288,N_45150);
nor U49919 (N_49919,N_47464,N_46427);
nand U49920 (N_49920,N_46197,N_46443);
nand U49921 (N_49921,N_46431,N_45630);
or U49922 (N_49922,N_46121,N_47020);
nor U49923 (N_49923,N_45818,N_46459);
nand U49924 (N_49924,N_45741,N_46836);
nand U49925 (N_49925,N_46023,N_45951);
nand U49926 (N_49926,N_47018,N_46741);
nand U49927 (N_49927,N_45756,N_45029);
or U49928 (N_49928,N_45403,N_47076);
xor U49929 (N_49929,N_46714,N_47479);
and U49930 (N_49930,N_46423,N_45606);
nor U49931 (N_49931,N_45433,N_45060);
nor U49932 (N_49932,N_46093,N_47266);
or U49933 (N_49933,N_46304,N_46160);
or U49934 (N_49934,N_46850,N_46165);
nand U49935 (N_49935,N_46698,N_46293);
nor U49936 (N_49936,N_46490,N_46667);
nor U49937 (N_49937,N_46807,N_46064);
and U49938 (N_49938,N_46767,N_46102);
xor U49939 (N_49939,N_46764,N_47396);
and U49940 (N_49940,N_47210,N_45937);
nand U49941 (N_49941,N_45772,N_46257);
xnor U49942 (N_49942,N_46579,N_46474);
nand U49943 (N_49943,N_47046,N_46104);
or U49944 (N_49944,N_46756,N_46075);
or U49945 (N_49945,N_46530,N_45148);
nor U49946 (N_49946,N_46186,N_47216);
nand U49947 (N_49947,N_47488,N_46021);
nand U49948 (N_49948,N_46731,N_47426);
nand U49949 (N_49949,N_46652,N_46803);
nor U49950 (N_49950,N_46403,N_46508);
and U49951 (N_49951,N_47336,N_47024);
nor U49952 (N_49952,N_45834,N_47138);
nand U49953 (N_49953,N_47243,N_46975);
or U49954 (N_49954,N_46366,N_47372);
and U49955 (N_49955,N_45697,N_46497);
and U49956 (N_49956,N_46751,N_45605);
or U49957 (N_49957,N_45197,N_45807);
and U49958 (N_49958,N_45935,N_46220);
and U49959 (N_49959,N_46128,N_46343);
and U49960 (N_49960,N_47075,N_46066);
nand U49961 (N_49961,N_45654,N_46578);
nand U49962 (N_49962,N_47081,N_45199);
nor U49963 (N_49963,N_45073,N_47136);
and U49964 (N_49964,N_46203,N_45065);
and U49965 (N_49965,N_46321,N_46972);
and U49966 (N_49966,N_45651,N_47273);
nand U49967 (N_49967,N_47214,N_45745);
nor U49968 (N_49968,N_46415,N_45901);
nand U49969 (N_49969,N_45613,N_47144);
and U49970 (N_49970,N_45935,N_46270);
nand U49971 (N_49971,N_46696,N_45876);
nand U49972 (N_49972,N_46682,N_45583);
xor U49973 (N_49973,N_46360,N_47071);
xnor U49974 (N_49974,N_46389,N_45493);
and U49975 (N_49975,N_47446,N_45807);
nand U49976 (N_49976,N_45221,N_46085);
xor U49977 (N_49977,N_45995,N_47284);
xnor U49978 (N_49978,N_45580,N_46844);
or U49979 (N_49979,N_47271,N_46532);
and U49980 (N_49980,N_45535,N_46053);
or U49981 (N_49981,N_46781,N_45614);
or U49982 (N_49982,N_46463,N_47414);
and U49983 (N_49983,N_45129,N_46960);
xor U49984 (N_49984,N_47326,N_45208);
or U49985 (N_49985,N_47140,N_45966);
xor U49986 (N_49986,N_47125,N_46574);
xnor U49987 (N_49987,N_46413,N_45331);
and U49988 (N_49988,N_45631,N_47352);
nor U49989 (N_49989,N_45387,N_46149);
xnor U49990 (N_49990,N_46656,N_46182);
and U49991 (N_49991,N_45076,N_46362);
or U49992 (N_49992,N_45561,N_46818);
and U49993 (N_49993,N_45877,N_46968);
nand U49994 (N_49994,N_47498,N_46195);
xnor U49995 (N_49995,N_46364,N_47049);
or U49996 (N_49996,N_47209,N_47044);
or U49997 (N_49997,N_46320,N_46121);
and U49998 (N_49998,N_46793,N_46361);
or U49999 (N_49999,N_47395,N_45577);
or UO_0 (O_0,N_48172,N_49415);
or UO_1 (O_1,N_49808,N_49610);
xor UO_2 (O_2,N_48189,N_49779);
xnor UO_3 (O_3,N_47734,N_49380);
nand UO_4 (O_4,N_49177,N_48432);
and UO_5 (O_5,N_49298,N_48804);
and UO_6 (O_6,N_47821,N_49401);
xnor UO_7 (O_7,N_49885,N_48501);
xor UO_8 (O_8,N_48291,N_49927);
xnor UO_9 (O_9,N_48798,N_47731);
nand UO_10 (O_10,N_49082,N_48465);
nand UO_11 (O_11,N_47977,N_47833);
nor UO_12 (O_12,N_49299,N_49780);
nor UO_13 (O_13,N_48483,N_49828);
xor UO_14 (O_14,N_49463,N_48310);
nor UO_15 (O_15,N_48005,N_49941);
and UO_16 (O_16,N_49497,N_48645);
and UO_17 (O_17,N_49252,N_49963);
and UO_18 (O_18,N_49353,N_47640);
nor UO_19 (O_19,N_48195,N_48082);
or UO_20 (O_20,N_49293,N_49996);
and UO_21 (O_21,N_49702,N_48306);
xor UO_22 (O_22,N_47824,N_48075);
nor UO_23 (O_23,N_49510,N_47781);
and UO_24 (O_24,N_49768,N_49373);
or UO_25 (O_25,N_48974,N_47930);
and UO_26 (O_26,N_48167,N_48695);
nand UO_27 (O_27,N_48790,N_49660);
nor UO_28 (O_28,N_48757,N_49578);
nand UO_29 (O_29,N_48472,N_49931);
nand UO_30 (O_30,N_49844,N_48540);
xor UO_31 (O_31,N_49449,N_48103);
nand UO_32 (O_32,N_47865,N_49980);
xor UO_33 (O_33,N_48754,N_48872);
xor UO_34 (O_34,N_49753,N_48234);
or UO_35 (O_35,N_47732,N_49146);
and UO_36 (O_36,N_49048,N_49511);
nand UO_37 (O_37,N_47700,N_48666);
xor UO_38 (O_38,N_47686,N_49688);
nand UO_39 (O_39,N_49607,N_49478);
xor UO_40 (O_40,N_47931,N_48841);
nor UO_41 (O_41,N_47815,N_49906);
nor UO_42 (O_42,N_47762,N_49235);
nand UO_43 (O_43,N_49932,N_49358);
nand UO_44 (O_44,N_49872,N_49646);
or UO_45 (O_45,N_49149,N_48358);
or UO_46 (O_46,N_48218,N_49655);
nand UO_47 (O_47,N_47757,N_48409);
xor UO_48 (O_48,N_47982,N_48773);
or UO_49 (O_49,N_47979,N_48111);
xnor UO_50 (O_50,N_48400,N_49131);
xor UO_51 (O_51,N_47631,N_49769);
nor UO_52 (O_52,N_49862,N_49217);
and UO_53 (O_53,N_49133,N_49671);
or UO_54 (O_54,N_48426,N_49331);
and UO_55 (O_55,N_47605,N_49632);
or UO_56 (O_56,N_49124,N_48289);
or UO_57 (O_57,N_49583,N_49046);
and UO_58 (O_58,N_48343,N_47510);
nor UO_59 (O_59,N_47905,N_49122);
and UO_60 (O_60,N_49759,N_47825);
and UO_61 (O_61,N_48392,N_49413);
nand UO_62 (O_62,N_48613,N_47683);
xnor UO_63 (O_63,N_49002,N_48003);
xor UO_64 (O_64,N_48920,N_48131);
or UO_65 (O_65,N_49717,N_48647);
or UO_66 (O_66,N_48593,N_49487);
nand UO_67 (O_67,N_48599,N_49575);
and UO_68 (O_68,N_49917,N_47654);
or UO_69 (O_69,N_48661,N_49153);
xnor UO_70 (O_70,N_47594,N_48406);
and UO_71 (O_71,N_47780,N_49335);
nor UO_72 (O_72,N_48524,N_48255);
nor UO_73 (O_73,N_48242,N_49110);
and UO_74 (O_74,N_47790,N_49870);
nand UO_75 (O_75,N_49563,N_48579);
or UO_76 (O_76,N_48534,N_48575);
and UO_77 (O_77,N_49956,N_49363);
and UO_78 (O_78,N_49374,N_47990);
and UO_79 (O_79,N_49159,N_49633);
nand UO_80 (O_80,N_48717,N_48527);
nand UO_81 (O_81,N_49275,N_49945);
and UO_82 (O_82,N_49831,N_49129);
nand UO_83 (O_83,N_49522,N_48238);
or UO_84 (O_84,N_48839,N_49326);
xnor UO_85 (O_85,N_48097,N_47832);
nor UO_86 (O_86,N_47848,N_48084);
and UO_87 (O_87,N_49384,N_49710);
xor UO_88 (O_88,N_49545,N_48022);
or UO_89 (O_89,N_48759,N_48700);
and UO_90 (O_90,N_49071,N_48794);
nor UO_91 (O_91,N_47627,N_48685);
nand UO_92 (O_92,N_49183,N_49553);
nor UO_93 (O_93,N_48824,N_48982);
or UO_94 (O_94,N_48994,N_48591);
nand UO_95 (O_95,N_49623,N_48679);
nand UO_96 (O_96,N_49645,N_47554);
nand UO_97 (O_97,N_48269,N_47634);
or UO_98 (O_98,N_48987,N_47808);
and UO_99 (O_99,N_48514,N_48037);
nand UO_100 (O_100,N_49277,N_49695);
nand UO_101 (O_101,N_49791,N_49954);
nand UO_102 (O_102,N_48014,N_47957);
or UO_103 (O_103,N_49976,N_48651);
xnor UO_104 (O_104,N_49044,N_47692);
nor UO_105 (O_105,N_48251,N_49852);
nor UO_106 (O_106,N_48240,N_49083);
nor UO_107 (O_107,N_47942,N_49765);
nand UO_108 (O_108,N_49892,N_48417);
xor UO_109 (O_109,N_47657,N_49547);
nand UO_110 (O_110,N_48021,N_48129);
or UO_111 (O_111,N_48668,N_49115);
or UO_112 (O_112,N_49014,N_49795);
or UO_113 (O_113,N_49261,N_48249);
nand UO_114 (O_114,N_47818,N_47630);
nor UO_115 (O_115,N_49050,N_48962);
or UO_116 (O_116,N_48142,N_47948);
nand UO_117 (O_117,N_49657,N_49724);
nand UO_118 (O_118,N_48891,N_49809);
nand UO_119 (O_119,N_48074,N_49108);
nor UO_120 (O_120,N_48963,N_48487);
or UO_121 (O_121,N_48282,N_49191);
and UO_122 (O_122,N_49447,N_49772);
nor UO_123 (O_123,N_48944,N_47590);
and UO_124 (O_124,N_49425,N_49987);
xnor UO_125 (O_125,N_48710,N_47584);
and UO_126 (O_126,N_49738,N_49306);
xor UO_127 (O_127,N_49601,N_49006);
nor UO_128 (O_128,N_49243,N_48319);
and UO_129 (O_129,N_47792,N_48040);
nor UO_130 (O_130,N_49784,N_47917);
and UO_131 (O_131,N_47847,N_47677);
xor UO_132 (O_132,N_48612,N_47711);
nand UO_133 (O_133,N_48544,N_48394);
and UO_134 (O_134,N_49584,N_48217);
and UO_135 (O_135,N_48069,N_48945);
nor UO_136 (O_136,N_48276,N_48985);
xnor UO_137 (O_137,N_48758,N_48870);
and UO_138 (O_138,N_47876,N_48976);
and UO_139 (O_139,N_48862,N_49145);
nor UO_140 (O_140,N_49340,N_47927);
nor UO_141 (O_141,N_48092,N_48328);
or UO_142 (O_142,N_48363,N_49405);
nor UO_143 (O_143,N_49749,N_48865);
or UO_144 (O_144,N_48342,N_49682);
and UO_145 (O_145,N_49643,N_48315);
nand UO_146 (O_146,N_49169,N_47563);
nor UO_147 (O_147,N_47937,N_49546);
xor UO_148 (O_148,N_48653,N_48546);
or UO_149 (O_149,N_47884,N_48590);
xnor UO_150 (O_150,N_48485,N_48478);
nand UO_151 (O_151,N_47761,N_49496);
or UO_152 (O_152,N_48634,N_49286);
xor UO_153 (O_153,N_48529,N_49250);
xor UO_154 (O_154,N_48890,N_49075);
xnor UO_155 (O_155,N_49818,N_48012);
xor UO_156 (O_156,N_49838,N_49567);
nand UO_157 (O_157,N_49391,N_48229);
or UO_158 (O_158,N_49198,N_48340);
xor UO_159 (O_159,N_47669,N_49403);
xor UO_160 (O_160,N_49411,N_49562);
nor UO_161 (O_161,N_49782,N_49664);
nand UO_162 (O_162,N_48563,N_48620);
or UO_163 (O_163,N_49744,N_48638);
or UO_164 (O_164,N_49857,N_48606);
or UO_165 (O_165,N_47813,N_49961);
nor UO_166 (O_166,N_48702,N_48813);
or UO_167 (O_167,N_49850,N_49897);
and UO_168 (O_168,N_49246,N_47585);
or UO_169 (O_169,N_49788,N_48497);
xnor UO_170 (O_170,N_48712,N_47858);
xnor UO_171 (O_171,N_49477,N_48854);
or UO_172 (O_172,N_48280,N_49541);
and UO_173 (O_173,N_47527,N_49459);
and UO_174 (O_174,N_47795,N_49792);
nor UO_175 (O_175,N_49034,N_48852);
and UO_176 (O_176,N_47500,N_48762);
nor UO_177 (O_177,N_48678,N_48808);
nand UO_178 (O_178,N_47663,N_47685);
xnor UO_179 (O_179,N_49849,N_48148);
or UO_180 (O_180,N_47863,N_49057);
nor UO_181 (O_181,N_48267,N_48745);
and UO_182 (O_182,N_48635,N_49348);
nand UO_183 (O_183,N_47609,N_49011);
nand UO_184 (O_184,N_48382,N_49408);
xor UO_185 (O_185,N_49543,N_49232);
nor UO_186 (O_186,N_49733,N_47501);
or UO_187 (O_187,N_49821,N_48515);
nor UO_188 (O_188,N_48309,N_47633);
xnor UO_189 (O_189,N_49616,N_47870);
nor UO_190 (O_190,N_47737,N_47976);
nor UO_191 (O_191,N_48895,N_49407);
and UO_192 (O_192,N_48397,N_49983);
and UO_193 (O_193,N_49495,N_48761);
or UO_194 (O_194,N_49958,N_47598);
nand UO_195 (O_195,N_49182,N_48299);
nand UO_196 (O_196,N_47643,N_48652);
xor UO_197 (O_197,N_48107,N_48477);
nand UO_198 (O_198,N_47577,N_49879);
or UO_199 (O_199,N_47610,N_49851);
or UO_200 (O_200,N_47749,N_48995);
or UO_201 (O_201,N_47955,N_47529);
nor UO_202 (O_202,N_49735,N_49536);
or UO_203 (O_203,N_48733,N_47759);
nand UO_204 (O_204,N_49533,N_48272);
and UO_205 (O_205,N_49585,N_49923);
nand UO_206 (O_206,N_47509,N_48126);
nand UO_207 (O_207,N_49040,N_47655);
nand UO_208 (O_208,N_48191,N_48959);
and UO_209 (O_209,N_47600,N_48327);
nand UO_210 (O_210,N_47629,N_49196);
nor UO_211 (O_211,N_49539,N_48338);
or UO_212 (O_212,N_48860,N_47772);
xnor UO_213 (O_213,N_49066,N_47557);
or UO_214 (O_214,N_47933,N_49924);
nand UO_215 (O_215,N_48031,N_49648);
xnor UO_216 (O_216,N_48175,N_49909);
nor UO_217 (O_217,N_48499,N_47862);
and UO_218 (O_218,N_49666,N_47713);
xnor UO_219 (O_219,N_47922,N_49992);
or UO_220 (O_220,N_49550,N_47779);
xor UO_221 (O_221,N_47932,N_47622);
and UO_222 (O_222,N_49801,N_49910);
and UO_223 (O_223,N_49908,N_48732);
and UO_224 (O_224,N_48709,N_49900);
or UO_225 (O_225,N_48973,N_48505);
nor UO_226 (O_226,N_48654,N_48004);
and UO_227 (O_227,N_47969,N_48064);
nor UO_228 (O_228,N_47688,N_49171);
and UO_229 (O_229,N_48099,N_49935);
xor UO_230 (O_230,N_48821,N_48248);
xor UO_231 (O_231,N_49835,N_48346);
or UO_232 (O_232,N_47588,N_49450);
or UO_233 (O_233,N_49309,N_48876);
nand UO_234 (O_234,N_47910,N_48106);
and UO_235 (O_235,N_49895,N_48859);
or UO_236 (O_236,N_48051,N_49292);
nand UO_237 (O_237,N_48531,N_49319);
xnor UO_238 (O_238,N_47934,N_47507);
nor UO_239 (O_239,N_48155,N_47964);
xnor UO_240 (O_240,N_49609,N_49767);
or UO_241 (O_241,N_48689,N_48368);
nand UO_242 (O_242,N_49558,N_49242);
and UO_243 (O_243,N_49134,N_48179);
or UO_244 (O_244,N_49042,N_48512);
and UO_245 (O_245,N_48916,N_48707);
nor UO_246 (O_246,N_48204,N_48245);
nor UO_247 (O_247,N_48354,N_49989);
nor UO_248 (O_248,N_48781,N_47562);
nor UO_249 (O_249,N_49868,N_47788);
or UO_250 (O_250,N_48969,N_47599);
xnor UO_251 (O_251,N_49869,N_47637);
and UO_252 (O_252,N_48079,N_47907);
or UO_253 (O_253,N_48027,N_47973);
nand UO_254 (O_254,N_48940,N_48493);
nor UO_255 (O_255,N_47889,N_49969);
and UO_256 (O_256,N_48318,N_49675);
nand UO_257 (O_257,N_49622,N_49499);
nand UO_258 (O_258,N_49836,N_48894);
and UO_259 (O_259,N_49775,N_48096);
nor UO_260 (O_260,N_48128,N_49344);
or UO_261 (O_261,N_48536,N_49460);
or UO_262 (O_262,N_48313,N_48185);
xnor UO_263 (O_263,N_49858,N_48122);
xor UO_264 (O_264,N_48461,N_49760);
nand UO_265 (O_265,N_49197,N_48362);
nand UO_266 (O_266,N_49757,N_49955);
or UO_267 (O_267,N_49631,N_49611);
and UO_268 (O_268,N_49883,N_47668);
nand UO_269 (O_269,N_48482,N_47911);
and UO_270 (O_270,N_49126,N_49053);
nor UO_271 (O_271,N_47791,N_48058);
or UO_272 (O_272,N_48323,N_48113);
or UO_273 (O_273,N_49940,N_48674);
nor UO_274 (O_274,N_47589,N_48750);
xor UO_275 (O_275,N_49445,N_49804);
nand UO_276 (O_276,N_49451,N_49297);
nor UO_277 (O_277,N_47893,N_48441);
or UO_278 (O_278,N_48152,N_48981);
nor UO_279 (O_279,N_49922,N_47623);
nor UO_280 (O_280,N_47604,N_47597);
and UO_281 (O_281,N_48246,N_48035);
nand UO_282 (O_282,N_49178,N_49117);
nand UO_283 (O_283,N_48223,N_49711);
or UO_284 (O_284,N_48873,N_47929);
xnor UO_285 (O_285,N_48206,N_48412);
or UO_286 (O_286,N_49412,N_48202);
or UO_287 (O_287,N_49934,N_49342);
nand UO_288 (O_288,N_49555,N_48151);
nand UO_289 (O_289,N_49520,N_49679);
xor UO_290 (O_290,N_48548,N_48506);
nand UO_291 (O_291,N_47582,N_47816);
nor UO_292 (O_292,N_47850,N_48334);
and UO_293 (O_293,N_48519,N_49314);
nand UO_294 (O_294,N_47648,N_48853);
or UO_295 (O_295,N_47671,N_49708);
nand UO_296 (O_296,N_48110,N_48468);
nand UO_297 (O_297,N_49901,N_48384);
xor UO_298 (O_298,N_49826,N_48370);
xor UO_299 (O_299,N_48573,N_48576);
nor UO_300 (O_300,N_49300,N_48207);
xor UO_301 (O_301,N_48596,N_48583);
nand UO_302 (O_302,N_49696,N_49698);
and UO_303 (O_303,N_49725,N_48210);
nand UO_304 (O_304,N_49840,N_47658);
nor UO_305 (O_305,N_49074,N_47550);
or UO_306 (O_306,N_48680,N_48927);
nand UO_307 (O_307,N_48383,N_48366);
nand UO_308 (O_308,N_48756,N_48632);
and UO_309 (O_309,N_49005,N_49957);
or UO_310 (O_310,N_48802,N_48067);
xor UO_311 (O_311,N_48855,N_48211);
and UO_312 (O_312,N_49164,N_49274);
nor UO_313 (O_313,N_49077,N_49301);
xor UO_314 (O_314,N_49204,N_48164);
and UO_315 (O_315,N_47768,N_48112);
nor UO_316 (O_316,N_49998,N_48949);
nor UO_317 (O_317,N_48329,N_48522);
nand UO_318 (O_318,N_48715,N_49316);
and UO_319 (O_319,N_49263,N_49336);
nor UO_320 (O_320,N_48119,N_48900);
xor UO_321 (O_321,N_47817,N_47804);
and UO_322 (O_322,N_49526,N_49685);
or UO_323 (O_323,N_47705,N_48013);
or UO_324 (O_324,N_47941,N_49026);
xnor UO_325 (O_325,N_49069,N_49328);
nor UO_326 (O_326,N_49490,N_49853);
xor UO_327 (O_327,N_49534,N_49111);
or UO_328 (O_328,N_49990,N_49639);
nand UO_329 (O_329,N_49233,N_48157);
xor UO_330 (O_330,N_48922,N_48102);
or UO_331 (O_331,N_48261,N_48029);
xor UO_332 (O_332,N_48034,N_48297);
nand UO_333 (O_333,N_49021,N_49942);
nor UO_334 (O_334,N_49078,N_47803);
or UO_335 (O_335,N_49742,N_47851);
and UO_336 (O_336,N_47972,N_49439);
and UO_337 (O_337,N_48684,N_49670);
nand UO_338 (O_338,N_48930,N_48800);
xor UO_339 (O_339,N_48589,N_49093);
nor UO_340 (O_340,N_49973,N_49148);
xor UO_341 (O_341,N_48834,N_49579);
or UO_342 (O_342,N_49588,N_48597);
nand UO_343 (O_343,N_49701,N_49023);
nor UO_344 (O_344,N_48349,N_49874);
nor UO_345 (O_345,N_47620,N_48050);
or UO_346 (O_346,N_49891,N_49059);
nand UO_347 (O_347,N_48615,N_47837);
nand UO_348 (O_348,N_49338,N_48311);
nand UO_349 (O_349,N_49523,N_49694);
and UO_350 (O_350,N_48026,N_48015);
nor UO_351 (O_351,N_48275,N_47614);
nand UO_352 (O_352,N_49448,N_49677);
nand UO_353 (O_353,N_49513,N_49476);
and UO_354 (O_354,N_48782,N_48221);
nor UO_355 (O_355,N_48988,N_49947);
and UO_356 (O_356,N_48060,N_49429);
xnor UO_357 (O_357,N_49847,N_48376);
nor UO_358 (O_358,N_48183,N_47756);
nor UO_359 (O_359,N_47727,N_49521);
xor UO_360 (O_360,N_48190,N_48550);
nor UO_361 (O_361,N_49970,N_48033);
and UO_362 (O_362,N_49193,N_48233);
xor UO_363 (O_363,N_48322,N_47784);
nand UO_364 (O_364,N_48510,N_48729);
xor UO_365 (O_365,N_48716,N_49746);
nand UO_366 (O_366,N_48828,N_47836);
or UO_367 (O_367,N_49615,N_49247);
xnor UO_368 (O_368,N_47699,N_49919);
nand UO_369 (O_369,N_49602,N_49525);
or UO_370 (O_370,N_49498,N_48101);
nor UO_371 (O_371,N_48120,N_49152);
nor UO_372 (O_372,N_48650,N_49729);
nand UO_373 (O_373,N_47698,N_48134);
nor UO_374 (O_374,N_49488,N_47827);
and UO_375 (O_375,N_48455,N_49995);
nor UO_376 (O_376,N_48147,N_49916);
and UO_377 (O_377,N_48078,N_49007);
and UO_378 (O_378,N_48177,N_48213);
xor UO_379 (O_379,N_48814,N_49067);
nor UO_380 (O_380,N_47971,N_49127);
or UO_381 (O_381,N_48044,N_47595);
and UO_382 (O_382,N_48431,N_49636);
and UO_383 (O_383,N_47601,N_48796);
xor UO_384 (O_384,N_49830,N_49282);
and UO_385 (O_385,N_49466,N_48325);
xor UO_386 (O_386,N_47938,N_48696);
or UO_387 (O_387,N_49022,N_49320);
and UO_388 (O_388,N_47548,N_47846);
nand UO_389 (O_389,N_49930,N_49430);
nand UO_390 (O_390,N_47914,N_49226);
nor UO_391 (O_391,N_47515,N_48942);
and UO_392 (O_392,N_49088,N_48742);
xor UO_393 (O_393,N_48184,N_47552);
nor UO_394 (O_394,N_49154,N_49912);
or UO_395 (O_395,N_47793,N_48619);
nor UO_396 (O_396,N_47693,N_49683);
nand UO_397 (O_397,N_49103,N_48705);
nand UO_398 (O_398,N_49166,N_49829);
and UO_399 (O_399,N_49333,N_49595);
and UO_400 (O_400,N_48656,N_48241);
or UO_401 (O_401,N_48357,N_48961);
and UO_402 (O_402,N_48292,N_48105);
nor UO_403 (O_403,N_48294,N_49206);
xor UO_404 (O_404,N_48398,N_49573);
and UO_405 (O_405,N_48007,N_49410);
nand UO_406 (O_406,N_49364,N_48630);
nor UO_407 (O_407,N_49586,N_47912);
nand UO_408 (O_408,N_47586,N_49750);
or UO_409 (O_409,N_47962,N_49345);
nor UO_410 (O_410,N_47526,N_48681);
nor UO_411 (O_411,N_49456,N_48445);
nor UO_412 (O_412,N_48020,N_49886);
nand UO_413 (O_413,N_48250,N_48751);
xnor UO_414 (O_414,N_48085,N_47532);
and UO_415 (O_415,N_49231,N_47823);
nand UO_416 (O_416,N_47799,N_48396);
xor UO_417 (O_417,N_48925,N_49518);
xnor UO_418 (O_418,N_49051,N_49649);
nand UO_419 (O_419,N_48955,N_47812);
nand UO_420 (O_420,N_47730,N_49921);
and UO_421 (O_421,N_47545,N_47720);
nor UO_422 (O_422,N_49876,N_49386);
xnor UO_423 (O_423,N_49352,N_48649);
xnor UO_424 (O_424,N_48879,N_48807);
or UO_425 (O_425,N_49531,N_49276);
nand UO_426 (O_426,N_48386,N_47565);
and UO_427 (O_427,N_49630,N_47615);
and UO_428 (O_428,N_49707,N_48877);
nor UO_429 (O_429,N_48424,N_48491);
or UO_430 (O_430,N_48466,N_48433);
nand UO_431 (O_431,N_47952,N_49125);
xor UO_432 (O_432,N_48956,N_48391);
or UO_433 (O_433,N_49863,N_49387);
nand UO_434 (O_434,N_49112,N_47994);
nand UO_435 (O_435,N_48525,N_49004);
nand UO_436 (O_436,N_48197,N_48301);
nand UO_437 (O_437,N_48224,N_48149);
or UO_438 (O_438,N_47619,N_49052);
nor UO_439 (O_439,N_48820,N_49418);
nor UO_440 (O_440,N_49985,N_47714);
and UO_441 (O_441,N_48595,N_49486);
nor UO_442 (O_442,N_47729,N_47747);
xor UO_443 (O_443,N_48772,N_49884);
nor UO_444 (O_444,N_47543,N_48582);
nand UO_445 (O_445,N_47897,N_49106);
nand UO_446 (O_446,N_48056,N_49102);
or UO_447 (O_447,N_49745,N_49176);
nand UO_448 (O_448,N_48565,N_49604);
nand UO_449 (O_449,N_48626,N_48699);
or UO_450 (O_450,N_48232,N_47514);
or UO_451 (O_451,N_49272,N_47879);
xor UO_452 (O_452,N_47659,N_48369);
or UO_453 (O_453,N_48998,N_49903);
or UO_454 (O_454,N_49266,N_48010);
nand UO_455 (O_455,N_49043,N_48011);
xor UO_456 (O_456,N_47834,N_48518);
nor UO_457 (O_457,N_48081,N_49218);
or UO_458 (O_458,N_49860,N_49285);
xor UO_459 (O_459,N_49417,N_49965);
nand UO_460 (O_460,N_49480,N_49819);
nand UO_461 (O_461,N_48305,N_49592);
nand UO_462 (O_462,N_49686,N_47770);
nand UO_463 (O_463,N_49442,N_48471);
xnor UO_464 (O_464,N_48427,N_49704);
nand UO_465 (O_465,N_49271,N_47920);
nand UO_466 (O_466,N_48627,N_49085);
nor UO_467 (O_467,N_48144,N_49215);
and UO_468 (O_468,N_49062,N_48032);
nor UO_469 (O_469,N_48585,N_48264);
and UO_470 (O_470,N_48320,N_49501);
nand UO_471 (O_471,N_48801,N_48330);
or UO_472 (O_472,N_49260,N_48553);
nor UO_473 (O_473,N_47660,N_49096);
nor UO_474 (O_474,N_49347,N_47987);
nand UO_475 (O_475,N_49249,N_48260);
xor UO_476 (O_476,N_48088,N_47765);
or UO_477 (O_477,N_49150,N_47763);
nor UO_478 (O_478,N_49723,N_49899);
nand UO_479 (O_479,N_49419,N_48186);
nor UO_480 (O_480,N_49599,N_47531);
and UO_481 (O_481,N_49255,N_49280);
or UO_482 (O_482,N_48816,N_48784);
xor UO_483 (O_483,N_48557,N_47647);
or UO_484 (O_484,N_49494,N_49329);
xnor UO_485 (O_485,N_49848,N_49458);
or UO_486 (O_486,N_48293,N_49013);
and UO_487 (O_487,N_48947,N_49596);
and UO_488 (O_488,N_49485,N_48139);
or UO_489 (O_489,N_47764,N_47886);
xnor UO_490 (O_490,N_47923,N_47733);
nor UO_491 (O_491,N_48049,N_49933);
or UO_492 (O_492,N_48452,N_48840);
or UO_493 (O_493,N_48533,N_47894);
nor UO_494 (O_494,N_49928,N_49740);
or UO_495 (O_495,N_49190,N_48953);
nand UO_496 (O_496,N_49267,N_49503);
or UO_497 (O_497,N_48124,N_48990);
nor UO_498 (O_498,N_48193,N_47904);
xnor UO_499 (O_499,N_48690,N_48569);
nand UO_500 (O_500,N_49187,N_48024);
nor UO_501 (O_501,N_49135,N_47961);
and UO_502 (O_502,N_48728,N_48542);
nor UO_503 (O_503,N_49789,N_49114);
and UO_504 (O_504,N_48002,N_47608);
or UO_505 (O_505,N_47575,N_49506);
nand UO_506 (O_506,N_49049,N_49427);
and UO_507 (O_507,N_47544,N_47709);
or UO_508 (O_508,N_48819,N_48803);
or UO_509 (O_509,N_49672,N_49944);
and UO_510 (O_510,N_48932,N_47644);
nand UO_511 (O_511,N_48109,N_49339);
or UO_512 (O_512,N_49199,N_49397);
xnor UO_513 (O_513,N_48592,N_49504);
and UO_514 (O_514,N_47696,N_47624);
nor UO_515 (O_515,N_48335,N_49378);
nand UO_516 (O_516,N_48365,N_49362);
nand UO_517 (O_517,N_49960,N_48835);
nor UO_518 (O_518,N_48132,N_47872);
nand UO_519 (O_519,N_48817,N_48298);
nand UO_520 (O_520,N_49845,N_49437);
or UO_521 (O_521,N_47568,N_48997);
and UO_522 (O_522,N_48795,N_47771);
nor UO_523 (O_523,N_48622,N_48809);
nand UO_524 (O_524,N_48324,N_49039);
nand UO_525 (O_525,N_48950,N_48450);
or UO_526 (O_526,N_48885,N_47744);
xnor UO_527 (O_527,N_47628,N_48364);
or UO_528 (O_528,N_49483,N_48984);
and UO_529 (O_529,N_49156,N_48806);
nor UO_530 (O_530,N_49047,N_48637);
nand UO_531 (O_531,N_49978,N_49349);
xnor UO_532 (O_532,N_49321,N_49283);
nor UO_533 (O_533,N_47641,N_49337);
nor UO_534 (O_534,N_47887,N_47895);
xnor UO_535 (O_535,N_49076,N_48559);
and UO_536 (O_536,N_48931,N_49140);
nand UO_537 (O_537,N_49718,N_49195);
nand UO_538 (O_538,N_48739,N_48827);
and UO_539 (O_539,N_48849,N_48952);
nand UO_540 (O_540,N_48832,N_49659);
and UO_541 (O_541,N_49720,N_47676);
nand UO_542 (O_542,N_48494,N_49530);
and UO_543 (O_543,N_47603,N_47782);
and UO_544 (O_544,N_48747,N_49877);
and UO_545 (O_545,N_48571,N_48605);
or UO_546 (O_546,N_49493,N_47502);
nand UO_547 (O_547,N_49141,N_47571);
and UO_548 (O_548,N_48837,N_47551);
nor UO_549 (O_549,N_49155,N_47708);
or UO_550 (O_550,N_49385,N_48588);
nor UO_551 (O_551,N_47712,N_47726);
or UO_552 (O_552,N_48484,N_49139);
nand UO_553 (O_553,N_49303,N_48815);
nand UO_554 (O_554,N_47831,N_48161);
nor UO_555 (O_555,N_47989,N_49953);
nor UO_556 (O_556,N_47820,N_48928);
or UO_557 (O_557,N_49369,N_48664);
and UO_558 (O_558,N_49270,N_47574);
or UO_559 (O_559,N_48381,N_49777);
nor UO_560 (O_560,N_48375,N_49165);
nand UO_561 (O_561,N_49988,N_49179);
and UO_562 (O_562,N_48537,N_48672);
or UO_563 (O_563,N_48065,N_48863);
or UO_564 (O_564,N_49461,N_48783);
nor UO_565 (O_565,N_48208,N_48216);
nor UO_566 (O_566,N_49479,N_47721);
and UO_567 (O_567,N_48867,N_48567);
xnor UO_568 (O_568,N_48401,N_47906);
xor UO_569 (O_569,N_49943,N_49295);
xnor UO_570 (O_570,N_49812,N_48621);
xor UO_571 (O_571,N_49502,N_49505);
nand UO_572 (O_572,N_48331,N_48030);
xnor UO_573 (O_573,N_49428,N_49109);
xnor UO_574 (O_574,N_47809,N_48978);
and UO_575 (O_575,N_48901,N_49719);
nor UO_576 (O_576,N_49406,N_48682);
or UO_577 (O_577,N_48001,N_49766);
nor UO_578 (O_578,N_47583,N_49515);
nand UO_579 (O_579,N_47561,N_47579);
and UO_580 (O_580,N_48378,N_49161);
and UO_581 (O_581,N_47988,N_48104);
and UO_582 (O_582,N_48697,N_48066);
nand UO_583 (O_583,N_49920,N_48316);
or UO_584 (O_584,N_49624,N_47703);
nand UO_585 (O_585,N_48736,N_47975);
xor UO_586 (O_586,N_47691,N_48473);
nor UO_587 (O_587,N_48910,N_47891);
xnor UO_588 (O_588,N_49409,N_49443);
or UO_589 (O_589,N_48117,N_48116);
and UO_590 (O_590,N_49580,N_49727);
xor UO_591 (O_591,N_48792,N_49012);
nor UO_592 (O_592,N_48486,N_47839);
xnor UO_593 (O_593,N_48847,N_49888);
and UO_594 (O_594,N_49396,N_48960);
or UO_595 (O_595,N_48640,N_47774);
xor UO_596 (O_596,N_49946,N_48284);
and UO_597 (O_597,N_49834,N_47519);
and UO_598 (O_598,N_47866,N_49399);
nand UO_599 (O_599,N_47993,N_48379);
or UO_600 (O_600,N_49031,N_49265);
nor UO_601 (O_601,N_47755,N_48419);
nand UO_602 (O_602,N_48633,N_48957);
nand UO_603 (O_603,N_47798,N_49327);
and UO_604 (O_604,N_48848,N_49431);
and UO_605 (O_605,N_47828,N_48991);
nor UO_606 (O_606,N_48496,N_47681);
nor UO_607 (O_607,N_48258,N_48259);
and UO_608 (O_608,N_48673,N_48345);
xor UO_609 (O_609,N_47796,N_48688);
nor UO_610 (O_610,N_47880,N_49350);
or UO_611 (O_611,N_48115,N_48000);
and UO_612 (O_612,N_49587,N_49180);
or UO_613 (O_613,N_48902,N_49142);
and UO_614 (O_614,N_49236,N_48926);
and UO_615 (O_615,N_48711,N_48380);
nand UO_616 (O_616,N_49209,N_48610);
and UO_617 (O_617,N_49548,N_47567);
and UO_618 (O_618,N_48393,N_47968);
xor UO_619 (O_619,N_49296,N_48474);
xnor UO_620 (O_620,N_48915,N_48153);
and UO_621 (O_621,N_49887,N_48449);
and UO_622 (O_622,N_49542,N_49778);
nand UO_623 (O_623,N_49090,N_48740);
nor UO_624 (O_624,N_49619,N_47881);
nor UO_625 (O_625,N_49758,N_49612);
nand UO_626 (O_626,N_48799,N_48476);
nand UO_627 (O_627,N_48265,N_48886);
nor UO_628 (O_628,N_48489,N_48787);
or UO_629 (O_629,N_48935,N_48989);
nand UO_630 (O_630,N_49099,N_48108);
and UO_631 (O_631,N_47580,N_49221);
or UO_632 (O_632,N_49121,N_48600);
and UO_633 (O_633,N_48314,N_48481);
nor UO_634 (O_634,N_48438,N_48061);
xor UO_635 (O_635,N_49684,N_48624);
or UO_636 (O_636,N_47844,N_47892);
and UO_637 (O_637,N_48749,N_47947);
and UO_638 (O_638,N_49259,N_49143);
and UO_639 (O_639,N_49123,N_48866);
and UO_640 (O_640,N_48212,N_47958);
nor UO_641 (O_641,N_49571,N_49737);
or UO_642 (O_642,N_48584,N_48435);
nor UO_643 (O_643,N_48256,N_47687);
or UO_644 (O_644,N_47750,N_47919);
nand UO_645 (O_645,N_48665,N_47666);
and UO_646 (O_646,N_49873,N_49572);
and UO_647 (O_647,N_49436,N_48899);
xor UO_648 (O_648,N_49621,N_48572);
or UO_649 (O_649,N_48601,N_49855);
nand UO_650 (O_650,N_48421,N_49398);
and UO_651 (O_651,N_49762,N_48200);
or UO_652 (O_652,N_48683,N_48541);
or UO_653 (O_653,N_48225,N_47801);
nand UO_654 (O_654,N_47835,N_48703);
or UO_655 (O_655,N_48018,N_49310);
and UO_656 (O_656,N_48222,N_49680);
or UO_657 (O_657,N_49324,N_48448);
or UO_658 (O_658,N_48287,N_47873);
xor UO_659 (O_659,N_49290,N_48169);
nor UO_660 (O_660,N_48490,N_48039);
and UO_661 (O_661,N_47569,N_49289);
xor UO_662 (O_662,N_48833,N_48239);
or UO_663 (O_663,N_49952,N_49101);
and UO_664 (O_664,N_47888,N_49825);
nor UO_665 (O_665,N_48077,N_48826);
nor UO_666 (O_666,N_49185,N_48838);
or UO_667 (O_667,N_48411,N_48986);
nand UO_668 (O_668,N_47786,N_47965);
nor UO_669 (O_669,N_48607,N_47974);
and UO_670 (O_670,N_49709,N_48521);
nand UO_671 (O_671,N_49716,N_48517);
nand UO_672 (O_672,N_48150,N_48552);
nor UO_673 (O_673,N_47890,N_47859);
nor UO_674 (O_674,N_47536,N_49871);
nand UO_675 (O_675,N_47596,N_48423);
nand UO_676 (O_676,N_49790,N_47704);
or UO_677 (O_677,N_49186,N_49644);
nor UO_678 (O_678,N_49175,N_47753);
and UO_679 (O_679,N_49785,N_48387);
nor UO_680 (O_680,N_48719,N_49764);
or UO_681 (O_681,N_48162,N_48236);
xnor UO_682 (O_682,N_48237,N_47985);
or UO_683 (O_683,N_48407,N_49414);
xor UO_684 (O_684,N_48954,N_47651);
or UO_685 (O_685,N_49824,N_48850);
xnor UO_686 (O_686,N_48447,N_48326);
nor UO_687 (O_687,N_49210,N_49747);
and UO_688 (O_688,N_48574,N_49392);
nand UO_689 (O_689,N_48123,N_48913);
nand UO_690 (O_690,N_49207,N_48475);
and UO_691 (O_691,N_47983,N_49582);
or UO_692 (O_692,N_49763,N_49800);
or UO_693 (O_693,N_48687,N_47902);
nor UO_694 (O_694,N_48045,N_47675);
nand UO_695 (O_695,N_49841,N_48203);
nand UO_696 (O_696,N_49229,N_47503);
nand UO_697 (O_697,N_48924,N_48972);
nand UO_698 (O_698,N_47538,N_48130);
nand UO_699 (O_699,N_49524,N_48999);
nor UO_700 (O_700,N_48036,N_49371);
and UO_701 (O_701,N_49691,N_49402);
and UO_702 (O_702,N_49212,N_48464);
xnor UO_703 (O_703,N_48353,N_48503);
xor UO_704 (O_704,N_48372,N_48446);
nor UO_705 (O_705,N_49654,N_48090);
and UO_706 (O_706,N_47611,N_49781);
and UO_707 (O_707,N_49667,N_48046);
or UO_708 (O_708,N_48577,N_48154);
and UO_709 (O_709,N_48625,N_48727);
nand UO_710 (O_710,N_48921,N_48934);
or UO_711 (O_711,N_49446,N_47618);
and UO_712 (O_712,N_49089,N_47723);
or UO_713 (O_713,N_47921,N_49514);
or UO_714 (O_714,N_48566,N_48479);
and UO_715 (O_715,N_49540,N_49311);
nor UO_716 (O_716,N_47540,N_48887);
nand UO_717 (O_717,N_48270,N_47903);
nand UO_718 (O_718,N_49713,N_49157);
and UO_719 (O_719,N_49200,N_48263);
and UO_720 (O_720,N_47524,N_48410);
nor UO_721 (O_721,N_48460,N_48415);
nand UO_722 (O_722,N_49925,N_48893);
or UO_723 (O_723,N_49999,N_48230);
and UO_724 (O_724,N_49366,N_49471);
and UO_725 (O_725,N_49544,N_48892);
nand UO_726 (O_726,N_47736,N_47505);
and UO_727 (O_727,N_47673,N_48764);
or UO_728 (O_728,N_49561,N_49971);
and UO_729 (O_729,N_48135,N_48016);
xor UO_730 (O_730,N_49591,N_48159);
and UO_731 (O_731,N_48068,N_48923);
nand UO_732 (O_732,N_48543,N_49465);
nand UO_733 (O_733,N_47707,N_49975);
nor UO_734 (O_734,N_48884,N_47775);
nand UO_735 (O_735,N_48513,N_49317);
or UO_736 (O_736,N_49351,N_49662);
and UO_737 (O_737,N_47998,N_47701);
or UO_738 (O_738,N_49393,N_47769);
nand UO_739 (O_739,N_49019,N_49291);
nor UO_740 (O_740,N_48125,N_49381);
nand UO_741 (O_741,N_48070,N_49706);
and UO_742 (O_742,N_48857,N_48422);
and UO_743 (O_743,N_48734,N_48738);
xnor UO_744 (O_744,N_48951,N_47797);
or UO_745 (O_745,N_47778,N_48785);
nand UO_746 (O_746,N_48114,N_48793);
and UO_747 (O_747,N_48166,N_47984);
and UO_748 (O_748,N_49227,N_48786);
and UO_749 (O_749,N_48205,N_47950);
and UO_750 (O_750,N_48788,N_49752);
xnor UO_751 (O_751,N_49589,N_48958);
and UO_752 (O_752,N_48701,N_49641);
or UO_753 (O_753,N_49205,N_48430);
and UO_754 (O_754,N_47899,N_47697);
or UO_755 (O_755,N_47625,N_48062);
nor UO_756 (O_756,N_49372,N_49839);
or UO_757 (O_757,N_47665,N_49070);
nor UO_758 (O_758,N_47874,N_47715);
and UO_759 (O_759,N_47559,N_47740);
or UO_760 (O_760,N_49228,N_49628);
and UO_761 (O_761,N_49130,N_48971);
xnor UO_762 (O_762,N_48779,N_48303);
and UO_763 (O_763,N_48187,N_48708);
nand UO_764 (O_764,N_49793,N_47572);
xnor UO_765 (O_765,N_49128,N_48532);
and UO_766 (O_766,N_48830,N_49783);
xor UO_767 (O_767,N_49674,N_48508);
nand UO_768 (O_768,N_47549,N_48285);
nor UO_769 (O_769,N_49001,N_47960);
xor UO_770 (O_770,N_48797,N_49086);
and UO_771 (O_771,N_49058,N_49832);
and UO_772 (O_772,N_48965,N_49015);
nand UO_773 (O_773,N_47954,N_49668);
nor UO_774 (O_774,N_47591,N_47811);
or UO_775 (O_775,N_49722,N_47845);
nand UO_776 (O_776,N_49244,N_47805);
nor UO_777 (O_777,N_48454,N_48385);
nand UO_778 (O_778,N_49846,N_49507);
xnor UO_779 (O_779,N_48199,N_49332);
or UO_780 (O_780,N_47838,N_49474);
or UO_781 (O_781,N_47646,N_49565);
nand UO_782 (O_782,N_49875,N_48706);
or UO_783 (O_783,N_49681,N_49269);
and UO_784 (O_784,N_48670,N_47909);
or UO_785 (O_785,N_47868,N_47678);
or UO_786 (O_786,N_49625,N_48882);
nor UO_787 (O_787,N_48098,N_47534);
nand UO_788 (O_788,N_47995,N_48403);
nand UO_789 (O_789,N_49512,N_48442);
nand UO_790 (O_790,N_48281,N_49898);
or UO_791 (O_791,N_48086,N_48822);
nor UO_792 (O_792,N_49568,N_48941);
or UO_793 (O_793,N_49676,N_49938);
or UO_794 (O_794,N_48723,N_49756);
xnor UO_795 (O_795,N_48278,N_49323);
nand UO_796 (O_796,N_49281,N_47842);
or UO_797 (O_797,N_49951,N_48547);
xor UO_798 (O_798,N_48405,N_49278);
xnor UO_799 (O_799,N_48616,N_49803);
xor UO_800 (O_800,N_47621,N_49867);
nor UO_801 (O_801,N_47656,N_47945);
and UO_802 (O_802,N_48283,N_49254);
or UO_803 (O_803,N_49959,N_47558);
and UO_804 (O_804,N_47857,N_49304);
xor UO_805 (O_805,N_49253,N_48671);
nor UO_806 (O_806,N_47777,N_47915);
or UO_807 (O_807,N_47943,N_49605);
xor UO_808 (O_808,N_47822,N_49967);
nand UO_809 (O_809,N_49330,N_49854);
and UO_810 (O_810,N_48562,N_47814);
or UO_811 (O_811,N_49305,N_49225);
xor UO_812 (O_812,N_49251,N_48608);
and UO_813 (O_813,N_47936,N_47926);
xnor UO_814 (O_814,N_49214,N_49726);
nor UO_815 (O_815,N_48254,N_47967);
nand UO_816 (O_816,N_49508,N_47849);
or UO_817 (O_817,N_48118,N_47794);
nand UO_818 (O_818,N_47739,N_48805);
xor UO_819 (O_819,N_49500,N_49626);
or UO_820 (O_820,N_49360,N_49652);
nand UO_821 (O_821,N_49661,N_49741);
or UO_822 (O_822,N_47959,N_48226);
nor UO_823 (O_823,N_47680,N_48648);
nor UO_824 (O_824,N_48906,N_48842);
xnor UO_825 (O_825,N_49453,N_49455);
nand UO_826 (O_826,N_47662,N_49433);
and UO_827 (O_827,N_49593,N_47896);
xnor UO_828 (O_828,N_49950,N_49693);
and UO_829 (O_829,N_48889,N_49098);
nor UO_830 (O_830,N_49367,N_48458);
and UO_831 (O_831,N_47670,N_49211);
or UO_832 (O_832,N_49346,N_49736);
nand UO_833 (O_833,N_47875,N_47539);
or UO_834 (O_834,N_49984,N_48578);
nor UO_835 (O_835,N_49697,N_48979);
xnor UO_836 (O_836,N_49484,N_47682);
nor UO_837 (O_837,N_49913,N_49084);
or UO_838 (O_838,N_49491,N_49056);
nand UO_839 (O_839,N_49234,N_48038);
xnor UO_840 (O_840,N_48636,N_47664);
and UO_841 (O_841,N_48196,N_48371);
and UO_842 (O_842,N_49273,N_48389);
or UO_843 (O_843,N_48617,N_48526);
or UO_844 (O_844,N_49467,N_48726);
xor UO_845 (O_845,N_48642,N_47986);
nor UO_846 (O_846,N_48659,N_49029);
or UO_847 (O_847,N_48861,N_49669);
and UO_848 (O_848,N_47511,N_48352);
and UO_849 (O_849,N_48094,N_49473);
and UO_850 (O_850,N_48076,N_48444);
nand UO_851 (O_851,N_49334,N_48929);
nand UO_852 (O_852,N_47754,N_47748);
nand UO_853 (O_853,N_47953,N_48048);
xor UO_854 (O_854,N_49557,N_48523);
and UO_855 (O_855,N_49383,N_49404);
and UO_856 (O_856,N_48883,N_48660);
xnor UO_857 (O_857,N_48127,N_48692);
or UO_858 (O_858,N_47533,N_49805);
and UO_859 (O_859,N_48629,N_48388);
nor UO_860 (O_860,N_49787,N_49962);
nor UO_861 (O_861,N_49532,N_49147);
or UO_862 (O_862,N_49118,N_49390);
nand UO_863 (O_863,N_48667,N_48439);
or UO_864 (O_864,N_49773,N_48903);
and UO_865 (O_865,N_49262,N_49638);
nor UO_866 (O_866,N_48434,N_49377);
and UO_867 (O_867,N_49627,N_48091);
nor UO_868 (O_868,N_47626,N_47843);
nor UO_869 (O_869,N_47639,N_48413);
or UO_870 (O_870,N_48996,N_49564);
nor UO_871 (O_871,N_49692,N_47853);
nor UO_872 (O_872,N_49734,N_47612);
or UO_873 (O_873,N_49569,N_49032);
nor UO_874 (O_874,N_47728,N_47645);
nand UO_875 (O_875,N_48133,N_48911);
and UO_876 (O_876,N_48373,N_48639);
or UO_877 (O_877,N_48215,N_48504);
and UO_878 (O_878,N_48561,N_48168);
or UO_879 (O_879,N_49240,N_49037);
and UO_880 (O_880,N_47717,N_48231);
xor UO_881 (O_881,N_48367,N_49432);
and UO_882 (O_882,N_49482,N_47946);
nor UO_883 (O_883,N_48500,N_49629);
xor UO_884 (O_884,N_48975,N_49288);
or UO_885 (O_885,N_49640,N_49008);
xnor UO_886 (O_886,N_49979,N_49878);
or UO_887 (O_887,N_49815,N_49016);
nor UO_888 (O_888,N_48469,N_49094);
and UO_889 (O_889,N_48219,N_49370);
nand UO_890 (O_890,N_49814,N_49423);
nor UO_891 (O_891,N_48905,N_48560);
xnor UO_892 (O_892,N_49203,N_49469);
or UO_893 (O_893,N_48480,N_47854);
and UO_894 (O_894,N_48771,N_49170);
xnor UO_895 (O_895,N_49343,N_49797);
xnor UO_896 (O_896,N_49560,N_48182);
nor UO_897 (O_897,N_48351,N_48789);
or UO_898 (O_898,N_49132,N_49837);
nand UO_899 (O_899,N_47918,N_47512);
nand UO_900 (O_900,N_49355,N_47908);
and UO_901 (O_901,N_49308,N_48871);
or UO_902 (O_902,N_48247,N_48279);
or UO_903 (O_903,N_48404,N_48374);
nand UO_904 (O_904,N_49703,N_49379);
and UO_905 (O_905,N_47649,N_48776);
or UO_906 (O_906,N_48603,N_47913);
nand UO_907 (O_907,N_48535,N_48201);
nand UO_908 (O_908,N_48170,N_47992);
or UO_909 (O_909,N_49614,N_48063);
and UO_910 (O_910,N_48775,N_47674);
or UO_911 (O_911,N_47898,N_49368);
or UO_912 (O_912,N_47773,N_49470);
nand UO_913 (O_913,N_49743,N_49861);
nor UO_914 (O_914,N_47885,N_48918);
nand UO_915 (O_915,N_48308,N_48744);
xnor UO_916 (O_916,N_49000,N_48746);
xor UO_917 (O_917,N_47741,N_47719);
and UO_918 (O_918,N_48355,N_48451);
and UO_919 (O_919,N_47883,N_48509);
nor UO_920 (O_920,N_48810,N_49116);
and UO_921 (O_921,N_48992,N_49551);
nor UO_922 (O_922,N_47802,N_47776);
and UO_923 (O_923,N_48456,N_48643);
and UO_924 (O_924,N_48657,N_49208);
xor UO_925 (O_925,N_47506,N_48165);
or UO_926 (O_926,N_47924,N_48869);
or UO_927 (O_927,N_49911,N_49313);
nand UO_928 (O_928,N_49820,N_47616);
nor UO_929 (O_929,N_48006,N_48158);
xor UO_930 (O_930,N_47861,N_48618);
or UO_931 (O_931,N_48156,N_49986);
or UO_932 (O_932,N_48348,N_48008);
nor UO_933 (O_933,N_47738,N_48936);
or UO_934 (O_934,N_49163,N_49650);
and UO_935 (O_935,N_48558,N_49230);
nor UO_936 (O_936,N_49063,N_49222);
or UO_937 (O_937,N_48053,N_48220);
nand UO_938 (O_938,N_49162,N_49302);
xor UO_939 (O_939,N_47940,N_49949);
xnor UO_940 (O_940,N_48395,N_49721);
and UO_941 (O_941,N_47689,N_47935);
nor UO_942 (O_942,N_49268,N_49219);
nand UO_943 (O_943,N_49120,N_49144);
and UO_944 (O_944,N_48770,N_47516);
and UO_945 (O_945,N_49770,N_48691);
and UO_946 (O_946,N_49816,N_49566);
xor UO_947 (O_947,N_49426,N_49843);
nor UO_948 (O_948,N_48677,N_49618);
xor UO_949 (O_949,N_49376,N_48360);
and UO_950 (O_950,N_47530,N_48704);
nand UO_951 (O_951,N_48868,N_49097);
nor UO_952 (O_952,N_48977,N_47566);
nand UO_953 (O_953,N_49400,N_48507);
nor UO_954 (O_954,N_48399,N_47635);
xor UO_955 (O_955,N_47504,N_49248);
xnor UO_956 (O_956,N_47513,N_49137);
nor UO_957 (O_957,N_48555,N_48145);
nand UO_958 (O_958,N_47592,N_48669);
nor UO_959 (O_959,N_48072,N_48312);
nor UO_960 (O_960,N_49864,N_49600);
and UO_961 (O_961,N_48093,N_48896);
nor UO_962 (O_962,N_47541,N_48390);
xnor UO_963 (O_963,N_49570,N_49994);
xor UO_964 (O_964,N_48880,N_47546);
nand UO_965 (O_965,N_49981,N_47706);
nor UO_966 (O_966,N_48288,N_49010);
nand UO_967 (O_967,N_48080,N_49224);
and UO_968 (O_968,N_48912,N_48420);
nand UO_969 (O_969,N_48730,N_49151);
nand UO_970 (O_970,N_49689,N_47856);
or UO_971 (O_971,N_49312,N_49651);
and UO_972 (O_972,N_48453,N_48598);
nor UO_973 (O_973,N_48993,N_49167);
nand UO_974 (O_974,N_48581,N_49181);
xnor UO_975 (O_975,N_47694,N_49027);
xnor UO_976 (O_976,N_49905,N_47819);
nand UO_977 (O_977,N_49105,N_48470);
and UO_978 (O_978,N_48344,N_48336);
xnor UO_979 (O_979,N_49528,N_49896);
nand UO_980 (O_980,N_48937,N_48812);
xnor UO_981 (O_981,N_49974,N_49492);
and UO_982 (O_982,N_47991,N_47570);
and UO_983 (O_983,N_49620,N_48071);
xor UO_984 (O_984,N_49732,N_49751);
nand UO_985 (O_985,N_48042,N_47617);
nand UO_986 (O_986,N_49160,N_47661);
nand UO_987 (O_987,N_48663,N_49827);
or UO_988 (O_988,N_49817,N_49065);
nor UO_989 (O_989,N_48243,N_49189);
and UO_990 (O_990,N_47725,N_49073);
xnor UO_991 (O_991,N_48914,N_49823);
nand UO_992 (O_992,N_48163,N_48658);
xor UO_993 (O_993,N_49918,N_47783);
or UO_994 (O_994,N_48858,N_49997);
nor UO_995 (O_995,N_47517,N_48089);
nor UO_996 (O_996,N_49421,N_48693);
and UO_997 (O_997,N_47806,N_49174);
nor UO_998 (O_998,N_47716,N_47869);
and UO_999 (O_999,N_49454,N_48321);
or UO_1000 (O_1000,N_49095,N_48768);
nor UO_1001 (O_1001,N_49881,N_47667);
or UO_1002 (O_1002,N_47787,N_49842);
and UO_1003 (O_1003,N_48549,N_49475);
nor UO_1004 (O_1004,N_48146,N_47556);
nor UO_1005 (O_1005,N_47978,N_48823);
and UO_1006 (O_1006,N_48073,N_48137);
or UO_1007 (O_1007,N_47746,N_49113);
xnor UO_1008 (O_1008,N_48271,N_48646);
nor UO_1009 (O_1009,N_49033,N_47560);
and UO_1010 (O_1010,N_48227,N_49481);
or UO_1011 (O_1011,N_48244,N_49357);
xnor UO_1012 (O_1012,N_48377,N_48530);
or UO_1013 (O_1013,N_49194,N_48462);
nand UO_1014 (O_1014,N_47956,N_47999);
xnor UO_1015 (O_1015,N_49577,N_47523);
nand UO_1016 (O_1016,N_49315,N_49018);
and UO_1017 (O_1017,N_49893,N_49519);
and UO_1018 (O_1018,N_48980,N_47522);
or UO_1019 (O_1019,N_48556,N_49907);
xnor UO_1020 (O_1020,N_49444,N_47966);
or UO_1021 (O_1021,N_48966,N_49991);
xnor UO_1022 (O_1022,N_48317,N_48694);
or UO_1023 (O_1023,N_49715,N_49081);
and UO_1024 (O_1024,N_49926,N_49354);
and UO_1025 (O_1025,N_47758,N_49220);
xor UO_1026 (O_1026,N_49993,N_49138);
and UO_1027 (O_1027,N_49937,N_49714);
and UO_1028 (O_1028,N_49598,N_48614);
or UO_1029 (O_1029,N_49794,N_48888);
xor UO_1030 (O_1030,N_48897,N_49647);
and UO_1031 (O_1031,N_48587,N_48087);
xor UO_1032 (O_1032,N_48429,N_49464);
and UO_1033 (O_1033,N_49798,N_49813);
and UO_1034 (O_1034,N_48825,N_48917);
and UO_1035 (O_1035,N_48721,N_49658);
nand UO_1036 (O_1036,N_48028,N_49136);
and UO_1037 (O_1037,N_48720,N_48054);
nor UO_1038 (O_1038,N_49158,N_49761);
xor UO_1039 (O_1039,N_49294,N_48844);
and UO_1040 (O_1040,N_49241,N_49635);
nor UO_1041 (O_1041,N_48511,N_49202);
nor UO_1042 (O_1042,N_49810,N_48009);
xor UO_1043 (O_1043,N_48545,N_47745);
and UO_1044 (O_1044,N_49258,N_49822);
nand UO_1045 (O_1045,N_49754,N_48845);
and UO_1046 (O_1046,N_48864,N_48253);
nand UO_1047 (O_1047,N_49356,N_49359);
nor UO_1048 (O_1048,N_49608,N_49656);
nor UO_1049 (O_1049,N_47939,N_48856);
and UO_1050 (O_1050,N_47867,N_49972);
and UO_1051 (O_1051,N_48843,N_48713);
or UO_1052 (O_1052,N_47718,N_49420);
nand UO_1053 (O_1053,N_49915,N_48564);
nor UO_1054 (O_1054,N_49003,N_47528);
or UO_1055 (O_1055,N_48722,N_49192);
and UO_1056 (O_1056,N_49904,N_47695);
nor UO_1057 (O_1057,N_48339,N_48252);
nor UO_1058 (O_1058,N_47690,N_48350);
xnor UO_1059 (O_1059,N_49438,N_49529);
nand UO_1060 (O_1060,N_49201,N_48528);
xnor UO_1061 (O_1061,N_48436,N_48811);
nand UO_1062 (O_1062,N_48769,N_49739);
and UO_1063 (O_1063,N_49223,N_47652);
or UO_1064 (O_1064,N_48047,N_49341);
nor UO_1065 (O_1065,N_49653,N_48686);
xnor UO_1066 (O_1066,N_47642,N_49771);
and UO_1067 (O_1067,N_48520,N_49866);
or UO_1068 (O_1068,N_47997,N_49395);
nor UO_1069 (O_1069,N_48724,N_48943);
or UO_1070 (O_1070,N_48964,N_48296);
xor UO_1071 (O_1071,N_47829,N_47564);
or UO_1072 (O_1072,N_48919,N_47810);
nand UO_1073 (O_1073,N_49041,N_49172);
xor UO_1074 (O_1074,N_47760,N_48516);
xnor UO_1075 (O_1075,N_49796,N_49859);
and UO_1076 (O_1076,N_48777,N_48361);
or UO_1077 (O_1077,N_47860,N_48554);
xor UO_1078 (O_1078,N_49948,N_48052);
xor UO_1079 (O_1079,N_49322,N_49434);
or UO_1080 (O_1080,N_48628,N_47537);
or UO_1081 (O_1081,N_48743,N_47980);
nand UO_1082 (O_1082,N_47679,N_49213);
nor UO_1083 (O_1083,N_49389,N_49574);
nor UO_1084 (O_1084,N_49581,N_49889);
and UO_1085 (O_1085,N_48194,N_49517);
and UO_1086 (O_1086,N_49936,N_47724);
xor UO_1087 (O_1087,N_49435,N_48408);
nand UO_1088 (O_1088,N_48121,N_47916);
xor UO_1089 (O_1089,N_48641,N_48939);
nor UO_1090 (O_1090,N_47864,N_48698);
nand UO_1091 (O_1091,N_48302,N_49468);
nand UO_1092 (O_1092,N_49375,N_48333);
nand UO_1093 (O_1093,N_48017,N_49472);
nand UO_1094 (O_1094,N_48290,N_47840);
and UO_1095 (O_1095,N_47613,N_49556);
and UO_1096 (O_1096,N_48492,N_49489);
and UO_1097 (O_1097,N_49690,N_49509);
xor UO_1098 (O_1098,N_49968,N_48160);
and UO_1099 (O_1099,N_48141,N_49914);
xnor UO_1100 (O_1100,N_48778,N_49045);
nand UO_1101 (O_1101,N_48909,N_49603);
nor UO_1102 (O_1102,N_48570,N_49559);
or UO_1103 (O_1103,N_48459,N_48262);
xnor UO_1104 (O_1104,N_48878,N_49665);
or UO_1105 (O_1105,N_48818,N_48898);
or UO_1106 (O_1106,N_48180,N_49617);
nand UO_1107 (O_1107,N_49576,N_47951);
xnor UO_1108 (O_1108,N_47602,N_49642);
or UO_1109 (O_1109,N_48631,N_48938);
and UO_1110 (O_1110,N_47807,N_49038);
or UO_1111 (O_1111,N_48059,N_49554);
nand UO_1112 (O_1112,N_49024,N_48908);
nor UO_1113 (O_1113,N_48277,N_48488);
and UO_1114 (O_1114,N_49072,N_47542);
nand UO_1115 (O_1115,N_48907,N_49705);
nand UO_1116 (O_1116,N_48604,N_48829);
xnor UO_1117 (O_1117,N_48457,N_49087);
nor UO_1118 (O_1118,N_47882,N_48970);
or UO_1119 (O_1119,N_47752,N_48948);
and UO_1120 (O_1120,N_49068,N_47852);
nor UO_1121 (O_1121,N_47789,N_49939);
xor UO_1122 (O_1122,N_49552,N_48968);
xnor UO_1123 (O_1123,N_49325,N_49287);
nand UO_1124 (O_1124,N_48359,N_48273);
xnor UO_1125 (O_1125,N_48425,N_48307);
nor UO_1126 (O_1126,N_49264,N_47767);
or UO_1127 (O_1127,N_48874,N_48414);
and UO_1128 (O_1128,N_47521,N_49238);
nand UO_1129 (O_1129,N_47949,N_47508);
nand UO_1130 (O_1130,N_49424,N_49422);
or UO_1131 (O_1131,N_48662,N_49549);
and UO_1132 (O_1132,N_49774,N_49982);
and UO_1133 (O_1133,N_48143,N_49880);
xor UO_1134 (O_1134,N_47996,N_47632);
nor UO_1135 (O_1135,N_48623,N_48502);
xor UO_1136 (O_1136,N_48714,N_49902);
and UO_1137 (O_1137,N_49441,N_49361);
or UO_1138 (O_1138,N_48498,N_49457);
and UO_1139 (O_1139,N_48933,N_47636);
nand UO_1140 (O_1140,N_48440,N_49245);
nand UO_1141 (O_1141,N_48767,N_48495);
nand UO_1142 (O_1142,N_47743,N_48337);
or UO_1143 (O_1143,N_48214,N_49239);
nor UO_1144 (O_1144,N_48718,N_48402);
and UO_1145 (O_1145,N_47735,N_47650);
xor UO_1146 (O_1146,N_48173,N_49537);
nand UO_1147 (O_1147,N_48181,N_49606);
nor UO_1148 (O_1148,N_47766,N_48418);
and UO_1149 (O_1149,N_48463,N_49966);
and UO_1150 (O_1150,N_48356,N_49678);
nand UO_1151 (O_1151,N_49929,N_49527);
nor UO_1152 (O_1152,N_48025,N_49856);
or UO_1153 (O_1153,N_48437,N_48341);
nor UO_1154 (O_1154,N_48946,N_48881);
and UO_1155 (O_1155,N_48140,N_49079);
nand UO_1156 (O_1156,N_49091,N_48286);
nand UO_1157 (O_1157,N_48765,N_47547);
or UO_1158 (O_1158,N_48836,N_47841);
xnor UO_1159 (O_1159,N_49516,N_48735);
nand UO_1160 (O_1160,N_48846,N_47587);
xnor UO_1161 (O_1161,N_49092,N_47963);
nor UO_1162 (O_1162,N_48019,N_49673);
or UO_1163 (O_1163,N_49284,N_47581);
and UO_1164 (O_1164,N_49009,N_48138);
or UO_1165 (O_1165,N_49440,N_48568);
or UO_1166 (O_1166,N_48192,N_48176);
xor UO_1167 (O_1167,N_48268,N_49699);
nand UO_1168 (O_1168,N_49188,N_49806);
xor UO_1169 (O_1169,N_48753,N_49882);
nand UO_1170 (O_1170,N_47900,N_48178);
or UO_1171 (O_1171,N_48043,N_47525);
or UO_1172 (O_1172,N_49054,N_49279);
or UO_1173 (O_1173,N_49535,N_48774);
nand UO_1174 (O_1174,N_47684,N_47710);
and UO_1175 (O_1175,N_48228,N_48136);
xnor UO_1176 (O_1176,N_48257,N_49104);
nand UO_1177 (O_1177,N_47702,N_48467);
or UO_1178 (O_1178,N_47855,N_49663);
nand UO_1179 (O_1179,N_48266,N_48209);
xor UO_1180 (O_1180,N_48737,N_49365);
nor UO_1181 (O_1181,N_48295,N_47520);
xnor UO_1182 (O_1182,N_47742,N_48171);
nand UO_1183 (O_1183,N_47826,N_49257);
nor UO_1184 (O_1184,N_48023,N_49590);
nand UO_1185 (O_1185,N_47800,N_48760);
nand UO_1186 (O_1186,N_47578,N_48655);
or UO_1187 (O_1187,N_47638,N_49833);
and UO_1188 (O_1188,N_48188,N_48332);
xnor UO_1189 (O_1189,N_48443,N_47901);
xor UO_1190 (O_1190,N_47593,N_48675);
and UO_1191 (O_1191,N_48100,N_49890);
or UO_1192 (O_1192,N_49318,N_49080);
and UO_1193 (O_1193,N_49538,N_49865);
and UO_1194 (O_1194,N_48611,N_47751);
nor UO_1195 (O_1195,N_48967,N_49462);
and UO_1196 (O_1196,N_49807,N_47871);
and UO_1197 (O_1197,N_49064,N_49687);
or UO_1198 (O_1198,N_49025,N_47535);
nor UO_1199 (O_1199,N_48300,N_48875);
nand UO_1200 (O_1200,N_49307,N_48731);
and UO_1201 (O_1201,N_49416,N_49061);
or UO_1202 (O_1202,N_48198,N_48904);
nand UO_1203 (O_1203,N_47518,N_48602);
and UO_1204 (O_1204,N_48347,N_47606);
nand UO_1205 (O_1205,N_49728,N_48791);
or UO_1206 (O_1206,N_48780,N_49977);
and UO_1207 (O_1207,N_48725,N_49637);
nor UO_1208 (O_1208,N_49452,N_49394);
xor UO_1209 (O_1209,N_48551,N_48676);
nor UO_1210 (O_1210,N_47672,N_49786);
or UO_1211 (O_1211,N_47653,N_48831);
nand UO_1212 (O_1212,N_48594,N_47553);
xnor UO_1213 (O_1213,N_48763,N_49712);
nor UO_1214 (O_1214,N_49168,N_47785);
xnor UO_1215 (O_1215,N_48609,N_48539);
xnor UO_1216 (O_1216,N_47722,N_48416);
xnor UO_1217 (O_1217,N_49731,N_49613);
xnor UO_1218 (O_1218,N_48752,N_47576);
or UO_1219 (O_1219,N_49964,N_49811);
xnor UO_1220 (O_1220,N_47830,N_49382);
xor UO_1221 (O_1221,N_48748,N_48174);
or UO_1222 (O_1222,N_49730,N_48083);
nand UO_1223 (O_1223,N_47878,N_48095);
nand UO_1224 (O_1224,N_49216,N_48274);
xor UO_1225 (O_1225,N_48766,N_49036);
and UO_1226 (O_1226,N_48055,N_49256);
nor UO_1227 (O_1227,N_47607,N_49028);
xor UO_1228 (O_1228,N_49594,N_47925);
nor UO_1229 (O_1229,N_47573,N_48580);
nor UO_1230 (O_1230,N_48235,N_47970);
nand UO_1231 (O_1231,N_49100,N_48538);
or UO_1232 (O_1232,N_48851,N_48041);
nor UO_1233 (O_1233,N_49020,N_48428);
or UO_1234 (O_1234,N_47555,N_49388);
nand UO_1235 (O_1235,N_49030,N_49055);
nand UO_1236 (O_1236,N_49017,N_47877);
nor UO_1237 (O_1237,N_47928,N_48586);
or UO_1238 (O_1238,N_49700,N_48057);
nor UO_1239 (O_1239,N_49597,N_49802);
and UO_1240 (O_1240,N_48741,N_48644);
or UO_1241 (O_1241,N_49060,N_49237);
nand UO_1242 (O_1242,N_48304,N_49799);
xor UO_1243 (O_1243,N_49184,N_49035);
xnor UO_1244 (O_1244,N_49107,N_49634);
or UO_1245 (O_1245,N_48755,N_49894);
and UO_1246 (O_1246,N_47944,N_49776);
nor UO_1247 (O_1247,N_47981,N_48983);
or UO_1248 (O_1248,N_49755,N_49173);
xnor UO_1249 (O_1249,N_49748,N_49119);
and UO_1250 (O_1250,N_48403,N_49419);
xnor UO_1251 (O_1251,N_49057,N_49094);
and UO_1252 (O_1252,N_47713,N_47805);
nor UO_1253 (O_1253,N_47698,N_47727);
xnor UO_1254 (O_1254,N_48516,N_48864);
xor UO_1255 (O_1255,N_47874,N_48996);
or UO_1256 (O_1256,N_48057,N_47514);
nor UO_1257 (O_1257,N_47550,N_48358);
and UO_1258 (O_1258,N_49985,N_48118);
nand UO_1259 (O_1259,N_49653,N_49325);
nor UO_1260 (O_1260,N_49193,N_48788);
nand UO_1261 (O_1261,N_48611,N_49501);
xor UO_1262 (O_1262,N_49907,N_48345);
nand UO_1263 (O_1263,N_48730,N_48936);
nand UO_1264 (O_1264,N_49043,N_48191);
nor UO_1265 (O_1265,N_49214,N_49926);
or UO_1266 (O_1266,N_48529,N_48794);
xor UO_1267 (O_1267,N_48169,N_49225);
or UO_1268 (O_1268,N_48084,N_48232);
and UO_1269 (O_1269,N_47509,N_48484);
nand UO_1270 (O_1270,N_48483,N_48973);
and UO_1271 (O_1271,N_49740,N_49519);
xor UO_1272 (O_1272,N_48716,N_49286);
or UO_1273 (O_1273,N_49177,N_49599);
or UO_1274 (O_1274,N_48552,N_48937);
and UO_1275 (O_1275,N_48305,N_48065);
or UO_1276 (O_1276,N_48964,N_49041);
xor UO_1277 (O_1277,N_49797,N_47850);
or UO_1278 (O_1278,N_48573,N_48988);
or UO_1279 (O_1279,N_47812,N_48156);
or UO_1280 (O_1280,N_47743,N_48778);
nand UO_1281 (O_1281,N_49585,N_47646);
nor UO_1282 (O_1282,N_47891,N_47824);
or UO_1283 (O_1283,N_49573,N_49222);
or UO_1284 (O_1284,N_48032,N_48083);
and UO_1285 (O_1285,N_49582,N_47690);
or UO_1286 (O_1286,N_49666,N_49454);
and UO_1287 (O_1287,N_48647,N_48970);
and UO_1288 (O_1288,N_48654,N_48138);
nand UO_1289 (O_1289,N_48011,N_48021);
xor UO_1290 (O_1290,N_49304,N_47560);
nand UO_1291 (O_1291,N_49495,N_48788);
nor UO_1292 (O_1292,N_48992,N_48659);
nand UO_1293 (O_1293,N_49246,N_49821);
nand UO_1294 (O_1294,N_47944,N_49146);
nor UO_1295 (O_1295,N_48755,N_48631);
nand UO_1296 (O_1296,N_48442,N_49260);
nand UO_1297 (O_1297,N_49742,N_49503);
or UO_1298 (O_1298,N_49116,N_49149);
nor UO_1299 (O_1299,N_49659,N_49856);
nor UO_1300 (O_1300,N_49513,N_48630);
and UO_1301 (O_1301,N_48644,N_48453);
and UO_1302 (O_1302,N_48749,N_49727);
and UO_1303 (O_1303,N_48703,N_47947);
or UO_1304 (O_1304,N_49395,N_48242);
nor UO_1305 (O_1305,N_47770,N_47543);
and UO_1306 (O_1306,N_48144,N_48306);
nor UO_1307 (O_1307,N_48689,N_49976);
nand UO_1308 (O_1308,N_48220,N_49762);
and UO_1309 (O_1309,N_49435,N_48596);
nor UO_1310 (O_1310,N_48915,N_48557);
and UO_1311 (O_1311,N_49909,N_49350);
or UO_1312 (O_1312,N_48265,N_48463);
nand UO_1313 (O_1313,N_48487,N_48129);
xnor UO_1314 (O_1314,N_47903,N_49538);
nand UO_1315 (O_1315,N_47621,N_47631);
xnor UO_1316 (O_1316,N_48332,N_49481);
nor UO_1317 (O_1317,N_47965,N_49528);
nor UO_1318 (O_1318,N_47645,N_48318);
or UO_1319 (O_1319,N_49529,N_47836);
nand UO_1320 (O_1320,N_47842,N_47665);
nand UO_1321 (O_1321,N_47993,N_49347);
nand UO_1322 (O_1322,N_48209,N_49984);
nand UO_1323 (O_1323,N_47714,N_48651);
and UO_1324 (O_1324,N_48358,N_49645);
or UO_1325 (O_1325,N_48413,N_49230);
xnor UO_1326 (O_1326,N_48525,N_49078);
xor UO_1327 (O_1327,N_49449,N_47885);
and UO_1328 (O_1328,N_48531,N_49933);
and UO_1329 (O_1329,N_48318,N_47928);
nor UO_1330 (O_1330,N_49455,N_48233);
xnor UO_1331 (O_1331,N_47581,N_47964);
or UO_1332 (O_1332,N_48517,N_48237);
nor UO_1333 (O_1333,N_48924,N_49653);
xnor UO_1334 (O_1334,N_47920,N_48159);
and UO_1335 (O_1335,N_47968,N_49155);
nand UO_1336 (O_1336,N_49101,N_49991);
nor UO_1337 (O_1337,N_49270,N_49892);
nor UO_1338 (O_1338,N_48658,N_48061);
xnor UO_1339 (O_1339,N_48094,N_49583);
xor UO_1340 (O_1340,N_48936,N_49698);
xnor UO_1341 (O_1341,N_48686,N_48159);
nand UO_1342 (O_1342,N_49836,N_47726);
nor UO_1343 (O_1343,N_48800,N_49003);
nor UO_1344 (O_1344,N_49156,N_48486);
nor UO_1345 (O_1345,N_48174,N_48701);
and UO_1346 (O_1346,N_48388,N_48979);
or UO_1347 (O_1347,N_49406,N_49213);
nor UO_1348 (O_1348,N_49412,N_48222);
xor UO_1349 (O_1349,N_48935,N_48081);
and UO_1350 (O_1350,N_49586,N_48373);
and UO_1351 (O_1351,N_49196,N_47609);
and UO_1352 (O_1352,N_49247,N_49822);
xnor UO_1353 (O_1353,N_48284,N_49234);
and UO_1354 (O_1354,N_49204,N_48644);
nor UO_1355 (O_1355,N_48929,N_47964);
nor UO_1356 (O_1356,N_49024,N_47959);
or UO_1357 (O_1357,N_49634,N_48160);
or UO_1358 (O_1358,N_47943,N_49022);
and UO_1359 (O_1359,N_49239,N_47861);
nor UO_1360 (O_1360,N_49431,N_49887);
nor UO_1361 (O_1361,N_49912,N_49942);
and UO_1362 (O_1362,N_49480,N_49254);
nand UO_1363 (O_1363,N_48250,N_49517);
nand UO_1364 (O_1364,N_48132,N_47989);
xnor UO_1365 (O_1365,N_48770,N_49406);
or UO_1366 (O_1366,N_47586,N_48693);
and UO_1367 (O_1367,N_47740,N_49770);
and UO_1368 (O_1368,N_48597,N_49291);
nand UO_1369 (O_1369,N_47531,N_48344);
nor UO_1370 (O_1370,N_48578,N_49255);
or UO_1371 (O_1371,N_47590,N_47660);
nor UO_1372 (O_1372,N_48278,N_48010);
and UO_1373 (O_1373,N_48059,N_47977);
or UO_1374 (O_1374,N_48608,N_49909);
and UO_1375 (O_1375,N_47870,N_48390);
xnor UO_1376 (O_1376,N_49488,N_48662);
nor UO_1377 (O_1377,N_49736,N_48823);
nor UO_1378 (O_1378,N_48496,N_48884);
or UO_1379 (O_1379,N_48157,N_49480);
or UO_1380 (O_1380,N_48584,N_49237);
and UO_1381 (O_1381,N_49879,N_49109);
and UO_1382 (O_1382,N_49529,N_49175);
xnor UO_1383 (O_1383,N_47834,N_49973);
xnor UO_1384 (O_1384,N_48361,N_48949);
xor UO_1385 (O_1385,N_49039,N_47653);
xnor UO_1386 (O_1386,N_49012,N_48284);
and UO_1387 (O_1387,N_47708,N_47532);
or UO_1388 (O_1388,N_48734,N_49332);
or UO_1389 (O_1389,N_49833,N_49134);
or UO_1390 (O_1390,N_49115,N_49996);
and UO_1391 (O_1391,N_49353,N_48487);
or UO_1392 (O_1392,N_49254,N_49415);
nand UO_1393 (O_1393,N_48573,N_48672);
xnor UO_1394 (O_1394,N_48170,N_47763);
and UO_1395 (O_1395,N_48940,N_48179);
xor UO_1396 (O_1396,N_48751,N_48080);
and UO_1397 (O_1397,N_48220,N_49600);
and UO_1398 (O_1398,N_48816,N_48326);
and UO_1399 (O_1399,N_49534,N_48436);
nor UO_1400 (O_1400,N_47712,N_48017);
xnor UO_1401 (O_1401,N_47914,N_47572);
and UO_1402 (O_1402,N_49362,N_48783);
nand UO_1403 (O_1403,N_47742,N_47643);
nand UO_1404 (O_1404,N_48667,N_47998);
nor UO_1405 (O_1405,N_48933,N_48279);
or UO_1406 (O_1406,N_47661,N_48389);
or UO_1407 (O_1407,N_47976,N_47550);
xor UO_1408 (O_1408,N_48004,N_47627);
and UO_1409 (O_1409,N_49602,N_49087);
or UO_1410 (O_1410,N_48885,N_49490);
xor UO_1411 (O_1411,N_48759,N_49103);
and UO_1412 (O_1412,N_48313,N_48996);
and UO_1413 (O_1413,N_49765,N_47663);
and UO_1414 (O_1414,N_47979,N_47658);
and UO_1415 (O_1415,N_49232,N_48642);
nor UO_1416 (O_1416,N_49869,N_49632);
nor UO_1417 (O_1417,N_48992,N_49894);
and UO_1418 (O_1418,N_47903,N_47660);
nand UO_1419 (O_1419,N_49802,N_49497);
xnor UO_1420 (O_1420,N_47779,N_47649);
nand UO_1421 (O_1421,N_48244,N_49072);
xor UO_1422 (O_1422,N_48266,N_49940);
nand UO_1423 (O_1423,N_47766,N_48508);
and UO_1424 (O_1424,N_47758,N_48342);
or UO_1425 (O_1425,N_49091,N_49135);
nor UO_1426 (O_1426,N_48593,N_48472);
xnor UO_1427 (O_1427,N_47538,N_49813);
or UO_1428 (O_1428,N_49965,N_49387);
nand UO_1429 (O_1429,N_48858,N_47980);
or UO_1430 (O_1430,N_48501,N_49125);
nand UO_1431 (O_1431,N_48679,N_49084);
nand UO_1432 (O_1432,N_48937,N_48292);
nor UO_1433 (O_1433,N_47890,N_47851);
or UO_1434 (O_1434,N_49456,N_48119);
and UO_1435 (O_1435,N_48127,N_48493);
nand UO_1436 (O_1436,N_47613,N_48054);
or UO_1437 (O_1437,N_48746,N_48753);
nor UO_1438 (O_1438,N_49353,N_49872);
xnor UO_1439 (O_1439,N_47826,N_48458);
or UO_1440 (O_1440,N_47822,N_48310);
or UO_1441 (O_1441,N_49763,N_48392);
or UO_1442 (O_1442,N_47795,N_49865);
nand UO_1443 (O_1443,N_49260,N_48446);
nor UO_1444 (O_1444,N_47734,N_49476);
or UO_1445 (O_1445,N_49596,N_49882);
xor UO_1446 (O_1446,N_47579,N_47707);
nor UO_1447 (O_1447,N_48391,N_49069);
xnor UO_1448 (O_1448,N_48430,N_49783);
and UO_1449 (O_1449,N_48961,N_49734);
and UO_1450 (O_1450,N_49187,N_48753);
and UO_1451 (O_1451,N_48130,N_48102);
nor UO_1452 (O_1452,N_48442,N_47602);
or UO_1453 (O_1453,N_49690,N_47942);
and UO_1454 (O_1454,N_48228,N_49658);
xor UO_1455 (O_1455,N_49942,N_48682);
xnor UO_1456 (O_1456,N_48263,N_48001);
xnor UO_1457 (O_1457,N_49509,N_49492);
or UO_1458 (O_1458,N_49080,N_47767);
nor UO_1459 (O_1459,N_49092,N_48378);
xnor UO_1460 (O_1460,N_49561,N_49306);
nor UO_1461 (O_1461,N_49285,N_48434);
xnor UO_1462 (O_1462,N_48470,N_48237);
xnor UO_1463 (O_1463,N_48869,N_49709);
nand UO_1464 (O_1464,N_49244,N_49938);
nor UO_1465 (O_1465,N_48652,N_49860);
xor UO_1466 (O_1466,N_48350,N_48390);
xnor UO_1467 (O_1467,N_47735,N_48529);
or UO_1468 (O_1468,N_48516,N_48948);
nor UO_1469 (O_1469,N_48154,N_49053);
or UO_1470 (O_1470,N_49425,N_49939);
xor UO_1471 (O_1471,N_49352,N_49109);
xnor UO_1472 (O_1472,N_48148,N_49786);
or UO_1473 (O_1473,N_49328,N_49816);
or UO_1474 (O_1474,N_49025,N_49202);
xnor UO_1475 (O_1475,N_47608,N_49177);
or UO_1476 (O_1476,N_48627,N_47514);
and UO_1477 (O_1477,N_48805,N_49708);
nand UO_1478 (O_1478,N_48412,N_48584);
nor UO_1479 (O_1479,N_48451,N_48386);
xnor UO_1480 (O_1480,N_49708,N_49824);
nand UO_1481 (O_1481,N_48842,N_48105);
or UO_1482 (O_1482,N_48656,N_49806);
and UO_1483 (O_1483,N_49398,N_49664);
xor UO_1484 (O_1484,N_49175,N_49869);
and UO_1485 (O_1485,N_49571,N_49867);
nor UO_1486 (O_1486,N_48404,N_49965);
nor UO_1487 (O_1487,N_49365,N_49994);
xnor UO_1488 (O_1488,N_48216,N_49321);
nand UO_1489 (O_1489,N_48169,N_48180);
xor UO_1490 (O_1490,N_49717,N_47775);
and UO_1491 (O_1491,N_48641,N_48807);
or UO_1492 (O_1492,N_48690,N_48228);
or UO_1493 (O_1493,N_49322,N_48338);
nand UO_1494 (O_1494,N_49311,N_48953);
nand UO_1495 (O_1495,N_48060,N_49479);
and UO_1496 (O_1496,N_49622,N_49913);
or UO_1497 (O_1497,N_48187,N_49762);
xnor UO_1498 (O_1498,N_47547,N_47922);
nor UO_1499 (O_1499,N_47778,N_48202);
xnor UO_1500 (O_1500,N_48441,N_49987);
nor UO_1501 (O_1501,N_47769,N_47691);
xor UO_1502 (O_1502,N_47712,N_49320);
or UO_1503 (O_1503,N_49496,N_49727);
and UO_1504 (O_1504,N_49135,N_48780);
nor UO_1505 (O_1505,N_48085,N_49816);
or UO_1506 (O_1506,N_49936,N_47670);
xor UO_1507 (O_1507,N_48910,N_48003);
or UO_1508 (O_1508,N_47989,N_48666);
or UO_1509 (O_1509,N_48974,N_48038);
and UO_1510 (O_1510,N_48892,N_48413);
nor UO_1511 (O_1511,N_48833,N_49496);
nor UO_1512 (O_1512,N_49554,N_47500);
or UO_1513 (O_1513,N_49782,N_47538);
or UO_1514 (O_1514,N_49439,N_47886);
or UO_1515 (O_1515,N_49682,N_49646);
xor UO_1516 (O_1516,N_49266,N_48687);
nand UO_1517 (O_1517,N_48421,N_47826);
or UO_1518 (O_1518,N_49179,N_48399);
nor UO_1519 (O_1519,N_49528,N_49987);
nand UO_1520 (O_1520,N_48950,N_49073);
nand UO_1521 (O_1521,N_48239,N_49786);
nor UO_1522 (O_1522,N_49057,N_49960);
xnor UO_1523 (O_1523,N_48885,N_48990);
and UO_1524 (O_1524,N_48197,N_49082);
nand UO_1525 (O_1525,N_49271,N_47510);
or UO_1526 (O_1526,N_49036,N_48624);
nor UO_1527 (O_1527,N_49723,N_49677);
and UO_1528 (O_1528,N_49396,N_48232);
nor UO_1529 (O_1529,N_49273,N_49744);
xnor UO_1530 (O_1530,N_48810,N_49245);
xnor UO_1531 (O_1531,N_49945,N_48460);
or UO_1532 (O_1532,N_47992,N_48360);
nand UO_1533 (O_1533,N_49241,N_48439);
and UO_1534 (O_1534,N_48361,N_48934);
xnor UO_1535 (O_1535,N_49928,N_49438);
nor UO_1536 (O_1536,N_47620,N_49054);
or UO_1537 (O_1537,N_49833,N_48131);
xnor UO_1538 (O_1538,N_49776,N_49581);
xnor UO_1539 (O_1539,N_47618,N_48940);
or UO_1540 (O_1540,N_48019,N_49149);
xnor UO_1541 (O_1541,N_48318,N_49174);
xor UO_1542 (O_1542,N_48270,N_49130);
nand UO_1543 (O_1543,N_49020,N_49042);
xnor UO_1544 (O_1544,N_49006,N_47644);
nor UO_1545 (O_1545,N_48388,N_47621);
or UO_1546 (O_1546,N_49274,N_48043);
nor UO_1547 (O_1547,N_49737,N_49797);
nor UO_1548 (O_1548,N_49981,N_48198);
and UO_1549 (O_1549,N_49786,N_48316);
nor UO_1550 (O_1550,N_49247,N_49965);
and UO_1551 (O_1551,N_48973,N_49250);
or UO_1552 (O_1552,N_47648,N_48233);
and UO_1553 (O_1553,N_49493,N_49660);
xnor UO_1554 (O_1554,N_49510,N_47823);
and UO_1555 (O_1555,N_49936,N_49059);
and UO_1556 (O_1556,N_49003,N_49310);
or UO_1557 (O_1557,N_47513,N_47803);
nor UO_1558 (O_1558,N_48693,N_47929);
xor UO_1559 (O_1559,N_48132,N_48495);
nand UO_1560 (O_1560,N_49132,N_48655);
or UO_1561 (O_1561,N_49238,N_47942);
nor UO_1562 (O_1562,N_48167,N_47632);
xor UO_1563 (O_1563,N_49532,N_49950);
or UO_1564 (O_1564,N_49636,N_49533);
nor UO_1565 (O_1565,N_49338,N_49226);
xor UO_1566 (O_1566,N_49721,N_47528);
or UO_1567 (O_1567,N_49003,N_48587);
and UO_1568 (O_1568,N_47846,N_47983);
and UO_1569 (O_1569,N_48211,N_48403);
and UO_1570 (O_1570,N_48792,N_48549);
nor UO_1571 (O_1571,N_48376,N_49649);
nand UO_1572 (O_1572,N_47750,N_48378);
nand UO_1573 (O_1573,N_49201,N_48504);
xor UO_1574 (O_1574,N_48401,N_48419);
and UO_1575 (O_1575,N_49736,N_48351);
and UO_1576 (O_1576,N_49649,N_47845);
xor UO_1577 (O_1577,N_47512,N_48525);
xnor UO_1578 (O_1578,N_49869,N_47847);
or UO_1579 (O_1579,N_49478,N_49929);
or UO_1580 (O_1580,N_49515,N_48642);
and UO_1581 (O_1581,N_48610,N_49295);
xnor UO_1582 (O_1582,N_48515,N_48203);
or UO_1583 (O_1583,N_48161,N_49689);
and UO_1584 (O_1584,N_49802,N_49962);
or UO_1585 (O_1585,N_48721,N_47585);
nand UO_1586 (O_1586,N_48227,N_49358);
or UO_1587 (O_1587,N_49098,N_48456);
xor UO_1588 (O_1588,N_47653,N_48627);
and UO_1589 (O_1589,N_49661,N_49094);
or UO_1590 (O_1590,N_48741,N_49762);
and UO_1591 (O_1591,N_49124,N_48749);
xnor UO_1592 (O_1592,N_49235,N_48436);
xnor UO_1593 (O_1593,N_48687,N_48333);
nand UO_1594 (O_1594,N_48036,N_48295);
nand UO_1595 (O_1595,N_49122,N_49867);
nor UO_1596 (O_1596,N_48404,N_48761);
xnor UO_1597 (O_1597,N_47688,N_49597);
nor UO_1598 (O_1598,N_49071,N_49301);
xnor UO_1599 (O_1599,N_49085,N_47727);
nand UO_1600 (O_1600,N_47701,N_48501);
xnor UO_1601 (O_1601,N_48976,N_48592);
nand UO_1602 (O_1602,N_47535,N_48348);
or UO_1603 (O_1603,N_49907,N_47891);
nor UO_1604 (O_1604,N_49965,N_49917);
and UO_1605 (O_1605,N_47810,N_47892);
nor UO_1606 (O_1606,N_47706,N_48164);
xor UO_1607 (O_1607,N_48626,N_47711);
or UO_1608 (O_1608,N_48915,N_49775);
and UO_1609 (O_1609,N_48667,N_47577);
or UO_1610 (O_1610,N_49761,N_48191);
nor UO_1611 (O_1611,N_48636,N_49487);
nor UO_1612 (O_1612,N_49016,N_49111);
and UO_1613 (O_1613,N_47527,N_48821);
or UO_1614 (O_1614,N_48841,N_48654);
or UO_1615 (O_1615,N_49073,N_48271);
nand UO_1616 (O_1616,N_49304,N_48714);
or UO_1617 (O_1617,N_49861,N_47648);
nand UO_1618 (O_1618,N_48960,N_49859);
or UO_1619 (O_1619,N_48712,N_49322);
nand UO_1620 (O_1620,N_49003,N_48552);
nor UO_1621 (O_1621,N_48134,N_47889);
xor UO_1622 (O_1622,N_48615,N_49722);
or UO_1623 (O_1623,N_49781,N_48854);
and UO_1624 (O_1624,N_48635,N_48120);
or UO_1625 (O_1625,N_47968,N_48260);
nand UO_1626 (O_1626,N_47897,N_48377);
nor UO_1627 (O_1627,N_47946,N_48763);
nor UO_1628 (O_1628,N_47869,N_48383);
nand UO_1629 (O_1629,N_49819,N_49439);
nor UO_1630 (O_1630,N_49817,N_47763);
or UO_1631 (O_1631,N_49634,N_49851);
nor UO_1632 (O_1632,N_48779,N_48818);
or UO_1633 (O_1633,N_49459,N_48006);
or UO_1634 (O_1634,N_48025,N_48670);
xnor UO_1635 (O_1635,N_49652,N_47577);
xor UO_1636 (O_1636,N_49293,N_47845);
nand UO_1637 (O_1637,N_49752,N_47725);
or UO_1638 (O_1638,N_48818,N_48832);
and UO_1639 (O_1639,N_49341,N_49413);
nor UO_1640 (O_1640,N_48381,N_48277);
and UO_1641 (O_1641,N_49072,N_48412);
and UO_1642 (O_1642,N_47712,N_47860);
nand UO_1643 (O_1643,N_48678,N_49068);
or UO_1644 (O_1644,N_48546,N_47991);
xor UO_1645 (O_1645,N_49720,N_48464);
xnor UO_1646 (O_1646,N_49204,N_48166);
xor UO_1647 (O_1647,N_48341,N_48097);
nor UO_1648 (O_1648,N_49349,N_49132);
nor UO_1649 (O_1649,N_49824,N_49507);
nand UO_1650 (O_1650,N_49839,N_48508);
xnor UO_1651 (O_1651,N_47896,N_48140);
nand UO_1652 (O_1652,N_48105,N_49200);
nor UO_1653 (O_1653,N_49621,N_48043);
nand UO_1654 (O_1654,N_49461,N_49782);
xor UO_1655 (O_1655,N_49879,N_47937);
and UO_1656 (O_1656,N_49980,N_48201);
nor UO_1657 (O_1657,N_48536,N_49863);
and UO_1658 (O_1658,N_49826,N_48571);
nor UO_1659 (O_1659,N_48643,N_48599);
nand UO_1660 (O_1660,N_49259,N_48456);
or UO_1661 (O_1661,N_48328,N_49777);
nor UO_1662 (O_1662,N_47937,N_49551);
or UO_1663 (O_1663,N_48048,N_48034);
nand UO_1664 (O_1664,N_48879,N_47643);
nand UO_1665 (O_1665,N_49526,N_48147);
and UO_1666 (O_1666,N_49028,N_47884);
xnor UO_1667 (O_1667,N_49684,N_49328);
nand UO_1668 (O_1668,N_49869,N_49486);
and UO_1669 (O_1669,N_47570,N_48902);
nor UO_1670 (O_1670,N_49013,N_48181);
nor UO_1671 (O_1671,N_49149,N_49835);
or UO_1672 (O_1672,N_48306,N_49311);
xnor UO_1673 (O_1673,N_47603,N_47999);
and UO_1674 (O_1674,N_48314,N_48237);
nand UO_1675 (O_1675,N_47956,N_48514);
nand UO_1676 (O_1676,N_49865,N_48156);
and UO_1677 (O_1677,N_47726,N_49342);
nand UO_1678 (O_1678,N_49922,N_48081);
nand UO_1679 (O_1679,N_49593,N_48546);
nand UO_1680 (O_1680,N_48270,N_48817);
nand UO_1681 (O_1681,N_48539,N_48103);
and UO_1682 (O_1682,N_48026,N_49869);
and UO_1683 (O_1683,N_49864,N_48187);
nor UO_1684 (O_1684,N_47533,N_48928);
or UO_1685 (O_1685,N_48674,N_49733);
xor UO_1686 (O_1686,N_49562,N_49956);
xnor UO_1687 (O_1687,N_49202,N_49156);
nand UO_1688 (O_1688,N_48908,N_48403);
xnor UO_1689 (O_1689,N_48708,N_49336);
and UO_1690 (O_1690,N_47700,N_47705);
nand UO_1691 (O_1691,N_47969,N_47732);
nor UO_1692 (O_1692,N_49541,N_48458);
xor UO_1693 (O_1693,N_49438,N_47749);
or UO_1694 (O_1694,N_49309,N_47666);
and UO_1695 (O_1695,N_49903,N_49516);
xnor UO_1696 (O_1696,N_47741,N_47836);
and UO_1697 (O_1697,N_48034,N_48563);
or UO_1698 (O_1698,N_49362,N_49072);
nand UO_1699 (O_1699,N_47861,N_47949);
and UO_1700 (O_1700,N_48366,N_48747);
and UO_1701 (O_1701,N_48096,N_49957);
nand UO_1702 (O_1702,N_49804,N_49641);
and UO_1703 (O_1703,N_48053,N_49652);
nor UO_1704 (O_1704,N_48838,N_48311);
nor UO_1705 (O_1705,N_48686,N_48136);
nand UO_1706 (O_1706,N_47954,N_48300);
nor UO_1707 (O_1707,N_47598,N_49294);
or UO_1708 (O_1708,N_47763,N_48686);
or UO_1709 (O_1709,N_47985,N_48230);
xnor UO_1710 (O_1710,N_49315,N_47931);
xnor UO_1711 (O_1711,N_49541,N_49302);
nor UO_1712 (O_1712,N_49658,N_47539);
xor UO_1713 (O_1713,N_47672,N_49273);
nand UO_1714 (O_1714,N_48031,N_48420);
xnor UO_1715 (O_1715,N_48675,N_48863);
or UO_1716 (O_1716,N_49473,N_49425);
and UO_1717 (O_1717,N_49794,N_49292);
nor UO_1718 (O_1718,N_48002,N_47610);
and UO_1719 (O_1719,N_48385,N_47591);
nor UO_1720 (O_1720,N_49924,N_48585);
nand UO_1721 (O_1721,N_49261,N_48085);
or UO_1722 (O_1722,N_49086,N_47699);
and UO_1723 (O_1723,N_49991,N_49198);
or UO_1724 (O_1724,N_49353,N_48463);
xnor UO_1725 (O_1725,N_49675,N_47973);
and UO_1726 (O_1726,N_47763,N_49005);
or UO_1727 (O_1727,N_48129,N_48380);
xor UO_1728 (O_1728,N_48175,N_47712);
nor UO_1729 (O_1729,N_48952,N_48137);
nand UO_1730 (O_1730,N_48770,N_48555);
and UO_1731 (O_1731,N_48199,N_49055);
or UO_1732 (O_1732,N_48640,N_48916);
nor UO_1733 (O_1733,N_48539,N_48676);
and UO_1734 (O_1734,N_47578,N_48824);
xnor UO_1735 (O_1735,N_47854,N_48514);
and UO_1736 (O_1736,N_49896,N_48410);
and UO_1737 (O_1737,N_47841,N_49932);
or UO_1738 (O_1738,N_48509,N_47941);
nor UO_1739 (O_1739,N_49703,N_47879);
nor UO_1740 (O_1740,N_48600,N_48904);
nor UO_1741 (O_1741,N_48244,N_48376);
and UO_1742 (O_1742,N_48914,N_47822);
nor UO_1743 (O_1743,N_49013,N_49851);
nand UO_1744 (O_1744,N_47854,N_48599);
nand UO_1745 (O_1745,N_48920,N_48753);
or UO_1746 (O_1746,N_48391,N_47649);
nor UO_1747 (O_1747,N_48037,N_49669);
nand UO_1748 (O_1748,N_49795,N_47673);
nand UO_1749 (O_1749,N_49388,N_49434);
xor UO_1750 (O_1750,N_49247,N_49540);
nor UO_1751 (O_1751,N_47768,N_48317);
nand UO_1752 (O_1752,N_49089,N_49921);
and UO_1753 (O_1753,N_49619,N_47882);
nand UO_1754 (O_1754,N_49380,N_48843);
nor UO_1755 (O_1755,N_48909,N_49432);
nand UO_1756 (O_1756,N_48183,N_49887);
or UO_1757 (O_1757,N_48114,N_49263);
and UO_1758 (O_1758,N_48146,N_49955);
nor UO_1759 (O_1759,N_49220,N_49348);
xnor UO_1760 (O_1760,N_48425,N_47526);
xnor UO_1761 (O_1761,N_48686,N_49689);
and UO_1762 (O_1762,N_49266,N_47565);
and UO_1763 (O_1763,N_48808,N_47627);
nor UO_1764 (O_1764,N_47557,N_48745);
xnor UO_1765 (O_1765,N_48394,N_48523);
xor UO_1766 (O_1766,N_48737,N_49150);
and UO_1767 (O_1767,N_47679,N_48176);
and UO_1768 (O_1768,N_47725,N_49307);
nand UO_1769 (O_1769,N_49691,N_49260);
and UO_1770 (O_1770,N_47515,N_48475);
or UO_1771 (O_1771,N_49674,N_49776);
nand UO_1772 (O_1772,N_48596,N_47815);
or UO_1773 (O_1773,N_48372,N_48548);
nand UO_1774 (O_1774,N_48785,N_49698);
or UO_1775 (O_1775,N_49701,N_47508);
nand UO_1776 (O_1776,N_49664,N_47783);
xor UO_1777 (O_1777,N_48154,N_49645);
and UO_1778 (O_1778,N_49361,N_48245);
nand UO_1779 (O_1779,N_49023,N_47548);
and UO_1780 (O_1780,N_49602,N_49188);
nand UO_1781 (O_1781,N_47525,N_48753);
xnor UO_1782 (O_1782,N_48745,N_47723);
and UO_1783 (O_1783,N_48730,N_48676);
and UO_1784 (O_1784,N_48797,N_47747);
nand UO_1785 (O_1785,N_47937,N_49688);
xnor UO_1786 (O_1786,N_49245,N_47815);
xnor UO_1787 (O_1787,N_48329,N_48888);
and UO_1788 (O_1788,N_49212,N_48299);
nand UO_1789 (O_1789,N_49039,N_49796);
xor UO_1790 (O_1790,N_48261,N_48488);
nand UO_1791 (O_1791,N_47914,N_48155);
xnor UO_1792 (O_1792,N_48161,N_49579);
and UO_1793 (O_1793,N_49975,N_48665);
nor UO_1794 (O_1794,N_49692,N_48433);
nand UO_1795 (O_1795,N_49936,N_49944);
or UO_1796 (O_1796,N_49544,N_49804);
xnor UO_1797 (O_1797,N_47710,N_49446);
nand UO_1798 (O_1798,N_48244,N_49829);
and UO_1799 (O_1799,N_48093,N_49061);
xor UO_1800 (O_1800,N_49461,N_48298);
and UO_1801 (O_1801,N_48890,N_49967);
and UO_1802 (O_1802,N_48713,N_47552);
and UO_1803 (O_1803,N_47781,N_48352);
or UO_1804 (O_1804,N_49005,N_49301);
and UO_1805 (O_1805,N_49913,N_49583);
nand UO_1806 (O_1806,N_48170,N_49058);
nor UO_1807 (O_1807,N_48446,N_47719);
xor UO_1808 (O_1808,N_48030,N_49256);
and UO_1809 (O_1809,N_49703,N_49125);
nor UO_1810 (O_1810,N_48043,N_48598);
and UO_1811 (O_1811,N_49582,N_48550);
xor UO_1812 (O_1812,N_47508,N_49866);
nand UO_1813 (O_1813,N_49043,N_48564);
nand UO_1814 (O_1814,N_49945,N_49843);
nand UO_1815 (O_1815,N_48176,N_49844);
nand UO_1816 (O_1816,N_49240,N_48081);
and UO_1817 (O_1817,N_49192,N_48110);
or UO_1818 (O_1818,N_49601,N_49125);
nor UO_1819 (O_1819,N_48860,N_48041);
nor UO_1820 (O_1820,N_49091,N_48318);
or UO_1821 (O_1821,N_49945,N_48924);
nand UO_1822 (O_1822,N_49473,N_48148);
nor UO_1823 (O_1823,N_49923,N_49790);
and UO_1824 (O_1824,N_49859,N_48589);
or UO_1825 (O_1825,N_48178,N_49969);
xnor UO_1826 (O_1826,N_49674,N_48972);
and UO_1827 (O_1827,N_47994,N_49349);
xnor UO_1828 (O_1828,N_48194,N_48877);
xnor UO_1829 (O_1829,N_49188,N_48590);
nand UO_1830 (O_1830,N_49809,N_47964);
and UO_1831 (O_1831,N_49050,N_47606);
nand UO_1832 (O_1832,N_49999,N_47902);
nor UO_1833 (O_1833,N_48955,N_48673);
nand UO_1834 (O_1834,N_49411,N_48532);
nor UO_1835 (O_1835,N_49702,N_49134);
nor UO_1836 (O_1836,N_47816,N_48738);
nor UO_1837 (O_1837,N_49027,N_48515);
or UO_1838 (O_1838,N_48232,N_49553);
nor UO_1839 (O_1839,N_48773,N_49108);
xnor UO_1840 (O_1840,N_48595,N_49839);
nand UO_1841 (O_1841,N_47873,N_48622);
or UO_1842 (O_1842,N_47937,N_49592);
nor UO_1843 (O_1843,N_49049,N_48036);
nand UO_1844 (O_1844,N_49712,N_49277);
or UO_1845 (O_1845,N_47760,N_47820);
or UO_1846 (O_1846,N_49411,N_47702);
xor UO_1847 (O_1847,N_47807,N_47742);
xor UO_1848 (O_1848,N_49012,N_49756);
nand UO_1849 (O_1849,N_47868,N_49374);
and UO_1850 (O_1850,N_47938,N_49821);
or UO_1851 (O_1851,N_48720,N_48221);
or UO_1852 (O_1852,N_49401,N_48209);
or UO_1853 (O_1853,N_47687,N_49316);
nand UO_1854 (O_1854,N_48396,N_48977);
xor UO_1855 (O_1855,N_47667,N_48731);
or UO_1856 (O_1856,N_49419,N_49669);
and UO_1857 (O_1857,N_48900,N_47843);
and UO_1858 (O_1858,N_48055,N_47923);
nor UO_1859 (O_1859,N_48759,N_49511);
or UO_1860 (O_1860,N_49185,N_48751);
and UO_1861 (O_1861,N_48433,N_47896);
nor UO_1862 (O_1862,N_48644,N_48348);
nand UO_1863 (O_1863,N_48218,N_49021);
and UO_1864 (O_1864,N_49129,N_48965);
nand UO_1865 (O_1865,N_49893,N_49632);
xor UO_1866 (O_1866,N_49508,N_48315);
and UO_1867 (O_1867,N_48052,N_48984);
xor UO_1868 (O_1868,N_47736,N_47612);
or UO_1869 (O_1869,N_49173,N_48471);
or UO_1870 (O_1870,N_47741,N_47691);
and UO_1871 (O_1871,N_48644,N_47837);
or UO_1872 (O_1872,N_49568,N_47755);
or UO_1873 (O_1873,N_47667,N_48614);
xnor UO_1874 (O_1874,N_49589,N_49902);
xor UO_1875 (O_1875,N_49352,N_47993);
nor UO_1876 (O_1876,N_47801,N_48414);
xor UO_1877 (O_1877,N_49017,N_47605);
nand UO_1878 (O_1878,N_48131,N_47865);
nand UO_1879 (O_1879,N_48591,N_49920);
or UO_1880 (O_1880,N_47999,N_48754);
nand UO_1881 (O_1881,N_49129,N_48344);
or UO_1882 (O_1882,N_49596,N_49341);
nor UO_1883 (O_1883,N_48050,N_49139);
xnor UO_1884 (O_1884,N_48365,N_47555);
nand UO_1885 (O_1885,N_48289,N_48413);
nor UO_1886 (O_1886,N_49790,N_48112);
xnor UO_1887 (O_1887,N_49378,N_49600);
and UO_1888 (O_1888,N_48900,N_48537);
nor UO_1889 (O_1889,N_48197,N_49080);
or UO_1890 (O_1890,N_49756,N_47718);
or UO_1891 (O_1891,N_48726,N_47570);
nor UO_1892 (O_1892,N_47575,N_47727);
nand UO_1893 (O_1893,N_47584,N_48795);
xor UO_1894 (O_1894,N_48786,N_48293);
xnor UO_1895 (O_1895,N_48180,N_48995);
xnor UO_1896 (O_1896,N_48318,N_48360);
or UO_1897 (O_1897,N_48395,N_47839);
xnor UO_1898 (O_1898,N_49603,N_49929);
nand UO_1899 (O_1899,N_47849,N_48541);
xor UO_1900 (O_1900,N_49651,N_48442);
xor UO_1901 (O_1901,N_48002,N_49273);
and UO_1902 (O_1902,N_47985,N_49403);
and UO_1903 (O_1903,N_48215,N_49012);
or UO_1904 (O_1904,N_48151,N_48199);
and UO_1905 (O_1905,N_49179,N_49364);
nand UO_1906 (O_1906,N_48036,N_49737);
xor UO_1907 (O_1907,N_49296,N_47886);
and UO_1908 (O_1908,N_49672,N_47826);
and UO_1909 (O_1909,N_49601,N_48940);
xnor UO_1910 (O_1910,N_47760,N_48542);
and UO_1911 (O_1911,N_49677,N_48953);
nand UO_1912 (O_1912,N_48633,N_47656);
or UO_1913 (O_1913,N_48392,N_48786);
or UO_1914 (O_1914,N_48773,N_49319);
xor UO_1915 (O_1915,N_47935,N_49462);
nor UO_1916 (O_1916,N_48335,N_48109);
or UO_1917 (O_1917,N_49251,N_48826);
or UO_1918 (O_1918,N_47936,N_48341);
nand UO_1919 (O_1919,N_49471,N_48629);
nand UO_1920 (O_1920,N_49527,N_48842);
nand UO_1921 (O_1921,N_48424,N_47921);
nor UO_1922 (O_1922,N_49078,N_47931);
nor UO_1923 (O_1923,N_47655,N_47883);
or UO_1924 (O_1924,N_48003,N_48737);
nand UO_1925 (O_1925,N_47757,N_48834);
or UO_1926 (O_1926,N_49362,N_49594);
nor UO_1927 (O_1927,N_49956,N_49939);
nor UO_1928 (O_1928,N_47507,N_48337);
xnor UO_1929 (O_1929,N_49762,N_49197);
xnor UO_1930 (O_1930,N_49930,N_48814);
xnor UO_1931 (O_1931,N_48939,N_47920);
nand UO_1932 (O_1932,N_49669,N_49318);
nor UO_1933 (O_1933,N_47891,N_48377);
xor UO_1934 (O_1934,N_48948,N_48282);
or UO_1935 (O_1935,N_49919,N_49625);
nand UO_1936 (O_1936,N_48875,N_48128);
nand UO_1937 (O_1937,N_48300,N_48166);
and UO_1938 (O_1938,N_47524,N_48788);
and UO_1939 (O_1939,N_49121,N_48442);
nand UO_1940 (O_1940,N_47966,N_48458);
or UO_1941 (O_1941,N_48307,N_48313);
xnor UO_1942 (O_1942,N_48270,N_48242);
and UO_1943 (O_1943,N_47712,N_49687);
or UO_1944 (O_1944,N_48770,N_49787);
and UO_1945 (O_1945,N_47901,N_49481);
nand UO_1946 (O_1946,N_49755,N_47658);
and UO_1947 (O_1947,N_49674,N_48976);
nor UO_1948 (O_1948,N_48716,N_48194);
nand UO_1949 (O_1949,N_48660,N_49294);
or UO_1950 (O_1950,N_48415,N_49106);
xnor UO_1951 (O_1951,N_48399,N_48710);
and UO_1952 (O_1952,N_48364,N_47691);
or UO_1953 (O_1953,N_47736,N_47504);
nor UO_1954 (O_1954,N_49869,N_48543);
nand UO_1955 (O_1955,N_48555,N_47692);
and UO_1956 (O_1956,N_49784,N_47708);
nor UO_1957 (O_1957,N_48778,N_48130);
nor UO_1958 (O_1958,N_48224,N_47773);
or UO_1959 (O_1959,N_49826,N_48540);
or UO_1960 (O_1960,N_48498,N_47525);
and UO_1961 (O_1961,N_47577,N_48693);
xor UO_1962 (O_1962,N_48057,N_48436);
and UO_1963 (O_1963,N_47513,N_47949);
or UO_1964 (O_1964,N_48832,N_48130);
and UO_1965 (O_1965,N_48709,N_48851);
and UO_1966 (O_1966,N_48852,N_48424);
xnor UO_1967 (O_1967,N_49636,N_47718);
and UO_1968 (O_1968,N_48320,N_48403);
and UO_1969 (O_1969,N_48564,N_48286);
nor UO_1970 (O_1970,N_49926,N_49324);
and UO_1971 (O_1971,N_49283,N_49457);
or UO_1972 (O_1972,N_49211,N_49520);
xnor UO_1973 (O_1973,N_48535,N_48900);
xor UO_1974 (O_1974,N_49501,N_47578);
xor UO_1975 (O_1975,N_49468,N_47811);
or UO_1976 (O_1976,N_49988,N_49230);
nor UO_1977 (O_1977,N_49535,N_48835);
nor UO_1978 (O_1978,N_47640,N_49162);
nand UO_1979 (O_1979,N_48937,N_48458);
and UO_1980 (O_1980,N_49933,N_48802);
nand UO_1981 (O_1981,N_49769,N_47776);
or UO_1982 (O_1982,N_49439,N_49080);
xnor UO_1983 (O_1983,N_49964,N_47719);
nor UO_1984 (O_1984,N_49330,N_49245);
nor UO_1985 (O_1985,N_49115,N_48202);
xor UO_1986 (O_1986,N_49230,N_48479);
xor UO_1987 (O_1987,N_49866,N_49212);
nand UO_1988 (O_1988,N_49374,N_49350);
and UO_1989 (O_1989,N_49529,N_47643);
nand UO_1990 (O_1990,N_49467,N_47768);
and UO_1991 (O_1991,N_49888,N_49393);
nand UO_1992 (O_1992,N_47668,N_48719);
nand UO_1993 (O_1993,N_48257,N_48093);
or UO_1994 (O_1994,N_47876,N_49970);
or UO_1995 (O_1995,N_48946,N_49891);
nor UO_1996 (O_1996,N_48909,N_49747);
xnor UO_1997 (O_1997,N_49222,N_49002);
or UO_1998 (O_1998,N_47774,N_48954);
and UO_1999 (O_1999,N_49101,N_48563);
nand UO_2000 (O_2000,N_48423,N_48889);
xnor UO_2001 (O_2001,N_49450,N_49554);
xor UO_2002 (O_2002,N_49169,N_48509);
or UO_2003 (O_2003,N_48176,N_48836);
or UO_2004 (O_2004,N_49812,N_48104);
nand UO_2005 (O_2005,N_49482,N_48061);
nor UO_2006 (O_2006,N_48677,N_49729);
nand UO_2007 (O_2007,N_48925,N_49800);
xnor UO_2008 (O_2008,N_47790,N_49608);
nand UO_2009 (O_2009,N_47836,N_47794);
and UO_2010 (O_2010,N_48939,N_49372);
or UO_2011 (O_2011,N_49144,N_48311);
and UO_2012 (O_2012,N_49377,N_48740);
or UO_2013 (O_2013,N_48419,N_48535);
xnor UO_2014 (O_2014,N_48332,N_49813);
and UO_2015 (O_2015,N_47751,N_48817);
nor UO_2016 (O_2016,N_49632,N_48887);
and UO_2017 (O_2017,N_49355,N_48539);
nand UO_2018 (O_2018,N_48024,N_47735);
or UO_2019 (O_2019,N_48496,N_47624);
nor UO_2020 (O_2020,N_49479,N_48946);
xnor UO_2021 (O_2021,N_49247,N_48625);
and UO_2022 (O_2022,N_49428,N_49896);
nand UO_2023 (O_2023,N_49909,N_48515);
and UO_2024 (O_2024,N_47507,N_48493);
xor UO_2025 (O_2025,N_49326,N_49342);
or UO_2026 (O_2026,N_49691,N_49524);
or UO_2027 (O_2027,N_48160,N_48182);
nor UO_2028 (O_2028,N_47635,N_49542);
or UO_2029 (O_2029,N_47791,N_47935);
or UO_2030 (O_2030,N_48150,N_49087);
nor UO_2031 (O_2031,N_48783,N_48083);
nand UO_2032 (O_2032,N_47956,N_48743);
and UO_2033 (O_2033,N_48059,N_49155);
xor UO_2034 (O_2034,N_48972,N_48777);
xnor UO_2035 (O_2035,N_49192,N_47684);
nor UO_2036 (O_2036,N_49179,N_47990);
nand UO_2037 (O_2037,N_49780,N_48738);
or UO_2038 (O_2038,N_48514,N_48876);
nor UO_2039 (O_2039,N_48964,N_48342);
and UO_2040 (O_2040,N_49255,N_48895);
or UO_2041 (O_2041,N_48168,N_47552);
and UO_2042 (O_2042,N_48355,N_49256);
nor UO_2043 (O_2043,N_48727,N_49569);
or UO_2044 (O_2044,N_49863,N_49896);
or UO_2045 (O_2045,N_48021,N_47512);
nor UO_2046 (O_2046,N_49025,N_48708);
nand UO_2047 (O_2047,N_49149,N_48283);
nand UO_2048 (O_2048,N_48837,N_47999);
nand UO_2049 (O_2049,N_48262,N_48139);
nand UO_2050 (O_2050,N_48714,N_49392);
xor UO_2051 (O_2051,N_48060,N_47917);
nand UO_2052 (O_2052,N_48409,N_49131);
nand UO_2053 (O_2053,N_49063,N_49293);
xnor UO_2054 (O_2054,N_49680,N_49302);
nor UO_2055 (O_2055,N_48400,N_47735);
nand UO_2056 (O_2056,N_48677,N_48534);
and UO_2057 (O_2057,N_48212,N_47524);
nor UO_2058 (O_2058,N_49116,N_49573);
nand UO_2059 (O_2059,N_49788,N_48266);
nor UO_2060 (O_2060,N_48549,N_48820);
or UO_2061 (O_2061,N_48798,N_49339);
nor UO_2062 (O_2062,N_49832,N_49662);
nand UO_2063 (O_2063,N_48188,N_49439);
or UO_2064 (O_2064,N_48934,N_48970);
xnor UO_2065 (O_2065,N_48850,N_48180);
and UO_2066 (O_2066,N_49642,N_48865);
nand UO_2067 (O_2067,N_48183,N_48628);
xnor UO_2068 (O_2068,N_49446,N_48882);
xor UO_2069 (O_2069,N_47770,N_48930);
and UO_2070 (O_2070,N_49230,N_49754);
and UO_2071 (O_2071,N_48017,N_47894);
or UO_2072 (O_2072,N_48037,N_47840);
nor UO_2073 (O_2073,N_48331,N_49188);
or UO_2074 (O_2074,N_49150,N_47822);
and UO_2075 (O_2075,N_48500,N_49756);
or UO_2076 (O_2076,N_49078,N_49852);
nor UO_2077 (O_2077,N_48456,N_49913);
nor UO_2078 (O_2078,N_49361,N_47822);
nand UO_2079 (O_2079,N_48702,N_48904);
nand UO_2080 (O_2080,N_48795,N_48400);
nor UO_2081 (O_2081,N_47533,N_49434);
xor UO_2082 (O_2082,N_47986,N_48390);
xor UO_2083 (O_2083,N_47877,N_48121);
xnor UO_2084 (O_2084,N_48289,N_47625);
and UO_2085 (O_2085,N_47644,N_48739);
nor UO_2086 (O_2086,N_47780,N_47637);
or UO_2087 (O_2087,N_48856,N_49137);
xnor UO_2088 (O_2088,N_49051,N_47940);
xnor UO_2089 (O_2089,N_47775,N_49477);
and UO_2090 (O_2090,N_49734,N_49348);
and UO_2091 (O_2091,N_48538,N_49921);
nor UO_2092 (O_2092,N_47966,N_47828);
nand UO_2093 (O_2093,N_47617,N_47862);
xnor UO_2094 (O_2094,N_48830,N_49077);
nor UO_2095 (O_2095,N_48013,N_48915);
or UO_2096 (O_2096,N_48344,N_48801);
and UO_2097 (O_2097,N_48789,N_49280);
nand UO_2098 (O_2098,N_49850,N_48691);
or UO_2099 (O_2099,N_49572,N_48949);
nand UO_2100 (O_2100,N_49720,N_48147);
nor UO_2101 (O_2101,N_49797,N_48715);
xor UO_2102 (O_2102,N_49685,N_48798);
or UO_2103 (O_2103,N_48457,N_48420);
nand UO_2104 (O_2104,N_47750,N_49689);
and UO_2105 (O_2105,N_48531,N_48878);
or UO_2106 (O_2106,N_48979,N_48982);
nand UO_2107 (O_2107,N_47840,N_48176);
nor UO_2108 (O_2108,N_48278,N_49479);
nand UO_2109 (O_2109,N_48436,N_48829);
or UO_2110 (O_2110,N_48670,N_49939);
nor UO_2111 (O_2111,N_49264,N_47672);
nor UO_2112 (O_2112,N_47954,N_47771);
and UO_2113 (O_2113,N_48241,N_49122);
or UO_2114 (O_2114,N_48224,N_47796);
nor UO_2115 (O_2115,N_49879,N_48812);
nor UO_2116 (O_2116,N_48318,N_48760);
or UO_2117 (O_2117,N_47837,N_48226);
nor UO_2118 (O_2118,N_48386,N_49960);
xnor UO_2119 (O_2119,N_49440,N_48626);
xnor UO_2120 (O_2120,N_48392,N_48280);
nor UO_2121 (O_2121,N_48268,N_49543);
or UO_2122 (O_2122,N_47974,N_48529);
and UO_2123 (O_2123,N_48555,N_49485);
xor UO_2124 (O_2124,N_49531,N_48566);
and UO_2125 (O_2125,N_48476,N_48579);
nor UO_2126 (O_2126,N_49682,N_49757);
and UO_2127 (O_2127,N_49339,N_49103);
nor UO_2128 (O_2128,N_49277,N_47724);
nand UO_2129 (O_2129,N_49915,N_47836);
or UO_2130 (O_2130,N_49620,N_48467);
nand UO_2131 (O_2131,N_47748,N_49488);
or UO_2132 (O_2132,N_49661,N_48947);
and UO_2133 (O_2133,N_48689,N_48859);
nand UO_2134 (O_2134,N_49337,N_48331);
and UO_2135 (O_2135,N_49907,N_47500);
nor UO_2136 (O_2136,N_47550,N_48476);
xor UO_2137 (O_2137,N_49587,N_48334);
and UO_2138 (O_2138,N_49828,N_49291);
and UO_2139 (O_2139,N_48141,N_47684);
nand UO_2140 (O_2140,N_48293,N_47886);
nor UO_2141 (O_2141,N_49700,N_47917);
or UO_2142 (O_2142,N_48220,N_48792);
nand UO_2143 (O_2143,N_49948,N_48267);
or UO_2144 (O_2144,N_49409,N_48391);
nor UO_2145 (O_2145,N_49587,N_48417);
and UO_2146 (O_2146,N_47709,N_47831);
nand UO_2147 (O_2147,N_47951,N_48668);
and UO_2148 (O_2148,N_49205,N_47593);
xor UO_2149 (O_2149,N_49014,N_47508);
xor UO_2150 (O_2150,N_48120,N_47830);
xnor UO_2151 (O_2151,N_49089,N_47992);
xor UO_2152 (O_2152,N_48578,N_47520);
and UO_2153 (O_2153,N_49603,N_49605);
nor UO_2154 (O_2154,N_47864,N_48217);
nor UO_2155 (O_2155,N_49465,N_48013);
nor UO_2156 (O_2156,N_48812,N_49066);
and UO_2157 (O_2157,N_48885,N_48766);
nand UO_2158 (O_2158,N_49085,N_48233);
nor UO_2159 (O_2159,N_47911,N_48577);
or UO_2160 (O_2160,N_49501,N_49749);
or UO_2161 (O_2161,N_48106,N_49736);
or UO_2162 (O_2162,N_47817,N_48483);
and UO_2163 (O_2163,N_48602,N_48989);
nor UO_2164 (O_2164,N_47586,N_48048);
or UO_2165 (O_2165,N_49280,N_49502);
nand UO_2166 (O_2166,N_47835,N_49409);
nor UO_2167 (O_2167,N_48001,N_48564);
nand UO_2168 (O_2168,N_47864,N_49579);
nor UO_2169 (O_2169,N_48259,N_48316);
xnor UO_2170 (O_2170,N_49178,N_49972);
or UO_2171 (O_2171,N_49382,N_48000);
or UO_2172 (O_2172,N_48582,N_48709);
nand UO_2173 (O_2173,N_49664,N_48516);
and UO_2174 (O_2174,N_49992,N_48886);
nand UO_2175 (O_2175,N_47827,N_49826);
xor UO_2176 (O_2176,N_49935,N_48031);
or UO_2177 (O_2177,N_49498,N_48942);
and UO_2178 (O_2178,N_49894,N_48444);
xor UO_2179 (O_2179,N_48897,N_49997);
nor UO_2180 (O_2180,N_49669,N_48335);
xnor UO_2181 (O_2181,N_49025,N_48301);
and UO_2182 (O_2182,N_48445,N_48328);
or UO_2183 (O_2183,N_49652,N_48733);
xor UO_2184 (O_2184,N_48364,N_48296);
and UO_2185 (O_2185,N_48629,N_48338);
nor UO_2186 (O_2186,N_48757,N_48371);
xnor UO_2187 (O_2187,N_48919,N_49731);
nand UO_2188 (O_2188,N_49014,N_49993);
nand UO_2189 (O_2189,N_49378,N_49563);
and UO_2190 (O_2190,N_48127,N_49958);
or UO_2191 (O_2191,N_47650,N_48069);
nand UO_2192 (O_2192,N_47637,N_49636);
nor UO_2193 (O_2193,N_49661,N_49719);
or UO_2194 (O_2194,N_49541,N_49455);
nor UO_2195 (O_2195,N_49971,N_48421);
nor UO_2196 (O_2196,N_47612,N_49120);
xnor UO_2197 (O_2197,N_48709,N_47826);
or UO_2198 (O_2198,N_49348,N_49591);
xnor UO_2199 (O_2199,N_49005,N_49504);
nor UO_2200 (O_2200,N_49344,N_49588);
xnor UO_2201 (O_2201,N_47978,N_47724);
and UO_2202 (O_2202,N_49942,N_49325);
or UO_2203 (O_2203,N_49268,N_48437);
or UO_2204 (O_2204,N_48787,N_49891);
nor UO_2205 (O_2205,N_48804,N_48256);
or UO_2206 (O_2206,N_47532,N_49544);
xor UO_2207 (O_2207,N_47730,N_49042);
nor UO_2208 (O_2208,N_48211,N_49588);
and UO_2209 (O_2209,N_47860,N_47783);
nand UO_2210 (O_2210,N_48915,N_47886);
nor UO_2211 (O_2211,N_47989,N_47790);
nor UO_2212 (O_2212,N_47615,N_47842);
and UO_2213 (O_2213,N_49705,N_49577);
nand UO_2214 (O_2214,N_49313,N_49364);
nand UO_2215 (O_2215,N_49624,N_47632);
nand UO_2216 (O_2216,N_47886,N_48402);
nand UO_2217 (O_2217,N_49684,N_49727);
xor UO_2218 (O_2218,N_49242,N_49060);
nand UO_2219 (O_2219,N_48149,N_49527);
or UO_2220 (O_2220,N_49371,N_49457);
or UO_2221 (O_2221,N_49034,N_48235);
and UO_2222 (O_2222,N_49593,N_47720);
nor UO_2223 (O_2223,N_49239,N_49306);
nor UO_2224 (O_2224,N_49678,N_49367);
and UO_2225 (O_2225,N_48942,N_48741);
and UO_2226 (O_2226,N_48393,N_47629);
xnor UO_2227 (O_2227,N_48226,N_49677);
or UO_2228 (O_2228,N_49751,N_49293);
or UO_2229 (O_2229,N_48990,N_47977);
xor UO_2230 (O_2230,N_49620,N_47966);
or UO_2231 (O_2231,N_47825,N_48016);
or UO_2232 (O_2232,N_48408,N_48388);
and UO_2233 (O_2233,N_48426,N_47779);
and UO_2234 (O_2234,N_49209,N_49158);
xor UO_2235 (O_2235,N_49696,N_47694);
nand UO_2236 (O_2236,N_49366,N_48115);
or UO_2237 (O_2237,N_47568,N_49342);
and UO_2238 (O_2238,N_49104,N_47993);
nand UO_2239 (O_2239,N_48130,N_47687);
nand UO_2240 (O_2240,N_49412,N_49850);
xnor UO_2241 (O_2241,N_49659,N_48428);
or UO_2242 (O_2242,N_49486,N_48851);
nand UO_2243 (O_2243,N_48918,N_48475);
or UO_2244 (O_2244,N_47629,N_48332);
nand UO_2245 (O_2245,N_48484,N_48424);
nor UO_2246 (O_2246,N_47576,N_47960);
nor UO_2247 (O_2247,N_48302,N_49816);
nor UO_2248 (O_2248,N_47881,N_48712);
and UO_2249 (O_2249,N_48385,N_49371);
nor UO_2250 (O_2250,N_48914,N_47612);
xor UO_2251 (O_2251,N_49490,N_48134);
and UO_2252 (O_2252,N_47769,N_49395);
nor UO_2253 (O_2253,N_49384,N_47960);
or UO_2254 (O_2254,N_49006,N_48962);
or UO_2255 (O_2255,N_47656,N_49628);
or UO_2256 (O_2256,N_48555,N_49551);
and UO_2257 (O_2257,N_48138,N_49030);
nor UO_2258 (O_2258,N_48272,N_48244);
or UO_2259 (O_2259,N_49055,N_47901);
nand UO_2260 (O_2260,N_48574,N_48054);
nand UO_2261 (O_2261,N_48750,N_49962);
and UO_2262 (O_2262,N_48236,N_47553);
and UO_2263 (O_2263,N_48017,N_48054);
nor UO_2264 (O_2264,N_48814,N_48282);
or UO_2265 (O_2265,N_48541,N_49858);
and UO_2266 (O_2266,N_49313,N_49274);
nor UO_2267 (O_2267,N_48733,N_49747);
or UO_2268 (O_2268,N_48412,N_49489);
and UO_2269 (O_2269,N_48506,N_49818);
and UO_2270 (O_2270,N_47665,N_47716);
xor UO_2271 (O_2271,N_49893,N_48857);
or UO_2272 (O_2272,N_48656,N_49000);
nor UO_2273 (O_2273,N_47846,N_48436);
nand UO_2274 (O_2274,N_48965,N_48137);
nand UO_2275 (O_2275,N_49863,N_48441);
nor UO_2276 (O_2276,N_49848,N_48897);
nor UO_2277 (O_2277,N_48216,N_49902);
xnor UO_2278 (O_2278,N_48896,N_47553);
nor UO_2279 (O_2279,N_47899,N_48347);
nor UO_2280 (O_2280,N_49981,N_48653);
nand UO_2281 (O_2281,N_48365,N_47547);
or UO_2282 (O_2282,N_49215,N_49574);
nor UO_2283 (O_2283,N_49639,N_48936);
and UO_2284 (O_2284,N_48451,N_48958);
nand UO_2285 (O_2285,N_49184,N_49544);
and UO_2286 (O_2286,N_49292,N_47916);
nand UO_2287 (O_2287,N_48509,N_49595);
nor UO_2288 (O_2288,N_47629,N_47909);
xnor UO_2289 (O_2289,N_48145,N_49378);
or UO_2290 (O_2290,N_48897,N_49467);
nor UO_2291 (O_2291,N_49538,N_48566);
or UO_2292 (O_2292,N_49829,N_48765);
nor UO_2293 (O_2293,N_48106,N_48324);
or UO_2294 (O_2294,N_49652,N_49592);
nor UO_2295 (O_2295,N_48032,N_48306);
xor UO_2296 (O_2296,N_49420,N_47806);
xor UO_2297 (O_2297,N_47931,N_47871);
nand UO_2298 (O_2298,N_49921,N_48587);
nand UO_2299 (O_2299,N_49379,N_49760);
nand UO_2300 (O_2300,N_49181,N_49919);
xor UO_2301 (O_2301,N_49194,N_48698);
xnor UO_2302 (O_2302,N_48976,N_49600);
and UO_2303 (O_2303,N_48845,N_49054);
or UO_2304 (O_2304,N_49264,N_49122);
nand UO_2305 (O_2305,N_49352,N_48867);
nor UO_2306 (O_2306,N_49308,N_49678);
xnor UO_2307 (O_2307,N_48295,N_49438);
nand UO_2308 (O_2308,N_48957,N_49530);
nor UO_2309 (O_2309,N_49956,N_49456);
and UO_2310 (O_2310,N_49385,N_49827);
and UO_2311 (O_2311,N_48094,N_48701);
nor UO_2312 (O_2312,N_47522,N_47743);
nand UO_2313 (O_2313,N_47707,N_49107);
or UO_2314 (O_2314,N_48511,N_48507);
nor UO_2315 (O_2315,N_48662,N_49928);
xnor UO_2316 (O_2316,N_48947,N_47548);
or UO_2317 (O_2317,N_47713,N_47548);
nand UO_2318 (O_2318,N_48777,N_49568);
nor UO_2319 (O_2319,N_48613,N_49475);
xnor UO_2320 (O_2320,N_48912,N_47526);
nand UO_2321 (O_2321,N_48128,N_48052);
nand UO_2322 (O_2322,N_49505,N_49500);
nand UO_2323 (O_2323,N_47846,N_48798);
or UO_2324 (O_2324,N_48511,N_49262);
and UO_2325 (O_2325,N_49003,N_49716);
nor UO_2326 (O_2326,N_49476,N_49734);
nor UO_2327 (O_2327,N_49843,N_47774);
xor UO_2328 (O_2328,N_48947,N_49286);
or UO_2329 (O_2329,N_48667,N_48942);
or UO_2330 (O_2330,N_49435,N_49342);
nor UO_2331 (O_2331,N_48653,N_49932);
and UO_2332 (O_2332,N_48598,N_48415);
xnor UO_2333 (O_2333,N_48900,N_49800);
nand UO_2334 (O_2334,N_48609,N_48153);
nor UO_2335 (O_2335,N_49538,N_49806);
xor UO_2336 (O_2336,N_49472,N_49325);
or UO_2337 (O_2337,N_48880,N_47580);
or UO_2338 (O_2338,N_49411,N_48681);
xor UO_2339 (O_2339,N_49960,N_48258);
and UO_2340 (O_2340,N_49149,N_47616);
or UO_2341 (O_2341,N_48480,N_49193);
and UO_2342 (O_2342,N_49862,N_48023);
nor UO_2343 (O_2343,N_48850,N_49383);
and UO_2344 (O_2344,N_49685,N_48740);
xor UO_2345 (O_2345,N_49674,N_48792);
or UO_2346 (O_2346,N_49951,N_47510);
nand UO_2347 (O_2347,N_48182,N_48762);
and UO_2348 (O_2348,N_48540,N_49029);
or UO_2349 (O_2349,N_48448,N_48936);
or UO_2350 (O_2350,N_48065,N_47744);
nor UO_2351 (O_2351,N_49193,N_47863);
or UO_2352 (O_2352,N_47751,N_49135);
nor UO_2353 (O_2353,N_47658,N_48554);
nor UO_2354 (O_2354,N_49660,N_47921);
xnor UO_2355 (O_2355,N_49495,N_48580);
nand UO_2356 (O_2356,N_48430,N_47648);
and UO_2357 (O_2357,N_49284,N_48293);
and UO_2358 (O_2358,N_49828,N_48214);
xnor UO_2359 (O_2359,N_47910,N_48867);
nand UO_2360 (O_2360,N_49873,N_49976);
nand UO_2361 (O_2361,N_48451,N_48069);
and UO_2362 (O_2362,N_49464,N_48698);
or UO_2363 (O_2363,N_48879,N_49416);
xor UO_2364 (O_2364,N_48568,N_47932);
xnor UO_2365 (O_2365,N_49183,N_49627);
nor UO_2366 (O_2366,N_49240,N_49271);
xor UO_2367 (O_2367,N_48145,N_49937);
nand UO_2368 (O_2368,N_48110,N_48204);
or UO_2369 (O_2369,N_47796,N_48172);
xor UO_2370 (O_2370,N_49934,N_48702);
and UO_2371 (O_2371,N_48941,N_47960);
or UO_2372 (O_2372,N_49890,N_47914);
or UO_2373 (O_2373,N_49064,N_49397);
nor UO_2374 (O_2374,N_48006,N_48675);
xnor UO_2375 (O_2375,N_48191,N_48821);
nand UO_2376 (O_2376,N_49455,N_48277);
nand UO_2377 (O_2377,N_49861,N_49901);
or UO_2378 (O_2378,N_47770,N_48620);
and UO_2379 (O_2379,N_48653,N_49526);
nand UO_2380 (O_2380,N_49035,N_47517);
nand UO_2381 (O_2381,N_47568,N_47903);
or UO_2382 (O_2382,N_48573,N_49738);
xor UO_2383 (O_2383,N_48572,N_47656);
or UO_2384 (O_2384,N_48776,N_48066);
and UO_2385 (O_2385,N_49688,N_48017);
or UO_2386 (O_2386,N_48373,N_48011);
nand UO_2387 (O_2387,N_47584,N_49575);
xor UO_2388 (O_2388,N_47841,N_49445);
and UO_2389 (O_2389,N_48764,N_49125);
nor UO_2390 (O_2390,N_48372,N_47576);
nand UO_2391 (O_2391,N_48611,N_47790);
nor UO_2392 (O_2392,N_49234,N_47538);
nand UO_2393 (O_2393,N_49296,N_48309);
nor UO_2394 (O_2394,N_48512,N_49237);
xor UO_2395 (O_2395,N_47848,N_48430);
nand UO_2396 (O_2396,N_49240,N_48170);
xnor UO_2397 (O_2397,N_48382,N_49851);
xor UO_2398 (O_2398,N_47596,N_47571);
xor UO_2399 (O_2399,N_48469,N_47703);
and UO_2400 (O_2400,N_48399,N_47761);
nand UO_2401 (O_2401,N_49200,N_48957);
and UO_2402 (O_2402,N_47774,N_48274);
or UO_2403 (O_2403,N_47527,N_49220);
or UO_2404 (O_2404,N_48074,N_48987);
and UO_2405 (O_2405,N_48681,N_48324);
or UO_2406 (O_2406,N_49990,N_48416);
nand UO_2407 (O_2407,N_47758,N_47680);
nor UO_2408 (O_2408,N_48623,N_47908);
nand UO_2409 (O_2409,N_48499,N_47564);
nand UO_2410 (O_2410,N_49221,N_49780);
or UO_2411 (O_2411,N_47606,N_47551);
or UO_2412 (O_2412,N_49931,N_48538);
nand UO_2413 (O_2413,N_49795,N_48140);
nor UO_2414 (O_2414,N_48067,N_49543);
nor UO_2415 (O_2415,N_49192,N_47828);
nor UO_2416 (O_2416,N_49785,N_49945);
nor UO_2417 (O_2417,N_49849,N_48687);
nand UO_2418 (O_2418,N_48463,N_47544);
xnor UO_2419 (O_2419,N_47674,N_49488);
and UO_2420 (O_2420,N_48101,N_49645);
and UO_2421 (O_2421,N_49331,N_47794);
nand UO_2422 (O_2422,N_48384,N_49592);
nor UO_2423 (O_2423,N_49403,N_47835);
nor UO_2424 (O_2424,N_49886,N_49859);
xor UO_2425 (O_2425,N_49157,N_49089);
or UO_2426 (O_2426,N_47821,N_48031);
and UO_2427 (O_2427,N_48986,N_49409);
nor UO_2428 (O_2428,N_47867,N_48731);
and UO_2429 (O_2429,N_48399,N_48063);
nor UO_2430 (O_2430,N_48283,N_47721);
or UO_2431 (O_2431,N_49758,N_48658);
nand UO_2432 (O_2432,N_49968,N_48886);
or UO_2433 (O_2433,N_49637,N_48212);
xor UO_2434 (O_2434,N_47794,N_48232);
and UO_2435 (O_2435,N_48142,N_48915);
nor UO_2436 (O_2436,N_49218,N_49970);
nor UO_2437 (O_2437,N_47592,N_49189);
or UO_2438 (O_2438,N_49797,N_48148);
or UO_2439 (O_2439,N_47953,N_47515);
and UO_2440 (O_2440,N_48509,N_49292);
or UO_2441 (O_2441,N_48998,N_48749);
or UO_2442 (O_2442,N_49434,N_49821);
xnor UO_2443 (O_2443,N_49568,N_49982);
xnor UO_2444 (O_2444,N_49989,N_49072);
xnor UO_2445 (O_2445,N_49786,N_47668);
nor UO_2446 (O_2446,N_48999,N_47899);
and UO_2447 (O_2447,N_48291,N_47586);
or UO_2448 (O_2448,N_47749,N_49835);
or UO_2449 (O_2449,N_49284,N_49376);
and UO_2450 (O_2450,N_49878,N_49221);
nand UO_2451 (O_2451,N_49657,N_49094);
and UO_2452 (O_2452,N_48993,N_49450);
and UO_2453 (O_2453,N_49939,N_49153);
xnor UO_2454 (O_2454,N_49438,N_49878);
nand UO_2455 (O_2455,N_49644,N_48300);
or UO_2456 (O_2456,N_49350,N_49480);
nand UO_2457 (O_2457,N_49571,N_49458);
xnor UO_2458 (O_2458,N_47611,N_48941);
nand UO_2459 (O_2459,N_48613,N_49483);
or UO_2460 (O_2460,N_49969,N_48097);
nor UO_2461 (O_2461,N_48451,N_49162);
nand UO_2462 (O_2462,N_47703,N_47948);
or UO_2463 (O_2463,N_49448,N_49336);
nand UO_2464 (O_2464,N_48603,N_49444);
or UO_2465 (O_2465,N_47571,N_48345);
nand UO_2466 (O_2466,N_48654,N_48829);
xor UO_2467 (O_2467,N_48359,N_49112);
nor UO_2468 (O_2468,N_48260,N_49579);
xnor UO_2469 (O_2469,N_48980,N_49394);
or UO_2470 (O_2470,N_49647,N_49935);
or UO_2471 (O_2471,N_49809,N_49552);
nand UO_2472 (O_2472,N_48453,N_48697);
nor UO_2473 (O_2473,N_49036,N_49040);
nand UO_2474 (O_2474,N_47658,N_49313);
and UO_2475 (O_2475,N_49688,N_47656);
or UO_2476 (O_2476,N_49803,N_48531);
xnor UO_2477 (O_2477,N_48863,N_49962);
or UO_2478 (O_2478,N_49802,N_48467);
xnor UO_2479 (O_2479,N_49262,N_47559);
nor UO_2480 (O_2480,N_47906,N_47964);
nor UO_2481 (O_2481,N_48315,N_48668);
or UO_2482 (O_2482,N_48460,N_49307);
and UO_2483 (O_2483,N_47680,N_48730);
or UO_2484 (O_2484,N_49721,N_49806);
nor UO_2485 (O_2485,N_48554,N_48990);
nor UO_2486 (O_2486,N_48197,N_49816);
xnor UO_2487 (O_2487,N_49859,N_48263);
or UO_2488 (O_2488,N_49951,N_49990);
or UO_2489 (O_2489,N_47548,N_49427);
nor UO_2490 (O_2490,N_48428,N_48651);
xor UO_2491 (O_2491,N_48858,N_48632);
or UO_2492 (O_2492,N_49487,N_48210);
and UO_2493 (O_2493,N_47973,N_47884);
or UO_2494 (O_2494,N_48039,N_49050);
nor UO_2495 (O_2495,N_49581,N_49504);
and UO_2496 (O_2496,N_48369,N_49024);
nor UO_2497 (O_2497,N_49374,N_49412);
and UO_2498 (O_2498,N_48167,N_49512);
xnor UO_2499 (O_2499,N_47962,N_47756);
nor UO_2500 (O_2500,N_49749,N_48807);
and UO_2501 (O_2501,N_48817,N_48016);
nand UO_2502 (O_2502,N_49846,N_48406);
or UO_2503 (O_2503,N_49140,N_49737);
and UO_2504 (O_2504,N_49880,N_48215);
or UO_2505 (O_2505,N_48591,N_49441);
and UO_2506 (O_2506,N_48597,N_49572);
and UO_2507 (O_2507,N_48622,N_47715);
xor UO_2508 (O_2508,N_49180,N_48146);
nor UO_2509 (O_2509,N_48226,N_49520);
and UO_2510 (O_2510,N_47577,N_49177);
xor UO_2511 (O_2511,N_48892,N_48380);
nor UO_2512 (O_2512,N_49927,N_48405);
nand UO_2513 (O_2513,N_49919,N_49897);
nor UO_2514 (O_2514,N_47872,N_48355);
or UO_2515 (O_2515,N_47522,N_48233);
nand UO_2516 (O_2516,N_49723,N_47722);
nor UO_2517 (O_2517,N_49273,N_49865);
nor UO_2518 (O_2518,N_48615,N_49896);
xor UO_2519 (O_2519,N_47942,N_48712);
nor UO_2520 (O_2520,N_48961,N_49838);
nand UO_2521 (O_2521,N_47891,N_47991);
and UO_2522 (O_2522,N_49139,N_49733);
and UO_2523 (O_2523,N_49149,N_48238);
xnor UO_2524 (O_2524,N_49809,N_47723);
nor UO_2525 (O_2525,N_49450,N_47934);
nand UO_2526 (O_2526,N_48504,N_47541);
and UO_2527 (O_2527,N_49918,N_47730);
and UO_2528 (O_2528,N_47526,N_49274);
nand UO_2529 (O_2529,N_48594,N_49908);
nor UO_2530 (O_2530,N_49494,N_48899);
or UO_2531 (O_2531,N_48597,N_48551);
and UO_2532 (O_2532,N_49997,N_47748);
nor UO_2533 (O_2533,N_49633,N_49177);
nand UO_2534 (O_2534,N_49138,N_49242);
xnor UO_2535 (O_2535,N_49356,N_49519);
or UO_2536 (O_2536,N_48106,N_49247);
nand UO_2537 (O_2537,N_49865,N_48598);
xor UO_2538 (O_2538,N_49215,N_48271);
or UO_2539 (O_2539,N_49751,N_49078);
or UO_2540 (O_2540,N_49853,N_47797);
and UO_2541 (O_2541,N_49407,N_49439);
xnor UO_2542 (O_2542,N_48267,N_49683);
nand UO_2543 (O_2543,N_47606,N_49992);
xor UO_2544 (O_2544,N_47815,N_48486);
or UO_2545 (O_2545,N_48622,N_49528);
and UO_2546 (O_2546,N_48197,N_48531);
xor UO_2547 (O_2547,N_48771,N_48911);
nand UO_2548 (O_2548,N_49703,N_48925);
xnor UO_2549 (O_2549,N_48960,N_48921);
and UO_2550 (O_2550,N_49096,N_48965);
nor UO_2551 (O_2551,N_49860,N_49548);
and UO_2552 (O_2552,N_49375,N_48271);
nor UO_2553 (O_2553,N_48195,N_48882);
and UO_2554 (O_2554,N_49741,N_49674);
nor UO_2555 (O_2555,N_48962,N_49373);
nand UO_2556 (O_2556,N_48444,N_49650);
xnor UO_2557 (O_2557,N_48089,N_49537);
xor UO_2558 (O_2558,N_49821,N_48187);
or UO_2559 (O_2559,N_49403,N_48547);
nand UO_2560 (O_2560,N_48281,N_47600);
xnor UO_2561 (O_2561,N_48335,N_48982);
and UO_2562 (O_2562,N_48506,N_49412);
nand UO_2563 (O_2563,N_49065,N_48761);
or UO_2564 (O_2564,N_49998,N_49778);
or UO_2565 (O_2565,N_48705,N_48976);
xor UO_2566 (O_2566,N_47595,N_49781);
or UO_2567 (O_2567,N_49640,N_49246);
nand UO_2568 (O_2568,N_47698,N_48376);
and UO_2569 (O_2569,N_49815,N_48097);
or UO_2570 (O_2570,N_48569,N_48762);
nand UO_2571 (O_2571,N_48609,N_47738);
nor UO_2572 (O_2572,N_49282,N_47684);
and UO_2573 (O_2573,N_48734,N_49244);
and UO_2574 (O_2574,N_48481,N_47819);
nand UO_2575 (O_2575,N_48329,N_47925);
or UO_2576 (O_2576,N_49075,N_47744);
nor UO_2577 (O_2577,N_49197,N_48902);
nor UO_2578 (O_2578,N_48549,N_48398);
or UO_2579 (O_2579,N_49354,N_48769);
nor UO_2580 (O_2580,N_48745,N_49931);
xor UO_2581 (O_2581,N_47753,N_48139);
nor UO_2582 (O_2582,N_48201,N_48268);
nand UO_2583 (O_2583,N_47720,N_49930);
xor UO_2584 (O_2584,N_48814,N_48944);
nand UO_2585 (O_2585,N_48549,N_49036);
nor UO_2586 (O_2586,N_48037,N_48878);
xor UO_2587 (O_2587,N_49484,N_47688);
or UO_2588 (O_2588,N_48293,N_47941);
nor UO_2589 (O_2589,N_47949,N_49682);
and UO_2590 (O_2590,N_48720,N_49476);
nand UO_2591 (O_2591,N_48577,N_47894);
or UO_2592 (O_2592,N_48649,N_49811);
and UO_2593 (O_2593,N_49940,N_48092);
or UO_2594 (O_2594,N_49360,N_49318);
xor UO_2595 (O_2595,N_49500,N_49700);
or UO_2596 (O_2596,N_48124,N_49576);
nand UO_2597 (O_2597,N_49939,N_49953);
xnor UO_2598 (O_2598,N_48275,N_49780);
nor UO_2599 (O_2599,N_48868,N_49513);
nor UO_2600 (O_2600,N_48105,N_49140);
nand UO_2601 (O_2601,N_49444,N_49854);
nor UO_2602 (O_2602,N_49039,N_49054);
xnor UO_2603 (O_2603,N_48698,N_48631);
nor UO_2604 (O_2604,N_48975,N_48808);
and UO_2605 (O_2605,N_49171,N_49873);
nand UO_2606 (O_2606,N_48059,N_47964);
xnor UO_2607 (O_2607,N_49018,N_49174);
or UO_2608 (O_2608,N_49975,N_47909);
nor UO_2609 (O_2609,N_49462,N_47938);
and UO_2610 (O_2610,N_48602,N_49145);
xor UO_2611 (O_2611,N_48908,N_48983);
nor UO_2612 (O_2612,N_48907,N_49743);
or UO_2613 (O_2613,N_47626,N_47797);
xor UO_2614 (O_2614,N_49272,N_47539);
and UO_2615 (O_2615,N_48744,N_48091);
and UO_2616 (O_2616,N_49658,N_48398);
nor UO_2617 (O_2617,N_49031,N_48615);
nor UO_2618 (O_2618,N_49103,N_48058);
xnor UO_2619 (O_2619,N_48066,N_48087);
and UO_2620 (O_2620,N_47968,N_48019);
xor UO_2621 (O_2621,N_48107,N_48644);
nand UO_2622 (O_2622,N_48151,N_48318);
or UO_2623 (O_2623,N_48176,N_48128);
or UO_2624 (O_2624,N_48318,N_47831);
xor UO_2625 (O_2625,N_47686,N_49448);
and UO_2626 (O_2626,N_47585,N_48863);
nand UO_2627 (O_2627,N_48683,N_48547);
nand UO_2628 (O_2628,N_48117,N_47714);
xor UO_2629 (O_2629,N_47697,N_48111);
xor UO_2630 (O_2630,N_49914,N_47746);
xor UO_2631 (O_2631,N_48633,N_49211);
or UO_2632 (O_2632,N_48009,N_49488);
nand UO_2633 (O_2633,N_49151,N_47665);
nor UO_2634 (O_2634,N_49230,N_49019);
nand UO_2635 (O_2635,N_48843,N_48399);
or UO_2636 (O_2636,N_49825,N_48994);
nand UO_2637 (O_2637,N_48445,N_48833);
and UO_2638 (O_2638,N_49151,N_49247);
xnor UO_2639 (O_2639,N_48188,N_48335);
nand UO_2640 (O_2640,N_48915,N_48787);
xor UO_2641 (O_2641,N_47550,N_47957);
and UO_2642 (O_2642,N_47725,N_49846);
and UO_2643 (O_2643,N_47881,N_48602);
nand UO_2644 (O_2644,N_49001,N_47803);
or UO_2645 (O_2645,N_49214,N_48535);
nor UO_2646 (O_2646,N_49955,N_49703);
nand UO_2647 (O_2647,N_48094,N_48500);
and UO_2648 (O_2648,N_49735,N_47739);
nand UO_2649 (O_2649,N_48121,N_48756);
and UO_2650 (O_2650,N_48759,N_49476);
xor UO_2651 (O_2651,N_47898,N_49465);
and UO_2652 (O_2652,N_47609,N_48305);
or UO_2653 (O_2653,N_49119,N_49088);
or UO_2654 (O_2654,N_49215,N_49508);
nor UO_2655 (O_2655,N_48460,N_48485);
xnor UO_2656 (O_2656,N_47635,N_48238);
nor UO_2657 (O_2657,N_49488,N_47833);
and UO_2658 (O_2658,N_49906,N_48746);
or UO_2659 (O_2659,N_48071,N_47927);
nor UO_2660 (O_2660,N_48640,N_49504);
nand UO_2661 (O_2661,N_49558,N_48923);
nor UO_2662 (O_2662,N_48890,N_49561);
or UO_2663 (O_2663,N_49788,N_48738);
nor UO_2664 (O_2664,N_47972,N_48732);
nor UO_2665 (O_2665,N_48133,N_49684);
nand UO_2666 (O_2666,N_48480,N_49614);
and UO_2667 (O_2667,N_48750,N_49192);
nor UO_2668 (O_2668,N_49736,N_49452);
or UO_2669 (O_2669,N_47764,N_49648);
and UO_2670 (O_2670,N_49070,N_47617);
or UO_2671 (O_2671,N_47976,N_47631);
nor UO_2672 (O_2672,N_49875,N_48666);
nor UO_2673 (O_2673,N_47917,N_47868);
and UO_2674 (O_2674,N_48979,N_47696);
xnor UO_2675 (O_2675,N_48900,N_48044);
or UO_2676 (O_2676,N_47925,N_47764);
xor UO_2677 (O_2677,N_48242,N_47541);
nand UO_2678 (O_2678,N_49781,N_49289);
and UO_2679 (O_2679,N_47899,N_48614);
or UO_2680 (O_2680,N_49125,N_47580);
nor UO_2681 (O_2681,N_48265,N_49428);
nand UO_2682 (O_2682,N_47686,N_48128);
or UO_2683 (O_2683,N_49855,N_48055);
and UO_2684 (O_2684,N_48895,N_47902);
nand UO_2685 (O_2685,N_48693,N_49118);
and UO_2686 (O_2686,N_48635,N_49458);
nand UO_2687 (O_2687,N_48294,N_49697);
xnor UO_2688 (O_2688,N_47565,N_47757);
nor UO_2689 (O_2689,N_49973,N_49620);
xor UO_2690 (O_2690,N_48269,N_49138);
xnor UO_2691 (O_2691,N_48884,N_49874);
nor UO_2692 (O_2692,N_49065,N_48865);
nor UO_2693 (O_2693,N_48880,N_49360);
nor UO_2694 (O_2694,N_49143,N_49862);
and UO_2695 (O_2695,N_47982,N_48210);
nor UO_2696 (O_2696,N_48001,N_48943);
and UO_2697 (O_2697,N_48753,N_48169);
nand UO_2698 (O_2698,N_48403,N_49021);
nor UO_2699 (O_2699,N_49693,N_47694);
nor UO_2700 (O_2700,N_48765,N_47897);
nand UO_2701 (O_2701,N_48716,N_48681);
xor UO_2702 (O_2702,N_49835,N_47880);
or UO_2703 (O_2703,N_49615,N_49437);
nor UO_2704 (O_2704,N_47727,N_49629);
nor UO_2705 (O_2705,N_49711,N_48052);
nor UO_2706 (O_2706,N_49980,N_48627);
and UO_2707 (O_2707,N_48382,N_48149);
nand UO_2708 (O_2708,N_49499,N_49805);
and UO_2709 (O_2709,N_49740,N_49888);
xnor UO_2710 (O_2710,N_49174,N_49932);
xor UO_2711 (O_2711,N_47988,N_49237);
xor UO_2712 (O_2712,N_49866,N_49935);
and UO_2713 (O_2713,N_47566,N_48276);
and UO_2714 (O_2714,N_47506,N_48873);
nand UO_2715 (O_2715,N_47730,N_49401);
and UO_2716 (O_2716,N_48099,N_48501);
nand UO_2717 (O_2717,N_48828,N_49148);
nand UO_2718 (O_2718,N_49649,N_48266);
or UO_2719 (O_2719,N_48575,N_49853);
xor UO_2720 (O_2720,N_47994,N_49136);
nor UO_2721 (O_2721,N_49317,N_47948);
or UO_2722 (O_2722,N_49834,N_48458);
or UO_2723 (O_2723,N_48910,N_49761);
nand UO_2724 (O_2724,N_48289,N_48073);
xor UO_2725 (O_2725,N_49732,N_47947);
and UO_2726 (O_2726,N_48041,N_49173);
xnor UO_2727 (O_2727,N_48350,N_49839);
xnor UO_2728 (O_2728,N_49827,N_49620);
and UO_2729 (O_2729,N_48846,N_49141);
or UO_2730 (O_2730,N_48209,N_49394);
nor UO_2731 (O_2731,N_48280,N_49392);
and UO_2732 (O_2732,N_48577,N_49263);
nor UO_2733 (O_2733,N_48147,N_48070);
nor UO_2734 (O_2734,N_47786,N_48430);
nand UO_2735 (O_2735,N_49419,N_48878);
nor UO_2736 (O_2736,N_48603,N_49235);
nor UO_2737 (O_2737,N_49711,N_48990);
nand UO_2738 (O_2738,N_49066,N_47760);
nor UO_2739 (O_2739,N_49028,N_49123);
xnor UO_2740 (O_2740,N_47562,N_48714);
or UO_2741 (O_2741,N_48925,N_48251);
xor UO_2742 (O_2742,N_49063,N_49866);
xnor UO_2743 (O_2743,N_47600,N_49897);
nor UO_2744 (O_2744,N_49793,N_47578);
and UO_2745 (O_2745,N_47875,N_48526);
nand UO_2746 (O_2746,N_49150,N_49063);
nor UO_2747 (O_2747,N_49007,N_48889);
or UO_2748 (O_2748,N_47916,N_49074);
nand UO_2749 (O_2749,N_49395,N_48977);
or UO_2750 (O_2750,N_49573,N_49875);
xor UO_2751 (O_2751,N_49125,N_47867);
nor UO_2752 (O_2752,N_49516,N_47988);
nor UO_2753 (O_2753,N_47722,N_49206);
or UO_2754 (O_2754,N_49772,N_48524);
or UO_2755 (O_2755,N_47766,N_48087);
nand UO_2756 (O_2756,N_48934,N_48420);
nand UO_2757 (O_2757,N_49946,N_48775);
and UO_2758 (O_2758,N_47899,N_48927);
or UO_2759 (O_2759,N_48208,N_48875);
nor UO_2760 (O_2760,N_49346,N_48250);
and UO_2761 (O_2761,N_47741,N_49826);
nand UO_2762 (O_2762,N_49209,N_49658);
nor UO_2763 (O_2763,N_48943,N_47869);
or UO_2764 (O_2764,N_48452,N_49364);
nand UO_2765 (O_2765,N_49457,N_47831);
nand UO_2766 (O_2766,N_49593,N_49148);
and UO_2767 (O_2767,N_48445,N_48819);
xnor UO_2768 (O_2768,N_48207,N_48677);
xnor UO_2769 (O_2769,N_48470,N_49726);
nand UO_2770 (O_2770,N_49796,N_48805);
and UO_2771 (O_2771,N_49455,N_49422);
and UO_2772 (O_2772,N_49664,N_48624);
nor UO_2773 (O_2773,N_48538,N_48343);
nor UO_2774 (O_2774,N_49375,N_48493);
xor UO_2775 (O_2775,N_48717,N_48614);
xnor UO_2776 (O_2776,N_49429,N_49751);
and UO_2777 (O_2777,N_49925,N_48902);
nand UO_2778 (O_2778,N_49214,N_49037);
nor UO_2779 (O_2779,N_49449,N_48009);
or UO_2780 (O_2780,N_49662,N_47825);
nand UO_2781 (O_2781,N_47794,N_48685);
xnor UO_2782 (O_2782,N_49079,N_49825);
nand UO_2783 (O_2783,N_47643,N_49097);
nand UO_2784 (O_2784,N_49192,N_49680);
nor UO_2785 (O_2785,N_49316,N_48748);
xor UO_2786 (O_2786,N_49734,N_47597);
nand UO_2787 (O_2787,N_49838,N_48026);
nor UO_2788 (O_2788,N_49849,N_47738);
nor UO_2789 (O_2789,N_49660,N_49925);
nor UO_2790 (O_2790,N_49217,N_49805);
nand UO_2791 (O_2791,N_48079,N_49509);
xnor UO_2792 (O_2792,N_48103,N_48654);
or UO_2793 (O_2793,N_47806,N_48232);
xnor UO_2794 (O_2794,N_48435,N_48640);
xnor UO_2795 (O_2795,N_47724,N_49153);
nand UO_2796 (O_2796,N_48852,N_49158);
nor UO_2797 (O_2797,N_49435,N_49264);
and UO_2798 (O_2798,N_47997,N_48147);
or UO_2799 (O_2799,N_49039,N_49196);
or UO_2800 (O_2800,N_48003,N_48828);
xor UO_2801 (O_2801,N_49850,N_47741);
nor UO_2802 (O_2802,N_49647,N_48894);
and UO_2803 (O_2803,N_48953,N_49368);
and UO_2804 (O_2804,N_48213,N_48850);
xor UO_2805 (O_2805,N_49619,N_48164);
nor UO_2806 (O_2806,N_49261,N_49995);
nor UO_2807 (O_2807,N_48422,N_47703);
and UO_2808 (O_2808,N_49842,N_48528);
or UO_2809 (O_2809,N_49249,N_48640);
xnor UO_2810 (O_2810,N_49859,N_47511);
nand UO_2811 (O_2811,N_49832,N_49961);
and UO_2812 (O_2812,N_47880,N_48227);
nor UO_2813 (O_2813,N_48786,N_48627);
nor UO_2814 (O_2814,N_47717,N_49162);
and UO_2815 (O_2815,N_49042,N_49521);
nor UO_2816 (O_2816,N_47660,N_49717);
and UO_2817 (O_2817,N_48966,N_48241);
or UO_2818 (O_2818,N_47983,N_47715);
nand UO_2819 (O_2819,N_49295,N_49775);
xor UO_2820 (O_2820,N_47511,N_47816);
nor UO_2821 (O_2821,N_49420,N_49569);
nand UO_2822 (O_2822,N_48129,N_49407);
or UO_2823 (O_2823,N_49425,N_49292);
nand UO_2824 (O_2824,N_48882,N_49815);
and UO_2825 (O_2825,N_47804,N_49220);
xnor UO_2826 (O_2826,N_48449,N_47668);
nor UO_2827 (O_2827,N_48717,N_48087);
nand UO_2828 (O_2828,N_47704,N_47569);
xor UO_2829 (O_2829,N_49583,N_49675);
and UO_2830 (O_2830,N_48676,N_49749);
xnor UO_2831 (O_2831,N_48879,N_48511);
and UO_2832 (O_2832,N_49443,N_48834);
nor UO_2833 (O_2833,N_47904,N_47764);
xnor UO_2834 (O_2834,N_49941,N_48900);
nand UO_2835 (O_2835,N_47904,N_47512);
xor UO_2836 (O_2836,N_48209,N_48499);
nand UO_2837 (O_2837,N_47565,N_48061);
nand UO_2838 (O_2838,N_47654,N_49616);
and UO_2839 (O_2839,N_49056,N_47546);
or UO_2840 (O_2840,N_49586,N_48787);
or UO_2841 (O_2841,N_49715,N_48946);
nand UO_2842 (O_2842,N_49016,N_48072);
or UO_2843 (O_2843,N_48457,N_49006);
and UO_2844 (O_2844,N_48232,N_48570);
nand UO_2845 (O_2845,N_49674,N_47805);
nor UO_2846 (O_2846,N_48606,N_49387);
or UO_2847 (O_2847,N_49429,N_48531);
and UO_2848 (O_2848,N_48939,N_49653);
or UO_2849 (O_2849,N_47549,N_49835);
xor UO_2850 (O_2850,N_49181,N_47795);
xnor UO_2851 (O_2851,N_49984,N_48986);
nor UO_2852 (O_2852,N_49198,N_48511);
nor UO_2853 (O_2853,N_48428,N_49566);
nand UO_2854 (O_2854,N_47516,N_49214);
nand UO_2855 (O_2855,N_48838,N_49259);
and UO_2856 (O_2856,N_47684,N_49743);
nand UO_2857 (O_2857,N_49777,N_47653);
xnor UO_2858 (O_2858,N_47576,N_48262);
xnor UO_2859 (O_2859,N_48379,N_49267);
or UO_2860 (O_2860,N_48397,N_49720);
nand UO_2861 (O_2861,N_48053,N_48013);
or UO_2862 (O_2862,N_49015,N_47616);
nor UO_2863 (O_2863,N_47518,N_49911);
or UO_2864 (O_2864,N_47655,N_49861);
or UO_2865 (O_2865,N_48039,N_48095);
and UO_2866 (O_2866,N_48764,N_48647);
and UO_2867 (O_2867,N_49131,N_48943);
xnor UO_2868 (O_2868,N_48094,N_48273);
and UO_2869 (O_2869,N_49971,N_48740);
nand UO_2870 (O_2870,N_48690,N_48634);
xor UO_2871 (O_2871,N_48761,N_48341);
or UO_2872 (O_2872,N_47793,N_48698);
xor UO_2873 (O_2873,N_48886,N_48355);
and UO_2874 (O_2874,N_48153,N_47720);
nand UO_2875 (O_2875,N_48649,N_48887);
and UO_2876 (O_2876,N_48821,N_49776);
or UO_2877 (O_2877,N_47751,N_49741);
nand UO_2878 (O_2878,N_48482,N_47791);
nor UO_2879 (O_2879,N_49906,N_47876);
or UO_2880 (O_2880,N_48560,N_49749);
xnor UO_2881 (O_2881,N_48434,N_49097);
and UO_2882 (O_2882,N_48075,N_49303);
xor UO_2883 (O_2883,N_48112,N_47520);
xor UO_2884 (O_2884,N_47848,N_48899);
xnor UO_2885 (O_2885,N_49903,N_47767);
or UO_2886 (O_2886,N_49054,N_48818);
xor UO_2887 (O_2887,N_47905,N_48336);
or UO_2888 (O_2888,N_48979,N_48652);
and UO_2889 (O_2889,N_49887,N_48503);
nor UO_2890 (O_2890,N_49653,N_47964);
and UO_2891 (O_2891,N_47520,N_49788);
xor UO_2892 (O_2892,N_47858,N_47601);
nor UO_2893 (O_2893,N_48648,N_48473);
xnor UO_2894 (O_2894,N_48048,N_49522);
nor UO_2895 (O_2895,N_49054,N_47908);
nand UO_2896 (O_2896,N_48579,N_48996);
nand UO_2897 (O_2897,N_48388,N_49243);
or UO_2898 (O_2898,N_47706,N_47885);
nor UO_2899 (O_2899,N_48257,N_49044);
nand UO_2900 (O_2900,N_49236,N_49968);
or UO_2901 (O_2901,N_49094,N_49895);
nor UO_2902 (O_2902,N_48672,N_49474);
and UO_2903 (O_2903,N_49146,N_48443);
xor UO_2904 (O_2904,N_47549,N_48983);
and UO_2905 (O_2905,N_47556,N_49253);
and UO_2906 (O_2906,N_49813,N_48058);
nand UO_2907 (O_2907,N_47634,N_48104);
xnor UO_2908 (O_2908,N_48649,N_49931);
xor UO_2909 (O_2909,N_47621,N_48186);
nor UO_2910 (O_2910,N_48745,N_47762);
nor UO_2911 (O_2911,N_49996,N_47958);
nand UO_2912 (O_2912,N_49505,N_48329);
or UO_2913 (O_2913,N_49891,N_47988);
nand UO_2914 (O_2914,N_48944,N_48853);
and UO_2915 (O_2915,N_48019,N_48164);
xnor UO_2916 (O_2916,N_49168,N_49251);
nor UO_2917 (O_2917,N_48191,N_47754);
nand UO_2918 (O_2918,N_49393,N_49983);
xor UO_2919 (O_2919,N_48526,N_47971);
or UO_2920 (O_2920,N_47769,N_47917);
xor UO_2921 (O_2921,N_49124,N_48062);
nand UO_2922 (O_2922,N_48338,N_47512);
nand UO_2923 (O_2923,N_48612,N_47907);
nand UO_2924 (O_2924,N_49985,N_48354);
and UO_2925 (O_2925,N_47963,N_48837);
nand UO_2926 (O_2926,N_47972,N_49464);
nand UO_2927 (O_2927,N_49486,N_49576);
and UO_2928 (O_2928,N_49341,N_49102);
xnor UO_2929 (O_2929,N_49275,N_47735);
and UO_2930 (O_2930,N_49015,N_47610);
and UO_2931 (O_2931,N_48900,N_47868);
and UO_2932 (O_2932,N_47809,N_48826);
xnor UO_2933 (O_2933,N_48820,N_49913);
or UO_2934 (O_2934,N_49100,N_49180);
nor UO_2935 (O_2935,N_48242,N_49543);
nand UO_2936 (O_2936,N_48228,N_49129);
and UO_2937 (O_2937,N_47665,N_49105);
nand UO_2938 (O_2938,N_47500,N_47651);
nor UO_2939 (O_2939,N_48050,N_48362);
and UO_2940 (O_2940,N_49682,N_48719);
xnor UO_2941 (O_2941,N_48112,N_48382);
nor UO_2942 (O_2942,N_48395,N_48056);
nor UO_2943 (O_2943,N_49736,N_48792);
nor UO_2944 (O_2944,N_49336,N_48838);
nor UO_2945 (O_2945,N_47829,N_49039);
xor UO_2946 (O_2946,N_49684,N_47519);
or UO_2947 (O_2947,N_48843,N_49724);
nand UO_2948 (O_2948,N_47587,N_48054);
nor UO_2949 (O_2949,N_48272,N_47558);
or UO_2950 (O_2950,N_49864,N_48346);
or UO_2951 (O_2951,N_49759,N_48109);
and UO_2952 (O_2952,N_49578,N_48299);
and UO_2953 (O_2953,N_47585,N_49136);
nor UO_2954 (O_2954,N_47634,N_49593);
nand UO_2955 (O_2955,N_48223,N_48126);
and UO_2956 (O_2956,N_49143,N_49521);
nand UO_2957 (O_2957,N_49096,N_48785);
or UO_2958 (O_2958,N_48223,N_48505);
nand UO_2959 (O_2959,N_49880,N_48027);
or UO_2960 (O_2960,N_47815,N_48480);
or UO_2961 (O_2961,N_49847,N_48082);
nor UO_2962 (O_2962,N_47707,N_47742);
or UO_2963 (O_2963,N_48779,N_49670);
and UO_2964 (O_2964,N_48657,N_49552);
or UO_2965 (O_2965,N_49298,N_49513);
and UO_2966 (O_2966,N_48384,N_49622);
and UO_2967 (O_2967,N_49122,N_49210);
nand UO_2968 (O_2968,N_49267,N_48937);
and UO_2969 (O_2969,N_49659,N_47763);
xnor UO_2970 (O_2970,N_48776,N_47939);
xnor UO_2971 (O_2971,N_47847,N_48655);
or UO_2972 (O_2972,N_48290,N_48177);
nand UO_2973 (O_2973,N_48327,N_49678);
and UO_2974 (O_2974,N_48080,N_47589);
xor UO_2975 (O_2975,N_48760,N_49210);
or UO_2976 (O_2976,N_47909,N_49720);
xnor UO_2977 (O_2977,N_48613,N_47656);
or UO_2978 (O_2978,N_49461,N_48438);
and UO_2979 (O_2979,N_49287,N_48687);
nor UO_2980 (O_2980,N_49410,N_49649);
nor UO_2981 (O_2981,N_49472,N_47526);
nand UO_2982 (O_2982,N_49813,N_49872);
nand UO_2983 (O_2983,N_49361,N_48685);
xor UO_2984 (O_2984,N_48923,N_47963);
xnor UO_2985 (O_2985,N_48545,N_48035);
and UO_2986 (O_2986,N_48632,N_48994);
nand UO_2987 (O_2987,N_49407,N_48976);
xnor UO_2988 (O_2988,N_48574,N_48658);
nand UO_2989 (O_2989,N_48317,N_49143);
xnor UO_2990 (O_2990,N_49841,N_47703);
nor UO_2991 (O_2991,N_48662,N_48078);
xor UO_2992 (O_2992,N_48095,N_48486);
and UO_2993 (O_2993,N_49091,N_48936);
and UO_2994 (O_2994,N_48522,N_49538);
nor UO_2995 (O_2995,N_48265,N_48262);
and UO_2996 (O_2996,N_47526,N_48049);
nor UO_2997 (O_2997,N_48393,N_47748);
nor UO_2998 (O_2998,N_48226,N_49271);
or UO_2999 (O_2999,N_49418,N_48682);
or UO_3000 (O_3000,N_49051,N_49974);
nor UO_3001 (O_3001,N_48442,N_48701);
xor UO_3002 (O_3002,N_47740,N_48157);
and UO_3003 (O_3003,N_49664,N_49110);
nand UO_3004 (O_3004,N_48337,N_47689);
nand UO_3005 (O_3005,N_47764,N_47501);
nand UO_3006 (O_3006,N_48315,N_49671);
or UO_3007 (O_3007,N_48852,N_48723);
nand UO_3008 (O_3008,N_48330,N_49285);
and UO_3009 (O_3009,N_49492,N_49018);
and UO_3010 (O_3010,N_48734,N_49877);
and UO_3011 (O_3011,N_49993,N_49927);
or UO_3012 (O_3012,N_48208,N_49502);
nand UO_3013 (O_3013,N_49198,N_48053);
xnor UO_3014 (O_3014,N_47586,N_48352);
and UO_3015 (O_3015,N_49040,N_47643);
nand UO_3016 (O_3016,N_47869,N_48672);
or UO_3017 (O_3017,N_49796,N_49550);
and UO_3018 (O_3018,N_48752,N_49029);
nor UO_3019 (O_3019,N_49177,N_48967);
xnor UO_3020 (O_3020,N_49807,N_49059);
or UO_3021 (O_3021,N_49111,N_48401);
xor UO_3022 (O_3022,N_48603,N_47884);
xor UO_3023 (O_3023,N_49580,N_48342);
nand UO_3024 (O_3024,N_48547,N_49712);
or UO_3025 (O_3025,N_48262,N_49336);
or UO_3026 (O_3026,N_48158,N_47591);
nor UO_3027 (O_3027,N_49133,N_47703);
and UO_3028 (O_3028,N_48674,N_47569);
nand UO_3029 (O_3029,N_48762,N_48410);
xor UO_3030 (O_3030,N_49980,N_48123);
nand UO_3031 (O_3031,N_48360,N_49991);
and UO_3032 (O_3032,N_47644,N_47739);
xnor UO_3033 (O_3033,N_47931,N_49819);
nor UO_3034 (O_3034,N_49274,N_48851);
nand UO_3035 (O_3035,N_48441,N_49385);
nand UO_3036 (O_3036,N_49131,N_49655);
nor UO_3037 (O_3037,N_49898,N_48291);
xnor UO_3038 (O_3038,N_48452,N_48931);
or UO_3039 (O_3039,N_47556,N_48380);
xnor UO_3040 (O_3040,N_48809,N_48551);
or UO_3041 (O_3041,N_49915,N_47827);
and UO_3042 (O_3042,N_48715,N_48908);
xnor UO_3043 (O_3043,N_49111,N_47898);
nand UO_3044 (O_3044,N_48796,N_48076);
nand UO_3045 (O_3045,N_47589,N_49881);
nor UO_3046 (O_3046,N_48261,N_48297);
nor UO_3047 (O_3047,N_49220,N_48676);
or UO_3048 (O_3048,N_48295,N_49136);
nor UO_3049 (O_3049,N_49942,N_49156);
and UO_3050 (O_3050,N_49437,N_49349);
or UO_3051 (O_3051,N_49592,N_48767);
nor UO_3052 (O_3052,N_47814,N_49807);
nand UO_3053 (O_3053,N_49645,N_49060);
and UO_3054 (O_3054,N_48287,N_49365);
or UO_3055 (O_3055,N_48661,N_47525);
or UO_3056 (O_3056,N_49513,N_48486);
nor UO_3057 (O_3057,N_49267,N_49934);
and UO_3058 (O_3058,N_48901,N_49137);
nor UO_3059 (O_3059,N_48187,N_49361);
or UO_3060 (O_3060,N_48376,N_49128);
xnor UO_3061 (O_3061,N_48498,N_48079);
nor UO_3062 (O_3062,N_49732,N_47904);
and UO_3063 (O_3063,N_48643,N_48167);
nand UO_3064 (O_3064,N_49223,N_49532);
nand UO_3065 (O_3065,N_48702,N_47855);
xnor UO_3066 (O_3066,N_47541,N_47601);
or UO_3067 (O_3067,N_47579,N_48895);
nor UO_3068 (O_3068,N_48195,N_47943);
nor UO_3069 (O_3069,N_48232,N_49417);
and UO_3070 (O_3070,N_49392,N_49294);
nand UO_3071 (O_3071,N_49086,N_49824);
xnor UO_3072 (O_3072,N_49718,N_48760);
nand UO_3073 (O_3073,N_47682,N_49368);
and UO_3074 (O_3074,N_48440,N_49384);
or UO_3075 (O_3075,N_49439,N_49022);
and UO_3076 (O_3076,N_49575,N_48433);
nor UO_3077 (O_3077,N_48819,N_49576);
and UO_3078 (O_3078,N_48215,N_49842);
xor UO_3079 (O_3079,N_48487,N_49950);
and UO_3080 (O_3080,N_49083,N_47564);
nor UO_3081 (O_3081,N_48442,N_49661);
xor UO_3082 (O_3082,N_49975,N_48379);
and UO_3083 (O_3083,N_49736,N_48078);
xor UO_3084 (O_3084,N_47965,N_49654);
or UO_3085 (O_3085,N_49340,N_49982);
nand UO_3086 (O_3086,N_49223,N_48503);
nand UO_3087 (O_3087,N_48894,N_48944);
nor UO_3088 (O_3088,N_49553,N_48767);
xnor UO_3089 (O_3089,N_48305,N_48203);
nor UO_3090 (O_3090,N_48915,N_49449);
xor UO_3091 (O_3091,N_49330,N_47788);
nor UO_3092 (O_3092,N_48174,N_49111);
and UO_3093 (O_3093,N_47645,N_49685);
xor UO_3094 (O_3094,N_49593,N_49028);
or UO_3095 (O_3095,N_47992,N_48340);
and UO_3096 (O_3096,N_48434,N_49784);
nor UO_3097 (O_3097,N_48752,N_49848);
and UO_3098 (O_3098,N_49510,N_48129);
nor UO_3099 (O_3099,N_48889,N_47964);
and UO_3100 (O_3100,N_49593,N_48359);
or UO_3101 (O_3101,N_49051,N_48006);
nand UO_3102 (O_3102,N_48104,N_48637);
and UO_3103 (O_3103,N_49781,N_47635);
and UO_3104 (O_3104,N_48854,N_48308);
nor UO_3105 (O_3105,N_49289,N_48153);
or UO_3106 (O_3106,N_48570,N_48381);
xor UO_3107 (O_3107,N_48207,N_49992);
nand UO_3108 (O_3108,N_47656,N_47977);
xor UO_3109 (O_3109,N_49372,N_48613);
or UO_3110 (O_3110,N_48205,N_48593);
and UO_3111 (O_3111,N_49274,N_48921);
nor UO_3112 (O_3112,N_48105,N_48618);
or UO_3113 (O_3113,N_47506,N_49667);
nand UO_3114 (O_3114,N_49920,N_49154);
nor UO_3115 (O_3115,N_49757,N_48870);
xnor UO_3116 (O_3116,N_48267,N_48772);
or UO_3117 (O_3117,N_49108,N_47541);
xor UO_3118 (O_3118,N_48754,N_48951);
nor UO_3119 (O_3119,N_48114,N_49371);
and UO_3120 (O_3120,N_49160,N_48142);
and UO_3121 (O_3121,N_47987,N_47633);
xor UO_3122 (O_3122,N_48308,N_47966);
nand UO_3123 (O_3123,N_49116,N_49267);
and UO_3124 (O_3124,N_49942,N_47569);
or UO_3125 (O_3125,N_47826,N_48397);
xor UO_3126 (O_3126,N_49458,N_47878);
or UO_3127 (O_3127,N_49139,N_49161);
xor UO_3128 (O_3128,N_49386,N_48487);
nand UO_3129 (O_3129,N_49815,N_49181);
xnor UO_3130 (O_3130,N_47703,N_48731);
and UO_3131 (O_3131,N_47847,N_47651);
xnor UO_3132 (O_3132,N_48274,N_49649);
nor UO_3133 (O_3133,N_47595,N_49744);
nor UO_3134 (O_3134,N_49419,N_48405);
xor UO_3135 (O_3135,N_49361,N_49629);
nor UO_3136 (O_3136,N_49619,N_49761);
and UO_3137 (O_3137,N_48609,N_48015);
nand UO_3138 (O_3138,N_49458,N_47748);
nand UO_3139 (O_3139,N_49633,N_49561);
or UO_3140 (O_3140,N_48788,N_48407);
or UO_3141 (O_3141,N_49833,N_47940);
nand UO_3142 (O_3142,N_49354,N_48414);
and UO_3143 (O_3143,N_47693,N_47537);
xor UO_3144 (O_3144,N_48052,N_48214);
nand UO_3145 (O_3145,N_48835,N_49825);
xor UO_3146 (O_3146,N_48533,N_49293);
nand UO_3147 (O_3147,N_47803,N_48804);
or UO_3148 (O_3148,N_48479,N_48727);
and UO_3149 (O_3149,N_48048,N_49475);
and UO_3150 (O_3150,N_47777,N_49981);
or UO_3151 (O_3151,N_49154,N_48262);
nor UO_3152 (O_3152,N_48979,N_49506);
xor UO_3153 (O_3153,N_49084,N_48933);
xnor UO_3154 (O_3154,N_49639,N_49537);
and UO_3155 (O_3155,N_49179,N_47794);
or UO_3156 (O_3156,N_48335,N_47508);
or UO_3157 (O_3157,N_49938,N_49755);
and UO_3158 (O_3158,N_48189,N_49853);
and UO_3159 (O_3159,N_48188,N_47938);
and UO_3160 (O_3160,N_49111,N_49277);
and UO_3161 (O_3161,N_49824,N_48079);
or UO_3162 (O_3162,N_47763,N_47905);
xnor UO_3163 (O_3163,N_49148,N_48053);
xnor UO_3164 (O_3164,N_48033,N_48731);
and UO_3165 (O_3165,N_47803,N_49209);
nor UO_3166 (O_3166,N_49529,N_47719);
or UO_3167 (O_3167,N_47616,N_47551);
xor UO_3168 (O_3168,N_48692,N_47549);
xnor UO_3169 (O_3169,N_48262,N_47945);
nor UO_3170 (O_3170,N_49060,N_47593);
nand UO_3171 (O_3171,N_49675,N_49994);
nand UO_3172 (O_3172,N_48462,N_49216);
nand UO_3173 (O_3173,N_49594,N_47621);
nor UO_3174 (O_3174,N_48479,N_48283);
nor UO_3175 (O_3175,N_47717,N_48948);
or UO_3176 (O_3176,N_47649,N_48016);
nor UO_3177 (O_3177,N_49911,N_48147);
nor UO_3178 (O_3178,N_49466,N_48936);
or UO_3179 (O_3179,N_49457,N_48496);
nor UO_3180 (O_3180,N_48845,N_48813);
or UO_3181 (O_3181,N_48358,N_48938);
xnor UO_3182 (O_3182,N_49386,N_48752);
nand UO_3183 (O_3183,N_48630,N_48080);
nand UO_3184 (O_3184,N_47855,N_48679);
xor UO_3185 (O_3185,N_49174,N_47901);
and UO_3186 (O_3186,N_48908,N_48984);
xnor UO_3187 (O_3187,N_47717,N_47551);
or UO_3188 (O_3188,N_49052,N_48339);
nand UO_3189 (O_3189,N_49041,N_48485);
nor UO_3190 (O_3190,N_48242,N_47766);
nor UO_3191 (O_3191,N_49483,N_49033);
or UO_3192 (O_3192,N_49049,N_48181);
nand UO_3193 (O_3193,N_48329,N_49159);
or UO_3194 (O_3194,N_48763,N_49057);
or UO_3195 (O_3195,N_48384,N_47655);
nand UO_3196 (O_3196,N_47841,N_49414);
and UO_3197 (O_3197,N_49238,N_48062);
or UO_3198 (O_3198,N_49565,N_49756);
and UO_3199 (O_3199,N_49885,N_49931);
or UO_3200 (O_3200,N_47547,N_49700);
xor UO_3201 (O_3201,N_47835,N_48599);
and UO_3202 (O_3202,N_48296,N_47869);
xor UO_3203 (O_3203,N_49841,N_49727);
nand UO_3204 (O_3204,N_49255,N_48666);
nor UO_3205 (O_3205,N_48027,N_48455);
nand UO_3206 (O_3206,N_47744,N_48872);
xor UO_3207 (O_3207,N_49417,N_47528);
nand UO_3208 (O_3208,N_48769,N_49758);
or UO_3209 (O_3209,N_48710,N_49273);
and UO_3210 (O_3210,N_48499,N_49890);
or UO_3211 (O_3211,N_48385,N_48850);
and UO_3212 (O_3212,N_49140,N_48580);
nand UO_3213 (O_3213,N_49530,N_48130);
or UO_3214 (O_3214,N_48274,N_48386);
nor UO_3215 (O_3215,N_48347,N_48654);
and UO_3216 (O_3216,N_49933,N_48157);
or UO_3217 (O_3217,N_47877,N_47874);
nand UO_3218 (O_3218,N_47565,N_48736);
nor UO_3219 (O_3219,N_49194,N_47910);
nor UO_3220 (O_3220,N_48003,N_49336);
nand UO_3221 (O_3221,N_47923,N_49859);
or UO_3222 (O_3222,N_47525,N_48952);
and UO_3223 (O_3223,N_48775,N_49056);
xnor UO_3224 (O_3224,N_48594,N_49968);
and UO_3225 (O_3225,N_47648,N_49768);
nor UO_3226 (O_3226,N_49036,N_47726);
and UO_3227 (O_3227,N_48325,N_49744);
xnor UO_3228 (O_3228,N_48616,N_49487);
or UO_3229 (O_3229,N_48612,N_48287);
and UO_3230 (O_3230,N_49331,N_48296);
and UO_3231 (O_3231,N_49455,N_47701);
xnor UO_3232 (O_3232,N_49381,N_48893);
nand UO_3233 (O_3233,N_48764,N_48232);
nor UO_3234 (O_3234,N_49996,N_47737);
and UO_3235 (O_3235,N_49236,N_49923);
or UO_3236 (O_3236,N_49115,N_49396);
nor UO_3237 (O_3237,N_48322,N_49996);
xor UO_3238 (O_3238,N_47602,N_48634);
nor UO_3239 (O_3239,N_49914,N_48868);
nand UO_3240 (O_3240,N_48108,N_49547);
and UO_3241 (O_3241,N_49254,N_47991);
xor UO_3242 (O_3242,N_49643,N_49994);
or UO_3243 (O_3243,N_49793,N_48983);
nand UO_3244 (O_3244,N_48274,N_48628);
nor UO_3245 (O_3245,N_48944,N_48081);
xnor UO_3246 (O_3246,N_49264,N_49041);
and UO_3247 (O_3247,N_49521,N_49961);
nand UO_3248 (O_3248,N_49483,N_48543);
nand UO_3249 (O_3249,N_49594,N_49373);
and UO_3250 (O_3250,N_49219,N_49004);
or UO_3251 (O_3251,N_48822,N_49935);
nand UO_3252 (O_3252,N_48661,N_48948);
or UO_3253 (O_3253,N_48145,N_48472);
and UO_3254 (O_3254,N_48913,N_49844);
nor UO_3255 (O_3255,N_48062,N_47746);
nor UO_3256 (O_3256,N_48776,N_48469);
xor UO_3257 (O_3257,N_48657,N_48832);
or UO_3258 (O_3258,N_48020,N_48605);
and UO_3259 (O_3259,N_48801,N_48787);
or UO_3260 (O_3260,N_48944,N_49037);
nand UO_3261 (O_3261,N_48093,N_48876);
or UO_3262 (O_3262,N_49717,N_49893);
or UO_3263 (O_3263,N_48678,N_49735);
and UO_3264 (O_3264,N_49912,N_47758);
and UO_3265 (O_3265,N_48597,N_48464);
nor UO_3266 (O_3266,N_48888,N_49481);
xnor UO_3267 (O_3267,N_49925,N_48524);
or UO_3268 (O_3268,N_48363,N_47530);
and UO_3269 (O_3269,N_49372,N_49633);
and UO_3270 (O_3270,N_48135,N_49802);
nor UO_3271 (O_3271,N_48826,N_49038);
or UO_3272 (O_3272,N_47809,N_48932);
nor UO_3273 (O_3273,N_47518,N_49436);
nor UO_3274 (O_3274,N_49058,N_49867);
nor UO_3275 (O_3275,N_48496,N_49755);
and UO_3276 (O_3276,N_48190,N_48899);
xnor UO_3277 (O_3277,N_48675,N_49272);
nor UO_3278 (O_3278,N_47801,N_49220);
nor UO_3279 (O_3279,N_48390,N_49518);
xnor UO_3280 (O_3280,N_48272,N_48295);
nand UO_3281 (O_3281,N_49994,N_49671);
and UO_3282 (O_3282,N_48936,N_48867);
xnor UO_3283 (O_3283,N_47911,N_48860);
nand UO_3284 (O_3284,N_47916,N_47512);
and UO_3285 (O_3285,N_49840,N_48133);
or UO_3286 (O_3286,N_48044,N_48815);
nor UO_3287 (O_3287,N_48836,N_48532);
xnor UO_3288 (O_3288,N_49077,N_48296);
nor UO_3289 (O_3289,N_47645,N_48476);
nand UO_3290 (O_3290,N_48550,N_48127);
nor UO_3291 (O_3291,N_48163,N_49492);
xnor UO_3292 (O_3292,N_48714,N_49232);
nand UO_3293 (O_3293,N_47810,N_47643);
xor UO_3294 (O_3294,N_49089,N_49825);
nand UO_3295 (O_3295,N_49671,N_48264);
nand UO_3296 (O_3296,N_48357,N_49923);
and UO_3297 (O_3297,N_47958,N_48660);
nand UO_3298 (O_3298,N_47614,N_48146);
xnor UO_3299 (O_3299,N_49216,N_49799);
and UO_3300 (O_3300,N_48881,N_49023);
or UO_3301 (O_3301,N_49553,N_48182);
or UO_3302 (O_3302,N_48611,N_49208);
or UO_3303 (O_3303,N_49048,N_49576);
nand UO_3304 (O_3304,N_48232,N_47759);
xnor UO_3305 (O_3305,N_48448,N_48686);
nor UO_3306 (O_3306,N_49014,N_49351);
and UO_3307 (O_3307,N_48156,N_49241);
nand UO_3308 (O_3308,N_48601,N_48763);
nand UO_3309 (O_3309,N_49302,N_47662);
nor UO_3310 (O_3310,N_49025,N_48454);
nand UO_3311 (O_3311,N_47718,N_47502);
and UO_3312 (O_3312,N_48206,N_48427);
xor UO_3313 (O_3313,N_49134,N_48655);
and UO_3314 (O_3314,N_49031,N_48268);
or UO_3315 (O_3315,N_47617,N_49019);
and UO_3316 (O_3316,N_49169,N_48274);
and UO_3317 (O_3317,N_49489,N_47638);
nand UO_3318 (O_3318,N_49611,N_49449);
and UO_3319 (O_3319,N_47657,N_49293);
or UO_3320 (O_3320,N_49085,N_49419);
nand UO_3321 (O_3321,N_48151,N_49443);
nand UO_3322 (O_3322,N_48585,N_49509);
nand UO_3323 (O_3323,N_48313,N_47673);
xnor UO_3324 (O_3324,N_47787,N_49972);
or UO_3325 (O_3325,N_49333,N_48026);
xnor UO_3326 (O_3326,N_48012,N_48522);
or UO_3327 (O_3327,N_47641,N_49193);
nand UO_3328 (O_3328,N_49396,N_48687);
and UO_3329 (O_3329,N_49179,N_47925);
nor UO_3330 (O_3330,N_48540,N_48158);
or UO_3331 (O_3331,N_48843,N_48272);
and UO_3332 (O_3332,N_49707,N_47785);
and UO_3333 (O_3333,N_47606,N_49052);
and UO_3334 (O_3334,N_48470,N_47892);
nand UO_3335 (O_3335,N_49525,N_48181);
or UO_3336 (O_3336,N_49538,N_49689);
or UO_3337 (O_3337,N_48943,N_48328);
or UO_3338 (O_3338,N_49282,N_48731);
or UO_3339 (O_3339,N_49978,N_49830);
xor UO_3340 (O_3340,N_49827,N_48838);
and UO_3341 (O_3341,N_48242,N_48147);
nor UO_3342 (O_3342,N_49817,N_48628);
nand UO_3343 (O_3343,N_47515,N_48977);
and UO_3344 (O_3344,N_48575,N_48549);
or UO_3345 (O_3345,N_48143,N_49704);
nand UO_3346 (O_3346,N_47760,N_48641);
and UO_3347 (O_3347,N_48616,N_49554);
xnor UO_3348 (O_3348,N_48810,N_49143);
or UO_3349 (O_3349,N_49437,N_49838);
xor UO_3350 (O_3350,N_48630,N_49389);
and UO_3351 (O_3351,N_47630,N_48460);
xnor UO_3352 (O_3352,N_49739,N_48081);
nand UO_3353 (O_3353,N_48729,N_49437);
nand UO_3354 (O_3354,N_49647,N_49941);
xnor UO_3355 (O_3355,N_49366,N_49452);
nor UO_3356 (O_3356,N_48176,N_49540);
nor UO_3357 (O_3357,N_49884,N_49298);
and UO_3358 (O_3358,N_48079,N_48295);
nand UO_3359 (O_3359,N_48933,N_49356);
and UO_3360 (O_3360,N_49066,N_47647);
xnor UO_3361 (O_3361,N_48858,N_49419);
xor UO_3362 (O_3362,N_48636,N_48650);
nor UO_3363 (O_3363,N_48450,N_48184);
nor UO_3364 (O_3364,N_48824,N_47555);
or UO_3365 (O_3365,N_48750,N_49132);
nor UO_3366 (O_3366,N_48865,N_48551);
nand UO_3367 (O_3367,N_48761,N_48494);
xnor UO_3368 (O_3368,N_49450,N_48726);
or UO_3369 (O_3369,N_48344,N_48565);
nand UO_3370 (O_3370,N_49479,N_49991);
xnor UO_3371 (O_3371,N_48210,N_48733);
and UO_3372 (O_3372,N_49505,N_49399);
or UO_3373 (O_3373,N_49265,N_48888);
and UO_3374 (O_3374,N_47508,N_49221);
nand UO_3375 (O_3375,N_47742,N_48405);
nor UO_3376 (O_3376,N_48033,N_48208);
and UO_3377 (O_3377,N_48646,N_49275);
and UO_3378 (O_3378,N_48463,N_48538);
nor UO_3379 (O_3379,N_47614,N_47612);
xor UO_3380 (O_3380,N_48319,N_48474);
or UO_3381 (O_3381,N_48514,N_47824);
xnor UO_3382 (O_3382,N_48994,N_49604);
and UO_3383 (O_3383,N_49971,N_49114);
and UO_3384 (O_3384,N_49478,N_48821);
nor UO_3385 (O_3385,N_48801,N_48790);
and UO_3386 (O_3386,N_48324,N_49467);
and UO_3387 (O_3387,N_48749,N_49947);
xor UO_3388 (O_3388,N_49295,N_49727);
nand UO_3389 (O_3389,N_47782,N_47915);
nand UO_3390 (O_3390,N_48334,N_47952);
xnor UO_3391 (O_3391,N_47892,N_49788);
and UO_3392 (O_3392,N_49235,N_47977);
or UO_3393 (O_3393,N_48338,N_47867);
nand UO_3394 (O_3394,N_49117,N_48663);
nor UO_3395 (O_3395,N_49929,N_49622);
xnor UO_3396 (O_3396,N_49631,N_48596);
nor UO_3397 (O_3397,N_49645,N_47900);
and UO_3398 (O_3398,N_49417,N_48637);
or UO_3399 (O_3399,N_49714,N_49419);
and UO_3400 (O_3400,N_47792,N_49023);
nor UO_3401 (O_3401,N_49144,N_49428);
or UO_3402 (O_3402,N_49826,N_48731);
nor UO_3403 (O_3403,N_48041,N_49075);
and UO_3404 (O_3404,N_49514,N_49173);
and UO_3405 (O_3405,N_49469,N_49738);
nand UO_3406 (O_3406,N_49572,N_48909);
nand UO_3407 (O_3407,N_48284,N_48115);
nand UO_3408 (O_3408,N_49990,N_47765);
xor UO_3409 (O_3409,N_48267,N_49811);
and UO_3410 (O_3410,N_49304,N_48463);
or UO_3411 (O_3411,N_48546,N_49301);
or UO_3412 (O_3412,N_49942,N_49916);
and UO_3413 (O_3413,N_48827,N_47868);
nand UO_3414 (O_3414,N_49282,N_49280);
and UO_3415 (O_3415,N_49025,N_48916);
or UO_3416 (O_3416,N_48320,N_47676);
nand UO_3417 (O_3417,N_48838,N_48430);
and UO_3418 (O_3418,N_49541,N_49268);
and UO_3419 (O_3419,N_49546,N_48583);
nand UO_3420 (O_3420,N_47664,N_48310);
nand UO_3421 (O_3421,N_47850,N_48080);
xnor UO_3422 (O_3422,N_49348,N_49184);
nor UO_3423 (O_3423,N_48311,N_49293);
xor UO_3424 (O_3424,N_49497,N_49109);
or UO_3425 (O_3425,N_49064,N_47633);
nand UO_3426 (O_3426,N_48839,N_48879);
nor UO_3427 (O_3427,N_48759,N_47588);
and UO_3428 (O_3428,N_49845,N_48121);
and UO_3429 (O_3429,N_48382,N_47636);
xor UO_3430 (O_3430,N_47750,N_49468);
or UO_3431 (O_3431,N_49707,N_48836);
xor UO_3432 (O_3432,N_49353,N_48566);
or UO_3433 (O_3433,N_48699,N_48046);
or UO_3434 (O_3434,N_49245,N_48911);
xnor UO_3435 (O_3435,N_49808,N_49959);
or UO_3436 (O_3436,N_49453,N_48311);
nor UO_3437 (O_3437,N_49214,N_48276);
nand UO_3438 (O_3438,N_49446,N_49461);
nand UO_3439 (O_3439,N_47946,N_49747);
or UO_3440 (O_3440,N_49875,N_49672);
nor UO_3441 (O_3441,N_48361,N_48809);
xnor UO_3442 (O_3442,N_48273,N_48073);
nand UO_3443 (O_3443,N_48452,N_48878);
and UO_3444 (O_3444,N_49421,N_49590);
or UO_3445 (O_3445,N_48327,N_49382);
xor UO_3446 (O_3446,N_48645,N_49958);
or UO_3447 (O_3447,N_47711,N_48876);
nand UO_3448 (O_3448,N_48568,N_47645);
or UO_3449 (O_3449,N_49318,N_48899);
nor UO_3450 (O_3450,N_49046,N_49225);
nand UO_3451 (O_3451,N_48677,N_48595);
and UO_3452 (O_3452,N_49150,N_49910);
nor UO_3453 (O_3453,N_48846,N_49473);
nor UO_3454 (O_3454,N_48570,N_48289);
nand UO_3455 (O_3455,N_47717,N_47900);
nand UO_3456 (O_3456,N_49793,N_48540);
and UO_3457 (O_3457,N_49531,N_48346);
xor UO_3458 (O_3458,N_48875,N_49443);
nor UO_3459 (O_3459,N_49763,N_47854);
nand UO_3460 (O_3460,N_48215,N_48685);
xor UO_3461 (O_3461,N_47882,N_49805);
and UO_3462 (O_3462,N_48640,N_47743);
nand UO_3463 (O_3463,N_49112,N_49482);
nor UO_3464 (O_3464,N_47838,N_47577);
and UO_3465 (O_3465,N_49948,N_48045);
and UO_3466 (O_3466,N_47569,N_49091);
nand UO_3467 (O_3467,N_47627,N_47584);
nor UO_3468 (O_3468,N_49927,N_49821);
xor UO_3469 (O_3469,N_47590,N_49343);
nand UO_3470 (O_3470,N_49065,N_47601);
nand UO_3471 (O_3471,N_48080,N_48146);
and UO_3472 (O_3472,N_48886,N_47786);
nand UO_3473 (O_3473,N_49997,N_48103);
and UO_3474 (O_3474,N_49614,N_48860);
or UO_3475 (O_3475,N_48618,N_48478);
and UO_3476 (O_3476,N_48504,N_49492);
and UO_3477 (O_3477,N_47655,N_47667);
xnor UO_3478 (O_3478,N_49554,N_48800);
or UO_3479 (O_3479,N_47963,N_49602);
and UO_3480 (O_3480,N_48394,N_49153);
nor UO_3481 (O_3481,N_49599,N_48195);
xnor UO_3482 (O_3482,N_49014,N_47681);
or UO_3483 (O_3483,N_49901,N_48421);
xor UO_3484 (O_3484,N_48597,N_49650);
or UO_3485 (O_3485,N_48931,N_48892);
xnor UO_3486 (O_3486,N_49282,N_49297);
and UO_3487 (O_3487,N_49805,N_48009);
xnor UO_3488 (O_3488,N_48499,N_47944);
nor UO_3489 (O_3489,N_48619,N_48896);
nand UO_3490 (O_3490,N_48521,N_49604);
or UO_3491 (O_3491,N_47637,N_47557);
or UO_3492 (O_3492,N_48791,N_48772);
nand UO_3493 (O_3493,N_48226,N_49228);
or UO_3494 (O_3494,N_47888,N_49452);
or UO_3495 (O_3495,N_49670,N_47708);
or UO_3496 (O_3496,N_48005,N_48693);
or UO_3497 (O_3497,N_49131,N_49039);
nor UO_3498 (O_3498,N_49466,N_49385);
or UO_3499 (O_3499,N_48462,N_47929);
and UO_3500 (O_3500,N_48365,N_48690);
xor UO_3501 (O_3501,N_47626,N_49412);
or UO_3502 (O_3502,N_48865,N_48953);
nor UO_3503 (O_3503,N_47671,N_49232);
nand UO_3504 (O_3504,N_48584,N_47748);
nor UO_3505 (O_3505,N_49433,N_47742);
nor UO_3506 (O_3506,N_47946,N_49655);
xnor UO_3507 (O_3507,N_47705,N_47733);
and UO_3508 (O_3508,N_48422,N_49875);
nor UO_3509 (O_3509,N_49882,N_49119);
nand UO_3510 (O_3510,N_48252,N_48713);
xor UO_3511 (O_3511,N_48336,N_48478);
or UO_3512 (O_3512,N_47917,N_48595);
nor UO_3513 (O_3513,N_48979,N_49570);
nor UO_3514 (O_3514,N_48172,N_47962);
or UO_3515 (O_3515,N_48495,N_49420);
nor UO_3516 (O_3516,N_49371,N_48810);
xor UO_3517 (O_3517,N_49760,N_49156);
and UO_3518 (O_3518,N_49045,N_47855);
nand UO_3519 (O_3519,N_47523,N_49294);
xnor UO_3520 (O_3520,N_48249,N_49144);
nor UO_3521 (O_3521,N_49683,N_49701);
xnor UO_3522 (O_3522,N_47974,N_49089);
nand UO_3523 (O_3523,N_47674,N_48144);
nand UO_3524 (O_3524,N_48621,N_49407);
xnor UO_3525 (O_3525,N_49919,N_49251);
or UO_3526 (O_3526,N_47658,N_49400);
nand UO_3527 (O_3527,N_48110,N_48342);
and UO_3528 (O_3528,N_48635,N_49505);
or UO_3529 (O_3529,N_48598,N_47904);
nor UO_3530 (O_3530,N_48372,N_48899);
nand UO_3531 (O_3531,N_48769,N_49628);
or UO_3532 (O_3532,N_48891,N_49174);
nor UO_3533 (O_3533,N_48998,N_49068);
nand UO_3534 (O_3534,N_49888,N_48821);
and UO_3535 (O_3535,N_49211,N_48203);
or UO_3536 (O_3536,N_47813,N_48695);
nor UO_3537 (O_3537,N_49410,N_49273);
nor UO_3538 (O_3538,N_49232,N_47813);
nand UO_3539 (O_3539,N_47901,N_49468);
xor UO_3540 (O_3540,N_48481,N_48317);
and UO_3541 (O_3541,N_49377,N_49198);
nor UO_3542 (O_3542,N_49140,N_47849);
nor UO_3543 (O_3543,N_47718,N_48966);
nor UO_3544 (O_3544,N_49020,N_47794);
xor UO_3545 (O_3545,N_47721,N_47915);
xor UO_3546 (O_3546,N_49633,N_49715);
and UO_3547 (O_3547,N_48364,N_49341);
or UO_3548 (O_3548,N_49623,N_48135);
nor UO_3549 (O_3549,N_49211,N_47784);
or UO_3550 (O_3550,N_49457,N_48489);
xnor UO_3551 (O_3551,N_48447,N_49135);
and UO_3552 (O_3552,N_48950,N_49859);
nor UO_3553 (O_3553,N_48903,N_48601);
nor UO_3554 (O_3554,N_49220,N_49883);
nand UO_3555 (O_3555,N_47788,N_49442);
and UO_3556 (O_3556,N_48503,N_48033);
and UO_3557 (O_3557,N_48223,N_47679);
nand UO_3558 (O_3558,N_49128,N_49611);
nor UO_3559 (O_3559,N_49546,N_49173);
nand UO_3560 (O_3560,N_48619,N_49753);
or UO_3561 (O_3561,N_49012,N_48944);
nor UO_3562 (O_3562,N_49380,N_47814);
nand UO_3563 (O_3563,N_49348,N_47706);
or UO_3564 (O_3564,N_49046,N_49839);
nor UO_3565 (O_3565,N_48808,N_49429);
nand UO_3566 (O_3566,N_48433,N_49949);
nand UO_3567 (O_3567,N_48053,N_47870);
or UO_3568 (O_3568,N_48235,N_48888);
nand UO_3569 (O_3569,N_48479,N_48627);
nand UO_3570 (O_3570,N_47829,N_49221);
xor UO_3571 (O_3571,N_48039,N_48118);
nor UO_3572 (O_3572,N_49130,N_49319);
or UO_3573 (O_3573,N_49069,N_49477);
xor UO_3574 (O_3574,N_48212,N_47929);
nor UO_3575 (O_3575,N_48852,N_48042);
xnor UO_3576 (O_3576,N_49767,N_48142);
xnor UO_3577 (O_3577,N_49682,N_48372);
xor UO_3578 (O_3578,N_49301,N_47720);
and UO_3579 (O_3579,N_47713,N_48195);
xnor UO_3580 (O_3580,N_48692,N_47681);
xor UO_3581 (O_3581,N_49705,N_48638);
nor UO_3582 (O_3582,N_49347,N_47768);
and UO_3583 (O_3583,N_49445,N_49421);
nor UO_3584 (O_3584,N_49198,N_48996);
xnor UO_3585 (O_3585,N_47557,N_49219);
xor UO_3586 (O_3586,N_49189,N_48149);
nor UO_3587 (O_3587,N_49660,N_49176);
nand UO_3588 (O_3588,N_49882,N_47897);
nand UO_3589 (O_3589,N_48296,N_49886);
and UO_3590 (O_3590,N_48712,N_48432);
nor UO_3591 (O_3591,N_49224,N_49025);
and UO_3592 (O_3592,N_48159,N_48595);
xor UO_3593 (O_3593,N_47670,N_47850);
xnor UO_3594 (O_3594,N_48124,N_47873);
and UO_3595 (O_3595,N_49546,N_48177);
and UO_3596 (O_3596,N_47886,N_49036);
nand UO_3597 (O_3597,N_48230,N_47857);
nor UO_3598 (O_3598,N_47683,N_48549);
xor UO_3599 (O_3599,N_47785,N_48650);
xnor UO_3600 (O_3600,N_49805,N_49067);
or UO_3601 (O_3601,N_48702,N_48212);
nor UO_3602 (O_3602,N_48718,N_48879);
xor UO_3603 (O_3603,N_48402,N_49819);
nand UO_3604 (O_3604,N_48328,N_49074);
nand UO_3605 (O_3605,N_48870,N_48022);
or UO_3606 (O_3606,N_48878,N_48120);
and UO_3607 (O_3607,N_48054,N_47882);
xnor UO_3608 (O_3608,N_49216,N_49885);
xnor UO_3609 (O_3609,N_48514,N_49293);
or UO_3610 (O_3610,N_48791,N_47949);
and UO_3611 (O_3611,N_48838,N_49705);
and UO_3612 (O_3612,N_48379,N_49654);
nand UO_3613 (O_3613,N_48280,N_48122);
nor UO_3614 (O_3614,N_48374,N_48028);
and UO_3615 (O_3615,N_48545,N_47679);
nor UO_3616 (O_3616,N_49325,N_49148);
or UO_3617 (O_3617,N_49241,N_48414);
nand UO_3618 (O_3618,N_49004,N_49935);
nor UO_3619 (O_3619,N_49855,N_48387);
nand UO_3620 (O_3620,N_49686,N_48969);
and UO_3621 (O_3621,N_49906,N_49285);
xnor UO_3622 (O_3622,N_48530,N_48162);
nor UO_3623 (O_3623,N_48814,N_48551);
nand UO_3624 (O_3624,N_48927,N_49175);
or UO_3625 (O_3625,N_48485,N_48861);
nor UO_3626 (O_3626,N_47600,N_48192);
nor UO_3627 (O_3627,N_47870,N_48251);
nor UO_3628 (O_3628,N_48534,N_49542);
xnor UO_3629 (O_3629,N_48059,N_48054);
and UO_3630 (O_3630,N_48285,N_49454);
nand UO_3631 (O_3631,N_49762,N_48326);
and UO_3632 (O_3632,N_49454,N_49818);
or UO_3633 (O_3633,N_49040,N_49985);
nand UO_3634 (O_3634,N_49092,N_48038);
nor UO_3635 (O_3635,N_49429,N_49652);
or UO_3636 (O_3636,N_49321,N_49469);
nand UO_3637 (O_3637,N_49063,N_48272);
and UO_3638 (O_3638,N_47502,N_48499);
xnor UO_3639 (O_3639,N_48493,N_48512);
nor UO_3640 (O_3640,N_47955,N_48818);
xor UO_3641 (O_3641,N_49443,N_48326);
nor UO_3642 (O_3642,N_49194,N_48222);
and UO_3643 (O_3643,N_48330,N_49251);
nand UO_3644 (O_3644,N_48157,N_49362);
or UO_3645 (O_3645,N_49280,N_48671);
and UO_3646 (O_3646,N_48257,N_49405);
nand UO_3647 (O_3647,N_48044,N_48825);
and UO_3648 (O_3648,N_49094,N_48740);
and UO_3649 (O_3649,N_49462,N_49024);
nand UO_3650 (O_3650,N_48168,N_48086);
nand UO_3651 (O_3651,N_48259,N_49076);
xnor UO_3652 (O_3652,N_47632,N_48101);
and UO_3653 (O_3653,N_49326,N_49791);
or UO_3654 (O_3654,N_49231,N_49720);
and UO_3655 (O_3655,N_49456,N_48413);
nand UO_3656 (O_3656,N_48038,N_49491);
or UO_3657 (O_3657,N_48108,N_47775);
xnor UO_3658 (O_3658,N_49760,N_48164);
xor UO_3659 (O_3659,N_49024,N_47927);
xor UO_3660 (O_3660,N_49372,N_48823);
xor UO_3661 (O_3661,N_48477,N_48045);
or UO_3662 (O_3662,N_47967,N_48690);
and UO_3663 (O_3663,N_48432,N_49601);
nand UO_3664 (O_3664,N_48981,N_48164);
xor UO_3665 (O_3665,N_48239,N_49494);
xor UO_3666 (O_3666,N_48418,N_49334);
or UO_3667 (O_3667,N_48900,N_47984);
nor UO_3668 (O_3668,N_49029,N_48977);
and UO_3669 (O_3669,N_49179,N_48499);
nand UO_3670 (O_3670,N_49475,N_49216);
nand UO_3671 (O_3671,N_49925,N_48264);
xor UO_3672 (O_3672,N_48439,N_49191);
nor UO_3673 (O_3673,N_49507,N_49730);
and UO_3674 (O_3674,N_49760,N_48842);
xor UO_3675 (O_3675,N_48847,N_47708);
nor UO_3676 (O_3676,N_47859,N_49333);
and UO_3677 (O_3677,N_49104,N_49945);
or UO_3678 (O_3678,N_49876,N_48553);
nand UO_3679 (O_3679,N_47814,N_49797);
and UO_3680 (O_3680,N_47500,N_49946);
and UO_3681 (O_3681,N_48990,N_49203);
or UO_3682 (O_3682,N_47928,N_48208);
and UO_3683 (O_3683,N_48361,N_49567);
nand UO_3684 (O_3684,N_48810,N_47794);
or UO_3685 (O_3685,N_48326,N_48594);
nor UO_3686 (O_3686,N_48729,N_47871);
xnor UO_3687 (O_3687,N_47973,N_49571);
and UO_3688 (O_3688,N_48438,N_48288);
xor UO_3689 (O_3689,N_47775,N_49106);
and UO_3690 (O_3690,N_49093,N_49441);
nand UO_3691 (O_3691,N_47949,N_49295);
and UO_3692 (O_3692,N_49650,N_48806);
nand UO_3693 (O_3693,N_49618,N_49464);
xor UO_3694 (O_3694,N_48167,N_48369);
nor UO_3695 (O_3695,N_49231,N_49498);
and UO_3696 (O_3696,N_48411,N_47772);
nand UO_3697 (O_3697,N_48827,N_49906);
nor UO_3698 (O_3698,N_49299,N_47558);
or UO_3699 (O_3699,N_47810,N_48879);
or UO_3700 (O_3700,N_48173,N_47953);
and UO_3701 (O_3701,N_48209,N_49205);
and UO_3702 (O_3702,N_47571,N_47714);
or UO_3703 (O_3703,N_48491,N_49456);
xnor UO_3704 (O_3704,N_48402,N_48779);
nand UO_3705 (O_3705,N_49648,N_48926);
and UO_3706 (O_3706,N_49868,N_48376);
xnor UO_3707 (O_3707,N_49461,N_49495);
nand UO_3708 (O_3708,N_48127,N_47542);
nand UO_3709 (O_3709,N_48653,N_47556);
or UO_3710 (O_3710,N_49245,N_49849);
and UO_3711 (O_3711,N_48156,N_47753);
or UO_3712 (O_3712,N_49052,N_49711);
and UO_3713 (O_3713,N_47701,N_47654);
nor UO_3714 (O_3714,N_48187,N_47671);
nand UO_3715 (O_3715,N_48095,N_48415);
or UO_3716 (O_3716,N_48484,N_48340);
nor UO_3717 (O_3717,N_48518,N_49416);
or UO_3718 (O_3718,N_48987,N_48900);
nand UO_3719 (O_3719,N_49220,N_47908);
xor UO_3720 (O_3720,N_49342,N_49953);
or UO_3721 (O_3721,N_48186,N_49654);
and UO_3722 (O_3722,N_49302,N_48300);
or UO_3723 (O_3723,N_47530,N_49857);
or UO_3724 (O_3724,N_48976,N_47588);
nor UO_3725 (O_3725,N_49783,N_49297);
or UO_3726 (O_3726,N_49489,N_49602);
xnor UO_3727 (O_3727,N_47882,N_48155);
nor UO_3728 (O_3728,N_49376,N_48435);
or UO_3729 (O_3729,N_49227,N_49915);
nor UO_3730 (O_3730,N_47709,N_48133);
nand UO_3731 (O_3731,N_49682,N_48354);
nand UO_3732 (O_3732,N_48165,N_49430);
nand UO_3733 (O_3733,N_49263,N_47543);
and UO_3734 (O_3734,N_49606,N_47529);
xor UO_3735 (O_3735,N_48310,N_48190);
and UO_3736 (O_3736,N_49304,N_48550);
and UO_3737 (O_3737,N_47528,N_49575);
and UO_3738 (O_3738,N_47611,N_49768);
xnor UO_3739 (O_3739,N_48106,N_47735);
or UO_3740 (O_3740,N_48662,N_47770);
or UO_3741 (O_3741,N_48437,N_49470);
xor UO_3742 (O_3742,N_49547,N_49074);
and UO_3743 (O_3743,N_48592,N_48114);
nor UO_3744 (O_3744,N_47550,N_49747);
nand UO_3745 (O_3745,N_49684,N_48336);
nor UO_3746 (O_3746,N_47964,N_47667);
xor UO_3747 (O_3747,N_48510,N_47903);
xor UO_3748 (O_3748,N_49457,N_48493);
and UO_3749 (O_3749,N_49585,N_48207);
nor UO_3750 (O_3750,N_49850,N_47800);
or UO_3751 (O_3751,N_49405,N_49025);
or UO_3752 (O_3752,N_49766,N_49504);
and UO_3753 (O_3753,N_49359,N_48782);
nor UO_3754 (O_3754,N_47956,N_47655);
and UO_3755 (O_3755,N_48913,N_47537);
nand UO_3756 (O_3756,N_48886,N_49584);
and UO_3757 (O_3757,N_47664,N_49256);
xor UO_3758 (O_3758,N_48579,N_47789);
nor UO_3759 (O_3759,N_49370,N_48216);
or UO_3760 (O_3760,N_49580,N_49492);
xor UO_3761 (O_3761,N_49593,N_49340);
or UO_3762 (O_3762,N_49228,N_49830);
xnor UO_3763 (O_3763,N_49162,N_49477);
nor UO_3764 (O_3764,N_49742,N_48592);
or UO_3765 (O_3765,N_48148,N_48613);
nor UO_3766 (O_3766,N_48016,N_48014);
and UO_3767 (O_3767,N_49299,N_48664);
or UO_3768 (O_3768,N_47659,N_49841);
xnor UO_3769 (O_3769,N_47925,N_47740);
and UO_3770 (O_3770,N_49374,N_49558);
nor UO_3771 (O_3771,N_48737,N_49499);
nand UO_3772 (O_3772,N_49157,N_47841);
or UO_3773 (O_3773,N_47685,N_47582);
and UO_3774 (O_3774,N_48575,N_48759);
nand UO_3775 (O_3775,N_47894,N_48222);
xor UO_3776 (O_3776,N_49606,N_49817);
and UO_3777 (O_3777,N_49783,N_49149);
nand UO_3778 (O_3778,N_49194,N_48919);
xnor UO_3779 (O_3779,N_49692,N_47707);
xor UO_3780 (O_3780,N_47895,N_49330);
nand UO_3781 (O_3781,N_49634,N_49720);
xnor UO_3782 (O_3782,N_49475,N_49557);
nand UO_3783 (O_3783,N_48096,N_49240);
or UO_3784 (O_3784,N_48247,N_49686);
xnor UO_3785 (O_3785,N_49720,N_49228);
nor UO_3786 (O_3786,N_47593,N_49497);
xor UO_3787 (O_3787,N_48656,N_49847);
nand UO_3788 (O_3788,N_49649,N_49983);
and UO_3789 (O_3789,N_49261,N_49082);
or UO_3790 (O_3790,N_49972,N_49680);
nor UO_3791 (O_3791,N_48335,N_48801);
nand UO_3792 (O_3792,N_49086,N_49188);
or UO_3793 (O_3793,N_49540,N_49364);
nor UO_3794 (O_3794,N_49345,N_47573);
nand UO_3795 (O_3795,N_47880,N_47929);
and UO_3796 (O_3796,N_49586,N_48644);
xor UO_3797 (O_3797,N_49657,N_47660);
xnor UO_3798 (O_3798,N_49096,N_49658);
or UO_3799 (O_3799,N_49774,N_49359);
nand UO_3800 (O_3800,N_47762,N_48573);
or UO_3801 (O_3801,N_49062,N_49257);
nor UO_3802 (O_3802,N_48296,N_47726);
or UO_3803 (O_3803,N_49158,N_49171);
nor UO_3804 (O_3804,N_49757,N_49061);
nor UO_3805 (O_3805,N_49646,N_48174);
xor UO_3806 (O_3806,N_49166,N_49033);
or UO_3807 (O_3807,N_48517,N_49949);
nor UO_3808 (O_3808,N_47622,N_48196);
nand UO_3809 (O_3809,N_48783,N_49732);
nand UO_3810 (O_3810,N_48522,N_49320);
nand UO_3811 (O_3811,N_48486,N_48001);
nand UO_3812 (O_3812,N_49527,N_47607);
and UO_3813 (O_3813,N_48258,N_49974);
xnor UO_3814 (O_3814,N_49553,N_49656);
nand UO_3815 (O_3815,N_48921,N_47627);
or UO_3816 (O_3816,N_49375,N_48438);
or UO_3817 (O_3817,N_47823,N_49988);
and UO_3818 (O_3818,N_48595,N_48394);
nor UO_3819 (O_3819,N_48586,N_47818);
or UO_3820 (O_3820,N_47944,N_49060);
or UO_3821 (O_3821,N_49358,N_47924);
and UO_3822 (O_3822,N_48243,N_48087);
nand UO_3823 (O_3823,N_48167,N_49676);
xnor UO_3824 (O_3824,N_49332,N_48510);
nand UO_3825 (O_3825,N_48643,N_49714);
nor UO_3826 (O_3826,N_49247,N_48568);
nor UO_3827 (O_3827,N_49531,N_49844);
nor UO_3828 (O_3828,N_49293,N_48464);
nor UO_3829 (O_3829,N_48953,N_49207);
or UO_3830 (O_3830,N_48867,N_49101);
and UO_3831 (O_3831,N_48466,N_49744);
and UO_3832 (O_3832,N_47646,N_49338);
and UO_3833 (O_3833,N_48817,N_48693);
or UO_3834 (O_3834,N_49212,N_49236);
or UO_3835 (O_3835,N_49301,N_48938);
nor UO_3836 (O_3836,N_48630,N_49912);
or UO_3837 (O_3837,N_49461,N_49909);
or UO_3838 (O_3838,N_48307,N_48410);
nand UO_3839 (O_3839,N_47946,N_48433);
nand UO_3840 (O_3840,N_47928,N_47826);
and UO_3841 (O_3841,N_49640,N_48188);
and UO_3842 (O_3842,N_49885,N_49034);
xor UO_3843 (O_3843,N_48519,N_49043);
or UO_3844 (O_3844,N_48435,N_49948);
and UO_3845 (O_3845,N_48483,N_48112);
nand UO_3846 (O_3846,N_49276,N_49414);
nor UO_3847 (O_3847,N_49682,N_48883);
xor UO_3848 (O_3848,N_48208,N_49757);
nand UO_3849 (O_3849,N_47768,N_47536);
and UO_3850 (O_3850,N_49750,N_48999);
nor UO_3851 (O_3851,N_49354,N_48344);
xor UO_3852 (O_3852,N_49052,N_48549);
nand UO_3853 (O_3853,N_48650,N_48810);
or UO_3854 (O_3854,N_48237,N_48434);
nor UO_3855 (O_3855,N_47964,N_49010);
and UO_3856 (O_3856,N_49163,N_48363);
and UO_3857 (O_3857,N_49074,N_49611);
and UO_3858 (O_3858,N_48417,N_49399);
or UO_3859 (O_3859,N_47643,N_48427);
nand UO_3860 (O_3860,N_47866,N_48384);
nor UO_3861 (O_3861,N_48361,N_48006);
or UO_3862 (O_3862,N_49203,N_49632);
xnor UO_3863 (O_3863,N_49913,N_48313);
or UO_3864 (O_3864,N_47961,N_47938);
xnor UO_3865 (O_3865,N_49069,N_49430);
xor UO_3866 (O_3866,N_47539,N_49047);
xor UO_3867 (O_3867,N_48247,N_47829);
nand UO_3868 (O_3868,N_48001,N_47767);
and UO_3869 (O_3869,N_49000,N_48395);
xor UO_3870 (O_3870,N_47753,N_49172);
nand UO_3871 (O_3871,N_49330,N_47988);
and UO_3872 (O_3872,N_49307,N_48111);
nor UO_3873 (O_3873,N_49845,N_49499);
xnor UO_3874 (O_3874,N_48269,N_47821);
or UO_3875 (O_3875,N_49464,N_47923);
xor UO_3876 (O_3876,N_47754,N_48394);
xnor UO_3877 (O_3877,N_48589,N_48377);
xnor UO_3878 (O_3878,N_48238,N_49550);
and UO_3879 (O_3879,N_47554,N_49885);
nand UO_3880 (O_3880,N_48782,N_48148);
nand UO_3881 (O_3881,N_48229,N_48687);
or UO_3882 (O_3882,N_48345,N_49604);
nor UO_3883 (O_3883,N_48825,N_49083);
or UO_3884 (O_3884,N_48864,N_47760);
xor UO_3885 (O_3885,N_49186,N_49326);
nor UO_3886 (O_3886,N_48429,N_48413);
nand UO_3887 (O_3887,N_47590,N_49326);
nand UO_3888 (O_3888,N_47615,N_47757);
and UO_3889 (O_3889,N_49774,N_49233);
or UO_3890 (O_3890,N_48344,N_47575);
nor UO_3891 (O_3891,N_49722,N_48822);
or UO_3892 (O_3892,N_48004,N_48106);
nand UO_3893 (O_3893,N_48746,N_48235);
nand UO_3894 (O_3894,N_49374,N_49960);
xor UO_3895 (O_3895,N_48664,N_48315);
nor UO_3896 (O_3896,N_48140,N_48385);
nand UO_3897 (O_3897,N_49828,N_47963);
nor UO_3898 (O_3898,N_49368,N_48395);
and UO_3899 (O_3899,N_47635,N_49473);
nand UO_3900 (O_3900,N_47542,N_48421);
and UO_3901 (O_3901,N_48819,N_49176);
and UO_3902 (O_3902,N_47565,N_49048);
nand UO_3903 (O_3903,N_49985,N_49569);
xor UO_3904 (O_3904,N_49197,N_47667);
and UO_3905 (O_3905,N_49262,N_49583);
or UO_3906 (O_3906,N_49744,N_49517);
nor UO_3907 (O_3907,N_48579,N_49167);
nor UO_3908 (O_3908,N_48110,N_49756);
and UO_3909 (O_3909,N_48078,N_48699);
nor UO_3910 (O_3910,N_48061,N_48187);
nand UO_3911 (O_3911,N_48407,N_48533);
nor UO_3912 (O_3912,N_49125,N_49854);
xor UO_3913 (O_3913,N_49174,N_49517);
and UO_3914 (O_3914,N_48263,N_48209);
xnor UO_3915 (O_3915,N_48956,N_48210);
nor UO_3916 (O_3916,N_48134,N_48556);
and UO_3917 (O_3917,N_48755,N_49770);
xor UO_3918 (O_3918,N_49677,N_49791);
or UO_3919 (O_3919,N_49784,N_49381);
xnor UO_3920 (O_3920,N_49724,N_49545);
and UO_3921 (O_3921,N_49714,N_49537);
or UO_3922 (O_3922,N_47983,N_49290);
or UO_3923 (O_3923,N_47928,N_49530);
nor UO_3924 (O_3924,N_49904,N_49713);
nand UO_3925 (O_3925,N_48980,N_49683);
or UO_3926 (O_3926,N_48808,N_49419);
xnor UO_3927 (O_3927,N_48138,N_49240);
nor UO_3928 (O_3928,N_48868,N_48186);
nand UO_3929 (O_3929,N_48362,N_49389);
and UO_3930 (O_3930,N_48937,N_48739);
and UO_3931 (O_3931,N_48292,N_48452);
nor UO_3932 (O_3932,N_48640,N_48053);
nand UO_3933 (O_3933,N_48130,N_47814);
nor UO_3934 (O_3934,N_49201,N_49362);
nand UO_3935 (O_3935,N_48922,N_47521);
or UO_3936 (O_3936,N_49844,N_49536);
nand UO_3937 (O_3937,N_47935,N_48848);
and UO_3938 (O_3938,N_48233,N_49042);
nor UO_3939 (O_3939,N_49160,N_48762);
or UO_3940 (O_3940,N_49082,N_47623);
or UO_3941 (O_3941,N_48775,N_49982);
xnor UO_3942 (O_3942,N_48891,N_49608);
xor UO_3943 (O_3943,N_49785,N_49192);
or UO_3944 (O_3944,N_49594,N_49234);
xnor UO_3945 (O_3945,N_47959,N_47774);
nand UO_3946 (O_3946,N_49564,N_49309);
xnor UO_3947 (O_3947,N_49837,N_49008);
or UO_3948 (O_3948,N_49363,N_47903);
nand UO_3949 (O_3949,N_48491,N_49602);
nor UO_3950 (O_3950,N_49259,N_49474);
xor UO_3951 (O_3951,N_48470,N_48920);
xnor UO_3952 (O_3952,N_48141,N_47701);
nand UO_3953 (O_3953,N_49030,N_49290);
or UO_3954 (O_3954,N_47806,N_48498);
nor UO_3955 (O_3955,N_47563,N_49836);
or UO_3956 (O_3956,N_47623,N_48546);
xnor UO_3957 (O_3957,N_49955,N_48393);
nor UO_3958 (O_3958,N_48245,N_47554);
nor UO_3959 (O_3959,N_47840,N_49479);
xnor UO_3960 (O_3960,N_49704,N_48046);
xor UO_3961 (O_3961,N_49508,N_48635);
nor UO_3962 (O_3962,N_47605,N_47720);
xor UO_3963 (O_3963,N_47556,N_48940);
xnor UO_3964 (O_3964,N_47670,N_48088);
xor UO_3965 (O_3965,N_48947,N_47696);
and UO_3966 (O_3966,N_48883,N_49904);
nor UO_3967 (O_3967,N_48909,N_48687);
and UO_3968 (O_3968,N_47600,N_47969);
xor UO_3969 (O_3969,N_48294,N_49464);
xnor UO_3970 (O_3970,N_49365,N_49081);
nor UO_3971 (O_3971,N_48879,N_49803);
or UO_3972 (O_3972,N_48287,N_49648);
and UO_3973 (O_3973,N_48921,N_49401);
or UO_3974 (O_3974,N_49544,N_48650);
and UO_3975 (O_3975,N_47688,N_48911);
and UO_3976 (O_3976,N_48744,N_48927);
and UO_3977 (O_3977,N_47669,N_48660);
xnor UO_3978 (O_3978,N_49730,N_49796);
xnor UO_3979 (O_3979,N_49425,N_48959);
xor UO_3980 (O_3980,N_49333,N_48082);
xnor UO_3981 (O_3981,N_49760,N_49601);
nand UO_3982 (O_3982,N_47976,N_47715);
xnor UO_3983 (O_3983,N_49825,N_48022);
nor UO_3984 (O_3984,N_48269,N_48150);
xnor UO_3985 (O_3985,N_48948,N_48486);
xor UO_3986 (O_3986,N_49513,N_48529);
or UO_3987 (O_3987,N_47844,N_49201);
xnor UO_3988 (O_3988,N_49400,N_49304);
and UO_3989 (O_3989,N_48153,N_48464);
nand UO_3990 (O_3990,N_48753,N_48343);
xnor UO_3991 (O_3991,N_47531,N_48276);
nor UO_3992 (O_3992,N_48495,N_47690);
nor UO_3993 (O_3993,N_48615,N_48062);
nand UO_3994 (O_3994,N_48603,N_47775);
and UO_3995 (O_3995,N_49402,N_49587);
nor UO_3996 (O_3996,N_49905,N_48394);
nand UO_3997 (O_3997,N_47723,N_47501);
nand UO_3998 (O_3998,N_47950,N_47595);
nand UO_3999 (O_3999,N_47621,N_49045);
xor UO_4000 (O_4000,N_47549,N_49347);
and UO_4001 (O_4001,N_49596,N_49992);
nand UO_4002 (O_4002,N_49636,N_47523);
nand UO_4003 (O_4003,N_49533,N_48512);
and UO_4004 (O_4004,N_47879,N_48742);
or UO_4005 (O_4005,N_49995,N_48895);
xnor UO_4006 (O_4006,N_49597,N_48458);
and UO_4007 (O_4007,N_48930,N_48837);
and UO_4008 (O_4008,N_48734,N_49031);
and UO_4009 (O_4009,N_48969,N_49753);
nor UO_4010 (O_4010,N_49315,N_49725);
nand UO_4011 (O_4011,N_49104,N_48807);
xnor UO_4012 (O_4012,N_49588,N_49881);
xnor UO_4013 (O_4013,N_47556,N_49486);
xnor UO_4014 (O_4014,N_48187,N_48710);
nor UO_4015 (O_4015,N_49480,N_49995);
and UO_4016 (O_4016,N_48226,N_48990);
nor UO_4017 (O_4017,N_47884,N_49274);
nand UO_4018 (O_4018,N_48476,N_48363);
or UO_4019 (O_4019,N_49321,N_47779);
and UO_4020 (O_4020,N_49462,N_49440);
or UO_4021 (O_4021,N_49228,N_48830);
or UO_4022 (O_4022,N_49483,N_47701);
nand UO_4023 (O_4023,N_48973,N_48127);
nor UO_4024 (O_4024,N_49298,N_47571);
xor UO_4025 (O_4025,N_48093,N_47871);
or UO_4026 (O_4026,N_48152,N_49809);
and UO_4027 (O_4027,N_48475,N_49245);
nand UO_4028 (O_4028,N_48549,N_48001);
xor UO_4029 (O_4029,N_47892,N_47634);
or UO_4030 (O_4030,N_48174,N_47627);
and UO_4031 (O_4031,N_49512,N_48000);
nand UO_4032 (O_4032,N_48732,N_47623);
or UO_4033 (O_4033,N_49666,N_48609);
nand UO_4034 (O_4034,N_48856,N_49610);
xnor UO_4035 (O_4035,N_49164,N_48490);
and UO_4036 (O_4036,N_48309,N_47906);
nand UO_4037 (O_4037,N_49706,N_49236);
or UO_4038 (O_4038,N_48848,N_47557);
or UO_4039 (O_4039,N_47896,N_49477);
nand UO_4040 (O_4040,N_49440,N_47907);
nand UO_4041 (O_4041,N_47562,N_49495);
or UO_4042 (O_4042,N_49288,N_49701);
nand UO_4043 (O_4043,N_49166,N_49290);
and UO_4044 (O_4044,N_47816,N_47630);
nand UO_4045 (O_4045,N_47816,N_49040);
nand UO_4046 (O_4046,N_48804,N_47617);
and UO_4047 (O_4047,N_49068,N_49897);
and UO_4048 (O_4048,N_48593,N_48507);
or UO_4049 (O_4049,N_47529,N_48100);
and UO_4050 (O_4050,N_47643,N_49004);
nor UO_4051 (O_4051,N_49728,N_48142);
and UO_4052 (O_4052,N_48468,N_48149);
nor UO_4053 (O_4053,N_49410,N_48021);
and UO_4054 (O_4054,N_47832,N_49104);
nor UO_4055 (O_4055,N_48896,N_49443);
nand UO_4056 (O_4056,N_48509,N_49029);
nand UO_4057 (O_4057,N_48817,N_47651);
xor UO_4058 (O_4058,N_48351,N_49742);
nor UO_4059 (O_4059,N_49008,N_49160);
or UO_4060 (O_4060,N_48114,N_49273);
or UO_4061 (O_4061,N_49937,N_48063);
xor UO_4062 (O_4062,N_49713,N_47636);
nand UO_4063 (O_4063,N_49145,N_47817);
nand UO_4064 (O_4064,N_49141,N_49811);
nor UO_4065 (O_4065,N_48568,N_49489);
or UO_4066 (O_4066,N_48617,N_48289);
and UO_4067 (O_4067,N_47715,N_48049);
xor UO_4068 (O_4068,N_49862,N_48993);
xor UO_4069 (O_4069,N_49033,N_48814);
nor UO_4070 (O_4070,N_49978,N_48343);
or UO_4071 (O_4071,N_49477,N_49036);
nor UO_4072 (O_4072,N_47688,N_49934);
xnor UO_4073 (O_4073,N_49229,N_49897);
or UO_4074 (O_4074,N_49427,N_49845);
or UO_4075 (O_4075,N_47910,N_47679);
xnor UO_4076 (O_4076,N_47620,N_48439);
or UO_4077 (O_4077,N_47820,N_47704);
xnor UO_4078 (O_4078,N_47563,N_49491);
nor UO_4079 (O_4079,N_49754,N_48962);
and UO_4080 (O_4080,N_49667,N_48535);
nand UO_4081 (O_4081,N_48496,N_49136);
xnor UO_4082 (O_4082,N_49649,N_47804);
xnor UO_4083 (O_4083,N_48139,N_48626);
xnor UO_4084 (O_4084,N_48119,N_48797);
and UO_4085 (O_4085,N_49840,N_49149);
nand UO_4086 (O_4086,N_48438,N_49268);
nand UO_4087 (O_4087,N_49292,N_48631);
and UO_4088 (O_4088,N_48972,N_49737);
nand UO_4089 (O_4089,N_48664,N_47689);
xnor UO_4090 (O_4090,N_49970,N_49211);
nor UO_4091 (O_4091,N_49233,N_48928);
nor UO_4092 (O_4092,N_47736,N_49758);
and UO_4093 (O_4093,N_47509,N_49534);
and UO_4094 (O_4094,N_47590,N_49966);
and UO_4095 (O_4095,N_48788,N_48448);
xnor UO_4096 (O_4096,N_48176,N_48520);
nand UO_4097 (O_4097,N_49351,N_47688);
or UO_4098 (O_4098,N_47570,N_48743);
xor UO_4099 (O_4099,N_48227,N_48301);
nand UO_4100 (O_4100,N_49022,N_49862);
or UO_4101 (O_4101,N_49850,N_49918);
xor UO_4102 (O_4102,N_49317,N_47978);
xor UO_4103 (O_4103,N_49745,N_48213);
xor UO_4104 (O_4104,N_49312,N_49443);
nor UO_4105 (O_4105,N_49515,N_47894);
xnor UO_4106 (O_4106,N_48478,N_48151);
nand UO_4107 (O_4107,N_48454,N_47562);
or UO_4108 (O_4108,N_48809,N_48295);
or UO_4109 (O_4109,N_48438,N_47865);
nor UO_4110 (O_4110,N_48474,N_49309);
and UO_4111 (O_4111,N_49637,N_48926);
xnor UO_4112 (O_4112,N_49424,N_49400);
xor UO_4113 (O_4113,N_48236,N_49917);
nor UO_4114 (O_4114,N_49267,N_47840);
and UO_4115 (O_4115,N_48787,N_48805);
and UO_4116 (O_4116,N_48526,N_49871);
nor UO_4117 (O_4117,N_48860,N_49674);
nor UO_4118 (O_4118,N_49812,N_48416);
nand UO_4119 (O_4119,N_47970,N_47980);
or UO_4120 (O_4120,N_49558,N_49081);
nor UO_4121 (O_4121,N_49042,N_48744);
nand UO_4122 (O_4122,N_49290,N_47731);
nor UO_4123 (O_4123,N_49362,N_48256);
nand UO_4124 (O_4124,N_48840,N_49347);
or UO_4125 (O_4125,N_49175,N_48717);
xor UO_4126 (O_4126,N_48731,N_48158);
xor UO_4127 (O_4127,N_48901,N_48445);
xnor UO_4128 (O_4128,N_49693,N_49961);
xor UO_4129 (O_4129,N_49837,N_49812);
xor UO_4130 (O_4130,N_48299,N_49543);
nor UO_4131 (O_4131,N_48965,N_49687);
nand UO_4132 (O_4132,N_48458,N_48649);
xor UO_4133 (O_4133,N_48564,N_49750);
or UO_4134 (O_4134,N_49123,N_49455);
nand UO_4135 (O_4135,N_47672,N_48715);
nor UO_4136 (O_4136,N_48523,N_48618);
nand UO_4137 (O_4137,N_49767,N_47588);
xnor UO_4138 (O_4138,N_49905,N_49700);
or UO_4139 (O_4139,N_47856,N_48593);
nand UO_4140 (O_4140,N_48725,N_49808);
or UO_4141 (O_4141,N_49370,N_49888);
and UO_4142 (O_4142,N_48067,N_49318);
xor UO_4143 (O_4143,N_49716,N_47583);
xnor UO_4144 (O_4144,N_48424,N_47715);
nor UO_4145 (O_4145,N_49286,N_47550);
or UO_4146 (O_4146,N_49577,N_47702);
nor UO_4147 (O_4147,N_48709,N_47868);
and UO_4148 (O_4148,N_48117,N_47971);
nor UO_4149 (O_4149,N_47643,N_47716);
and UO_4150 (O_4150,N_49882,N_47858);
nor UO_4151 (O_4151,N_49138,N_49976);
nand UO_4152 (O_4152,N_47725,N_49242);
xor UO_4153 (O_4153,N_48322,N_49463);
nand UO_4154 (O_4154,N_48690,N_49077);
xor UO_4155 (O_4155,N_47652,N_49659);
or UO_4156 (O_4156,N_49366,N_49350);
and UO_4157 (O_4157,N_49975,N_49232);
and UO_4158 (O_4158,N_48848,N_48663);
or UO_4159 (O_4159,N_48535,N_49863);
nand UO_4160 (O_4160,N_49952,N_49346);
nand UO_4161 (O_4161,N_47613,N_47538);
and UO_4162 (O_4162,N_49990,N_48531);
xor UO_4163 (O_4163,N_47898,N_49877);
and UO_4164 (O_4164,N_49331,N_48186);
and UO_4165 (O_4165,N_48706,N_49414);
or UO_4166 (O_4166,N_48993,N_47629);
nor UO_4167 (O_4167,N_49206,N_48553);
nand UO_4168 (O_4168,N_48204,N_48051);
nand UO_4169 (O_4169,N_49584,N_48000);
nor UO_4170 (O_4170,N_49345,N_49240);
nand UO_4171 (O_4171,N_49818,N_47957);
xor UO_4172 (O_4172,N_48475,N_48858);
nand UO_4173 (O_4173,N_47581,N_49845);
and UO_4174 (O_4174,N_48305,N_48529);
or UO_4175 (O_4175,N_48875,N_49621);
or UO_4176 (O_4176,N_49836,N_49759);
xnor UO_4177 (O_4177,N_47968,N_49077);
or UO_4178 (O_4178,N_47827,N_47862);
or UO_4179 (O_4179,N_48824,N_48567);
nand UO_4180 (O_4180,N_49481,N_49470);
xnor UO_4181 (O_4181,N_47943,N_48740);
or UO_4182 (O_4182,N_48154,N_49192);
nor UO_4183 (O_4183,N_47677,N_49731);
nor UO_4184 (O_4184,N_48869,N_48598);
xnor UO_4185 (O_4185,N_49817,N_48626);
nor UO_4186 (O_4186,N_48505,N_49328);
and UO_4187 (O_4187,N_48862,N_48055);
or UO_4188 (O_4188,N_49009,N_49666);
nor UO_4189 (O_4189,N_49347,N_49797);
xor UO_4190 (O_4190,N_49673,N_49255);
or UO_4191 (O_4191,N_49984,N_49285);
nor UO_4192 (O_4192,N_49061,N_48223);
and UO_4193 (O_4193,N_47738,N_47832);
nand UO_4194 (O_4194,N_49307,N_49732);
nand UO_4195 (O_4195,N_49301,N_49698);
nand UO_4196 (O_4196,N_47539,N_49402);
or UO_4197 (O_4197,N_48655,N_47830);
nand UO_4198 (O_4198,N_48361,N_49919);
or UO_4199 (O_4199,N_47892,N_48467);
xor UO_4200 (O_4200,N_47564,N_49050);
or UO_4201 (O_4201,N_49193,N_48994);
and UO_4202 (O_4202,N_49150,N_47611);
xor UO_4203 (O_4203,N_49750,N_48304);
xor UO_4204 (O_4204,N_49683,N_47667);
nand UO_4205 (O_4205,N_47966,N_48457);
nor UO_4206 (O_4206,N_49321,N_47784);
xor UO_4207 (O_4207,N_49621,N_47843);
nand UO_4208 (O_4208,N_48974,N_49649);
or UO_4209 (O_4209,N_49097,N_48938);
and UO_4210 (O_4210,N_48114,N_48269);
and UO_4211 (O_4211,N_49165,N_49149);
or UO_4212 (O_4212,N_49134,N_47776);
or UO_4213 (O_4213,N_48953,N_49597);
nor UO_4214 (O_4214,N_49199,N_49990);
xor UO_4215 (O_4215,N_48213,N_49877);
nor UO_4216 (O_4216,N_48782,N_49831);
nor UO_4217 (O_4217,N_49885,N_49929);
nor UO_4218 (O_4218,N_47640,N_48078);
nor UO_4219 (O_4219,N_47985,N_47777);
and UO_4220 (O_4220,N_49818,N_49544);
xor UO_4221 (O_4221,N_48279,N_48306);
xnor UO_4222 (O_4222,N_48265,N_49011);
or UO_4223 (O_4223,N_47692,N_49169);
nand UO_4224 (O_4224,N_48587,N_48297);
nor UO_4225 (O_4225,N_48037,N_48456);
and UO_4226 (O_4226,N_49253,N_49912);
or UO_4227 (O_4227,N_48792,N_47743);
nor UO_4228 (O_4228,N_49333,N_48287);
xor UO_4229 (O_4229,N_48321,N_49587);
or UO_4230 (O_4230,N_49076,N_49656);
nor UO_4231 (O_4231,N_47628,N_49107);
nand UO_4232 (O_4232,N_49727,N_49067);
and UO_4233 (O_4233,N_48330,N_47708);
and UO_4234 (O_4234,N_47744,N_48893);
nand UO_4235 (O_4235,N_47677,N_47936);
nand UO_4236 (O_4236,N_48148,N_47512);
and UO_4237 (O_4237,N_47972,N_49182);
and UO_4238 (O_4238,N_48421,N_47973);
nor UO_4239 (O_4239,N_47530,N_48821);
xnor UO_4240 (O_4240,N_47933,N_48339);
nor UO_4241 (O_4241,N_47576,N_47746);
nor UO_4242 (O_4242,N_48206,N_48004);
nor UO_4243 (O_4243,N_49212,N_47521);
or UO_4244 (O_4244,N_47687,N_48440);
nor UO_4245 (O_4245,N_47837,N_47514);
or UO_4246 (O_4246,N_48077,N_48560);
nor UO_4247 (O_4247,N_48420,N_48244);
nand UO_4248 (O_4248,N_48677,N_49123);
nand UO_4249 (O_4249,N_49298,N_49817);
or UO_4250 (O_4250,N_48180,N_48491);
xor UO_4251 (O_4251,N_48544,N_48029);
or UO_4252 (O_4252,N_48360,N_47841);
nand UO_4253 (O_4253,N_48427,N_49017);
nor UO_4254 (O_4254,N_48425,N_47638);
nor UO_4255 (O_4255,N_48402,N_49918);
nand UO_4256 (O_4256,N_49073,N_49020);
xor UO_4257 (O_4257,N_49270,N_49272);
xnor UO_4258 (O_4258,N_48575,N_49789);
xor UO_4259 (O_4259,N_49033,N_47548);
or UO_4260 (O_4260,N_49948,N_49144);
or UO_4261 (O_4261,N_47648,N_47560);
nand UO_4262 (O_4262,N_49727,N_48753);
or UO_4263 (O_4263,N_49236,N_48022);
nor UO_4264 (O_4264,N_47589,N_49646);
nor UO_4265 (O_4265,N_49322,N_49584);
or UO_4266 (O_4266,N_49804,N_49231);
nor UO_4267 (O_4267,N_48563,N_49074);
and UO_4268 (O_4268,N_48999,N_48539);
nand UO_4269 (O_4269,N_49263,N_49785);
nor UO_4270 (O_4270,N_49763,N_48407);
nand UO_4271 (O_4271,N_49576,N_49154);
nor UO_4272 (O_4272,N_49214,N_47548);
nand UO_4273 (O_4273,N_49597,N_47597);
nand UO_4274 (O_4274,N_49610,N_49396);
and UO_4275 (O_4275,N_48356,N_49320);
and UO_4276 (O_4276,N_48934,N_49412);
xnor UO_4277 (O_4277,N_48494,N_48283);
nor UO_4278 (O_4278,N_49641,N_48905);
xor UO_4279 (O_4279,N_49403,N_49023);
nand UO_4280 (O_4280,N_47930,N_49388);
or UO_4281 (O_4281,N_48206,N_48300);
xor UO_4282 (O_4282,N_49775,N_49972);
nand UO_4283 (O_4283,N_47631,N_49883);
or UO_4284 (O_4284,N_48947,N_49242);
nor UO_4285 (O_4285,N_48893,N_49265);
or UO_4286 (O_4286,N_48797,N_48882);
xnor UO_4287 (O_4287,N_47978,N_49610);
xor UO_4288 (O_4288,N_47756,N_49138);
nand UO_4289 (O_4289,N_47957,N_47719);
nand UO_4290 (O_4290,N_48296,N_49522);
xnor UO_4291 (O_4291,N_48334,N_49021);
nor UO_4292 (O_4292,N_48464,N_49361);
and UO_4293 (O_4293,N_49042,N_47764);
xnor UO_4294 (O_4294,N_49150,N_49277);
and UO_4295 (O_4295,N_47734,N_47817);
xor UO_4296 (O_4296,N_47886,N_48842);
nor UO_4297 (O_4297,N_47742,N_49950);
xor UO_4298 (O_4298,N_49224,N_49288);
and UO_4299 (O_4299,N_48549,N_49014);
xor UO_4300 (O_4300,N_48340,N_48681);
nor UO_4301 (O_4301,N_47808,N_48312);
xnor UO_4302 (O_4302,N_48522,N_47668);
nor UO_4303 (O_4303,N_48438,N_47671);
and UO_4304 (O_4304,N_48352,N_48334);
or UO_4305 (O_4305,N_49498,N_48350);
or UO_4306 (O_4306,N_48619,N_48573);
nand UO_4307 (O_4307,N_49714,N_48080);
nor UO_4308 (O_4308,N_47682,N_49847);
nor UO_4309 (O_4309,N_49311,N_47927);
nand UO_4310 (O_4310,N_48812,N_47645);
nand UO_4311 (O_4311,N_49510,N_47605);
xor UO_4312 (O_4312,N_47581,N_48094);
and UO_4313 (O_4313,N_49612,N_48780);
or UO_4314 (O_4314,N_48499,N_49492);
or UO_4315 (O_4315,N_48257,N_48647);
xor UO_4316 (O_4316,N_49561,N_47722);
nand UO_4317 (O_4317,N_49358,N_49924);
nand UO_4318 (O_4318,N_49177,N_48953);
nand UO_4319 (O_4319,N_49764,N_48128);
or UO_4320 (O_4320,N_49606,N_49561);
or UO_4321 (O_4321,N_48659,N_49205);
nand UO_4322 (O_4322,N_48328,N_48079);
xnor UO_4323 (O_4323,N_48268,N_48343);
nand UO_4324 (O_4324,N_48516,N_49881);
nand UO_4325 (O_4325,N_48467,N_47820);
and UO_4326 (O_4326,N_47768,N_48719);
xnor UO_4327 (O_4327,N_47532,N_49732);
and UO_4328 (O_4328,N_48567,N_48866);
nand UO_4329 (O_4329,N_49384,N_47671);
or UO_4330 (O_4330,N_48988,N_48648);
nand UO_4331 (O_4331,N_49911,N_49059);
xnor UO_4332 (O_4332,N_49627,N_49796);
and UO_4333 (O_4333,N_48214,N_49378);
xor UO_4334 (O_4334,N_48224,N_48279);
or UO_4335 (O_4335,N_48800,N_49130);
nand UO_4336 (O_4336,N_48003,N_48340);
nand UO_4337 (O_4337,N_48527,N_48422);
nand UO_4338 (O_4338,N_48316,N_47551);
and UO_4339 (O_4339,N_48493,N_49380);
or UO_4340 (O_4340,N_48711,N_48110);
or UO_4341 (O_4341,N_47878,N_49181);
and UO_4342 (O_4342,N_49012,N_47649);
xor UO_4343 (O_4343,N_49626,N_47514);
nand UO_4344 (O_4344,N_49361,N_48218);
nor UO_4345 (O_4345,N_47825,N_48387);
or UO_4346 (O_4346,N_47600,N_48905);
nor UO_4347 (O_4347,N_47785,N_49391);
nor UO_4348 (O_4348,N_47644,N_49768);
nor UO_4349 (O_4349,N_47686,N_48845);
nor UO_4350 (O_4350,N_49135,N_48869);
nor UO_4351 (O_4351,N_48360,N_49241);
and UO_4352 (O_4352,N_48760,N_47670);
nand UO_4353 (O_4353,N_48108,N_49712);
and UO_4354 (O_4354,N_48781,N_48711);
xor UO_4355 (O_4355,N_49381,N_47958);
or UO_4356 (O_4356,N_49737,N_49566);
or UO_4357 (O_4357,N_47961,N_49530);
xnor UO_4358 (O_4358,N_47811,N_49317);
and UO_4359 (O_4359,N_47704,N_47848);
nor UO_4360 (O_4360,N_47753,N_48588);
xnor UO_4361 (O_4361,N_49532,N_48811);
or UO_4362 (O_4362,N_48218,N_47525);
or UO_4363 (O_4363,N_48816,N_47978);
or UO_4364 (O_4364,N_47838,N_49615);
nand UO_4365 (O_4365,N_48178,N_49107);
nand UO_4366 (O_4366,N_49743,N_47974);
xor UO_4367 (O_4367,N_47769,N_48032);
and UO_4368 (O_4368,N_48110,N_48876);
xnor UO_4369 (O_4369,N_48419,N_48552);
or UO_4370 (O_4370,N_48766,N_49584);
xnor UO_4371 (O_4371,N_48654,N_49748);
or UO_4372 (O_4372,N_48854,N_49420);
nand UO_4373 (O_4373,N_48386,N_47937);
xnor UO_4374 (O_4374,N_49039,N_49266);
nand UO_4375 (O_4375,N_49469,N_49176);
nand UO_4376 (O_4376,N_48867,N_49338);
nor UO_4377 (O_4377,N_48597,N_48433);
and UO_4378 (O_4378,N_48777,N_48582);
xnor UO_4379 (O_4379,N_48520,N_47924);
xor UO_4380 (O_4380,N_48510,N_48491);
and UO_4381 (O_4381,N_48681,N_48291);
or UO_4382 (O_4382,N_48644,N_48279);
nand UO_4383 (O_4383,N_48496,N_48337);
or UO_4384 (O_4384,N_48178,N_48859);
nor UO_4385 (O_4385,N_48977,N_49639);
nor UO_4386 (O_4386,N_48972,N_47835);
nor UO_4387 (O_4387,N_49329,N_48568);
nor UO_4388 (O_4388,N_48000,N_49471);
nand UO_4389 (O_4389,N_49344,N_49119);
or UO_4390 (O_4390,N_47816,N_49447);
and UO_4391 (O_4391,N_48556,N_49346);
or UO_4392 (O_4392,N_49771,N_48400);
nand UO_4393 (O_4393,N_49376,N_48067);
xnor UO_4394 (O_4394,N_49124,N_48417);
and UO_4395 (O_4395,N_48367,N_48201);
nand UO_4396 (O_4396,N_47548,N_49656);
or UO_4397 (O_4397,N_49280,N_49339);
and UO_4398 (O_4398,N_47944,N_47687);
xor UO_4399 (O_4399,N_48212,N_48786);
and UO_4400 (O_4400,N_49201,N_48353);
nand UO_4401 (O_4401,N_47740,N_49390);
or UO_4402 (O_4402,N_48632,N_49755);
xor UO_4403 (O_4403,N_49980,N_48325);
xor UO_4404 (O_4404,N_49215,N_49935);
nor UO_4405 (O_4405,N_47795,N_49403);
or UO_4406 (O_4406,N_48151,N_48214);
xor UO_4407 (O_4407,N_49615,N_48282);
nor UO_4408 (O_4408,N_48566,N_49203);
nand UO_4409 (O_4409,N_48266,N_49489);
or UO_4410 (O_4410,N_47606,N_48865);
xor UO_4411 (O_4411,N_48725,N_49580);
nor UO_4412 (O_4412,N_47686,N_48413);
or UO_4413 (O_4413,N_49072,N_48842);
xor UO_4414 (O_4414,N_48723,N_47526);
or UO_4415 (O_4415,N_49746,N_49536);
nand UO_4416 (O_4416,N_49654,N_47811);
nor UO_4417 (O_4417,N_49660,N_49271);
or UO_4418 (O_4418,N_47803,N_47662);
nor UO_4419 (O_4419,N_48444,N_49567);
xor UO_4420 (O_4420,N_48721,N_49859);
nor UO_4421 (O_4421,N_48972,N_48639);
nand UO_4422 (O_4422,N_48163,N_48612);
nand UO_4423 (O_4423,N_47984,N_47907);
nand UO_4424 (O_4424,N_47684,N_49504);
or UO_4425 (O_4425,N_48190,N_49231);
nor UO_4426 (O_4426,N_49948,N_47775);
xor UO_4427 (O_4427,N_47547,N_48771);
xnor UO_4428 (O_4428,N_49282,N_48238);
and UO_4429 (O_4429,N_47540,N_47985);
or UO_4430 (O_4430,N_48534,N_49715);
xor UO_4431 (O_4431,N_47790,N_47828);
or UO_4432 (O_4432,N_47923,N_47824);
nand UO_4433 (O_4433,N_47748,N_48300);
xor UO_4434 (O_4434,N_48824,N_49777);
xor UO_4435 (O_4435,N_49642,N_48260);
nor UO_4436 (O_4436,N_48368,N_49047);
and UO_4437 (O_4437,N_48380,N_47792);
nor UO_4438 (O_4438,N_48270,N_47523);
and UO_4439 (O_4439,N_48303,N_49884);
or UO_4440 (O_4440,N_48035,N_49363);
nor UO_4441 (O_4441,N_49888,N_48749);
and UO_4442 (O_4442,N_48253,N_48430);
nor UO_4443 (O_4443,N_48351,N_49479);
xnor UO_4444 (O_4444,N_48912,N_47511);
and UO_4445 (O_4445,N_48160,N_49756);
xnor UO_4446 (O_4446,N_48136,N_49486);
nor UO_4447 (O_4447,N_47793,N_48402);
or UO_4448 (O_4448,N_48351,N_48032);
or UO_4449 (O_4449,N_48651,N_49214);
or UO_4450 (O_4450,N_48323,N_49289);
nor UO_4451 (O_4451,N_48284,N_48704);
or UO_4452 (O_4452,N_48614,N_49227);
nand UO_4453 (O_4453,N_47791,N_49758);
nand UO_4454 (O_4454,N_48939,N_49475);
nand UO_4455 (O_4455,N_49052,N_49515);
or UO_4456 (O_4456,N_49118,N_48060);
or UO_4457 (O_4457,N_48774,N_48711);
xnor UO_4458 (O_4458,N_49725,N_49687);
nor UO_4459 (O_4459,N_49851,N_49506);
nor UO_4460 (O_4460,N_49390,N_47867);
nand UO_4461 (O_4461,N_48988,N_49402);
and UO_4462 (O_4462,N_49250,N_48196);
and UO_4463 (O_4463,N_48111,N_48529);
and UO_4464 (O_4464,N_49912,N_49965);
and UO_4465 (O_4465,N_47860,N_49089);
xor UO_4466 (O_4466,N_48074,N_48300);
nand UO_4467 (O_4467,N_48744,N_49429);
or UO_4468 (O_4468,N_47870,N_49914);
and UO_4469 (O_4469,N_49170,N_48015);
and UO_4470 (O_4470,N_48245,N_48109);
and UO_4471 (O_4471,N_49078,N_49581);
xor UO_4472 (O_4472,N_48204,N_48227);
or UO_4473 (O_4473,N_48013,N_49525);
nand UO_4474 (O_4474,N_48964,N_48676);
nor UO_4475 (O_4475,N_49104,N_48339);
or UO_4476 (O_4476,N_48391,N_48143);
and UO_4477 (O_4477,N_49452,N_47901);
nor UO_4478 (O_4478,N_48684,N_48147);
or UO_4479 (O_4479,N_48608,N_48692);
nor UO_4480 (O_4480,N_49096,N_48304);
xnor UO_4481 (O_4481,N_48336,N_48252);
or UO_4482 (O_4482,N_49623,N_49023);
and UO_4483 (O_4483,N_48817,N_49868);
nand UO_4484 (O_4484,N_49018,N_49172);
and UO_4485 (O_4485,N_47623,N_49783);
xnor UO_4486 (O_4486,N_47941,N_48995);
and UO_4487 (O_4487,N_48402,N_49142);
and UO_4488 (O_4488,N_47684,N_49107);
xor UO_4489 (O_4489,N_48248,N_49922);
and UO_4490 (O_4490,N_48101,N_47967);
nor UO_4491 (O_4491,N_48262,N_47760);
or UO_4492 (O_4492,N_48860,N_49109);
nor UO_4493 (O_4493,N_48193,N_49720);
and UO_4494 (O_4494,N_49151,N_47864);
and UO_4495 (O_4495,N_47841,N_48470);
xor UO_4496 (O_4496,N_49945,N_47976);
xnor UO_4497 (O_4497,N_49154,N_48923);
nor UO_4498 (O_4498,N_48118,N_47933);
or UO_4499 (O_4499,N_49411,N_49740);
nand UO_4500 (O_4500,N_49897,N_48315);
nor UO_4501 (O_4501,N_48639,N_49643);
or UO_4502 (O_4502,N_48304,N_47934);
or UO_4503 (O_4503,N_49788,N_49875);
or UO_4504 (O_4504,N_49009,N_49869);
or UO_4505 (O_4505,N_48085,N_47571);
or UO_4506 (O_4506,N_49897,N_48546);
xor UO_4507 (O_4507,N_49853,N_49818);
and UO_4508 (O_4508,N_48262,N_49244);
nor UO_4509 (O_4509,N_49077,N_47703);
or UO_4510 (O_4510,N_49572,N_47630);
xor UO_4511 (O_4511,N_47707,N_49190);
and UO_4512 (O_4512,N_48303,N_49798);
xnor UO_4513 (O_4513,N_48813,N_48705);
xor UO_4514 (O_4514,N_49537,N_49242);
nor UO_4515 (O_4515,N_48278,N_49315);
nor UO_4516 (O_4516,N_47800,N_48691);
xor UO_4517 (O_4517,N_49800,N_49107);
or UO_4518 (O_4518,N_48235,N_48056);
or UO_4519 (O_4519,N_49299,N_48857);
or UO_4520 (O_4520,N_48404,N_47693);
xnor UO_4521 (O_4521,N_47663,N_49488);
nor UO_4522 (O_4522,N_48315,N_49049);
nand UO_4523 (O_4523,N_48724,N_48428);
and UO_4524 (O_4524,N_49029,N_49857);
xor UO_4525 (O_4525,N_47890,N_49353);
or UO_4526 (O_4526,N_48631,N_48292);
nand UO_4527 (O_4527,N_49186,N_48901);
nand UO_4528 (O_4528,N_48671,N_49483);
xor UO_4529 (O_4529,N_48411,N_47631);
and UO_4530 (O_4530,N_47917,N_47638);
and UO_4531 (O_4531,N_48379,N_49727);
or UO_4532 (O_4532,N_48675,N_48583);
or UO_4533 (O_4533,N_49394,N_49915);
and UO_4534 (O_4534,N_47697,N_49292);
nand UO_4535 (O_4535,N_49851,N_47630);
nor UO_4536 (O_4536,N_48011,N_49783);
or UO_4537 (O_4537,N_48673,N_49968);
xnor UO_4538 (O_4538,N_47684,N_48593);
nor UO_4539 (O_4539,N_47699,N_47564);
or UO_4540 (O_4540,N_47555,N_49182);
xor UO_4541 (O_4541,N_49901,N_48641);
nand UO_4542 (O_4542,N_49828,N_47606);
xor UO_4543 (O_4543,N_47953,N_48974);
xnor UO_4544 (O_4544,N_47853,N_48391);
nand UO_4545 (O_4545,N_49646,N_48789);
or UO_4546 (O_4546,N_49084,N_49757);
or UO_4547 (O_4547,N_48433,N_49452);
and UO_4548 (O_4548,N_48406,N_47821);
xor UO_4549 (O_4549,N_49839,N_48060);
or UO_4550 (O_4550,N_48504,N_49421);
nor UO_4551 (O_4551,N_49675,N_49644);
xor UO_4552 (O_4552,N_48911,N_49124);
nor UO_4553 (O_4553,N_47571,N_49138);
and UO_4554 (O_4554,N_48194,N_49256);
xor UO_4555 (O_4555,N_49319,N_49849);
nand UO_4556 (O_4556,N_48129,N_47876);
xor UO_4557 (O_4557,N_48715,N_47760);
xnor UO_4558 (O_4558,N_47624,N_48209);
nand UO_4559 (O_4559,N_47737,N_48929);
nor UO_4560 (O_4560,N_48892,N_48210);
and UO_4561 (O_4561,N_49366,N_47699);
nor UO_4562 (O_4562,N_49729,N_48780);
and UO_4563 (O_4563,N_49965,N_49964);
or UO_4564 (O_4564,N_48090,N_48477);
nand UO_4565 (O_4565,N_49352,N_48074);
or UO_4566 (O_4566,N_49554,N_47870);
or UO_4567 (O_4567,N_47876,N_49780);
and UO_4568 (O_4568,N_48209,N_48244);
xnor UO_4569 (O_4569,N_49704,N_49894);
or UO_4570 (O_4570,N_49999,N_47860);
and UO_4571 (O_4571,N_47663,N_49741);
xnor UO_4572 (O_4572,N_49746,N_47778);
nand UO_4573 (O_4573,N_47810,N_49871);
or UO_4574 (O_4574,N_48255,N_48099);
nor UO_4575 (O_4575,N_49313,N_47976);
nand UO_4576 (O_4576,N_49631,N_48342);
nor UO_4577 (O_4577,N_49885,N_48377);
or UO_4578 (O_4578,N_48745,N_47825);
xnor UO_4579 (O_4579,N_47884,N_47989);
and UO_4580 (O_4580,N_49167,N_49824);
and UO_4581 (O_4581,N_47952,N_49994);
and UO_4582 (O_4582,N_49404,N_49922);
or UO_4583 (O_4583,N_48603,N_47827);
and UO_4584 (O_4584,N_47509,N_48171);
nor UO_4585 (O_4585,N_47802,N_48936);
and UO_4586 (O_4586,N_49759,N_49832);
and UO_4587 (O_4587,N_49111,N_47793);
nor UO_4588 (O_4588,N_49306,N_48472);
nor UO_4589 (O_4589,N_49063,N_49270);
or UO_4590 (O_4590,N_49769,N_48388);
xor UO_4591 (O_4591,N_49970,N_49783);
nor UO_4592 (O_4592,N_48071,N_47982);
xor UO_4593 (O_4593,N_48046,N_48566);
or UO_4594 (O_4594,N_47915,N_47786);
nand UO_4595 (O_4595,N_48382,N_49644);
nand UO_4596 (O_4596,N_49028,N_49032);
nor UO_4597 (O_4597,N_49675,N_48019);
nor UO_4598 (O_4598,N_47996,N_48851);
nand UO_4599 (O_4599,N_49215,N_48330);
nor UO_4600 (O_4600,N_48785,N_47538);
and UO_4601 (O_4601,N_49252,N_49917);
nand UO_4602 (O_4602,N_47579,N_49417);
xnor UO_4603 (O_4603,N_49097,N_48740);
nor UO_4604 (O_4604,N_48063,N_49728);
or UO_4605 (O_4605,N_49322,N_49456);
and UO_4606 (O_4606,N_47983,N_48484);
nor UO_4607 (O_4607,N_47783,N_49327);
and UO_4608 (O_4608,N_49438,N_48339);
nor UO_4609 (O_4609,N_48397,N_48881);
and UO_4610 (O_4610,N_48354,N_49519);
and UO_4611 (O_4611,N_48656,N_49873);
nor UO_4612 (O_4612,N_49302,N_49868);
or UO_4613 (O_4613,N_49673,N_48428);
nand UO_4614 (O_4614,N_49390,N_49317);
or UO_4615 (O_4615,N_48549,N_48505);
or UO_4616 (O_4616,N_49531,N_47942);
nand UO_4617 (O_4617,N_48175,N_49907);
and UO_4618 (O_4618,N_48187,N_49269);
or UO_4619 (O_4619,N_48178,N_48835);
nand UO_4620 (O_4620,N_49769,N_47954);
and UO_4621 (O_4621,N_49871,N_47593);
or UO_4622 (O_4622,N_49669,N_49250);
nand UO_4623 (O_4623,N_48026,N_48172);
or UO_4624 (O_4624,N_47542,N_47722);
xnor UO_4625 (O_4625,N_49209,N_47619);
and UO_4626 (O_4626,N_48219,N_49936);
xnor UO_4627 (O_4627,N_48376,N_47746);
and UO_4628 (O_4628,N_49734,N_47811);
xor UO_4629 (O_4629,N_49719,N_47600);
or UO_4630 (O_4630,N_49700,N_49144);
nand UO_4631 (O_4631,N_49311,N_48488);
xnor UO_4632 (O_4632,N_49508,N_48442);
nor UO_4633 (O_4633,N_48682,N_49829);
xor UO_4634 (O_4634,N_49096,N_49345);
nor UO_4635 (O_4635,N_48767,N_48130);
or UO_4636 (O_4636,N_49340,N_48447);
nor UO_4637 (O_4637,N_48254,N_48621);
and UO_4638 (O_4638,N_49604,N_49273);
nand UO_4639 (O_4639,N_47986,N_48660);
or UO_4640 (O_4640,N_49115,N_49966);
and UO_4641 (O_4641,N_49368,N_48783);
nor UO_4642 (O_4642,N_49746,N_47974);
nor UO_4643 (O_4643,N_49568,N_47871);
nor UO_4644 (O_4644,N_47825,N_48268);
nand UO_4645 (O_4645,N_47817,N_47585);
or UO_4646 (O_4646,N_49521,N_49574);
nor UO_4647 (O_4647,N_48968,N_49301);
or UO_4648 (O_4648,N_49438,N_48663);
or UO_4649 (O_4649,N_49610,N_47898);
nor UO_4650 (O_4650,N_48703,N_48834);
nand UO_4651 (O_4651,N_47717,N_48090);
or UO_4652 (O_4652,N_49023,N_49376);
nand UO_4653 (O_4653,N_49255,N_49581);
nor UO_4654 (O_4654,N_49609,N_49316);
nand UO_4655 (O_4655,N_49505,N_47524);
xnor UO_4656 (O_4656,N_49073,N_49727);
nand UO_4657 (O_4657,N_48790,N_48827);
and UO_4658 (O_4658,N_47897,N_47637);
nand UO_4659 (O_4659,N_49389,N_48393);
nor UO_4660 (O_4660,N_47551,N_49253);
nand UO_4661 (O_4661,N_49317,N_48125);
xor UO_4662 (O_4662,N_47988,N_49737);
xnor UO_4663 (O_4663,N_49637,N_49788);
or UO_4664 (O_4664,N_48719,N_49712);
or UO_4665 (O_4665,N_49493,N_49459);
xnor UO_4666 (O_4666,N_48275,N_47707);
or UO_4667 (O_4667,N_49232,N_49052);
nand UO_4668 (O_4668,N_49274,N_48575);
nand UO_4669 (O_4669,N_49967,N_47538);
nand UO_4670 (O_4670,N_47597,N_49070);
and UO_4671 (O_4671,N_47767,N_47952);
and UO_4672 (O_4672,N_48945,N_48605);
and UO_4673 (O_4673,N_48503,N_47937);
and UO_4674 (O_4674,N_47807,N_49033);
nor UO_4675 (O_4675,N_48095,N_49995);
or UO_4676 (O_4676,N_48979,N_48677);
nand UO_4677 (O_4677,N_48637,N_48976);
nor UO_4678 (O_4678,N_47523,N_49624);
nor UO_4679 (O_4679,N_48312,N_49328);
xor UO_4680 (O_4680,N_49993,N_48893);
and UO_4681 (O_4681,N_48025,N_48090);
or UO_4682 (O_4682,N_47874,N_49292);
nand UO_4683 (O_4683,N_49929,N_49834);
nand UO_4684 (O_4684,N_48213,N_49820);
and UO_4685 (O_4685,N_49775,N_49344);
xor UO_4686 (O_4686,N_48619,N_47943);
nand UO_4687 (O_4687,N_49860,N_47555);
nand UO_4688 (O_4688,N_47845,N_49897);
or UO_4689 (O_4689,N_48724,N_49347);
nor UO_4690 (O_4690,N_49747,N_49646);
nor UO_4691 (O_4691,N_48205,N_48201);
and UO_4692 (O_4692,N_47740,N_49705);
nand UO_4693 (O_4693,N_49379,N_49454);
nand UO_4694 (O_4694,N_48522,N_49313);
nand UO_4695 (O_4695,N_49229,N_48418);
or UO_4696 (O_4696,N_48879,N_48615);
nand UO_4697 (O_4697,N_48690,N_48848);
nor UO_4698 (O_4698,N_49656,N_47886);
nand UO_4699 (O_4699,N_47897,N_49561);
or UO_4700 (O_4700,N_49382,N_48152);
and UO_4701 (O_4701,N_48290,N_49746);
or UO_4702 (O_4702,N_47652,N_48553);
or UO_4703 (O_4703,N_48917,N_49193);
xnor UO_4704 (O_4704,N_49322,N_48541);
xor UO_4705 (O_4705,N_49119,N_48550);
nand UO_4706 (O_4706,N_48423,N_47786);
and UO_4707 (O_4707,N_48518,N_49210);
or UO_4708 (O_4708,N_48788,N_48782);
xnor UO_4709 (O_4709,N_47560,N_49584);
or UO_4710 (O_4710,N_48899,N_48640);
or UO_4711 (O_4711,N_48509,N_49012);
and UO_4712 (O_4712,N_48910,N_49105);
nand UO_4713 (O_4713,N_47642,N_49191);
nand UO_4714 (O_4714,N_48215,N_48748);
nand UO_4715 (O_4715,N_48968,N_49952);
and UO_4716 (O_4716,N_48099,N_47612);
xor UO_4717 (O_4717,N_49029,N_47864);
nor UO_4718 (O_4718,N_48090,N_48037);
nor UO_4719 (O_4719,N_49321,N_48121);
nor UO_4720 (O_4720,N_49219,N_49171);
or UO_4721 (O_4721,N_47818,N_49983);
nand UO_4722 (O_4722,N_49715,N_49109);
xor UO_4723 (O_4723,N_48373,N_48185);
nand UO_4724 (O_4724,N_49021,N_48751);
or UO_4725 (O_4725,N_48930,N_49344);
xor UO_4726 (O_4726,N_47646,N_49452);
or UO_4727 (O_4727,N_49182,N_47917);
and UO_4728 (O_4728,N_49138,N_49409);
and UO_4729 (O_4729,N_48822,N_49338);
or UO_4730 (O_4730,N_49373,N_49615);
nand UO_4731 (O_4731,N_48411,N_48862);
nand UO_4732 (O_4732,N_48512,N_49988);
or UO_4733 (O_4733,N_47515,N_49390);
nand UO_4734 (O_4734,N_49076,N_49550);
nor UO_4735 (O_4735,N_47634,N_48795);
nand UO_4736 (O_4736,N_49180,N_48339);
xnor UO_4737 (O_4737,N_48557,N_49047);
and UO_4738 (O_4738,N_47511,N_47619);
nor UO_4739 (O_4739,N_49333,N_49598);
and UO_4740 (O_4740,N_49215,N_48334);
xnor UO_4741 (O_4741,N_47968,N_49891);
or UO_4742 (O_4742,N_48379,N_48279);
nor UO_4743 (O_4743,N_49349,N_48545);
nand UO_4744 (O_4744,N_48518,N_47915);
and UO_4745 (O_4745,N_49049,N_48231);
xor UO_4746 (O_4746,N_49390,N_49319);
xnor UO_4747 (O_4747,N_49643,N_48661);
and UO_4748 (O_4748,N_48274,N_49257);
xor UO_4749 (O_4749,N_47729,N_48045);
xor UO_4750 (O_4750,N_47589,N_47757);
nor UO_4751 (O_4751,N_48482,N_49012);
or UO_4752 (O_4752,N_47948,N_49458);
xor UO_4753 (O_4753,N_48369,N_48035);
or UO_4754 (O_4754,N_47749,N_48654);
and UO_4755 (O_4755,N_48060,N_47946);
or UO_4756 (O_4756,N_49174,N_47579);
or UO_4757 (O_4757,N_48020,N_48949);
nor UO_4758 (O_4758,N_48648,N_47975);
and UO_4759 (O_4759,N_49161,N_49503);
xnor UO_4760 (O_4760,N_49012,N_48827);
or UO_4761 (O_4761,N_48928,N_49105);
or UO_4762 (O_4762,N_48167,N_49854);
xnor UO_4763 (O_4763,N_47949,N_49807);
and UO_4764 (O_4764,N_48414,N_49483);
and UO_4765 (O_4765,N_48858,N_49568);
xor UO_4766 (O_4766,N_47822,N_49728);
nor UO_4767 (O_4767,N_49836,N_49921);
nor UO_4768 (O_4768,N_48933,N_48271);
and UO_4769 (O_4769,N_48351,N_49932);
nor UO_4770 (O_4770,N_49033,N_49757);
nand UO_4771 (O_4771,N_49853,N_48129);
and UO_4772 (O_4772,N_49971,N_48114);
xnor UO_4773 (O_4773,N_49398,N_48198);
nor UO_4774 (O_4774,N_47617,N_49955);
nand UO_4775 (O_4775,N_49920,N_48126);
and UO_4776 (O_4776,N_48274,N_49903);
nand UO_4777 (O_4777,N_47939,N_49689);
nand UO_4778 (O_4778,N_48509,N_49579);
and UO_4779 (O_4779,N_48678,N_49527);
xor UO_4780 (O_4780,N_47915,N_48397);
xnor UO_4781 (O_4781,N_47637,N_49621);
xnor UO_4782 (O_4782,N_48659,N_49176);
xnor UO_4783 (O_4783,N_47600,N_47628);
nor UO_4784 (O_4784,N_49275,N_48850);
xnor UO_4785 (O_4785,N_47703,N_49627);
xnor UO_4786 (O_4786,N_49426,N_49572);
or UO_4787 (O_4787,N_49036,N_48215);
xnor UO_4788 (O_4788,N_47826,N_49305);
nand UO_4789 (O_4789,N_48671,N_49329);
nor UO_4790 (O_4790,N_49044,N_49021);
nand UO_4791 (O_4791,N_48434,N_48077);
nor UO_4792 (O_4792,N_49554,N_49789);
xnor UO_4793 (O_4793,N_48972,N_49964);
xor UO_4794 (O_4794,N_48369,N_49087);
and UO_4795 (O_4795,N_47831,N_49342);
and UO_4796 (O_4796,N_48349,N_48524);
or UO_4797 (O_4797,N_49989,N_48153);
nor UO_4798 (O_4798,N_48010,N_48151);
xnor UO_4799 (O_4799,N_47658,N_48871);
nor UO_4800 (O_4800,N_48353,N_49441);
xnor UO_4801 (O_4801,N_48575,N_48285);
or UO_4802 (O_4802,N_49884,N_49967);
xor UO_4803 (O_4803,N_47592,N_48499);
nor UO_4804 (O_4804,N_49258,N_49029);
xnor UO_4805 (O_4805,N_49243,N_49542);
nand UO_4806 (O_4806,N_47655,N_49157);
nand UO_4807 (O_4807,N_49405,N_48713);
or UO_4808 (O_4808,N_49060,N_48635);
nand UO_4809 (O_4809,N_48487,N_48820);
or UO_4810 (O_4810,N_47998,N_49904);
nor UO_4811 (O_4811,N_48398,N_49042);
and UO_4812 (O_4812,N_49324,N_49143);
xor UO_4813 (O_4813,N_47752,N_49605);
and UO_4814 (O_4814,N_48305,N_49613);
and UO_4815 (O_4815,N_49296,N_49550);
xor UO_4816 (O_4816,N_47790,N_49769);
nand UO_4817 (O_4817,N_49865,N_49746);
xor UO_4818 (O_4818,N_49004,N_49438);
xnor UO_4819 (O_4819,N_48893,N_48962);
nor UO_4820 (O_4820,N_48171,N_47951);
or UO_4821 (O_4821,N_48763,N_48125);
nand UO_4822 (O_4822,N_49729,N_49061);
or UO_4823 (O_4823,N_49725,N_49205);
xnor UO_4824 (O_4824,N_49282,N_47922);
xor UO_4825 (O_4825,N_48353,N_48947);
and UO_4826 (O_4826,N_47964,N_47871);
and UO_4827 (O_4827,N_48905,N_49465);
or UO_4828 (O_4828,N_47998,N_48941);
and UO_4829 (O_4829,N_49147,N_48042);
nand UO_4830 (O_4830,N_47881,N_49712);
or UO_4831 (O_4831,N_48607,N_49172);
nand UO_4832 (O_4832,N_48613,N_48143);
nor UO_4833 (O_4833,N_48999,N_48167);
or UO_4834 (O_4834,N_49619,N_47839);
nor UO_4835 (O_4835,N_48118,N_49826);
xor UO_4836 (O_4836,N_48000,N_49890);
nor UO_4837 (O_4837,N_47990,N_47817);
nand UO_4838 (O_4838,N_49455,N_47943);
nand UO_4839 (O_4839,N_49174,N_49580);
xor UO_4840 (O_4840,N_49397,N_49705);
or UO_4841 (O_4841,N_48395,N_49273);
or UO_4842 (O_4842,N_49194,N_47714);
and UO_4843 (O_4843,N_48507,N_49064);
and UO_4844 (O_4844,N_48417,N_49674);
and UO_4845 (O_4845,N_49430,N_49401);
or UO_4846 (O_4846,N_48035,N_47926);
nor UO_4847 (O_4847,N_48716,N_49505);
or UO_4848 (O_4848,N_48790,N_48082);
or UO_4849 (O_4849,N_49727,N_47981);
or UO_4850 (O_4850,N_49912,N_47725);
nand UO_4851 (O_4851,N_47788,N_49445);
and UO_4852 (O_4852,N_48434,N_48809);
and UO_4853 (O_4853,N_48719,N_49694);
nor UO_4854 (O_4854,N_48902,N_49859);
xor UO_4855 (O_4855,N_48118,N_48850);
xor UO_4856 (O_4856,N_49468,N_47541);
xor UO_4857 (O_4857,N_48926,N_49428);
nor UO_4858 (O_4858,N_48590,N_48034);
or UO_4859 (O_4859,N_49576,N_48677);
and UO_4860 (O_4860,N_48818,N_48829);
and UO_4861 (O_4861,N_48548,N_49024);
or UO_4862 (O_4862,N_48943,N_49326);
nand UO_4863 (O_4863,N_47573,N_48989);
xor UO_4864 (O_4864,N_47696,N_48778);
or UO_4865 (O_4865,N_48713,N_48558);
and UO_4866 (O_4866,N_47865,N_49079);
or UO_4867 (O_4867,N_48446,N_49499);
and UO_4868 (O_4868,N_48367,N_48172);
or UO_4869 (O_4869,N_47741,N_48242);
nand UO_4870 (O_4870,N_49474,N_49843);
or UO_4871 (O_4871,N_49722,N_47769);
xor UO_4872 (O_4872,N_49322,N_48297);
and UO_4873 (O_4873,N_48065,N_49359);
and UO_4874 (O_4874,N_49106,N_49624);
xor UO_4875 (O_4875,N_47630,N_48725);
nor UO_4876 (O_4876,N_49694,N_48684);
nand UO_4877 (O_4877,N_48643,N_48521);
nand UO_4878 (O_4878,N_47740,N_48793);
and UO_4879 (O_4879,N_49822,N_48802);
or UO_4880 (O_4880,N_47523,N_49493);
or UO_4881 (O_4881,N_48039,N_48025);
nand UO_4882 (O_4882,N_47624,N_48521);
and UO_4883 (O_4883,N_47814,N_49248);
xor UO_4884 (O_4884,N_49792,N_48025);
and UO_4885 (O_4885,N_48041,N_47991);
nor UO_4886 (O_4886,N_48291,N_49469);
xor UO_4887 (O_4887,N_48792,N_49323);
nor UO_4888 (O_4888,N_49865,N_49978);
xnor UO_4889 (O_4889,N_48072,N_49617);
and UO_4890 (O_4890,N_47619,N_49202);
and UO_4891 (O_4891,N_49753,N_49410);
or UO_4892 (O_4892,N_49072,N_49082);
or UO_4893 (O_4893,N_47997,N_49328);
and UO_4894 (O_4894,N_48506,N_48713);
and UO_4895 (O_4895,N_48290,N_49581);
or UO_4896 (O_4896,N_48415,N_48653);
nor UO_4897 (O_4897,N_48106,N_49788);
or UO_4898 (O_4898,N_47846,N_49094);
nor UO_4899 (O_4899,N_49174,N_48391);
xnor UO_4900 (O_4900,N_49439,N_47579);
xor UO_4901 (O_4901,N_48104,N_48948);
xnor UO_4902 (O_4902,N_49648,N_47755);
or UO_4903 (O_4903,N_47929,N_49085);
nor UO_4904 (O_4904,N_49381,N_49604);
nor UO_4905 (O_4905,N_47718,N_48110);
nand UO_4906 (O_4906,N_48611,N_48996);
or UO_4907 (O_4907,N_49718,N_49210);
nor UO_4908 (O_4908,N_48564,N_49497);
and UO_4909 (O_4909,N_48033,N_49496);
xor UO_4910 (O_4910,N_48451,N_48683);
xor UO_4911 (O_4911,N_48148,N_48343);
xnor UO_4912 (O_4912,N_49196,N_49527);
nor UO_4913 (O_4913,N_49903,N_49581);
or UO_4914 (O_4914,N_48298,N_48567);
or UO_4915 (O_4915,N_47925,N_48521);
and UO_4916 (O_4916,N_48094,N_48137);
xnor UO_4917 (O_4917,N_48892,N_48407);
xnor UO_4918 (O_4918,N_49515,N_49005);
nand UO_4919 (O_4919,N_49221,N_48614);
and UO_4920 (O_4920,N_49985,N_49487);
xnor UO_4921 (O_4921,N_48753,N_48066);
or UO_4922 (O_4922,N_49987,N_48158);
nor UO_4923 (O_4923,N_48786,N_47639);
nor UO_4924 (O_4924,N_49689,N_49449);
xnor UO_4925 (O_4925,N_49633,N_47531);
nand UO_4926 (O_4926,N_47624,N_49155);
and UO_4927 (O_4927,N_49214,N_48420);
xnor UO_4928 (O_4928,N_49204,N_47581);
or UO_4929 (O_4929,N_47795,N_49913);
nand UO_4930 (O_4930,N_49869,N_48078);
xnor UO_4931 (O_4931,N_48956,N_47705);
xor UO_4932 (O_4932,N_48417,N_49285);
nand UO_4933 (O_4933,N_49747,N_48822);
nor UO_4934 (O_4934,N_48099,N_49150);
nand UO_4935 (O_4935,N_48208,N_48095);
nand UO_4936 (O_4936,N_47782,N_49784);
nor UO_4937 (O_4937,N_47956,N_48032);
or UO_4938 (O_4938,N_49610,N_49221);
xor UO_4939 (O_4939,N_47618,N_49708);
nor UO_4940 (O_4940,N_49067,N_47928);
nand UO_4941 (O_4941,N_49158,N_49011);
or UO_4942 (O_4942,N_48197,N_49044);
or UO_4943 (O_4943,N_48424,N_47637);
or UO_4944 (O_4944,N_49730,N_47633);
nor UO_4945 (O_4945,N_49999,N_48693);
xor UO_4946 (O_4946,N_48422,N_49132);
nand UO_4947 (O_4947,N_48036,N_49311);
or UO_4948 (O_4948,N_49769,N_49669);
and UO_4949 (O_4949,N_47769,N_47752);
nor UO_4950 (O_4950,N_48091,N_48268);
nor UO_4951 (O_4951,N_49275,N_47929);
or UO_4952 (O_4952,N_48580,N_49733);
nor UO_4953 (O_4953,N_48897,N_47939);
or UO_4954 (O_4954,N_48892,N_49519);
nand UO_4955 (O_4955,N_48304,N_47710);
and UO_4956 (O_4956,N_48364,N_49662);
nor UO_4957 (O_4957,N_49855,N_49132);
nor UO_4958 (O_4958,N_47572,N_47595);
and UO_4959 (O_4959,N_47847,N_48205);
or UO_4960 (O_4960,N_49132,N_47734);
and UO_4961 (O_4961,N_48168,N_48771);
or UO_4962 (O_4962,N_48113,N_47954);
or UO_4963 (O_4963,N_49270,N_48979);
nor UO_4964 (O_4964,N_49734,N_49249);
and UO_4965 (O_4965,N_47953,N_49269);
nor UO_4966 (O_4966,N_49103,N_48076);
nor UO_4967 (O_4967,N_48348,N_49398);
or UO_4968 (O_4968,N_47896,N_48798);
nand UO_4969 (O_4969,N_49601,N_47512);
and UO_4970 (O_4970,N_48510,N_49513);
nand UO_4971 (O_4971,N_47574,N_49266);
or UO_4972 (O_4972,N_47883,N_47500);
nand UO_4973 (O_4973,N_49786,N_48394);
and UO_4974 (O_4974,N_48635,N_49814);
nand UO_4975 (O_4975,N_48573,N_48069);
nor UO_4976 (O_4976,N_49834,N_48644);
nor UO_4977 (O_4977,N_48618,N_47965);
and UO_4978 (O_4978,N_49527,N_47973);
or UO_4979 (O_4979,N_48759,N_48927);
nand UO_4980 (O_4980,N_48829,N_48949);
nand UO_4981 (O_4981,N_47881,N_48940);
xnor UO_4982 (O_4982,N_47630,N_49080);
or UO_4983 (O_4983,N_48291,N_48303);
nor UO_4984 (O_4984,N_48351,N_49552);
or UO_4985 (O_4985,N_49467,N_47501);
or UO_4986 (O_4986,N_49309,N_47521);
or UO_4987 (O_4987,N_48665,N_48959);
nor UO_4988 (O_4988,N_49820,N_48842);
nand UO_4989 (O_4989,N_49003,N_47982);
or UO_4990 (O_4990,N_49563,N_49821);
and UO_4991 (O_4991,N_48363,N_49567);
or UO_4992 (O_4992,N_48968,N_49697);
and UO_4993 (O_4993,N_49986,N_47558);
and UO_4994 (O_4994,N_49206,N_48721);
xor UO_4995 (O_4995,N_48336,N_48596);
or UO_4996 (O_4996,N_49669,N_47990);
nor UO_4997 (O_4997,N_48645,N_48616);
nand UO_4998 (O_4998,N_48060,N_48781);
or UO_4999 (O_4999,N_47911,N_48872);
endmodule