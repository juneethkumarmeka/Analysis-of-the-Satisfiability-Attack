module basic_750_5000_1000_2_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2503,N_2504,N_2505,N_2506,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2525,N_2526,N_2527,N_2528,N_2530,N_2532,N_2533,N_2534,N_2535,N_2537,N_2538,N_2540,N_2541,N_2542,N_2543,N_2545,N_2547,N_2548,N_2549,N_2551,N_2552,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2582,N_2585,N_2586,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2602,N_2603,N_2606,N_2607,N_2608,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2626,N_2627,N_2630,N_2631,N_2632,N_2634,N_2636,N_2637,N_2638,N_2639,N_2640,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2660,N_2661,N_2662,N_2664,N_2665,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2687,N_2688,N_2689,N_2691,N_2692,N_2693,N_2696,N_2697,N_2698,N_2699,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2709,N_2710,N_2713,N_2714,N_2715,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2724,N_2725,N_2726,N_2727,N_2728,N_2730,N_2733,N_2734,N_2735,N_2736,N_2738,N_2739,N_2740,N_2741,N_2742,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2752,N_2754,N_2756,N_2757,N_2758,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2783,N_2784,N_2786,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2798,N_2799,N_2800,N_2803,N_2805,N_2807,N_2808,N_2809,N_2810,N_2813,N_2814,N_2815,N_2816,N_2817,N_2819,N_2821,N_2823,N_2824,N_2825,N_2827,N_2829,N_2831,N_2832,N_2833,N_2834,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2882,N_2887,N_2888,N_2889,N_2890,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2903,N_2904,N_2905,N_2906,N_2908,N_2909,N_2910,N_2912,N_2913,N_2914,N_2915,N_2917,N_2918,N_2919,N_2920,N_2923,N_2924,N_2926,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2963,N_2964,N_2965,N_2967,N_2969,N_2970,N_2971,N_2972,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2987,N_2988,N_2989,N_2990,N_2991,N_2993,N_2995,N_2996,N_2998,N_3000,N_3001,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3012,N_3013,N_3014,N_3017,N_3018,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3027,N_3028,N_3030,N_3032,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3072,N_3073,N_3074,N_3075,N_3076,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3123,N_3124,N_3125,N_3126,N_3128,N_3129,N_3130,N_3131,N_3133,N_3135,N_3136,N_3137,N_3138,N_3139,N_3141,N_3142,N_3143,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3155,N_3156,N_3157,N_3158,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3171,N_3172,N_3173,N_3174,N_3177,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3195,N_3196,N_3198,N_3200,N_3201,N_3202,N_3204,N_3205,N_3206,N_3208,N_3211,N_3212,N_3213,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3239,N_3240,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3250,N_3251,N_3252,N_3253,N_3254,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3270,N_3271,N_3272,N_3273,N_3275,N_3276,N_3277,N_3278,N_3279,N_3281,N_3282,N_3283,N_3284,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3299,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3312,N_3313,N_3314,N_3316,N_3317,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3328,N_3329,N_3330,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3341,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3370,N_3371,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3415,N_3416,N_3417,N_3418,N_3420,N_3421,N_3422,N_3424,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3462,N_3463,N_3464,N_3465,N_3467,N_3468,N_3469,N_3470,N_3471,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3489,N_3490,N_3491,N_3493,N_3495,N_3496,N_3497,N_3501,N_3502,N_3503,N_3504,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3536,N_3537,N_3538,N_3539,N_3540,N_3542,N_3544,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3561,N_3562,N_3563,N_3564,N_3565,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3574,N_3575,N_3576,N_3577,N_3579,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3592,N_3593,N_3594,N_3595,N_3596,N_3598,N_3599,N_3600,N_3601,N_3602,N_3605,N_3606,N_3608,N_3609,N_3610,N_3611,N_3613,N_3614,N_3615,N_3617,N_3619,N_3620,N_3621,N_3622,N_3624,N_3625,N_3626,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3637,N_3638,N_3639,N_3643,N_3644,N_3645,N_3646,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3667,N_3669,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3679,N_3680,N_3681,N_3682,N_3684,N_3685,N_3686,N_3688,N_3689,N_3690,N_3692,N_3693,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3704,N_3705,N_3706,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3730,N_3731,N_3732,N_3734,N_3735,N_3736,N_3738,N_3739,N_3740,N_3741,N_3743,N_3744,N_3745,N_3746,N_3747,N_3749,N_3750,N_3751,N_3752,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3765,N_3766,N_3767,N_3768,N_3769,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3782,N_3783,N_3784,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3795,N_3796,N_3797,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3808,N_3810,N_3811,N_3813,N_3814,N_3815,N_3816,N_3817,N_3819,N_3820,N_3821,N_3823,N_3824,N_3828,N_3829,N_3830,N_3831,N_3832,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3845,N_3847,N_3849,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3870,N_3872,N_3874,N_3876,N_3877,N_3878,N_3879,N_3881,N_3883,N_3885,N_3886,N_3888,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3909,N_3910,N_3913,N_3915,N_3916,N_3917,N_3918,N_3921,N_3922,N_3923,N_3925,N_3926,N_3927,N_3929,N_3930,N_3931,N_3933,N_3935,N_3936,N_3938,N_3939,N_3941,N_3943,N_3944,N_3945,N_3946,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3960,N_3961,N_3962,N_3963,N_3965,N_3966,N_3967,N_3969,N_3970,N_3974,N_3975,N_3976,N_3977,N_3979,N_3980,N_3981,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3995,N_3996,N_3997,N_3998,N_4000,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4010,N_4013,N_4014,N_4016,N_4017,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4026,N_4027,N_4028,N_4029,N_4030,N_4032,N_4033,N_4034,N_4035,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4053,N_4054,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4086,N_4087,N_4089,N_4090,N_4091,N_4092,N_4094,N_4095,N_4096,N_4098,N_4099,N_4100,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4109,N_4110,N_4111,N_4112,N_4113,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4127,N_4128,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4138,N_4139,N_4141,N_4142,N_4143,N_4144,N_4145,N_4147,N_4148,N_4149,N_4150,N_4151,N_4153,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4176,N_4177,N_4178,N_4180,N_4181,N_4182,N_4183,N_4184,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4199,N_4200,N_4201,N_4202,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4211,N_4212,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4232,N_4233,N_4236,N_4238,N_4239,N_4240,N_4241,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4275,N_4277,N_4278,N_4279,N_4280,N_4284,N_4285,N_4286,N_4287,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4299,N_4301,N_4302,N_4303,N_4304,N_4305,N_4307,N_4308,N_4309,N_4312,N_4313,N_4315,N_4316,N_4318,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4336,N_4337,N_4338,N_4339,N_4340,N_4342,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4353,N_4354,N_4355,N_4357,N_4358,N_4359,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4378,N_4379,N_4380,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4391,N_4392,N_4393,N_4395,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4406,N_4407,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4418,N_4419,N_4421,N_4422,N_4423,N_4425,N_4426,N_4427,N_4430,N_4431,N_4434,N_4435,N_4436,N_4437,N_4439,N_4440,N_4441,N_4444,N_4446,N_4447,N_4449,N_4451,N_4453,N_4455,N_4456,N_4458,N_4459,N_4460,N_4462,N_4465,N_4466,N_4468,N_4469,N_4470,N_4472,N_4473,N_4474,N_4475,N_4478,N_4479,N_4480,N_4482,N_4483,N_4484,N_4485,N_4487,N_4488,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4515,N_4516,N_4518,N_4519,N_4520,N_4522,N_4523,N_4524,N_4525,N_4527,N_4528,N_4529,N_4530,N_4532,N_4533,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4543,N_4544,N_4546,N_4547,N_4548,N_4550,N_4552,N_4553,N_4554,N_4555,N_4556,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4606,N_4608,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4619,N_4620,N_4623,N_4624,N_4625,N_4626,N_4629,N_4630,N_4631,N_4633,N_4634,N_4635,N_4636,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4646,N_4647,N_4649,N_4650,N_4651,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4683,N_4687,N_4688,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4698,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4708,N_4709,N_4710,N_4711,N_4714,N_4716,N_4717,N_4718,N_4721,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4731,N_4732,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4744,N_4745,N_4746,N_4747,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4758,N_4759,N_4760,N_4761,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4781,N_4782,N_4783,N_4784,N_4785,N_4787,N_4788,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4800,N_4801,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4811,N_4812,N_4814,N_4815,N_4817,N_4819,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4836,N_4838,N_4839,N_4840,N_4842,N_4843,N_4844,N_4845,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4871,N_4872,N_4874,N_4875,N_4877,N_4879,N_4880,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4908,N_4909,N_4911,N_4912,N_4913,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4952,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4962,N_4963,N_4964,N_4965,N_4967,N_4968,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4977,N_4979,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4997,N_4998,N_4999;
nor U0 (N_0,In_367,In_280);
nor U1 (N_1,In_3,In_702);
nor U2 (N_2,In_549,In_176);
and U3 (N_3,In_246,In_46);
nor U4 (N_4,In_97,In_34);
nand U5 (N_5,In_264,In_158);
xnor U6 (N_6,In_378,In_64);
nand U7 (N_7,In_385,In_295);
nand U8 (N_8,In_533,In_372);
nor U9 (N_9,In_574,In_610);
and U10 (N_10,In_279,In_683);
xor U11 (N_11,In_735,In_149);
nand U12 (N_12,In_408,In_81);
nor U13 (N_13,In_67,In_369);
or U14 (N_14,In_336,In_698);
or U15 (N_15,In_204,In_255);
xnor U16 (N_16,In_422,In_444);
xnor U17 (N_17,In_113,In_99);
xnor U18 (N_18,In_145,In_89);
nor U19 (N_19,In_441,In_381);
nand U20 (N_20,In_712,In_0);
or U21 (N_21,In_183,In_592);
nor U22 (N_22,In_479,In_440);
xnor U23 (N_23,In_605,In_314);
and U24 (N_24,In_392,In_516);
or U25 (N_25,In_359,In_565);
nand U26 (N_26,In_497,In_687);
nand U27 (N_27,In_306,In_254);
nor U28 (N_28,In_648,In_54);
nor U29 (N_29,In_748,In_631);
nor U30 (N_30,In_288,In_73);
and U31 (N_31,In_339,In_107);
nor U32 (N_32,In_318,In_347);
nor U33 (N_33,In_351,In_507);
nor U34 (N_34,In_63,In_705);
nand U35 (N_35,In_739,In_483);
nor U36 (N_36,In_364,In_78);
or U37 (N_37,In_266,In_701);
and U38 (N_38,In_285,In_606);
nor U39 (N_39,In_40,In_162);
or U40 (N_40,In_305,In_691);
or U41 (N_41,In_404,In_12);
nor U42 (N_42,In_562,In_337);
nor U43 (N_43,In_690,In_116);
and U44 (N_44,In_414,In_538);
and U45 (N_45,In_83,In_317);
or U46 (N_46,In_172,In_212);
xor U47 (N_47,In_45,In_390);
and U48 (N_48,In_124,In_684);
or U49 (N_49,In_720,In_323);
xor U50 (N_50,In_420,In_543);
and U51 (N_51,In_44,In_341);
xor U52 (N_52,In_692,In_60);
xnor U53 (N_53,In_135,In_394);
nand U54 (N_54,In_730,In_608);
and U55 (N_55,In_510,In_48);
xor U56 (N_56,In_58,In_438);
nor U57 (N_57,In_644,In_108);
or U58 (N_58,In_519,In_56);
or U59 (N_59,In_612,In_699);
and U60 (N_60,In_348,In_437);
nor U61 (N_61,In_621,In_708);
and U62 (N_62,In_506,In_589);
and U63 (N_63,In_39,In_628);
and U64 (N_64,In_342,In_94);
and U65 (N_65,In_96,In_227);
or U66 (N_66,In_100,In_294);
nand U67 (N_67,In_627,In_356);
or U68 (N_68,In_27,In_250);
nor U69 (N_69,In_578,In_368);
xor U70 (N_70,In_586,In_402);
nor U71 (N_71,In_388,In_71);
nor U72 (N_72,In_459,In_482);
nand U73 (N_73,In_535,In_603);
and U74 (N_74,In_594,In_76);
nand U75 (N_75,In_84,In_544);
xor U76 (N_76,In_361,In_649);
nand U77 (N_77,In_273,In_238);
nand U78 (N_78,In_407,In_163);
or U79 (N_79,In_741,In_292);
xor U80 (N_80,In_171,In_6);
nand U81 (N_81,In_198,In_595);
nor U82 (N_82,In_576,In_106);
and U83 (N_83,In_480,In_241);
nand U84 (N_84,In_332,In_201);
nor U85 (N_85,In_148,In_467);
nand U86 (N_86,In_278,In_258);
nor U87 (N_87,In_453,In_47);
nand U88 (N_88,In_445,In_207);
nand U89 (N_89,In_520,In_380);
and U90 (N_90,In_680,In_512);
nand U91 (N_91,In_518,In_303);
nor U92 (N_92,In_231,In_377);
nand U93 (N_93,In_349,In_726);
nor U94 (N_94,In_736,In_251);
and U95 (N_95,In_749,In_117);
or U96 (N_96,In_617,In_308);
and U97 (N_97,In_715,In_2);
nand U98 (N_98,In_209,In_234);
xnor U99 (N_99,In_620,In_744);
xor U100 (N_100,In_25,In_421);
and U101 (N_101,In_182,In_714);
and U102 (N_102,In_276,In_706);
nor U103 (N_103,In_98,In_62);
nor U104 (N_104,In_340,In_287);
nor U105 (N_105,In_469,In_167);
nor U106 (N_106,In_443,In_307);
xnor U107 (N_107,In_366,In_740);
xor U108 (N_108,In_387,In_104);
and U109 (N_109,In_127,In_493);
nand U110 (N_110,In_464,In_524);
and U111 (N_111,In_213,In_373);
or U112 (N_112,In_661,In_43);
or U113 (N_113,In_637,In_232);
nor U114 (N_114,In_728,In_299);
and U115 (N_115,In_501,In_564);
nor U116 (N_116,In_284,In_406);
and U117 (N_117,In_395,In_600);
and U118 (N_118,In_202,In_618);
xor U119 (N_119,In_547,In_523);
nor U120 (N_120,In_442,In_707);
nand U121 (N_121,In_334,In_147);
nand U122 (N_122,In_671,In_345);
and U123 (N_123,In_10,In_325);
or U124 (N_124,In_322,In_19);
nor U125 (N_125,In_129,In_330);
and U126 (N_126,In_721,In_169);
nor U127 (N_127,In_105,In_331);
and U128 (N_128,In_33,In_537);
nor U129 (N_129,In_642,In_693);
nand U130 (N_130,In_473,In_432);
nor U131 (N_131,In_528,In_174);
and U132 (N_132,In_678,In_24);
nor U133 (N_133,In_50,In_188);
nand U134 (N_134,In_168,In_742);
or U135 (N_135,In_240,In_32);
xnor U136 (N_136,In_393,In_87);
nand U137 (N_137,In_203,In_451);
or U138 (N_138,In_7,In_666);
nand U139 (N_139,In_622,In_522);
and U140 (N_140,In_681,In_70);
nor U141 (N_141,In_585,In_546);
nand U142 (N_142,In_599,In_477);
nand U143 (N_143,In_570,In_91);
or U144 (N_144,In_180,In_624);
or U145 (N_145,In_737,In_270);
and U146 (N_146,In_181,In_677);
and U147 (N_147,In_607,In_190);
and U148 (N_148,In_685,In_256);
nor U149 (N_149,In_654,In_615);
nor U150 (N_150,In_556,In_249);
or U151 (N_151,In_418,In_553);
and U152 (N_152,In_230,In_352);
xor U153 (N_153,In_670,In_625);
and U154 (N_154,In_268,In_655);
xor U155 (N_155,In_511,In_324);
nand U156 (N_156,In_725,In_478);
and U157 (N_157,In_379,In_192);
or U158 (N_158,In_499,In_696);
nor U159 (N_159,In_311,In_426);
nand U160 (N_160,In_300,In_494);
xnor U161 (N_161,In_577,In_557);
nand U162 (N_162,In_672,In_566);
or U163 (N_163,In_738,In_614);
nand U164 (N_164,In_115,In_466);
and U165 (N_165,In_111,In_515);
nor U166 (N_166,In_312,In_132);
nor U167 (N_167,In_66,In_509);
or U168 (N_168,In_718,In_141);
nand U169 (N_169,In_686,In_85);
or U170 (N_170,In_568,In_496);
xor U171 (N_171,In_456,In_355);
xnor U172 (N_172,In_344,In_245);
and U173 (N_173,In_668,In_481);
xor U174 (N_174,In_112,In_187);
or U175 (N_175,In_102,In_650);
nor U176 (N_176,In_346,In_109);
nor U177 (N_177,In_651,In_92);
nor U178 (N_178,In_237,In_362);
nor U179 (N_179,In_659,In_123);
and U180 (N_180,In_667,In_552);
nor U181 (N_181,In_383,In_277);
nor U182 (N_182,In_601,In_598);
and U183 (N_183,In_689,In_450);
nand U184 (N_184,In_186,In_134);
nand U185 (N_185,In_52,In_271);
nand U186 (N_186,In_315,In_248);
nand U187 (N_187,In_199,In_674);
nand U188 (N_188,In_320,In_80);
or U189 (N_189,In_252,In_452);
xnor U190 (N_190,In_175,In_401);
nor U191 (N_191,In_222,In_283);
nor U192 (N_192,In_36,In_118);
nand U193 (N_193,In_210,In_139);
xnor U194 (N_194,In_590,In_643);
and U195 (N_195,In_584,In_711);
or U196 (N_196,In_413,In_461);
xor U197 (N_197,In_504,In_214);
xnor U198 (N_198,In_110,In_121);
xor U199 (N_199,In_662,In_724);
xnor U200 (N_200,In_272,In_65);
and U201 (N_201,In_136,In_28);
nor U202 (N_202,In_59,In_243);
xor U203 (N_203,In_120,In_69);
nor U204 (N_204,In_409,In_709);
xor U205 (N_205,In_42,In_211);
xnor U206 (N_206,In_173,In_150);
nor U207 (N_207,In_449,In_267);
and U208 (N_208,In_122,In_593);
xor U209 (N_209,In_242,In_688);
or U210 (N_210,In_727,In_194);
xor U211 (N_211,In_573,In_486);
nand U212 (N_212,In_425,In_17);
nor U213 (N_213,In_632,In_669);
and U214 (N_214,In_530,In_660);
nand U215 (N_215,In_154,In_428);
nor U216 (N_216,In_411,In_508);
or U217 (N_217,In_257,In_376);
xnor U218 (N_218,In_675,In_178);
and U219 (N_219,In_732,In_21);
nor U220 (N_220,In_144,In_555);
or U221 (N_221,In_695,In_218);
nor U222 (N_222,In_220,In_531);
xnor U223 (N_223,In_604,In_559);
or U224 (N_224,In_673,In_733);
and U225 (N_225,In_191,In_560);
xnor U226 (N_226,In_391,In_338);
and U227 (N_227,In_143,In_458);
nand U228 (N_228,In_462,In_572);
and U229 (N_229,In_580,In_641);
xor U230 (N_230,In_233,In_128);
or U231 (N_231,In_219,In_567);
or U232 (N_232,In_457,In_554);
nor U233 (N_233,In_472,In_485);
xor U234 (N_234,In_57,In_261);
nor U235 (N_235,In_260,In_471);
or U236 (N_236,In_263,In_639);
and U237 (N_237,In_498,In_151);
nor U238 (N_238,In_489,In_247);
or U239 (N_239,In_156,In_454);
nand U240 (N_240,In_354,In_448);
nor U241 (N_241,In_658,In_374);
and U242 (N_242,In_281,In_534);
and U243 (N_243,In_527,In_31);
nand U244 (N_244,In_88,In_229);
nor U245 (N_245,In_517,In_30);
nor U246 (N_246,In_636,In_14);
and U247 (N_247,In_446,In_638);
nand U248 (N_248,In_545,In_343);
xor U249 (N_249,In_5,In_298);
nor U250 (N_250,In_196,In_131);
xnor U251 (N_251,In_126,In_503);
and U252 (N_252,In_51,In_13);
and U253 (N_253,In_304,In_22);
xnor U254 (N_254,In_130,In_429);
or U255 (N_255,In_309,In_412);
xor U256 (N_256,In_95,In_205);
and U257 (N_257,In_114,In_646);
or U258 (N_258,In_743,In_226);
or U259 (N_259,In_403,In_396);
xor U260 (N_260,In_291,In_540);
xnor U261 (N_261,In_18,In_133);
nor U262 (N_262,In_551,In_676);
and U263 (N_263,In_236,In_184);
nand U264 (N_264,In_611,In_74);
or U265 (N_265,In_716,In_37);
xor U266 (N_266,In_189,In_137);
or U267 (N_267,In_329,In_384);
and U268 (N_268,In_79,In_206);
or U269 (N_269,In_635,In_682);
or U270 (N_270,In_370,In_244);
xor U271 (N_271,In_155,In_289);
or U272 (N_272,In_282,In_302);
and U273 (N_273,In_4,In_623);
xor U274 (N_274,In_259,In_177);
or U275 (N_275,In_613,In_587);
and U276 (N_276,In_26,In_398);
or U277 (N_277,In_399,In_571);
xor U278 (N_278,In_433,In_596);
or U279 (N_279,In_328,In_125);
nor U280 (N_280,In_93,In_274);
and U281 (N_281,In_195,In_400);
nor U282 (N_282,In_435,In_29);
xnor U283 (N_283,In_616,In_8);
nand U284 (N_284,In_694,In_217);
nor U285 (N_285,In_16,In_296);
xor U286 (N_286,In_558,In_275);
xor U287 (N_287,In_72,In_526);
or U288 (N_288,In_253,In_61);
xor U289 (N_289,In_645,In_363);
nor U290 (N_290,In_164,In_626);
and U291 (N_291,In_389,In_729);
xor U292 (N_292,In_719,In_474);
nand U293 (N_293,In_23,In_439);
nand U294 (N_294,In_165,In_542);
xor U295 (N_295,In_665,In_375);
nor U296 (N_296,In_1,In_321);
nand U297 (N_297,In_539,In_200);
xor U298 (N_298,In_140,In_460);
and U299 (N_299,In_333,In_713);
or U300 (N_300,In_161,In_488);
and U301 (N_301,In_652,In_166);
nand U302 (N_302,In_262,In_633);
and U303 (N_303,In_316,In_228);
and U304 (N_304,In_653,In_313);
nor U305 (N_305,In_463,In_717);
nor U306 (N_306,In_53,In_582);
and U307 (N_307,In_157,In_476);
xnor U308 (N_308,In_215,In_82);
xor U309 (N_309,In_77,In_704);
nand U310 (N_310,In_360,In_185);
xor U311 (N_311,In_583,In_495);
xnor U312 (N_312,In_423,In_216);
nor U313 (N_313,In_224,In_427);
nor U314 (N_314,In_647,In_75);
and U315 (N_315,In_548,In_529);
nor U316 (N_316,In_170,In_357);
or U317 (N_317,In_101,In_747);
xnor U318 (N_318,In_301,In_710);
or U319 (N_319,In_436,In_416);
nor U320 (N_320,In_146,In_563);
and U321 (N_321,In_492,In_629);
and U322 (N_322,In_9,In_86);
and U323 (N_323,In_327,In_11);
nor U324 (N_324,In_397,In_38);
xor U325 (N_325,In_41,In_269);
xor U326 (N_326,In_265,In_335);
and U327 (N_327,In_597,In_634);
nand U328 (N_328,In_697,In_159);
nor U329 (N_329,In_700,In_221);
or U330 (N_330,In_197,In_468);
and U331 (N_331,In_703,In_470);
and U332 (N_332,In_319,In_430);
and U333 (N_333,In_663,In_208);
and U334 (N_334,In_521,In_179);
nand U335 (N_335,In_293,In_591);
or U336 (N_336,In_290,In_455);
nor U337 (N_337,In_575,In_569);
xnor U338 (N_338,In_550,In_664);
xnor U339 (N_339,In_505,In_500);
nor U340 (N_340,In_415,In_417);
or U341 (N_341,In_286,In_579);
nor U342 (N_342,In_119,In_225);
or U343 (N_343,In_90,In_640);
nor U344 (N_344,In_353,In_386);
and U345 (N_345,In_193,In_49);
xor U346 (N_346,In_536,In_630);
xnor U347 (N_347,In_223,In_152);
and U348 (N_348,In_487,In_138);
xor U349 (N_349,In_465,In_310);
or U350 (N_350,In_358,In_410);
xnor U351 (N_351,In_722,In_55);
and U352 (N_352,In_502,In_541);
or U353 (N_353,In_514,In_447);
or U354 (N_354,In_525,In_491);
or U355 (N_355,In_513,In_588);
nor U356 (N_356,In_239,In_297);
or U357 (N_357,In_20,In_532);
xor U358 (N_358,In_723,In_490);
nand U359 (N_359,In_365,In_68);
nor U360 (N_360,In_15,In_160);
nor U361 (N_361,In_424,In_561);
xnor U362 (N_362,In_609,In_431);
xnor U363 (N_363,In_103,In_581);
nor U364 (N_364,In_475,In_731);
and U365 (N_365,In_434,In_382);
nor U366 (N_366,In_734,In_602);
nor U367 (N_367,In_484,In_142);
xor U368 (N_368,In_419,In_657);
nor U369 (N_369,In_235,In_35);
xor U370 (N_370,In_619,In_405);
nand U371 (N_371,In_745,In_679);
or U372 (N_372,In_153,In_350);
and U373 (N_373,In_746,In_326);
nand U374 (N_374,In_371,In_656);
or U375 (N_375,In_113,In_131);
and U376 (N_376,In_683,In_670);
and U377 (N_377,In_293,In_715);
nor U378 (N_378,In_686,In_423);
and U379 (N_379,In_24,In_311);
nor U380 (N_380,In_322,In_472);
nand U381 (N_381,In_733,In_556);
nand U382 (N_382,In_508,In_179);
xnor U383 (N_383,In_138,In_155);
or U384 (N_384,In_598,In_744);
nand U385 (N_385,In_176,In_731);
or U386 (N_386,In_596,In_525);
and U387 (N_387,In_69,In_539);
or U388 (N_388,In_87,In_168);
and U389 (N_389,In_480,In_528);
or U390 (N_390,In_383,In_560);
nor U391 (N_391,In_188,In_200);
nand U392 (N_392,In_659,In_418);
nand U393 (N_393,In_343,In_597);
xnor U394 (N_394,In_624,In_188);
nand U395 (N_395,In_460,In_695);
xor U396 (N_396,In_245,In_1);
or U397 (N_397,In_702,In_89);
xor U398 (N_398,In_282,In_725);
nor U399 (N_399,In_456,In_17);
or U400 (N_400,In_345,In_584);
xnor U401 (N_401,In_211,In_264);
xor U402 (N_402,In_83,In_4);
nand U403 (N_403,In_186,In_129);
xor U404 (N_404,In_405,In_628);
xnor U405 (N_405,In_529,In_510);
or U406 (N_406,In_406,In_729);
xnor U407 (N_407,In_514,In_670);
and U408 (N_408,In_189,In_308);
and U409 (N_409,In_509,In_341);
nand U410 (N_410,In_207,In_374);
or U411 (N_411,In_713,In_102);
nand U412 (N_412,In_391,In_633);
nand U413 (N_413,In_451,In_47);
and U414 (N_414,In_172,In_386);
nor U415 (N_415,In_507,In_296);
or U416 (N_416,In_572,In_727);
nor U417 (N_417,In_541,In_503);
nand U418 (N_418,In_461,In_625);
or U419 (N_419,In_604,In_306);
xor U420 (N_420,In_514,In_164);
nand U421 (N_421,In_162,In_415);
nand U422 (N_422,In_507,In_526);
and U423 (N_423,In_9,In_285);
and U424 (N_424,In_724,In_616);
nand U425 (N_425,In_26,In_628);
and U426 (N_426,In_742,In_167);
or U427 (N_427,In_227,In_554);
and U428 (N_428,In_479,In_320);
and U429 (N_429,In_688,In_267);
nand U430 (N_430,In_641,In_73);
nand U431 (N_431,In_132,In_454);
or U432 (N_432,In_473,In_447);
nand U433 (N_433,In_706,In_631);
and U434 (N_434,In_159,In_465);
and U435 (N_435,In_538,In_85);
nand U436 (N_436,In_112,In_583);
nand U437 (N_437,In_481,In_244);
and U438 (N_438,In_614,In_711);
nand U439 (N_439,In_347,In_196);
nor U440 (N_440,In_654,In_421);
or U441 (N_441,In_628,In_183);
and U442 (N_442,In_96,In_223);
and U443 (N_443,In_175,In_246);
nor U444 (N_444,In_159,In_203);
xnor U445 (N_445,In_319,In_46);
nor U446 (N_446,In_570,In_666);
nor U447 (N_447,In_240,In_582);
nor U448 (N_448,In_615,In_626);
nor U449 (N_449,In_124,In_566);
nand U450 (N_450,In_122,In_645);
xnor U451 (N_451,In_598,In_409);
xor U452 (N_452,In_122,In_134);
nor U453 (N_453,In_236,In_144);
and U454 (N_454,In_9,In_437);
xor U455 (N_455,In_376,In_340);
nor U456 (N_456,In_389,In_661);
or U457 (N_457,In_534,In_118);
and U458 (N_458,In_267,In_536);
xnor U459 (N_459,In_155,In_616);
nand U460 (N_460,In_385,In_733);
nand U461 (N_461,In_459,In_367);
or U462 (N_462,In_553,In_129);
nand U463 (N_463,In_552,In_656);
and U464 (N_464,In_440,In_252);
nor U465 (N_465,In_479,In_347);
nor U466 (N_466,In_193,In_433);
xor U467 (N_467,In_625,In_521);
and U468 (N_468,In_320,In_373);
xnor U469 (N_469,In_745,In_742);
nand U470 (N_470,In_343,In_149);
nand U471 (N_471,In_311,In_395);
nor U472 (N_472,In_477,In_299);
xnor U473 (N_473,In_263,In_391);
nand U474 (N_474,In_539,In_373);
nand U475 (N_475,In_66,In_139);
and U476 (N_476,In_91,In_646);
nand U477 (N_477,In_81,In_79);
and U478 (N_478,In_4,In_610);
and U479 (N_479,In_432,In_451);
and U480 (N_480,In_198,In_509);
nor U481 (N_481,In_654,In_454);
nor U482 (N_482,In_669,In_151);
nor U483 (N_483,In_701,In_106);
xnor U484 (N_484,In_689,In_77);
xor U485 (N_485,In_3,In_109);
and U486 (N_486,In_427,In_599);
nor U487 (N_487,In_482,In_269);
nand U488 (N_488,In_223,In_613);
nor U489 (N_489,In_708,In_2);
nor U490 (N_490,In_604,In_635);
nand U491 (N_491,In_298,In_704);
nor U492 (N_492,In_453,In_494);
xnor U493 (N_493,In_399,In_248);
nand U494 (N_494,In_30,In_644);
nand U495 (N_495,In_448,In_310);
nand U496 (N_496,In_715,In_343);
nor U497 (N_497,In_427,In_731);
or U498 (N_498,In_348,In_426);
and U499 (N_499,In_385,In_405);
or U500 (N_500,In_28,In_51);
xor U501 (N_501,In_71,In_340);
xnor U502 (N_502,In_470,In_660);
xnor U503 (N_503,In_346,In_115);
or U504 (N_504,In_21,In_727);
nand U505 (N_505,In_295,In_338);
nand U506 (N_506,In_698,In_718);
and U507 (N_507,In_638,In_533);
nand U508 (N_508,In_9,In_639);
or U509 (N_509,In_397,In_710);
and U510 (N_510,In_235,In_612);
nand U511 (N_511,In_474,In_576);
nor U512 (N_512,In_393,In_217);
and U513 (N_513,In_325,In_462);
nand U514 (N_514,In_642,In_353);
and U515 (N_515,In_9,In_210);
nor U516 (N_516,In_616,In_673);
and U517 (N_517,In_355,In_122);
xnor U518 (N_518,In_676,In_267);
nand U519 (N_519,In_531,In_452);
xnor U520 (N_520,In_285,In_660);
nand U521 (N_521,In_117,In_609);
or U522 (N_522,In_666,In_684);
and U523 (N_523,In_301,In_58);
nand U524 (N_524,In_411,In_581);
and U525 (N_525,In_556,In_623);
nand U526 (N_526,In_342,In_386);
or U527 (N_527,In_305,In_496);
or U528 (N_528,In_225,In_648);
nor U529 (N_529,In_69,In_487);
nor U530 (N_530,In_33,In_332);
and U531 (N_531,In_305,In_88);
xnor U532 (N_532,In_413,In_611);
xnor U533 (N_533,In_416,In_66);
or U534 (N_534,In_478,In_38);
and U535 (N_535,In_89,In_32);
xnor U536 (N_536,In_317,In_74);
nor U537 (N_537,In_707,In_408);
nor U538 (N_538,In_151,In_187);
nand U539 (N_539,In_665,In_284);
nor U540 (N_540,In_39,In_518);
and U541 (N_541,In_121,In_733);
nor U542 (N_542,In_358,In_395);
nor U543 (N_543,In_546,In_381);
nand U544 (N_544,In_257,In_205);
xnor U545 (N_545,In_122,In_369);
or U546 (N_546,In_438,In_730);
and U547 (N_547,In_493,In_651);
xor U548 (N_548,In_346,In_212);
or U549 (N_549,In_388,In_204);
nand U550 (N_550,In_438,In_447);
xnor U551 (N_551,In_538,In_109);
nor U552 (N_552,In_640,In_18);
or U553 (N_553,In_224,In_111);
nor U554 (N_554,In_108,In_24);
xor U555 (N_555,In_403,In_87);
and U556 (N_556,In_240,In_522);
xor U557 (N_557,In_406,In_484);
nor U558 (N_558,In_161,In_635);
and U559 (N_559,In_53,In_130);
nand U560 (N_560,In_591,In_719);
or U561 (N_561,In_513,In_457);
or U562 (N_562,In_340,In_104);
nand U563 (N_563,In_692,In_572);
nor U564 (N_564,In_360,In_626);
or U565 (N_565,In_79,In_582);
or U566 (N_566,In_313,In_613);
and U567 (N_567,In_124,In_648);
or U568 (N_568,In_274,In_498);
nand U569 (N_569,In_705,In_618);
or U570 (N_570,In_335,In_738);
nor U571 (N_571,In_162,In_303);
nand U572 (N_572,In_295,In_391);
or U573 (N_573,In_195,In_182);
nor U574 (N_574,In_660,In_526);
or U575 (N_575,In_746,In_501);
or U576 (N_576,In_76,In_195);
nand U577 (N_577,In_272,In_562);
nand U578 (N_578,In_505,In_28);
or U579 (N_579,In_195,In_582);
and U580 (N_580,In_41,In_602);
xnor U581 (N_581,In_48,In_25);
xor U582 (N_582,In_329,In_421);
nand U583 (N_583,In_555,In_6);
xor U584 (N_584,In_164,In_527);
or U585 (N_585,In_640,In_212);
xnor U586 (N_586,In_601,In_346);
nor U587 (N_587,In_505,In_393);
and U588 (N_588,In_86,In_355);
xnor U589 (N_589,In_378,In_676);
nand U590 (N_590,In_378,In_649);
and U591 (N_591,In_51,In_351);
nor U592 (N_592,In_443,In_721);
xnor U593 (N_593,In_445,In_189);
xnor U594 (N_594,In_312,In_452);
nor U595 (N_595,In_624,In_362);
nand U596 (N_596,In_661,In_624);
nor U597 (N_597,In_457,In_575);
nor U598 (N_598,In_468,In_316);
and U599 (N_599,In_421,In_248);
or U600 (N_600,In_599,In_402);
and U601 (N_601,In_250,In_708);
and U602 (N_602,In_62,In_267);
nor U603 (N_603,In_235,In_88);
and U604 (N_604,In_522,In_70);
nor U605 (N_605,In_433,In_443);
nand U606 (N_606,In_99,In_611);
or U607 (N_607,In_431,In_235);
xnor U608 (N_608,In_77,In_475);
xor U609 (N_609,In_480,In_562);
nand U610 (N_610,In_719,In_437);
nor U611 (N_611,In_147,In_730);
xnor U612 (N_612,In_14,In_312);
or U613 (N_613,In_27,In_424);
nor U614 (N_614,In_303,In_641);
nand U615 (N_615,In_576,In_519);
nand U616 (N_616,In_502,In_425);
nand U617 (N_617,In_149,In_355);
xor U618 (N_618,In_220,In_86);
or U619 (N_619,In_351,In_243);
xor U620 (N_620,In_84,In_735);
nand U621 (N_621,In_728,In_331);
xnor U622 (N_622,In_644,In_329);
and U623 (N_623,In_551,In_471);
nand U624 (N_624,In_713,In_498);
and U625 (N_625,In_140,In_224);
or U626 (N_626,In_331,In_673);
or U627 (N_627,In_55,In_678);
and U628 (N_628,In_566,In_517);
and U629 (N_629,In_28,In_241);
nand U630 (N_630,In_596,In_182);
xor U631 (N_631,In_392,In_287);
and U632 (N_632,In_672,In_736);
or U633 (N_633,In_402,In_189);
and U634 (N_634,In_490,In_346);
nor U635 (N_635,In_749,In_738);
and U636 (N_636,In_524,In_287);
or U637 (N_637,In_629,In_514);
nand U638 (N_638,In_398,In_358);
or U639 (N_639,In_216,In_329);
nand U640 (N_640,In_322,In_35);
nand U641 (N_641,In_238,In_175);
xnor U642 (N_642,In_190,In_653);
and U643 (N_643,In_479,In_577);
nor U644 (N_644,In_649,In_514);
and U645 (N_645,In_542,In_682);
nor U646 (N_646,In_312,In_392);
nor U647 (N_647,In_532,In_356);
nor U648 (N_648,In_740,In_5);
xor U649 (N_649,In_578,In_546);
nand U650 (N_650,In_125,In_226);
nor U651 (N_651,In_689,In_260);
or U652 (N_652,In_615,In_214);
or U653 (N_653,In_563,In_455);
xnor U654 (N_654,In_246,In_326);
nand U655 (N_655,In_619,In_71);
nand U656 (N_656,In_404,In_268);
nor U657 (N_657,In_199,In_326);
and U658 (N_658,In_400,In_529);
nand U659 (N_659,In_143,In_499);
nand U660 (N_660,In_387,In_63);
nand U661 (N_661,In_375,In_361);
nand U662 (N_662,In_3,In_97);
nor U663 (N_663,In_25,In_680);
or U664 (N_664,In_547,In_686);
or U665 (N_665,In_565,In_260);
and U666 (N_666,In_265,In_721);
xor U667 (N_667,In_229,In_20);
and U668 (N_668,In_598,In_486);
xor U669 (N_669,In_248,In_37);
nor U670 (N_670,In_308,In_508);
nand U671 (N_671,In_315,In_513);
and U672 (N_672,In_531,In_604);
or U673 (N_673,In_597,In_355);
nor U674 (N_674,In_547,In_457);
and U675 (N_675,In_308,In_43);
xor U676 (N_676,In_518,In_631);
and U677 (N_677,In_566,In_623);
nand U678 (N_678,In_521,In_257);
nand U679 (N_679,In_93,In_276);
xor U680 (N_680,In_1,In_247);
and U681 (N_681,In_499,In_722);
nor U682 (N_682,In_151,In_723);
xor U683 (N_683,In_381,In_333);
nand U684 (N_684,In_735,In_300);
and U685 (N_685,In_503,In_543);
and U686 (N_686,In_472,In_621);
nor U687 (N_687,In_237,In_443);
or U688 (N_688,In_31,In_177);
nor U689 (N_689,In_236,In_500);
nor U690 (N_690,In_740,In_95);
nand U691 (N_691,In_301,In_688);
or U692 (N_692,In_352,In_73);
xor U693 (N_693,In_343,In_1);
and U694 (N_694,In_731,In_264);
nand U695 (N_695,In_276,In_322);
xnor U696 (N_696,In_558,In_421);
or U697 (N_697,In_521,In_723);
and U698 (N_698,In_63,In_579);
xnor U699 (N_699,In_691,In_310);
nand U700 (N_700,In_318,In_10);
and U701 (N_701,In_314,In_439);
nor U702 (N_702,In_108,In_8);
and U703 (N_703,In_382,In_300);
and U704 (N_704,In_215,In_219);
nand U705 (N_705,In_385,In_62);
or U706 (N_706,In_617,In_382);
xnor U707 (N_707,In_742,In_77);
nand U708 (N_708,In_691,In_498);
or U709 (N_709,In_704,In_578);
or U710 (N_710,In_330,In_84);
nor U711 (N_711,In_354,In_374);
and U712 (N_712,In_604,In_337);
or U713 (N_713,In_344,In_729);
xnor U714 (N_714,In_727,In_211);
or U715 (N_715,In_540,In_249);
xor U716 (N_716,In_708,In_591);
and U717 (N_717,In_412,In_261);
nor U718 (N_718,In_59,In_576);
nor U719 (N_719,In_680,In_152);
and U720 (N_720,In_319,In_611);
or U721 (N_721,In_612,In_179);
or U722 (N_722,In_475,In_88);
xor U723 (N_723,In_75,In_229);
nand U724 (N_724,In_123,In_248);
and U725 (N_725,In_682,In_246);
and U726 (N_726,In_444,In_215);
and U727 (N_727,In_490,In_272);
nand U728 (N_728,In_473,In_18);
or U729 (N_729,In_308,In_218);
nand U730 (N_730,In_666,In_423);
nor U731 (N_731,In_161,In_462);
nand U732 (N_732,In_263,In_582);
nor U733 (N_733,In_446,In_82);
and U734 (N_734,In_407,In_347);
or U735 (N_735,In_577,In_414);
xnor U736 (N_736,In_352,In_242);
xnor U737 (N_737,In_631,In_607);
and U738 (N_738,In_143,In_356);
xnor U739 (N_739,In_361,In_430);
xor U740 (N_740,In_700,In_600);
and U741 (N_741,In_267,In_283);
or U742 (N_742,In_220,In_594);
nor U743 (N_743,In_613,In_285);
nor U744 (N_744,In_200,In_126);
xnor U745 (N_745,In_707,In_169);
and U746 (N_746,In_20,In_92);
nand U747 (N_747,In_154,In_326);
or U748 (N_748,In_661,In_524);
or U749 (N_749,In_216,In_610);
nor U750 (N_750,In_588,In_346);
and U751 (N_751,In_108,In_133);
and U752 (N_752,In_570,In_28);
and U753 (N_753,In_96,In_502);
nor U754 (N_754,In_363,In_75);
nor U755 (N_755,In_185,In_100);
or U756 (N_756,In_110,In_365);
nand U757 (N_757,In_555,In_127);
and U758 (N_758,In_409,In_233);
nand U759 (N_759,In_126,In_21);
xnor U760 (N_760,In_289,In_527);
or U761 (N_761,In_266,In_333);
or U762 (N_762,In_103,In_410);
or U763 (N_763,In_296,In_30);
and U764 (N_764,In_492,In_695);
xor U765 (N_765,In_743,In_209);
or U766 (N_766,In_517,In_447);
and U767 (N_767,In_292,In_592);
or U768 (N_768,In_468,In_95);
and U769 (N_769,In_379,In_572);
xnor U770 (N_770,In_732,In_726);
and U771 (N_771,In_381,In_345);
xnor U772 (N_772,In_63,In_196);
xor U773 (N_773,In_395,In_570);
nand U774 (N_774,In_251,In_30);
nand U775 (N_775,In_83,In_61);
and U776 (N_776,In_346,In_183);
nor U777 (N_777,In_677,In_618);
nor U778 (N_778,In_218,In_305);
and U779 (N_779,In_76,In_276);
nand U780 (N_780,In_725,In_483);
and U781 (N_781,In_355,In_694);
nor U782 (N_782,In_486,In_364);
and U783 (N_783,In_138,In_245);
nand U784 (N_784,In_7,In_274);
nor U785 (N_785,In_79,In_275);
nand U786 (N_786,In_572,In_504);
or U787 (N_787,In_661,In_26);
and U788 (N_788,In_53,In_33);
nand U789 (N_789,In_651,In_174);
xnor U790 (N_790,In_178,In_538);
nand U791 (N_791,In_153,In_473);
nor U792 (N_792,In_399,In_658);
or U793 (N_793,In_677,In_565);
nor U794 (N_794,In_672,In_32);
nor U795 (N_795,In_563,In_515);
or U796 (N_796,In_296,In_428);
and U797 (N_797,In_566,In_579);
or U798 (N_798,In_534,In_265);
or U799 (N_799,In_591,In_244);
nor U800 (N_800,In_620,In_339);
xnor U801 (N_801,In_728,In_21);
xnor U802 (N_802,In_544,In_4);
nor U803 (N_803,In_279,In_203);
or U804 (N_804,In_99,In_654);
nand U805 (N_805,In_221,In_714);
nor U806 (N_806,In_632,In_297);
nor U807 (N_807,In_681,In_7);
or U808 (N_808,In_76,In_706);
nand U809 (N_809,In_43,In_564);
and U810 (N_810,In_63,In_508);
xor U811 (N_811,In_685,In_679);
nand U812 (N_812,In_385,In_510);
or U813 (N_813,In_655,In_664);
xnor U814 (N_814,In_581,In_111);
xor U815 (N_815,In_202,In_507);
xor U816 (N_816,In_707,In_607);
and U817 (N_817,In_602,In_238);
and U818 (N_818,In_76,In_692);
nor U819 (N_819,In_238,In_336);
nand U820 (N_820,In_197,In_113);
nor U821 (N_821,In_622,In_743);
nor U822 (N_822,In_747,In_113);
nor U823 (N_823,In_86,In_127);
nor U824 (N_824,In_38,In_47);
nor U825 (N_825,In_108,In_136);
and U826 (N_826,In_576,In_161);
nand U827 (N_827,In_692,In_125);
and U828 (N_828,In_484,In_502);
nor U829 (N_829,In_1,In_381);
nor U830 (N_830,In_160,In_473);
xnor U831 (N_831,In_275,In_200);
or U832 (N_832,In_23,In_387);
xor U833 (N_833,In_329,In_643);
or U834 (N_834,In_313,In_80);
nand U835 (N_835,In_329,In_64);
nand U836 (N_836,In_459,In_610);
xnor U837 (N_837,In_391,In_57);
or U838 (N_838,In_308,In_72);
nand U839 (N_839,In_722,In_230);
nor U840 (N_840,In_371,In_226);
or U841 (N_841,In_683,In_128);
or U842 (N_842,In_368,In_628);
nor U843 (N_843,In_311,In_149);
and U844 (N_844,In_82,In_707);
nor U845 (N_845,In_472,In_204);
and U846 (N_846,In_467,In_506);
nor U847 (N_847,In_304,In_324);
nor U848 (N_848,In_51,In_395);
xor U849 (N_849,In_91,In_46);
nor U850 (N_850,In_320,In_619);
and U851 (N_851,In_198,In_497);
xnor U852 (N_852,In_682,In_461);
nor U853 (N_853,In_659,In_485);
nor U854 (N_854,In_240,In_619);
and U855 (N_855,In_334,In_717);
or U856 (N_856,In_192,In_666);
xnor U857 (N_857,In_83,In_150);
or U858 (N_858,In_668,In_421);
xor U859 (N_859,In_248,In_539);
or U860 (N_860,In_131,In_115);
nor U861 (N_861,In_513,In_352);
nor U862 (N_862,In_80,In_643);
xor U863 (N_863,In_242,In_710);
nand U864 (N_864,In_478,In_678);
and U865 (N_865,In_699,In_326);
or U866 (N_866,In_293,In_371);
nand U867 (N_867,In_61,In_273);
nor U868 (N_868,In_593,In_443);
and U869 (N_869,In_530,In_141);
and U870 (N_870,In_6,In_679);
or U871 (N_871,In_598,In_31);
and U872 (N_872,In_207,In_18);
nand U873 (N_873,In_679,In_154);
xnor U874 (N_874,In_689,In_384);
xor U875 (N_875,In_657,In_206);
nor U876 (N_876,In_566,In_721);
and U877 (N_877,In_310,In_61);
nor U878 (N_878,In_207,In_162);
nand U879 (N_879,In_708,In_392);
and U880 (N_880,In_6,In_259);
nor U881 (N_881,In_93,In_471);
nand U882 (N_882,In_198,In_661);
nand U883 (N_883,In_529,In_711);
xor U884 (N_884,In_128,In_584);
nor U885 (N_885,In_402,In_244);
xor U886 (N_886,In_51,In_248);
xnor U887 (N_887,In_112,In_596);
and U888 (N_888,In_462,In_375);
nor U889 (N_889,In_542,In_37);
or U890 (N_890,In_520,In_591);
nand U891 (N_891,In_210,In_333);
nor U892 (N_892,In_565,In_712);
xor U893 (N_893,In_440,In_396);
xnor U894 (N_894,In_444,In_564);
xor U895 (N_895,In_41,In_64);
or U896 (N_896,In_696,In_446);
nor U897 (N_897,In_522,In_709);
nor U898 (N_898,In_469,In_423);
and U899 (N_899,In_413,In_671);
or U900 (N_900,In_495,In_382);
or U901 (N_901,In_747,In_228);
and U902 (N_902,In_439,In_159);
nor U903 (N_903,In_31,In_136);
or U904 (N_904,In_142,In_598);
nand U905 (N_905,In_720,In_138);
and U906 (N_906,In_244,In_478);
nor U907 (N_907,In_397,In_381);
or U908 (N_908,In_708,In_37);
nand U909 (N_909,In_698,In_533);
or U910 (N_910,In_743,In_619);
nor U911 (N_911,In_466,In_299);
and U912 (N_912,In_120,In_123);
xor U913 (N_913,In_473,In_61);
or U914 (N_914,In_565,In_566);
nand U915 (N_915,In_677,In_104);
xor U916 (N_916,In_93,In_651);
xnor U917 (N_917,In_531,In_274);
nand U918 (N_918,In_163,In_521);
or U919 (N_919,In_634,In_22);
or U920 (N_920,In_240,In_478);
or U921 (N_921,In_398,In_428);
nand U922 (N_922,In_372,In_609);
and U923 (N_923,In_333,In_487);
xnor U924 (N_924,In_402,In_356);
nand U925 (N_925,In_134,In_615);
or U926 (N_926,In_471,In_277);
and U927 (N_927,In_351,In_216);
xor U928 (N_928,In_80,In_670);
nand U929 (N_929,In_392,In_492);
nand U930 (N_930,In_355,In_243);
xnor U931 (N_931,In_253,In_114);
nand U932 (N_932,In_99,In_746);
or U933 (N_933,In_684,In_354);
nor U934 (N_934,In_306,In_481);
nor U935 (N_935,In_199,In_85);
nor U936 (N_936,In_314,In_173);
and U937 (N_937,In_104,In_193);
or U938 (N_938,In_597,In_636);
nor U939 (N_939,In_66,In_332);
nor U940 (N_940,In_511,In_188);
nand U941 (N_941,In_570,In_189);
or U942 (N_942,In_619,In_175);
xor U943 (N_943,In_290,In_687);
xnor U944 (N_944,In_428,In_588);
nor U945 (N_945,In_423,In_413);
xnor U946 (N_946,In_662,In_444);
nand U947 (N_947,In_27,In_565);
nor U948 (N_948,In_105,In_521);
xnor U949 (N_949,In_499,In_537);
nand U950 (N_950,In_684,In_735);
or U951 (N_951,In_107,In_666);
nand U952 (N_952,In_739,In_43);
and U953 (N_953,In_482,In_7);
nor U954 (N_954,In_408,In_370);
nor U955 (N_955,In_12,In_530);
and U956 (N_956,In_124,In_533);
xnor U957 (N_957,In_65,In_239);
xnor U958 (N_958,In_717,In_13);
nand U959 (N_959,In_16,In_497);
nor U960 (N_960,In_422,In_477);
nand U961 (N_961,In_505,In_206);
and U962 (N_962,In_561,In_392);
and U963 (N_963,In_523,In_379);
xor U964 (N_964,In_710,In_123);
xor U965 (N_965,In_456,In_228);
or U966 (N_966,In_231,In_192);
nand U967 (N_967,In_583,In_630);
nand U968 (N_968,In_559,In_534);
and U969 (N_969,In_512,In_458);
xnor U970 (N_970,In_316,In_561);
xnor U971 (N_971,In_426,In_433);
nor U972 (N_972,In_576,In_434);
nand U973 (N_973,In_391,In_749);
and U974 (N_974,In_302,In_332);
nor U975 (N_975,In_47,In_325);
nor U976 (N_976,In_12,In_343);
xor U977 (N_977,In_249,In_431);
nor U978 (N_978,In_203,In_183);
and U979 (N_979,In_732,In_728);
nand U980 (N_980,In_70,In_257);
and U981 (N_981,In_583,In_702);
nor U982 (N_982,In_551,In_112);
nand U983 (N_983,In_545,In_342);
or U984 (N_984,In_63,In_665);
nand U985 (N_985,In_560,In_318);
xor U986 (N_986,In_379,In_153);
nor U987 (N_987,In_585,In_125);
and U988 (N_988,In_531,In_448);
nor U989 (N_989,In_707,In_733);
or U990 (N_990,In_443,In_38);
nand U991 (N_991,In_346,In_221);
and U992 (N_992,In_58,In_498);
xor U993 (N_993,In_596,In_214);
nor U994 (N_994,In_566,In_335);
nand U995 (N_995,In_5,In_605);
nor U996 (N_996,In_707,In_91);
nor U997 (N_997,In_311,In_369);
xnor U998 (N_998,In_635,In_689);
nand U999 (N_999,In_274,In_655);
nor U1000 (N_1000,In_78,In_194);
or U1001 (N_1001,In_736,In_216);
nand U1002 (N_1002,In_736,In_282);
xnor U1003 (N_1003,In_506,In_470);
nand U1004 (N_1004,In_649,In_448);
nor U1005 (N_1005,In_507,In_638);
nor U1006 (N_1006,In_412,In_580);
xor U1007 (N_1007,In_698,In_737);
nor U1008 (N_1008,In_625,In_471);
nand U1009 (N_1009,In_376,In_239);
and U1010 (N_1010,In_478,In_234);
or U1011 (N_1011,In_147,In_296);
or U1012 (N_1012,In_169,In_233);
and U1013 (N_1013,In_66,In_609);
nand U1014 (N_1014,In_747,In_334);
or U1015 (N_1015,In_372,In_143);
nor U1016 (N_1016,In_636,In_612);
and U1017 (N_1017,In_50,In_413);
and U1018 (N_1018,In_88,In_158);
or U1019 (N_1019,In_740,In_149);
xor U1020 (N_1020,In_693,In_32);
or U1021 (N_1021,In_709,In_549);
xor U1022 (N_1022,In_291,In_370);
xnor U1023 (N_1023,In_118,In_711);
xor U1024 (N_1024,In_438,In_41);
or U1025 (N_1025,In_549,In_744);
nand U1026 (N_1026,In_122,In_491);
or U1027 (N_1027,In_123,In_379);
and U1028 (N_1028,In_635,In_463);
xor U1029 (N_1029,In_406,In_91);
nor U1030 (N_1030,In_211,In_240);
xnor U1031 (N_1031,In_424,In_673);
nor U1032 (N_1032,In_440,In_520);
xnor U1033 (N_1033,In_89,In_705);
and U1034 (N_1034,In_322,In_520);
or U1035 (N_1035,In_447,In_464);
nor U1036 (N_1036,In_119,In_493);
and U1037 (N_1037,In_662,In_664);
nand U1038 (N_1038,In_267,In_457);
nand U1039 (N_1039,In_436,In_710);
nor U1040 (N_1040,In_265,In_526);
nand U1041 (N_1041,In_341,In_725);
or U1042 (N_1042,In_605,In_76);
xor U1043 (N_1043,In_534,In_486);
or U1044 (N_1044,In_248,In_198);
and U1045 (N_1045,In_445,In_64);
nor U1046 (N_1046,In_732,In_423);
xor U1047 (N_1047,In_66,In_67);
xor U1048 (N_1048,In_353,In_693);
nor U1049 (N_1049,In_675,In_243);
or U1050 (N_1050,In_195,In_427);
xor U1051 (N_1051,In_42,In_631);
nand U1052 (N_1052,In_585,In_447);
and U1053 (N_1053,In_482,In_69);
nand U1054 (N_1054,In_472,In_341);
and U1055 (N_1055,In_633,In_477);
xor U1056 (N_1056,In_234,In_107);
and U1057 (N_1057,In_209,In_190);
xnor U1058 (N_1058,In_503,In_364);
nor U1059 (N_1059,In_167,In_237);
and U1060 (N_1060,In_524,In_610);
nand U1061 (N_1061,In_628,In_613);
xnor U1062 (N_1062,In_44,In_15);
nor U1063 (N_1063,In_545,In_186);
nand U1064 (N_1064,In_661,In_302);
and U1065 (N_1065,In_150,In_676);
or U1066 (N_1066,In_13,In_120);
or U1067 (N_1067,In_268,In_146);
or U1068 (N_1068,In_618,In_52);
or U1069 (N_1069,In_296,In_591);
or U1070 (N_1070,In_259,In_309);
nand U1071 (N_1071,In_247,In_569);
nor U1072 (N_1072,In_218,In_666);
and U1073 (N_1073,In_340,In_590);
or U1074 (N_1074,In_433,In_12);
nor U1075 (N_1075,In_505,In_601);
and U1076 (N_1076,In_257,In_22);
nor U1077 (N_1077,In_381,In_290);
and U1078 (N_1078,In_526,In_173);
nor U1079 (N_1079,In_2,In_742);
and U1080 (N_1080,In_277,In_473);
nor U1081 (N_1081,In_591,In_340);
xor U1082 (N_1082,In_42,In_28);
or U1083 (N_1083,In_622,In_31);
xnor U1084 (N_1084,In_84,In_702);
nor U1085 (N_1085,In_630,In_270);
and U1086 (N_1086,In_366,In_135);
xnor U1087 (N_1087,In_60,In_342);
nor U1088 (N_1088,In_27,In_120);
and U1089 (N_1089,In_280,In_738);
and U1090 (N_1090,In_29,In_57);
nor U1091 (N_1091,In_258,In_442);
and U1092 (N_1092,In_166,In_244);
xnor U1093 (N_1093,In_694,In_583);
nor U1094 (N_1094,In_543,In_276);
or U1095 (N_1095,In_525,In_114);
and U1096 (N_1096,In_669,In_523);
xnor U1097 (N_1097,In_135,In_20);
nor U1098 (N_1098,In_86,In_493);
nand U1099 (N_1099,In_329,In_703);
nand U1100 (N_1100,In_153,In_195);
nor U1101 (N_1101,In_139,In_22);
nand U1102 (N_1102,In_110,In_223);
nand U1103 (N_1103,In_52,In_296);
or U1104 (N_1104,In_491,In_426);
and U1105 (N_1105,In_204,In_420);
nand U1106 (N_1106,In_292,In_508);
nor U1107 (N_1107,In_103,In_0);
or U1108 (N_1108,In_47,In_72);
and U1109 (N_1109,In_10,In_199);
xor U1110 (N_1110,In_232,In_207);
and U1111 (N_1111,In_255,In_85);
and U1112 (N_1112,In_54,In_148);
or U1113 (N_1113,In_78,In_502);
nand U1114 (N_1114,In_106,In_36);
nor U1115 (N_1115,In_638,In_359);
nand U1116 (N_1116,In_564,In_430);
or U1117 (N_1117,In_229,In_7);
xnor U1118 (N_1118,In_449,In_414);
and U1119 (N_1119,In_590,In_625);
xor U1120 (N_1120,In_312,In_460);
and U1121 (N_1121,In_185,In_237);
and U1122 (N_1122,In_335,In_556);
or U1123 (N_1123,In_707,In_111);
xor U1124 (N_1124,In_422,In_663);
xor U1125 (N_1125,In_454,In_267);
xor U1126 (N_1126,In_367,In_548);
nor U1127 (N_1127,In_50,In_130);
xnor U1128 (N_1128,In_232,In_128);
and U1129 (N_1129,In_495,In_67);
nor U1130 (N_1130,In_71,In_707);
or U1131 (N_1131,In_74,In_363);
and U1132 (N_1132,In_408,In_446);
nand U1133 (N_1133,In_563,In_481);
nand U1134 (N_1134,In_69,In_179);
and U1135 (N_1135,In_595,In_150);
or U1136 (N_1136,In_630,In_202);
or U1137 (N_1137,In_193,In_365);
nand U1138 (N_1138,In_366,In_587);
or U1139 (N_1139,In_207,In_397);
nor U1140 (N_1140,In_626,In_715);
nand U1141 (N_1141,In_292,In_135);
nand U1142 (N_1142,In_421,In_188);
xor U1143 (N_1143,In_2,In_185);
xnor U1144 (N_1144,In_363,In_232);
nand U1145 (N_1145,In_446,In_36);
nand U1146 (N_1146,In_71,In_20);
or U1147 (N_1147,In_30,In_208);
and U1148 (N_1148,In_382,In_349);
nand U1149 (N_1149,In_249,In_44);
nor U1150 (N_1150,In_601,In_218);
nand U1151 (N_1151,In_301,In_162);
or U1152 (N_1152,In_373,In_620);
or U1153 (N_1153,In_642,In_285);
nor U1154 (N_1154,In_151,In_640);
nand U1155 (N_1155,In_205,In_265);
xnor U1156 (N_1156,In_42,In_99);
nand U1157 (N_1157,In_60,In_510);
nand U1158 (N_1158,In_507,In_133);
xnor U1159 (N_1159,In_659,In_291);
nand U1160 (N_1160,In_282,In_313);
nand U1161 (N_1161,In_236,In_379);
or U1162 (N_1162,In_324,In_501);
nor U1163 (N_1163,In_644,In_626);
nor U1164 (N_1164,In_171,In_85);
or U1165 (N_1165,In_661,In_680);
xor U1166 (N_1166,In_40,In_10);
and U1167 (N_1167,In_615,In_367);
nand U1168 (N_1168,In_406,In_219);
nand U1169 (N_1169,In_693,In_696);
nand U1170 (N_1170,In_606,In_667);
or U1171 (N_1171,In_560,In_664);
nand U1172 (N_1172,In_167,In_325);
xnor U1173 (N_1173,In_497,In_138);
nand U1174 (N_1174,In_167,In_4);
and U1175 (N_1175,In_368,In_609);
xor U1176 (N_1176,In_56,In_688);
nand U1177 (N_1177,In_2,In_140);
or U1178 (N_1178,In_153,In_128);
or U1179 (N_1179,In_407,In_126);
xor U1180 (N_1180,In_667,In_589);
and U1181 (N_1181,In_458,In_378);
nor U1182 (N_1182,In_290,In_299);
or U1183 (N_1183,In_573,In_173);
nor U1184 (N_1184,In_649,In_146);
and U1185 (N_1185,In_744,In_292);
nor U1186 (N_1186,In_22,In_274);
nor U1187 (N_1187,In_403,In_412);
nand U1188 (N_1188,In_377,In_153);
xnor U1189 (N_1189,In_615,In_46);
and U1190 (N_1190,In_54,In_604);
or U1191 (N_1191,In_138,In_210);
nand U1192 (N_1192,In_637,In_653);
or U1193 (N_1193,In_658,In_419);
and U1194 (N_1194,In_5,In_541);
or U1195 (N_1195,In_2,In_266);
xor U1196 (N_1196,In_74,In_248);
or U1197 (N_1197,In_307,In_502);
xnor U1198 (N_1198,In_28,In_326);
or U1199 (N_1199,In_421,In_715);
or U1200 (N_1200,In_329,In_441);
nor U1201 (N_1201,In_334,In_184);
nand U1202 (N_1202,In_302,In_274);
and U1203 (N_1203,In_287,In_688);
nor U1204 (N_1204,In_160,In_462);
nand U1205 (N_1205,In_500,In_541);
nand U1206 (N_1206,In_200,In_554);
or U1207 (N_1207,In_219,In_491);
xor U1208 (N_1208,In_744,In_676);
nand U1209 (N_1209,In_10,In_652);
xor U1210 (N_1210,In_158,In_578);
and U1211 (N_1211,In_503,In_660);
or U1212 (N_1212,In_333,In_126);
nor U1213 (N_1213,In_594,In_5);
and U1214 (N_1214,In_118,In_731);
nand U1215 (N_1215,In_712,In_681);
xnor U1216 (N_1216,In_707,In_188);
nor U1217 (N_1217,In_588,In_615);
xnor U1218 (N_1218,In_240,In_12);
xnor U1219 (N_1219,In_102,In_387);
and U1220 (N_1220,In_53,In_706);
nor U1221 (N_1221,In_123,In_246);
xnor U1222 (N_1222,In_482,In_682);
or U1223 (N_1223,In_510,In_735);
nand U1224 (N_1224,In_271,In_489);
nor U1225 (N_1225,In_215,In_562);
or U1226 (N_1226,In_470,In_185);
nand U1227 (N_1227,In_65,In_258);
nand U1228 (N_1228,In_601,In_624);
or U1229 (N_1229,In_450,In_302);
xor U1230 (N_1230,In_314,In_118);
nand U1231 (N_1231,In_591,In_427);
nand U1232 (N_1232,In_587,In_98);
nor U1233 (N_1233,In_296,In_358);
or U1234 (N_1234,In_246,In_323);
xor U1235 (N_1235,In_503,In_654);
nand U1236 (N_1236,In_174,In_165);
xor U1237 (N_1237,In_56,In_508);
nor U1238 (N_1238,In_692,In_188);
nor U1239 (N_1239,In_492,In_425);
nand U1240 (N_1240,In_221,In_51);
or U1241 (N_1241,In_169,In_612);
nor U1242 (N_1242,In_729,In_489);
or U1243 (N_1243,In_691,In_398);
and U1244 (N_1244,In_704,In_211);
xnor U1245 (N_1245,In_574,In_365);
nand U1246 (N_1246,In_611,In_156);
xor U1247 (N_1247,In_570,In_266);
nand U1248 (N_1248,In_452,In_349);
nand U1249 (N_1249,In_435,In_574);
or U1250 (N_1250,In_16,In_39);
nor U1251 (N_1251,In_188,In_315);
or U1252 (N_1252,In_526,In_444);
and U1253 (N_1253,In_634,In_739);
or U1254 (N_1254,In_77,In_592);
xnor U1255 (N_1255,In_338,In_540);
nor U1256 (N_1256,In_225,In_421);
and U1257 (N_1257,In_728,In_388);
and U1258 (N_1258,In_323,In_487);
or U1259 (N_1259,In_340,In_189);
nand U1260 (N_1260,In_255,In_390);
or U1261 (N_1261,In_31,In_213);
nand U1262 (N_1262,In_52,In_715);
xor U1263 (N_1263,In_42,In_125);
and U1264 (N_1264,In_49,In_281);
or U1265 (N_1265,In_393,In_378);
nand U1266 (N_1266,In_455,In_379);
nand U1267 (N_1267,In_530,In_470);
and U1268 (N_1268,In_414,In_316);
xnor U1269 (N_1269,In_293,In_520);
nor U1270 (N_1270,In_254,In_352);
nand U1271 (N_1271,In_90,In_211);
and U1272 (N_1272,In_61,In_504);
or U1273 (N_1273,In_529,In_41);
nand U1274 (N_1274,In_290,In_609);
nor U1275 (N_1275,In_9,In_372);
and U1276 (N_1276,In_605,In_618);
or U1277 (N_1277,In_700,In_722);
xnor U1278 (N_1278,In_121,In_708);
or U1279 (N_1279,In_302,In_36);
nand U1280 (N_1280,In_619,In_627);
xor U1281 (N_1281,In_703,In_424);
and U1282 (N_1282,In_198,In_734);
and U1283 (N_1283,In_511,In_294);
and U1284 (N_1284,In_358,In_580);
or U1285 (N_1285,In_661,In_603);
and U1286 (N_1286,In_296,In_84);
nand U1287 (N_1287,In_238,In_214);
or U1288 (N_1288,In_195,In_645);
nor U1289 (N_1289,In_560,In_715);
and U1290 (N_1290,In_131,In_317);
or U1291 (N_1291,In_747,In_7);
nor U1292 (N_1292,In_77,In_38);
xor U1293 (N_1293,In_661,In_153);
and U1294 (N_1294,In_15,In_615);
nand U1295 (N_1295,In_611,In_150);
nor U1296 (N_1296,In_540,In_390);
and U1297 (N_1297,In_413,In_151);
or U1298 (N_1298,In_695,In_388);
xnor U1299 (N_1299,In_210,In_513);
xnor U1300 (N_1300,In_478,In_499);
nor U1301 (N_1301,In_107,In_199);
xnor U1302 (N_1302,In_744,In_546);
and U1303 (N_1303,In_594,In_54);
and U1304 (N_1304,In_679,In_428);
or U1305 (N_1305,In_193,In_429);
nand U1306 (N_1306,In_632,In_747);
and U1307 (N_1307,In_287,In_283);
xor U1308 (N_1308,In_464,In_549);
nor U1309 (N_1309,In_626,In_609);
nor U1310 (N_1310,In_319,In_393);
nor U1311 (N_1311,In_655,In_665);
and U1312 (N_1312,In_259,In_681);
or U1313 (N_1313,In_743,In_431);
and U1314 (N_1314,In_602,In_700);
xor U1315 (N_1315,In_475,In_519);
nand U1316 (N_1316,In_469,In_114);
or U1317 (N_1317,In_439,In_553);
or U1318 (N_1318,In_489,In_201);
nor U1319 (N_1319,In_527,In_683);
nor U1320 (N_1320,In_191,In_706);
or U1321 (N_1321,In_642,In_385);
or U1322 (N_1322,In_377,In_89);
xor U1323 (N_1323,In_319,In_90);
or U1324 (N_1324,In_465,In_86);
xnor U1325 (N_1325,In_746,In_267);
nand U1326 (N_1326,In_442,In_467);
and U1327 (N_1327,In_311,In_627);
and U1328 (N_1328,In_664,In_450);
and U1329 (N_1329,In_201,In_431);
or U1330 (N_1330,In_392,In_542);
nor U1331 (N_1331,In_422,In_645);
nor U1332 (N_1332,In_551,In_249);
and U1333 (N_1333,In_151,In_163);
nor U1334 (N_1334,In_95,In_733);
xnor U1335 (N_1335,In_158,In_86);
or U1336 (N_1336,In_264,In_86);
and U1337 (N_1337,In_127,In_345);
and U1338 (N_1338,In_51,In_659);
nand U1339 (N_1339,In_262,In_727);
or U1340 (N_1340,In_302,In_122);
or U1341 (N_1341,In_197,In_460);
nor U1342 (N_1342,In_459,In_654);
xnor U1343 (N_1343,In_221,In_504);
nand U1344 (N_1344,In_244,In_698);
and U1345 (N_1345,In_368,In_714);
nand U1346 (N_1346,In_717,In_348);
xor U1347 (N_1347,In_339,In_245);
and U1348 (N_1348,In_281,In_261);
xnor U1349 (N_1349,In_688,In_511);
and U1350 (N_1350,In_177,In_455);
nand U1351 (N_1351,In_746,In_472);
or U1352 (N_1352,In_123,In_610);
and U1353 (N_1353,In_706,In_11);
nand U1354 (N_1354,In_514,In_331);
nor U1355 (N_1355,In_681,In_64);
nor U1356 (N_1356,In_267,In_494);
and U1357 (N_1357,In_429,In_543);
and U1358 (N_1358,In_232,In_246);
or U1359 (N_1359,In_318,In_710);
xor U1360 (N_1360,In_623,In_309);
or U1361 (N_1361,In_605,In_282);
nor U1362 (N_1362,In_129,In_213);
xnor U1363 (N_1363,In_424,In_299);
or U1364 (N_1364,In_371,In_151);
xor U1365 (N_1365,In_552,In_173);
or U1366 (N_1366,In_256,In_337);
or U1367 (N_1367,In_509,In_104);
nor U1368 (N_1368,In_658,In_649);
and U1369 (N_1369,In_592,In_96);
nor U1370 (N_1370,In_621,In_388);
and U1371 (N_1371,In_645,In_558);
nor U1372 (N_1372,In_604,In_6);
or U1373 (N_1373,In_603,In_442);
and U1374 (N_1374,In_170,In_203);
and U1375 (N_1375,In_304,In_483);
and U1376 (N_1376,In_583,In_708);
xor U1377 (N_1377,In_348,In_225);
nor U1378 (N_1378,In_53,In_343);
nand U1379 (N_1379,In_511,In_387);
xnor U1380 (N_1380,In_611,In_38);
or U1381 (N_1381,In_553,In_25);
or U1382 (N_1382,In_303,In_293);
nand U1383 (N_1383,In_69,In_665);
and U1384 (N_1384,In_331,In_522);
xor U1385 (N_1385,In_265,In_569);
and U1386 (N_1386,In_196,In_331);
nand U1387 (N_1387,In_6,In_265);
nand U1388 (N_1388,In_516,In_99);
and U1389 (N_1389,In_81,In_443);
and U1390 (N_1390,In_236,In_396);
nor U1391 (N_1391,In_723,In_43);
and U1392 (N_1392,In_365,In_67);
nor U1393 (N_1393,In_82,In_88);
nand U1394 (N_1394,In_662,In_435);
nor U1395 (N_1395,In_399,In_101);
and U1396 (N_1396,In_468,In_252);
or U1397 (N_1397,In_624,In_509);
nor U1398 (N_1398,In_324,In_534);
and U1399 (N_1399,In_52,In_246);
xor U1400 (N_1400,In_410,In_695);
or U1401 (N_1401,In_597,In_662);
nand U1402 (N_1402,In_94,In_701);
and U1403 (N_1403,In_494,In_173);
nand U1404 (N_1404,In_395,In_169);
and U1405 (N_1405,In_366,In_733);
xnor U1406 (N_1406,In_71,In_494);
or U1407 (N_1407,In_409,In_238);
nand U1408 (N_1408,In_708,In_414);
nand U1409 (N_1409,In_408,In_320);
and U1410 (N_1410,In_636,In_13);
xnor U1411 (N_1411,In_426,In_494);
nor U1412 (N_1412,In_47,In_631);
and U1413 (N_1413,In_301,In_662);
nor U1414 (N_1414,In_615,In_380);
and U1415 (N_1415,In_90,In_36);
nand U1416 (N_1416,In_601,In_371);
and U1417 (N_1417,In_708,In_359);
nand U1418 (N_1418,In_536,In_512);
and U1419 (N_1419,In_455,In_375);
xor U1420 (N_1420,In_579,In_733);
and U1421 (N_1421,In_97,In_255);
or U1422 (N_1422,In_6,In_69);
nor U1423 (N_1423,In_261,In_357);
or U1424 (N_1424,In_199,In_316);
xor U1425 (N_1425,In_352,In_356);
and U1426 (N_1426,In_404,In_22);
or U1427 (N_1427,In_614,In_263);
and U1428 (N_1428,In_2,In_628);
xnor U1429 (N_1429,In_490,In_729);
nor U1430 (N_1430,In_524,In_400);
or U1431 (N_1431,In_566,In_604);
and U1432 (N_1432,In_60,In_31);
nand U1433 (N_1433,In_217,In_154);
or U1434 (N_1434,In_531,In_14);
nand U1435 (N_1435,In_670,In_633);
nand U1436 (N_1436,In_484,In_369);
nor U1437 (N_1437,In_359,In_686);
nand U1438 (N_1438,In_353,In_155);
nor U1439 (N_1439,In_235,In_608);
and U1440 (N_1440,In_565,In_369);
and U1441 (N_1441,In_252,In_460);
xor U1442 (N_1442,In_43,In_158);
or U1443 (N_1443,In_585,In_325);
nor U1444 (N_1444,In_526,In_447);
or U1445 (N_1445,In_74,In_90);
or U1446 (N_1446,In_295,In_84);
xor U1447 (N_1447,In_676,In_262);
or U1448 (N_1448,In_194,In_709);
xnor U1449 (N_1449,In_351,In_579);
xor U1450 (N_1450,In_315,In_463);
and U1451 (N_1451,In_270,In_424);
nand U1452 (N_1452,In_545,In_346);
nor U1453 (N_1453,In_465,In_615);
and U1454 (N_1454,In_251,In_143);
xnor U1455 (N_1455,In_630,In_470);
xor U1456 (N_1456,In_418,In_592);
or U1457 (N_1457,In_508,In_620);
xor U1458 (N_1458,In_43,In_663);
nor U1459 (N_1459,In_215,In_117);
xnor U1460 (N_1460,In_704,In_8);
xnor U1461 (N_1461,In_4,In_316);
or U1462 (N_1462,In_40,In_707);
and U1463 (N_1463,In_318,In_44);
xnor U1464 (N_1464,In_390,In_68);
nor U1465 (N_1465,In_277,In_730);
nor U1466 (N_1466,In_646,In_513);
nand U1467 (N_1467,In_619,In_686);
or U1468 (N_1468,In_565,In_137);
or U1469 (N_1469,In_417,In_678);
nand U1470 (N_1470,In_711,In_718);
and U1471 (N_1471,In_28,In_450);
xor U1472 (N_1472,In_28,In_458);
xor U1473 (N_1473,In_154,In_439);
or U1474 (N_1474,In_380,In_704);
nor U1475 (N_1475,In_521,In_115);
nand U1476 (N_1476,In_349,In_560);
and U1477 (N_1477,In_385,In_354);
and U1478 (N_1478,In_181,In_718);
xor U1479 (N_1479,In_748,In_398);
nand U1480 (N_1480,In_594,In_730);
xnor U1481 (N_1481,In_336,In_72);
xnor U1482 (N_1482,In_718,In_607);
nor U1483 (N_1483,In_137,In_567);
and U1484 (N_1484,In_232,In_540);
and U1485 (N_1485,In_210,In_90);
xor U1486 (N_1486,In_42,In_157);
or U1487 (N_1487,In_300,In_420);
nor U1488 (N_1488,In_140,In_207);
and U1489 (N_1489,In_206,In_310);
nand U1490 (N_1490,In_258,In_573);
xor U1491 (N_1491,In_531,In_179);
nor U1492 (N_1492,In_388,In_260);
or U1493 (N_1493,In_0,In_317);
and U1494 (N_1494,In_659,In_409);
nand U1495 (N_1495,In_383,In_698);
or U1496 (N_1496,In_313,In_508);
nor U1497 (N_1497,In_457,In_1);
nor U1498 (N_1498,In_556,In_20);
xor U1499 (N_1499,In_132,In_150);
nand U1500 (N_1500,In_608,In_271);
or U1501 (N_1501,In_704,In_57);
or U1502 (N_1502,In_110,In_320);
nor U1503 (N_1503,In_468,In_138);
and U1504 (N_1504,In_525,In_260);
nand U1505 (N_1505,In_639,In_544);
xor U1506 (N_1506,In_78,In_592);
or U1507 (N_1507,In_582,In_639);
nand U1508 (N_1508,In_503,In_677);
nand U1509 (N_1509,In_122,In_113);
or U1510 (N_1510,In_282,In_326);
nand U1511 (N_1511,In_727,In_120);
xor U1512 (N_1512,In_544,In_164);
or U1513 (N_1513,In_741,In_278);
xnor U1514 (N_1514,In_421,In_64);
nand U1515 (N_1515,In_411,In_175);
xnor U1516 (N_1516,In_15,In_308);
xnor U1517 (N_1517,In_295,In_102);
nand U1518 (N_1518,In_303,In_337);
nand U1519 (N_1519,In_683,In_358);
and U1520 (N_1520,In_32,In_15);
or U1521 (N_1521,In_401,In_324);
and U1522 (N_1522,In_384,In_108);
nand U1523 (N_1523,In_53,In_300);
and U1524 (N_1524,In_433,In_398);
and U1525 (N_1525,In_214,In_286);
and U1526 (N_1526,In_644,In_678);
nand U1527 (N_1527,In_645,In_154);
xor U1528 (N_1528,In_668,In_173);
nor U1529 (N_1529,In_93,In_293);
xnor U1530 (N_1530,In_83,In_231);
or U1531 (N_1531,In_456,In_251);
xnor U1532 (N_1532,In_648,In_685);
xor U1533 (N_1533,In_336,In_699);
xnor U1534 (N_1534,In_364,In_594);
nand U1535 (N_1535,In_23,In_425);
nor U1536 (N_1536,In_84,In_233);
and U1537 (N_1537,In_510,In_715);
and U1538 (N_1538,In_662,In_539);
xor U1539 (N_1539,In_137,In_702);
nand U1540 (N_1540,In_368,In_338);
or U1541 (N_1541,In_407,In_213);
or U1542 (N_1542,In_270,In_625);
xor U1543 (N_1543,In_90,In_378);
nor U1544 (N_1544,In_349,In_563);
or U1545 (N_1545,In_340,In_363);
or U1546 (N_1546,In_313,In_579);
nor U1547 (N_1547,In_265,In_59);
nand U1548 (N_1548,In_630,In_453);
nand U1549 (N_1549,In_54,In_285);
or U1550 (N_1550,In_76,In_559);
nand U1551 (N_1551,In_382,In_564);
or U1552 (N_1552,In_651,In_395);
or U1553 (N_1553,In_100,In_740);
or U1554 (N_1554,In_235,In_489);
nor U1555 (N_1555,In_533,In_116);
nand U1556 (N_1556,In_506,In_193);
nor U1557 (N_1557,In_312,In_375);
nand U1558 (N_1558,In_594,In_294);
and U1559 (N_1559,In_338,In_483);
nor U1560 (N_1560,In_334,In_561);
nor U1561 (N_1561,In_11,In_223);
nand U1562 (N_1562,In_29,In_744);
nand U1563 (N_1563,In_170,In_642);
nand U1564 (N_1564,In_645,In_356);
xnor U1565 (N_1565,In_154,In_601);
nand U1566 (N_1566,In_381,In_202);
or U1567 (N_1567,In_577,In_346);
and U1568 (N_1568,In_530,In_410);
and U1569 (N_1569,In_482,In_292);
or U1570 (N_1570,In_179,In_255);
xnor U1571 (N_1571,In_162,In_382);
or U1572 (N_1572,In_665,In_402);
nor U1573 (N_1573,In_529,In_649);
nand U1574 (N_1574,In_322,In_711);
or U1575 (N_1575,In_119,In_528);
nand U1576 (N_1576,In_745,In_79);
or U1577 (N_1577,In_541,In_174);
or U1578 (N_1578,In_280,In_576);
and U1579 (N_1579,In_716,In_108);
and U1580 (N_1580,In_242,In_616);
xnor U1581 (N_1581,In_454,In_385);
xor U1582 (N_1582,In_120,In_126);
and U1583 (N_1583,In_459,In_678);
xnor U1584 (N_1584,In_693,In_158);
xor U1585 (N_1585,In_65,In_14);
nand U1586 (N_1586,In_203,In_8);
xnor U1587 (N_1587,In_208,In_601);
and U1588 (N_1588,In_320,In_180);
nor U1589 (N_1589,In_93,In_292);
or U1590 (N_1590,In_741,In_686);
and U1591 (N_1591,In_211,In_34);
nor U1592 (N_1592,In_122,In_298);
xnor U1593 (N_1593,In_45,In_698);
and U1594 (N_1594,In_714,In_118);
nand U1595 (N_1595,In_432,In_408);
xnor U1596 (N_1596,In_173,In_431);
nor U1597 (N_1597,In_455,In_619);
or U1598 (N_1598,In_560,In_518);
xnor U1599 (N_1599,In_601,In_279);
nand U1600 (N_1600,In_590,In_125);
and U1601 (N_1601,In_297,In_322);
nor U1602 (N_1602,In_203,In_109);
nor U1603 (N_1603,In_535,In_310);
and U1604 (N_1604,In_260,In_177);
and U1605 (N_1605,In_293,In_575);
nor U1606 (N_1606,In_573,In_428);
xor U1607 (N_1607,In_441,In_701);
nor U1608 (N_1608,In_365,In_18);
nor U1609 (N_1609,In_273,In_63);
nor U1610 (N_1610,In_289,In_574);
and U1611 (N_1611,In_262,In_188);
nor U1612 (N_1612,In_15,In_588);
nand U1613 (N_1613,In_338,In_202);
or U1614 (N_1614,In_641,In_490);
and U1615 (N_1615,In_700,In_311);
or U1616 (N_1616,In_335,In_209);
and U1617 (N_1617,In_346,In_424);
or U1618 (N_1618,In_115,In_225);
nand U1619 (N_1619,In_251,In_16);
nor U1620 (N_1620,In_746,In_167);
and U1621 (N_1621,In_72,In_552);
nor U1622 (N_1622,In_54,In_644);
nand U1623 (N_1623,In_95,In_514);
or U1624 (N_1624,In_237,In_468);
nand U1625 (N_1625,In_497,In_390);
or U1626 (N_1626,In_496,In_597);
or U1627 (N_1627,In_319,In_330);
and U1628 (N_1628,In_683,In_563);
nand U1629 (N_1629,In_111,In_404);
and U1630 (N_1630,In_388,In_103);
nor U1631 (N_1631,In_276,In_505);
or U1632 (N_1632,In_334,In_520);
xor U1633 (N_1633,In_409,In_94);
xnor U1634 (N_1634,In_516,In_639);
and U1635 (N_1635,In_150,In_245);
nor U1636 (N_1636,In_282,In_503);
or U1637 (N_1637,In_297,In_123);
nor U1638 (N_1638,In_145,In_28);
or U1639 (N_1639,In_450,In_262);
xor U1640 (N_1640,In_1,In_144);
or U1641 (N_1641,In_165,In_324);
or U1642 (N_1642,In_304,In_589);
or U1643 (N_1643,In_426,In_307);
nand U1644 (N_1644,In_352,In_285);
nand U1645 (N_1645,In_567,In_598);
nand U1646 (N_1646,In_84,In_737);
or U1647 (N_1647,In_344,In_728);
and U1648 (N_1648,In_153,In_99);
xor U1649 (N_1649,In_432,In_537);
xor U1650 (N_1650,In_17,In_296);
nand U1651 (N_1651,In_162,In_211);
nand U1652 (N_1652,In_496,In_413);
xnor U1653 (N_1653,In_455,In_85);
nor U1654 (N_1654,In_695,In_331);
nor U1655 (N_1655,In_740,In_475);
or U1656 (N_1656,In_739,In_373);
or U1657 (N_1657,In_69,In_96);
and U1658 (N_1658,In_504,In_372);
or U1659 (N_1659,In_158,In_71);
xor U1660 (N_1660,In_31,In_650);
nand U1661 (N_1661,In_293,In_264);
nand U1662 (N_1662,In_539,In_552);
or U1663 (N_1663,In_509,In_628);
and U1664 (N_1664,In_565,In_197);
or U1665 (N_1665,In_378,In_546);
and U1666 (N_1666,In_392,In_189);
nand U1667 (N_1667,In_698,In_73);
nand U1668 (N_1668,In_104,In_158);
or U1669 (N_1669,In_396,In_25);
nor U1670 (N_1670,In_432,In_653);
or U1671 (N_1671,In_259,In_175);
and U1672 (N_1672,In_276,In_185);
xnor U1673 (N_1673,In_370,In_221);
xnor U1674 (N_1674,In_533,In_388);
nand U1675 (N_1675,In_253,In_655);
or U1676 (N_1676,In_730,In_244);
or U1677 (N_1677,In_548,In_318);
or U1678 (N_1678,In_83,In_429);
nand U1679 (N_1679,In_681,In_267);
xor U1680 (N_1680,In_412,In_413);
nor U1681 (N_1681,In_511,In_84);
or U1682 (N_1682,In_175,In_57);
nor U1683 (N_1683,In_383,In_682);
or U1684 (N_1684,In_671,In_716);
or U1685 (N_1685,In_523,In_355);
xor U1686 (N_1686,In_423,In_373);
xor U1687 (N_1687,In_130,In_382);
nor U1688 (N_1688,In_528,In_491);
and U1689 (N_1689,In_135,In_2);
nand U1690 (N_1690,In_688,In_66);
nor U1691 (N_1691,In_744,In_642);
and U1692 (N_1692,In_139,In_231);
and U1693 (N_1693,In_482,In_731);
nor U1694 (N_1694,In_463,In_311);
or U1695 (N_1695,In_689,In_103);
xnor U1696 (N_1696,In_251,In_188);
nand U1697 (N_1697,In_140,In_523);
and U1698 (N_1698,In_198,In_171);
nand U1699 (N_1699,In_96,In_452);
and U1700 (N_1700,In_426,In_474);
and U1701 (N_1701,In_156,In_441);
or U1702 (N_1702,In_615,In_202);
or U1703 (N_1703,In_676,In_655);
xor U1704 (N_1704,In_107,In_245);
and U1705 (N_1705,In_667,In_129);
nand U1706 (N_1706,In_405,In_199);
and U1707 (N_1707,In_110,In_138);
nor U1708 (N_1708,In_153,In_165);
or U1709 (N_1709,In_527,In_492);
nand U1710 (N_1710,In_5,In_393);
nor U1711 (N_1711,In_163,In_745);
nor U1712 (N_1712,In_612,In_126);
or U1713 (N_1713,In_665,In_274);
and U1714 (N_1714,In_1,In_420);
and U1715 (N_1715,In_203,In_4);
nand U1716 (N_1716,In_184,In_82);
nand U1717 (N_1717,In_383,In_386);
xor U1718 (N_1718,In_182,In_386);
nand U1719 (N_1719,In_457,In_388);
xor U1720 (N_1720,In_8,In_115);
and U1721 (N_1721,In_613,In_204);
xnor U1722 (N_1722,In_612,In_15);
nand U1723 (N_1723,In_8,In_49);
or U1724 (N_1724,In_343,In_505);
and U1725 (N_1725,In_363,In_73);
xnor U1726 (N_1726,In_91,In_312);
or U1727 (N_1727,In_525,In_286);
nand U1728 (N_1728,In_538,In_361);
and U1729 (N_1729,In_681,In_664);
nand U1730 (N_1730,In_152,In_114);
or U1731 (N_1731,In_272,In_184);
nor U1732 (N_1732,In_476,In_324);
xnor U1733 (N_1733,In_216,In_709);
nand U1734 (N_1734,In_269,In_424);
nand U1735 (N_1735,In_478,In_604);
or U1736 (N_1736,In_404,In_342);
or U1737 (N_1737,In_111,In_325);
nand U1738 (N_1738,In_34,In_445);
and U1739 (N_1739,In_602,In_103);
nand U1740 (N_1740,In_636,In_516);
or U1741 (N_1741,In_463,In_140);
and U1742 (N_1742,In_574,In_379);
and U1743 (N_1743,In_328,In_392);
nand U1744 (N_1744,In_408,In_184);
xnor U1745 (N_1745,In_454,In_534);
or U1746 (N_1746,In_63,In_495);
nand U1747 (N_1747,In_727,In_583);
and U1748 (N_1748,In_710,In_684);
nor U1749 (N_1749,In_674,In_185);
nor U1750 (N_1750,In_165,In_203);
nand U1751 (N_1751,In_55,In_504);
nand U1752 (N_1752,In_733,In_493);
and U1753 (N_1753,In_465,In_658);
nand U1754 (N_1754,In_417,In_66);
and U1755 (N_1755,In_605,In_660);
or U1756 (N_1756,In_49,In_355);
nor U1757 (N_1757,In_412,In_44);
and U1758 (N_1758,In_334,In_64);
or U1759 (N_1759,In_373,In_406);
nor U1760 (N_1760,In_616,In_142);
nand U1761 (N_1761,In_630,In_3);
nor U1762 (N_1762,In_628,In_632);
nor U1763 (N_1763,In_721,In_728);
nand U1764 (N_1764,In_143,In_575);
xor U1765 (N_1765,In_691,In_563);
nand U1766 (N_1766,In_392,In_599);
nand U1767 (N_1767,In_9,In_139);
nor U1768 (N_1768,In_551,In_299);
nand U1769 (N_1769,In_581,In_277);
xor U1770 (N_1770,In_717,In_516);
or U1771 (N_1771,In_677,In_732);
nand U1772 (N_1772,In_667,In_149);
xor U1773 (N_1773,In_504,In_267);
or U1774 (N_1774,In_526,In_450);
and U1775 (N_1775,In_55,In_429);
and U1776 (N_1776,In_379,In_295);
nand U1777 (N_1777,In_693,In_405);
or U1778 (N_1778,In_22,In_348);
nand U1779 (N_1779,In_31,In_109);
or U1780 (N_1780,In_103,In_542);
nand U1781 (N_1781,In_57,In_515);
or U1782 (N_1782,In_180,In_537);
xnor U1783 (N_1783,In_222,In_324);
and U1784 (N_1784,In_304,In_497);
or U1785 (N_1785,In_664,In_682);
xnor U1786 (N_1786,In_8,In_477);
and U1787 (N_1787,In_306,In_555);
nor U1788 (N_1788,In_210,In_250);
nand U1789 (N_1789,In_73,In_403);
or U1790 (N_1790,In_185,In_552);
and U1791 (N_1791,In_332,In_517);
xor U1792 (N_1792,In_389,In_739);
xor U1793 (N_1793,In_609,In_488);
nand U1794 (N_1794,In_105,In_181);
or U1795 (N_1795,In_687,In_122);
nor U1796 (N_1796,In_469,In_579);
nor U1797 (N_1797,In_49,In_537);
and U1798 (N_1798,In_658,In_475);
or U1799 (N_1799,In_420,In_50);
nand U1800 (N_1800,In_122,In_76);
nand U1801 (N_1801,In_178,In_37);
or U1802 (N_1802,In_355,In_496);
nor U1803 (N_1803,In_39,In_613);
and U1804 (N_1804,In_735,In_188);
or U1805 (N_1805,In_471,In_364);
or U1806 (N_1806,In_695,In_154);
xnor U1807 (N_1807,In_665,In_249);
xor U1808 (N_1808,In_422,In_585);
or U1809 (N_1809,In_704,In_93);
xor U1810 (N_1810,In_108,In_278);
nor U1811 (N_1811,In_193,In_55);
nand U1812 (N_1812,In_720,In_457);
xnor U1813 (N_1813,In_4,In_572);
and U1814 (N_1814,In_372,In_720);
xor U1815 (N_1815,In_354,In_473);
nand U1816 (N_1816,In_336,In_66);
xor U1817 (N_1817,In_450,In_108);
nor U1818 (N_1818,In_609,In_132);
and U1819 (N_1819,In_96,In_482);
nand U1820 (N_1820,In_741,In_270);
and U1821 (N_1821,In_705,In_318);
nand U1822 (N_1822,In_249,In_122);
nor U1823 (N_1823,In_3,In_187);
xor U1824 (N_1824,In_738,In_314);
or U1825 (N_1825,In_599,In_730);
nor U1826 (N_1826,In_313,In_275);
and U1827 (N_1827,In_393,In_622);
xor U1828 (N_1828,In_434,In_60);
or U1829 (N_1829,In_125,In_451);
and U1830 (N_1830,In_366,In_175);
and U1831 (N_1831,In_6,In_54);
nor U1832 (N_1832,In_30,In_717);
or U1833 (N_1833,In_545,In_635);
or U1834 (N_1834,In_740,In_581);
nor U1835 (N_1835,In_126,In_483);
and U1836 (N_1836,In_551,In_185);
nand U1837 (N_1837,In_342,In_112);
xnor U1838 (N_1838,In_222,In_58);
or U1839 (N_1839,In_18,In_200);
nand U1840 (N_1840,In_302,In_342);
nand U1841 (N_1841,In_572,In_415);
nand U1842 (N_1842,In_33,In_88);
and U1843 (N_1843,In_591,In_270);
nand U1844 (N_1844,In_587,In_210);
and U1845 (N_1845,In_366,In_249);
xnor U1846 (N_1846,In_348,In_527);
or U1847 (N_1847,In_536,In_312);
nand U1848 (N_1848,In_14,In_102);
nor U1849 (N_1849,In_55,In_488);
or U1850 (N_1850,In_643,In_523);
or U1851 (N_1851,In_742,In_376);
nor U1852 (N_1852,In_244,In_448);
nor U1853 (N_1853,In_628,In_448);
nand U1854 (N_1854,In_211,In_66);
xnor U1855 (N_1855,In_386,In_331);
xor U1856 (N_1856,In_84,In_590);
nor U1857 (N_1857,In_36,In_157);
nor U1858 (N_1858,In_360,In_667);
xor U1859 (N_1859,In_680,In_448);
nor U1860 (N_1860,In_542,In_511);
nand U1861 (N_1861,In_668,In_225);
and U1862 (N_1862,In_325,In_291);
nand U1863 (N_1863,In_700,In_617);
xor U1864 (N_1864,In_203,In_662);
and U1865 (N_1865,In_709,In_220);
and U1866 (N_1866,In_521,In_351);
and U1867 (N_1867,In_346,In_83);
xnor U1868 (N_1868,In_55,In_108);
nand U1869 (N_1869,In_354,In_671);
nor U1870 (N_1870,In_99,In_216);
nor U1871 (N_1871,In_497,In_634);
xnor U1872 (N_1872,In_243,In_435);
nand U1873 (N_1873,In_73,In_318);
or U1874 (N_1874,In_265,In_367);
or U1875 (N_1875,In_402,In_9);
nor U1876 (N_1876,In_370,In_526);
xor U1877 (N_1877,In_460,In_300);
xor U1878 (N_1878,In_83,In_368);
and U1879 (N_1879,In_745,In_557);
nor U1880 (N_1880,In_635,In_370);
or U1881 (N_1881,In_308,In_483);
xnor U1882 (N_1882,In_411,In_456);
nor U1883 (N_1883,In_737,In_64);
nand U1884 (N_1884,In_303,In_272);
xnor U1885 (N_1885,In_42,In_709);
and U1886 (N_1886,In_367,In_512);
or U1887 (N_1887,In_250,In_725);
nand U1888 (N_1888,In_381,In_528);
and U1889 (N_1889,In_207,In_309);
nor U1890 (N_1890,In_331,In_197);
and U1891 (N_1891,In_165,In_297);
or U1892 (N_1892,In_612,In_208);
or U1893 (N_1893,In_3,In_215);
nor U1894 (N_1894,In_178,In_195);
or U1895 (N_1895,In_61,In_96);
and U1896 (N_1896,In_674,In_556);
or U1897 (N_1897,In_571,In_418);
nor U1898 (N_1898,In_682,In_579);
or U1899 (N_1899,In_423,In_319);
nor U1900 (N_1900,In_512,In_304);
or U1901 (N_1901,In_466,In_472);
or U1902 (N_1902,In_166,In_591);
and U1903 (N_1903,In_204,In_250);
and U1904 (N_1904,In_413,In_728);
nor U1905 (N_1905,In_279,In_718);
xnor U1906 (N_1906,In_32,In_355);
xor U1907 (N_1907,In_505,In_619);
xor U1908 (N_1908,In_208,In_57);
nand U1909 (N_1909,In_647,In_162);
and U1910 (N_1910,In_93,In_612);
nor U1911 (N_1911,In_11,In_337);
and U1912 (N_1912,In_285,In_428);
nand U1913 (N_1913,In_98,In_521);
and U1914 (N_1914,In_95,In_123);
xnor U1915 (N_1915,In_488,In_518);
xnor U1916 (N_1916,In_37,In_539);
xnor U1917 (N_1917,In_720,In_303);
nor U1918 (N_1918,In_75,In_523);
or U1919 (N_1919,In_217,In_557);
or U1920 (N_1920,In_581,In_95);
nor U1921 (N_1921,In_450,In_414);
and U1922 (N_1922,In_424,In_468);
and U1923 (N_1923,In_704,In_372);
and U1924 (N_1924,In_683,In_419);
xnor U1925 (N_1925,In_288,In_434);
or U1926 (N_1926,In_300,In_69);
and U1927 (N_1927,In_511,In_693);
nand U1928 (N_1928,In_311,In_199);
nand U1929 (N_1929,In_474,In_581);
or U1930 (N_1930,In_732,In_181);
and U1931 (N_1931,In_385,In_567);
nor U1932 (N_1932,In_5,In_451);
nor U1933 (N_1933,In_373,In_153);
and U1934 (N_1934,In_188,In_737);
or U1935 (N_1935,In_490,In_362);
nor U1936 (N_1936,In_78,In_213);
and U1937 (N_1937,In_219,In_351);
and U1938 (N_1938,In_42,In_280);
nand U1939 (N_1939,In_727,In_679);
nand U1940 (N_1940,In_514,In_47);
nand U1941 (N_1941,In_68,In_56);
nand U1942 (N_1942,In_236,In_655);
nor U1943 (N_1943,In_614,In_248);
xnor U1944 (N_1944,In_227,In_361);
or U1945 (N_1945,In_501,In_532);
xnor U1946 (N_1946,In_432,In_292);
or U1947 (N_1947,In_415,In_189);
nand U1948 (N_1948,In_712,In_722);
nand U1949 (N_1949,In_248,In_624);
xnor U1950 (N_1950,In_582,In_239);
and U1951 (N_1951,In_233,In_156);
or U1952 (N_1952,In_47,In_96);
nor U1953 (N_1953,In_366,In_508);
and U1954 (N_1954,In_487,In_215);
or U1955 (N_1955,In_273,In_393);
and U1956 (N_1956,In_272,In_104);
nand U1957 (N_1957,In_731,In_227);
nor U1958 (N_1958,In_331,In_486);
nand U1959 (N_1959,In_486,In_551);
nor U1960 (N_1960,In_34,In_241);
xnor U1961 (N_1961,In_387,In_444);
and U1962 (N_1962,In_96,In_461);
and U1963 (N_1963,In_203,In_306);
nand U1964 (N_1964,In_412,In_260);
nor U1965 (N_1965,In_29,In_728);
or U1966 (N_1966,In_546,In_657);
nor U1967 (N_1967,In_658,In_499);
or U1968 (N_1968,In_336,In_205);
xnor U1969 (N_1969,In_158,In_90);
or U1970 (N_1970,In_29,In_574);
xor U1971 (N_1971,In_114,In_79);
xnor U1972 (N_1972,In_526,In_283);
nand U1973 (N_1973,In_596,In_323);
and U1974 (N_1974,In_693,In_610);
nand U1975 (N_1975,In_413,In_98);
xor U1976 (N_1976,In_745,In_291);
or U1977 (N_1977,In_532,In_38);
nor U1978 (N_1978,In_632,In_494);
or U1979 (N_1979,In_473,In_399);
or U1980 (N_1980,In_588,In_484);
nand U1981 (N_1981,In_364,In_42);
xor U1982 (N_1982,In_255,In_357);
nor U1983 (N_1983,In_139,In_505);
or U1984 (N_1984,In_260,In_109);
xor U1985 (N_1985,In_462,In_152);
and U1986 (N_1986,In_555,In_521);
nor U1987 (N_1987,In_336,In_693);
or U1988 (N_1988,In_271,In_13);
nor U1989 (N_1989,In_668,In_66);
or U1990 (N_1990,In_483,In_554);
nand U1991 (N_1991,In_82,In_445);
or U1992 (N_1992,In_84,In_749);
xnor U1993 (N_1993,In_256,In_217);
nor U1994 (N_1994,In_563,In_443);
or U1995 (N_1995,In_658,In_274);
nor U1996 (N_1996,In_304,In_52);
or U1997 (N_1997,In_681,In_418);
and U1998 (N_1998,In_605,In_537);
and U1999 (N_1999,In_633,In_715);
or U2000 (N_2000,In_361,In_287);
xnor U2001 (N_2001,In_407,In_733);
and U2002 (N_2002,In_141,In_49);
and U2003 (N_2003,In_201,In_484);
and U2004 (N_2004,In_497,In_596);
and U2005 (N_2005,In_524,In_26);
xor U2006 (N_2006,In_53,In_368);
and U2007 (N_2007,In_320,In_333);
xor U2008 (N_2008,In_614,In_47);
nor U2009 (N_2009,In_370,In_437);
nor U2010 (N_2010,In_314,In_224);
or U2011 (N_2011,In_123,In_140);
nor U2012 (N_2012,In_11,In_419);
nor U2013 (N_2013,In_276,In_367);
and U2014 (N_2014,In_64,In_459);
nor U2015 (N_2015,In_356,In_199);
nand U2016 (N_2016,In_39,In_261);
nor U2017 (N_2017,In_254,In_236);
and U2018 (N_2018,In_289,In_56);
xnor U2019 (N_2019,In_332,In_211);
xnor U2020 (N_2020,In_66,In_345);
and U2021 (N_2021,In_454,In_281);
or U2022 (N_2022,In_236,In_292);
or U2023 (N_2023,In_601,In_201);
nand U2024 (N_2024,In_659,In_632);
or U2025 (N_2025,In_385,In_170);
xor U2026 (N_2026,In_88,In_670);
nor U2027 (N_2027,In_676,In_503);
nor U2028 (N_2028,In_297,In_659);
and U2029 (N_2029,In_729,In_51);
nand U2030 (N_2030,In_681,In_629);
nand U2031 (N_2031,In_387,In_159);
nand U2032 (N_2032,In_615,In_87);
or U2033 (N_2033,In_355,In_467);
nor U2034 (N_2034,In_525,In_536);
nand U2035 (N_2035,In_494,In_78);
or U2036 (N_2036,In_116,In_284);
or U2037 (N_2037,In_214,In_584);
nor U2038 (N_2038,In_539,In_448);
nor U2039 (N_2039,In_335,In_186);
and U2040 (N_2040,In_700,In_615);
and U2041 (N_2041,In_145,In_326);
nor U2042 (N_2042,In_589,In_356);
or U2043 (N_2043,In_328,In_537);
nand U2044 (N_2044,In_283,In_382);
nand U2045 (N_2045,In_358,In_558);
and U2046 (N_2046,In_503,In_455);
or U2047 (N_2047,In_122,In_664);
nor U2048 (N_2048,In_732,In_619);
and U2049 (N_2049,In_499,In_554);
and U2050 (N_2050,In_104,In_311);
and U2051 (N_2051,In_598,In_645);
and U2052 (N_2052,In_125,In_504);
nor U2053 (N_2053,In_332,In_309);
or U2054 (N_2054,In_632,In_287);
or U2055 (N_2055,In_719,In_304);
xor U2056 (N_2056,In_310,In_698);
nor U2057 (N_2057,In_29,In_673);
or U2058 (N_2058,In_506,In_373);
and U2059 (N_2059,In_248,In_297);
or U2060 (N_2060,In_9,In_586);
nand U2061 (N_2061,In_282,In_338);
xor U2062 (N_2062,In_442,In_580);
or U2063 (N_2063,In_25,In_721);
xor U2064 (N_2064,In_548,In_516);
nand U2065 (N_2065,In_743,In_218);
nor U2066 (N_2066,In_190,In_245);
or U2067 (N_2067,In_467,In_627);
or U2068 (N_2068,In_647,In_731);
and U2069 (N_2069,In_167,In_575);
xor U2070 (N_2070,In_256,In_306);
xnor U2071 (N_2071,In_706,In_396);
or U2072 (N_2072,In_497,In_76);
and U2073 (N_2073,In_367,In_293);
xor U2074 (N_2074,In_538,In_733);
nor U2075 (N_2075,In_117,In_548);
nor U2076 (N_2076,In_231,In_596);
or U2077 (N_2077,In_90,In_712);
nand U2078 (N_2078,In_645,In_688);
nor U2079 (N_2079,In_748,In_701);
nor U2080 (N_2080,In_626,In_590);
nor U2081 (N_2081,In_177,In_2);
and U2082 (N_2082,In_568,In_738);
nand U2083 (N_2083,In_587,In_250);
xor U2084 (N_2084,In_372,In_72);
or U2085 (N_2085,In_266,In_455);
xnor U2086 (N_2086,In_672,In_363);
nor U2087 (N_2087,In_257,In_150);
nand U2088 (N_2088,In_531,In_450);
xnor U2089 (N_2089,In_397,In_659);
nor U2090 (N_2090,In_210,In_473);
nand U2091 (N_2091,In_159,In_347);
and U2092 (N_2092,In_101,In_318);
nor U2093 (N_2093,In_227,In_716);
nor U2094 (N_2094,In_663,In_648);
nand U2095 (N_2095,In_655,In_590);
nand U2096 (N_2096,In_256,In_3);
xor U2097 (N_2097,In_561,In_126);
nor U2098 (N_2098,In_537,In_618);
or U2099 (N_2099,In_504,In_34);
nor U2100 (N_2100,In_688,In_660);
and U2101 (N_2101,In_527,In_465);
nor U2102 (N_2102,In_53,In_671);
and U2103 (N_2103,In_465,In_492);
xor U2104 (N_2104,In_594,In_584);
xor U2105 (N_2105,In_67,In_26);
nor U2106 (N_2106,In_97,In_471);
nand U2107 (N_2107,In_664,In_334);
xnor U2108 (N_2108,In_460,In_565);
and U2109 (N_2109,In_502,In_622);
nand U2110 (N_2110,In_188,In_728);
or U2111 (N_2111,In_489,In_66);
xnor U2112 (N_2112,In_307,In_471);
and U2113 (N_2113,In_352,In_1);
or U2114 (N_2114,In_459,In_247);
xor U2115 (N_2115,In_320,In_625);
or U2116 (N_2116,In_423,In_616);
and U2117 (N_2117,In_412,In_396);
nor U2118 (N_2118,In_185,In_450);
xor U2119 (N_2119,In_107,In_349);
nand U2120 (N_2120,In_340,In_62);
and U2121 (N_2121,In_71,In_230);
nand U2122 (N_2122,In_606,In_542);
xor U2123 (N_2123,In_465,In_404);
nand U2124 (N_2124,In_166,In_457);
nand U2125 (N_2125,In_124,In_62);
or U2126 (N_2126,In_289,In_610);
and U2127 (N_2127,In_354,In_453);
or U2128 (N_2128,In_649,In_459);
or U2129 (N_2129,In_79,In_99);
nand U2130 (N_2130,In_354,In_721);
or U2131 (N_2131,In_330,In_150);
nand U2132 (N_2132,In_46,In_454);
and U2133 (N_2133,In_606,In_744);
xnor U2134 (N_2134,In_717,In_454);
nand U2135 (N_2135,In_213,In_418);
and U2136 (N_2136,In_716,In_688);
nor U2137 (N_2137,In_430,In_79);
and U2138 (N_2138,In_495,In_353);
nand U2139 (N_2139,In_484,In_640);
or U2140 (N_2140,In_22,In_573);
nand U2141 (N_2141,In_612,In_2);
and U2142 (N_2142,In_222,In_108);
or U2143 (N_2143,In_133,In_566);
nand U2144 (N_2144,In_70,In_435);
nand U2145 (N_2145,In_702,In_358);
and U2146 (N_2146,In_448,In_728);
nand U2147 (N_2147,In_553,In_520);
and U2148 (N_2148,In_10,In_540);
or U2149 (N_2149,In_670,In_326);
nand U2150 (N_2150,In_203,In_601);
and U2151 (N_2151,In_457,In_7);
nor U2152 (N_2152,In_678,In_231);
or U2153 (N_2153,In_615,In_618);
xor U2154 (N_2154,In_75,In_63);
nor U2155 (N_2155,In_478,In_35);
xor U2156 (N_2156,In_617,In_27);
or U2157 (N_2157,In_685,In_247);
nand U2158 (N_2158,In_510,In_629);
xnor U2159 (N_2159,In_234,In_401);
nor U2160 (N_2160,In_170,In_489);
nor U2161 (N_2161,In_684,In_321);
xor U2162 (N_2162,In_512,In_566);
and U2163 (N_2163,In_108,In_478);
nor U2164 (N_2164,In_699,In_733);
xnor U2165 (N_2165,In_606,In_428);
nor U2166 (N_2166,In_293,In_689);
nor U2167 (N_2167,In_425,In_321);
xor U2168 (N_2168,In_104,In_744);
or U2169 (N_2169,In_469,In_735);
xor U2170 (N_2170,In_249,In_115);
xor U2171 (N_2171,In_468,In_610);
nor U2172 (N_2172,In_251,In_572);
nand U2173 (N_2173,In_317,In_514);
xnor U2174 (N_2174,In_399,In_336);
xor U2175 (N_2175,In_105,In_641);
nor U2176 (N_2176,In_0,In_518);
or U2177 (N_2177,In_397,In_299);
nor U2178 (N_2178,In_494,In_645);
and U2179 (N_2179,In_409,In_429);
nand U2180 (N_2180,In_719,In_17);
and U2181 (N_2181,In_708,In_362);
nor U2182 (N_2182,In_617,In_147);
and U2183 (N_2183,In_19,In_379);
nor U2184 (N_2184,In_470,In_369);
xor U2185 (N_2185,In_410,In_515);
nand U2186 (N_2186,In_314,In_42);
nor U2187 (N_2187,In_426,In_243);
nand U2188 (N_2188,In_187,In_655);
nor U2189 (N_2189,In_469,In_293);
xnor U2190 (N_2190,In_408,In_306);
and U2191 (N_2191,In_457,In_728);
nor U2192 (N_2192,In_316,In_589);
nand U2193 (N_2193,In_530,In_377);
and U2194 (N_2194,In_215,In_232);
and U2195 (N_2195,In_31,In_364);
xor U2196 (N_2196,In_53,In_252);
or U2197 (N_2197,In_397,In_159);
nor U2198 (N_2198,In_62,In_206);
xor U2199 (N_2199,In_606,In_372);
or U2200 (N_2200,In_447,In_386);
nand U2201 (N_2201,In_412,In_256);
and U2202 (N_2202,In_417,In_371);
nand U2203 (N_2203,In_599,In_719);
xnor U2204 (N_2204,In_461,In_619);
nor U2205 (N_2205,In_467,In_701);
or U2206 (N_2206,In_238,In_103);
nand U2207 (N_2207,In_103,In_167);
xor U2208 (N_2208,In_201,In_596);
or U2209 (N_2209,In_296,In_707);
xnor U2210 (N_2210,In_719,In_592);
nand U2211 (N_2211,In_9,In_347);
nand U2212 (N_2212,In_370,In_652);
and U2213 (N_2213,In_543,In_331);
or U2214 (N_2214,In_179,In_89);
nand U2215 (N_2215,In_305,In_25);
and U2216 (N_2216,In_78,In_26);
nor U2217 (N_2217,In_381,In_374);
and U2218 (N_2218,In_545,In_268);
and U2219 (N_2219,In_64,In_90);
xnor U2220 (N_2220,In_705,In_426);
nand U2221 (N_2221,In_126,In_221);
nand U2222 (N_2222,In_377,In_36);
and U2223 (N_2223,In_66,In_536);
or U2224 (N_2224,In_145,In_155);
nor U2225 (N_2225,In_220,In_695);
xor U2226 (N_2226,In_36,In_105);
and U2227 (N_2227,In_606,In_148);
xnor U2228 (N_2228,In_562,In_589);
or U2229 (N_2229,In_492,In_304);
or U2230 (N_2230,In_523,In_22);
nand U2231 (N_2231,In_167,In_53);
and U2232 (N_2232,In_252,In_24);
or U2233 (N_2233,In_304,In_44);
xnor U2234 (N_2234,In_531,In_726);
nand U2235 (N_2235,In_408,In_393);
xor U2236 (N_2236,In_99,In_404);
nor U2237 (N_2237,In_227,In_552);
xor U2238 (N_2238,In_287,In_212);
nand U2239 (N_2239,In_295,In_152);
nand U2240 (N_2240,In_522,In_569);
nand U2241 (N_2241,In_14,In_326);
and U2242 (N_2242,In_304,In_131);
nand U2243 (N_2243,In_117,In_269);
or U2244 (N_2244,In_369,In_266);
nand U2245 (N_2245,In_559,In_149);
nand U2246 (N_2246,In_289,In_508);
nor U2247 (N_2247,In_669,In_158);
and U2248 (N_2248,In_509,In_567);
and U2249 (N_2249,In_220,In_391);
or U2250 (N_2250,In_674,In_582);
nand U2251 (N_2251,In_101,In_257);
xor U2252 (N_2252,In_599,In_570);
or U2253 (N_2253,In_14,In_115);
nor U2254 (N_2254,In_544,In_222);
nand U2255 (N_2255,In_284,In_705);
xor U2256 (N_2256,In_604,In_419);
nor U2257 (N_2257,In_512,In_142);
nand U2258 (N_2258,In_482,In_741);
and U2259 (N_2259,In_33,In_432);
nand U2260 (N_2260,In_662,In_699);
nand U2261 (N_2261,In_26,In_135);
xor U2262 (N_2262,In_133,In_266);
and U2263 (N_2263,In_727,In_312);
xor U2264 (N_2264,In_194,In_305);
and U2265 (N_2265,In_565,In_478);
xnor U2266 (N_2266,In_314,In_218);
or U2267 (N_2267,In_497,In_372);
or U2268 (N_2268,In_738,In_169);
xnor U2269 (N_2269,In_238,In_545);
nor U2270 (N_2270,In_229,In_475);
nor U2271 (N_2271,In_75,In_739);
nor U2272 (N_2272,In_398,In_260);
or U2273 (N_2273,In_523,In_534);
nand U2274 (N_2274,In_355,In_327);
nand U2275 (N_2275,In_502,In_675);
nand U2276 (N_2276,In_741,In_81);
xnor U2277 (N_2277,In_212,In_223);
xor U2278 (N_2278,In_682,In_97);
nor U2279 (N_2279,In_637,In_48);
nor U2280 (N_2280,In_59,In_339);
xnor U2281 (N_2281,In_145,In_188);
and U2282 (N_2282,In_108,In_330);
and U2283 (N_2283,In_422,In_281);
and U2284 (N_2284,In_237,In_639);
or U2285 (N_2285,In_358,In_708);
or U2286 (N_2286,In_499,In_449);
nor U2287 (N_2287,In_525,In_523);
xnor U2288 (N_2288,In_49,In_683);
or U2289 (N_2289,In_592,In_478);
nor U2290 (N_2290,In_320,In_310);
and U2291 (N_2291,In_221,In_46);
nor U2292 (N_2292,In_474,In_17);
nor U2293 (N_2293,In_364,In_658);
nor U2294 (N_2294,In_711,In_132);
nor U2295 (N_2295,In_306,In_197);
nor U2296 (N_2296,In_144,In_82);
nand U2297 (N_2297,In_38,In_424);
nor U2298 (N_2298,In_46,In_25);
nand U2299 (N_2299,In_395,In_443);
nor U2300 (N_2300,In_300,In_201);
xnor U2301 (N_2301,In_736,In_715);
nand U2302 (N_2302,In_690,In_597);
nor U2303 (N_2303,In_152,In_488);
nand U2304 (N_2304,In_311,In_182);
and U2305 (N_2305,In_414,In_495);
xor U2306 (N_2306,In_183,In_304);
nand U2307 (N_2307,In_515,In_678);
xnor U2308 (N_2308,In_93,In_748);
nor U2309 (N_2309,In_618,In_381);
and U2310 (N_2310,In_570,In_527);
xnor U2311 (N_2311,In_544,In_555);
or U2312 (N_2312,In_637,In_448);
nor U2313 (N_2313,In_595,In_424);
nor U2314 (N_2314,In_404,In_172);
or U2315 (N_2315,In_705,In_74);
xor U2316 (N_2316,In_642,In_537);
or U2317 (N_2317,In_542,In_395);
nor U2318 (N_2318,In_328,In_485);
xnor U2319 (N_2319,In_443,In_441);
nor U2320 (N_2320,In_686,In_146);
xor U2321 (N_2321,In_112,In_157);
nand U2322 (N_2322,In_166,In_83);
or U2323 (N_2323,In_479,In_552);
xor U2324 (N_2324,In_124,In_471);
and U2325 (N_2325,In_127,In_554);
and U2326 (N_2326,In_48,In_625);
nor U2327 (N_2327,In_652,In_397);
nand U2328 (N_2328,In_694,In_319);
and U2329 (N_2329,In_442,In_713);
and U2330 (N_2330,In_257,In_669);
and U2331 (N_2331,In_611,In_19);
xnor U2332 (N_2332,In_505,In_277);
nor U2333 (N_2333,In_389,In_597);
nor U2334 (N_2334,In_35,In_207);
nor U2335 (N_2335,In_655,In_387);
nand U2336 (N_2336,In_722,In_524);
or U2337 (N_2337,In_221,In_459);
nor U2338 (N_2338,In_31,In_699);
nand U2339 (N_2339,In_341,In_636);
or U2340 (N_2340,In_384,In_749);
nand U2341 (N_2341,In_495,In_465);
nand U2342 (N_2342,In_346,In_341);
nor U2343 (N_2343,In_590,In_325);
xnor U2344 (N_2344,In_638,In_725);
xnor U2345 (N_2345,In_568,In_651);
nand U2346 (N_2346,In_440,In_739);
nor U2347 (N_2347,In_506,In_127);
or U2348 (N_2348,In_330,In_384);
nand U2349 (N_2349,In_310,In_490);
or U2350 (N_2350,In_441,In_170);
and U2351 (N_2351,In_444,In_222);
xnor U2352 (N_2352,In_641,In_469);
nor U2353 (N_2353,In_350,In_194);
or U2354 (N_2354,In_640,In_63);
nand U2355 (N_2355,In_80,In_369);
nor U2356 (N_2356,In_110,In_619);
or U2357 (N_2357,In_416,In_85);
nand U2358 (N_2358,In_707,In_263);
nand U2359 (N_2359,In_219,In_22);
and U2360 (N_2360,In_24,In_204);
nor U2361 (N_2361,In_731,In_327);
nand U2362 (N_2362,In_725,In_561);
xnor U2363 (N_2363,In_731,In_584);
nand U2364 (N_2364,In_737,In_252);
nor U2365 (N_2365,In_283,In_399);
xnor U2366 (N_2366,In_636,In_621);
nor U2367 (N_2367,In_676,In_539);
nand U2368 (N_2368,In_622,In_571);
nor U2369 (N_2369,In_46,In_616);
nor U2370 (N_2370,In_534,In_299);
and U2371 (N_2371,In_307,In_251);
or U2372 (N_2372,In_349,In_559);
nand U2373 (N_2373,In_632,In_329);
nor U2374 (N_2374,In_128,In_59);
nand U2375 (N_2375,In_249,In_274);
nand U2376 (N_2376,In_63,In_10);
and U2377 (N_2377,In_478,In_129);
and U2378 (N_2378,In_119,In_577);
nand U2379 (N_2379,In_460,In_213);
nor U2380 (N_2380,In_468,In_394);
nor U2381 (N_2381,In_216,In_514);
xnor U2382 (N_2382,In_696,In_565);
xor U2383 (N_2383,In_559,In_6);
or U2384 (N_2384,In_477,In_174);
nor U2385 (N_2385,In_342,In_268);
nand U2386 (N_2386,In_567,In_586);
nand U2387 (N_2387,In_73,In_682);
and U2388 (N_2388,In_239,In_227);
and U2389 (N_2389,In_508,In_243);
and U2390 (N_2390,In_356,In_432);
and U2391 (N_2391,In_365,In_676);
or U2392 (N_2392,In_513,In_502);
and U2393 (N_2393,In_206,In_331);
xor U2394 (N_2394,In_354,In_1);
xor U2395 (N_2395,In_199,In_512);
nand U2396 (N_2396,In_253,In_200);
or U2397 (N_2397,In_392,In_197);
or U2398 (N_2398,In_142,In_592);
nand U2399 (N_2399,In_211,In_150);
nand U2400 (N_2400,In_501,In_613);
or U2401 (N_2401,In_546,In_41);
xor U2402 (N_2402,In_73,In_59);
xor U2403 (N_2403,In_242,In_376);
or U2404 (N_2404,In_248,In_70);
nand U2405 (N_2405,In_590,In_485);
nand U2406 (N_2406,In_26,In_529);
nor U2407 (N_2407,In_411,In_167);
nand U2408 (N_2408,In_700,In_292);
xor U2409 (N_2409,In_108,In_553);
and U2410 (N_2410,In_236,In_689);
nand U2411 (N_2411,In_174,In_296);
nand U2412 (N_2412,In_31,In_621);
nand U2413 (N_2413,In_105,In_156);
xor U2414 (N_2414,In_304,In_313);
nor U2415 (N_2415,In_572,In_723);
xnor U2416 (N_2416,In_146,In_702);
nand U2417 (N_2417,In_323,In_237);
or U2418 (N_2418,In_446,In_19);
nor U2419 (N_2419,In_343,In_147);
or U2420 (N_2420,In_217,In_558);
nor U2421 (N_2421,In_150,In_454);
nand U2422 (N_2422,In_460,In_557);
nor U2423 (N_2423,In_257,In_524);
nand U2424 (N_2424,In_184,In_522);
or U2425 (N_2425,In_59,In_429);
nand U2426 (N_2426,In_183,In_726);
and U2427 (N_2427,In_220,In_701);
nor U2428 (N_2428,In_456,In_552);
or U2429 (N_2429,In_531,In_655);
xor U2430 (N_2430,In_102,In_174);
nand U2431 (N_2431,In_293,In_534);
nand U2432 (N_2432,In_416,In_631);
and U2433 (N_2433,In_638,In_633);
xor U2434 (N_2434,In_33,In_713);
nand U2435 (N_2435,In_636,In_357);
nand U2436 (N_2436,In_193,In_663);
nand U2437 (N_2437,In_199,In_551);
or U2438 (N_2438,In_105,In_447);
xor U2439 (N_2439,In_470,In_329);
nand U2440 (N_2440,In_93,In_562);
or U2441 (N_2441,In_462,In_630);
and U2442 (N_2442,In_30,In_39);
xor U2443 (N_2443,In_31,In_0);
nand U2444 (N_2444,In_724,In_431);
nand U2445 (N_2445,In_407,In_314);
nand U2446 (N_2446,In_696,In_360);
nand U2447 (N_2447,In_111,In_416);
nor U2448 (N_2448,In_536,In_143);
nand U2449 (N_2449,In_601,In_84);
and U2450 (N_2450,In_284,In_122);
and U2451 (N_2451,In_11,In_258);
nor U2452 (N_2452,In_679,In_644);
or U2453 (N_2453,In_645,In_214);
or U2454 (N_2454,In_623,In_46);
or U2455 (N_2455,In_628,In_15);
nand U2456 (N_2456,In_365,In_66);
nor U2457 (N_2457,In_49,In_58);
and U2458 (N_2458,In_514,In_347);
or U2459 (N_2459,In_711,In_527);
xnor U2460 (N_2460,In_143,In_96);
nor U2461 (N_2461,In_237,In_162);
or U2462 (N_2462,In_408,In_78);
or U2463 (N_2463,In_102,In_592);
nand U2464 (N_2464,In_288,In_147);
or U2465 (N_2465,In_665,In_16);
xor U2466 (N_2466,In_544,In_204);
or U2467 (N_2467,In_11,In_422);
nor U2468 (N_2468,In_75,In_623);
and U2469 (N_2469,In_31,In_321);
and U2470 (N_2470,In_488,In_217);
or U2471 (N_2471,In_157,In_460);
and U2472 (N_2472,In_296,In_595);
xnor U2473 (N_2473,In_519,In_211);
nor U2474 (N_2474,In_240,In_227);
nor U2475 (N_2475,In_471,In_526);
nor U2476 (N_2476,In_347,In_493);
or U2477 (N_2477,In_70,In_338);
and U2478 (N_2478,In_438,In_201);
nand U2479 (N_2479,In_294,In_136);
or U2480 (N_2480,In_148,In_425);
nor U2481 (N_2481,In_397,In_421);
or U2482 (N_2482,In_24,In_600);
or U2483 (N_2483,In_201,In_462);
xor U2484 (N_2484,In_481,In_420);
or U2485 (N_2485,In_547,In_481);
and U2486 (N_2486,In_643,In_206);
nor U2487 (N_2487,In_513,In_663);
and U2488 (N_2488,In_156,In_245);
and U2489 (N_2489,In_42,In_325);
nand U2490 (N_2490,In_279,In_88);
nor U2491 (N_2491,In_146,In_305);
and U2492 (N_2492,In_480,In_534);
xnor U2493 (N_2493,In_360,In_461);
or U2494 (N_2494,In_414,In_443);
and U2495 (N_2495,In_276,In_325);
xnor U2496 (N_2496,In_502,In_215);
nor U2497 (N_2497,In_739,In_459);
nand U2498 (N_2498,In_174,In_103);
nand U2499 (N_2499,In_282,In_703);
nand U2500 (N_2500,N_293,N_1616);
nand U2501 (N_2501,N_478,N_2404);
xor U2502 (N_2502,N_848,N_1921);
nand U2503 (N_2503,N_1061,N_509);
and U2504 (N_2504,N_2191,N_1947);
and U2505 (N_2505,N_2115,N_82);
or U2506 (N_2506,N_1938,N_2302);
nor U2507 (N_2507,N_500,N_323);
nor U2508 (N_2508,N_1309,N_667);
or U2509 (N_2509,N_1101,N_1467);
nor U2510 (N_2510,N_391,N_2132);
nor U2511 (N_2511,N_1991,N_1338);
and U2512 (N_2512,N_1943,N_1385);
nand U2513 (N_2513,N_1151,N_1202);
nand U2514 (N_2514,N_2300,N_1303);
xor U2515 (N_2515,N_1875,N_2279);
xor U2516 (N_2516,N_1416,N_2079);
nand U2517 (N_2517,N_2004,N_370);
nand U2518 (N_2518,N_1756,N_829);
nand U2519 (N_2519,N_807,N_1482);
or U2520 (N_2520,N_2495,N_1659);
nand U2521 (N_2521,N_78,N_2261);
xnor U2522 (N_2522,N_46,N_277);
and U2523 (N_2523,N_2246,N_2036);
and U2524 (N_2524,N_1314,N_2110);
or U2525 (N_2525,N_56,N_2044);
and U2526 (N_2526,N_115,N_719);
and U2527 (N_2527,N_275,N_1236);
and U2528 (N_2528,N_1284,N_642);
or U2529 (N_2529,N_709,N_746);
nor U2530 (N_2530,N_104,N_1026);
or U2531 (N_2531,N_1739,N_862);
and U2532 (N_2532,N_1665,N_1924);
nand U2533 (N_2533,N_2170,N_577);
and U2534 (N_2534,N_1644,N_2135);
or U2535 (N_2535,N_2193,N_269);
and U2536 (N_2536,N_1941,N_2217);
nand U2537 (N_2537,N_1071,N_1187);
nand U2538 (N_2538,N_1152,N_1724);
and U2539 (N_2539,N_1751,N_346);
nand U2540 (N_2540,N_805,N_1598);
and U2541 (N_2541,N_2321,N_700);
or U2542 (N_2542,N_1046,N_1534);
nor U2543 (N_2543,N_295,N_1400);
or U2544 (N_2544,N_303,N_936);
xnor U2545 (N_2545,N_716,N_1851);
nand U2546 (N_2546,N_237,N_555);
nand U2547 (N_2547,N_2424,N_59);
xnor U2548 (N_2548,N_2209,N_2165);
or U2549 (N_2549,N_2204,N_1181);
nor U2550 (N_2550,N_1406,N_224);
nand U2551 (N_2551,N_1411,N_1402);
xnor U2552 (N_2552,N_1819,N_1683);
or U2553 (N_2553,N_145,N_1239);
or U2554 (N_2554,N_2050,N_2011);
nand U2555 (N_2555,N_1953,N_1667);
and U2556 (N_2556,N_502,N_2393);
and U2557 (N_2557,N_148,N_1126);
xor U2558 (N_2558,N_904,N_36);
or U2559 (N_2559,N_388,N_521);
nand U2560 (N_2560,N_2453,N_2155);
nand U2561 (N_2561,N_192,N_2144);
xnor U2562 (N_2562,N_1701,N_1716);
or U2563 (N_2563,N_1237,N_2466);
or U2564 (N_2564,N_2130,N_1240);
nand U2565 (N_2565,N_909,N_479);
xor U2566 (N_2566,N_1632,N_567);
nand U2567 (N_2567,N_1618,N_1717);
or U2568 (N_2568,N_200,N_2277);
nand U2569 (N_2569,N_21,N_390);
or U2570 (N_2570,N_2356,N_1143);
and U2571 (N_2571,N_621,N_1049);
and U2572 (N_2572,N_1356,N_1353);
nand U2573 (N_2573,N_125,N_1355);
xor U2574 (N_2574,N_216,N_1347);
and U2575 (N_2575,N_445,N_619);
nand U2576 (N_2576,N_2381,N_2377);
nand U2577 (N_2577,N_1317,N_1579);
and U2578 (N_2578,N_1144,N_1692);
nor U2579 (N_2579,N_15,N_1937);
nand U2580 (N_2580,N_1611,N_2203);
nor U2581 (N_2581,N_332,N_1700);
and U2582 (N_2582,N_434,N_1377);
nand U2583 (N_2583,N_1562,N_874);
nand U2584 (N_2584,N_414,N_2208);
xnor U2585 (N_2585,N_2387,N_331);
nand U2586 (N_2586,N_832,N_1379);
nand U2587 (N_2587,N_261,N_1962);
or U2588 (N_2588,N_289,N_1639);
and U2589 (N_2589,N_2497,N_1981);
or U2590 (N_2590,N_1384,N_1858);
nand U2591 (N_2591,N_2270,N_671);
nand U2592 (N_2592,N_1863,N_1220);
nor U2593 (N_2593,N_1271,N_534);
or U2594 (N_2594,N_1620,N_2197);
and U2595 (N_2595,N_1653,N_622);
and U2596 (N_2596,N_1262,N_30);
nand U2597 (N_2597,N_219,N_325);
or U2598 (N_2598,N_206,N_1276);
nor U2599 (N_2599,N_1588,N_67);
nand U2600 (N_2600,N_1758,N_1925);
xnor U2601 (N_2601,N_7,N_236);
xnor U2602 (N_2602,N_1580,N_1612);
nor U2603 (N_2603,N_1154,N_1081);
and U2604 (N_2604,N_92,N_2425);
or U2605 (N_2605,N_1866,N_260);
nor U2606 (N_2606,N_2026,N_1902);
and U2607 (N_2607,N_288,N_1440);
and U2608 (N_2608,N_2375,N_1749);
or U2609 (N_2609,N_1329,N_801);
and U2610 (N_2610,N_150,N_959);
xor U2611 (N_2611,N_2491,N_2337);
nor U2612 (N_2612,N_788,N_1547);
xnor U2613 (N_2613,N_785,N_302);
nand U2614 (N_2614,N_1939,N_993);
nand U2615 (N_2615,N_230,N_396);
nor U2616 (N_2616,N_8,N_1231);
or U2617 (N_2617,N_2299,N_94);
nor U2618 (N_2618,N_2329,N_1668);
and U2619 (N_2619,N_1483,N_2174);
or U2620 (N_2620,N_1374,N_871);
and U2621 (N_2621,N_490,N_547);
and U2622 (N_2622,N_1072,N_1854);
and U2623 (N_2623,N_2370,N_2462);
nor U2624 (N_2624,N_2061,N_2219);
and U2625 (N_2625,N_2126,N_3);
or U2626 (N_2626,N_854,N_468);
or U2627 (N_2627,N_605,N_1058);
or U2628 (N_2628,N_2484,N_404);
and U2629 (N_2629,N_1104,N_2233);
xor U2630 (N_2630,N_1980,N_2463);
xnor U2631 (N_2631,N_1967,N_2474);
nor U2632 (N_2632,N_2196,N_307);
and U2633 (N_2633,N_1032,N_930);
nand U2634 (N_2634,N_1387,N_1090);
nand U2635 (N_2635,N_2345,N_1292);
nand U2636 (N_2636,N_609,N_839);
and U2637 (N_2637,N_637,N_533);
and U2638 (N_2638,N_1559,N_470);
or U2639 (N_2639,N_556,N_428);
or U2640 (N_2640,N_2017,N_751);
nor U2641 (N_2641,N_935,N_1556);
nor U2642 (N_2642,N_1435,N_2091);
xor U2643 (N_2643,N_377,N_1209);
xnor U2644 (N_2644,N_301,N_2069);
xor U2645 (N_2645,N_1843,N_2290);
nor U2646 (N_2646,N_1363,N_1246);
nand U2647 (N_2647,N_2432,N_2060);
or U2648 (N_2648,N_727,N_2365);
and U2649 (N_2649,N_1578,N_2301);
and U2650 (N_2650,N_1555,N_382);
nor U2651 (N_2651,N_763,N_941);
and U2652 (N_2652,N_1987,N_652);
and U2653 (N_2653,N_342,N_744);
nor U2654 (N_2654,N_2210,N_2023);
xnor U2655 (N_2655,N_1802,N_672);
xor U2656 (N_2656,N_1272,N_1219);
or U2657 (N_2657,N_1218,N_1465);
nor U2658 (N_2658,N_83,N_2222);
xor U2659 (N_2659,N_1684,N_1872);
and U2660 (N_2660,N_1336,N_1456);
and U2661 (N_2661,N_2092,N_1931);
and U2662 (N_2662,N_1162,N_157);
nand U2663 (N_2663,N_1063,N_187);
or U2664 (N_2664,N_484,N_863);
xnor U2665 (N_2665,N_897,N_2105);
and U2666 (N_2666,N_866,N_2189);
nand U2667 (N_2667,N_1381,N_1059);
nor U2668 (N_2668,N_2131,N_398);
nand U2669 (N_2669,N_314,N_531);
and U2670 (N_2670,N_2447,N_1122);
or U2671 (N_2671,N_1901,N_475);
xor U2672 (N_2672,N_1983,N_724);
and U2673 (N_2673,N_1771,N_90);
nor U2674 (N_2674,N_1422,N_778);
and U2675 (N_2675,N_895,N_461);
xnor U2676 (N_2676,N_1666,N_513);
xnor U2677 (N_2677,N_877,N_2228);
or U2678 (N_2678,N_1608,N_1321);
and U2679 (N_2679,N_2326,N_933);
or U2680 (N_2680,N_2402,N_2035);
and U2681 (N_2681,N_1737,N_582);
and U2682 (N_2682,N_195,N_1473);
nor U2683 (N_2683,N_251,N_110);
or U2684 (N_2684,N_139,N_334);
nand U2685 (N_2685,N_1573,N_1222);
or U2686 (N_2686,N_74,N_2499);
nand U2687 (N_2687,N_433,N_655);
xnor U2688 (N_2688,N_1848,N_519);
nand U2689 (N_2689,N_2033,N_629);
and U2690 (N_2690,N_227,N_2243);
nand U2691 (N_2691,N_1429,N_2494);
nor U2692 (N_2692,N_628,N_2423);
and U2693 (N_2693,N_1341,N_907);
or U2694 (N_2694,N_2320,N_204);
or U2695 (N_2695,N_100,N_810);
nand U2696 (N_2696,N_123,N_1935);
xnor U2697 (N_2697,N_339,N_2258);
nor U2698 (N_2698,N_732,N_1265);
nor U2699 (N_2699,N_77,N_198);
and U2700 (N_2700,N_818,N_1775);
nor U2701 (N_2701,N_830,N_2363);
xor U2702 (N_2702,N_1092,N_1793);
and U2703 (N_2703,N_2224,N_645);
or U2704 (N_2704,N_1076,N_1164);
nand U2705 (N_2705,N_387,N_633);
or U2706 (N_2706,N_1805,N_715);
and U2707 (N_2707,N_765,N_2392);
nand U2708 (N_2708,N_1114,N_313);
or U2709 (N_2709,N_872,N_287);
xnor U2710 (N_2710,N_202,N_352);
xor U2711 (N_2711,N_823,N_962);
xnor U2712 (N_2712,N_2444,N_472);
nor U2713 (N_2713,N_1337,N_117);
nand U2714 (N_2714,N_559,N_2291);
and U2715 (N_2715,N_774,N_2239);
nor U2716 (N_2716,N_57,N_2124);
and U2717 (N_2717,N_1631,N_229);
nor U2718 (N_2718,N_1965,N_193);
xor U2719 (N_2719,N_26,N_2469);
xnor U2720 (N_2720,N_1677,N_498);
nor U2721 (N_2721,N_1936,N_2010);
xnor U2722 (N_2722,N_2134,N_2293);
xor U2723 (N_2723,N_2051,N_1105);
and U2724 (N_2724,N_349,N_2448);
nand U2725 (N_2725,N_789,N_1776);
nor U2726 (N_2726,N_248,N_460);
or U2727 (N_2727,N_1954,N_1452);
and U2728 (N_2728,N_601,N_1089);
nor U2729 (N_2729,N_721,N_119);
or U2730 (N_2730,N_2351,N_838);
nand U2731 (N_2731,N_782,N_345);
and U2732 (N_2732,N_2112,N_1763);
and U2733 (N_2733,N_1755,N_730);
xor U2734 (N_2734,N_2238,N_1312);
nor U2735 (N_2735,N_1324,N_1157);
nand U2736 (N_2736,N_121,N_600);
and U2737 (N_2737,N_2223,N_38);
or U2738 (N_2738,N_1821,N_263);
xnor U2739 (N_2739,N_981,N_1177);
or U2740 (N_2740,N_2029,N_894);
nand U2741 (N_2741,N_1413,N_285);
or U2742 (N_2742,N_1955,N_958);
nand U2743 (N_2743,N_365,N_2169);
and U2744 (N_2744,N_634,N_2089);
nor U2745 (N_2745,N_1275,N_2236);
or U2746 (N_2746,N_1887,N_2213);
xor U2747 (N_2747,N_31,N_1548);
or U2748 (N_2748,N_143,N_1922);
nand U2749 (N_2749,N_1648,N_1487);
xor U2750 (N_2750,N_266,N_2156);
or U2751 (N_2751,N_108,N_1464);
xnor U2752 (N_2752,N_2158,N_430);
xor U2753 (N_2753,N_2085,N_2160);
nor U2754 (N_2754,N_944,N_977);
nor U2755 (N_2755,N_1917,N_16);
and U2756 (N_2756,N_568,N_1426);
nand U2757 (N_2757,N_1077,N_1801);
or U2758 (N_2758,N_1301,N_1358);
nor U2759 (N_2759,N_1185,N_201);
or U2760 (N_2760,N_477,N_913);
xor U2761 (N_2761,N_1886,N_1302);
and U2762 (N_2762,N_1070,N_174);
or U2763 (N_2763,N_1780,N_1223);
nor U2764 (N_2764,N_2355,N_713);
and U2765 (N_2765,N_358,N_1946);
or U2766 (N_2766,N_1360,N_598);
or U2767 (N_2767,N_1053,N_574);
nand U2768 (N_2768,N_1012,N_347);
and U2769 (N_2769,N_2308,N_2353);
nor U2770 (N_2770,N_2482,N_2489);
or U2771 (N_2771,N_1715,N_133);
nand U2772 (N_2772,N_1148,N_1690);
xor U2773 (N_2773,N_794,N_623);
nand U2774 (N_2774,N_28,N_2176);
xnor U2775 (N_2775,N_1028,N_1822);
and U2776 (N_2776,N_681,N_2366);
and U2777 (N_2777,N_1626,N_882);
and U2778 (N_2778,N_1335,N_2359);
nand U2779 (N_2779,N_2347,N_833);
or U2780 (N_2780,N_2218,N_1581);
nand U2781 (N_2781,N_1586,N_1551);
nand U2782 (N_2782,N_20,N_32);
and U2783 (N_2783,N_954,N_1718);
nor U2784 (N_2784,N_284,N_1785);
xnor U2785 (N_2785,N_60,N_1405);
or U2786 (N_2786,N_1136,N_2206);
xnor U2787 (N_2787,N_69,N_2161);
nand U2788 (N_2788,N_2098,N_2262);
nor U2789 (N_2789,N_890,N_1508);
nor U2790 (N_2790,N_247,N_617);
or U2791 (N_2791,N_1019,N_1740);
nand U2792 (N_2792,N_999,N_154);
nand U2793 (N_2793,N_2207,N_290);
nand U2794 (N_2794,N_421,N_2212);
or U2795 (N_2795,N_220,N_1361);
xor U2796 (N_2796,N_1257,N_2249);
xor U2797 (N_2797,N_4,N_1180);
nand U2798 (N_2798,N_1609,N_2350);
and U2799 (N_2799,N_1910,N_1307);
or U2800 (N_2800,N_1277,N_714);
nor U2801 (N_2801,N_1259,N_1876);
xnor U2802 (N_2802,N_523,N_1602);
xnor U2803 (N_2803,N_1830,N_2339);
or U2804 (N_2804,N_793,N_2150);
or U2805 (N_2805,N_1825,N_2412);
xnor U2806 (N_2806,N_1146,N_817);
or U2807 (N_2807,N_1582,N_1054);
and U2808 (N_2808,N_1037,N_80);
or U2809 (N_2809,N_1134,N_508);
and U2810 (N_2810,N_2431,N_581);
nor U2811 (N_2811,N_1959,N_243);
or U2812 (N_2812,N_1506,N_1787);
nand U2813 (N_2813,N_548,N_995);
or U2814 (N_2814,N_693,N_1795);
xor U2815 (N_2815,N_899,N_47);
xor U2816 (N_2816,N_997,N_2314);
nand U2817 (N_2817,N_2120,N_837);
nor U2818 (N_2818,N_367,N_903);
nor U2819 (N_2819,N_2030,N_134);
nor U2820 (N_2820,N_759,N_1643);
nor U2821 (N_2821,N_2162,N_2153);
nor U2822 (N_2822,N_2002,N_2014);
and U2823 (N_2823,N_2127,N_492);
and U2824 (N_2824,N_809,N_786);
nor U2825 (N_2825,N_1132,N_783);
or U2826 (N_2826,N_680,N_282);
nor U2827 (N_2827,N_1078,N_503);
xnor U2828 (N_2828,N_1509,N_122);
and U2829 (N_2829,N_1603,N_1888);
or U2830 (N_2830,N_530,N_1651);
xnor U2831 (N_2831,N_965,N_663);
and U2832 (N_2832,N_1884,N_665);
or U2833 (N_2833,N_1928,N_1810);
xor U2834 (N_2834,N_161,N_1100);
or U2835 (N_2835,N_221,N_297);
or U2836 (N_2836,N_1735,N_2226);
xor U2837 (N_2837,N_1367,N_2006);
xor U2838 (N_2838,N_1827,N_2216);
or U2839 (N_2839,N_87,N_1885);
nor U2840 (N_2840,N_1201,N_912);
and U2841 (N_2841,N_2455,N_2286);
nand U2842 (N_2842,N_983,N_169);
xnor U2843 (N_2843,N_2295,N_1907);
or U2844 (N_2844,N_846,N_1727);
nor U2845 (N_2845,N_1044,N_1682);
or U2846 (N_2846,N_1362,N_185);
nor U2847 (N_2847,N_1904,N_1705);
nand U2848 (N_2848,N_979,N_102);
nand U2849 (N_2849,N_180,N_2283);
xnor U2850 (N_2850,N_675,N_1905);
nand U2851 (N_2851,N_939,N_666);
or U2852 (N_2852,N_550,N_1045);
nand U2853 (N_2853,N_405,N_79);
nand U2854 (N_2854,N_61,N_1807);
nand U2855 (N_2855,N_1899,N_613);
and U2856 (N_2856,N_2182,N_673);
xnor U2857 (N_2857,N_366,N_1158);
nor U2858 (N_2858,N_1485,N_480);
xnor U2859 (N_2859,N_552,N_1194);
nand U2860 (N_2860,N_773,N_733);
and U2861 (N_2861,N_2009,N_1828);
or U2862 (N_2862,N_971,N_1798);
nand U2863 (N_2863,N_760,N_1592);
nand U2864 (N_2864,N_1867,N_1641);
xnor U2865 (N_2865,N_1438,N_1544);
or U2866 (N_2866,N_964,N_940);
xnor U2867 (N_2867,N_1649,N_1330);
nand U2868 (N_2868,N_1129,N_1784);
nand U2869 (N_2869,N_880,N_1062);
nor U2870 (N_2870,N_2485,N_397);
nand U2871 (N_2871,N_2486,N_1777);
nor U2872 (N_2872,N_902,N_780);
and U2873 (N_2873,N_11,N_2056);
nand U2874 (N_2874,N_1661,N_1929);
nor U2875 (N_2875,N_1961,N_2405);
nand U2876 (N_2876,N_708,N_640);
nor U2877 (N_2877,N_113,N_1210);
nand U2878 (N_2878,N_987,N_869);
nor U2879 (N_2879,N_1165,N_2341);
nand U2880 (N_2880,N_1514,N_1537);
and U2881 (N_2881,N_1192,N_1001);
or U2882 (N_2882,N_2067,N_931);
or U2883 (N_2883,N_624,N_1428);
or U2884 (N_2884,N_2260,N_636);
nor U2885 (N_2885,N_511,N_368);
xor U2886 (N_2886,N_1765,N_643);
nand U2887 (N_2887,N_1283,N_611);
and U2888 (N_2888,N_1671,N_542);
nand U2889 (N_2889,N_2214,N_1532);
xor U2890 (N_2890,N_1820,N_2016);
xor U2891 (N_2891,N_1593,N_2096);
nor U2892 (N_2892,N_2235,N_2330);
nand U2893 (N_2893,N_2244,N_1110);
or U2894 (N_2894,N_2118,N_710);
or U2895 (N_2895,N_35,N_2241);
xor U2896 (N_2896,N_1920,N_85);
nor U2897 (N_2897,N_1849,N_5);
nor U2898 (N_2898,N_1856,N_2177);
or U2899 (N_2899,N_544,N_725);
nand U2900 (N_2900,N_153,N_1357);
nor U2901 (N_2901,N_168,N_2097);
nand U2902 (N_2902,N_29,N_757);
xnor U2903 (N_2903,N_2361,N_967);
nand U2904 (N_2904,N_1490,N_481);
or U2905 (N_2905,N_1968,N_144);
nor U2906 (N_2906,N_1280,N_1408);
nor U2907 (N_2907,N_2103,N_1503);
nor U2908 (N_2908,N_167,N_1075);
nand U2909 (N_2909,N_1957,N_1655);
xor U2910 (N_2910,N_856,N_1117);
nor U2911 (N_2911,N_2317,N_137);
nand U2912 (N_2912,N_1125,N_597);
xnor U2913 (N_2913,N_1680,N_10);
or U2914 (N_2914,N_594,N_1736);
nand U2915 (N_2915,N_2245,N_420);
and U2916 (N_2916,N_1085,N_379);
xnor U2917 (N_2917,N_186,N_1726);
nor U2918 (N_2918,N_2184,N_417);
nand U2919 (N_2919,N_2171,N_510);
and U2920 (N_2920,N_1191,N_1672);
nor U2921 (N_2921,N_813,N_1167);
xor U2922 (N_2922,N_1051,N_1663);
nand U2923 (N_2923,N_25,N_2149);
and U2924 (N_2924,N_1447,N_1782);
xnor U2925 (N_2925,N_452,N_1211);
or U2926 (N_2926,N_2357,N_1698);
nor U2927 (N_2927,N_1000,N_1778);
or U2928 (N_2928,N_1471,N_1729);
xor U2929 (N_2929,N_658,N_411);
nor U2930 (N_2930,N_1809,N_791);
nand U2931 (N_2931,N_705,N_286);
and U2932 (N_2932,N_1007,N_177);
nor U2933 (N_2933,N_1956,N_831);
nand U2934 (N_2934,N_207,N_819);
and U2935 (N_2935,N_1748,N_1119);
and U2936 (N_2936,N_853,N_1903);
xor U2937 (N_2937,N_1617,N_2376);
nor U2938 (N_2938,N_1891,N_1461);
or U2939 (N_2939,N_1021,N_1803);
nand U2940 (N_2940,N_386,N_1817);
nand U2941 (N_2941,N_2360,N_588);
nand U2942 (N_2942,N_2322,N_1944);
or U2943 (N_2943,N_1861,N_938);
nand U2944 (N_2944,N_1747,N_473);
and U2945 (N_2945,N_1510,N_1459);
and U2946 (N_2946,N_1606,N_887);
nor U2947 (N_2947,N_1171,N_1566);
xnor U2948 (N_2948,N_446,N_1370);
or U2949 (N_2949,N_2114,N_124);
and U2950 (N_2950,N_1150,N_1523);
or U2951 (N_2951,N_1500,N_1103);
nand U2952 (N_2952,N_142,N_250);
nor U2953 (N_2953,N_2159,N_2072);
nand U2954 (N_2954,N_1267,N_33);
or U2955 (N_2955,N_2417,N_2335);
or U2956 (N_2956,N_741,N_578);
nand U2957 (N_2957,N_240,N_1399);
nand U2958 (N_2958,N_151,N_1882);
and U2959 (N_2959,N_1505,N_341);
nand U2960 (N_2960,N_1658,N_1241);
nand U2961 (N_2961,N_50,N_678);
xor U2962 (N_2962,N_156,N_822);
and U2963 (N_2963,N_612,N_2095);
nand U2964 (N_2964,N_176,N_957);
nor U2965 (N_2965,N_272,N_441);
xnor U2966 (N_2966,N_2410,N_1881);
or U2967 (N_2967,N_1933,N_1999);
and U2968 (N_2968,N_149,N_811);
or U2969 (N_2969,N_1446,N_1997);
nand U2970 (N_2970,N_175,N_2076);
nand U2971 (N_2971,N_1113,N_651);
nand U2972 (N_2972,N_2048,N_1650);
xnor U2973 (N_2973,N_1952,N_1145);
or U2974 (N_2974,N_264,N_2145);
nor U2975 (N_2975,N_1840,N_706);
nand U2976 (N_2976,N_1299,N_921);
nand U2977 (N_2977,N_1804,N_2265);
or U2978 (N_2978,N_1607,N_857);
nor U2979 (N_2979,N_953,N_383);
xnor U2980 (N_2980,N_132,N_1372);
xor U2981 (N_2981,N_335,N_265);
and U2982 (N_2982,N_497,N_65);
or U2983 (N_2983,N_1226,N_1789);
nand U2984 (N_2984,N_908,N_1216);
nand U2985 (N_2985,N_1712,N_2088);
nand U2986 (N_2986,N_2054,N_1536);
nor U2987 (N_2987,N_1811,N_1325);
xor U2988 (N_2988,N_560,N_2388);
xor U2989 (N_2989,N_1365,N_2111);
nor U2990 (N_2990,N_1468,N_998);
nand U2991 (N_2991,N_1808,N_2318);
and U2992 (N_2992,N_2305,N_27);
xnor U2993 (N_2993,N_1528,N_2385);
xor U2994 (N_2994,N_2230,N_1589);
and U2995 (N_2995,N_1781,N_1111);
nor U2996 (N_2996,N_607,N_1250);
nor U2997 (N_2997,N_2136,N_178);
or U2998 (N_2998,N_1786,N_2312);
nand U2999 (N_2999,N_1331,N_42);
nor U3000 (N_3000,N_1344,N_1591);
or U3001 (N_3001,N_1229,N_182);
xnor U3002 (N_3002,N_1153,N_2167);
xor U3003 (N_3003,N_281,N_2316);
nand U3004 (N_3004,N_676,N_1082);
nor U3005 (N_3005,N_2139,N_380);
xnor U3006 (N_3006,N_1120,N_2278);
or U3007 (N_3007,N_1833,N_639);
nor U3008 (N_3008,N_37,N_2254);
or U3009 (N_3009,N_2075,N_1689);
nand U3010 (N_3010,N_1326,N_360);
nand U3011 (N_3011,N_952,N_1149);
or U3012 (N_3012,N_1974,N_2229);
nor U3013 (N_3013,N_489,N_322);
xor U3014 (N_3014,N_1711,N_259);
nor U3015 (N_3015,N_753,N_321);
nand U3016 (N_3016,N_2419,N_2394);
and U3017 (N_3017,N_62,N_563);
nand U3018 (N_3018,N_1264,N_231);
nand U3019 (N_3019,N_919,N_522);
nand U3020 (N_3020,N_1225,N_435);
and U3021 (N_3021,N_2013,N_1868);
nand U3022 (N_3022,N_1744,N_1652);
or U3023 (N_3023,N_211,N_564);
nand U3024 (N_3024,N_2266,N_467);
xor U3025 (N_3025,N_2227,N_2215);
and U3026 (N_3026,N_1960,N_1834);
xor U3027 (N_3027,N_1245,N_2173);
nor U3028 (N_3028,N_1513,N_127);
xnor U3029 (N_3029,N_39,N_412);
nand U3030 (N_3030,N_864,N_1750);
or U3031 (N_3031,N_1688,N_1141);
nor U3032 (N_3032,N_726,N_738);
or U3033 (N_3033,N_371,N_562);
or U3034 (N_3034,N_491,N_992);
and U3035 (N_3035,N_755,N_2451);
and U3036 (N_3036,N_946,N_2440);
xor U3037 (N_3037,N_2340,N_926);
or U3038 (N_3038,N_2498,N_276);
and U3039 (N_3039,N_2022,N_898);
xnor U3040 (N_3040,N_1130,N_761);
and U3041 (N_3041,N_1870,N_2211);
nor U3042 (N_3042,N_516,N_1025);
and U3043 (N_3043,N_1048,N_920);
and U3044 (N_3044,N_2040,N_1992);
or U3045 (N_3045,N_164,N_494);
or U3046 (N_3046,N_239,N_1969);
nand U3047 (N_3047,N_2192,N_1003);
nor U3048 (N_3048,N_1812,N_424);
nor U3049 (N_3049,N_1173,N_526);
and U3050 (N_3050,N_1499,N_2058);
xnor U3051 (N_3051,N_1930,N_188);
nor U3052 (N_3052,N_2107,N_111);
and U3053 (N_3053,N_1306,N_1382);
and U3054 (N_3054,N_2178,N_795);
and U3055 (N_3055,N_2128,N_1183);
or U3056 (N_3056,N_306,N_1334);
nand U3057 (N_3057,N_768,N_1142);
or U3058 (N_3058,N_469,N_1349);
nand U3059 (N_3059,N_1212,N_1945);
nand U3060 (N_3060,N_1660,N_1873);
nand U3061 (N_3061,N_328,N_2433);
xor U3062 (N_3062,N_431,N_1086);
xnor U3063 (N_3063,N_197,N_586);
nor U3064 (N_3064,N_2166,N_608);
nor U3065 (N_3065,N_1627,N_1743);
and U3066 (N_3066,N_541,N_1206);
and U3067 (N_3067,N_2267,N_947);
xor U3068 (N_3068,N_1091,N_128);
or U3069 (N_3069,N_1409,N_1635);
xnor U3070 (N_3070,N_2102,N_1430);
and U3071 (N_3071,N_267,N_499);
or U3072 (N_3072,N_949,N_1696);
and U3073 (N_3073,N_1074,N_76);
nand U3074 (N_3074,N_1837,N_2152);
nand U3075 (N_3075,N_875,N_2221);
xor U3076 (N_3076,N_1376,N_1721);
xor U3077 (N_3077,N_1320,N_2049);
nand U3078 (N_3078,N_1137,N_1348);
nor U3079 (N_3079,N_1714,N_1697);
xor U3080 (N_3080,N_569,N_1450);
nor U3081 (N_3081,N_1610,N_969);
xnor U3082 (N_3082,N_1417,N_843);
nor U3083 (N_3083,N_415,N_466);
and U3084 (N_3084,N_2231,N_418);
nand U3085 (N_3085,N_1199,N_1488);
nor U3086 (N_3086,N_86,N_804);
xor U3087 (N_3087,N_599,N_1507);
or U3088 (N_3088,N_1332,N_2395);
or U3089 (N_3089,N_585,N_406);
xnor U3090 (N_3090,N_2275,N_2242);
nor U3091 (N_3091,N_438,N_1249);
nor U3092 (N_3092,N_1102,N_1168);
xor U3093 (N_3093,N_1599,N_1140);
xor U3094 (N_3094,N_1390,N_1484);
nand U3095 (N_3095,N_889,N_1979);
and U3096 (N_3096,N_790,N_1520);
and U3097 (N_3097,N_9,N_1594);
nor U3098 (N_3098,N_1541,N_2146);
nor U3099 (N_3099,N_1538,N_1339);
and U3100 (N_3100,N_851,N_1002);
and U3101 (N_3101,N_1254,N_214);
xor U3102 (N_3102,N_318,N_1874);
xnor U3103 (N_3103,N_879,N_910);
or U3104 (N_3104,N_764,N_554);
xnor U3105 (N_3105,N_603,N_208);
and U3106 (N_3106,N_553,N_2195);
and U3107 (N_3107,N_828,N_1766);
or U3108 (N_3108,N_1350,N_2426);
nor U3109 (N_3109,N_543,N_1552);
nand U3110 (N_3110,N_1287,N_2493);
nor U3111 (N_3111,N_1575,N_723);
nand U3112 (N_3112,N_2436,N_695);
xnor U3113 (N_3113,N_858,N_194);
nor U3114 (N_3114,N_1816,N_308);
nor U3115 (N_3115,N_1806,N_2);
nor U3116 (N_3116,N_483,N_2476);
nand U3117 (N_3117,N_986,N_354);
or U3118 (N_3118,N_859,N_703);
or U3119 (N_3119,N_2306,N_771);
nor U3120 (N_3120,N_2407,N_408);
or U3121 (N_3121,N_2113,N_769);
xor U3122 (N_3122,N_226,N_881);
xor U3123 (N_3123,N_2430,N_1480);
xor U3124 (N_3124,N_2479,N_71);
nand U3125 (N_3125,N_23,N_1491);
or U3126 (N_3126,N_2101,N_458);
nor U3127 (N_3127,N_1208,N_1539);
xnor U3128 (N_3128,N_1359,N_2090);
nand U3129 (N_3129,N_1964,N_2403);
nor U3130 (N_3130,N_1549,N_2464);
nor U3131 (N_3131,N_344,N_429);
or U3132 (N_3132,N_253,N_1702);
nand U3133 (N_3133,N_1410,N_1184);
nor U3134 (N_3134,N_1879,N_107);
and U3135 (N_3135,N_234,N_432);
or U3136 (N_3136,N_834,N_1752);
xnor U3137 (N_3137,N_316,N_495);
and U3138 (N_3138,N_989,N_66);
nor U3139 (N_3139,N_2294,N_1121);
nand U3140 (N_3140,N_849,N_2108);
or U3141 (N_3141,N_927,N_847);
xnor U3142 (N_3142,N_1629,N_1831);
or U3143 (N_3143,N_1414,N_241);
and U3144 (N_3144,N_1919,N_1251);
xnor U3145 (N_3145,N_618,N_2399);
xnor U3146 (N_3146,N_18,N_1345);
nor U3147 (N_3147,N_2041,N_1247);
and U3148 (N_3148,N_1553,N_135);
nor U3149 (N_3149,N_679,N_1783);
nor U3150 (N_3150,N_1685,N_2078);
or U3151 (N_3151,N_796,N_1900);
nand U3152 (N_3152,N_2348,N_1458);
nor U3153 (N_3153,N_1695,N_2005);
or U3154 (N_3154,N_413,N_2125);
or U3155 (N_3155,N_1050,N_659);
nor U3156 (N_3156,N_72,N_2452);
nor U3157 (N_3157,N_2422,N_1083);
or U3158 (N_3158,N_1217,N_1190);
and U3159 (N_3159,N_238,N_1260);
or U3160 (N_3160,N_1545,N_280);
nor U3161 (N_3161,N_305,N_2374);
nor U3162 (N_3162,N_2490,N_2461);
or U3163 (N_3163,N_1386,N_1139);
nand U3164 (N_3164,N_1389,N_1797);
nand U3165 (N_3165,N_268,N_81);
xor U3166 (N_3166,N_1673,N_1978);
nor U3167 (N_3167,N_507,N_784);
nor U3168 (N_3168,N_1628,N_2188);
or U3169 (N_3169,N_943,N_1982);
nand U3170 (N_3170,N_402,N_165);
or U3171 (N_3171,N_1170,N_1397);
and U3172 (N_3172,N_1286,N_687);
or U3173 (N_3173,N_2389,N_1511);
nor U3174 (N_3174,N_131,N_2342);
nand U3175 (N_3175,N_1232,N_2175);
xnor U3176 (N_3176,N_1038,N_2332);
xor U3177 (N_3177,N_1769,N_1017);
and U3178 (N_3178,N_2117,N_968);
nor U3179 (N_3179,N_463,N_1115);
and U3180 (N_3180,N_329,N_1990);
and U3181 (N_3181,N_1625,N_49);
xor U3182 (N_3182,N_2119,N_855);
or U3183 (N_3183,N_179,N_1892);
or U3184 (N_3184,N_2104,N_2019);
nor U3185 (N_3185,N_422,N_487);
nor U3186 (N_3186,N_14,N_450);
or U3187 (N_3187,N_669,N_451);
or U3188 (N_3188,N_2481,N_1574);
xor U3189 (N_3189,N_1517,N_1027);
nor U3190 (N_3190,N_728,N_410);
nor U3191 (N_3191,N_2164,N_41);
xor U3192 (N_3192,N_797,N_584);
and U3193 (N_3193,N_465,N_464);
and U3194 (N_3194,N_1709,N_1322);
or U3195 (N_3195,N_1033,N_1394);
and U3196 (N_3196,N_112,N_566);
nor U3197 (N_3197,N_1215,N_2398);
or U3198 (N_3198,N_116,N_2100);
nand U3199 (N_3199,N_130,N_1754);
nand U3200 (N_3200,N_535,N_754);
xnor U3201 (N_3201,N_1300,N_2478);
or U3202 (N_3202,N_232,N_1569);
and U3203 (N_3203,N_749,N_1515);
or U3204 (N_3204,N_970,N_758);
nor U3205 (N_3205,N_2368,N_615);
or U3206 (N_3206,N_2015,N_906);
xnor U3207 (N_3207,N_209,N_925);
nand U3208 (N_3208,N_2059,N_1131);
xor U3209 (N_3209,N_646,N_2073);
xnor U3210 (N_3210,N_1996,N_1779);
and U3211 (N_3211,N_610,N_183);
xor U3212 (N_3212,N_1421,N_376);
nand U3213 (N_3213,N_2141,N_1404);
and U3214 (N_3214,N_95,N_1583);
nor U3215 (N_3215,N_2411,N_924);
and U3216 (N_3216,N_93,N_2449);
or U3217 (N_3217,N_686,N_2083);
and U3218 (N_3218,N_2190,N_1601);
or U3219 (N_3219,N_1871,N_1279);
nor U3220 (N_3220,N_1746,N_800);
nor U3221 (N_3221,N_2429,N_278);
xor U3222 (N_3222,N_2255,N_1407);
nand U3223 (N_3223,N_1311,N_2379);
or U3224 (N_3224,N_565,N_684);
nor U3225 (N_3225,N_1460,N_1378);
and U3226 (N_3226,N_1890,N_1238);
nand U3227 (N_3227,N_2247,N_527);
nand U3228 (N_3228,N_52,N_792);
xnor U3229 (N_3229,N_980,N_106);
and U3230 (N_3230,N_1388,N_1313);
nand U3231 (N_3231,N_1699,N_1518);
xor U3232 (N_3232,N_1455,N_1147);
nor U3233 (N_3233,N_2296,N_850);
nor U3234 (N_3234,N_752,N_2047);
and U3235 (N_3235,N_1554,N_891);
nor U3236 (N_3236,N_892,N_160);
and U3237 (N_3237,N_1343,N_1169);
xor U3238 (N_3238,N_311,N_1159);
and U3239 (N_3239,N_199,N_737);
xor U3240 (N_3240,N_2304,N_1093);
and U3241 (N_3241,N_664,N_1773);
and U3242 (N_3242,N_1570,N_99);
nand U3243 (N_3243,N_2185,N_279);
nand U3244 (N_3244,N_2483,N_2094);
xnor U3245 (N_3245,N_638,N_873);
or U3246 (N_3246,N_1847,N_1916);
nor U3247 (N_3247,N_1525,N_140);
nor U3248 (N_3248,N_1175,N_1590);
and U3249 (N_3249,N_2349,N_1864);
nor U3250 (N_3250,N_1637,N_2080);
nor U3251 (N_3251,N_262,N_816);
or U3252 (N_3252,N_1691,N_1800);
and U3253 (N_3253,N_439,N_1951);
or U3254 (N_3254,N_1268,N_2445);
nand U3255 (N_3255,N_1762,N_1266);
and U3256 (N_3256,N_1571,N_448);
nand U3257 (N_3257,N_486,N_1694);
nor U3258 (N_3258,N_1971,N_244);
nand U3259 (N_3259,N_2382,N_170);
nand U3260 (N_3260,N_369,N_427);
xnor U3261 (N_3261,N_453,N_966);
nor U3262 (N_3262,N_2408,N_1501);
or U3263 (N_3263,N_24,N_1498);
nand U3264 (N_3264,N_1118,N_228);
or U3265 (N_3265,N_775,N_2303);
nand U3266 (N_3266,N_1679,N_699);
xor U3267 (N_3267,N_399,N_338);
or U3268 (N_3268,N_2358,N_1662);
or U3269 (N_3269,N_1495,N_592);
nand U3270 (N_3270,N_2383,N_1862);
or U3271 (N_3271,N_1761,N_2310);
nand U3272 (N_3272,N_1745,N_1434);
xor U3273 (N_3273,N_1479,N_1055);
or U3274 (N_3274,N_878,N_1188);
nand U3275 (N_3275,N_361,N_114);
xor U3276 (N_3276,N_2220,N_1818);
or U3277 (N_3277,N_163,N_1432);
nor U3278 (N_3278,N_545,N_2057);
or U3279 (N_3279,N_900,N_654);
xor U3280 (N_3280,N_1010,N_1889);
xor U3281 (N_3281,N_2240,N_1865);
nand U3282 (N_3282,N_1195,N_691);
or U3283 (N_3283,N_1731,N_1561);
nand U3284 (N_3284,N_2137,N_326);
nand U3285 (N_3285,N_1242,N_1442);
and U3286 (N_3286,N_2268,N_425);
nand U3287 (N_3287,N_225,N_1123);
and U3288 (N_3288,N_841,N_606);
nand U3289 (N_3289,N_1258,N_2148);
or U3290 (N_3290,N_2401,N_394);
nor U3291 (N_3291,N_2180,N_353);
xnor U3292 (N_3292,N_1646,N_756);
or U3293 (N_3293,N_2346,N_63);
nand U3294 (N_3294,N_1088,N_340);
and U3295 (N_3295,N_2027,N_1516);
nand U3296 (N_3296,N_2391,N_1654);
nor U3297 (N_3297,N_1419,N_1163);
or U3298 (N_3298,N_1687,N_697);
nor U3299 (N_3299,N_2163,N_2338);
nor U3300 (N_3300,N_1030,N_242);
or U3301 (N_3301,N_217,N_1310);
nor U3302 (N_3302,N_1563,N_688);
xnor U3303 (N_3303,N_1064,N_2000);
or U3304 (N_3304,N_1970,N_1730);
and U3305 (N_3305,N_1308,N_403);
nor U3306 (N_3306,N_1630,N_474);
xnor U3307 (N_3307,N_2071,N_501);
nand U3308 (N_3308,N_2116,N_1883);
xor U3309 (N_3309,N_2354,N_1706);
nor U3310 (N_3310,N_304,N_2336);
nand U3311 (N_3311,N_476,N_75);
or U3312 (N_3312,N_1597,N_662);
nor U3313 (N_3313,N_1636,N_101);
or U3314 (N_3314,N_1504,N_454);
and U3315 (N_3315,N_1634,N_1333);
nand U3316 (N_3316,N_166,N_1657);
and U3317 (N_3317,N_2480,N_1393);
or U3318 (N_3318,N_1546,N_558);
xor U3319 (N_3319,N_2284,N_1527);
xnor U3320 (N_3320,N_1068,N_504);
nand U3321 (N_3321,N_2472,N_750);
or U3322 (N_3322,N_824,N_1832);
xnor U3323 (N_3323,N_1760,N_449);
nor U3324 (N_3324,N_436,N_51);
and U3325 (N_3325,N_2168,N_1057);
nor U3326 (N_3326,N_914,N_1252);
nor U3327 (N_3327,N_576,N_827);
and U3328 (N_3328,N_310,N_1774);
nand U3329 (N_3329,N_587,N_141);
or U3330 (N_3330,N_1441,N_524);
xnor U3331 (N_3331,N_1342,N_34);
xnor U3332 (N_3332,N_670,N_718);
nor U3333 (N_3333,N_2437,N_1108);
and U3334 (N_3334,N_73,N_2202);
or U3335 (N_3335,N_1244,N_291);
or U3336 (N_3336,N_1640,N_89);
nor U3337 (N_3337,N_1444,N_1281);
nor U3338 (N_3338,N_233,N_994);
and U3339 (N_3339,N_978,N_1734);
nand U3340 (N_3340,N_1069,N_1815);
and U3341 (N_3341,N_1039,N_1040);
nor U3342 (N_3342,N_580,N_1124);
or U3343 (N_3343,N_1470,N_1906);
nor U3344 (N_3344,N_1790,N_1995);
and U3345 (N_3345,N_1519,N_896);
nor U3346 (N_3346,N_2143,N_2077);
nor U3347 (N_3347,N_2179,N_64);
and U3348 (N_3348,N_1844,N_1642);
nand U3349 (N_3349,N_720,N_766);
xnor U3350 (N_3350,N_53,N_867);
or U3351 (N_3351,N_96,N_711);
nor U3352 (N_3352,N_996,N_975);
nand U3353 (N_3353,N_886,N_1476);
and U3354 (N_3354,N_19,N_2288);
nand U3355 (N_3355,N_2413,N_776);
xnor U3356 (N_3356,N_2292,N_1615);
xor U3357 (N_3357,N_1243,N_1638);
xor U3358 (N_3358,N_2093,N_2038);
nor U3359 (N_3359,N_745,N_1248);
and U3360 (N_3360,N_1923,N_283);
or U3361 (N_3361,N_620,N_400);
nor U3362 (N_3362,N_893,N_1799);
and U3363 (N_3363,N_1738,N_255);
or U3364 (N_3364,N_1624,N_1087);
nand U3365 (N_3365,N_2311,N_1439);
and U3366 (N_3366,N_950,N_689);
nand U3367 (N_3367,N_2280,N_320);
xor U3368 (N_3368,N_1383,N_973);
or U3369 (N_3369,N_2380,N_319);
and U3370 (N_3370,N_742,N_1814);
nand U3371 (N_3371,N_683,N_2253);
or U3372 (N_3372,N_1567,N_2441);
or U3373 (N_3373,N_1469,N_252);
nor U3374 (N_3374,N_2415,N_190);
nor U3375 (N_3375,N_1788,N_1477);
xor U3376 (N_3376,N_1304,N_1412);
xor U3377 (N_3377,N_868,N_355);
nor U3378 (N_3378,N_223,N_1425);
nor U3379 (N_3379,N_203,N_1669);
xor U3380 (N_3380,N_1156,N_1619);
xor U3381 (N_3381,N_2442,N_298);
or U3382 (N_3382,N_1829,N_2025);
nand U3383 (N_3383,N_364,N_1859);
or U3384 (N_3384,N_865,N_2042);
nand U3385 (N_3385,N_918,N_717);
nand U3386 (N_3386,N_2039,N_539);
nor U3387 (N_3387,N_1794,N_660);
xnor U3388 (N_3388,N_812,N_2257);
nand U3389 (N_3389,N_1558,N_2434);
nor U3390 (N_3390,N_1454,N_1966);
or U3391 (N_3391,N_1535,N_392);
and U3392 (N_3392,N_2264,N_602);
or U3393 (N_3393,N_515,N_1296);
nand U3394 (N_3394,N_2384,N_762);
nor U3395 (N_3395,N_1719,N_2151);
nand U3396 (N_3396,N_2438,N_570);
xnor U3397 (N_3397,N_1674,N_842);
and U3398 (N_3398,N_1989,N_1023);
and U3399 (N_3399,N_2319,N_271);
and U3400 (N_3400,N_1572,N_146);
xor U3401 (N_3401,N_1949,N_2186);
nor U3402 (N_3402,N_147,N_561);
xor U3403 (N_3403,N_1723,N_1116);
and U3404 (N_3404,N_2414,N_1621);
nand U3405 (N_3405,N_1912,N_1155);
or U3406 (N_3406,N_740,N_1496);
nor U3407 (N_3407,N_1369,N_1481);
nand U3408 (N_3408,N_1605,N_2281);
xor U3409 (N_3409,N_1096,N_2082);
xor U3410 (N_3410,N_327,N_835);
nor U3411 (N_3411,N_814,N_2276);
or U3412 (N_3412,N_1733,N_722);
nand U3413 (N_3413,N_136,N_315);
nand U3414 (N_3414,N_1486,N_440);
and U3415 (N_3415,N_1328,N_378);
xor U3416 (N_3416,N_2087,N_988);
nand U3417 (N_3417,N_1233,N_649);
xor U3418 (N_3418,N_1197,N_1060);
and U3419 (N_3419,N_1443,N_1200);
nand U3420 (N_3420,N_625,N_447);
nand U3421 (N_3421,N_2477,N_901);
xor U3422 (N_3422,N_58,N_385);
nand U3423 (N_3423,N_395,N_2324);
or U3424 (N_3424,N_1845,N_2045);
xnor U3425 (N_3425,N_1392,N_1767);
nand U3426 (N_3426,N_690,N_330);
xor U3427 (N_3427,N_1494,N_70);
and U3428 (N_3428,N_1079,N_374);
and U3429 (N_3429,N_245,N_888);
nand U3430 (N_3430,N_1728,N_1204);
xnor U3431 (N_3431,N_1351,N_915);
and U3432 (N_3432,N_1230,N_1492);
and U3433 (N_3433,N_105,N_1253);
and U3434 (N_3434,N_2443,N_2400);
or U3435 (N_3435,N_1396,N_808);
nand U3436 (N_3436,N_2269,N_437);
or U3437 (N_3437,N_911,N_677);
nand U3438 (N_3438,N_1047,N_1988);
nor U3439 (N_3439,N_1319,N_2052);
nor U3440 (N_3440,N_212,N_2199);
nor U3441 (N_3441,N_2435,N_246);
nor U3442 (N_3442,N_951,N_1445);
and U3443 (N_3443,N_1256,N_845);
or U3444 (N_3444,N_1448,N_496);
nor U3445 (N_3445,N_1693,N_1366);
nor U3446 (N_3446,N_1676,N_1042);
and U3447 (N_3447,N_2129,N_2263);
nor U3448 (N_3448,N_1401,N_2475);
and U3449 (N_3449,N_337,N_274);
nor U3450 (N_3450,N_1542,N_614);
nand U3451 (N_3451,N_1768,N_2372);
xor U3452 (N_3452,N_2467,N_2021);
and U3453 (N_3453,N_627,N_348);
nand U3454 (N_3454,N_1826,N_1305);
xnor U3455 (N_3455,N_1976,N_2084);
nand U3456 (N_3456,N_1524,N_1792);
nand U3457 (N_3457,N_300,N_43);
nand U3458 (N_3458,N_2488,N_767);
nand U3459 (N_3459,N_735,N_444);
or U3460 (N_3460,N_591,N_961);
and U3461 (N_3461,N_1178,N_1824);
and U3462 (N_3462,N_423,N_1986);
and U3463 (N_3463,N_1722,N_120);
or U3464 (N_3464,N_2409,N_1564);
nand U3465 (N_3465,N_1013,N_1176);
nor U3466 (N_3466,N_2065,N_1645);
nand U3467 (N_3467,N_1015,N_573);
nand U3468 (N_3468,N_2037,N_97);
and U3469 (N_3469,N_1913,N_1877);
or U3470 (N_3470,N_1099,N_1041);
and U3471 (N_3471,N_1963,N_1052);
nand U3472 (N_3472,N_44,N_1274);
nand U3473 (N_3473,N_707,N_443);
xor U3474 (N_3474,N_668,N_1994);
and U3475 (N_3475,N_2274,N_1029);
and U3476 (N_3476,N_2421,N_1869);
or U3477 (N_3477,N_1681,N_884);
nand U3478 (N_3478,N_1323,N_1295);
nor U3479 (N_3479,N_1853,N_2297);
and U3480 (N_3480,N_1166,N_88);
or U3481 (N_3481,N_181,N_363);
and U3482 (N_3482,N_1596,N_1489);
or U3483 (N_3483,N_557,N_1006);
xor U3484 (N_3484,N_825,N_2007);
and U3485 (N_3485,N_138,N_2237);
nor U3486 (N_3486,N_546,N_1403);
and U3487 (N_3487,N_2454,N_296);
or U3488 (N_3488,N_1927,N_373);
and U3489 (N_3489,N_292,N_799);
and U3490 (N_3490,N_1172,N_1035);
xnor U3491 (N_3491,N_2046,N_551);
xor U3492 (N_3492,N_517,N_1291);
or U3493 (N_3493,N_1227,N_1823);
nor U3494 (N_3494,N_2378,N_1493);
and U3495 (N_3495,N_2248,N_84);
and U3496 (N_3496,N_1462,N_1835);
and U3497 (N_3497,N_2373,N_1531);
and U3498 (N_3498,N_2121,N_2086);
or U3499 (N_3499,N_729,N_91);
nand U3500 (N_3500,N_1623,N_2068);
nor U3501 (N_3501,N_1364,N_222);
xor U3502 (N_3502,N_2138,N_457);
or U3503 (N_3503,N_1497,N_1066);
or U3504 (N_3504,N_1203,N_779);
nor U3505 (N_3505,N_932,N_1457);
and U3506 (N_3506,N_694,N_1073);
and U3507 (N_3507,N_158,N_1633);
xnor U3508 (N_3508,N_840,N_419);
nand U3509 (N_3509,N_929,N_529);
or U3510 (N_3510,N_1234,N_1855);
or U3511 (N_3511,N_6,N_1415);
nor U3512 (N_3512,N_1741,N_2140);
or U3513 (N_3513,N_1138,N_798);
xor U3514 (N_3514,N_196,N_1427);
xor U3515 (N_3515,N_40,N_1067);
nand U3516 (N_3516,N_1533,N_1024);
nand U3517 (N_3517,N_1850,N_1878);
nand U3518 (N_3518,N_1420,N_631);
or U3519 (N_3519,N_1095,N_2157);
nor U3520 (N_3520,N_1373,N_2142);
and U3521 (N_3521,N_734,N_604);
or U3522 (N_3522,N_657,N_324);
or U3523 (N_3523,N_976,N_1418);
nor U3524 (N_3524,N_820,N_1568);
nand U3525 (N_3525,N_1543,N_1725);
xnor U3526 (N_3526,N_2225,N_2386);
xnor U3527 (N_3527,N_536,N_2313);
or U3528 (N_3528,N_2420,N_1704);
or U3529 (N_3529,N_1918,N_2427);
or U3530 (N_3530,N_1600,N_1261);
nand U3531 (N_3531,N_2446,N_12);
nand U3532 (N_3532,N_1043,N_528);
and U3533 (N_3533,N_1,N_126);
nor U3534 (N_3534,N_549,N_1294);
nand U3535 (N_3535,N_456,N_2099);
and U3536 (N_3536,N_54,N_1288);
nor U3537 (N_3537,N_626,N_1127);
xnor U3538 (N_3538,N_1014,N_1942);
nor U3539 (N_3539,N_205,N_257);
or U3540 (N_3540,N_2457,N_2272);
or U3541 (N_3541,N_173,N_2390);
nand U3542 (N_3542,N_2106,N_213);
and U3543 (N_3543,N_1909,N_1278);
xor U3544 (N_3544,N_375,N_1675);
xnor U3545 (N_3545,N_2333,N_1720);
nor U3546 (N_3546,N_426,N_1893);
or U3547 (N_3547,N_770,N_630);
xnor U3548 (N_3548,N_661,N_518);
nor U3549 (N_3549,N_2232,N_189);
xor U3550 (N_3550,N_1897,N_273);
nand U3551 (N_3551,N_806,N_590);
or U3552 (N_3552,N_1926,N_159);
nand U3553 (N_3553,N_1431,N_459);
xnor U3554 (N_3554,N_1375,N_1269);
nand U3555 (N_3555,N_1213,N_1433);
nor U3556 (N_3556,N_948,N_650);
nand U3557 (N_3557,N_1207,N_1174);
xor U3558 (N_3558,N_579,N_1056);
and U3559 (N_3559,N_350,N_1908);
or U3560 (N_3560,N_2371,N_781);
and U3561 (N_3561,N_22,N_1841);
or U3562 (N_3562,N_1474,N_1950);
nand U3563 (N_3563,N_942,N_2487);
and U3564 (N_3564,N_595,N_462);
or U3565 (N_3565,N_1772,N_1522);
or U3566 (N_3566,N_1193,N_2063);
nor U3567 (N_3567,N_2327,N_2282);
xnor U3568 (N_3568,N_1895,N_299);
xnor U3569 (N_3569,N_682,N_2181);
and U3570 (N_3570,N_674,N_1005);
nor U3571 (N_3571,N_118,N_2123);
nor U3572 (N_3572,N_13,N_739);
or U3573 (N_3573,N_1224,N_1036);
or U3574 (N_3574,N_1732,N_1587);
and U3575 (N_3575,N_1622,N_2331);
and U3576 (N_3576,N_1911,N_1958);
xor U3577 (N_3577,N_653,N_351);
and U3578 (N_3578,N_270,N_748);
xor U3579 (N_3579,N_336,N_1424);
nor U3580 (N_3580,N_1759,N_1710);
or U3581 (N_3581,N_2020,N_2122);
nand U3582 (N_3582,N_1098,N_1368);
and U3583 (N_3583,N_883,N_2133);
xnor U3584 (N_3584,N_2470,N_152);
nor U3585 (N_3585,N_916,N_2008);
nand U3586 (N_3586,N_1133,N_945);
nand U3587 (N_3587,N_1478,N_2406);
and U3588 (N_3588,N_1975,N_1273);
or U3589 (N_3589,N_1189,N_960);
nor U3590 (N_3590,N_2309,N_1932);
nor U3591 (N_3591,N_861,N_1423);
and U3592 (N_3592,N_1934,N_2471);
xnor U3593 (N_3593,N_1880,N_1998);
xnor U3594 (N_3594,N_616,N_2397);
xor U3595 (N_3595,N_1984,N_1080);
or U3596 (N_3596,N_826,N_254);
nor U3597 (N_3597,N_256,N_2328);
nor U3598 (N_3598,N_685,N_191);
nor U3599 (N_3599,N_1757,N_648);
nand U3600 (N_3600,N_381,N_2250);
and U3601 (N_3601,N_1034,N_2325);
nor U3602 (N_3602,N_917,N_2187);
or U3603 (N_3603,N_2183,N_372);
and U3604 (N_3604,N_2456,N_963);
nand U3605 (N_3605,N_537,N_852);
nor U3606 (N_3606,N_583,N_2062);
or U3607 (N_3607,N_2298,N_1451);
nand U3608 (N_3608,N_1550,N_572);
and U3609 (N_3609,N_1713,N_1018);
and U3610 (N_3610,N_2053,N_1318);
or U3611 (N_3611,N_698,N_249);
and U3612 (N_3612,N_1993,N_1179);
xor U3613 (N_3613,N_2109,N_777);
xnor U3614 (N_3614,N_1263,N_172);
nand U3615 (N_3615,N_1221,N_1791);
or U3616 (N_3616,N_1664,N_1796);
or U3617 (N_3617,N_656,N_1678);
xnor U3618 (N_3618,N_2154,N_2287);
nor U3619 (N_3619,N_876,N_704);
xor U3620 (N_3620,N_393,N_803);
nand U3621 (N_3621,N_1182,N_409);
or U3622 (N_3622,N_2364,N_1914);
and U3623 (N_3623,N_1205,N_2473);
nor U3624 (N_3624,N_1770,N_1112);
nor U3625 (N_3625,N_1613,N_407);
and U3626 (N_3626,N_2043,N_1022);
or U3627 (N_3627,N_1836,N_506);
and U3628 (N_3628,N_1391,N_2251);
xor U3629 (N_3629,N_294,N_2460);
xnor U3630 (N_3630,N_1813,N_514);
and U3631 (N_3631,N_1708,N_2001);
xnor U3632 (N_3632,N_1595,N_1297);
or U3633 (N_3633,N_1031,N_2066);
nand U3634 (N_3634,N_2252,N_505);
and U3635 (N_3635,N_972,N_1466);
nand U3636 (N_3636,N_1857,N_772);
xor U3637 (N_3637,N_442,N_68);
nor U3638 (N_3638,N_1475,N_1529);
and U3639 (N_3639,N_333,N_956);
and U3640 (N_3640,N_974,N_589);
nand U3641 (N_3641,N_1196,N_2034);
and U3642 (N_3642,N_1282,N_701);
and U3643 (N_3643,N_362,N_1016);
nor U3644 (N_3644,N_991,N_1540);
or U3645 (N_3645,N_2323,N_692);
xor U3646 (N_3646,N_1838,N_2012);
and U3647 (N_3647,N_1449,N_2362);
xor U3648 (N_3648,N_471,N_2028);
nand U3649 (N_3649,N_384,N_357);
or U3650 (N_3650,N_1228,N_1346);
xnor U3651 (N_3651,N_712,N_2315);
or U3652 (N_3652,N_1255,N_1316);
or U3653 (N_3653,N_632,N_1285);
nor U3654 (N_3654,N_1084,N_2396);
or U3655 (N_3655,N_171,N_1852);
or U3656 (N_3656,N_48,N_1235);
nor U3657 (N_3657,N_1011,N_2307);
nor U3658 (N_3658,N_2344,N_2416);
or U3659 (N_3659,N_218,N_1985);
xnor U3660 (N_3660,N_1398,N_1604);
or U3661 (N_3661,N_210,N_1352);
or U3662 (N_3662,N_696,N_1161);
nor U3663 (N_3663,N_2234,N_2439);
nand U3664 (N_3664,N_2070,N_571);
nand U3665 (N_3665,N_1521,N_2273);
nand U3666 (N_3666,N_2064,N_644);
nand U3667 (N_3667,N_702,N_2147);
nor U3668 (N_3668,N_309,N_1753);
nand U3669 (N_3669,N_1270,N_1214);
nand U3670 (N_3670,N_2032,N_1656);
nor U3671 (N_3671,N_1186,N_103);
xnor U3672 (N_3672,N_985,N_821);
xor U3673 (N_3673,N_258,N_1128);
nor U3674 (N_3674,N_2496,N_593);
xnor U3675 (N_3675,N_493,N_525);
xor U3676 (N_3676,N_1020,N_1896);
nor U3677 (N_3677,N_1437,N_2201);
and U3678 (N_3678,N_1560,N_1160);
nor U3679 (N_3679,N_2003,N_787);
and U3680 (N_3680,N_1898,N_0);
or U3681 (N_3681,N_1290,N_870);
nand U3682 (N_3682,N_2450,N_955);
and U3683 (N_3683,N_1298,N_2492);
nand U3684 (N_3684,N_844,N_45);
nand U3685 (N_3685,N_2172,N_2200);
nor U3686 (N_3686,N_647,N_1109);
or U3687 (N_3687,N_1977,N_2194);
or U3688 (N_3688,N_184,N_2343);
xor U3689 (N_3689,N_2271,N_635);
and U3690 (N_3690,N_731,N_416);
nand U3691 (N_3691,N_937,N_1565);
nor U3692 (N_3692,N_1106,N_356);
nor U3693 (N_3693,N_2369,N_1004);
nor U3694 (N_3694,N_1557,N_1135);
nor U3695 (N_3695,N_1293,N_1502);
or U3696 (N_3696,N_2198,N_1380);
or U3697 (N_3697,N_1839,N_109);
or U3698 (N_3698,N_1948,N_2055);
nor U3699 (N_3699,N_982,N_1846);
xor U3700 (N_3700,N_2459,N_1742);
nand U3701 (N_3701,N_1094,N_359);
nor U3702 (N_3702,N_984,N_1972);
nor U3703 (N_3703,N_1327,N_1463);
or U3704 (N_3704,N_1354,N_1860);
nand U3705 (N_3705,N_1915,N_1584);
nand U3706 (N_3706,N_1436,N_482);
xnor U3707 (N_3707,N_1289,N_235);
nor U3708 (N_3708,N_1614,N_2465);
and U3709 (N_3709,N_485,N_1526);
nand U3710 (N_3710,N_922,N_2367);
or U3711 (N_3711,N_1453,N_1472);
xnor U3712 (N_3712,N_312,N_1395);
and U3713 (N_3713,N_1647,N_1315);
nand U3714 (N_3714,N_1065,N_2418);
or U3715 (N_3715,N_455,N_1842);
nor U3716 (N_3716,N_990,N_802);
or U3717 (N_3717,N_743,N_1340);
nand U3718 (N_3718,N_1576,N_1940);
or U3719 (N_3719,N_2256,N_1894);
nand U3720 (N_3720,N_1097,N_2285);
nand U3721 (N_3721,N_747,N_2018);
xnor U3722 (N_3722,N_540,N_1585);
and U3723 (N_3723,N_2352,N_815);
xnor U3724 (N_3724,N_129,N_1008);
nor U3725 (N_3725,N_1009,N_1530);
nor U3726 (N_3726,N_860,N_2289);
xor U3727 (N_3727,N_1670,N_488);
nor U3728 (N_3728,N_1198,N_885);
nand U3729 (N_3729,N_215,N_162);
or U3730 (N_3730,N_2081,N_1107);
or U3731 (N_3731,N_1707,N_1577);
and U3732 (N_3732,N_596,N_512);
nand U3733 (N_3733,N_532,N_317);
or U3734 (N_3734,N_2468,N_836);
nor U3735 (N_3735,N_389,N_520);
or U3736 (N_3736,N_1973,N_1703);
xnor U3737 (N_3737,N_17,N_575);
or U3738 (N_3738,N_2205,N_1371);
nand U3739 (N_3739,N_2334,N_401);
or U3740 (N_3740,N_2074,N_2024);
or U3741 (N_3741,N_923,N_2259);
xor U3742 (N_3742,N_905,N_1686);
xor U3743 (N_3743,N_155,N_928);
nand U3744 (N_3744,N_641,N_55);
nor U3745 (N_3745,N_1512,N_2031);
or U3746 (N_3746,N_2458,N_736);
and U3747 (N_3747,N_2428,N_538);
nand U3748 (N_3748,N_934,N_1764);
or U3749 (N_3749,N_98,N_343);
nor U3750 (N_3750,N_1256,N_1133);
nor U3751 (N_3751,N_729,N_2206);
or U3752 (N_3752,N_967,N_974);
xor U3753 (N_3753,N_1285,N_696);
xnor U3754 (N_3754,N_2023,N_540);
or U3755 (N_3755,N_1456,N_2035);
nand U3756 (N_3756,N_114,N_710);
nand U3757 (N_3757,N_177,N_596);
xnor U3758 (N_3758,N_1339,N_2483);
nor U3759 (N_3759,N_816,N_391);
nor U3760 (N_3760,N_2481,N_517);
and U3761 (N_3761,N_2414,N_818);
nand U3762 (N_3762,N_400,N_1301);
nand U3763 (N_3763,N_2152,N_1442);
and U3764 (N_3764,N_2060,N_2034);
nor U3765 (N_3765,N_982,N_1315);
nor U3766 (N_3766,N_1658,N_1704);
and U3767 (N_3767,N_541,N_322);
nor U3768 (N_3768,N_1528,N_822);
xnor U3769 (N_3769,N_707,N_463);
or U3770 (N_3770,N_784,N_1123);
xor U3771 (N_3771,N_183,N_865);
or U3772 (N_3772,N_183,N_1668);
nand U3773 (N_3773,N_580,N_1349);
nor U3774 (N_3774,N_420,N_2188);
or U3775 (N_3775,N_287,N_465);
or U3776 (N_3776,N_1516,N_1292);
nand U3777 (N_3777,N_1387,N_968);
or U3778 (N_3778,N_2101,N_413);
xnor U3779 (N_3779,N_533,N_1998);
nor U3780 (N_3780,N_2469,N_63);
xnor U3781 (N_3781,N_127,N_1122);
nor U3782 (N_3782,N_551,N_95);
or U3783 (N_3783,N_1556,N_58);
nor U3784 (N_3784,N_713,N_1602);
xor U3785 (N_3785,N_1167,N_1322);
or U3786 (N_3786,N_2282,N_772);
or U3787 (N_3787,N_225,N_1490);
or U3788 (N_3788,N_906,N_1646);
nand U3789 (N_3789,N_1690,N_1668);
nand U3790 (N_3790,N_1070,N_2245);
and U3791 (N_3791,N_2045,N_1725);
nand U3792 (N_3792,N_1619,N_1393);
xor U3793 (N_3793,N_1437,N_1155);
xor U3794 (N_3794,N_2134,N_1976);
and U3795 (N_3795,N_2391,N_1723);
and U3796 (N_3796,N_704,N_1648);
or U3797 (N_3797,N_1418,N_1128);
nor U3798 (N_3798,N_1476,N_49);
nor U3799 (N_3799,N_1394,N_1508);
xnor U3800 (N_3800,N_331,N_453);
nor U3801 (N_3801,N_165,N_265);
or U3802 (N_3802,N_876,N_2453);
or U3803 (N_3803,N_840,N_2481);
or U3804 (N_3804,N_1386,N_848);
or U3805 (N_3805,N_1352,N_1552);
xnor U3806 (N_3806,N_1059,N_1855);
and U3807 (N_3807,N_2104,N_2322);
nor U3808 (N_3808,N_1650,N_2221);
nand U3809 (N_3809,N_1988,N_329);
or U3810 (N_3810,N_371,N_407);
nor U3811 (N_3811,N_287,N_288);
nand U3812 (N_3812,N_2030,N_3);
nor U3813 (N_3813,N_2115,N_1143);
and U3814 (N_3814,N_1609,N_1724);
nand U3815 (N_3815,N_1684,N_1048);
nor U3816 (N_3816,N_1062,N_1064);
or U3817 (N_3817,N_1108,N_824);
nand U3818 (N_3818,N_2374,N_2158);
nor U3819 (N_3819,N_2241,N_622);
and U3820 (N_3820,N_1011,N_545);
and U3821 (N_3821,N_1527,N_2089);
or U3822 (N_3822,N_1673,N_2229);
nor U3823 (N_3823,N_2097,N_2283);
and U3824 (N_3824,N_1132,N_620);
nor U3825 (N_3825,N_703,N_2073);
nand U3826 (N_3826,N_89,N_2484);
nand U3827 (N_3827,N_2060,N_1070);
and U3828 (N_3828,N_1599,N_625);
nor U3829 (N_3829,N_598,N_429);
and U3830 (N_3830,N_183,N_1101);
and U3831 (N_3831,N_1888,N_453);
nand U3832 (N_3832,N_1361,N_2266);
nor U3833 (N_3833,N_1145,N_198);
nor U3834 (N_3834,N_98,N_286);
xnor U3835 (N_3835,N_1264,N_363);
and U3836 (N_3836,N_1533,N_953);
xor U3837 (N_3837,N_2018,N_551);
nand U3838 (N_3838,N_532,N_1434);
nand U3839 (N_3839,N_1630,N_2152);
and U3840 (N_3840,N_851,N_1077);
or U3841 (N_3841,N_1289,N_197);
nor U3842 (N_3842,N_914,N_1146);
nor U3843 (N_3843,N_1504,N_289);
nor U3844 (N_3844,N_457,N_1911);
nor U3845 (N_3845,N_1286,N_1416);
and U3846 (N_3846,N_81,N_1600);
and U3847 (N_3847,N_1371,N_2114);
nor U3848 (N_3848,N_620,N_1522);
nand U3849 (N_3849,N_1555,N_1566);
xor U3850 (N_3850,N_362,N_212);
xor U3851 (N_3851,N_2255,N_843);
nor U3852 (N_3852,N_227,N_2480);
or U3853 (N_3853,N_1899,N_1620);
and U3854 (N_3854,N_1945,N_1412);
xor U3855 (N_3855,N_1737,N_220);
or U3856 (N_3856,N_9,N_2476);
nand U3857 (N_3857,N_1039,N_2393);
or U3858 (N_3858,N_1269,N_2141);
or U3859 (N_3859,N_1841,N_1976);
or U3860 (N_3860,N_1086,N_1066);
nand U3861 (N_3861,N_340,N_931);
nand U3862 (N_3862,N_749,N_96);
and U3863 (N_3863,N_2251,N_2207);
and U3864 (N_3864,N_2290,N_1258);
nor U3865 (N_3865,N_2326,N_17);
or U3866 (N_3866,N_1886,N_1543);
xor U3867 (N_3867,N_349,N_215);
xnor U3868 (N_3868,N_2169,N_1990);
and U3869 (N_3869,N_2474,N_1565);
or U3870 (N_3870,N_2096,N_692);
or U3871 (N_3871,N_1312,N_506);
and U3872 (N_3872,N_318,N_2445);
and U3873 (N_3873,N_215,N_2485);
xnor U3874 (N_3874,N_1262,N_158);
or U3875 (N_3875,N_975,N_342);
nand U3876 (N_3876,N_1615,N_1119);
or U3877 (N_3877,N_411,N_155);
and U3878 (N_3878,N_550,N_1137);
nand U3879 (N_3879,N_2366,N_114);
nand U3880 (N_3880,N_2331,N_314);
nor U3881 (N_3881,N_765,N_2372);
nand U3882 (N_3882,N_646,N_2496);
and U3883 (N_3883,N_2469,N_2304);
nor U3884 (N_3884,N_1032,N_249);
xnor U3885 (N_3885,N_2339,N_2275);
and U3886 (N_3886,N_1903,N_115);
nand U3887 (N_3887,N_2099,N_1405);
nor U3888 (N_3888,N_530,N_1373);
or U3889 (N_3889,N_1761,N_494);
xor U3890 (N_3890,N_2376,N_301);
xor U3891 (N_3891,N_1374,N_363);
and U3892 (N_3892,N_2496,N_1212);
nor U3893 (N_3893,N_392,N_1450);
xnor U3894 (N_3894,N_80,N_205);
and U3895 (N_3895,N_434,N_1743);
xnor U3896 (N_3896,N_1606,N_1258);
and U3897 (N_3897,N_744,N_893);
xnor U3898 (N_3898,N_2248,N_814);
or U3899 (N_3899,N_337,N_2489);
or U3900 (N_3900,N_1063,N_1414);
or U3901 (N_3901,N_1867,N_2312);
or U3902 (N_3902,N_1660,N_2394);
nand U3903 (N_3903,N_2178,N_2102);
xor U3904 (N_3904,N_628,N_324);
nand U3905 (N_3905,N_1956,N_1375);
nor U3906 (N_3906,N_673,N_1171);
and U3907 (N_3907,N_506,N_2451);
nor U3908 (N_3908,N_466,N_1917);
xor U3909 (N_3909,N_2447,N_2499);
and U3910 (N_3910,N_2046,N_197);
and U3911 (N_3911,N_2461,N_2408);
nand U3912 (N_3912,N_442,N_291);
nor U3913 (N_3913,N_741,N_2132);
nor U3914 (N_3914,N_1910,N_463);
and U3915 (N_3915,N_211,N_1434);
and U3916 (N_3916,N_1259,N_643);
and U3917 (N_3917,N_145,N_1729);
nor U3918 (N_3918,N_612,N_871);
and U3919 (N_3919,N_2087,N_399);
nand U3920 (N_3920,N_443,N_1255);
nor U3921 (N_3921,N_528,N_1698);
nand U3922 (N_3922,N_568,N_137);
or U3923 (N_3923,N_2021,N_894);
and U3924 (N_3924,N_602,N_629);
nor U3925 (N_3925,N_2477,N_1470);
and U3926 (N_3926,N_334,N_1241);
nand U3927 (N_3927,N_1672,N_10);
xnor U3928 (N_3928,N_2167,N_2098);
and U3929 (N_3929,N_2104,N_696);
nor U3930 (N_3930,N_2369,N_2233);
xor U3931 (N_3931,N_395,N_265);
and U3932 (N_3932,N_1714,N_1095);
nor U3933 (N_3933,N_2109,N_149);
and U3934 (N_3934,N_924,N_564);
nand U3935 (N_3935,N_2258,N_166);
or U3936 (N_3936,N_478,N_934);
or U3937 (N_3937,N_1001,N_673);
or U3938 (N_3938,N_2314,N_79);
xnor U3939 (N_3939,N_2230,N_272);
and U3940 (N_3940,N_2166,N_1996);
nor U3941 (N_3941,N_641,N_1573);
or U3942 (N_3942,N_813,N_1717);
xnor U3943 (N_3943,N_678,N_6);
or U3944 (N_3944,N_1920,N_1938);
nor U3945 (N_3945,N_69,N_1046);
and U3946 (N_3946,N_603,N_1581);
and U3947 (N_3947,N_240,N_1180);
nor U3948 (N_3948,N_1437,N_618);
nor U3949 (N_3949,N_1868,N_1801);
xnor U3950 (N_3950,N_2199,N_836);
xnor U3951 (N_3951,N_2151,N_2343);
or U3952 (N_3952,N_518,N_484);
or U3953 (N_3953,N_1437,N_426);
nor U3954 (N_3954,N_2249,N_22);
nand U3955 (N_3955,N_2415,N_293);
or U3956 (N_3956,N_1462,N_812);
nand U3957 (N_3957,N_319,N_1481);
nand U3958 (N_3958,N_2101,N_2438);
and U3959 (N_3959,N_1884,N_2385);
nand U3960 (N_3960,N_1010,N_383);
xor U3961 (N_3961,N_332,N_2231);
and U3962 (N_3962,N_627,N_618);
nand U3963 (N_3963,N_2345,N_777);
xor U3964 (N_3964,N_998,N_313);
or U3965 (N_3965,N_1411,N_2362);
and U3966 (N_3966,N_1340,N_382);
nor U3967 (N_3967,N_2166,N_1293);
and U3968 (N_3968,N_232,N_1669);
or U3969 (N_3969,N_553,N_1462);
nand U3970 (N_3970,N_1411,N_1245);
or U3971 (N_3971,N_1808,N_495);
or U3972 (N_3972,N_41,N_1793);
nand U3973 (N_3973,N_1281,N_2105);
xor U3974 (N_3974,N_1094,N_1951);
and U3975 (N_3975,N_2246,N_2390);
xor U3976 (N_3976,N_469,N_653);
and U3977 (N_3977,N_1402,N_39);
or U3978 (N_3978,N_1707,N_1005);
xnor U3979 (N_3979,N_1110,N_255);
nor U3980 (N_3980,N_1323,N_2315);
and U3981 (N_3981,N_1378,N_2423);
xor U3982 (N_3982,N_2204,N_500);
and U3983 (N_3983,N_770,N_1430);
nor U3984 (N_3984,N_690,N_1103);
and U3985 (N_3985,N_1486,N_1772);
nor U3986 (N_3986,N_688,N_1756);
nor U3987 (N_3987,N_1543,N_1724);
and U3988 (N_3988,N_1634,N_1200);
and U3989 (N_3989,N_381,N_1593);
nand U3990 (N_3990,N_1640,N_1367);
or U3991 (N_3991,N_2090,N_1615);
and U3992 (N_3992,N_1445,N_1319);
and U3993 (N_3993,N_853,N_365);
or U3994 (N_3994,N_119,N_1628);
xnor U3995 (N_3995,N_2482,N_740);
nand U3996 (N_3996,N_1979,N_938);
and U3997 (N_3997,N_360,N_2287);
or U3998 (N_3998,N_901,N_2235);
or U3999 (N_3999,N_330,N_1854);
nor U4000 (N_4000,N_1279,N_1258);
and U4001 (N_4001,N_1149,N_1101);
nand U4002 (N_4002,N_584,N_303);
or U4003 (N_4003,N_250,N_1887);
and U4004 (N_4004,N_1816,N_752);
xor U4005 (N_4005,N_917,N_585);
nor U4006 (N_4006,N_1221,N_614);
xnor U4007 (N_4007,N_154,N_1546);
or U4008 (N_4008,N_297,N_1531);
or U4009 (N_4009,N_870,N_719);
xnor U4010 (N_4010,N_2179,N_969);
nor U4011 (N_4011,N_2210,N_1356);
and U4012 (N_4012,N_2397,N_50);
or U4013 (N_4013,N_86,N_2331);
nand U4014 (N_4014,N_389,N_1346);
nor U4015 (N_4015,N_964,N_1092);
nor U4016 (N_4016,N_1771,N_511);
and U4017 (N_4017,N_735,N_2021);
nand U4018 (N_4018,N_1672,N_2070);
xnor U4019 (N_4019,N_1631,N_386);
nor U4020 (N_4020,N_2386,N_934);
xor U4021 (N_4021,N_959,N_794);
or U4022 (N_4022,N_2258,N_868);
nand U4023 (N_4023,N_1998,N_754);
xnor U4024 (N_4024,N_2492,N_1402);
and U4025 (N_4025,N_1891,N_2121);
nor U4026 (N_4026,N_2345,N_381);
nor U4027 (N_4027,N_2269,N_1262);
nor U4028 (N_4028,N_2068,N_834);
xnor U4029 (N_4029,N_1732,N_2298);
nor U4030 (N_4030,N_337,N_662);
and U4031 (N_4031,N_146,N_2410);
or U4032 (N_4032,N_679,N_2009);
nor U4033 (N_4033,N_715,N_976);
or U4034 (N_4034,N_1567,N_432);
xnor U4035 (N_4035,N_2016,N_1192);
nor U4036 (N_4036,N_2017,N_1573);
xnor U4037 (N_4037,N_236,N_2149);
nand U4038 (N_4038,N_1410,N_2009);
or U4039 (N_4039,N_870,N_1625);
nor U4040 (N_4040,N_438,N_1707);
or U4041 (N_4041,N_1069,N_1327);
nand U4042 (N_4042,N_1422,N_611);
nor U4043 (N_4043,N_1624,N_2104);
nor U4044 (N_4044,N_801,N_1445);
xor U4045 (N_4045,N_1279,N_296);
nor U4046 (N_4046,N_1187,N_424);
and U4047 (N_4047,N_1008,N_1562);
nand U4048 (N_4048,N_1085,N_340);
and U4049 (N_4049,N_632,N_1499);
nand U4050 (N_4050,N_2192,N_277);
nor U4051 (N_4051,N_1131,N_1746);
nor U4052 (N_4052,N_761,N_2393);
or U4053 (N_4053,N_913,N_655);
nor U4054 (N_4054,N_271,N_2314);
or U4055 (N_4055,N_1608,N_2490);
or U4056 (N_4056,N_2006,N_1954);
or U4057 (N_4057,N_126,N_1459);
and U4058 (N_4058,N_802,N_164);
nor U4059 (N_4059,N_424,N_577);
or U4060 (N_4060,N_26,N_1693);
xor U4061 (N_4061,N_2263,N_1397);
nor U4062 (N_4062,N_661,N_621);
or U4063 (N_4063,N_2231,N_1715);
or U4064 (N_4064,N_1576,N_1334);
or U4065 (N_4065,N_19,N_506);
and U4066 (N_4066,N_2214,N_1041);
nor U4067 (N_4067,N_1421,N_1574);
or U4068 (N_4068,N_2082,N_1092);
and U4069 (N_4069,N_625,N_364);
and U4070 (N_4070,N_2249,N_484);
nor U4071 (N_4071,N_447,N_696);
xor U4072 (N_4072,N_197,N_1556);
nor U4073 (N_4073,N_1849,N_1525);
nand U4074 (N_4074,N_1708,N_1047);
nor U4075 (N_4075,N_831,N_2300);
xor U4076 (N_4076,N_1428,N_2384);
nor U4077 (N_4077,N_56,N_1604);
nor U4078 (N_4078,N_955,N_894);
xnor U4079 (N_4079,N_1006,N_2439);
xnor U4080 (N_4080,N_241,N_879);
nand U4081 (N_4081,N_883,N_1377);
nand U4082 (N_4082,N_2329,N_567);
and U4083 (N_4083,N_1645,N_1263);
and U4084 (N_4084,N_222,N_885);
and U4085 (N_4085,N_258,N_1322);
or U4086 (N_4086,N_316,N_700);
and U4087 (N_4087,N_1957,N_286);
nand U4088 (N_4088,N_73,N_377);
nand U4089 (N_4089,N_2211,N_662);
or U4090 (N_4090,N_1189,N_1103);
nand U4091 (N_4091,N_298,N_2413);
nand U4092 (N_4092,N_1570,N_1455);
and U4093 (N_4093,N_153,N_1225);
and U4094 (N_4094,N_1550,N_1977);
nand U4095 (N_4095,N_506,N_1357);
and U4096 (N_4096,N_1752,N_182);
xnor U4097 (N_4097,N_945,N_759);
nand U4098 (N_4098,N_1372,N_1440);
or U4099 (N_4099,N_11,N_1363);
nand U4100 (N_4100,N_1804,N_1631);
and U4101 (N_4101,N_1913,N_250);
and U4102 (N_4102,N_353,N_343);
xnor U4103 (N_4103,N_255,N_1087);
and U4104 (N_4104,N_1178,N_1303);
or U4105 (N_4105,N_2067,N_526);
nor U4106 (N_4106,N_137,N_1615);
xnor U4107 (N_4107,N_23,N_1593);
and U4108 (N_4108,N_2309,N_455);
and U4109 (N_4109,N_1367,N_1823);
xnor U4110 (N_4110,N_323,N_1519);
xnor U4111 (N_4111,N_1534,N_867);
or U4112 (N_4112,N_1206,N_2243);
nand U4113 (N_4113,N_1980,N_1468);
xnor U4114 (N_4114,N_16,N_1611);
nand U4115 (N_4115,N_2156,N_999);
nor U4116 (N_4116,N_1627,N_1329);
nor U4117 (N_4117,N_1006,N_388);
nand U4118 (N_4118,N_1949,N_735);
nor U4119 (N_4119,N_610,N_1379);
nor U4120 (N_4120,N_1188,N_2383);
nor U4121 (N_4121,N_1422,N_2346);
or U4122 (N_4122,N_1715,N_1341);
and U4123 (N_4123,N_2268,N_420);
xnor U4124 (N_4124,N_1736,N_1018);
and U4125 (N_4125,N_903,N_2006);
nor U4126 (N_4126,N_1176,N_2239);
and U4127 (N_4127,N_1283,N_1583);
and U4128 (N_4128,N_2071,N_1666);
or U4129 (N_4129,N_1729,N_1316);
xor U4130 (N_4130,N_560,N_251);
and U4131 (N_4131,N_1010,N_579);
xor U4132 (N_4132,N_1328,N_2166);
or U4133 (N_4133,N_1259,N_1596);
and U4134 (N_4134,N_1394,N_1447);
nand U4135 (N_4135,N_1491,N_354);
or U4136 (N_4136,N_1763,N_1160);
or U4137 (N_4137,N_79,N_2008);
and U4138 (N_4138,N_1584,N_312);
nand U4139 (N_4139,N_168,N_346);
nand U4140 (N_4140,N_475,N_1756);
or U4141 (N_4141,N_2018,N_326);
xor U4142 (N_4142,N_1383,N_1050);
and U4143 (N_4143,N_309,N_1004);
or U4144 (N_4144,N_552,N_2242);
nor U4145 (N_4145,N_1056,N_1035);
and U4146 (N_4146,N_1309,N_389);
or U4147 (N_4147,N_467,N_415);
and U4148 (N_4148,N_627,N_1803);
nor U4149 (N_4149,N_1274,N_785);
nor U4150 (N_4150,N_2310,N_2087);
and U4151 (N_4151,N_1271,N_862);
nor U4152 (N_4152,N_354,N_1251);
xnor U4153 (N_4153,N_1277,N_532);
and U4154 (N_4154,N_1744,N_2465);
and U4155 (N_4155,N_308,N_1431);
nand U4156 (N_4156,N_2055,N_964);
or U4157 (N_4157,N_2133,N_609);
and U4158 (N_4158,N_1696,N_1907);
nand U4159 (N_4159,N_1753,N_663);
xor U4160 (N_4160,N_2191,N_106);
and U4161 (N_4161,N_1529,N_424);
and U4162 (N_4162,N_219,N_215);
nand U4163 (N_4163,N_177,N_1504);
xor U4164 (N_4164,N_864,N_915);
nor U4165 (N_4165,N_529,N_2322);
nor U4166 (N_4166,N_1555,N_2090);
xor U4167 (N_4167,N_615,N_292);
and U4168 (N_4168,N_1054,N_1340);
and U4169 (N_4169,N_822,N_281);
nand U4170 (N_4170,N_865,N_1601);
nand U4171 (N_4171,N_1529,N_1619);
or U4172 (N_4172,N_1893,N_998);
or U4173 (N_4173,N_1992,N_1593);
xor U4174 (N_4174,N_2402,N_1855);
and U4175 (N_4175,N_1956,N_340);
nor U4176 (N_4176,N_2343,N_1977);
xnor U4177 (N_4177,N_43,N_1124);
nor U4178 (N_4178,N_1511,N_1883);
or U4179 (N_4179,N_1428,N_1780);
nand U4180 (N_4180,N_1541,N_2011);
nor U4181 (N_4181,N_2429,N_1461);
nand U4182 (N_4182,N_1306,N_2399);
nor U4183 (N_4183,N_2289,N_1656);
and U4184 (N_4184,N_1766,N_1316);
and U4185 (N_4185,N_2318,N_992);
and U4186 (N_4186,N_2395,N_1944);
nand U4187 (N_4187,N_1097,N_805);
nand U4188 (N_4188,N_59,N_2290);
and U4189 (N_4189,N_1676,N_2473);
and U4190 (N_4190,N_1550,N_455);
xnor U4191 (N_4191,N_793,N_2356);
and U4192 (N_4192,N_580,N_118);
and U4193 (N_4193,N_1495,N_1336);
xor U4194 (N_4194,N_2437,N_1898);
nor U4195 (N_4195,N_1851,N_1805);
nand U4196 (N_4196,N_2277,N_481);
nor U4197 (N_4197,N_49,N_1524);
xor U4198 (N_4198,N_2275,N_612);
and U4199 (N_4199,N_577,N_2105);
nand U4200 (N_4200,N_2188,N_2054);
xor U4201 (N_4201,N_381,N_489);
xnor U4202 (N_4202,N_715,N_914);
nor U4203 (N_4203,N_499,N_1332);
nand U4204 (N_4204,N_1331,N_1515);
and U4205 (N_4205,N_1325,N_809);
xnor U4206 (N_4206,N_2002,N_899);
or U4207 (N_4207,N_2342,N_13);
nor U4208 (N_4208,N_380,N_529);
or U4209 (N_4209,N_1951,N_1919);
nand U4210 (N_4210,N_1106,N_1802);
and U4211 (N_4211,N_1171,N_1435);
nand U4212 (N_4212,N_602,N_1838);
nor U4213 (N_4213,N_2199,N_917);
xnor U4214 (N_4214,N_1083,N_1719);
or U4215 (N_4215,N_1070,N_2470);
xor U4216 (N_4216,N_1134,N_1023);
and U4217 (N_4217,N_368,N_1513);
nand U4218 (N_4218,N_477,N_2055);
or U4219 (N_4219,N_873,N_1275);
xor U4220 (N_4220,N_1233,N_1048);
nand U4221 (N_4221,N_793,N_790);
xor U4222 (N_4222,N_672,N_1717);
xnor U4223 (N_4223,N_2259,N_1032);
and U4224 (N_4224,N_1663,N_2154);
xnor U4225 (N_4225,N_2407,N_1848);
xnor U4226 (N_4226,N_350,N_1091);
xor U4227 (N_4227,N_1647,N_1979);
and U4228 (N_4228,N_1269,N_2322);
or U4229 (N_4229,N_1323,N_2089);
nand U4230 (N_4230,N_31,N_440);
xor U4231 (N_4231,N_964,N_1899);
or U4232 (N_4232,N_902,N_1228);
xor U4233 (N_4233,N_282,N_1795);
nand U4234 (N_4234,N_2470,N_875);
or U4235 (N_4235,N_2239,N_951);
or U4236 (N_4236,N_1795,N_201);
nor U4237 (N_4237,N_1931,N_578);
nor U4238 (N_4238,N_1782,N_2363);
nand U4239 (N_4239,N_2113,N_1304);
and U4240 (N_4240,N_2071,N_1133);
xor U4241 (N_4241,N_2137,N_1817);
or U4242 (N_4242,N_1337,N_1971);
and U4243 (N_4243,N_1768,N_227);
and U4244 (N_4244,N_1592,N_2249);
nand U4245 (N_4245,N_2103,N_1004);
or U4246 (N_4246,N_329,N_365);
xnor U4247 (N_4247,N_449,N_101);
nor U4248 (N_4248,N_1912,N_1322);
nand U4249 (N_4249,N_197,N_1892);
xnor U4250 (N_4250,N_1631,N_1977);
xnor U4251 (N_4251,N_1695,N_3);
nor U4252 (N_4252,N_158,N_630);
nand U4253 (N_4253,N_2358,N_1536);
and U4254 (N_4254,N_126,N_2);
nor U4255 (N_4255,N_2220,N_1784);
xor U4256 (N_4256,N_1992,N_94);
nor U4257 (N_4257,N_1840,N_2277);
or U4258 (N_4258,N_1359,N_1260);
xor U4259 (N_4259,N_456,N_640);
or U4260 (N_4260,N_1116,N_1350);
xnor U4261 (N_4261,N_758,N_874);
xor U4262 (N_4262,N_1627,N_1837);
or U4263 (N_4263,N_2385,N_1772);
nor U4264 (N_4264,N_612,N_801);
and U4265 (N_4265,N_1908,N_1867);
nor U4266 (N_4266,N_1683,N_1941);
nor U4267 (N_4267,N_381,N_1442);
and U4268 (N_4268,N_2049,N_1983);
or U4269 (N_4269,N_1475,N_2100);
nand U4270 (N_4270,N_649,N_2372);
or U4271 (N_4271,N_976,N_1513);
and U4272 (N_4272,N_901,N_619);
nor U4273 (N_4273,N_1642,N_200);
or U4274 (N_4274,N_2241,N_1995);
or U4275 (N_4275,N_1717,N_1512);
xor U4276 (N_4276,N_1522,N_1801);
or U4277 (N_4277,N_1164,N_2138);
nand U4278 (N_4278,N_398,N_676);
nor U4279 (N_4279,N_1816,N_67);
or U4280 (N_4280,N_2075,N_1482);
and U4281 (N_4281,N_1276,N_1256);
and U4282 (N_4282,N_1101,N_2291);
xor U4283 (N_4283,N_343,N_949);
or U4284 (N_4284,N_383,N_28);
or U4285 (N_4285,N_1957,N_636);
xnor U4286 (N_4286,N_637,N_1384);
or U4287 (N_4287,N_892,N_2354);
nand U4288 (N_4288,N_539,N_1032);
xor U4289 (N_4289,N_386,N_121);
xnor U4290 (N_4290,N_2490,N_1292);
nand U4291 (N_4291,N_2258,N_1694);
nand U4292 (N_4292,N_1966,N_1330);
nand U4293 (N_4293,N_1760,N_377);
nor U4294 (N_4294,N_1575,N_502);
nand U4295 (N_4295,N_1806,N_795);
and U4296 (N_4296,N_281,N_1502);
nand U4297 (N_4297,N_744,N_568);
nor U4298 (N_4298,N_2405,N_2320);
nor U4299 (N_4299,N_243,N_949);
and U4300 (N_4300,N_1351,N_83);
and U4301 (N_4301,N_707,N_2034);
or U4302 (N_4302,N_194,N_996);
nor U4303 (N_4303,N_1579,N_1123);
nand U4304 (N_4304,N_416,N_1315);
nand U4305 (N_4305,N_2437,N_751);
or U4306 (N_4306,N_1033,N_981);
nand U4307 (N_4307,N_137,N_376);
or U4308 (N_4308,N_327,N_1659);
xor U4309 (N_4309,N_486,N_1464);
xor U4310 (N_4310,N_1040,N_2118);
nand U4311 (N_4311,N_887,N_993);
or U4312 (N_4312,N_1319,N_741);
or U4313 (N_4313,N_9,N_1102);
or U4314 (N_4314,N_856,N_279);
and U4315 (N_4315,N_1449,N_211);
nor U4316 (N_4316,N_2466,N_2420);
nand U4317 (N_4317,N_1816,N_1411);
nand U4318 (N_4318,N_919,N_2101);
nand U4319 (N_4319,N_1987,N_1448);
nand U4320 (N_4320,N_214,N_1624);
xnor U4321 (N_4321,N_1154,N_1407);
nor U4322 (N_4322,N_435,N_2161);
nor U4323 (N_4323,N_105,N_835);
nand U4324 (N_4324,N_2367,N_496);
xnor U4325 (N_4325,N_811,N_1922);
nand U4326 (N_4326,N_443,N_2400);
and U4327 (N_4327,N_839,N_2078);
and U4328 (N_4328,N_317,N_2429);
and U4329 (N_4329,N_1519,N_2289);
or U4330 (N_4330,N_290,N_837);
nand U4331 (N_4331,N_2089,N_1178);
nor U4332 (N_4332,N_509,N_946);
xor U4333 (N_4333,N_1430,N_884);
nor U4334 (N_4334,N_1312,N_995);
or U4335 (N_4335,N_10,N_2452);
nor U4336 (N_4336,N_665,N_462);
xnor U4337 (N_4337,N_103,N_6);
and U4338 (N_4338,N_183,N_931);
nand U4339 (N_4339,N_492,N_2276);
xor U4340 (N_4340,N_1017,N_793);
and U4341 (N_4341,N_1561,N_2089);
xnor U4342 (N_4342,N_116,N_1339);
or U4343 (N_4343,N_790,N_1111);
nand U4344 (N_4344,N_131,N_1786);
nor U4345 (N_4345,N_2423,N_1878);
nand U4346 (N_4346,N_1304,N_2381);
nand U4347 (N_4347,N_791,N_593);
nand U4348 (N_4348,N_1079,N_536);
xor U4349 (N_4349,N_2216,N_82);
xor U4350 (N_4350,N_1594,N_2100);
and U4351 (N_4351,N_268,N_1177);
nor U4352 (N_4352,N_226,N_324);
or U4353 (N_4353,N_2279,N_426);
nand U4354 (N_4354,N_1748,N_536);
nand U4355 (N_4355,N_411,N_741);
nand U4356 (N_4356,N_1088,N_1810);
nand U4357 (N_4357,N_574,N_1918);
nor U4358 (N_4358,N_470,N_971);
nor U4359 (N_4359,N_1288,N_465);
nand U4360 (N_4360,N_2261,N_1727);
nor U4361 (N_4361,N_336,N_1445);
and U4362 (N_4362,N_70,N_2454);
or U4363 (N_4363,N_1378,N_2364);
or U4364 (N_4364,N_2175,N_1815);
nand U4365 (N_4365,N_686,N_1471);
nand U4366 (N_4366,N_461,N_454);
nor U4367 (N_4367,N_1422,N_1973);
or U4368 (N_4368,N_91,N_1935);
or U4369 (N_4369,N_2017,N_2476);
or U4370 (N_4370,N_817,N_1103);
and U4371 (N_4371,N_1676,N_486);
nand U4372 (N_4372,N_868,N_671);
or U4373 (N_4373,N_2195,N_1162);
xor U4374 (N_4374,N_1486,N_866);
or U4375 (N_4375,N_1716,N_784);
xnor U4376 (N_4376,N_174,N_1669);
or U4377 (N_4377,N_899,N_325);
nor U4378 (N_4378,N_500,N_1586);
nor U4379 (N_4379,N_1224,N_1800);
xor U4380 (N_4380,N_1891,N_138);
or U4381 (N_4381,N_190,N_1147);
or U4382 (N_4382,N_2267,N_84);
nand U4383 (N_4383,N_1716,N_1148);
nand U4384 (N_4384,N_1095,N_1485);
nand U4385 (N_4385,N_904,N_289);
nor U4386 (N_4386,N_2313,N_2339);
nor U4387 (N_4387,N_1974,N_373);
or U4388 (N_4388,N_285,N_1984);
nand U4389 (N_4389,N_889,N_2174);
nor U4390 (N_4390,N_1301,N_1746);
xor U4391 (N_4391,N_644,N_997);
nand U4392 (N_4392,N_1590,N_2414);
nor U4393 (N_4393,N_2244,N_2364);
and U4394 (N_4394,N_1299,N_8);
nor U4395 (N_4395,N_2182,N_1761);
or U4396 (N_4396,N_1677,N_126);
nor U4397 (N_4397,N_735,N_1969);
nor U4398 (N_4398,N_148,N_2440);
nor U4399 (N_4399,N_2470,N_1452);
xnor U4400 (N_4400,N_2070,N_1744);
or U4401 (N_4401,N_1129,N_339);
xor U4402 (N_4402,N_805,N_81);
or U4403 (N_4403,N_377,N_1452);
or U4404 (N_4404,N_1634,N_285);
xnor U4405 (N_4405,N_2242,N_2348);
nand U4406 (N_4406,N_710,N_2253);
or U4407 (N_4407,N_347,N_1563);
nor U4408 (N_4408,N_161,N_13);
xor U4409 (N_4409,N_2026,N_1072);
nand U4410 (N_4410,N_1084,N_650);
nand U4411 (N_4411,N_894,N_412);
xor U4412 (N_4412,N_390,N_2204);
xor U4413 (N_4413,N_1441,N_182);
nor U4414 (N_4414,N_720,N_1300);
nor U4415 (N_4415,N_1124,N_2257);
nand U4416 (N_4416,N_316,N_167);
xor U4417 (N_4417,N_1207,N_37);
nor U4418 (N_4418,N_1696,N_1842);
nand U4419 (N_4419,N_1987,N_334);
and U4420 (N_4420,N_1037,N_1690);
or U4421 (N_4421,N_346,N_881);
nand U4422 (N_4422,N_696,N_1625);
nand U4423 (N_4423,N_2487,N_1005);
and U4424 (N_4424,N_1804,N_1578);
or U4425 (N_4425,N_1680,N_1499);
xor U4426 (N_4426,N_2473,N_150);
or U4427 (N_4427,N_538,N_2087);
and U4428 (N_4428,N_396,N_2171);
or U4429 (N_4429,N_1278,N_480);
and U4430 (N_4430,N_1417,N_2409);
xor U4431 (N_4431,N_788,N_1651);
nor U4432 (N_4432,N_1603,N_118);
nor U4433 (N_4433,N_1230,N_2490);
nand U4434 (N_4434,N_1788,N_1524);
and U4435 (N_4435,N_1440,N_167);
xor U4436 (N_4436,N_224,N_1470);
nor U4437 (N_4437,N_1954,N_124);
xor U4438 (N_4438,N_2390,N_1288);
xnor U4439 (N_4439,N_2079,N_1611);
or U4440 (N_4440,N_2026,N_2323);
xnor U4441 (N_4441,N_790,N_631);
or U4442 (N_4442,N_758,N_44);
xor U4443 (N_4443,N_1339,N_1304);
nor U4444 (N_4444,N_618,N_1535);
nand U4445 (N_4445,N_1801,N_1776);
or U4446 (N_4446,N_2395,N_540);
or U4447 (N_4447,N_1465,N_22);
nand U4448 (N_4448,N_843,N_706);
nor U4449 (N_4449,N_209,N_2340);
or U4450 (N_4450,N_1164,N_372);
nand U4451 (N_4451,N_2227,N_486);
nor U4452 (N_4452,N_2426,N_1057);
nand U4453 (N_4453,N_345,N_2223);
or U4454 (N_4454,N_1974,N_1597);
xor U4455 (N_4455,N_310,N_1651);
nor U4456 (N_4456,N_236,N_159);
or U4457 (N_4457,N_924,N_673);
and U4458 (N_4458,N_402,N_940);
nor U4459 (N_4459,N_76,N_592);
and U4460 (N_4460,N_629,N_2465);
nand U4461 (N_4461,N_809,N_2237);
xor U4462 (N_4462,N_530,N_410);
or U4463 (N_4463,N_364,N_2084);
or U4464 (N_4464,N_1362,N_1000);
nor U4465 (N_4465,N_1788,N_2220);
xnor U4466 (N_4466,N_0,N_1248);
nor U4467 (N_4467,N_610,N_1206);
nand U4468 (N_4468,N_1617,N_1196);
nor U4469 (N_4469,N_1505,N_1435);
or U4470 (N_4470,N_1709,N_217);
or U4471 (N_4471,N_186,N_1462);
nor U4472 (N_4472,N_1674,N_1211);
nand U4473 (N_4473,N_2321,N_1395);
and U4474 (N_4474,N_826,N_443);
nand U4475 (N_4475,N_2486,N_2494);
xnor U4476 (N_4476,N_302,N_1632);
xor U4477 (N_4477,N_850,N_1378);
or U4478 (N_4478,N_897,N_46);
nor U4479 (N_4479,N_2403,N_60);
nand U4480 (N_4480,N_1390,N_2033);
nor U4481 (N_4481,N_2287,N_1684);
or U4482 (N_4482,N_197,N_2164);
nand U4483 (N_4483,N_771,N_1679);
nand U4484 (N_4484,N_2310,N_2104);
nand U4485 (N_4485,N_297,N_2416);
or U4486 (N_4486,N_234,N_1848);
nand U4487 (N_4487,N_1384,N_1336);
nand U4488 (N_4488,N_1478,N_329);
nor U4489 (N_4489,N_155,N_953);
nand U4490 (N_4490,N_114,N_552);
and U4491 (N_4491,N_1234,N_306);
nand U4492 (N_4492,N_881,N_882);
nor U4493 (N_4493,N_479,N_619);
nand U4494 (N_4494,N_1723,N_1527);
nor U4495 (N_4495,N_1046,N_502);
or U4496 (N_4496,N_1712,N_2416);
nor U4497 (N_4497,N_1676,N_2288);
and U4498 (N_4498,N_111,N_1193);
or U4499 (N_4499,N_783,N_2280);
nand U4500 (N_4500,N_1187,N_1407);
xor U4501 (N_4501,N_1624,N_669);
nor U4502 (N_4502,N_1467,N_1129);
or U4503 (N_4503,N_625,N_384);
xor U4504 (N_4504,N_1034,N_1123);
and U4505 (N_4505,N_2402,N_1389);
nand U4506 (N_4506,N_2315,N_344);
and U4507 (N_4507,N_996,N_420);
and U4508 (N_4508,N_1847,N_1435);
nand U4509 (N_4509,N_1702,N_241);
xnor U4510 (N_4510,N_99,N_1901);
or U4511 (N_4511,N_1621,N_563);
and U4512 (N_4512,N_649,N_273);
nor U4513 (N_4513,N_1542,N_1965);
and U4514 (N_4514,N_331,N_1001);
nand U4515 (N_4515,N_2092,N_1007);
or U4516 (N_4516,N_518,N_45);
nor U4517 (N_4517,N_2441,N_2036);
and U4518 (N_4518,N_2317,N_1950);
nor U4519 (N_4519,N_1500,N_369);
nor U4520 (N_4520,N_2313,N_2377);
or U4521 (N_4521,N_872,N_2214);
xor U4522 (N_4522,N_2464,N_1874);
xnor U4523 (N_4523,N_2059,N_1055);
nor U4524 (N_4524,N_2114,N_1743);
and U4525 (N_4525,N_1524,N_240);
xor U4526 (N_4526,N_2359,N_619);
or U4527 (N_4527,N_1036,N_1465);
xnor U4528 (N_4528,N_1528,N_2138);
nand U4529 (N_4529,N_776,N_2094);
nor U4530 (N_4530,N_1454,N_571);
nand U4531 (N_4531,N_913,N_430);
nor U4532 (N_4532,N_490,N_359);
xor U4533 (N_4533,N_1871,N_2080);
xor U4534 (N_4534,N_1800,N_381);
or U4535 (N_4535,N_793,N_35);
nand U4536 (N_4536,N_1899,N_1248);
xor U4537 (N_4537,N_2187,N_2311);
nand U4538 (N_4538,N_1894,N_1847);
nand U4539 (N_4539,N_1002,N_1864);
or U4540 (N_4540,N_1971,N_863);
nand U4541 (N_4541,N_902,N_525);
nor U4542 (N_4542,N_118,N_804);
xnor U4543 (N_4543,N_1541,N_219);
or U4544 (N_4544,N_1194,N_632);
and U4545 (N_4545,N_2146,N_2434);
xnor U4546 (N_4546,N_1671,N_1546);
xnor U4547 (N_4547,N_679,N_2366);
and U4548 (N_4548,N_1302,N_1771);
nor U4549 (N_4549,N_1510,N_544);
or U4550 (N_4550,N_2400,N_2237);
nor U4551 (N_4551,N_2003,N_418);
nand U4552 (N_4552,N_1811,N_1870);
nor U4553 (N_4553,N_549,N_431);
xnor U4554 (N_4554,N_96,N_82);
nor U4555 (N_4555,N_872,N_2341);
and U4556 (N_4556,N_258,N_1334);
nand U4557 (N_4557,N_1904,N_657);
and U4558 (N_4558,N_421,N_1623);
nor U4559 (N_4559,N_875,N_1299);
and U4560 (N_4560,N_1880,N_2429);
nor U4561 (N_4561,N_528,N_1343);
xnor U4562 (N_4562,N_400,N_1637);
or U4563 (N_4563,N_1975,N_1260);
nand U4564 (N_4564,N_775,N_1761);
or U4565 (N_4565,N_306,N_2266);
xnor U4566 (N_4566,N_2040,N_1028);
and U4567 (N_4567,N_1834,N_2337);
xnor U4568 (N_4568,N_116,N_2245);
and U4569 (N_4569,N_254,N_2207);
nor U4570 (N_4570,N_461,N_1475);
nand U4571 (N_4571,N_238,N_823);
xor U4572 (N_4572,N_890,N_1017);
and U4573 (N_4573,N_1084,N_2490);
and U4574 (N_4574,N_389,N_1208);
nor U4575 (N_4575,N_1804,N_1024);
xor U4576 (N_4576,N_2066,N_215);
nor U4577 (N_4577,N_574,N_595);
xor U4578 (N_4578,N_1905,N_331);
and U4579 (N_4579,N_1527,N_2171);
xor U4580 (N_4580,N_1200,N_372);
nand U4581 (N_4581,N_1830,N_2128);
nand U4582 (N_4582,N_1822,N_1111);
xnor U4583 (N_4583,N_1892,N_433);
or U4584 (N_4584,N_1449,N_185);
or U4585 (N_4585,N_537,N_1736);
xnor U4586 (N_4586,N_523,N_2305);
nand U4587 (N_4587,N_363,N_2481);
and U4588 (N_4588,N_1492,N_92);
nand U4589 (N_4589,N_1373,N_1737);
nand U4590 (N_4590,N_1295,N_1366);
and U4591 (N_4591,N_363,N_1600);
nor U4592 (N_4592,N_797,N_2026);
xnor U4593 (N_4593,N_1654,N_2335);
nor U4594 (N_4594,N_459,N_2143);
nor U4595 (N_4595,N_761,N_571);
xnor U4596 (N_4596,N_709,N_777);
or U4597 (N_4597,N_87,N_1966);
and U4598 (N_4598,N_112,N_781);
xor U4599 (N_4599,N_74,N_1249);
xnor U4600 (N_4600,N_134,N_923);
or U4601 (N_4601,N_784,N_1841);
or U4602 (N_4602,N_948,N_942);
or U4603 (N_4603,N_840,N_1417);
nand U4604 (N_4604,N_421,N_363);
nand U4605 (N_4605,N_2228,N_1672);
nand U4606 (N_4606,N_2384,N_872);
and U4607 (N_4607,N_1476,N_644);
nand U4608 (N_4608,N_1286,N_1889);
xnor U4609 (N_4609,N_1459,N_2210);
nor U4610 (N_4610,N_2389,N_1233);
or U4611 (N_4611,N_1314,N_948);
nand U4612 (N_4612,N_1252,N_2232);
or U4613 (N_4613,N_491,N_1830);
nand U4614 (N_4614,N_713,N_2180);
xor U4615 (N_4615,N_497,N_1593);
nor U4616 (N_4616,N_797,N_217);
nand U4617 (N_4617,N_1044,N_1225);
or U4618 (N_4618,N_530,N_1955);
or U4619 (N_4619,N_470,N_1746);
nor U4620 (N_4620,N_1720,N_1594);
nor U4621 (N_4621,N_1190,N_1492);
and U4622 (N_4622,N_299,N_207);
nand U4623 (N_4623,N_174,N_1011);
and U4624 (N_4624,N_2164,N_1525);
xnor U4625 (N_4625,N_1483,N_1493);
nor U4626 (N_4626,N_1962,N_2301);
and U4627 (N_4627,N_1505,N_1067);
nor U4628 (N_4628,N_1882,N_45);
nor U4629 (N_4629,N_1015,N_1154);
or U4630 (N_4630,N_1051,N_1025);
and U4631 (N_4631,N_1919,N_1809);
and U4632 (N_4632,N_312,N_1448);
and U4633 (N_4633,N_2242,N_103);
xnor U4634 (N_4634,N_193,N_261);
xor U4635 (N_4635,N_1923,N_2214);
nand U4636 (N_4636,N_1892,N_1583);
xnor U4637 (N_4637,N_657,N_897);
nor U4638 (N_4638,N_1600,N_2184);
nand U4639 (N_4639,N_374,N_1209);
and U4640 (N_4640,N_1957,N_2165);
nand U4641 (N_4641,N_469,N_795);
xor U4642 (N_4642,N_609,N_1175);
nand U4643 (N_4643,N_1168,N_817);
xor U4644 (N_4644,N_1855,N_1254);
nand U4645 (N_4645,N_710,N_2332);
nand U4646 (N_4646,N_960,N_812);
or U4647 (N_4647,N_1205,N_720);
or U4648 (N_4648,N_946,N_2362);
or U4649 (N_4649,N_2263,N_1822);
nand U4650 (N_4650,N_2000,N_1075);
nor U4651 (N_4651,N_754,N_310);
nor U4652 (N_4652,N_980,N_127);
nand U4653 (N_4653,N_1441,N_1963);
xor U4654 (N_4654,N_290,N_1162);
nor U4655 (N_4655,N_1508,N_136);
xor U4656 (N_4656,N_1155,N_1116);
nand U4657 (N_4657,N_313,N_1194);
nor U4658 (N_4658,N_813,N_807);
xor U4659 (N_4659,N_1845,N_1113);
xnor U4660 (N_4660,N_1489,N_354);
xor U4661 (N_4661,N_200,N_1074);
and U4662 (N_4662,N_2384,N_1625);
or U4663 (N_4663,N_1375,N_1092);
nor U4664 (N_4664,N_391,N_1821);
nor U4665 (N_4665,N_1697,N_1046);
and U4666 (N_4666,N_2021,N_749);
or U4667 (N_4667,N_724,N_2250);
nand U4668 (N_4668,N_593,N_486);
xnor U4669 (N_4669,N_321,N_565);
and U4670 (N_4670,N_401,N_2278);
nand U4671 (N_4671,N_2233,N_2042);
nor U4672 (N_4672,N_521,N_35);
nor U4673 (N_4673,N_2089,N_1283);
and U4674 (N_4674,N_717,N_1235);
nor U4675 (N_4675,N_181,N_396);
and U4676 (N_4676,N_1053,N_2088);
xnor U4677 (N_4677,N_94,N_1094);
and U4678 (N_4678,N_908,N_2252);
or U4679 (N_4679,N_787,N_523);
or U4680 (N_4680,N_1811,N_2175);
or U4681 (N_4681,N_1670,N_1017);
xor U4682 (N_4682,N_971,N_1621);
nand U4683 (N_4683,N_208,N_1077);
xor U4684 (N_4684,N_914,N_267);
nor U4685 (N_4685,N_2455,N_1227);
and U4686 (N_4686,N_2199,N_1589);
or U4687 (N_4687,N_796,N_1630);
nand U4688 (N_4688,N_1823,N_710);
nand U4689 (N_4689,N_2126,N_2251);
xnor U4690 (N_4690,N_2433,N_1944);
xnor U4691 (N_4691,N_1676,N_615);
nand U4692 (N_4692,N_75,N_1967);
nand U4693 (N_4693,N_499,N_568);
nand U4694 (N_4694,N_2408,N_1282);
nand U4695 (N_4695,N_58,N_1520);
and U4696 (N_4696,N_1293,N_106);
nand U4697 (N_4697,N_759,N_1678);
or U4698 (N_4698,N_1719,N_442);
and U4699 (N_4699,N_811,N_203);
and U4700 (N_4700,N_1315,N_1742);
or U4701 (N_4701,N_1516,N_2135);
nor U4702 (N_4702,N_664,N_1480);
nand U4703 (N_4703,N_1525,N_1618);
nor U4704 (N_4704,N_1773,N_1183);
or U4705 (N_4705,N_77,N_1270);
nor U4706 (N_4706,N_394,N_1355);
xnor U4707 (N_4707,N_111,N_2074);
nor U4708 (N_4708,N_672,N_228);
or U4709 (N_4709,N_1522,N_1874);
nand U4710 (N_4710,N_360,N_2468);
nand U4711 (N_4711,N_1943,N_1648);
xor U4712 (N_4712,N_30,N_20);
nand U4713 (N_4713,N_1190,N_240);
xnor U4714 (N_4714,N_1145,N_501);
or U4715 (N_4715,N_1620,N_960);
nand U4716 (N_4716,N_46,N_858);
nor U4717 (N_4717,N_2019,N_1807);
nor U4718 (N_4718,N_1111,N_1501);
xor U4719 (N_4719,N_2153,N_648);
xnor U4720 (N_4720,N_153,N_1278);
nor U4721 (N_4721,N_1964,N_1028);
nor U4722 (N_4722,N_1240,N_744);
and U4723 (N_4723,N_216,N_2143);
or U4724 (N_4724,N_2484,N_199);
nand U4725 (N_4725,N_2297,N_1437);
or U4726 (N_4726,N_1783,N_1607);
and U4727 (N_4727,N_356,N_1909);
nand U4728 (N_4728,N_2457,N_16);
or U4729 (N_4729,N_1863,N_854);
xor U4730 (N_4730,N_2121,N_1654);
and U4731 (N_4731,N_18,N_148);
or U4732 (N_4732,N_1131,N_1076);
or U4733 (N_4733,N_1665,N_2045);
or U4734 (N_4734,N_461,N_1347);
xnor U4735 (N_4735,N_973,N_310);
and U4736 (N_4736,N_266,N_2488);
and U4737 (N_4737,N_2157,N_1867);
or U4738 (N_4738,N_1717,N_1668);
or U4739 (N_4739,N_329,N_2219);
and U4740 (N_4740,N_1455,N_1276);
nor U4741 (N_4741,N_65,N_733);
or U4742 (N_4742,N_1073,N_1024);
nand U4743 (N_4743,N_1717,N_1779);
nor U4744 (N_4744,N_1762,N_1142);
or U4745 (N_4745,N_218,N_1236);
nor U4746 (N_4746,N_2086,N_1557);
nand U4747 (N_4747,N_1578,N_1169);
nand U4748 (N_4748,N_2063,N_1843);
nand U4749 (N_4749,N_2239,N_700);
nor U4750 (N_4750,N_2412,N_605);
xnor U4751 (N_4751,N_1229,N_2442);
xnor U4752 (N_4752,N_60,N_669);
xnor U4753 (N_4753,N_1651,N_1262);
or U4754 (N_4754,N_670,N_1231);
nor U4755 (N_4755,N_532,N_1137);
nand U4756 (N_4756,N_916,N_549);
and U4757 (N_4757,N_1244,N_1033);
xor U4758 (N_4758,N_2190,N_1854);
or U4759 (N_4759,N_1720,N_418);
xnor U4760 (N_4760,N_908,N_1922);
nand U4761 (N_4761,N_1577,N_1380);
and U4762 (N_4762,N_422,N_929);
or U4763 (N_4763,N_754,N_869);
nor U4764 (N_4764,N_1956,N_1035);
nor U4765 (N_4765,N_2007,N_2487);
nand U4766 (N_4766,N_934,N_1464);
nor U4767 (N_4767,N_2361,N_1377);
nand U4768 (N_4768,N_1474,N_453);
and U4769 (N_4769,N_2207,N_1860);
or U4770 (N_4770,N_2331,N_1683);
xor U4771 (N_4771,N_38,N_717);
nor U4772 (N_4772,N_625,N_1926);
and U4773 (N_4773,N_2470,N_1736);
or U4774 (N_4774,N_1877,N_1598);
xor U4775 (N_4775,N_1577,N_516);
xnor U4776 (N_4776,N_1117,N_706);
nand U4777 (N_4777,N_578,N_1997);
and U4778 (N_4778,N_600,N_468);
xor U4779 (N_4779,N_291,N_1908);
nor U4780 (N_4780,N_1202,N_1918);
nand U4781 (N_4781,N_267,N_1153);
nand U4782 (N_4782,N_727,N_948);
and U4783 (N_4783,N_516,N_500);
nand U4784 (N_4784,N_1818,N_1904);
nor U4785 (N_4785,N_2163,N_1242);
and U4786 (N_4786,N_806,N_1336);
or U4787 (N_4787,N_886,N_2413);
and U4788 (N_4788,N_1797,N_1616);
nand U4789 (N_4789,N_46,N_2389);
nor U4790 (N_4790,N_1060,N_899);
or U4791 (N_4791,N_1471,N_1289);
and U4792 (N_4792,N_667,N_1725);
nand U4793 (N_4793,N_1232,N_1293);
xnor U4794 (N_4794,N_653,N_1665);
nor U4795 (N_4795,N_915,N_2217);
nor U4796 (N_4796,N_106,N_1266);
nor U4797 (N_4797,N_1187,N_374);
nor U4798 (N_4798,N_146,N_480);
and U4799 (N_4799,N_1427,N_566);
nand U4800 (N_4800,N_2226,N_2403);
or U4801 (N_4801,N_958,N_1254);
and U4802 (N_4802,N_883,N_579);
xnor U4803 (N_4803,N_2320,N_1216);
nor U4804 (N_4804,N_169,N_1328);
or U4805 (N_4805,N_1002,N_166);
and U4806 (N_4806,N_1830,N_2424);
xnor U4807 (N_4807,N_419,N_1127);
xnor U4808 (N_4808,N_1787,N_773);
and U4809 (N_4809,N_1542,N_1626);
and U4810 (N_4810,N_545,N_2433);
nand U4811 (N_4811,N_742,N_1262);
nor U4812 (N_4812,N_1603,N_599);
nand U4813 (N_4813,N_2268,N_1887);
or U4814 (N_4814,N_893,N_1229);
nand U4815 (N_4815,N_1889,N_113);
nand U4816 (N_4816,N_2384,N_291);
and U4817 (N_4817,N_811,N_1200);
xnor U4818 (N_4818,N_1300,N_782);
nand U4819 (N_4819,N_2292,N_1472);
nand U4820 (N_4820,N_373,N_2398);
or U4821 (N_4821,N_1701,N_950);
nor U4822 (N_4822,N_612,N_1699);
or U4823 (N_4823,N_2206,N_1368);
xor U4824 (N_4824,N_2417,N_1917);
nand U4825 (N_4825,N_1333,N_1173);
nand U4826 (N_4826,N_1042,N_1585);
xor U4827 (N_4827,N_344,N_749);
nand U4828 (N_4828,N_1534,N_542);
and U4829 (N_4829,N_1117,N_1682);
xnor U4830 (N_4830,N_1074,N_1320);
or U4831 (N_4831,N_1737,N_957);
nor U4832 (N_4832,N_615,N_2019);
or U4833 (N_4833,N_183,N_2414);
nand U4834 (N_4834,N_454,N_2170);
nand U4835 (N_4835,N_1326,N_1569);
nor U4836 (N_4836,N_22,N_1025);
xor U4837 (N_4837,N_1644,N_1486);
or U4838 (N_4838,N_73,N_2430);
nand U4839 (N_4839,N_1799,N_2066);
nand U4840 (N_4840,N_585,N_1965);
nor U4841 (N_4841,N_2163,N_1298);
nor U4842 (N_4842,N_594,N_819);
nand U4843 (N_4843,N_1146,N_2127);
nand U4844 (N_4844,N_1232,N_158);
xnor U4845 (N_4845,N_1823,N_1112);
and U4846 (N_4846,N_1839,N_2237);
and U4847 (N_4847,N_587,N_736);
nand U4848 (N_4848,N_1225,N_1352);
and U4849 (N_4849,N_185,N_1050);
or U4850 (N_4850,N_832,N_1725);
xnor U4851 (N_4851,N_1351,N_1363);
and U4852 (N_4852,N_249,N_1479);
nor U4853 (N_4853,N_470,N_561);
nor U4854 (N_4854,N_275,N_376);
and U4855 (N_4855,N_563,N_1100);
nand U4856 (N_4856,N_2198,N_1483);
or U4857 (N_4857,N_1315,N_35);
nand U4858 (N_4858,N_1339,N_2096);
and U4859 (N_4859,N_1311,N_521);
nand U4860 (N_4860,N_759,N_1817);
xor U4861 (N_4861,N_933,N_1963);
xnor U4862 (N_4862,N_2348,N_1535);
nor U4863 (N_4863,N_46,N_1310);
or U4864 (N_4864,N_1437,N_377);
nand U4865 (N_4865,N_1773,N_2460);
or U4866 (N_4866,N_1992,N_2016);
or U4867 (N_4867,N_358,N_2252);
or U4868 (N_4868,N_2290,N_1589);
or U4869 (N_4869,N_1606,N_1729);
or U4870 (N_4870,N_888,N_1991);
and U4871 (N_4871,N_777,N_643);
and U4872 (N_4872,N_2446,N_872);
or U4873 (N_4873,N_1524,N_36);
xnor U4874 (N_4874,N_1899,N_309);
and U4875 (N_4875,N_1399,N_506);
xor U4876 (N_4876,N_2210,N_851);
or U4877 (N_4877,N_1923,N_1136);
and U4878 (N_4878,N_181,N_210);
nand U4879 (N_4879,N_1415,N_1316);
xnor U4880 (N_4880,N_1643,N_478);
and U4881 (N_4881,N_435,N_1136);
nand U4882 (N_4882,N_2245,N_2458);
or U4883 (N_4883,N_990,N_325);
and U4884 (N_4884,N_340,N_423);
nand U4885 (N_4885,N_580,N_1470);
and U4886 (N_4886,N_1548,N_1839);
nand U4887 (N_4887,N_377,N_2308);
nor U4888 (N_4888,N_2030,N_1505);
and U4889 (N_4889,N_836,N_768);
nand U4890 (N_4890,N_2472,N_1766);
xor U4891 (N_4891,N_190,N_1003);
nand U4892 (N_4892,N_1426,N_2289);
xnor U4893 (N_4893,N_2246,N_2028);
nor U4894 (N_4894,N_103,N_391);
xor U4895 (N_4895,N_65,N_468);
or U4896 (N_4896,N_1510,N_355);
or U4897 (N_4897,N_1464,N_189);
xor U4898 (N_4898,N_492,N_1614);
xnor U4899 (N_4899,N_700,N_995);
nor U4900 (N_4900,N_810,N_1539);
and U4901 (N_4901,N_253,N_2117);
and U4902 (N_4902,N_1447,N_852);
nor U4903 (N_4903,N_93,N_595);
or U4904 (N_4904,N_1257,N_797);
nor U4905 (N_4905,N_2201,N_1346);
xor U4906 (N_4906,N_77,N_250);
nand U4907 (N_4907,N_1215,N_361);
and U4908 (N_4908,N_1009,N_2404);
nand U4909 (N_4909,N_1381,N_108);
xor U4910 (N_4910,N_283,N_1797);
and U4911 (N_4911,N_954,N_1661);
nand U4912 (N_4912,N_2225,N_2038);
xor U4913 (N_4913,N_1727,N_1012);
and U4914 (N_4914,N_3,N_318);
nor U4915 (N_4915,N_781,N_1430);
or U4916 (N_4916,N_2229,N_1373);
nor U4917 (N_4917,N_865,N_2287);
nand U4918 (N_4918,N_293,N_2408);
nor U4919 (N_4919,N_1819,N_1323);
and U4920 (N_4920,N_2268,N_2323);
nor U4921 (N_4921,N_253,N_411);
xnor U4922 (N_4922,N_1555,N_506);
and U4923 (N_4923,N_989,N_291);
or U4924 (N_4924,N_928,N_2299);
nor U4925 (N_4925,N_1098,N_62);
or U4926 (N_4926,N_1295,N_664);
nand U4927 (N_4927,N_2445,N_2035);
nor U4928 (N_4928,N_1658,N_834);
or U4929 (N_4929,N_1399,N_702);
and U4930 (N_4930,N_2338,N_1693);
and U4931 (N_4931,N_134,N_2027);
nand U4932 (N_4932,N_1982,N_2398);
nand U4933 (N_4933,N_1524,N_1492);
and U4934 (N_4934,N_2188,N_1508);
xor U4935 (N_4935,N_1751,N_1143);
and U4936 (N_4936,N_1581,N_1302);
nor U4937 (N_4937,N_318,N_1161);
nor U4938 (N_4938,N_1276,N_1438);
xnor U4939 (N_4939,N_482,N_15);
nor U4940 (N_4940,N_1229,N_71);
nand U4941 (N_4941,N_1364,N_187);
nand U4942 (N_4942,N_1153,N_914);
and U4943 (N_4943,N_1937,N_1351);
nand U4944 (N_4944,N_2135,N_297);
nor U4945 (N_4945,N_2129,N_506);
and U4946 (N_4946,N_1262,N_1880);
or U4947 (N_4947,N_617,N_1320);
or U4948 (N_4948,N_649,N_1528);
nand U4949 (N_4949,N_985,N_1939);
or U4950 (N_4950,N_2356,N_9);
xor U4951 (N_4951,N_1869,N_64);
nor U4952 (N_4952,N_1181,N_1704);
nor U4953 (N_4953,N_1299,N_2148);
nand U4954 (N_4954,N_1566,N_454);
and U4955 (N_4955,N_267,N_314);
nor U4956 (N_4956,N_1912,N_2279);
nor U4957 (N_4957,N_1101,N_176);
nand U4958 (N_4958,N_1079,N_1340);
or U4959 (N_4959,N_1830,N_2323);
and U4960 (N_4960,N_836,N_2232);
nor U4961 (N_4961,N_2251,N_1967);
xor U4962 (N_4962,N_2041,N_1649);
or U4963 (N_4963,N_801,N_426);
nor U4964 (N_4964,N_284,N_1282);
or U4965 (N_4965,N_2101,N_1679);
nor U4966 (N_4966,N_120,N_173);
nand U4967 (N_4967,N_148,N_183);
nor U4968 (N_4968,N_978,N_397);
and U4969 (N_4969,N_18,N_427);
xor U4970 (N_4970,N_324,N_328);
xor U4971 (N_4971,N_1159,N_721);
nor U4972 (N_4972,N_1052,N_2070);
nor U4973 (N_4973,N_477,N_1191);
and U4974 (N_4974,N_2083,N_113);
or U4975 (N_4975,N_591,N_1819);
and U4976 (N_4976,N_659,N_470);
or U4977 (N_4977,N_2327,N_482);
xnor U4978 (N_4978,N_1802,N_182);
xor U4979 (N_4979,N_712,N_2335);
xnor U4980 (N_4980,N_1452,N_1594);
xnor U4981 (N_4981,N_774,N_2497);
and U4982 (N_4982,N_1941,N_1308);
nor U4983 (N_4983,N_1681,N_944);
or U4984 (N_4984,N_206,N_1407);
xor U4985 (N_4985,N_148,N_1410);
nor U4986 (N_4986,N_2178,N_1263);
and U4987 (N_4987,N_2100,N_923);
or U4988 (N_4988,N_1557,N_2097);
xor U4989 (N_4989,N_2028,N_1076);
xor U4990 (N_4990,N_678,N_1580);
xnor U4991 (N_4991,N_1360,N_1557);
nand U4992 (N_4992,N_2194,N_1382);
and U4993 (N_4993,N_470,N_1950);
xnor U4994 (N_4994,N_339,N_1504);
nor U4995 (N_4995,N_1896,N_619);
or U4996 (N_4996,N_2323,N_949);
nor U4997 (N_4997,N_435,N_1803);
and U4998 (N_4998,N_1090,N_744);
and U4999 (N_4999,N_2138,N_1165);
nand UO_0 (O_0,N_3631,N_3504);
or UO_1 (O_1,N_2778,N_3477);
nand UO_2 (O_2,N_3200,N_3365);
or UO_3 (O_3,N_3749,N_3542);
nor UO_4 (O_4,N_4946,N_4207);
or UO_5 (O_5,N_3202,N_3510);
or UO_6 (O_6,N_4155,N_4781);
nor UO_7 (O_7,N_3397,N_3162);
xor UO_8 (O_8,N_4815,N_4124);
or UO_9 (O_9,N_3611,N_3744);
or UO_10 (O_10,N_3553,N_2563);
xor UO_11 (O_11,N_4600,N_4104);
nor UO_12 (O_12,N_4375,N_2869);
and UO_13 (O_13,N_4950,N_3845);
xor UO_14 (O_14,N_4254,N_4026);
xor UO_15 (O_15,N_3592,N_2855);
nor UO_16 (O_16,N_4090,N_2547);
and UO_17 (O_17,N_4745,N_4788);
nor UO_18 (O_18,N_4511,N_2614);
or UO_19 (O_19,N_4496,N_4741);
nand UO_20 (O_20,N_3757,N_4672);
nor UO_21 (O_21,N_4422,N_3909);
nand UO_22 (O_22,N_3010,N_4116);
and UO_23 (O_23,N_4519,N_4641);
nand UO_24 (O_24,N_4602,N_3745);
nand UO_25 (O_25,N_4711,N_4359);
nand UO_26 (O_26,N_4512,N_4665);
xnor UO_27 (O_27,N_3440,N_3817);
xor UO_28 (O_28,N_3864,N_3225);
nor UO_29 (O_29,N_4379,N_2791);
and UO_30 (O_30,N_3984,N_3349);
nor UO_31 (O_31,N_3613,N_4239);
and UO_32 (O_32,N_2889,N_4916);
and UO_33 (O_33,N_3420,N_4933);
or UO_34 (O_34,N_2839,N_2590);
or UO_35 (O_35,N_4058,N_3532);
and UO_36 (O_36,N_3525,N_2738);
nor UO_37 (O_37,N_4934,N_2900);
nor UO_38 (O_38,N_3302,N_3007);
nor UO_39 (O_39,N_4159,N_2972);
and UO_40 (O_40,N_4014,N_4384);
or UO_41 (O_41,N_3621,N_4660);
xnor UO_42 (O_42,N_3997,N_4889);
xor UO_43 (O_43,N_3518,N_4985);
and UO_44 (O_44,N_3471,N_3392);
nor UO_45 (O_45,N_4478,N_2678);
xor UO_46 (O_46,N_4756,N_4764);
nand UO_47 (O_47,N_3533,N_2545);
or UO_48 (O_48,N_3431,N_4795);
or UO_49 (O_49,N_3782,N_3589);
or UO_50 (O_50,N_4839,N_3561);
and UO_51 (O_51,N_3305,N_3040);
and UO_52 (O_52,N_3145,N_4334);
nor UO_53 (O_53,N_3310,N_3074);
nand UO_54 (O_54,N_3890,N_2562);
nand UO_55 (O_55,N_4280,N_3177);
xor UO_56 (O_56,N_4455,N_3345);
nor UO_57 (O_57,N_4544,N_4004);
nor UO_58 (O_58,N_4825,N_4109);
and UO_59 (O_59,N_4638,N_2540);
xnor UO_60 (O_60,N_4079,N_3758);
or UO_61 (O_61,N_4939,N_2640);
xnor UO_62 (O_62,N_3171,N_4527);
or UO_63 (O_63,N_3926,N_2989);
nor UO_64 (O_64,N_2569,N_4157);
xor UO_65 (O_65,N_3445,N_3617);
or UO_66 (O_66,N_3313,N_4694);
nand UO_67 (O_67,N_2722,N_4800);
or UO_68 (O_68,N_4509,N_2765);
and UO_69 (O_69,N_2861,N_4853);
or UO_70 (O_70,N_3839,N_3157);
or UO_71 (O_71,N_3273,N_3629);
nor UO_72 (O_72,N_2845,N_2946);
and UO_73 (O_73,N_4158,N_3128);
nand UO_74 (O_74,N_3581,N_3969);
and UO_75 (O_75,N_3513,N_4120);
nand UO_76 (O_76,N_3679,N_4217);
and UO_77 (O_77,N_4230,N_3108);
nor UO_78 (O_78,N_2509,N_3131);
or UO_79 (O_79,N_2549,N_4960);
nor UO_80 (O_80,N_2896,N_3276);
xnor UO_81 (O_81,N_4761,N_3156);
xnor UO_82 (O_82,N_4565,N_3165);
nor UO_83 (O_83,N_3537,N_2894);
nand UO_84 (O_84,N_4830,N_4345);
xnor UO_85 (O_85,N_4110,N_3052);
nor UO_86 (O_86,N_2955,N_2682);
and UO_87 (O_87,N_4613,N_3316);
xnor UO_88 (O_88,N_4924,N_3201);
or UO_89 (O_89,N_3355,N_4619);
or UO_90 (O_90,N_3119,N_3776);
or UO_91 (O_91,N_4060,N_4669);
and UO_92 (O_92,N_3761,N_3859);
or UO_93 (O_93,N_2630,N_2566);
xor UO_94 (O_94,N_4382,N_2767);
nor UO_95 (O_95,N_3779,N_4184);
nor UO_96 (O_96,N_4983,N_4418);
and UO_97 (O_97,N_4925,N_2568);
nand UO_98 (O_98,N_4843,N_4123);
nor UO_99 (O_99,N_3669,N_4879);
xor UO_100 (O_100,N_4161,N_3696);
xnor UO_101 (O_101,N_4163,N_4331);
xnor UO_102 (O_102,N_2846,N_4100);
or UO_103 (O_103,N_2988,N_4528);
nor UO_104 (O_104,N_4706,N_4067);
nand UO_105 (O_105,N_4620,N_3852);
nor UO_106 (O_106,N_3759,N_2862);
or UO_107 (O_107,N_3286,N_4918);
xnor UO_108 (O_108,N_2703,N_3650);
xnor UO_109 (O_109,N_4787,N_4425);
xor UO_110 (O_110,N_4449,N_3367);
nor UO_111 (O_111,N_2679,N_4194);
or UO_112 (O_112,N_2577,N_4199);
or UO_113 (O_113,N_3223,N_3773);
xnor UO_114 (O_114,N_4214,N_3495);
or UO_115 (O_115,N_3424,N_3064);
and UO_116 (O_116,N_4347,N_2792);
and UO_117 (O_117,N_4913,N_4657);
nand UO_118 (O_118,N_3688,N_4411);
or UO_119 (O_119,N_4874,N_2949);
xor UO_120 (O_120,N_2572,N_3323);
xnor UO_121 (O_121,N_3232,N_4566);
nand UO_122 (O_122,N_4016,N_4387);
xnor UO_123 (O_123,N_4777,N_3320);
nor UO_124 (O_124,N_4039,N_4580);
and UO_125 (O_125,N_4831,N_4040);
and UO_126 (O_126,N_2574,N_3885);
and UO_127 (O_127,N_3393,N_2607);
xor UO_128 (O_128,N_4868,N_4753);
xor UO_129 (O_129,N_4416,N_4981);
or UO_130 (O_130,N_2895,N_4119);
nand UO_131 (O_131,N_3651,N_4965);
nand UO_132 (O_132,N_4482,N_2939);
xor UO_133 (O_133,N_4439,N_2871);
or UO_134 (O_134,N_4523,N_2523);
nor UO_135 (O_135,N_3003,N_2784);
nor UO_136 (O_136,N_2967,N_3409);
nor UO_137 (O_137,N_4727,N_4614);
xor UO_138 (O_138,N_2875,N_3916);
nand UO_139 (O_139,N_2953,N_2571);
nand UO_140 (O_140,N_3754,N_3529);
xnor UO_141 (O_141,N_3457,N_3325);
nor UO_142 (O_142,N_3490,N_4812);
xnor UO_143 (O_143,N_3251,N_3266);
and UO_144 (O_144,N_4739,N_4047);
and UO_145 (O_145,N_2942,N_4253);
xnor UO_146 (O_146,N_2613,N_2720);
nor UO_147 (O_147,N_3715,N_4007);
or UO_148 (O_148,N_4351,N_4912);
xor UO_149 (O_149,N_2654,N_3073);
nor UO_150 (O_150,N_3790,N_4671);
nor UO_151 (O_151,N_2632,N_3292);
nor UO_152 (O_152,N_3093,N_3667);
and UO_153 (O_153,N_3865,N_3112);
nor UO_154 (O_154,N_4373,N_3208);
or UO_155 (O_155,N_3443,N_3262);
and UO_156 (O_156,N_2616,N_3892);
and UO_157 (O_157,N_3354,N_3427);
xnor UO_158 (O_158,N_3017,N_3267);
nand UO_159 (O_159,N_3066,N_2912);
and UO_160 (O_160,N_2932,N_3469);
nor UO_161 (O_161,N_3479,N_3555);
xor UO_162 (O_162,N_3936,N_4144);
xor UO_163 (O_163,N_3596,N_4869);
and UO_164 (O_164,N_2752,N_3726);
xor UO_165 (O_165,N_4220,N_3192);
and UO_166 (O_166,N_3101,N_3855);
and UO_167 (O_167,N_4259,N_2693);
and UO_168 (O_168,N_3410,N_4229);
nand UO_169 (O_169,N_2876,N_3123);
nor UO_170 (O_170,N_4670,N_4823);
or UO_171 (O_171,N_3205,N_3700);
xnor UO_172 (O_172,N_3212,N_4105);
or UO_173 (O_173,N_3075,N_3341);
nor UO_174 (O_174,N_3465,N_3044);
nor UO_175 (O_175,N_4401,N_4502);
nand UO_176 (O_176,N_3554,N_4832);
xnor UO_177 (O_177,N_4244,N_3482);
xnor UO_178 (O_178,N_2983,N_3359);
or UO_179 (O_179,N_4147,N_4629);
or UO_180 (O_180,N_4061,N_4854);
or UO_181 (O_181,N_4947,N_3820);
nor UO_182 (O_182,N_3933,N_4987);
xnor UO_183 (O_183,N_3185,N_4664);
and UO_184 (O_184,N_2591,N_4516);
and UO_185 (O_185,N_2775,N_4885);
xnor UO_186 (O_186,N_3883,N_2760);
nand UO_187 (O_187,N_4397,N_3786);
or UO_188 (O_188,N_3906,N_4267);
nand UO_189 (O_189,N_4995,N_2564);
nand UO_190 (O_190,N_3861,N_4845);
or UO_191 (O_191,N_4264,N_4555);
nor UO_192 (O_192,N_4696,N_3559);
nor UO_193 (O_193,N_4647,N_3888);
and UO_194 (O_194,N_3268,N_3370);
nand UO_195 (O_195,N_3886,N_2824);
xor UO_196 (O_196,N_3849,N_3265);
and UO_197 (O_197,N_3734,N_3161);
nor UO_198 (O_198,N_4107,N_3092);
and UO_199 (O_199,N_3900,N_3042);
nand UO_200 (O_200,N_3810,N_2906);
and UO_201 (O_201,N_2593,N_4049);
xor UO_202 (O_202,N_4537,N_3377);
and UO_203 (O_203,N_4403,N_3035);
xor UO_204 (O_204,N_4746,N_4166);
or UO_205 (O_205,N_3780,N_3620);
xor UO_206 (O_206,N_4902,N_2516);
xnor UO_207 (O_207,N_3048,N_4059);
or UO_208 (O_208,N_3142,N_4543);
xor UO_209 (O_209,N_4182,N_3148);
nand UO_210 (O_210,N_3024,N_3455);
xnor UO_211 (O_211,N_4782,N_3439);
nor UO_212 (O_212,N_3184,N_2854);
xnor UO_213 (O_213,N_2651,N_4659);
nor UO_214 (O_214,N_4705,N_3701);
nand UO_215 (O_215,N_2905,N_3038);
xor UO_216 (O_216,N_3059,N_2926);
xnor UO_217 (O_217,N_4176,N_3049);
nand UO_218 (O_218,N_4410,N_4558);
and UO_219 (O_219,N_3730,N_2592);
and UO_220 (O_220,N_3364,N_4508);
nand UO_221 (O_221,N_3814,N_2834);
nor UO_222 (O_222,N_4860,N_3330);
or UO_223 (O_223,N_4847,N_4233);
or UO_224 (O_224,N_3638,N_2816);
nand UO_225 (O_225,N_2978,N_2696);
nor UO_226 (O_226,N_4301,N_3512);
or UO_227 (O_227,N_2652,N_3163);
or UO_228 (O_228,N_3248,N_4856);
xor UO_229 (O_229,N_3838,N_3953);
nand UO_230 (O_230,N_4312,N_4051);
xnor UO_231 (O_231,N_2669,N_2511);
or UO_232 (O_232,N_4247,N_3433);
and UO_233 (O_233,N_4595,N_4851);
and UO_234 (O_234,N_4848,N_3105);
or UO_235 (O_235,N_4456,N_3181);
nor UO_236 (O_236,N_2795,N_4738);
xnor UO_237 (O_237,N_4162,N_4855);
nand UO_238 (O_238,N_2878,N_4898);
and UO_239 (O_239,N_4768,N_3087);
and UO_240 (O_240,N_4008,N_2726);
nor UO_241 (O_241,N_3222,N_3078);
nor UO_242 (O_242,N_4434,N_3380);
or UO_243 (O_243,N_4524,N_3139);
nor UO_244 (O_244,N_4616,N_4474);
and UO_245 (O_245,N_2909,N_4391);
nor UO_246 (O_246,N_4042,N_3544);
or UO_247 (O_247,N_3254,N_4836);
or UO_248 (O_248,N_3018,N_2982);
or UO_249 (O_249,N_3685,N_2803);
nor UO_250 (O_250,N_2870,N_3795);
and UO_251 (O_251,N_3277,N_3841);
nand UO_252 (O_252,N_2844,N_3491);
nand UO_253 (O_253,N_3732,N_2504);
and UO_254 (O_254,N_4962,N_4068);
or UO_255 (O_255,N_4043,N_3980);
nor UO_256 (O_256,N_2951,N_4646);
nand UO_257 (O_257,N_3346,N_4295);
nor UO_258 (O_258,N_4466,N_4770);
nor UO_259 (O_259,N_2995,N_4993);
nand UO_260 (O_260,N_3417,N_3981);
nor UO_261 (O_261,N_3653,N_4826);
xor UO_262 (O_262,N_4273,N_3763);
nand UO_263 (O_263,N_3929,N_3407);
nor UO_264 (O_264,N_3778,N_2707);
xor UO_265 (O_265,N_4069,N_4216);
nand UO_266 (O_266,N_3987,N_4296);
nor UO_267 (O_267,N_4095,N_2774);
xnor UO_268 (O_268,N_4692,N_2598);
nand UO_269 (O_269,N_4535,N_3468);
xor UO_270 (O_270,N_4048,N_4631);
nor UO_271 (O_271,N_4611,N_3774);
nand UO_272 (O_272,N_3244,N_3271);
and UO_273 (O_273,N_4488,N_3008);
or UO_274 (O_274,N_2756,N_2819);
or UO_275 (O_275,N_3649,N_2928);
xnor UO_276 (O_276,N_4583,N_2758);
xnor UO_277 (O_277,N_4680,N_3360);
or UO_278 (O_278,N_4571,N_3762);
xor UO_279 (O_279,N_4044,N_3913);
and UO_280 (O_280,N_3467,N_4342);
or UO_281 (O_281,N_3366,N_3236);
nor UO_282 (O_282,N_3643,N_4361);
xor UO_283 (O_283,N_3576,N_4994);
nor UO_284 (O_284,N_3437,N_2639);
xnor UO_285 (O_285,N_4444,N_4693);
nand UO_286 (O_286,N_2897,N_3279);
xor UO_287 (O_287,N_3704,N_4115);
nor UO_288 (O_288,N_2914,N_3577);
xor UO_289 (O_289,N_4718,N_3497);
or UO_290 (O_290,N_4023,N_2829);
or UO_291 (O_291,N_3384,N_3923);
and UO_292 (O_292,N_2808,N_2918);
nor UO_293 (O_293,N_3056,N_4529);
and UO_294 (O_294,N_4172,N_3388);
nand UO_295 (O_295,N_3610,N_4075);
or UO_296 (O_296,N_4017,N_4982);
xnor UO_297 (O_297,N_4292,N_4374);
nor UO_298 (O_298,N_4594,N_4307);
nor UO_299 (O_299,N_3950,N_3245);
or UO_300 (O_300,N_3198,N_4167);
nor UO_301 (O_301,N_3293,N_4000);
nor UO_302 (O_302,N_3028,N_3032);
or UO_303 (O_303,N_3151,N_2699);
or UO_304 (O_304,N_2576,N_2815);
or UO_305 (O_305,N_2780,N_3784);
xor UO_306 (O_306,N_4970,N_4691);
nand UO_307 (O_307,N_3047,N_3684);
or UO_308 (O_308,N_4302,N_4193);
nor UO_309 (O_309,N_4056,N_3961);
nor UO_310 (O_310,N_4773,N_4737);
and UO_311 (O_311,N_2762,N_3719);
nand UO_312 (O_312,N_3317,N_2748);
nand UO_313 (O_313,N_4779,N_3282);
or UO_314 (O_314,N_3141,N_2961);
nand UO_315 (O_315,N_2923,N_4177);
or UO_316 (O_316,N_4575,N_4389);
nor UO_317 (O_317,N_4236,N_3760);
and UO_318 (O_318,N_2727,N_2683);
xnor UO_319 (O_319,N_2821,N_2958);
xor UO_320 (O_320,N_4656,N_4796);
or UO_321 (O_321,N_2580,N_3582);
or UO_322 (O_322,N_4112,N_4228);
xnor UO_323 (O_323,N_3705,N_3521);
nand UO_324 (O_324,N_2793,N_3012);
xor UO_325 (O_325,N_4590,N_3673);
nor UO_326 (O_326,N_2565,N_3314);
or UO_327 (O_327,N_4714,N_4130);
nand UO_328 (O_328,N_4897,N_4562);
nand UO_329 (O_329,N_4792,N_3270);
and UO_330 (O_330,N_3858,N_2954);
nor UO_331 (O_331,N_4398,N_4400);
or UO_332 (O_332,N_4462,N_2887);
xor UO_333 (O_333,N_4033,N_3030);
nor UO_334 (O_334,N_3086,N_4131);
nand UO_335 (O_335,N_3182,N_2920);
nor UO_336 (O_336,N_3363,N_4695);
nor UO_337 (O_337,N_2915,N_4336);
nand UO_338 (O_338,N_3333,N_3910);
or UO_339 (O_339,N_2930,N_4499);
or UO_340 (O_340,N_4451,N_3095);
nor UO_341 (O_341,N_4034,N_4877);
nor UO_342 (O_342,N_2681,N_4117);
or UO_343 (O_343,N_4678,N_4365);
nand UO_344 (O_344,N_4188,N_3189);
or UO_345 (O_345,N_3639,N_4353);
nand UO_346 (O_346,N_3138,N_3516);
xor UO_347 (O_347,N_4639,N_2763);
nand UO_348 (O_348,N_3219,N_4968);
nor UO_349 (O_349,N_2736,N_4633);
nor UO_350 (O_350,N_2850,N_2624);
nand UO_351 (O_351,N_4245,N_3637);
and UO_352 (O_352,N_4204,N_4838);
and UO_353 (O_353,N_4406,N_3503);
nand UO_354 (O_354,N_4308,N_3456);
and UO_355 (O_355,N_4383,N_4252);
or UO_356 (O_356,N_4518,N_3091);
and UO_357 (O_357,N_4708,N_4884);
xor UO_358 (O_358,N_3659,N_3432);
nor UO_359 (O_359,N_4473,N_2575);
or UO_360 (O_360,N_3935,N_2706);
nor UO_361 (O_361,N_3051,N_2987);
and UO_362 (O_362,N_4431,N_2676);
or UO_363 (O_363,N_4121,N_4173);
or UO_364 (O_364,N_4498,N_3813);
nand UO_365 (O_365,N_2541,N_3338);
xor UO_366 (O_366,N_3526,N_4900);
xnor UO_367 (O_367,N_2770,N_3698);
and UO_368 (O_368,N_4895,N_3847);
nor UO_369 (O_369,N_3966,N_4942);
and UO_370 (O_370,N_4078,N_4208);
nor UO_371 (O_371,N_4806,N_4728);
and UO_372 (O_372,N_4494,N_3728);
and UO_373 (O_373,N_2754,N_3930);
xor UO_374 (O_374,N_3475,N_2560);
xor UO_375 (O_375,N_4592,N_3309);
xnor UO_376 (O_376,N_3523,N_3041);
and UO_377 (O_377,N_3939,N_2619);
nand UO_378 (O_378,N_2656,N_4074);
and UO_379 (O_379,N_2522,N_2952);
nand UO_380 (O_380,N_2874,N_2691);
nor UO_381 (O_381,N_4755,N_4186);
xor UO_382 (O_382,N_3692,N_2513);
nor UO_383 (O_383,N_3037,N_3382);
or UO_384 (O_384,N_3569,N_2814);
nor UO_385 (O_385,N_3036,N_3164);
nand UO_386 (O_386,N_4209,N_3110);
and UO_387 (O_387,N_4998,N_4165);
xor UO_388 (O_388,N_4329,N_4700);
xor UO_389 (O_389,N_4844,N_2963);
xor UO_390 (O_390,N_4608,N_4350);
xor UO_391 (O_391,N_4080,N_4828);
nand UO_392 (O_392,N_3870,N_4701);
xnor UO_393 (O_393,N_4872,N_4568);
and UO_394 (O_394,N_3718,N_2742);
xnor UO_395 (O_395,N_2636,N_4407);
xor UO_396 (O_396,N_4019,N_4687);
nand UO_397 (O_397,N_4809,N_4937);
nor UO_398 (O_398,N_3050,N_3767);
nor UO_399 (O_399,N_3585,N_3663);
or UO_400 (O_400,N_3501,N_4959);
and UO_401 (O_401,N_2859,N_3570);
or UO_402 (O_402,N_3080,N_3675);
nor UO_403 (O_403,N_3283,N_2519);
nand UO_404 (O_404,N_3985,N_3451);
nand UO_405 (O_405,N_3090,N_4721);
nor UO_406 (O_406,N_4865,N_3702);
xor UO_407 (O_407,N_4362,N_2537);
xor UO_408 (O_408,N_3738,N_4598);
nand UO_409 (O_409,N_3107,N_4196);
and UO_410 (O_410,N_2867,N_2730);
nor UO_411 (O_411,N_4125,N_3741);
xnor UO_412 (O_412,N_3344,N_4928);
nand UO_413 (O_413,N_2660,N_3275);
xnor UO_414 (O_414,N_4772,N_4927);
xnor UO_415 (O_415,N_3598,N_2788);
or UO_416 (O_416,N_3307,N_4634);
and UO_417 (O_417,N_3129,N_4153);
nand UO_418 (O_418,N_2718,N_2991);
nand UO_419 (O_419,N_4585,N_3480);
or UO_420 (O_420,N_4977,N_2857);
nand UO_421 (O_421,N_4742,N_4294);
or UO_422 (O_422,N_3288,N_3628);
or UO_423 (O_423,N_3511,N_4064);
and UO_424 (O_424,N_3579,N_4459);
nor UO_425 (O_425,N_3717,N_2898);
and UO_426 (O_426,N_3699,N_3952);
xor UO_427 (O_427,N_2655,N_3614);
nand UO_428 (O_428,N_3258,N_2888);
and UO_429 (O_429,N_4197,N_3894);
and UO_430 (O_430,N_2934,N_3113);
nor UO_431 (O_431,N_3874,N_4178);
xor UO_432 (O_432,N_3188,N_4992);
nand UO_433 (O_433,N_4118,N_2578);
nor UO_434 (O_434,N_4191,N_4997);
xnor UO_435 (O_435,N_3104,N_4624);
and UO_436 (O_436,N_2744,N_3083);
xnor UO_437 (O_437,N_3735,N_4533);
xor UO_438 (O_438,N_4752,N_4584);
and UO_439 (O_439,N_4921,N_4525);
nand UO_440 (O_440,N_3771,N_4547);
or UO_441 (O_441,N_3046,N_2594);
nand UO_442 (O_442,N_3860,N_2713);
nor UO_443 (O_443,N_4644,N_3941);
and UO_444 (O_444,N_3600,N_4143);
or UO_445 (O_445,N_3043,N_2526);
and UO_446 (O_446,N_2747,N_3571);
and UO_447 (O_447,N_4378,N_4287);
nor UO_448 (O_448,N_3796,N_3789);
nand UO_449 (O_449,N_3062,N_4999);
xnor UO_450 (O_450,N_4160,N_2557);
and UO_451 (O_451,N_3487,N_3565);
xnor UO_452 (O_452,N_2600,N_3963);
nand UO_453 (O_453,N_3291,N_4472);
nand UO_454 (O_454,N_4419,N_4880);
and UO_455 (O_455,N_4402,N_3206);
nor UO_456 (O_456,N_4053,N_3326);
or UO_457 (O_457,N_4135,N_4785);
nor UO_458 (O_458,N_3593,N_3117);
or UO_459 (O_459,N_3353,N_3548);
nor UO_460 (O_460,N_3458,N_3100);
nand UO_461 (O_461,N_4736,N_3396);
nand UO_462 (O_462,N_3125,N_2570);
and UO_463 (O_463,N_3528,N_2956);
or UO_464 (O_464,N_2985,N_3564);
xnor UO_465 (O_465,N_4716,N_3398);
nor UO_466 (O_466,N_3452,N_4145);
and UO_467 (O_467,N_4842,N_3295);
nand UO_468 (O_468,N_4149,N_3633);
xnor UO_469 (O_469,N_4395,N_2827);
and UO_470 (O_470,N_4357,N_3211);
nor UO_471 (O_471,N_3674,N_4251);
and UO_472 (O_472,N_4975,N_3081);
or UO_473 (O_473,N_3829,N_4174);
or UO_474 (O_474,N_4763,N_3531);
nor UO_475 (O_475,N_2551,N_4990);
xor UO_476 (O_476,N_4945,N_4559);
and UO_477 (O_477,N_3568,N_3146);
or UO_478 (O_478,N_4683,N_2615);
or UO_479 (O_479,N_2702,N_4485);
nor UO_480 (O_480,N_3534,N_4704);
or UO_481 (O_481,N_3278,N_4372);
or UO_482 (O_482,N_4979,N_2929);
and UO_483 (O_483,N_3634,N_3856);
nor UO_484 (O_484,N_3460,N_4917);
and UO_485 (O_485,N_4908,N_4187);
or UO_486 (O_486,N_4089,N_4765);
nor UO_487 (O_487,N_4050,N_2647);
and UO_488 (O_488,N_4440,N_3103);
or UO_489 (O_489,N_3988,N_4581);
nand UO_490 (O_490,N_3230,N_4675);
and UO_491 (O_491,N_4886,N_3216);
nand UO_492 (O_492,N_3195,N_4817);
and UO_493 (O_493,N_4972,N_2515);
xor UO_494 (O_494,N_4349,N_4579);
xnor UO_495 (O_495,N_4666,N_4238);
or UO_496 (O_496,N_3102,N_3376);
nor UO_497 (O_497,N_4423,N_3588);
or UO_498 (O_498,N_3804,N_4510);
or UO_499 (O_499,N_3716,N_2950);
or UO_500 (O_500,N_4293,N_2627);
xnor UO_501 (O_501,N_4005,N_3901);
xor UO_502 (O_502,N_3661,N_3586);
nand UO_503 (O_503,N_4096,N_3013);
xor UO_504 (O_504,N_3851,N_2661);
nand UO_505 (O_505,N_2740,N_2503);
xor UO_506 (O_506,N_4190,N_3290);
xnor UO_507 (O_507,N_3805,N_2853);
nand UO_508 (O_508,N_2620,N_3943);
nand UO_509 (O_509,N_3005,N_4128);
or UO_510 (O_510,N_3955,N_4663);
and UO_511 (O_511,N_3312,N_4006);
nor UO_512 (O_512,N_4774,N_2879);
nor UO_513 (O_513,N_3068,N_3058);
nand UO_514 (O_514,N_3287,N_3977);
xor UO_515 (O_515,N_3927,N_3689);
nor UO_516 (O_516,N_3925,N_3783);
or UO_517 (O_517,N_2831,N_3133);
or UO_518 (O_518,N_3387,N_3945);
nor UO_519 (O_519,N_4366,N_4576);
xnor UO_520 (O_520,N_4679,N_4285);
and UO_521 (O_521,N_3562,N_3336);
nor UO_522 (O_522,N_4952,N_3976);
nand UO_523 (O_523,N_3992,N_4227);
nor UO_524 (O_524,N_4279,N_4170);
or UO_525 (O_525,N_3990,N_3399);
xnor UO_526 (O_526,N_3079,N_3808);
or UO_527 (O_527,N_2688,N_4150);
xor UO_528 (O_528,N_4915,N_3350);
xor UO_529 (O_529,N_4747,N_3239);
nand UO_530 (O_530,N_2662,N_3413);
nor UO_531 (O_531,N_2719,N_3084);
and UO_532 (O_532,N_4956,N_4325);
nor UO_533 (O_533,N_4320,N_2510);
xnor UO_534 (O_534,N_4321,N_4348);
and UO_535 (O_535,N_4991,N_3536);
nor UO_536 (O_536,N_2637,N_2892);
xnor UO_537 (O_537,N_4778,N_4435);
and UO_538 (O_538,N_3257,N_3606);
and UO_539 (O_539,N_3907,N_2561);
and UO_540 (O_540,N_2924,N_4541);
xnor UO_541 (O_541,N_4030,N_3962);
nor UO_542 (O_542,N_4305,N_2643);
and UO_543 (O_543,N_3551,N_2717);
nand UO_544 (O_544,N_3476,N_3098);
or UO_545 (O_545,N_3021,N_4324);
nor UO_546 (O_546,N_4386,N_3459);
nand UO_547 (O_547,N_3053,N_2768);
and UO_548 (O_548,N_3390,N_3803);
nor UO_549 (O_549,N_2979,N_3252);
nand UO_550 (O_550,N_3970,N_3115);
or UO_551 (O_551,N_3766,N_4552);
nand UO_552 (O_552,N_3727,N_4803);
xnor UO_553 (O_553,N_4673,N_2646);
nand UO_554 (O_554,N_2579,N_2936);
and UO_555 (O_555,N_3772,N_3289);
nor UO_556 (O_556,N_3957,N_4205);
nor UO_557 (O_557,N_2944,N_3449);
nand UO_558 (O_558,N_4635,N_3204);
and UO_559 (O_559,N_4938,N_3944);
xnor UO_560 (O_560,N_2552,N_3830);
nand UO_561 (O_561,N_3777,N_3264);
and UO_562 (O_562,N_4139,N_2984);
nand UO_563 (O_563,N_2933,N_3483);
or UO_564 (O_564,N_3329,N_2585);
and UO_565 (O_565,N_3878,N_3558);
nand UO_566 (O_566,N_3722,N_4278);
or UO_567 (O_567,N_2860,N_2783);
nor UO_568 (O_568,N_4376,N_4122);
nand UO_569 (O_569,N_2843,N_3824);
nor UO_570 (O_570,N_3821,N_4248);
or UO_571 (O_571,N_4437,N_3130);
or UO_572 (O_572,N_2710,N_2750);
nor UO_573 (O_573,N_4550,N_3463);
nand UO_574 (O_574,N_4224,N_2799);
and UO_575 (O_575,N_4487,N_3706);
nor UO_576 (O_576,N_4086,N_2622);
nand UO_577 (O_577,N_2882,N_3321);
or UO_578 (O_578,N_4491,N_4920);
or UO_579 (O_579,N_4867,N_4572);
and UO_580 (O_580,N_3429,N_2809);
and UO_581 (O_581,N_3247,N_3524);
nand UO_582 (O_582,N_4520,N_2612);
nand UO_583 (O_583,N_2500,N_2721);
nand UO_584 (O_584,N_3602,N_3284);
xnor UO_585 (O_585,N_3756,N_4304);
nand UO_586 (O_586,N_3368,N_3747);
or UO_587 (O_587,N_4313,N_4189);
nor UO_588 (O_588,N_4690,N_2938);
nand UO_589 (O_589,N_3389,N_3775);
or UO_590 (O_590,N_4556,N_2761);
nor UO_591 (O_591,N_4232,N_4046);
nand UO_592 (O_592,N_3448,N_3624);
and UO_593 (O_593,N_3601,N_4370);
nand UO_594 (O_594,N_2800,N_4141);
or UO_595 (O_595,N_4226,N_4582);
nand UO_596 (O_596,N_3351,N_4911);
nor UO_597 (O_597,N_3792,N_2734);
nor UO_598 (O_598,N_4003,N_2908);
and UO_599 (O_599,N_3902,N_4546);
nand UO_600 (O_600,N_4893,N_4949);
and UO_601 (O_601,N_4850,N_3802);
xor UO_602 (O_602,N_4899,N_3519);
nor UO_603 (O_603,N_3430,N_3891);
and UO_604 (O_604,N_3135,N_4943);
and UO_605 (O_605,N_2807,N_3335);
nor UO_606 (O_606,N_3263,N_3823);
nor UO_607 (O_607,N_3681,N_3520);
and UO_608 (O_608,N_3332,N_4859);
or UO_609 (O_609,N_2794,N_4964);
xnor UO_610 (O_610,N_2698,N_4642);
nand UO_611 (O_611,N_4218,N_3899);
xor UO_612 (O_612,N_4493,N_4775);
and UO_613 (O_613,N_4532,N_4901);
nand UO_614 (O_614,N_4989,N_2597);
nor UO_615 (O_615,N_2847,N_3442);
and UO_616 (O_616,N_2863,N_4814);
nor UO_617 (O_617,N_3725,N_2735);
nor UO_618 (O_618,N_4385,N_2825);
and UO_619 (O_619,N_4861,N_4032);
xnor UO_620 (O_620,N_4766,N_2877);
and UO_621 (O_621,N_2917,N_2595);
nand UO_622 (O_622,N_4504,N_4225);
nand UO_623 (O_623,N_2602,N_2971);
and UO_624 (O_624,N_2517,N_4271);
xor UO_625 (O_625,N_2534,N_4589);
and UO_626 (O_626,N_4681,N_3308);
xor UO_627 (O_627,N_2535,N_2611);
nor UO_628 (O_628,N_2692,N_3299);
or UO_629 (O_629,N_4587,N_4726);
and UO_630 (O_630,N_3746,N_4286);
xnor UO_631 (O_631,N_2623,N_2964);
nor UO_632 (O_632,N_4717,N_3022);
xor UO_633 (O_633,N_2671,N_2608);
xnor UO_634 (O_634,N_4783,N_3441);
nand UO_635 (O_635,N_2618,N_3379);
nand UO_636 (O_636,N_3546,N_4769);
and UO_637 (O_637,N_4667,N_3025);
nand UO_638 (O_638,N_3583,N_2626);
xnor UO_639 (O_639,N_3539,N_2508);
nor UO_640 (O_640,N_4066,N_4045);
xor UO_641 (O_641,N_3881,N_4984);
and UO_642 (O_642,N_3983,N_3998);
or UO_643 (O_643,N_4168,N_2542);
nor UO_644 (O_644,N_4599,N_2810);
nand UO_645 (O_645,N_3339,N_4303);
xor UO_646 (O_646,N_4246,N_2728);
or UO_647 (O_647,N_4490,N_4284);
and UO_648 (O_648,N_4270,N_3322);
nand UO_649 (O_649,N_3800,N_3474);
and UO_650 (O_650,N_2948,N_3502);
xor UO_651 (O_651,N_4536,N_2697);
nand UO_652 (O_652,N_4909,N_3951);
or UO_653 (O_653,N_3682,N_3166);
nand UO_654 (O_654,N_4725,N_4076);
and UO_655 (O_655,N_3872,N_3507);
xnor UO_656 (O_656,N_3218,N_3069);
or UO_657 (O_657,N_3383,N_2514);
nor UO_658 (O_658,N_4643,N_4181);
nor UO_659 (O_659,N_3224,N_4863);
nor UO_660 (O_660,N_4688,N_3281);
or UO_661 (O_661,N_4759,N_2842);
or UO_662 (O_662,N_4805,N_3938);
or UO_663 (O_663,N_4054,N_4241);
nor UO_664 (O_664,N_4967,N_4790);
or UO_665 (O_665,N_4930,N_3540);
and UO_666 (O_666,N_4243,N_4650);
or UO_667 (O_667,N_2650,N_4601);
nor UO_668 (O_668,N_4495,N_3527);
nand UO_669 (O_669,N_3004,N_3118);
and UO_670 (O_670,N_3485,N_3221);
or UO_671 (O_671,N_4791,N_3626);
xnor UO_672 (O_672,N_2866,N_3556);
nor UO_673 (O_673,N_2667,N_3347);
nor UO_674 (O_674,N_4206,N_3168);
nor UO_675 (O_675,N_2817,N_4771);
nand UO_676 (O_676,N_2823,N_4035);
and UO_677 (O_677,N_4588,N_3837);
nand UO_678 (O_678,N_2665,N_3009);
and UO_679 (O_679,N_4896,N_4219);
nand UO_680 (O_680,N_3712,N_3693);
nand UO_681 (O_681,N_2672,N_2505);
xor UO_682 (O_682,N_2638,N_2668);
or UO_683 (O_683,N_2725,N_2919);
nor UO_684 (O_684,N_3137,N_4538);
nor UO_685 (O_685,N_2789,N_3866);
or UO_686 (O_686,N_4468,N_2777);
nor UO_687 (O_687,N_3751,N_4890);
xnor UO_688 (O_688,N_4744,N_4171);
and UO_689 (O_689,N_3150,N_3109);
xnor UO_690 (O_690,N_3831,N_3478);
nand UO_691 (O_691,N_3572,N_3713);
or UO_692 (O_692,N_3220,N_3635);
and UO_693 (O_693,N_2559,N_3755);
nor UO_694 (O_694,N_3438,N_3509);
and UO_695 (O_695,N_4323,N_2543);
nor UO_696 (O_696,N_2913,N_3421);
nand UO_697 (O_697,N_4957,N_4904);
xor UO_698 (O_698,N_4651,N_4903);
or UO_699 (O_699,N_3575,N_3996);
or UO_700 (O_700,N_2586,N_3731);
nor UO_701 (O_701,N_3948,N_4729);
xor UO_702 (O_702,N_3508,N_4098);
nor UO_703 (O_703,N_4180,N_4954);
nand UO_704 (O_704,N_4421,N_4625);
xnor UO_705 (O_705,N_4358,N_2582);
or UO_706 (O_706,N_4084,N_4971);
xnor UO_707 (O_707,N_4480,N_3415);
nor UO_708 (O_708,N_4469,N_3517);
or UO_709 (O_709,N_4503,N_3723);
xnor UO_710 (O_710,N_4626,N_2525);
nor UO_711 (O_711,N_3599,N_3172);
or UO_712 (O_712,N_2910,N_3160);
nand UO_713 (O_713,N_4570,N_4940);
nand UO_714 (O_714,N_4427,N_3304);
or UO_715 (O_715,N_3190,N_3099);
nand UO_716 (O_716,N_3375,N_3147);
and UO_717 (O_717,N_4776,N_2996);
and UO_718 (O_718,N_2959,N_3630);
xnor UO_719 (O_719,N_4354,N_3045);
nand UO_720 (O_720,N_2532,N_3654);
and UO_721 (O_721,N_3954,N_4591);
nand UO_722 (O_722,N_4677,N_4299);
or UO_723 (O_723,N_4563,N_4309);
nand UO_724 (O_724,N_4327,N_4364);
nand UO_725 (O_725,N_3801,N_4606);
xnor UO_726 (O_726,N_4133,N_4326);
or UO_727 (O_727,N_3187,N_4460);
nand UO_728 (O_728,N_4029,N_2970);
xor UO_729 (O_729,N_4257,N_4192);
or UO_730 (O_730,N_4328,N_4392);
xnor UO_731 (O_731,N_3797,N_2684);
xnor UO_732 (O_732,N_3836,N_2739);
nor UO_733 (O_733,N_2981,N_4338);
nor UO_734 (O_734,N_3743,N_3085);
xnor UO_735 (O_735,N_2653,N_4399);
or UO_736 (O_736,N_4072,N_4077);
nor UO_737 (O_737,N_3337,N_3835);
nand UO_738 (O_738,N_3547,N_3868);
xor UO_739 (O_739,N_4530,N_3550);
or UO_740 (O_740,N_4255,N_2645);
nand UO_741 (O_741,N_2796,N_4010);
nand UO_742 (O_742,N_4028,N_2957);
xnor UO_743 (O_743,N_3714,N_3067);
and UO_744 (O_744,N_4065,N_3584);
or UO_745 (O_745,N_4501,N_4250);
or UO_746 (O_746,N_3958,N_2715);
and UO_747 (O_747,N_4734,N_4484);
or UO_748 (O_748,N_2872,N_3411);
and UO_749 (O_749,N_3348,N_3416);
or UO_750 (O_750,N_3956,N_4409);
nand UO_751 (O_751,N_3395,N_3303);
xnor UO_752 (O_752,N_4702,N_3893);
nor UO_753 (O_753,N_2556,N_3842);
or UO_754 (O_754,N_2776,N_3750);
or UO_755 (O_755,N_3357,N_4447);
and UO_756 (O_756,N_3111,N_3186);
and UO_757 (O_757,N_3356,N_3652);
xnor UO_758 (O_758,N_4211,N_3174);
xor UO_759 (O_759,N_4833,N_4164);
xnor UO_760 (O_760,N_2704,N_4623);
nand UO_761 (O_761,N_3243,N_2528);
and UO_762 (O_762,N_2904,N_2674);
nor UO_763 (O_763,N_4106,N_4102);
or UO_764 (O_764,N_4822,N_4492);
xnor UO_765 (O_765,N_2960,N_4829);
nor UO_766 (O_766,N_3234,N_3676);
and UO_767 (O_767,N_3680,N_4071);
xnor UO_768 (O_768,N_3001,N_3406);
and UO_769 (O_769,N_4804,N_3076);
nand UO_770 (O_770,N_2772,N_4808);
nand UO_771 (O_771,N_4258,N_2901);
xor UO_772 (O_772,N_4834,N_3788);
and UO_773 (O_773,N_3736,N_3240);
xnor UO_774 (O_774,N_4363,N_4475);
xor UO_775 (O_775,N_4955,N_3965);
nor UO_776 (O_776,N_4322,N_3371);
or UO_777 (O_777,N_3319,N_3054);
nor UO_778 (O_778,N_3724,N_2771);
xor UO_779 (O_779,N_4784,N_3710);
xor UO_780 (O_780,N_3422,N_4081);
xor UO_781 (O_781,N_2790,N_2687);
nand UO_782 (O_782,N_2538,N_3496);
xor UO_783 (O_783,N_4415,N_4497);
xnor UO_784 (O_784,N_4958,N_4703);
and UO_785 (O_785,N_2634,N_4760);
nor UO_786 (O_786,N_4603,N_2805);
or UO_787 (O_787,N_4798,N_2773);
nand UO_788 (O_788,N_4148,N_4291);
or UO_789 (O_789,N_2838,N_4082);
nor UO_790 (O_790,N_2599,N_4750);
nand UO_791 (O_791,N_3595,N_3453);
nand UO_792 (O_792,N_4215,N_3863);
nor UO_793 (O_793,N_4676,N_2798);
nor UO_794 (O_794,N_3563,N_3124);
nand UO_795 (O_795,N_4393,N_3769);
nand UO_796 (O_796,N_4658,N_4027);
nand UO_797 (O_797,N_3057,N_3615);
or UO_798 (O_798,N_4266,N_4269);
or UO_799 (O_799,N_4515,N_2975);
xor UO_800 (O_800,N_2947,N_4441);
and UO_801 (O_801,N_3975,N_4111);
or UO_802 (O_802,N_4201,N_3765);
nor UO_803 (O_803,N_4615,N_4022);
nor UO_804 (O_804,N_3522,N_2746);
or UO_805 (O_805,N_3253,N_3231);
nand UO_806 (O_806,N_3408,N_2781);
xnor UO_807 (O_807,N_3489,N_2976);
or UO_808 (O_808,N_3656,N_4212);
or UO_809 (O_809,N_3720,N_3306);
and UO_810 (O_810,N_4610,N_4797);
nor UO_811 (O_811,N_3272,N_4355);
nand UO_812 (O_812,N_3227,N_4824);
or UO_813 (O_813,N_4470,N_4263);
and UO_814 (O_814,N_4926,N_3619);
nor UO_815 (O_815,N_2993,N_3121);
or UO_816 (O_816,N_4513,N_2851);
nor UO_817 (O_817,N_3904,N_3493);
xnor UO_818 (O_818,N_4404,N_3296);
nand UO_819 (O_819,N_4986,N_3000);
nor UO_820 (O_820,N_2840,N_3481);
or UO_821 (O_821,N_3246,N_3840);
nand UO_822 (O_822,N_4662,N_3662);
or UO_823 (O_823,N_2832,N_3915);
xor UO_824 (O_824,N_3173,N_2530);
or UO_825 (O_825,N_3027,N_2512);
and UO_826 (O_826,N_3671,N_4369);
xnor UO_827 (O_827,N_3655,N_3587);
xor UO_828 (O_828,N_2724,N_4754);
nand UO_829 (O_829,N_3158,N_2980);
xor UO_830 (O_830,N_2852,N_4200);
and UO_831 (O_831,N_3632,N_4640);
or UO_832 (O_832,N_4862,N_4316);
nor UO_833 (O_833,N_2621,N_4919);
nand UO_834 (O_834,N_3014,N_2786);
or UO_835 (O_835,N_4655,N_3557);
nand UO_836 (O_836,N_4567,N_3120);
nand UO_837 (O_837,N_2937,N_3412);
nand UO_838 (O_838,N_3447,N_2965);
and UO_839 (O_839,N_4261,N_3179);
nand UO_840 (O_840,N_3226,N_3402);
xor UO_841 (O_841,N_2890,N_3334);
xor UO_842 (O_842,N_2990,N_4554);
nor UO_843 (O_843,N_4539,N_2677);
and UO_844 (O_844,N_3989,N_3097);
nor UO_845 (O_845,N_4151,N_4612);
and UO_846 (O_846,N_4963,N_4094);
and UO_847 (O_847,N_2558,N_3645);
and UO_848 (O_848,N_2864,N_4894);
or UO_849 (O_849,N_3931,N_3183);
and UO_850 (O_850,N_4932,N_4866);
or UO_851 (O_851,N_3143,N_4132);
nor UO_852 (O_852,N_3644,N_2675);
and UO_853 (O_853,N_3853,N_3854);
nor UO_854 (O_854,N_2893,N_2977);
nand UO_855 (O_855,N_4811,N_4974);
nand UO_856 (O_856,N_3401,N_3903);
xor UO_857 (O_857,N_4929,N_4636);
nor UO_858 (O_858,N_3405,N_4240);
nand UO_859 (O_859,N_3155,N_4413);
nand UO_860 (O_860,N_2664,N_4340);
xor UO_861 (O_861,N_2533,N_4561);
nand UO_862 (O_862,N_3378,N_3709);
xnor UO_863 (O_863,N_3515,N_2880);
or UO_864 (O_864,N_4871,N_4767);
or UO_865 (O_865,N_2858,N_2689);
or UO_866 (O_866,N_3922,N_2741);
or UO_867 (O_867,N_2779,N_4426);
nor UO_868 (O_868,N_4183,N_4277);
xor UO_869 (O_869,N_2709,N_2610);
and UO_870 (O_870,N_3324,N_3917);
nand UO_871 (O_871,N_4973,N_2714);
and UO_872 (O_872,N_4265,N_4380);
nand UO_873 (O_873,N_2935,N_3454);
nand UO_874 (O_874,N_2658,N_4617);
nand UO_875 (O_875,N_3506,N_2733);
or UO_876 (O_876,N_3622,N_4113);
nor UO_877 (O_877,N_3082,N_3089);
or UO_878 (O_878,N_4654,N_3949);
xnor UO_879 (O_879,N_4564,N_4849);
or UO_880 (O_880,N_4887,N_3816);
xor UO_881 (O_881,N_2899,N_3995);
xor UO_882 (O_882,N_3250,N_4710);
and UO_883 (O_883,N_3486,N_3391);
and UO_884 (O_884,N_3664,N_4134);
or UO_885 (O_885,N_3180,N_3294);
or UO_886 (O_886,N_3711,N_3444);
xnor UO_887 (O_887,N_3065,N_2567);
nor UO_888 (O_888,N_3167,N_4574);
nor UO_889 (O_889,N_3686,N_3979);
xor UO_890 (O_890,N_3233,N_4505);
nand UO_891 (O_891,N_4948,N_3386);
and UO_892 (O_892,N_2749,N_3857);
and UO_893 (O_893,N_3260,N_3898);
and UO_894 (O_894,N_2769,N_3876);
xor UO_895 (O_895,N_4483,N_4931);
xor UO_896 (O_896,N_3530,N_3149);
nor UO_897 (O_897,N_2631,N_2745);
or UO_898 (O_898,N_3538,N_4709);
or UO_899 (O_899,N_4540,N_2764);
nand UO_900 (O_900,N_4458,N_4758);
or UO_901 (O_901,N_4698,N_3213);
xnor UO_902 (O_902,N_4888,N_4339);
nand UO_903 (O_903,N_2865,N_3196);
xor UO_904 (O_904,N_3946,N_4794);
nor UO_905 (O_905,N_3834,N_3752);
nand UO_906 (O_906,N_4414,N_2931);
nor UO_907 (O_907,N_4732,N_3217);
nand UO_908 (O_908,N_4446,N_4367);
nand UO_909 (O_909,N_4821,N_4661);
xnor UO_910 (O_910,N_4202,N_4021);
xnor UO_911 (O_911,N_3381,N_4268);
or UO_912 (O_912,N_3791,N_3605);
xnor UO_913 (O_913,N_2518,N_4522);
or UO_914 (O_914,N_4013,N_4344);
and UO_915 (O_915,N_4195,N_3235);
xnor UO_916 (O_916,N_3690,N_3418);
xnor UO_917 (O_917,N_3136,N_2520);
and UO_918 (O_918,N_3259,N_4604);
or UO_919 (O_919,N_3986,N_4318);
xor UO_920 (O_920,N_2903,N_4553);
or UO_921 (O_921,N_3895,N_2642);
nand UO_922 (O_922,N_2596,N_2644);
nor UO_923 (O_923,N_4735,N_3867);
or UO_924 (O_924,N_2998,N_2848);
or UO_925 (O_925,N_3126,N_4892);
xnor UO_926 (O_926,N_4577,N_3061);
xnor UO_927 (O_927,N_3328,N_2685);
nand UO_928 (O_928,N_4724,N_4430);
or UO_929 (O_929,N_3063,N_4388);
and UO_930 (O_930,N_4668,N_3991);
xnor UO_931 (O_931,N_2873,N_2548);
and UO_932 (O_932,N_4840,N_3094);
nand UO_933 (O_933,N_3114,N_3464);
nand UO_934 (O_934,N_3039,N_2657);
nor UO_935 (O_935,N_4087,N_4819);
xor UO_936 (O_936,N_3428,N_3918);
xor UO_937 (O_937,N_4740,N_2969);
and UO_938 (O_938,N_2945,N_4260);
nor UO_939 (O_939,N_4453,N_3739);
nor UO_940 (O_940,N_3400,N_3567);
nor UO_941 (O_941,N_3549,N_3819);
or UO_942 (O_942,N_2606,N_3594);
or UO_943 (O_943,N_3832,N_4944);
or UO_944 (O_944,N_4793,N_4731);
xor UO_945 (O_945,N_4332,N_2943);
xor UO_946 (O_946,N_3896,N_3072);
and UO_947 (O_947,N_3228,N_4092);
and UO_948 (O_948,N_4091,N_3552);
or UO_949 (O_949,N_3215,N_3462);
and UO_950 (O_950,N_4593,N_4548);
xor UO_951 (O_951,N_3020,N_3811);
or UO_952 (O_952,N_4127,N_2603);
or UO_953 (O_953,N_4852,N_4346);
nor UO_954 (O_954,N_4099,N_4630);
xor UO_955 (O_955,N_3358,N_3695);
xnor UO_956 (O_956,N_3116,N_4041);
or UO_957 (O_957,N_4272,N_2701);
nor UO_958 (O_958,N_2940,N_4569);
nor UO_959 (O_959,N_2680,N_3921);
nor UO_960 (O_960,N_4169,N_3362);
and UO_961 (O_961,N_4262,N_4333);
xor UO_962 (O_962,N_4103,N_4073);
and UO_963 (O_963,N_4479,N_4578);
nor UO_964 (O_964,N_4436,N_3023);
nand UO_965 (O_965,N_3006,N_4506);
and UO_966 (O_966,N_4057,N_2527);
nor UO_967 (O_967,N_3625,N_3646);
xnor UO_968 (O_968,N_3905,N_3470);
or UO_969 (O_969,N_3877,N_3657);
and UO_970 (O_970,N_2555,N_4807);
and UO_971 (O_971,N_3609,N_2506);
nor UO_972 (O_972,N_3974,N_4156);
nor UO_973 (O_973,N_3660,N_3740);
and UO_974 (O_974,N_3574,N_4751);
nor UO_975 (O_975,N_4649,N_3879);
nor UO_976 (O_976,N_2670,N_4858);
xnor UO_977 (O_977,N_3191,N_2841);
nor UO_978 (O_978,N_4290,N_4138);
nor UO_979 (O_979,N_3297,N_3608);
or UO_980 (O_980,N_3843,N_3152);
or UO_981 (O_981,N_3721,N_3787);
or UO_982 (O_982,N_3967,N_4864);
xor UO_983 (O_983,N_2705,N_2521);
or UO_984 (O_984,N_4875,N_3672);
or UO_985 (O_985,N_3484,N_4465);
xor UO_986 (O_986,N_3828,N_3450);
or UO_987 (O_987,N_3960,N_4020);
and UO_988 (O_988,N_2833,N_4596);
and UO_989 (O_989,N_4315,N_3768);
or UO_990 (O_990,N_3055,N_3153);
and UO_991 (O_991,N_4412,N_4891);
xor UO_992 (O_992,N_4275,N_4142);
xnor UO_993 (O_993,N_4371,N_4330);
nor UO_994 (O_994,N_4024,N_2813);
nor UO_995 (O_995,N_3697,N_2757);
nor UO_996 (O_996,N_4941,N_4083);
or UO_997 (O_997,N_3815,N_4337);
and UO_998 (O_998,N_4560,N_4801);
or UO_999 (O_999,N_3088,N_3261);
endmodule