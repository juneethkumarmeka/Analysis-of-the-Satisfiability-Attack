module basic_500_3000_500_60_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_362,In_353);
or U1 (N_1,In_267,In_305);
or U2 (N_2,In_250,In_135);
nand U3 (N_3,In_319,In_396);
nand U4 (N_4,In_74,In_175);
or U5 (N_5,In_314,In_11);
nor U6 (N_6,In_132,In_251);
nand U7 (N_7,In_219,In_234);
and U8 (N_8,In_370,In_321);
nor U9 (N_9,In_156,In_63);
nor U10 (N_10,In_170,In_382);
nand U11 (N_11,In_298,In_96);
and U12 (N_12,In_242,In_105);
or U13 (N_13,In_245,In_150);
nand U14 (N_14,In_355,In_66);
nor U15 (N_15,In_118,In_241);
and U16 (N_16,In_248,In_142);
nand U17 (N_17,In_369,In_34);
nor U18 (N_18,In_306,In_164);
nand U19 (N_19,In_104,In_32);
and U20 (N_20,In_457,In_498);
nor U21 (N_21,In_217,In_100);
xor U22 (N_22,In_123,In_349);
nor U23 (N_23,In_304,In_317);
and U24 (N_24,In_431,In_180);
nor U25 (N_25,In_129,In_299);
nor U26 (N_26,In_162,In_140);
and U27 (N_27,In_54,In_433);
nor U28 (N_28,In_337,In_324);
nand U29 (N_29,In_15,In_436);
nor U30 (N_30,In_177,In_266);
or U31 (N_31,In_57,In_309);
and U32 (N_32,In_228,In_237);
and U33 (N_33,In_290,In_310);
nor U34 (N_34,In_192,In_410);
xor U35 (N_35,In_292,In_161);
and U36 (N_36,In_80,In_480);
nand U37 (N_37,In_199,In_130);
and U38 (N_38,In_218,In_332);
xor U39 (N_39,In_81,In_411);
nor U40 (N_40,In_271,In_0);
nor U41 (N_41,In_18,In_416);
nand U42 (N_42,In_184,In_351);
or U43 (N_43,In_29,In_405);
nor U44 (N_44,In_52,In_1);
and U45 (N_45,In_190,In_253);
nor U46 (N_46,In_222,In_195);
xor U47 (N_47,In_260,In_256);
nor U48 (N_48,In_268,In_201);
and U49 (N_49,In_126,In_285);
nor U50 (N_50,In_350,In_45);
nand U51 (N_51,In_191,In_196);
xnor U52 (N_52,In_70,In_51);
nor U53 (N_53,In_68,In_72);
nor U54 (N_54,In_3,In_209);
nor U55 (N_55,In_122,In_139);
nand U56 (N_56,N_18,In_363);
or U57 (N_57,In_42,In_345);
or U58 (N_58,In_97,In_4);
or U59 (N_59,In_303,In_79);
nand U60 (N_60,In_360,In_99);
nand U61 (N_61,In_327,In_106);
xor U62 (N_62,In_472,In_427);
nor U63 (N_63,In_87,N_28);
and U64 (N_64,In_451,In_24);
or U65 (N_65,In_459,In_417);
or U66 (N_66,In_274,In_36);
and U67 (N_67,In_422,N_9);
nor U68 (N_68,In_110,N_11);
nor U69 (N_69,In_65,In_124);
and U70 (N_70,In_38,In_92);
nand U71 (N_71,In_2,In_346);
nor U72 (N_72,In_372,In_394);
nand U73 (N_73,In_377,In_93);
nand U74 (N_74,In_240,In_426);
and U75 (N_75,In_226,In_211);
and U76 (N_76,In_408,In_465);
nor U77 (N_77,In_461,In_114);
nor U78 (N_78,In_295,In_280);
nand U79 (N_79,In_398,N_32);
nor U80 (N_80,In_149,In_26);
or U81 (N_81,In_82,In_155);
or U82 (N_82,N_4,In_313);
and U83 (N_83,In_341,In_232);
nand U84 (N_84,In_16,In_278);
or U85 (N_85,In_255,In_335);
and U86 (N_86,In_151,In_58);
xor U87 (N_87,In_183,N_0);
or U88 (N_88,In_352,In_478);
nor U89 (N_89,N_41,In_159);
and U90 (N_90,N_14,In_147);
and U91 (N_91,In_41,In_273);
or U92 (N_92,In_276,In_378);
or U93 (N_93,In_146,In_154);
or U94 (N_94,In_144,N_40);
and U95 (N_95,In_419,In_482);
nand U96 (N_96,In_358,In_308);
nor U97 (N_97,In_456,In_27);
and U98 (N_98,In_148,N_21);
and U99 (N_99,In_495,N_7);
and U100 (N_100,In_171,N_71);
nand U101 (N_101,In_270,In_445);
nor U102 (N_102,N_99,In_434);
nand U103 (N_103,In_400,In_94);
and U104 (N_104,In_37,In_432);
and U105 (N_105,In_261,In_55);
and U106 (N_106,In_282,In_357);
and U107 (N_107,In_474,N_58);
and U108 (N_108,In_447,In_395);
or U109 (N_109,In_33,In_107);
or U110 (N_110,In_404,In_203);
and U111 (N_111,In_13,N_86);
nand U112 (N_112,In_64,In_497);
xor U113 (N_113,In_152,N_13);
nand U114 (N_114,In_44,In_71);
and U115 (N_115,In_75,In_393);
xnor U116 (N_116,In_289,In_412);
and U117 (N_117,In_479,In_375);
nor U118 (N_118,N_35,In_86);
and U119 (N_119,In_389,In_281);
and U120 (N_120,In_444,In_249);
or U121 (N_121,In_202,In_43);
nand U122 (N_122,In_379,In_493);
or U123 (N_123,In_439,In_56);
nand U124 (N_124,In_287,N_48);
nand U125 (N_125,In_12,In_334);
and U126 (N_126,In_198,N_67);
and U127 (N_127,In_224,In_157);
nand U128 (N_128,In_23,In_207);
or U129 (N_129,In_338,In_294);
and U130 (N_130,In_22,N_93);
nand U131 (N_131,In_463,In_301);
nor U132 (N_132,N_73,N_68);
xor U133 (N_133,In_46,In_429);
or U134 (N_134,N_81,In_437);
nor U135 (N_135,N_80,N_47);
and U136 (N_136,In_264,In_197);
and U137 (N_137,In_297,In_257);
and U138 (N_138,N_88,In_325);
nor U139 (N_139,N_27,In_210);
nor U140 (N_140,In_399,In_61);
nand U141 (N_141,In_484,In_101);
nand U142 (N_142,In_8,In_316);
and U143 (N_143,N_97,In_247);
or U144 (N_144,In_259,N_52);
nor U145 (N_145,N_3,In_442);
and U146 (N_146,In_258,N_49);
xnor U147 (N_147,In_499,In_31);
nand U148 (N_148,In_39,In_361);
xor U149 (N_149,In_356,N_63);
nor U150 (N_150,N_10,In_409);
nand U151 (N_151,In_403,In_112);
and U152 (N_152,In_134,In_166);
or U153 (N_153,N_44,In_453);
and U154 (N_154,N_95,N_57);
nand U155 (N_155,In_418,In_89);
nor U156 (N_156,N_123,In_21);
nand U157 (N_157,In_113,N_113);
or U158 (N_158,N_20,N_61);
and U159 (N_159,In_236,In_486);
and U160 (N_160,In_30,N_105);
nor U161 (N_161,N_6,N_39);
nor U162 (N_162,In_359,In_141);
or U163 (N_163,N_45,In_187);
nor U164 (N_164,In_269,N_34);
or U165 (N_165,In_168,In_145);
and U166 (N_166,In_492,In_227);
nand U167 (N_167,In_230,In_212);
and U168 (N_168,N_94,N_79);
nand U169 (N_169,In_223,N_96);
nand U170 (N_170,In_208,In_488);
nand U171 (N_171,In_200,In_179);
and U172 (N_172,In_452,In_231);
and U173 (N_173,In_387,In_318);
and U174 (N_174,N_117,N_147);
and U175 (N_175,In_435,N_130);
nand U176 (N_176,N_125,In_19);
xnor U177 (N_177,N_103,In_464);
and U178 (N_178,In_476,In_414);
xnor U179 (N_179,In_333,In_60);
and U180 (N_180,In_6,In_181);
or U181 (N_181,In_215,N_33);
and U182 (N_182,In_388,In_471);
and U183 (N_183,N_129,In_455);
or U184 (N_184,N_72,In_178);
and U185 (N_185,N_148,In_494);
and U186 (N_186,In_119,In_322);
or U187 (N_187,N_142,In_401);
nand U188 (N_188,N_1,N_124);
nand U189 (N_189,In_205,N_70);
nand U190 (N_190,In_214,In_448);
or U191 (N_191,N_126,N_98);
xor U192 (N_192,In_172,In_291);
and U193 (N_193,In_50,N_109);
nand U194 (N_194,In_347,N_134);
nor U195 (N_195,N_12,In_169);
nor U196 (N_196,In_336,In_128);
or U197 (N_197,In_40,In_225);
and U198 (N_198,In_47,N_36);
or U199 (N_199,N_118,In_425);
and U200 (N_200,N_102,In_78);
and U201 (N_201,In_485,In_252);
and U202 (N_202,In_467,N_139);
xor U203 (N_203,N_76,In_279);
or U204 (N_204,In_138,N_145);
and U205 (N_205,In_213,In_206);
nand U206 (N_206,In_460,N_43);
and U207 (N_207,N_23,N_16);
or U208 (N_208,In_91,In_468);
and U209 (N_209,N_55,N_29);
nor U210 (N_210,N_132,In_9);
or U211 (N_211,N_112,In_329);
nor U212 (N_212,In_189,In_328);
and U213 (N_213,N_136,In_176);
nor U214 (N_214,In_420,N_164);
nor U215 (N_215,In_311,N_169);
nand U216 (N_216,In_302,N_192);
or U217 (N_217,N_101,N_150);
or U218 (N_218,In_406,In_477);
nor U219 (N_219,N_92,N_135);
nand U220 (N_220,In_496,N_189);
nand U221 (N_221,N_168,N_153);
nand U222 (N_222,In_173,In_193);
nor U223 (N_223,N_15,In_20);
or U224 (N_224,N_184,N_177);
nand U225 (N_225,In_342,In_343);
nor U226 (N_226,N_106,In_383);
nand U227 (N_227,N_42,In_143);
nand U228 (N_228,N_143,In_466);
and U229 (N_229,In_428,N_172);
or U230 (N_230,N_46,N_90);
or U231 (N_231,N_50,N_56);
xor U232 (N_232,In_421,N_2);
nand U233 (N_233,In_108,In_331);
nand U234 (N_234,In_424,N_115);
and U235 (N_235,In_158,N_194);
nor U236 (N_236,N_131,In_376);
xnor U237 (N_237,N_108,In_137);
or U238 (N_238,N_195,In_83);
and U239 (N_239,In_481,N_65);
nand U240 (N_240,In_449,In_374);
nand U241 (N_241,In_111,In_28);
or U242 (N_242,In_185,In_483);
and U243 (N_243,N_83,N_154);
nand U244 (N_244,N_158,In_454);
nor U245 (N_245,N_91,N_133);
and U246 (N_246,In_423,In_339);
nand U247 (N_247,In_262,N_119);
nor U248 (N_248,N_162,N_127);
and U249 (N_249,N_5,N_151);
nand U250 (N_250,In_392,In_62);
and U251 (N_251,In_293,N_87);
nor U252 (N_252,N_100,In_386);
nand U253 (N_253,In_263,In_233);
or U254 (N_254,In_216,N_38);
nand U255 (N_255,In_446,N_75);
nor U256 (N_256,N_204,N_211);
and U257 (N_257,In_73,In_265);
or U258 (N_258,In_443,In_49);
nor U259 (N_259,N_229,In_131);
xnor U260 (N_260,In_127,In_284);
and U261 (N_261,N_110,In_121);
nand U262 (N_262,N_219,In_136);
nand U263 (N_263,In_229,N_206);
xnor U264 (N_264,In_373,In_85);
or U265 (N_265,N_233,In_491);
and U266 (N_266,N_104,N_19);
or U267 (N_267,N_221,In_275);
xnor U268 (N_268,In_165,N_141);
and U269 (N_269,N_239,N_238);
nor U270 (N_270,N_173,N_160);
nand U271 (N_271,In_186,N_196);
or U272 (N_272,N_248,N_213);
nor U273 (N_273,In_330,In_153);
nor U274 (N_274,N_144,In_163);
or U275 (N_275,In_48,N_121);
nor U276 (N_276,In_7,N_171);
and U277 (N_277,N_234,N_181);
or U278 (N_278,N_242,In_371);
nor U279 (N_279,N_180,N_156);
or U280 (N_280,In_125,In_277);
nand U281 (N_281,N_66,N_185);
and U282 (N_282,N_237,In_239);
or U283 (N_283,In_390,N_8);
nand U284 (N_284,N_24,N_223);
nor U285 (N_285,N_163,N_54);
and U286 (N_286,N_51,In_120);
xor U287 (N_287,N_85,In_77);
or U288 (N_288,In_194,N_186);
xnor U289 (N_289,In_340,N_60);
nand U290 (N_290,N_235,In_235);
nand U291 (N_291,In_367,In_364);
nand U292 (N_292,N_152,N_208);
and U293 (N_293,N_77,N_247);
nand U294 (N_294,In_441,In_490);
nand U295 (N_295,N_62,N_122);
and U296 (N_296,In_402,In_53);
and U297 (N_297,In_254,N_69);
and U298 (N_298,In_221,N_199);
or U299 (N_299,N_198,N_17);
nor U300 (N_300,N_289,N_25);
nor U301 (N_301,In_67,N_297);
and U302 (N_302,N_78,N_203);
or U303 (N_303,In_365,In_109);
nand U304 (N_304,N_283,N_157);
and U305 (N_305,N_228,N_114);
and U306 (N_306,N_232,N_222);
xor U307 (N_307,N_165,In_102);
nor U308 (N_308,N_187,N_274);
or U309 (N_309,N_281,N_251);
or U310 (N_310,N_245,In_133);
or U311 (N_311,In_413,N_250);
nor U312 (N_312,N_269,In_470);
and U313 (N_313,N_53,N_292);
nand U314 (N_314,In_160,N_120);
nand U315 (N_315,N_246,In_246);
xnor U316 (N_316,N_64,In_238);
nand U317 (N_317,In_475,N_230);
and U318 (N_318,N_262,N_182);
and U319 (N_319,N_202,In_17);
nand U320 (N_320,N_266,N_30);
and U321 (N_321,In_380,N_161);
nor U322 (N_322,N_155,In_307);
nor U323 (N_323,N_243,In_300);
nand U324 (N_324,In_283,N_37);
nor U325 (N_325,In_286,N_271);
or U326 (N_326,N_259,N_278);
nand U327 (N_327,In_35,N_215);
xor U328 (N_328,In_397,In_407);
nor U329 (N_329,In_462,N_216);
nand U330 (N_330,N_298,N_31);
or U331 (N_331,N_295,In_440);
xnor U332 (N_332,N_210,In_326);
or U333 (N_333,In_366,N_270);
and U334 (N_334,N_137,In_116);
and U335 (N_335,N_107,In_391);
nor U336 (N_336,In_95,N_138);
or U337 (N_337,N_146,N_116);
nand U338 (N_338,N_260,In_296);
nand U339 (N_339,In_5,N_267);
xnor U340 (N_340,In_204,In_84);
nand U341 (N_341,N_175,In_174);
or U342 (N_342,N_290,N_201);
or U343 (N_343,In_354,N_299);
nor U344 (N_344,N_74,N_288);
and U345 (N_345,In_90,N_258);
and U346 (N_346,N_276,N_149);
nor U347 (N_347,N_257,In_88);
nand U348 (N_348,N_190,N_220);
nand U349 (N_349,N_256,N_84);
or U350 (N_350,N_82,N_227);
nand U351 (N_351,N_111,N_179);
nor U352 (N_352,N_217,N_218);
or U353 (N_353,N_291,N_348);
or U354 (N_354,N_212,N_303);
or U355 (N_355,N_302,N_275);
and U356 (N_356,N_261,N_301);
xor U357 (N_357,N_22,N_263);
nor U358 (N_358,N_323,N_191);
and U359 (N_359,In_415,N_59);
nand U360 (N_360,N_89,N_240);
or U361 (N_361,N_337,N_342);
nor U362 (N_362,N_322,N_285);
nand U363 (N_363,In_312,In_385);
or U364 (N_364,In_469,In_117);
nand U365 (N_365,N_345,N_335);
nor U366 (N_366,N_252,N_170);
nor U367 (N_367,In_69,N_310);
and U368 (N_368,N_254,In_76);
xnor U369 (N_369,In_368,In_489);
and U370 (N_370,N_319,In_272);
nand U371 (N_371,N_317,N_325);
or U372 (N_372,N_339,In_188);
nand U373 (N_373,N_316,N_277);
or U374 (N_374,N_286,In_220);
and U375 (N_375,N_296,N_308);
or U376 (N_376,N_330,In_381);
nand U377 (N_377,N_272,N_255);
or U378 (N_378,N_231,N_26);
nand U379 (N_379,N_329,In_244);
nor U380 (N_380,N_284,N_331);
nand U381 (N_381,N_140,N_324);
nand U382 (N_382,In_458,N_318);
xor U383 (N_383,In_25,In_10);
xor U384 (N_384,N_320,In_344);
or U385 (N_385,N_214,In_438);
and U386 (N_386,N_264,N_306);
nor U387 (N_387,In_487,N_315);
nor U388 (N_388,N_309,N_349);
nand U389 (N_389,In_182,N_279);
and U390 (N_390,N_209,In_167);
nor U391 (N_391,In_320,In_450);
or U392 (N_392,In_430,N_332);
nor U393 (N_393,In_288,N_236);
nand U394 (N_394,N_341,N_343);
nor U395 (N_395,N_336,N_293);
nor U396 (N_396,N_265,In_59);
or U397 (N_397,In_243,In_348);
and U398 (N_398,N_268,N_327);
xnor U399 (N_399,N_321,N_188);
nand U400 (N_400,In_384,N_241);
nand U401 (N_401,N_379,N_249);
nand U402 (N_402,N_344,N_361);
nor U403 (N_403,N_367,N_225);
or U404 (N_404,N_382,N_282);
xnor U405 (N_405,N_244,N_313);
or U406 (N_406,N_352,N_340);
and U407 (N_407,N_128,N_386);
xor U408 (N_408,N_287,N_311);
and U409 (N_409,N_334,N_385);
nor U410 (N_410,N_300,In_473);
nand U411 (N_411,N_366,N_328);
xor U412 (N_412,N_197,N_387);
and U413 (N_413,N_273,N_372);
nand U414 (N_414,N_395,N_312);
nor U415 (N_415,N_369,N_380);
nand U416 (N_416,N_384,N_388);
and U417 (N_417,In_323,N_370);
and U418 (N_418,N_376,N_378);
and U419 (N_419,N_374,N_314);
and U420 (N_420,N_397,N_176);
nand U421 (N_421,In_14,N_207);
nor U422 (N_422,N_159,In_98);
and U423 (N_423,N_305,N_166);
and U424 (N_424,N_375,In_115);
nor U425 (N_425,N_354,N_357);
or U426 (N_426,N_398,N_193);
or U427 (N_427,N_304,N_362);
nand U428 (N_428,N_381,N_347);
and U429 (N_429,N_307,N_356);
nor U430 (N_430,N_373,N_280);
and U431 (N_431,In_315,N_183);
and U432 (N_432,N_253,N_205);
and U433 (N_433,N_294,N_371);
and U434 (N_434,N_351,N_360);
and U435 (N_435,N_346,N_224);
xnor U436 (N_436,N_368,N_167);
nor U437 (N_437,N_392,N_226);
and U438 (N_438,N_396,N_389);
nor U439 (N_439,N_383,N_394);
nor U440 (N_440,N_399,N_350);
nor U441 (N_441,N_365,N_358);
nand U442 (N_442,N_377,N_178);
and U443 (N_443,N_390,N_364);
and U444 (N_444,N_200,N_359);
and U445 (N_445,N_393,N_333);
or U446 (N_446,N_338,N_355);
nand U447 (N_447,N_353,N_174);
and U448 (N_448,In_103,N_363);
or U449 (N_449,N_391,N_326);
nand U450 (N_450,N_423,N_424);
nand U451 (N_451,N_430,N_411);
nor U452 (N_452,N_432,N_413);
or U453 (N_453,N_406,N_402);
or U454 (N_454,N_415,N_418);
nand U455 (N_455,N_443,N_404);
nand U456 (N_456,N_449,N_440);
or U457 (N_457,N_435,N_436);
nand U458 (N_458,N_419,N_409);
or U459 (N_459,N_437,N_431);
xnor U460 (N_460,N_407,N_427);
nand U461 (N_461,N_448,N_434);
or U462 (N_462,N_414,N_410);
nand U463 (N_463,N_429,N_439);
or U464 (N_464,N_446,N_428);
nor U465 (N_465,N_420,N_417);
nor U466 (N_466,N_433,N_421);
or U467 (N_467,N_401,N_425);
and U468 (N_468,N_408,N_412);
or U469 (N_469,N_445,N_416);
nand U470 (N_470,N_441,N_447);
nand U471 (N_471,N_405,N_403);
or U472 (N_472,N_438,N_422);
nor U473 (N_473,N_426,N_442);
or U474 (N_474,N_444,N_400);
nand U475 (N_475,N_436,N_401);
xnor U476 (N_476,N_432,N_441);
nor U477 (N_477,N_442,N_405);
or U478 (N_478,N_415,N_448);
and U479 (N_479,N_410,N_447);
xnor U480 (N_480,N_410,N_428);
and U481 (N_481,N_419,N_421);
xnor U482 (N_482,N_439,N_400);
or U483 (N_483,N_439,N_408);
nor U484 (N_484,N_418,N_427);
and U485 (N_485,N_401,N_442);
and U486 (N_486,N_430,N_414);
nand U487 (N_487,N_407,N_445);
and U488 (N_488,N_414,N_433);
and U489 (N_489,N_448,N_412);
and U490 (N_490,N_436,N_420);
nand U491 (N_491,N_402,N_429);
nand U492 (N_492,N_405,N_421);
and U493 (N_493,N_417,N_412);
and U494 (N_494,N_427,N_428);
and U495 (N_495,N_414,N_418);
and U496 (N_496,N_449,N_428);
nor U497 (N_497,N_402,N_426);
and U498 (N_498,N_430,N_420);
and U499 (N_499,N_426,N_406);
nand U500 (N_500,N_487,N_477);
nand U501 (N_501,N_478,N_499);
or U502 (N_502,N_466,N_458);
or U503 (N_503,N_484,N_495);
or U504 (N_504,N_453,N_457);
and U505 (N_505,N_463,N_486);
xnor U506 (N_506,N_492,N_472);
nand U507 (N_507,N_459,N_493);
nor U508 (N_508,N_452,N_496);
and U509 (N_509,N_450,N_455);
nand U510 (N_510,N_470,N_473);
xor U511 (N_511,N_482,N_488);
nand U512 (N_512,N_489,N_467);
nand U513 (N_513,N_454,N_498);
nand U514 (N_514,N_474,N_461);
nor U515 (N_515,N_494,N_490);
xor U516 (N_516,N_491,N_485);
nand U517 (N_517,N_451,N_469);
xor U518 (N_518,N_475,N_471);
nor U519 (N_519,N_479,N_481);
nand U520 (N_520,N_476,N_483);
or U521 (N_521,N_468,N_497);
and U522 (N_522,N_460,N_462);
and U523 (N_523,N_464,N_480);
or U524 (N_524,N_465,N_456);
nor U525 (N_525,N_483,N_499);
nand U526 (N_526,N_483,N_454);
and U527 (N_527,N_462,N_498);
nor U528 (N_528,N_471,N_473);
nor U529 (N_529,N_467,N_469);
nand U530 (N_530,N_476,N_462);
nand U531 (N_531,N_461,N_467);
nand U532 (N_532,N_457,N_450);
and U533 (N_533,N_473,N_493);
nand U534 (N_534,N_470,N_486);
and U535 (N_535,N_489,N_493);
nand U536 (N_536,N_491,N_473);
nand U537 (N_537,N_488,N_477);
nand U538 (N_538,N_459,N_489);
nor U539 (N_539,N_479,N_470);
nor U540 (N_540,N_475,N_463);
or U541 (N_541,N_470,N_453);
nand U542 (N_542,N_476,N_452);
and U543 (N_543,N_463,N_471);
or U544 (N_544,N_488,N_461);
and U545 (N_545,N_450,N_483);
and U546 (N_546,N_485,N_460);
or U547 (N_547,N_478,N_453);
nor U548 (N_548,N_460,N_496);
xor U549 (N_549,N_478,N_479);
nand U550 (N_550,N_528,N_541);
or U551 (N_551,N_518,N_513);
or U552 (N_552,N_521,N_530);
or U553 (N_553,N_516,N_549);
nor U554 (N_554,N_531,N_509);
nor U555 (N_555,N_517,N_511);
or U556 (N_556,N_547,N_525);
and U557 (N_557,N_505,N_540);
nor U558 (N_558,N_510,N_519);
nor U559 (N_559,N_512,N_535);
and U560 (N_560,N_542,N_504);
and U561 (N_561,N_532,N_537);
nand U562 (N_562,N_506,N_523);
nand U563 (N_563,N_522,N_545);
or U564 (N_564,N_529,N_526);
nand U565 (N_565,N_500,N_539);
nor U566 (N_566,N_548,N_520);
or U567 (N_567,N_514,N_502);
or U568 (N_568,N_524,N_534);
or U569 (N_569,N_503,N_546);
nor U570 (N_570,N_538,N_536);
and U571 (N_571,N_501,N_527);
nand U572 (N_572,N_508,N_544);
or U573 (N_573,N_507,N_515);
nor U574 (N_574,N_533,N_543);
xor U575 (N_575,N_546,N_526);
nor U576 (N_576,N_511,N_504);
nand U577 (N_577,N_549,N_520);
nor U578 (N_578,N_510,N_542);
nor U579 (N_579,N_537,N_513);
or U580 (N_580,N_542,N_533);
or U581 (N_581,N_502,N_523);
nor U582 (N_582,N_514,N_526);
xnor U583 (N_583,N_538,N_515);
nand U584 (N_584,N_531,N_526);
and U585 (N_585,N_538,N_513);
nor U586 (N_586,N_521,N_535);
nand U587 (N_587,N_522,N_513);
xor U588 (N_588,N_513,N_526);
and U589 (N_589,N_517,N_503);
or U590 (N_590,N_515,N_545);
nor U591 (N_591,N_533,N_500);
and U592 (N_592,N_525,N_522);
or U593 (N_593,N_530,N_526);
and U594 (N_594,N_503,N_536);
or U595 (N_595,N_520,N_529);
xor U596 (N_596,N_523,N_518);
nand U597 (N_597,N_543,N_505);
xor U598 (N_598,N_524,N_547);
or U599 (N_599,N_534,N_526);
xor U600 (N_600,N_557,N_569);
or U601 (N_601,N_591,N_570);
nor U602 (N_602,N_597,N_556);
nand U603 (N_603,N_580,N_581);
nand U604 (N_604,N_595,N_592);
nand U605 (N_605,N_579,N_565);
nor U606 (N_606,N_566,N_551);
nor U607 (N_607,N_589,N_584);
or U608 (N_608,N_572,N_564);
and U609 (N_609,N_582,N_554);
or U610 (N_610,N_594,N_562);
and U611 (N_611,N_586,N_598);
and U612 (N_612,N_590,N_575);
nor U613 (N_613,N_555,N_587);
or U614 (N_614,N_577,N_573);
nand U615 (N_615,N_593,N_558);
and U616 (N_616,N_561,N_560);
xor U617 (N_617,N_553,N_550);
nor U618 (N_618,N_599,N_578);
nand U619 (N_619,N_571,N_576);
nand U620 (N_620,N_552,N_559);
or U621 (N_621,N_588,N_568);
and U622 (N_622,N_567,N_585);
or U623 (N_623,N_583,N_596);
nor U624 (N_624,N_574,N_563);
or U625 (N_625,N_551,N_572);
and U626 (N_626,N_579,N_568);
and U627 (N_627,N_570,N_565);
nor U628 (N_628,N_580,N_570);
nand U629 (N_629,N_559,N_567);
xnor U630 (N_630,N_571,N_584);
nand U631 (N_631,N_572,N_562);
nor U632 (N_632,N_552,N_597);
nand U633 (N_633,N_561,N_595);
and U634 (N_634,N_556,N_592);
nor U635 (N_635,N_554,N_583);
xor U636 (N_636,N_554,N_584);
nor U637 (N_637,N_597,N_599);
nor U638 (N_638,N_584,N_555);
nand U639 (N_639,N_554,N_553);
nand U640 (N_640,N_560,N_570);
nand U641 (N_641,N_550,N_566);
or U642 (N_642,N_561,N_567);
and U643 (N_643,N_553,N_593);
nor U644 (N_644,N_550,N_567);
or U645 (N_645,N_561,N_556);
nand U646 (N_646,N_576,N_581);
xnor U647 (N_647,N_596,N_560);
xnor U648 (N_648,N_598,N_571);
nand U649 (N_649,N_551,N_552);
or U650 (N_650,N_645,N_615);
nand U651 (N_651,N_640,N_625);
or U652 (N_652,N_638,N_602);
and U653 (N_653,N_611,N_614);
and U654 (N_654,N_608,N_637);
nand U655 (N_655,N_631,N_634);
or U656 (N_656,N_649,N_635);
nor U657 (N_657,N_621,N_606);
nor U658 (N_658,N_639,N_646);
and U659 (N_659,N_628,N_603);
or U660 (N_660,N_647,N_605);
nand U661 (N_661,N_623,N_636);
nand U662 (N_662,N_642,N_600);
nor U663 (N_663,N_616,N_619);
nor U664 (N_664,N_630,N_632);
or U665 (N_665,N_620,N_613);
xnor U666 (N_666,N_643,N_618);
nand U667 (N_667,N_629,N_627);
xnor U668 (N_668,N_607,N_633);
and U669 (N_669,N_604,N_609);
or U670 (N_670,N_641,N_624);
and U671 (N_671,N_626,N_617);
or U672 (N_672,N_622,N_610);
nor U673 (N_673,N_644,N_612);
nor U674 (N_674,N_648,N_601);
xor U675 (N_675,N_625,N_604);
nor U676 (N_676,N_628,N_636);
nand U677 (N_677,N_634,N_614);
nand U678 (N_678,N_639,N_628);
or U679 (N_679,N_600,N_613);
nor U680 (N_680,N_648,N_606);
xor U681 (N_681,N_624,N_636);
nand U682 (N_682,N_616,N_634);
nand U683 (N_683,N_648,N_636);
and U684 (N_684,N_619,N_642);
nor U685 (N_685,N_646,N_630);
xnor U686 (N_686,N_625,N_633);
or U687 (N_687,N_644,N_634);
nand U688 (N_688,N_629,N_625);
nand U689 (N_689,N_629,N_613);
nand U690 (N_690,N_613,N_639);
or U691 (N_691,N_637,N_623);
and U692 (N_692,N_602,N_643);
nor U693 (N_693,N_636,N_619);
or U694 (N_694,N_605,N_615);
nand U695 (N_695,N_638,N_642);
nand U696 (N_696,N_624,N_630);
xnor U697 (N_697,N_636,N_634);
xor U698 (N_698,N_645,N_606);
or U699 (N_699,N_635,N_600);
and U700 (N_700,N_678,N_684);
nor U701 (N_701,N_666,N_670);
nand U702 (N_702,N_660,N_694);
nor U703 (N_703,N_671,N_652);
xnor U704 (N_704,N_695,N_655);
nor U705 (N_705,N_682,N_650);
xnor U706 (N_706,N_672,N_685);
nand U707 (N_707,N_657,N_661);
nand U708 (N_708,N_692,N_683);
and U709 (N_709,N_680,N_658);
nand U710 (N_710,N_679,N_659);
and U711 (N_711,N_691,N_664);
and U712 (N_712,N_689,N_673);
nor U713 (N_713,N_698,N_665);
nor U714 (N_714,N_686,N_697);
nor U715 (N_715,N_693,N_699);
or U716 (N_716,N_668,N_663);
and U717 (N_717,N_667,N_656);
xor U718 (N_718,N_662,N_651);
or U719 (N_719,N_677,N_681);
nand U720 (N_720,N_654,N_675);
nand U721 (N_721,N_674,N_690);
nand U722 (N_722,N_687,N_688);
or U723 (N_723,N_696,N_676);
nand U724 (N_724,N_669,N_653);
nor U725 (N_725,N_666,N_694);
nand U726 (N_726,N_668,N_655);
nand U727 (N_727,N_660,N_675);
nand U728 (N_728,N_664,N_666);
nand U729 (N_729,N_651,N_676);
nor U730 (N_730,N_684,N_686);
nand U731 (N_731,N_662,N_654);
nand U732 (N_732,N_678,N_677);
nand U733 (N_733,N_651,N_654);
nand U734 (N_734,N_674,N_683);
and U735 (N_735,N_695,N_664);
or U736 (N_736,N_668,N_684);
and U737 (N_737,N_656,N_682);
nor U738 (N_738,N_659,N_652);
or U739 (N_739,N_670,N_656);
or U740 (N_740,N_653,N_671);
and U741 (N_741,N_673,N_663);
or U742 (N_742,N_678,N_680);
nor U743 (N_743,N_663,N_672);
xnor U744 (N_744,N_661,N_685);
nand U745 (N_745,N_669,N_693);
and U746 (N_746,N_676,N_679);
nor U747 (N_747,N_655,N_696);
nor U748 (N_748,N_658,N_672);
nor U749 (N_749,N_652,N_684);
and U750 (N_750,N_708,N_733);
nor U751 (N_751,N_740,N_712);
xor U752 (N_752,N_709,N_736);
nand U753 (N_753,N_747,N_745);
nand U754 (N_754,N_732,N_720);
nand U755 (N_755,N_706,N_710);
nor U756 (N_756,N_748,N_744);
nor U757 (N_757,N_734,N_716);
or U758 (N_758,N_713,N_707);
xor U759 (N_759,N_727,N_749);
or U760 (N_760,N_738,N_743);
xnor U761 (N_761,N_739,N_741);
and U762 (N_762,N_735,N_705);
and U763 (N_763,N_702,N_719);
nor U764 (N_764,N_746,N_724);
nand U765 (N_765,N_731,N_742);
or U766 (N_766,N_717,N_718);
nand U767 (N_767,N_726,N_729);
nand U768 (N_768,N_714,N_725);
or U769 (N_769,N_700,N_704);
and U770 (N_770,N_722,N_721);
nand U771 (N_771,N_723,N_715);
nand U772 (N_772,N_730,N_737);
or U773 (N_773,N_701,N_703);
nor U774 (N_774,N_711,N_728);
xor U775 (N_775,N_740,N_735);
and U776 (N_776,N_741,N_729);
xnor U777 (N_777,N_707,N_716);
and U778 (N_778,N_740,N_718);
nor U779 (N_779,N_748,N_710);
and U780 (N_780,N_730,N_726);
xnor U781 (N_781,N_712,N_742);
or U782 (N_782,N_714,N_727);
and U783 (N_783,N_719,N_744);
nor U784 (N_784,N_710,N_705);
nor U785 (N_785,N_742,N_744);
and U786 (N_786,N_702,N_747);
or U787 (N_787,N_700,N_707);
or U788 (N_788,N_732,N_707);
nor U789 (N_789,N_727,N_737);
and U790 (N_790,N_748,N_712);
or U791 (N_791,N_704,N_749);
and U792 (N_792,N_717,N_727);
nand U793 (N_793,N_718,N_749);
xor U794 (N_794,N_724,N_740);
or U795 (N_795,N_707,N_749);
nand U796 (N_796,N_709,N_708);
nand U797 (N_797,N_733,N_748);
nor U798 (N_798,N_716,N_747);
and U799 (N_799,N_749,N_744);
nand U800 (N_800,N_765,N_775);
nand U801 (N_801,N_785,N_780);
or U802 (N_802,N_786,N_773);
and U803 (N_803,N_768,N_750);
and U804 (N_804,N_792,N_756);
nand U805 (N_805,N_753,N_771);
nand U806 (N_806,N_793,N_794);
nand U807 (N_807,N_760,N_778);
and U808 (N_808,N_774,N_766);
or U809 (N_809,N_797,N_762);
or U810 (N_810,N_776,N_751);
nand U811 (N_811,N_798,N_795);
and U812 (N_812,N_777,N_781);
xor U813 (N_813,N_790,N_761);
and U814 (N_814,N_796,N_782);
nand U815 (N_815,N_791,N_764);
nor U816 (N_816,N_789,N_779);
and U817 (N_817,N_769,N_770);
nand U818 (N_818,N_767,N_799);
nor U819 (N_819,N_755,N_757);
nor U820 (N_820,N_763,N_752);
nor U821 (N_821,N_787,N_788);
nor U822 (N_822,N_783,N_754);
nand U823 (N_823,N_758,N_759);
xor U824 (N_824,N_772,N_784);
or U825 (N_825,N_799,N_790);
nand U826 (N_826,N_764,N_787);
nand U827 (N_827,N_755,N_784);
nor U828 (N_828,N_796,N_771);
or U829 (N_829,N_760,N_753);
nor U830 (N_830,N_762,N_756);
nand U831 (N_831,N_772,N_761);
nand U832 (N_832,N_790,N_779);
or U833 (N_833,N_778,N_752);
xor U834 (N_834,N_783,N_773);
and U835 (N_835,N_757,N_789);
nand U836 (N_836,N_750,N_758);
and U837 (N_837,N_770,N_765);
or U838 (N_838,N_757,N_768);
nand U839 (N_839,N_793,N_752);
nor U840 (N_840,N_792,N_768);
or U841 (N_841,N_752,N_754);
or U842 (N_842,N_761,N_777);
and U843 (N_843,N_794,N_774);
nor U844 (N_844,N_753,N_773);
and U845 (N_845,N_760,N_767);
nor U846 (N_846,N_766,N_764);
or U847 (N_847,N_763,N_762);
or U848 (N_848,N_752,N_760);
nor U849 (N_849,N_798,N_799);
or U850 (N_850,N_821,N_819);
xnor U851 (N_851,N_833,N_849);
or U852 (N_852,N_802,N_845);
nand U853 (N_853,N_837,N_809);
and U854 (N_854,N_822,N_801);
xnor U855 (N_855,N_805,N_836);
nor U856 (N_856,N_839,N_800);
nor U857 (N_857,N_825,N_831);
xor U858 (N_858,N_838,N_846);
or U859 (N_859,N_824,N_826);
nand U860 (N_860,N_827,N_812);
or U861 (N_861,N_830,N_807);
and U862 (N_862,N_840,N_803);
nor U863 (N_863,N_844,N_848);
nor U864 (N_864,N_817,N_847);
and U865 (N_865,N_832,N_829);
xor U866 (N_866,N_806,N_823);
nand U867 (N_867,N_804,N_843);
or U868 (N_868,N_813,N_816);
xnor U869 (N_869,N_841,N_810);
nor U870 (N_870,N_811,N_835);
or U871 (N_871,N_834,N_808);
nor U872 (N_872,N_814,N_828);
nand U873 (N_873,N_818,N_815);
or U874 (N_874,N_842,N_820);
nand U875 (N_875,N_846,N_841);
nand U876 (N_876,N_825,N_823);
nor U877 (N_877,N_841,N_828);
nor U878 (N_878,N_803,N_841);
nand U879 (N_879,N_821,N_806);
and U880 (N_880,N_840,N_813);
and U881 (N_881,N_832,N_807);
nand U882 (N_882,N_842,N_826);
nand U883 (N_883,N_832,N_808);
nand U884 (N_884,N_840,N_828);
nand U885 (N_885,N_830,N_848);
and U886 (N_886,N_837,N_816);
nand U887 (N_887,N_815,N_846);
nor U888 (N_888,N_821,N_849);
or U889 (N_889,N_848,N_840);
or U890 (N_890,N_827,N_834);
and U891 (N_891,N_822,N_811);
or U892 (N_892,N_846,N_843);
nor U893 (N_893,N_816,N_833);
or U894 (N_894,N_846,N_807);
nor U895 (N_895,N_809,N_802);
nor U896 (N_896,N_830,N_833);
or U897 (N_897,N_841,N_843);
nand U898 (N_898,N_813,N_839);
and U899 (N_899,N_848,N_806);
xor U900 (N_900,N_883,N_877);
nand U901 (N_901,N_865,N_862);
or U902 (N_902,N_899,N_864);
or U903 (N_903,N_876,N_889);
xnor U904 (N_904,N_891,N_884);
and U905 (N_905,N_888,N_857);
nand U906 (N_906,N_885,N_875);
nand U907 (N_907,N_863,N_892);
or U908 (N_908,N_855,N_869);
or U909 (N_909,N_890,N_868);
nand U910 (N_910,N_882,N_893);
or U911 (N_911,N_859,N_870);
or U912 (N_912,N_852,N_872);
nor U913 (N_913,N_860,N_871);
or U914 (N_914,N_861,N_856);
nand U915 (N_915,N_897,N_874);
or U916 (N_916,N_854,N_851);
and U917 (N_917,N_853,N_894);
nand U918 (N_918,N_850,N_866);
xor U919 (N_919,N_898,N_858);
nand U920 (N_920,N_878,N_887);
and U921 (N_921,N_896,N_881);
or U922 (N_922,N_867,N_873);
and U923 (N_923,N_886,N_879);
nor U924 (N_924,N_880,N_895);
or U925 (N_925,N_854,N_857);
or U926 (N_926,N_878,N_854);
nor U927 (N_927,N_896,N_886);
nand U928 (N_928,N_880,N_864);
and U929 (N_929,N_853,N_875);
and U930 (N_930,N_896,N_865);
nor U931 (N_931,N_870,N_885);
nor U932 (N_932,N_866,N_875);
nand U933 (N_933,N_867,N_865);
nor U934 (N_934,N_877,N_898);
xnor U935 (N_935,N_886,N_851);
or U936 (N_936,N_869,N_870);
nand U937 (N_937,N_857,N_874);
or U938 (N_938,N_867,N_895);
nor U939 (N_939,N_894,N_896);
nand U940 (N_940,N_867,N_871);
nor U941 (N_941,N_861,N_852);
and U942 (N_942,N_880,N_853);
and U943 (N_943,N_890,N_871);
xnor U944 (N_944,N_856,N_878);
and U945 (N_945,N_854,N_858);
or U946 (N_946,N_894,N_879);
nand U947 (N_947,N_889,N_859);
xor U948 (N_948,N_853,N_893);
or U949 (N_949,N_877,N_889);
nor U950 (N_950,N_942,N_914);
or U951 (N_951,N_935,N_933);
nand U952 (N_952,N_948,N_903);
nand U953 (N_953,N_909,N_949);
xnor U954 (N_954,N_922,N_943);
or U955 (N_955,N_908,N_930);
or U956 (N_956,N_915,N_927);
nand U957 (N_957,N_916,N_911);
nor U958 (N_958,N_910,N_929);
or U959 (N_959,N_934,N_925);
nand U960 (N_960,N_939,N_924);
and U961 (N_961,N_928,N_944);
xor U962 (N_962,N_905,N_923);
nand U963 (N_963,N_906,N_921);
nor U964 (N_964,N_920,N_919);
nor U965 (N_965,N_947,N_936);
or U966 (N_966,N_912,N_926);
or U967 (N_967,N_938,N_907);
and U968 (N_968,N_918,N_900);
or U969 (N_969,N_931,N_932);
xor U970 (N_970,N_940,N_937);
nand U971 (N_971,N_946,N_901);
xnor U972 (N_972,N_941,N_904);
or U973 (N_973,N_917,N_945);
nor U974 (N_974,N_913,N_902);
or U975 (N_975,N_911,N_933);
nand U976 (N_976,N_917,N_943);
and U977 (N_977,N_938,N_927);
or U978 (N_978,N_910,N_934);
nor U979 (N_979,N_926,N_930);
and U980 (N_980,N_937,N_935);
or U981 (N_981,N_908,N_943);
nor U982 (N_982,N_940,N_915);
nor U983 (N_983,N_922,N_941);
and U984 (N_984,N_901,N_931);
and U985 (N_985,N_928,N_936);
xor U986 (N_986,N_947,N_903);
or U987 (N_987,N_908,N_907);
or U988 (N_988,N_906,N_917);
or U989 (N_989,N_909,N_912);
nor U990 (N_990,N_919,N_917);
or U991 (N_991,N_921,N_929);
nand U992 (N_992,N_944,N_912);
nor U993 (N_993,N_904,N_911);
or U994 (N_994,N_927,N_930);
or U995 (N_995,N_900,N_934);
xnor U996 (N_996,N_901,N_924);
nor U997 (N_997,N_906,N_945);
nand U998 (N_998,N_917,N_913);
nand U999 (N_999,N_925,N_948);
and U1000 (N_1000,N_972,N_977);
nand U1001 (N_1001,N_989,N_994);
and U1002 (N_1002,N_984,N_992);
or U1003 (N_1003,N_990,N_970);
nor U1004 (N_1004,N_983,N_968);
or U1005 (N_1005,N_950,N_976);
nand U1006 (N_1006,N_986,N_978);
or U1007 (N_1007,N_952,N_960);
nand U1008 (N_1008,N_967,N_957);
nor U1009 (N_1009,N_962,N_999);
and U1010 (N_1010,N_963,N_966);
and U1011 (N_1011,N_965,N_988);
nand U1012 (N_1012,N_997,N_958);
and U1013 (N_1013,N_974,N_953);
or U1014 (N_1014,N_954,N_951);
nand U1015 (N_1015,N_996,N_979);
nor U1016 (N_1016,N_964,N_982);
and U1017 (N_1017,N_975,N_956);
and U1018 (N_1018,N_993,N_955);
or U1019 (N_1019,N_985,N_961);
or U1020 (N_1020,N_969,N_998);
and U1021 (N_1021,N_995,N_959);
xnor U1022 (N_1022,N_973,N_980);
or U1023 (N_1023,N_987,N_991);
nor U1024 (N_1024,N_971,N_981);
nand U1025 (N_1025,N_996,N_977);
xnor U1026 (N_1026,N_992,N_968);
or U1027 (N_1027,N_963,N_968);
and U1028 (N_1028,N_960,N_963);
nor U1029 (N_1029,N_978,N_980);
or U1030 (N_1030,N_951,N_950);
or U1031 (N_1031,N_975,N_965);
or U1032 (N_1032,N_964,N_993);
nor U1033 (N_1033,N_989,N_963);
and U1034 (N_1034,N_962,N_998);
or U1035 (N_1035,N_952,N_998);
nand U1036 (N_1036,N_961,N_994);
nor U1037 (N_1037,N_993,N_954);
and U1038 (N_1038,N_992,N_980);
and U1039 (N_1039,N_956,N_968);
or U1040 (N_1040,N_975,N_996);
xor U1041 (N_1041,N_982,N_951);
and U1042 (N_1042,N_958,N_966);
and U1043 (N_1043,N_978,N_957);
and U1044 (N_1044,N_972,N_996);
and U1045 (N_1045,N_975,N_983);
nor U1046 (N_1046,N_955,N_983);
and U1047 (N_1047,N_977,N_995);
and U1048 (N_1048,N_951,N_971);
or U1049 (N_1049,N_950,N_952);
and U1050 (N_1050,N_1024,N_1011);
xnor U1051 (N_1051,N_1018,N_1013);
nand U1052 (N_1052,N_1043,N_1045);
nor U1053 (N_1053,N_1030,N_1047);
or U1054 (N_1054,N_1029,N_1025);
or U1055 (N_1055,N_1017,N_1026);
nand U1056 (N_1056,N_1044,N_1023);
nor U1057 (N_1057,N_1021,N_1033);
nand U1058 (N_1058,N_1014,N_1041);
nand U1059 (N_1059,N_1016,N_1027);
or U1060 (N_1060,N_1005,N_1010);
nor U1061 (N_1061,N_1036,N_1006);
nand U1062 (N_1062,N_1042,N_1001);
nand U1063 (N_1063,N_1008,N_1012);
nand U1064 (N_1064,N_1046,N_1038);
nor U1065 (N_1065,N_1002,N_1004);
nand U1066 (N_1066,N_1000,N_1007);
xnor U1067 (N_1067,N_1028,N_1019);
nor U1068 (N_1068,N_1040,N_1031);
and U1069 (N_1069,N_1039,N_1003);
nor U1070 (N_1070,N_1049,N_1032);
nand U1071 (N_1071,N_1020,N_1037);
nand U1072 (N_1072,N_1022,N_1009);
and U1073 (N_1073,N_1015,N_1034);
or U1074 (N_1074,N_1035,N_1048);
nand U1075 (N_1075,N_1043,N_1037);
or U1076 (N_1076,N_1000,N_1040);
nand U1077 (N_1077,N_1035,N_1004);
nor U1078 (N_1078,N_1007,N_1002);
and U1079 (N_1079,N_1016,N_1018);
nor U1080 (N_1080,N_1044,N_1003);
nand U1081 (N_1081,N_1008,N_1034);
nor U1082 (N_1082,N_1013,N_1025);
or U1083 (N_1083,N_1021,N_1014);
xor U1084 (N_1084,N_1047,N_1046);
nand U1085 (N_1085,N_1021,N_1042);
or U1086 (N_1086,N_1016,N_1030);
or U1087 (N_1087,N_1020,N_1018);
or U1088 (N_1088,N_1034,N_1048);
nand U1089 (N_1089,N_1036,N_1041);
nor U1090 (N_1090,N_1049,N_1010);
nand U1091 (N_1091,N_1042,N_1034);
and U1092 (N_1092,N_1012,N_1044);
or U1093 (N_1093,N_1022,N_1021);
or U1094 (N_1094,N_1027,N_1009);
and U1095 (N_1095,N_1030,N_1044);
xor U1096 (N_1096,N_1029,N_1019);
nor U1097 (N_1097,N_1044,N_1037);
nand U1098 (N_1098,N_1036,N_1046);
and U1099 (N_1099,N_1040,N_1024);
xnor U1100 (N_1100,N_1097,N_1098);
and U1101 (N_1101,N_1095,N_1080);
and U1102 (N_1102,N_1050,N_1072);
nand U1103 (N_1103,N_1089,N_1063);
nand U1104 (N_1104,N_1082,N_1099);
xnor U1105 (N_1105,N_1071,N_1051);
nor U1106 (N_1106,N_1086,N_1078);
nor U1107 (N_1107,N_1077,N_1064);
nor U1108 (N_1108,N_1079,N_1094);
nor U1109 (N_1109,N_1076,N_1059);
xnor U1110 (N_1110,N_1074,N_1068);
or U1111 (N_1111,N_1075,N_1083);
nor U1112 (N_1112,N_1070,N_1084);
nand U1113 (N_1113,N_1081,N_1053);
nor U1114 (N_1114,N_1069,N_1073);
nand U1115 (N_1115,N_1054,N_1092);
and U1116 (N_1116,N_1052,N_1066);
nor U1117 (N_1117,N_1091,N_1087);
xnor U1118 (N_1118,N_1061,N_1096);
nor U1119 (N_1119,N_1085,N_1058);
nand U1120 (N_1120,N_1062,N_1067);
and U1121 (N_1121,N_1090,N_1065);
nor U1122 (N_1122,N_1093,N_1056);
nor U1123 (N_1123,N_1060,N_1055);
xor U1124 (N_1124,N_1088,N_1057);
nor U1125 (N_1125,N_1073,N_1099);
and U1126 (N_1126,N_1088,N_1050);
nor U1127 (N_1127,N_1061,N_1071);
or U1128 (N_1128,N_1056,N_1055);
nor U1129 (N_1129,N_1087,N_1095);
nand U1130 (N_1130,N_1064,N_1094);
nand U1131 (N_1131,N_1052,N_1084);
nand U1132 (N_1132,N_1070,N_1088);
nor U1133 (N_1133,N_1084,N_1092);
nor U1134 (N_1134,N_1064,N_1068);
nand U1135 (N_1135,N_1057,N_1055);
and U1136 (N_1136,N_1070,N_1053);
nand U1137 (N_1137,N_1052,N_1056);
or U1138 (N_1138,N_1091,N_1061);
and U1139 (N_1139,N_1083,N_1055);
and U1140 (N_1140,N_1055,N_1073);
or U1141 (N_1141,N_1065,N_1092);
or U1142 (N_1142,N_1054,N_1060);
nor U1143 (N_1143,N_1086,N_1085);
or U1144 (N_1144,N_1080,N_1055);
nand U1145 (N_1145,N_1078,N_1098);
and U1146 (N_1146,N_1071,N_1072);
xnor U1147 (N_1147,N_1051,N_1079);
nand U1148 (N_1148,N_1061,N_1068);
nor U1149 (N_1149,N_1099,N_1087);
nand U1150 (N_1150,N_1115,N_1135);
nand U1151 (N_1151,N_1118,N_1127);
nand U1152 (N_1152,N_1108,N_1116);
nor U1153 (N_1153,N_1141,N_1129);
nor U1154 (N_1154,N_1146,N_1110);
and U1155 (N_1155,N_1119,N_1101);
or U1156 (N_1156,N_1123,N_1102);
and U1157 (N_1157,N_1142,N_1138);
and U1158 (N_1158,N_1100,N_1120);
and U1159 (N_1159,N_1111,N_1145);
nor U1160 (N_1160,N_1149,N_1147);
and U1161 (N_1161,N_1137,N_1126);
nor U1162 (N_1162,N_1117,N_1130);
or U1163 (N_1163,N_1104,N_1109);
nor U1164 (N_1164,N_1128,N_1113);
and U1165 (N_1165,N_1148,N_1140);
and U1166 (N_1166,N_1125,N_1134);
or U1167 (N_1167,N_1132,N_1139);
nor U1168 (N_1168,N_1105,N_1112);
nand U1169 (N_1169,N_1131,N_1106);
or U1170 (N_1170,N_1114,N_1133);
nor U1171 (N_1171,N_1144,N_1107);
nand U1172 (N_1172,N_1124,N_1143);
nor U1173 (N_1173,N_1122,N_1121);
or U1174 (N_1174,N_1103,N_1136);
nand U1175 (N_1175,N_1120,N_1129);
or U1176 (N_1176,N_1133,N_1107);
nand U1177 (N_1177,N_1123,N_1149);
and U1178 (N_1178,N_1101,N_1132);
nor U1179 (N_1179,N_1102,N_1128);
and U1180 (N_1180,N_1105,N_1113);
nor U1181 (N_1181,N_1128,N_1110);
or U1182 (N_1182,N_1117,N_1149);
and U1183 (N_1183,N_1119,N_1143);
or U1184 (N_1184,N_1115,N_1104);
and U1185 (N_1185,N_1122,N_1111);
or U1186 (N_1186,N_1115,N_1134);
nand U1187 (N_1187,N_1148,N_1109);
nand U1188 (N_1188,N_1116,N_1124);
nand U1189 (N_1189,N_1117,N_1116);
xnor U1190 (N_1190,N_1125,N_1129);
and U1191 (N_1191,N_1102,N_1117);
nor U1192 (N_1192,N_1145,N_1100);
xor U1193 (N_1193,N_1140,N_1135);
xor U1194 (N_1194,N_1103,N_1125);
or U1195 (N_1195,N_1127,N_1123);
or U1196 (N_1196,N_1140,N_1117);
nor U1197 (N_1197,N_1116,N_1106);
and U1198 (N_1198,N_1135,N_1100);
and U1199 (N_1199,N_1148,N_1102);
or U1200 (N_1200,N_1179,N_1193);
nor U1201 (N_1201,N_1191,N_1194);
nand U1202 (N_1202,N_1187,N_1171);
and U1203 (N_1203,N_1174,N_1172);
nor U1204 (N_1204,N_1180,N_1150);
xnor U1205 (N_1205,N_1157,N_1159);
nand U1206 (N_1206,N_1198,N_1168);
nand U1207 (N_1207,N_1185,N_1165);
or U1208 (N_1208,N_1184,N_1182);
nor U1209 (N_1209,N_1166,N_1152);
or U1210 (N_1210,N_1151,N_1155);
nor U1211 (N_1211,N_1186,N_1153);
or U1212 (N_1212,N_1162,N_1178);
and U1213 (N_1213,N_1161,N_1189);
nor U1214 (N_1214,N_1163,N_1199);
or U1215 (N_1215,N_1170,N_1164);
or U1216 (N_1216,N_1195,N_1176);
or U1217 (N_1217,N_1197,N_1156);
or U1218 (N_1218,N_1169,N_1175);
nor U1219 (N_1219,N_1181,N_1183);
nand U1220 (N_1220,N_1167,N_1196);
and U1221 (N_1221,N_1160,N_1192);
nor U1222 (N_1222,N_1154,N_1177);
or U1223 (N_1223,N_1188,N_1158);
and U1224 (N_1224,N_1190,N_1173);
and U1225 (N_1225,N_1192,N_1181);
and U1226 (N_1226,N_1173,N_1198);
nor U1227 (N_1227,N_1192,N_1194);
xnor U1228 (N_1228,N_1176,N_1157);
and U1229 (N_1229,N_1194,N_1157);
and U1230 (N_1230,N_1180,N_1151);
xor U1231 (N_1231,N_1183,N_1158);
nor U1232 (N_1232,N_1185,N_1199);
nor U1233 (N_1233,N_1190,N_1182);
nand U1234 (N_1234,N_1180,N_1172);
and U1235 (N_1235,N_1185,N_1189);
or U1236 (N_1236,N_1182,N_1176);
and U1237 (N_1237,N_1178,N_1168);
and U1238 (N_1238,N_1197,N_1154);
or U1239 (N_1239,N_1192,N_1186);
xnor U1240 (N_1240,N_1184,N_1179);
and U1241 (N_1241,N_1167,N_1175);
nand U1242 (N_1242,N_1172,N_1182);
nand U1243 (N_1243,N_1172,N_1151);
xor U1244 (N_1244,N_1181,N_1191);
or U1245 (N_1245,N_1162,N_1151);
or U1246 (N_1246,N_1186,N_1180);
or U1247 (N_1247,N_1172,N_1192);
and U1248 (N_1248,N_1188,N_1194);
xnor U1249 (N_1249,N_1172,N_1167);
and U1250 (N_1250,N_1220,N_1221);
nand U1251 (N_1251,N_1212,N_1214);
nor U1252 (N_1252,N_1236,N_1223);
and U1253 (N_1253,N_1232,N_1203);
nor U1254 (N_1254,N_1244,N_1226);
or U1255 (N_1255,N_1225,N_1202);
nand U1256 (N_1256,N_1207,N_1235);
nand U1257 (N_1257,N_1231,N_1229);
or U1258 (N_1258,N_1241,N_1204);
nor U1259 (N_1259,N_1245,N_1222);
xor U1260 (N_1260,N_1215,N_1242);
or U1261 (N_1261,N_1219,N_1227);
or U1262 (N_1262,N_1210,N_1217);
xnor U1263 (N_1263,N_1239,N_1243);
xnor U1264 (N_1264,N_1246,N_1208);
nor U1265 (N_1265,N_1237,N_1249);
and U1266 (N_1266,N_1218,N_1234);
nand U1267 (N_1267,N_1206,N_1248);
and U1268 (N_1268,N_1216,N_1213);
nor U1269 (N_1269,N_1230,N_1247);
xor U1270 (N_1270,N_1200,N_1209);
or U1271 (N_1271,N_1201,N_1240);
nor U1272 (N_1272,N_1205,N_1224);
or U1273 (N_1273,N_1233,N_1238);
or U1274 (N_1274,N_1211,N_1228);
nor U1275 (N_1275,N_1240,N_1230);
nor U1276 (N_1276,N_1219,N_1243);
or U1277 (N_1277,N_1234,N_1205);
nand U1278 (N_1278,N_1248,N_1225);
and U1279 (N_1279,N_1200,N_1211);
nor U1280 (N_1280,N_1218,N_1216);
nor U1281 (N_1281,N_1208,N_1245);
nand U1282 (N_1282,N_1211,N_1236);
nor U1283 (N_1283,N_1241,N_1202);
nand U1284 (N_1284,N_1215,N_1220);
and U1285 (N_1285,N_1249,N_1239);
or U1286 (N_1286,N_1239,N_1237);
or U1287 (N_1287,N_1242,N_1231);
or U1288 (N_1288,N_1239,N_1229);
and U1289 (N_1289,N_1208,N_1205);
nor U1290 (N_1290,N_1236,N_1214);
nand U1291 (N_1291,N_1225,N_1204);
xor U1292 (N_1292,N_1241,N_1225);
nor U1293 (N_1293,N_1234,N_1209);
nand U1294 (N_1294,N_1238,N_1204);
nand U1295 (N_1295,N_1240,N_1242);
nand U1296 (N_1296,N_1216,N_1235);
or U1297 (N_1297,N_1248,N_1237);
and U1298 (N_1298,N_1227,N_1230);
nor U1299 (N_1299,N_1200,N_1236);
nor U1300 (N_1300,N_1282,N_1253);
nor U1301 (N_1301,N_1291,N_1264);
or U1302 (N_1302,N_1299,N_1250);
nor U1303 (N_1303,N_1258,N_1256);
and U1304 (N_1304,N_1271,N_1274);
nand U1305 (N_1305,N_1259,N_1290);
or U1306 (N_1306,N_1263,N_1260);
or U1307 (N_1307,N_1292,N_1297);
and U1308 (N_1308,N_1279,N_1294);
nor U1309 (N_1309,N_1289,N_1296);
or U1310 (N_1310,N_1265,N_1293);
and U1311 (N_1311,N_1269,N_1277);
or U1312 (N_1312,N_1266,N_1273);
or U1313 (N_1313,N_1272,N_1251);
or U1314 (N_1314,N_1295,N_1288);
or U1315 (N_1315,N_1281,N_1287);
and U1316 (N_1316,N_1298,N_1283);
nand U1317 (N_1317,N_1276,N_1262);
and U1318 (N_1318,N_1254,N_1267);
xnor U1319 (N_1319,N_1268,N_1285);
nor U1320 (N_1320,N_1261,N_1278);
and U1321 (N_1321,N_1270,N_1275);
nor U1322 (N_1322,N_1252,N_1284);
nand U1323 (N_1323,N_1286,N_1257);
xnor U1324 (N_1324,N_1255,N_1280);
nor U1325 (N_1325,N_1287,N_1264);
or U1326 (N_1326,N_1259,N_1257);
xor U1327 (N_1327,N_1277,N_1260);
nor U1328 (N_1328,N_1295,N_1264);
or U1329 (N_1329,N_1257,N_1253);
nand U1330 (N_1330,N_1296,N_1271);
xor U1331 (N_1331,N_1293,N_1277);
nor U1332 (N_1332,N_1285,N_1288);
nand U1333 (N_1333,N_1285,N_1256);
xor U1334 (N_1334,N_1291,N_1286);
and U1335 (N_1335,N_1298,N_1282);
xor U1336 (N_1336,N_1259,N_1296);
xnor U1337 (N_1337,N_1265,N_1281);
nand U1338 (N_1338,N_1284,N_1259);
nor U1339 (N_1339,N_1276,N_1272);
or U1340 (N_1340,N_1268,N_1255);
nand U1341 (N_1341,N_1268,N_1284);
nor U1342 (N_1342,N_1255,N_1289);
and U1343 (N_1343,N_1277,N_1294);
and U1344 (N_1344,N_1284,N_1296);
or U1345 (N_1345,N_1286,N_1295);
nand U1346 (N_1346,N_1293,N_1259);
nor U1347 (N_1347,N_1289,N_1284);
nand U1348 (N_1348,N_1262,N_1294);
and U1349 (N_1349,N_1269,N_1295);
and U1350 (N_1350,N_1317,N_1340);
nand U1351 (N_1351,N_1329,N_1314);
or U1352 (N_1352,N_1347,N_1308);
xor U1353 (N_1353,N_1310,N_1306);
and U1354 (N_1354,N_1311,N_1330);
and U1355 (N_1355,N_1328,N_1349);
nand U1356 (N_1356,N_1338,N_1305);
and U1357 (N_1357,N_1326,N_1324);
nand U1358 (N_1358,N_1316,N_1331);
or U1359 (N_1359,N_1346,N_1348);
or U1360 (N_1360,N_1333,N_1300);
nor U1361 (N_1361,N_1342,N_1343);
nor U1362 (N_1362,N_1337,N_1313);
nand U1363 (N_1363,N_1319,N_1341);
or U1364 (N_1364,N_1309,N_1321);
and U1365 (N_1365,N_1336,N_1322);
xor U1366 (N_1366,N_1325,N_1315);
nor U1367 (N_1367,N_1344,N_1335);
nand U1368 (N_1368,N_1318,N_1303);
nor U1369 (N_1369,N_1304,N_1332);
or U1370 (N_1370,N_1339,N_1345);
nor U1371 (N_1371,N_1302,N_1327);
or U1372 (N_1372,N_1307,N_1323);
nor U1373 (N_1373,N_1312,N_1301);
nor U1374 (N_1374,N_1320,N_1334);
and U1375 (N_1375,N_1303,N_1342);
nor U1376 (N_1376,N_1324,N_1304);
and U1377 (N_1377,N_1327,N_1305);
nor U1378 (N_1378,N_1341,N_1343);
xnor U1379 (N_1379,N_1334,N_1311);
nand U1380 (N_1380,N_1335,N_1333);
and U1381 (N_1381,N_1340,N_1308);
xnor U1382 (N_1382,N_1308,N_1318);
xor U1383 (N_1383,N_1339,N_1311);
or U1384 (N_1384,N_1313,N_1304);
or U1385 (N_1385,N_1331,N_1319);
nor U1386 (N_1386,N_1305,N_1335);
nor U1387 (N_1387,N_1316,N_1330);
nor U1388 (N_1388,N_1332,N_1347);
nor U1389 (N_1389,N_1315,N_1346);
nand U1390 (N_1390,N_1327,N_1321);
or U1391 (N_1391,N_1314,N_1333);
and U1392 (N_1392,N_1340,N_1339);
and U1393 (N_1393,N_1341,N_1335);
nor U1394 (N_1394,N_1336,N_1301);
nand U1395 (N_1395,N_1340,N_1320);
and U1396 (N_1396,N_1303,N_1330);
nor U1397 (N_1397,N_1331,N_1321);
nor U1398 (N_1398,N_1313,N_1303);
nor U1399 (N_1399,N_1301,N_1342);
nand U1400 (N_1400,N_1392,N_1380);
nor U1401 (N_1401,N_1362,N_1384);
and U1402 (N_1402,N_1351,N_1398);
or U1403 (N_1403,N_1357,N_1393);
nor U1404 (N_1404,N_1395,N_1355);
and U1405 (N_1405,N_1369,N_1383);
or U1406 (N_1406,N_1378,N_1390);
nor U1407 (N_1407,N_1368,N_1389);
or U1408 (N_1408,N_1370,N_1394);
or U1409 (N_1409,N_1397,N_1377);
nand U1410 (N_1410,N_1374,N_1387);
or U1411 (N_1411,N_1399,N_1385);
nor U1412 (N_1412,N_1365,N_1375);
nand U1413 (N_1413,N_1360,N_1391);
and U1414 (N_1414,N_1388,N_1364);
xor U1415 (N_1415,N_1366,N_1367);
and U1416 (N_1416,N_1371,N_1352);
xor U1417 (N_1417,N_1350,N_1396);
or U1418 (N_1418,N_1356,N_1381);
nand U1419 (N_1419,N_1361,N_1376);
and U1420 (N_1420,N_1359,N_1353);
nor U1421 (N_1421,N_1354,N_1358);
nor U1422 (N_1422,N_1372,N_1386);
xor U1423 (N_1423,N_1379,N_1382);
nor U1424 (N_1424,N_1373,N_1363);
and U1425 (N_1425,N_1397,N_1372);
or U1426 (N_1426,N_1367,N_1385);
nor U1427 (N_1427,N_1375,N_1373);
or U1428 (N_1428,N_1368,N_1384);
and U1429 (N_1429,N_1363,N_1380);
nor U1430 (N_1430,N_1378,N_1395);
nand U1431 (N_1431,N_1353,N_1395);
or U1432 (N_1432,N_1359,N_1397);
xor U1433 (N_1433,N_1388,N_1395);
or U1434 (N_1434,N_1379,N_1361);
nand U1435 (N_1435,N_1398,N_1386);
nor U1436 (N_1436,N_1379,N_1356);
or U1437 (N_1437,N_1390,N_1376);
nand U1438 (N_1438,N_1391,N_1383);
xor U1439 (N_1439,N_1393,N_1368);
or U1440 (N_1440,N_1362,N_1370);
nand U1441 (N_1441,N_1357,N_1396);
xnor U1442 (N_1442,N_1399,N_1375);
and U1443 (N_1443,N_1381,N_1379);
or U1444 (N_1444,N_1379,N_1390);
and U1445 (N_1445,N_1358,N_1384);
and U1446 (N_1446,N_1354,N_1393);
nand U1447 (N_1447,N_1366,N_1385);
nor U1448 (N_1448,N_1354,N_1395);
xor U1449 (N_1449,N_1380,N_1390);
nor U1450 (N_1450,N_1430,N_1425);
and U1451 (N_1451,N_1400,N_1446);
nor U1452 (N_1452,N_1407,N_1406);
or U1453 (N_1453,N_1436,N_1423);
and U1454 (N_1454,N_1438,N_1432);
and U1455 (N_1455,N_1443,N_1427);
and U1456 (N_1456,N_1416,N_1428);
and U1457 (N_1457,N_1405,N_1431);
nand U1458 (N_1458,N_1448,N_1424);
and U1459 (N_1459,N_1415,N_1447);
xor U1460 (N_1460,N_1414,N_1419);
nand U1461 (N_1461,N_1421,N_1412);
and U1462 (N_1462,N_1437,N_1404);
or U1463 (N_1463,N_1413,N_1439);
nand U1464 (N_1464,N_1442,N_1433);
and U1465 (N_1465,N_1417,N_1449);
nand U1466 (N_1466,N_1410,N_1422);
or U1467 (N_1467,N_1403,N_1408);
nand U1468 (N_1468,N_1409,N_1441);
and U1469 (N_1469,N_1434,N_1426);
or U1470 (N_1470,N_1411,N_1402);
nor U1471 (N_1471,N_1445,N_1435);
nor U1472 (N_1472,N_1440,N_1401);
nand U1473 (N_1473,N_1429,N_1418);
and U1474 (N_1474,N_1420,N_1444);
and U1475 (N_1475,N_1432,N_1435);
nand U1476 (N_1476,N_1440,N_1412);
nand U1477 (N_1477,N_1423,N_1412);
xnor U1478 (N_1478,N_1420,N_1437);
xnor U1479 (N_1479,N_1410,N_1448);
and U1480 (N_1480,N_1416,N_1400);
or U1481 (N_1481,N_1404,N_1413);
nand U1482 (N_1482,N_1401,N_1437);
nand U1483 (N_1483,N_1438,N_1431);
nand U1484 (N_1484,N_1447,N_1404);
or U1485 (N_1485,N_1426,N_1413);
or U1486 (N_1486,N_1433,N_1448);
and U1487 (N_1487,N_1415,N_1401);
or U1488 (N_1488,N_1443,N_1447);
and U1489 (N_1489,N_1424,N_1445);
nor U1490 (N_1490,N_1414,N_1400);
nand U1491 (N_1491,N_1438,N_1434);
or U1492 (N_1492,N_1429,N_1449);
nand U1493 (N_1493,N_1425,N_1433);
nand U1494 (N_1494,N_1447,N_1435);
and U1495 (N_1495,N_1406,N_1404);
and U1496 (N_1496,N_1444,N_1416);
nor U1497 (N_1497,N_1408,N_1418);
and U1498 (N_1498,N_1446,N_1440);
nand U1499 (N_1499,N_1443,N_1401);
nor U1500 (N_1500,N_1470,N_1472);
and U1501 (N_1501,N_1495,N_1476);
nand U1502 (N_1502,N_1450,N_1454);
and U1503 (N_1503,N_1469,N_1489);
nor U1504 (N_1504,N_1460,N_1456);
nand U1505 (N_1505,N_1468,N_1467);
or U1506 (N_1506,N_1484,N_1464);
and U1507 (N_1507,N_1478,N_1466);
xnor U1508 (N_1508,N_1485,N_1498);
and U1509 (N_1509,N_1475,N_1481);
nor U1510 (N_1510,N_1483,N_1473);
or U1511 (N_1511,N_1479,N_1477);
nand U1512 (N_1512,N_1492,N_1459);
nand U1513 (N_1513,N_1493,N_1458);
xor U1514 (N_1514,N_1499,N_1463);
and U1515 (N_1515,N_1497,N_1465);
or U1516 (N_1516,N_1471,N_1451);
or U1517 (N_1517,N_1486,N_1453);
xor U1518 (N_1518,N_1452,N_1457);
and U1519 (N_1519,N_1461,N_1462);
nor U1520 (N_1520,N_1494,N_1491);
or U1521 (N_1521,N_1482,N_1480);
or U1522 (N_1522,N_1490,N_1455);
or U1523 (N_1523,N_1487,N_1474);
nand U1524 (N_1524,N_1496,N_1488);
nor U1525 (N_1525,N_1481,N_1485);
and U1526 (N_1526,N_1487,N_1494);
nor U1527 (N_1527,N_1472,N_1478);
nand U1528 (N_1528,N_1486,N_1455);
and U1529 (N_1529,N_1459,N_1463);
nor U1530 (N_1530,N_1464,N_1483);
and U1531 (N_1531,N_1484,N_1482);
nor U1532 (N_1532,N_1452,N_1456);
or U1533 (N_1533,N_1474,N_1468);
xnor U1534 (N_1534,N_1494,N_1479);
nor U1535 (N_1535,N_1454,N_1459);
or U1536 (N_1536,N_1493,N_1481);
and U1537 (N_1537,N_1495,N_1460);
or U1538 (N_1538,N_1459,N_1494);
nand U1539 (N_1539,N_1454,N_1455);
or U1540 (N_1540,N_1499,N_1457);
nor U1541 (N_1541,N_1463,N_1490);
nand U1542 (N_1542,N_1458,N_1470);
and U1543 (N_1543,N_1477,N_1460);
xnor U1544 (N_1544,N_1476,N_1482);
or U1545 (N_1545,N_1466,N_1475);
nand U1546 (N_1546,N_1472,N_1466);
and U1547 (N_1547,N_1486,N_1461);
nor U1548 (N_1548,N_1473,N_1452);
or U1549 (N_1549,N_1489,N_1495);
nand U1550 (N_1550,N_1518,N_1549);
or U1551 (N_1551,N_1502,N_1519);
and U1552 (N_1552,N_1540,N_1539);
nor U1553 (N_1553,N_1528,N_1501);
and U1554 (N_1554,N_1531,N_1545);
nand U1555 (N_1555,N_1511,N_1505);
or U1556 (N_1556,N_1509,N_1547);
nor U1557 (N_1557,N_1533,N_1513);
nor U1558 (N_1558,N_1548,N_1517);
nor U1559 (N_1559,N_1514,N_1507);
or U1560 (N_1560,N_1535,N_1544);
or U1561 (N_1561,N_1512,N_1532);
or U1562 (N_1562,N_1536,N_1530);
nand U1563 (N_1563,N_1534,N_1515);
and U1564 (N_1564,N_1522,N_1541);
or U1565 (N_1565,N_1529,N_1503);
and U1566 (N_1566,N_1523,N_1526);
xnor U1567 (N_1567,N_1524,N_1506);
or U1568 (N_1568,N_1510,N_1500);
and U1569 (N_1569,N_1504,N_1508);
nor U1570 (N_1570,N_1525,N_1520);
nand U1571 (N_1571,N_1516,N_1543);
and U1572 (N_1572,N_1527,N_1521);
nand U1573 (N_1573,N_1546,N_1537);
nand U1574 (N_1574,N_1542,N_1538);
nor U1575 (N_1575,N_1512,N_1540);
nor U1576 (N_1576,N_1533,N_1543);
nor U1577 (N_1577,N_1534,N_1548);
nand U1578 (N_1578,N_1539,N_1513);
and U1579 (N_1579,N_1509,N_1518);
nor U1580 (N_1580,N_1542,N_1501);
xnor U1581 (N_1581,N_1535,N_1531);
or U1582 (N_1582,N_1512,N_1534);
nor U1583 (N_1583,N_1531,N_1536);
nand U1584 (N_1584,N_1526,N_1536);
or U1585 (N_1585,N_1511,N_1536);
and U1586 (N_1586,N_1509,N_1513);
or U1587 (N_1587,N_1517,N_1528);
or U1588 (N_1588,N_1514,N_1528);
nor U1589 (N_1589,N_1535,N_1539);
nand U1590 (N_1590,N_1511,N_1546);
or U1591 (N_1591,N_1516,N_1510);
nor U1592 (N_1592,N_1502,N_1505);
nor U1593 (N_1593,N_1526,N_1515);
nor U1594 (N_1594,N_1544,N_1501);
nor U1595 (N_1595,N_1532,N_1546);
nor U1596 (N_1596,N_1508,N_1524);
nand U1597 (N_1597,N_1526,N_1530);
or U1598 (N_1598,N_1505,N_1517);
xnor U1599 (N_1599,N_1538,N_1548);
or U1600 (N_1600,N_1577,N_1583);
and U1601 (N_1601,N_1560,N_1552);
or U1602 (N_1602,N_1571,N_1585);
nand U1603 (N_1603,N_1596,N_1557);
nand U1604 (N_1604,N_1584,N_1597);
nor U1605 (N_1605,N_1593,N_1569);
or U1606 (N_1606,N_1574,N_1587);
nor U1607 (N_1607,N_1565,N_1550);
nand U1608 (N_1608,N_1568,N_1586);
and U1609 (N_1609,N_1599,N_1561);
and U1610 (N_1610,N_1595,N_1562);
and U1611 (N_1611,N_1575,N_1564);
nand U1612 (N_1612,N_1556,N_1559);
or U1613 (N_1613,N_1581,N_1572);
nor U1614 (N_1614,N_1576,N_1580);
or U1615 (N_1615,N_1589,N_1598);
and U1616 (N_1616,N_1563,N_1555);
and U1617 (N_1617,N_1553,N_1551);
and U1618 (N_1618,N_1591,N_1566);
and U1619 (N_1619,N_1558,N_1594);
nand U1620 (N_1620,N_1578,N_1588);
and U1621 (N_1621,N_1579,N_1570);
nor U1622 (N_1622,N_1582,N_1590);
nor U1623 (N_1623,N_1592,N_1567);
or U1624 (N_1624,N_1554,N_1573);
xnor U1625 (N_1625,N_1597,N_1589);
xnor U1626 (N_1626,N_1574,N_1592);
nor U1627 (N_1627,N_1568,N_1550);
or U1628 (N_1628,N_1573,N_1593);
and U1629 (N_1629,N_1562,N_1574);
nand U1630 (N_1630,N_1598,N_1573);
nand U1631 (N_1631,N_1578,N_1568);
nand U1632 (N_1632,N_1564,N_1585);
nand U1633 (N_1633,N_1591,N_1582);
or U1634 (N_1634,N_1564,N_1557);
xor U1635 (N_1635,N_1563,N_1589);
nand U1636 (N_1636,N_1561,N_1566);
or U1637 (N_1637,N_1599,N_1580);
and U1638 (N_1638,N_1571,N_1587);
or U1639 (N_1639,N_1558,N_1572);
nor U1640 (N_1640,N_1556,N_1571);
or U1641 (N_1641,N_1553,N_1583);
nor U1642 (N_1642,N_1552,N_1591);
or U1643 (N_1643,N_1557,N_1554);
or U1644 (N_1644,N_1580,N_1569);
nor U1645 (N_1645,N_1569,N_1596);
nor U1646 (N_1646,N_1576,N_1594);
nand U1647 (N_1647,N_1590,N_1556);
nor U1648 (N_1648,N_1560,N_1569);
nand U1649 (N_1649,N_1574,N_1568);
and U1650 (N_1650,N_1602,N_1605);
xor U1651 (N_1651,N_1642,N_1620);
nand U1652 (N_1652,N_1608,N_1626);
and U1653 (N_1653,N_1629,N_1625);
and U1654 (N_1654,N_1606,N_1600);
nor U1655 (N_1655,N_1636,N_1648);
nand U1656 (N_1656,N_1641,N_1639);
or U1657 (N_1657,N_1638,N_1627);
or U1658 (N_1658,N_1617,N_1618);
and U1659 (N_1659,N_1644,N_1622);
nor U1660 (N_1660,N_1616,N_1647);
nand U1661 (N_1661,N_1635,N_1645);
or U1662 (N_1662,N_1604,N_1619);
and U1663 (N_1663,N_1610,N_1632);
and U1664 (N_1664,N_1646,N_1603);
nand U1665 (N_1665,N_1615,N_1640);
xnor U1666 (N_1666,N_1609,N_1601);
or U1667 (N_1667,N_1607,N_1611);
nor U1668 (N_1668,N_1613,N_1624);
and U1669 (N_1669,N_1634,N_1612);
nor U1670 (N_1670,N_1628,N_1623);
nand U1671 (N_1671,N_1614,N_1621);
xor U1672 (N_1672,N_1630,N_1631);
nand U1673 (N_1673,N_1633,N_1643);
nand U1674 (N_1674,N_1649,N_1637);
nor U1675 (N_1675,N_1631,N_1639);
and U1676 (N_1676,N_1625,N_1603);
xnor U1677 (N_1677,N_1606,N_1603);
or U1678 (N_1678,N_1607,N_1608);
and U1679 (N_1679,N_1610,N_1602);
or U1680 (N_1680,N_1632,N_1603);
nor U1681 (N_1681,N_1601,N_1630);
nor U1682 (N_1682,N_1632,N_1628);
and U1683 (N_1683,N_1602,N_1636);
xor U1684 (N_1684,N_1606,N_1637);
or U1685 (N_1685,N_1619,N_1600);
nand U1686 (N_1686,N_1636,N_1644);
or U1687 (N_1687,N_1611,N_1602);
nor U1688 (N_1688,N_1600,N_1628);
nor U1689 (N_1689,N_1629,N_1618);
nor U1690 (N_1690,N_1633,N_1612);
nor U1691 (N_1691,N_1616,N_1632);
xor U1692 (N_1692,N_1649,N_1646);
or U1693 (N_1693,N_1606,N_1649);
nor U1694 (N_1694,N_1601,N_1613);
and U1695 (N_1695,N_1634,N_1622);
and U1696 (N_1696,N_1609,N_1616);
nand U1697 (N_1697,N_1604,N_1643);
and U1698 (N_1698,N_1619,N_1615);
or U1699 (N_1699,N_1617,N_1636);
and U1700 (N_1700,N_1699,N_1682);
nor U1701 (N_1701,N_1657,N_1686);
nand U1702 (N_1702,N_1690,N_1674);
xnor U1703 (N_1703,N_1652,N_1656);
or U1704 (N_1704,N_1650,N_1663);
nor U1705 (N_1705,N_1664,N_1684);
nor U1706 (N_1706,N_1658,N_1683);
and U1707 (N_1707,N_1692,N_1668);
and U1708 (N_1708,N_1655,N_1680);
xor U1709 (N_1709,N_1676,N_1681);
nand U1710 (N_1710,N_1698,N_1677);
and U1711 (N_1711,N_1688,N_1661);
xnor U1712 (N_1712,N_1672,N_1697);
xor U1713 (N_1713,N_1685,N_1670);
nor U1714 (N_1714,N_1679,N_1675);
and U1715 (N_1715,N_1689,N_1667);
nor U1716 (N_1716,N_1654,N_1695);
nand U1717 (N_1717,N_1651,N_1665);
and U1718 (N_1718,N_1678,N_1659);
or U1719 (N_1719,N_1673,N_1687);
nor U1720 (N_1720,N_1669,N_1671);
or U1721 (N_1721,N_1696,N_1694);
nand U1722 (N_1722,N_1691,N_1666);
or U1723 (N_1723,N_1662,N_1693);
nor U1724 (N_1724,N_1660,N_1653);
nor U1725 (N_1725,N_1668,N_1665);
nand U1726 (N_1726,N_1661,N_1693);
and U1727 (N_1727,N_1658,N_1655);
nor U1728 (N_1728,N_1694,N_1673);
nor U1729 (N_1729,N_1663,N_1683);
and U1730 (N_1730,N_1654,N_1681);
and U1731 (N_1731,N_1673,N_1684);
nand U1732 (N_1732,N_1666,N_1670);
and U1733 (N_1733,N_1695,N_1662);
nand U1734 (N_1734,N_1668,N_1679);
nor U1735 (N_1735,N_1654,N_1671);
and U1736 (N_1736,N_1674,N_1688);
nand U1737 (N_1737,N_1656,N_1699);
and U1738 (N_1738,N_1657,N_1698);
nand U1739 (N_1739,N_1676,N_1693);
nand U1740 (N_1740,N_1693,N_1652);
nor U1741 (N_1741,N_1679,N_1653);
nand U1742 (N_1742,N_1699,N_1693);
nor U1743 (N_1743,N_1677,N_1693);
xnor U1744 (N_1744,N_1671,N_1678);
xor U1745 (N_1745,N_1688,N_1673);
and U1746 (N_1746,N_1686,N_1683);
nand U1747 (N_1747,N_1697,N_1666);
nor U1748 (N_1748,N_1661,N_1678);
or U1749 (N_1749,N_1673,N_1677);
nor U1750 (N_1750,N_1706,N_1716);
and U1751 (N_1751,N_1717,N_1744);
xnor U1752 (N_1752,N_1721,N_1748);
nor U1753 (N_1753,N_1726,N_1745);
xor U1754 (N_1754,N_1723,N_1747);
and U1755 (N_1755,N_1733,N_1705);
nor U1756 (N_1756,N_1708,N_1743);
xnor U1757 (N_1757,N_1739,N_1738);
nand U1758 (N_1758,N_1735,N_1711);
nand U1759 (N_1759,N_1727,N_1720);
xnor U1760 (N_1760,N_1730,N_1724);
nand U1761 (N_1761,N_1703,N_1707);
and U1762 (N_1762,N_1700,N_1712);
nand U1763 (N_1763,N_1725,N_1702);
nand U1764 (N_1764,N_1715,N_1731);
or U1765 (N_1765,N_1732,N_1722);
nand U1766 (N_1766,N_1728,N_1737);
nor U1767 (N_1767,N_1741,N_1704);
nand U1768 (N_1768,N_1719,N_1742);
nor U1769 (N_1769,N_1710,N_1709);
xor U1770 (N_1770,N_1718,N_1736);
or U1771 (N_1771,N_1714,N_1701);
and U1772 (N_1772,N_1746,N_1713);
xnor U1773 (N_1773,N_1740,N_1729);
xnor U1774 (N_1774,N_1749,N_1734);
or U1775 (N_1775,N_1701,N_1734);
or U1776 (N_1776,N_1722,N_1713);
or U1777 (N_1777,N_1718,N_1746);
nor U1778 (N_1778,N_1748,N_1744);
nand U1779 (N_1779,N_1729,N_1718);
nand U1780 (N_1780,N_1724,N_1705);
or U1781 (N_1781,N_1724,N_1721);
xor U1782 (N_1782,N_1737,N_1710);
nand U1783 (N_1783,N_1727,N_1706);
or U1784 (N_1784,N_1714,N_1729);
nor U1785 (N_1785,N_1737,N_1744);
nand U1786 (N_1786,N_1736,N_1728);
xor U1787 (N_1787,N_1724,N_1739);
nand U1788 (N_1788,N_1732,N_1723);
nor U1789 (N_1789,N_1718,N_1703);
and U1790 (N_1790,N_1706,N_1712);
or U1791 (N_1791,N_1704,N_1731);
nor U1792 (N_1792,N_1701,N_1710);
or U1793 (N_1793,N_1734,N_1711);
nand U1794 (N_1794,N_1702,N_1749);
nand U1795 (N_1795,N_1707,N_1701);
and U1796 (N_1796,N_1744,N_1742);
nor U1797 (N_1797,N_1703,N_1744);
nor U1798 (N_1798,N_1744,N_1727);
nand U1799 (N_1799,N_1706,N_1717);
nand U1800 (N_1800,N_1765,N_1752);
nor U1801 (N_1801,N_1766,N_1770);
or U1802 (N_1802,N_1779,N_1789);
nand U1803 (N_1803,N_1771,N_1776);
nor U1804 (N_1804,N_1788,N_1782);
or U1805 (N_1805,N_1755,N_1790);
or U1806 (N_1806,N_1778,N_1769);
and U1807 (N_1807,N_1768,N_1775);
xor U1808 (N_1808,N_1781,N_1757);
or U1809 (N_1809,N_1794,N_1774);
nor U1810 (N_1810,N_1750,N_1759);
and U1811 (N_1811,N_1763,N_1756);
nor U1812 (N_1812,N_1758,N_1761);
xnor U1813 (N_1813,N_1796,N_1783);
nor U1814 (N_1814,N_1797,N_1795);
and U1815 (N_1815,N_1754,N_1786);
and U1816 (N_1816,N_1777,N_1780);
or U1817 (N_1817,N_1751,N_1787);
xnor U1818 (N_1818,N_1762,N_1792);
nand U1819 (N_1819,N_1767,N_1760);
and U1820 (N_1820,N_1791,N_1785);
or U1821 (N_1821,N_1793,N_1773);
nand U1822 (N_1822,N_1772,N_1753);
or U1823 (N_1823,N_1784,N_1764);
nand U1824 (N_1824,N_1798,N_1799);
and U1825 (N_1825,N_1751,N_1754);
nor U1826 (N_1826,N_1754,N_1768);
nand U1827 (N_1827,N_1759,N_1768);
and U1828 (N_1828,N_1784,N_1797);
nor U1829 (N_1829,N_1793,N_1756);
and U1830 (N_1830,N_1771,N_1798);
nor U1831 (N_1831,N_1771,N_1778);
nand U1832 (N_1832,N_1779,N_1754);
nor U1833 (N_1833,N_1751,N_1770);
xor U1834 (N_1834,N_1790,N_1773);
nand U1835 (N_1835,N_1778,N_1752);
or U1836 (N_1836,N_1756,N_1753);
nor U1837 (N_1837,N_1795,N_1788);
and U1838 (N_1838,N_1777,N_1799);
and U1839 (N_1839,N_1786,N_1789);
or U1840 (N_1840,N_1763,N_1783);
nand U1841 (N_1841,N_1784,N_1786);
or U1842 (N_1842,N_1761,N_1759);
or U1843 (N_1843,N_1776,N_1787);
and U1844 (N_1844,N_1765,N_1791);
xor U1845 (N_1845,N_1759,N_1765);
or U1846 (N_1846,N_1766,N_1779);
or U1847 (N_1847,N_1756,N_1760);
xnor U1848 (N_1848,N_1782,N_1771);
or U1849 (N_1849,N_1774,N_1784);
xnor U1850 (N_1850,N_1833,N_1806);
nand U1851 (N_1851,N_1825,N_1827);
nor U1852 (N_1852,N_1818,N_1823);
nor U1853 (N_1853,N_1800,N_1822);
xnor U1854 (N_1854,N_1834,N_1832);
nand U1855 (N_1855,N_1847,N_1807);
and U1856 (N_1856,N_1802,N_1826);
nand U1857 (N_1857,N_1840,N_1842);
nor U1858 (N_1858,N_1805,N_1846);
or U1859 (N_1859,N_1815,N_1814);
or U1860 (N_1860,N_1819,N_1816);
nor U1861 (N_1861,N_1836,N_1824);
or U1862 (N_1862,N_1811,N_1830);
or U1863 (N_1863,N_1844,N_1808);
nand U1864 (N_1864,N_1801,N_1838);
xnor U1865 (N_1865,N_1845,N_1841);
nor U1866 (N_1866,N_1803,N_1829);
or U1867 (N_1867,N_1835,N_1849);
nor U1868 (N_1868,N_1831,N_1843);
nor U1869 (N_1869,N_1848,N_1809);
nand U1870 (N_1870,N_1817,N_1804);
and U1871 (N_1871,N_1839,N_1820);
and U1872 (N_1872,N_1812,N_1837);
nor U1873 (N_1873,N_1810,N_1821);
and U1874 (N_1874,N_1813,N_1828);
and U1875 (N_1875,N_1812,N_1818);
nand U1876 (N_1876,N_1801,N_1849);
nand U1877 (N_1877,N_1810,N_1834);
or U1878 (N_1878,N_1847,N_1817);
xnor U1879 (N_1879,N_1845,N_1840);
nand U1880 (N_1880,N_1844,N_1806);
nor U1881 (N_1881,N_1812,N_1833);
nand U1882 (N_1882,N_1831,N_1839);
nand U1883 (N_1883,N_1831,N_1828);
nand U1884 (N_1884,N_1808,N_1801);
and U1885 (N_1885,N_1805,N_1822);
nand U1886 (N_1886,N_1811,N_1806);
nor U1887 (N_1887,N_1845,N_1800);
nand U1888 (N_1888,N_1834,N_1820);
nor U1889 (N_1889,N_1816,N_1803);
nand U1890 (N_1890,N_1813,N_1832);
nor U1891 (N_1891,N_1828,N_1829);
nand U1892 (N_1892,N_1817,N_1838);
or U1893 (N_1893,N_1848,N_1818);
nand U1894 (N_1894,N_1841,N_1800);
or U1895 (N_1895,N_1807,N_1837);
nand U1896 (N_1896,N_1845,N_1843);
nand U1897 (N_1897,N_1812,N_1802);
nor U1898 (N_1898,N_1802,N_1813);
nor U1899 (N_1899,N_1820,N_1849);
xor U1900 (N_1900,N_1888,N_1861);
or U1901 (N_1901,N_1865,N_1858);
nor U1902 (N_1902,N_1885,N_1879);
and U1903 (N_1903,N_1891,N_1896);
and U1904 (N_1904,N_1869,N_1875);
nor U1905 (N_1905,N_1876,N_1872);
and U1906 (N_1906,N_1857,N_1852);
nor U1907 (N_1907,N_1894,N_1889);
xnor U1908 (N_1908,N_1851,N_1893);
nand U1909 (N_1909,N_1866,N_1898);
and U1910 (N_1910,N_1863,N_1868);
nand U1911 (N_1911,N_1856,N_1862);
nand U1912 (N_1912,N_1874,N_1883);
nand U1913 (N_1913,N_1853,N_1895);
nor U1914 (N_1914,N_1871,N_1890);
or U1915 (N_1915,N_1887,N_1873);
or U1916 (N_1916,N_1867,N_1850);
nand U1917 (N_1917,N_1880,N_1854);
or U1918 (N_1918,N_1884,N_1864);
and U1919 (N_1919,N_1878,N_1892);
and U1920 (N_1920,N_1886,N_1877);
xnor U1921 (N_1921,N_1882,N_1899);
or U1922 (N_1922,N_1870,N_1855);
and U1923 (N_1923,N_1859,N_1881);
nand U1924 (N_1924,N_1860,N_1897);
xor U1925 (N_1925,N_1878,N_1855);
nand U1926 (N_1926,N_1884,N_1863);
or U1927 (N_1927,N_1872,N_1865);
xor U1928 (N_1928,N_1875,N_1894);
nor U1929 (N_1929,N_1877,N_1896);
xor U1930 (N_1930,N_1872,N_1883);
xor U1931 (N_1931,N_1887,N_1860);
or U1932 (N_1932,N_1872,N_1857);
and U1933 (N_1933,N_1885,N_1876);
nor U1934 (N_1934,N_1853,N_1856);
or U1935 (N_1935,N_1883,N_1871);
nor U1936 (N_1936,N_1878,N_1890);
nand U1937 (N_1937,N_1894,N_1890);
or U1938 (N_1938,N_1877,N_1858);
or U1939 (N_1939,N_1874,N_1890);
and U1940 (N_1940,N_1875,N_1866);
or U1941 (N_1941,N_1895,N_1899);
or U1942 (N_1942,N_1862,N_1876);
and U1943 (N_1943,N_1857,N_1869);
nand U1944 (N_1944,N_1852,N_1875);
nand U1945 (N_1945,N_1876,N_1889);
or U1946 (N_1946,N_1879,N_1861);
nand U1947 (N_1947,N_1877,N_1885);
and U1948 (N_1948,N_1878,N_1874);
xor U1949 (N_1949,N_1864,N_1850);
nor U1950 (N_1950,N_1944,N_1946);
and U1951 (N_1951,N_1909,N_1903);
nand U1952 (N_1952,N_1929,N_1948);
nand U1953 (N_1953,N_1921,N_1925);
or U1954 (N_1954,N_1933,N_1927);
nor U1955 (N_1955,N_1926,N_1914);
nor U1956 (N_1956,N_1937,N_1924);
nand U1957 (N_1957,N_1932,N_1913);
and U1958 (N_1958,N_1906,N_1912);
and U1959 (N_1959,N_1916,N_1934);
nor U1960 (N_1960,N_1940,N_1900);
nor U1961 (N_1961,N_1908,N_1939);
xnor U1962 (N_1962,N_1935,N_1936);
or U1963 (N_1963,N_1947,N_1942);
nand U1964 (N_1964,N_1905,N_1923);
or U1965 (N_1965,N_1910,N_1930);
nor U1966 (N_1966,N_1917,N_1928);
and U1967 (N_1967,N_1901,N_1943);
or U1968 (N_1968,N_1931,N_1949);
nor U1969 (N_1969,N_1922,N_1920);
or U1970 (N_1970,N_1902,N_1941);
or U1971 (N_1971,N_1918,N_1919);
and U1972 (N_1972,N_1945,N_1904);
and U1973 (N_1973,N_1907,N_1915);
xor U1974 (N_1974,N_1911,N_1938);
and U1975 (N_1975,N_1943,N_1930);
xor U1976 (N_1976,N_1923,N_1940);
nor U1977 (N_1977,N_1903,N_1935);
and U1978 (N_1978,N_1936,N_1903);
and U1979 (N_1979,N_1904,N_1918);
and U1980 (N_1980,N_1946,N_1945);
or U1981 (N_1981,N_1948,N_1921);
and U1982 (N_1982,N_1921,N_1938);
or U1983 (N_1983,N_1943,N_1925);
nand U1984 (N_1984,N_1934,N_1941);
or U1985 (N_1985,N_1946,N_1940);
nand U1986 (N_1986,N_1916,N_1908);
or U1987 (N_1987,N_1914,N_1939);
xor U1988 (N_1988,N_1924,N_1916);
nor U1989 (N_1989,N_1948,N_1919);
nor U1990 (N_1990,N_1913,N_1912);
nor U1991 (N_1991,N_1948,N_1939);
nand U1992 (N_1992,N_1930,N_1909);
or U1993 (N_1993,N_1940,N_1942);
or U1994 (N_1994,N_1909,N_1907);
and U1995 (N_1995,N_1942,N_1909);
and U1996 (N_1996,N_1916,N_1932);
or U1997 (N_1997,N_1919,N_1935);
and U1998 (N_1998,N_1915,N_1905);
and U1999 (N_1999,N_1910,N_1920);
nor U2000 (N_2000,N_1997,N_1971);
nand U2001 (N_2001,N_1978,N_1994);
nand U2002 (N_2002,N_1962,N_1973);
or U2003 (N_2003,N_1960,N_1972);
xor U2004 (N_2004,N_1999,N_1979);
nor U2005 (N_2005,N_1958,N_1996);
nand U2006 (N_2006,N_1963,N_1970);
or U2007 (N_2007,N_1956,N_1953);
xor U2008 (N_2008,N_1954,N_1952);
or U2009 (N_2009,N_1966,N_1969);
nor U2010 (N_2010,N_1998,N_1959);
nor U2011 (N_2011,N_1989,N_1983);
nand U2012 (N_2012,N_1988,N_1995);
xor U2013 (N_2013,N_1986,N_1982);
and U2014 (N_2014,N_1984,N_1964);
xnor U2015 (N_2015,N_1981,N_1967);
nor U2016 (N_2016,N_1961,N_1990);
and U2017 (N_2017,N_1951,N_1957);
or U2018 (N_2018,N_1965,N_1991);
or U2019 (N_2019,N_1955,N_1975);
and U2020 (N_2020,N_1974,N_1985);
or U2021 (N_2021,N_1980,N_1968);
nand U2022 (N_2022,N_1976,N_1977);
and U2023 (N_2023,N_1993,N_1992);
and U2024 (N_2024,N_1987,N_1950);
and U2025 (N_2025,N_1989,N_1952);
or U2026 (N_2026,N_1998,N_1957);
nor U2027 (N_2027,N_1956,N_1957);
or U2028 (N_2028,N_1975,N_1994);
nand U2029 (N_2029,N_1966,N_1990);
or U2030 (N_2030,N_1980,N_1999);
and U2031 (N_2031,N_1958,N_1995);
nor U2032 (N_2032,N_1993,N_1991);
nor U2033 (N_2033,N_1964,N_1975);
xnor U2034 (N_2034,N_1991,N_1953);
nand U2035 (N_2035,N_1950,N_1994);
and U2036 (N_2036,N_1968,N_1979);
and U2037 (N_2037,N_1998,N_1973);
nand U2038 (N_2038,N_1952,N_1985);
nand U2039 (N_2039,N_1987,N_1964);
or U2040 (N_2040,N_1995,N_1991);
nor U2041 (N_2041,N_1997,N_1993);
and U2042 (N_2042,N_1974,N_1986);
nor U2043 (N_2043,N_1998,N_1960);
nor U2044 (N_2044,N_1980,N_1960);
nor U2045 (N_2045,N_1995,N_1983);
and U2046 (N_2046,N_1963,N_1983);
nand U2047 (N_2047,N_1960,N_1992);
and U2048 (N_2048,N_1969,N_1956);
nand U2049 (N_2049,N_1978,N_1992);
nand U2050 (N_2050,N_2033,N_2016);
and U2051 (N_2051,N_2018,N_2046);
and U2052 (N_2052,N_2019,N_2036);
and U2053 (N_2053,N_2038,N_2039);
and U2054 (N_2054,N_2049,N_2001);
nor U2055 (N_2055,N_2034,N_2042);
nor U2056 (N_2056,N_2043,N_2022);
or U2057 (N_2057,N_2021,N_2040);
nor U2058 (N_2058,N_2023,N_2047);
nor U2059 (N_2059,N_2029,N_2011);
nand U2060 (N_2060,N_2028,N_2037);
nor U2061 (N_2061,N_2044,N_2013);
and U2062 (N_2062,N_2035,N_2008);
nand U2063 (N_2063,N_2010,N_2017);
and U2064 (N_2064,N_2014,N_2004);
nand U2065 (N_2065,N_2002,N_2020);
or U2066 (N_2066,N_2045,N_2030);
xor U2067 (N_2067,N_2025,N_2027);
nand U2068 (N_2068,N_2003,N_2048);
nand U2069 (N_2069,N_2012,N_2006);
and U2070 (N_2070,N_2009,N_2026);
nand U2071 (N_2071,N_2041,N_2015);
nand U2072 (N_2072,N_2032,N_2031);
and U2073 (N_2073,N_2024,N_2005);
or U2074 (N_2074,N_2007,N_2000);
nor U2075 (N_2075,N_2027,N_2011);
xor U2076 (N_2076,N_2001,N_2047);
or U2077 (N_2077,N_2030,N_2022);
nor U2078 (N_2078,N_2035,N_2021);
or U2079 (N_2079,N_2048,N_2017);
nor U2080 (N_2080,N_2031,N_2015);
nand U2081 (N_2081,N_2044,N_2025);
or U2082 (N_2082,N_2025,N_2039);
nor U2083 (N_2083,N_2013,N_2008);
or U2084 (N_2084,N_2049,N_2038);
nand U2085 (N_2085,N_2040,N_2024);
nor U2086 (N_2086,N_2041,N_2049);
or U2087 (N_2087,N_2006,N_2023);
and U2088 (N_2088,N_2017,N_2049);
or U2089 (N_2089,N_2038,N_2013);
nand U2090 (N_2090,N_2019,N_2041);
nand U2091 (N_2091,N_2020,N_2019);
xor U2092 (N_2092,N_2034,N_2044);
nand U2093 (N_2093,N_2017,N_2001);
and U2094 (N_2094,N_2032,N_2012);
nor U2095 (N_2095,N_2044,N_2035);
nor U2096 (N_2096,N_2025,N_2040);
nand U2097 (N_2097,N_2042,N_2037);
or U2098 (N_2098,N_2010,N_2015);
and U2099 (N_2099,N_2040,N_2011);
and U2100 (N_2100,N_2097,N_2053);
nand U2101 (N_2101,N_2057,N_2098);
or U2102 (N_2102,N_2071,N_2070);
or U2103 (N_2103,N_2077,N_2092);
nor U2104 (N_2104,N_2054,N_2081);
or U2105 (N_2105,N_2055,N_2066);
and U2106 (N_2106,N_2052,N_2079);
or U2107 (N_2107,N_2089,N_2099);
nor U2108 (N_2108,N_2069,N_2056);
nor U2109 (N_2109,N_2060,N_2067);
xor U2110 (N_2110,N_2075,N_2062);
nand U2111 (N_2111,N_2064,N_2084);
nand U2112 (N_2112,N_2065,N_2063);
nor U2113 (N_2113,N_2090,N_2080);
and U2114 (N_2114,N_2087,N_2073);
and U2115 (N_2115,N_2078,N_2076);
xor U2116 (N_2116,N_2072,N_2050);
xor U2117 (N_2117,N_2093,N_2095);
and U2118 (N_2118,N_2096,N_2086);
nand U2119 (N_2119,N_2068,N_2088);
nand U2120 (N_2120,N_2082,N_2061);
nand U2121 (N_2121,N_2058,N_2085);
and U2122 (N_2122,N_2074,N_2051);
nand U2123 (N_2123,N_2059,N_2091);
nor U2124 (N_2124,N_2094,N_2083);
and U2125 (N_2125,N_2094,N_2062);
nor U2126 (N_2126,N_2091,N_2058);
and U2127 (N_2127,N_2093,N_2067);
nor U2128 (N_2128,N_2072,N_2095);
nor U2129 (N_2129,N_2053,N_2084);
or U2130 (N_2130,N_2096,N_2062);
or U2131 (N_2131,N_2071,N_2068);
nand U2132 (N_2132,N_2080,N_2055);
or U2133 (N_2133,N_2092,N_2073);
nand U2134 (N_2134,N_2063,N_2087);
nand U2135 (N_2135,N_2059,N_2089);
nor U2136 (N_2136,N_2079,N_2050);
nand U2137 (N_2137,N_2065,N_2072);
nand U2138 (N_2138,N_2085,N_2089);
and U2139 (N_2139,N_2073,N_2065);
xor U2140 (N_2140,N_2068,N_2084);
and U2141 (N_2141,N_2068,N_2085);
nand U2142 (N_2142,N_2068,N_2099);
nor U2143 (N_2143,N_2077,N_2080);
or U2144 (N_2144,N_2082,N_2098);
or U2145 (N_2145,N_2095,N_2076);
or U2146 (N_2146,N_2070,N_2097);
or U2147 (N_2147,N_2071,N_2067);
and U2148 (N_2148,N_2082,N_2067);
nand U2149 (N_2149,N_2079,N_2051);
nor U2150 (N_2150,N_2141,N_2134);
or U2151 (N_2151,N_2125,N_2130);
nor U2152 (N_2152,N_2102,N_2111);
or U2153 (N_2153,N_2139,N_2118);
and U2154 (N_2154,N_2140,N_2136);
or U2155 (N_2155,N_2143,N_2137);
nand U2156 (N_2156,N_2114,N_2132);
nand U2157 (N_2157,N_2145,N_2128);
and U2158 (N_2158,N_2124,N_2105);
or U2159 (N_2159,N_2104,N_2110);
and U2160 (N_2160,N_2101,N_2116);
nand U2161 (N_2161,N_2113,N_2115);
xor U2162 (N_2162,N_2109,N_2144);
or U2163 (N_2163,N_2149,N_2106);
or U2164 (N_2164,N_2142,N_2117);
nor U2165 (N_2165,N_2107,N_2108);
or U2166 (N_2166,N_2147,N_2120);
nand U2167 (N_2167,N_2119,N_2112);
or U2168 (N_2168,N_2123,N_2121);
nor U2169 (N_2169,N_2138,N_2127);
or U2170 (N_2170,N_2131,N_2129);
nor U2171 (N_2171,N_2126,N_2103);
and U2172 (N_2172,N_2122,N_2148);
xnor U2173 (N_2173,N_2133,N_2146);
and U2174 (N_2174,N_2135,N_2100);
or U2175 (N_2175,N_2145,N_2141);
xor U2176 (N_2176,N_2107,N_2116);
nor U2177 (N_2177,N_2109,N_2102);
nor U2178 (N_2178,N_2120,N_2104);
nor U2179 (N_2179,N_2130,N_2148);
and U2180 (N_2180,N_2148,N_2137);
and U2181 (N_2181,N_2143,N_2136);
and U2182 (N_2182,N_2129,N_2147);
and U2183 (N_2183,N_2120,N_2142);
xor U2184 (N_2184,N_2142,N_2138);
nand U2185 (N_2185,N_2135,N_2129);
nor U2186 (N_2186,N_2149,N_2143);
and U2187 (N_2187,N_2110,N_2147);
or U2188 (N_2188,N_2149,N_2115);
and U2189 (N_2189,N_2146,N_2126);
and U2190 (N_2190,N_2115,N_2117);
nor U2191 (N_2191,N_2141,N_2105);
or U2192 (N_2192,N_2144,N_2107);
or U2193 (N_2193,N_2137,N_2119);
and U2194 (N_2194,N_2147,N_2123);
or U2195 (N_2195,N_2109,N_2114);
or U2196 (N_2196,N_2135,N_2142);
nand U2197 (N_2197,N_2104,N_2102);
nor U2198 (N_2198,N_2106,N_2137);
and U2199 (N_2199,N_2147,N_2131);
and U2200 (N_2200,N_2170,N_2176);
nor U2201 (N_2201,N_2169,N_2193);
xnor U2202 (N_2202,N_2175,N_2171);
and U2203 (N_2203,N_2199,N_2166);
and U2204 (N_2204,N_2186,N_2183);
or U2205 (N_2205,N_2150,N_2191);
or U2206 (N_2206,N_2197,N_2158);
and U2207 (N_2207,N_2185,N_2160);
or U2208 (N_2208,N_2163,N_2167);
or U2209 (N_2209,N_2179,N_2153);
nand U2210 (N_2210,N_2189,N_2178);
nand U2211 (N_2211,N_2194,N_2162);
nor U2212 (N_2212,N_2190,N_2165);
nand U2213 (N_2213,N_2180,N_2168);
xnor U2214 (N_2214,N_2155,N_2154);
or U2215 (N_2215,N_2174,N_2151);
and U2216 (N_2216,N_2172,N_2173);
nor U2217 (N_2217,N_2184,N_2195);
nor U2218 (N_2218,N_2188,N_2159);
and U2219 (N_2219,N_2152,N_2156);
or U2220 (N_2220,N_2157,N_2164);
or U2221 (N_2221,N_2181,N_2198);
nand U2222 (N_2222,N_2161,N_2196);
nand U2223 (N_2223,N_2177,N_2182);
nand U2224 (N_2224,N_2192,N_2187);
nand U2225 (N_2225,N_2163,N_2171);
nor U2226 (N_2226,N_2177,N_2166);
nand U2227 (N_2227,N_2177,N_2168);
and U2228 (N_2228,N_2178,N_2155);
or U2229 (N_2229,N_2167,N_2191);
nand U2230 (N_2230,N_2173,N_2193);
or U2231 (N_2231,N_2155,N_2171);
or U2232 (N_2232,N_2187,N_2177);
and U2233 (N_2233,N_2169,N_2196);
nor U2234 (N_2234,N_2160,N_2165);
and U2235 (N_2235,N_2157,N_2197);
and U2236 (N_2236,N_2180,N_2199);
nand U2237 (N_2237,N_2154,N_2176);
or U2238 (N_2238,N_2186,N_2179);
nor U2239 (N_2239,N_2181,N_2179);
nand U2240 (N_2240,N_2155,N_2184);
xor U2241 (N_2241,N_2167,N_2177);
or U2242 (N_2242,N_2185,N_2181);
and U2243 (N_2243,N_2165,N_2151);
nand U2244 (N_2244,N_2153,N_2195);
or U2245 (N_2245,N_2183,N_2174);
or U2246 (N_2246,N_2173,N_2185);
nand U2247 (N_2247,N_2184,N_2175);
nor U2248 (N_2248,N_2178,N_2170);
and U2249 (N_2249,N_2154,N_2197);
and U2250 (N_2250,N_2204,N_2227);
or U2251 (N_2251,N_2202,N_2237);
nor U2252 (N_2252,N_2242,N_2215);
nand U2253 (N_2253,N_2201,N_2200);
nand U2254 (N_2254,N_2234,N_2205);
or U2255 (N_2255,N_2214,N_2225);
and U2256 (N_2256,N_2207,N_2245);
and U2257 (N_2257,N_2230,N_2222);
xnor U2258 (N_2258,N_2223,N_2209);
or U2259 (N_2259,N_2249,N_2208);
nand U2260 (N_2260,N_2248,N_2231);
nor U2261 (N_2261,N_2220,N_2240);
or U2262 (N_2262,N_2212,N_2219);
or U2263 (N_2263,N_2236,N_2213);
nor U2264 (N_2264,N_2241,N_2210);
and U2265 (N_2265,N_2221,N_2217);
nor U2266 (N_2266,N_2235,N_2226);
or U2267 (N_2267,N_2218,N_2203);
nand U2268 (N_2268,N_2244,N_2224);
and U2269 (N_2269,N_2243,N_2206);
nand U2270 (N_2270,N_2239,N_2229);
nor U2271 (N_2271,N_2246,N_2233);
or U2272 (N_2272,N_2238,N_2247);
nand U2273 (N_2273,N_2232,N_2216);
nor U2274 (N_2274,N_2228,N_2211);
nand U2275 (N_2275,N_2242,N_2210);
and U2276 (N_2276,N_2216,N_2219);
nand U2277 (N_2277,N_2236,N_2200);
or U2278 (N_2278,N_2225,N_2210);
xnor U2279 (N_2279,N_2203,N_2239);
nor U2280 (N_2280,N_2230,N_2249);
or U2281 (N_2281,N_2236,N_2217);
nand U2282 (N_2282,N_2225,N_2247);
and U2283 (N_2283,N_2227,N_2231);
nand U2284 (N_2284,N_2236,N_2220);
or U2285 (N_2285,N_2242,N_2245);
nand U2286 (N_2286,N_2233,N_2247);
or U2287 (N_2287,N_2245,N_2208);
nor U2288 (N_2288,N_2211,N_2209);
xnor U2289 (N_2289,N_2206,N_2218);
and U2290 (N_2290,N_2245,N_2235);
xnor U2291 (N_2291,N_2249,N_2233);
and U2292 (N_2292,N_2246,N_2226);
nor U2293 (N_2293,N_2238,N_2206);
nand U2294 (N_2294,N_2200,N_2249);
or U2295 (N_2295,N_2202,N_2224);
and U2296 (N_2296,N_2244,N_2242);
or U2297 (N_2297,N_2229,N_2211);
nor U2298 (N_2298,N_2225,N_2230);
or U2299 (N_2299,N_2230,N_2210);
nor U2300 (N_2300,N_2273,N_2265);
nand U2301 (N_2301,N_2268,N_2278);
nor U2302 (N_2302,N_2291,N_2254);
nor U2303 (N_2303,N_2255,N_2280);
or U2304 (N_2304,N_2275,N_2263);
and U2305 (N_2305,N_2288,N_2283);
nand U2306 (N_2306,N_2294,N_2258);
and U2307 (N_2307,N_2298,N_2269);
nand U2308 (N_2308,N_2297,N_2257);
nor U2309 (N_2309,N_2296,N_2281);
nand U2310 (N_2310,N_2266,N_2260);
xor U2311 (N_2311,N_2289,N_2272);
xor U2312 (N_2312,N_2290,N_2274);
and U2313 (N_2313,N_2253,N_2287);
and U2314 (N_2314,N_2256,N_2282);
and U2315 (N_2315,N_2284,N_2251);
and U2316 (N_2316,N_2279,N_2299);
nand U2317 (N_2317,N_2276,N_2285);
nor U2318 (N_2318,N_2261,N_2293);
or U2319 (N_2319,N_2262,N_2295);
xor U2320 (N_2320,N_2271,N_2252);
or U2321 (N_2321,N_2250,N_2277);
or U2322 (N_2322,N_2264,N_2270);
or U2323 (N_2323,N_2267,N_2286);
and U2324 (N_2324,N_2259,N_2292);
xor U2325 (N_2325,N_2274,N_2264);
nor U2326 (N_2326,N_2276,N_2283);
and U2327 (N_2327,N_2284,N_2294);
nand U2328 (N_2328,N_2285,N_2267);
nor U2329 (N_2329,N_2264,N_2296);
nor U2330 (N_2330,N_2296,N_2274);
nand U2331 (N_2331,N_2275,N_2297);
and U2332 (N_2332,N_2291,N_2292);
and U2333 (N_2333,N_2272,N_2263);
nand U2334 (N_2334,N_2289,N_2286);
or U2335 (N_2335,N_2260,N_2297);
nand U2336 (N_2336,N_2268,N_2263);
and U2337 (N_2337,N_2291,N_2275);
and U2338 (N_2338,N_2282,N_2278);
nand U2339 (N_2339,N_2256,N_2263);
xnor U2340 (N_2340,N_2297,N_2280);
xor U2341 (N_2341,N_2270,N_2283);
nor U2342 (N_2342,N_2270,N_2294);
or U2343 (N_2343,N_2265,N_2278);
nand U2344 (N_2344,N_2268,N_2298);
and U2345 (N_2345,N_2260,N_2281);
or U2346 (N_2346,N_2296,N_2280);
nor U2347 (N_2347,N_2278,N_2267);
and U2348 (N_2348,N_2275,N_2270);
and U2349 (N_2349,N_2250,N_2263);
nor U2350 (N_2350,N_2317,N_2328);
and U2351 (N_2351,N_2315,N_2324);
nand U2352 (N_2352,N_2300,N_2314);
or U2353 (N_2353,N_2344,N_2341);
nor U2354 (N_2354,N_2332,N_2343);
and U2355 (N_2355,N_2339,N_2345);
xnor U2356 (N_2356,N_2335,N_2322);
and U2357 (N_2357,N_2321,N_2336);
nand U2358 (N_2358,N_2342,N_2302);
and U2359 (N_2359,N_2311,N_2327);
or U2360 (N_2360,N_2318,N_2320);
nor U2361 (N_2361,N_2333,N_2331);
nor U2362 (N_2362,N_2301,N_2308);
nor U2363 (N_2363,N_2305,N_2348);
nor U2364 (N_2364,N_2349,N_2316);
and U2365 (N_2365,N_2326,N_2323);
or U2366 (N_2366,N_2307,N_2310);
nor U2367 (N_2367,N_2346,N_2337);
or U2368 (N_2368,N_2340,N_2338);
and U2369 (N_2369,N_2319,N_2334);
nor U2370 (N_2370,N_2313,N_2312);
nor U2371 (N_2371,N_2325,N_2329);
nand U2372 (N_2372,N_2303,N_2330);
nor U2373 (N_2373,N_2304,N_2306);
and U2374 (N_2374,N_2309,N_2347);
nor U2375 (N_2375,N_2324,N_2339);
or U2376 (N_2376,N_2309,N_2304);
and U2377 (N_2377,N_2318,N_2341);
and U2378 (N_2378,N_2339,N_2315);
xor U2379 (N_2379,N_2316,N_2339);
nand U2380 (N_2380,N_2301,N_2309);
or U2381 (N_2381,N_2337,N_2349);
and U2382 (N_2382,N_2346,N_2300);
nand U2383 (N_2383,N_2305,N_2303);
or U2384 (N_2384,N_2319,N_2346);
nand U2385 (N_2385,N_2348,N_2343);
xnor U2386 (N_2386,N_2308,N_2315);
nor U2387 (N_2387,N_2327,N_2316);
nand U2388 (N_2388,N_2301,N_2307);
and U2389 (N_2389,N_2319,N_2345);
or U2390 (N_2390,N_2340,N_2329);
or U2391 (N_2391,N_2332,N_2325);
nand U2392 (N_2392,N_2317,N_2315);
and U2393 (N_2393,N_2342,N_2344);
nand U2394 (N_2394,N_2300,N_2326);
nand U2395 (N_2395,N_2339,N_2311);
or U2396 (N_2396,N_2318,N_2335);
nor U2397 (N_2397,N_2348,N_2349);
nand U2398 (N_2398,N_2308,N_2321);
or U2399 (N_2399,N_2314,N_2320);
nand U2400 (N_2400,N_2366,N_2354);
and U2401 (N_2401,N_2370,N_2379);
nor U2402 (N_2402,N_2356,N_2399);
or U2403 (N_2403,N_2371,N_2359);
and U2404 (N_2404,N_2391,N_2369);
and U2405 (N_2405,N_2352,N_2388);
nor U2406 (N_2406,N_2384,N_2376);
nand U2407 (N_2407,N_2365,N_2375);
nand U2408 (N_2408,N_2350,N_2381);
nor U2409 (N_2409,N_2394,N_2398);
nor U2410 (N_2410,N_2382,N_2364);
and U2411 (N_2411,N_2380,N_2374);
nor U2412 (N_2412,N_2386,N_2353);
xor U2413 (N_2413,N_2368,N_2378);
nor U2414 (N_2414,N_2396,N_2389);
or U2415 (N_2415,N_2385,N_2387);
xnor U2416 (N_2416,N_2392,N_2395);
nor U2417 (N_2417,N_2372,N_2360);
nor U2418 (N_2418,N_2363,N_2383);
or U2419 (N_2419,N_2367,N_2361);
xor U2420 (N_2420,N_2358,N_2357);
and U2421 (N_2421,N_2351,N_2397);
nand U2422 (N_2422,N_2377,N_2362);
or U2423 (N_2423,N_2355,N_2393);
and U2424 (N_2424,N_2373,N_2390);
xnor U2425 (N_2425,N_2370,N_2398);
or U2426 (N_2426,N_2370,N_2369);
and U2427 (N_2427,N_2398,N_2366);
or U2428 (N_2428,N_2355,N_2376);
nand U2429 (N_2429,N_2354,N_2382);
nor U2430 (N_2430,N_2353,N_2391);
or U2431 (N_2431,N_2374,N_2358);
or U2432 (N_2432,N_2363,N_2373);
nor U2433 (N_2433,N_2370,N_2355);
and U2434 (N_2434,N_2378,N_2385);
nor U2435 (N_2435,N_2386,N_2385);
nor U2436 (N_2436,N_2385,N_2399);
and U2437 (N_2437,N_2394,N_2362);
and U2438 (N_2438,N_2370,N_2361);
and U2439 (N_2439,N_2370,N_2357);
xnor U2440 (N_2440,N_2361,N_2373);
and U2441 (N_2441,N_2368,N_2372);
and U2442 (N_2442,N_2399,N_2351);
nor U2443 (N_2443,N_2355,N_2367);
nand U2444 (N_2444,N_2396,N_2365);
xnor U2445 (N_2445,N_2352,N_2396);
and U2446 (N_2446,N_2351,N_2359);
or U2447 (N_2447,N_2398,N_2374);
nand U2448 (N_2448,N_2379,N_2398);
and U2449 (N_2449,N_2365,N_2353);
nand U2450 (N_2450,N_2416,N_2446);
nor U2451 (N_2451,N_2440,N_2402);
and U2452 (N_2452,N_2413,N_2445);
and U2453 (N_2453,N_2420,N_2410);
and U2454 (N_2454,N_2443,N_2426);
nor U2455 (N_2455,N_2444,N_2401);
nand U2456 (N_2456,N_2414,N_2422);
and U2457 (N_2457,N_2435,N_2406);
or U2458 (N_2458,N_2442,N_2412);
and U2459 (N_2459,N_2449,N_2404);
or U2460 (N_2460,N_2409,N_2428);
and U2461 (N_2461,N_2441,N_2431);
nor U2462 (N_2462,N_2448,N_2419);
and U2463 (N_2463,N_2423,N_2424);
or U2464 (N_2464,N_2430,N_2432);
nor U2465 (N_2465,N_2439,N_2408);
nor U2466 (N_2466,N_2433,N_2403);
and U2467 (N_2467,N_2407,N_2438);
nand U2468 (N_2468,N_2427,N_2421);
or U2469 (N_2469,N_2400,N_2436);
nor U2470 (N_2470,N_2405,N_2447);
or U2471 (N_2471,N_2425,N_2418);
nand U2472 (N_2472,N_2429,N_2437);
nand U2473 (N_2473,N_2417,N_2411);
nand U2474 (N_2474,N_2434,N_2415);
and U2475 (N_2475,N_2442,N_2406);
and U2476 (N_2476,N_2400,N_2416);
and U2477 (N_2477,N_2415,N_2403);
or U2478 (N_2478,N_2403,N_2406);
nor U2479 (N_2479,N_2412,N_2415);
and U2480 (N_2480,N_2431,N_2438);
and U2481 (N_2481,N_2449,N_2416);
or U2482 (N_2482,N_2434,N_2400);
nor U2483 (N_2483,N_2440,N_2403);
and U2484 (N_2484,N_2409,N_2402);
or U2485 (N_2485,N_2427,N_2401);
or U2486 (N_2486,N_2425,N_2433);
nor U2487 (N_2487,N_2433,N_2429);
and U2488 (N_2488,N_2428,N_2431);
nand U2489 (N_2489,N_2419,N_2406);
nor U2490 (N_2490,N_2424,N_2415);
nor U2491 (N_2491,N_2429,N_2423);
or U2492 (N_2492,N_2442,N_2426);
nand U2493 (N_2493,N_2443,N_2432);
xor U2494 (N_2494,N_2429,N_2442);
nand U2495 (N_2495,N_2414,N_2409);
nor U2496 (N_2496,N_2423,N_2422);
xnor U2497 (N_2497,N_2419,N_2415);
xnor U2498 (N_2498,N_2437,N_2447);
or U2499 (N_2499,N_2402,N_2428);
and U2500 (N_2500,N_2467,N_2471);
nor U2501 (N_2501,N_2483,N_2459);
nand U2502 (N_2502,N_2491,N_2461);
or U2503 (N_2503,N_2477,N_2475);
and U2504 (N_2504,N_2482,N_2474);
nand U2505 (N_2505,N_2495,N_2454);
and U2506 (N_2506,N_2457,N_2487);
nand U2507 (N_2507,N_2462,N_2498);
nand U2508 (N_2508,N_2486,N_2492);
nand U2509 (N_2509,N_2489,N_2496);
nand U2510 (N_2510,N_2452,N_2468);
nand U2511 (N_2511,N_2490,N_2485);
and U2512 (N_2512,N_2478,N_2456);
nand U2513 (N_2513,N_2480,N_2464);
nand U2514 (N_2514,N_2451,N_2455);
nand U2515 (N_2515,N_2458,N_2484);
or U2516 (N_2516,N_2463,N_2497);
nand U2517 (N_2517,N_2465,N_2499);
nor U2518 (N_2518,N_2472,N_2488);
or U2519 (N_2519,N_2460,N_2466);
nand U2520 (N_2520,N_2481,N_2479);
or U2521 (N_2521,N_2473,N_2470);
and U2522 (N_2522,N_2476,N_2450);
nand U2523 (N_2523,N_2494,N_2493);
nand U2524 (N_2524,N_2469,N_2453);
nand U2525 (N_2525,N_2464,N_2492);
nor U2526 (N_2526,N_2465,N_2494);
nor U2527 (N_2527,N_2456,N_2491);
and U2528 (N_2528,N_2456,N_2495);
nor U2529 (N_2529,N_2482,N_2458);
or U2530 (N_2530,N_2482,N_2471);
and U2531 (N_2531,N_2463,N_2468);
and U2532 (N_2532,N_2462,N_2451);
nor U2533 (N_2533,N_2479,N_2457);
nor U2534 (N_2534,N_2461,N_2475);
or U2535 (N_2535,N_2494,N_2480);
nor U2536 (N_2536,N_2488,N_2460);
xnor U2537 (N_2537,N_2496,N_2470);
nand U2538 (N_2538,N_2466,N_2480);
and U2539 (N_2539,N_2474,N_2450);
nor U2540 (N_2540,N_2487,N_2456);
xnor U2541 (N_2541,N_2475,N_2454);
nand U2542 (N_2542,N_2480,N_2460);
or U2543 (N_2543,N_2477,N_2481);
or U2544 (N_2544,N_2478,N_2492);
nand U2545 (N_2545,N_2475,N_2490);
or U2546 (N_2546,N_2455,N_2485);
nand U2547 (N_2547,N_2467,N_2464);
and U2548 (N_2548,N_2456,N_2492);
xnor U2549 (N_2549,N_2457,N_2450);
xor U2550 (N_2550,N_2541,N_2515);
or U2551 (N_2551,N_2535,N_2549);
nand U2552 (N_2552,N_2543,N_2523);
or U2553 (N_2553,N_2519,N_2518);
or U2554 (N_2554,N_2533,N_2527);
or U2555 (N_2555,N_2531,N_2534);
and U2556 (N_2556,N_2503,N_2505);
nand U2557 (N_2557,N_2524,N_2508);
or U2558 (N_2558,N_2522,N_2528);
or U2559 (N_2559,N_2545,N_2509);
and U2560 (N_2560,N_2500,N_2511);
xnor U2561 (N_2561,N_2539,N_2525);
nand U2562 (N_2562,N_2520,N_2529);
and U2563 (N_2563,N_2514,N_2526);
nand U2564 (N_2564,N_2502,N_2530);
xor U2565 (N_2565,N_2538,N_2537);
nor U2566 (N_2566,N_2547,N_2546);
nand U2567 (N_2567,N_2504,N_2516);
nand U2568 (N_2568,N_2506,N_2544);
nor U2569 (N_2569,N_2513,N_2501);
and U2570 (N_2570,N_2521,N_2540);
nand U2571 (N_2571,N_2532,N_2548);
nand U2572 (N_2572,N_2536,N_2517);
nor U2573 (N_2573,N_2512,N_2507);
and U2574 (N_2574,N_2542,N_2510);
and U2575 (N_2575,N_2537,N_2548);
nand U2576 (N_2576,N_2503,N_2527);
xor U2577 (N_2577,N_2523,N_2520);
or U2578 (N_2578,N_2547,N_2516);
or U2579 (N_2579,N_2544,N_2536);
nand U2580 (N_2580,N_2512,N_2538);
or U2581 (N_2581,N_2513,N_2525);
nand U2582 (N_2582,N_2548,N_2528);
and U2583 (N_2583,N_2521,N_2526);
xnor U2584 (N_2584,N_2547,N_2515);
nor U2585 (N_2585,N_2528,N_2545);
or U2586 (N_2586,N_2504,N_2536);
nand U2587 (N_2587,N_2545,N_2504);
nand U2588 (N_2588,N_2508,N_2545);
and U2589 (N_2589,N_2547,N_2545);
and U2590 (N_2590,N_2515,N_2526);
and U2591 (N_2591,N_2531,N_2510);
and U2592 (N_2592,N_2502,N_2544);
nand U2593 (N_2593,N_2511,N_2526);
nand U2594 (N_2594,N_2503,N_2544);
and U2595 (N_2595,N_2512,N_2518);
nand U2596 (N_2596,N_2511,N_2502);
or U2597 (N_2597,N_2510,N_2525);
nor U2598 (N_2598,N_2516,N_2514);
or U2599 (N_2599,N_2539,N_2542);
xnor U2600 (N_2600,N_2598,N_2591);
xnor U2601 (N_2601,N_2574,N_2564);
and U2602 (N_2602,N_2560,N_2572);
and U2603 (N_2603,N_2551,N_2565);
nor U2604 (N_2604,N_2562,N_2558);
xor U2605 (N_2605,N_2555,N_2559);
or U2606 (N_2606,N_2581,N_2577);
and U2607 (N_2607,N_2567,N_2585);
or U2608 (N_2608,N_2583,N_2576);
or U2609 (N_2609,N_2568,N_2561);
or U2610 (N_2610,N_2592,N_2557);
and U2611 (N_2611,N_2579,N_2586);
nor U2612 (N_2612,N_2573,N_2595);
or U2613 (N_2613,N_2578,N_2587);
nor U2614 (N_2614,N_2582,N_2597);
xnor U2615 (N_2615,N_2550,N_2554);
or U2616 (N_2616,N_2553,N_2589);
and U2617 (N_2617,N_2580,N_2566);
or U2618 (N_2618,N_2594,N_2596);
nor U2619 (N_2619,N_2556,N_2563);
and U2620 (N_2620,N_2588,N_2590);
nand U2621 (N_2621,N_2552,N_2593);
nand U2622 (N_2622,N_2584,N_2570);
or U2623 (N_2623,N_2599,N_2569);
and U2624 (N_2624,N_2575,N_2571);
xor U2625 (N_2625,N_2594,N_2575);
nor U2626 (N_2626,N_2566,N_2561);
nand U2627 (N_2627,N_2568,N_2575);
nand U2628 (N_2628,N_2556,N_2555);
xnor U2629 (N_2629,N_2599,N_2576);
or U2630 (N_2630,N_2582,N_2587);
nand U2631 (N_2631,N_2585,N_2551);
or U2632 (N_2632,N_2582,N_2589);
xor U2633 (N_2633,N_2564,N_2572);
nor U2634 (N_2634,N_2562,N_2585);
and U2635 (N_2635,N_2554,N_2560);
xnor U2636 (N_2636,N_2552,N_2586);
and U2637 (N_2637,N_2577,N_2566);
nor U2638 (N_2638,N_2572,N_2566);
nand U2639 (N_2639,N_2585,N_2553);
nand U2640 (N_2640,N_2595,N_2556);
nand U2641 (N_2641,N_2558,N_2552);
or U2642 (N_2642,N_2574,N_2585);
or U2643 (N_2643,N_2554,N_2596);
nand U2644 (N_2644,N_2576,N_2571);
xnor U2645 (N_2645,N_2562,N_2568);
nand U2646 (N_2646,N_2580,N_2596);
or U2647 (N_2647,N_2583,N_2560);
or U2648 (N_2648,N_2562,N_2551);
and U2649 (N_2649,N_2558,N_2564);
and U2650 (N_2650,N_2605,N_2628);
nor U2651 (N_2651,N_2610,N_2625);
or U2652 (N_2652,N_2642,N_2644);
nor U2653 (N_2653,N_2601,N_2613);
or U2654 (N_2654,N_2614,N_2649);
xor U2655 (N_2655,N_2647,N_2602);
xnor U2656 (N_2656,N_2626,N_2609);
nor U2657 (N_2657,N_2618,N_2627);
and U2658 (N_2658,N_2616,N_2639);
or U2659 (N_2659,N_2603,N_2608);
nand U2660 (N_2660,N_2623,N_2637);
nand U2661 (N_2661,N_2646,N_2615);
nor U2662 (N_2662,N_2641,N_2643);
nand U2663 (N_2663,N_2633,N_2622);
or U2664 (N_2664,N_2631,N_2635);
and U2665 (N_2665,N_2629,N_2607);
nor U2666 (N_2666,N_2612,N_2634);
nor U2667 (N_2667,N_2617,N_2620);
nand U2668 (N_2668,N_2624,N_2640);
or U2669 (N_2669,N_2645,N_2638);
nand U2670 (N_2670,N_2648,N_2604);
and U2671 (N_2671,N_2600,N_2621);
nand U2672 (N_2672,N_2606,N_2611);
nor U2673 (N_2673,N_2632,N_2619);
nand U2674 (N_2674,N_2630,N_2636);
or U2675 (N_2675,N_2621,N_2609);
and U2676 (N_2676,N_2642,N_2621);
or U2677 (N_2677,N_2602,N_2644);
nand U2678 (N_2678,N_2601,N_2612);
or U2679 (N_2679,N_2613,N_2600);
nand U2680 (N_2680,N_2610,N_2620);
nand U2681 (N_2681,N_2602,N_2611);
nor U2682 (N_2682,N_2621,N_2630);
nand U2683 (N_2683,N_2610,N_2617);
and U2684 (N_2684,N_2612,N_2626);
nor U2685 (N_2685,N_2612,N_2643);
and U2686 (N_2686,N_2614,N_2624);
nor U2687 (N_2687,N_2623,N_2621);
nand U2688 (N_2688,N_2603,N_2628);
and U2689 (N_2689,N_2636,N_2622);
nand U2690 (N_2690,N_2611,N_2628);
and U2691 (N_2691,N_2647,N_2627);
nor U2692 (N_2692,N_2624,N_2610);
nand U2693 (N_2693,N_2613,N_2624);
nor U2694 (N_2694,N_2629,N_2628);
or U2695 (N_2695,N_2638,N_2626);
nor U2696 (N_2696,N_2640,N_2648);
and U2697 (N_2697,N_2643,N_2610);
nand U2698 (N_2698,N_2648,N_2631);
and U2699 (N_2699,N_2645,N_2616);
or U2700 (N_2700,N_2668,N_2681);
nand U2701 (N_2701,N_2690,N_2672);
nor U2702 (N_2702,N_2652,N_2675);
or U2703 (N_2703,N_2650,N_2686);
nor U2704 (N_2704,N_2671,N_2666);
or U2705 (N_2705,N_2697,N_2678);
nor U2706 (N_2706,N_2688,N_2656);
nand U2707 (N_2707,N_2653,N_2696);
nand U2708 (N_2708,N_2677,N_2657);
and U2709 (N_2709,N_2655,N_2669);
nor U2710 (N_2710,N_2692,N_2654);
nand U2711 (N_2711,N_2694,N_2699);
xnor U2712 (N_2712,N_2661,N_2670);
or U2713 (N_2713,N_2662,N_2667);
and U2714 (N_2714,N_2685,N_2674);
and U2715 (N_2715,N_2698,N_2689);
xnor U2716 (N_2716,N_2691,N_2679);
xor U2717 (N_2717,N_2664,N_2660);
or U2718 (N_2718,N_2676,N_2687);
nand U2719 (N_2719,N_2658,N_2673);
or U2720 (N_2720,N_2659,N_2695);
nand U2721 (N_2721,N_2663,N_2665);
nor U2722 (N_2722,N_2683,N_2651);
nand U2723 (N_2723,N_2682,N_2684);
and U2724 (N_2724,N_2693,N_2680);
xor U2725 (N_2725,N_2651,N_2668);
or U2726 (N_2726,N_2675,N_2673);
or U2727 (N_2727,N_2654,N_2699);
xnor U2728 (N_2728,N_2674,N_2658);
and U2729 (N_2729,N_2683,N_2686);
nand U2730 (N_2730,N_2651,N_2655);
or U2731 (N_2731,N_2668,N_2659);
nand U2732 (N_2732,N_2686,N_2693);
nor U2733 (N_2733,N_2653,N_2698);
and U2734 (N_2734,N_2654,N_2688);
nor U2735 (N_2735,N_2661,N_2651);
xor U2736 (N_2736,N_2692,N_2680);
and U2737 (N_2737,N_2699,N_2686);
or U2738 (N_2738,N_2677,N_2654);
or U2739 (N_2739,N_2668,N_2694);
or U2740 (N_2740,N_2656,N_2665);
and U2741 (N_2741,N_2667,N_2694);
or U2742 (N_2742,N_2674,N_2664);
nand U2743 (N_2743,N_2698,N_2668);
and U2744 (N_2744,N_2691,N_2658);
or U2745 (N_2745,N_2699,N_2697);
or U2746 (N_2746,N_2658,N_2661);
nand U2747 (N_2747,N_2673,N_2693);
nand U2748 (N_2748,N_2678,N_2696);
xor U2749 (N_2749,N_2661,N_2685);
nor U2750 (N_2750,N_2714,N_2707);
and U2751 (N_2751,N_2717,N_2725);
nand U2752 (N_2752,N_2735,N_2738);
or U2753 (N_2753,N_2744,N_2721);
and U2754 (N_2754,N_2718,N_2704);
nor U2755 (N_2755,N_2743,N_2749);
nor U2756 (N_2756,N_2745,N_2739);
or U2757 (N_2757,N_2736,N_2734);
xor U2758 (N_2758,N_2710,N_2701);
or U2759 (N_2759,N_2715,N_2708);
nand U2760 (N_2760,N_2731,N_2737);
nand U2761 (N_2761,N_2742,N_2726);
nand U2762 (N_2762,N_2747,N_2730);
and U2763 (N_2763,N_2748,N_2702);
xnor U2764 (N_2764,N_2703,N_2740);
or U2765 (N_2765,N_2746,N_2719);
nor U2766 (N_2766,N_2741,N_2713);
and U2767 (N_2767,N_2705,N_2729);
and U2768 (N_2768,N_2700,N_2723);
nor U2769 (N_2769,N_2716,N_2706);
nand U2770 (N_2770,N_2720,N_2733);
and U2771 (N_2771,N_2722,N_2724);
or U2772 (N_2772,N_2712,N_2732);
xnor U2773 (N_2773,N_2728,N_2727);
or U2774 (N_2774,N_2709,N_2711);
nor U2775 (N_2775,N_2728,N_2700);
and U2776 (N_2776,N_2726,N_2739);
and U2777 (N_2777,N_2736,N_2742);
nand U2778 (N_2778,N_2700,N_2707);
nand U2779 (N_2779,N_2740,N_2717);
or U2780 (N_2780,N_2728,N_2722);
nor U2781 (N_2781,N_2740,N_2706);
or U2782 (N_2782,N_2721,N_2706);
or U2783 (N_2783,N_2734,N_2711);
and U2784 (N_2784,N_2711,N_2735);
nand U2785 (N_2785,N_2748,N_2726);
and U2786 (N_2786,N_2744,N_2727);
xor U2787 (N_2787,N_2715,N_2720);
or U2788 (N_2788,N_2711,N_2733);
or U2789 (N_2789,N_2710,N_2722);
and U2790 (N_2790,N_2720,N_2728);
nand U2791 (N_2791,N_2705,N_2715);
nor U2792 (N_2792,N_2726,N_2701);
and U2793 (N_2793,N_2712,N_2747);
nor U2794 (N_2794,N_2729,N_2728);
nor U2795 (N_2795,N_2741,N_2725);
or U2796 (N_2796,N_2715,N_2717);
nand U2797 (N_2797,N_2711,N_2700);
nand U2798 (N_2798,N_2700,N_2717);
nor U2799 (N_2799,N_2713,N_2749);
nand U2800 (N_2800,N_2754,N_2767);
xnor U2801 (N_2801,N_2786,N_2756);
or U2802 (N_2802,N_2752,N_2776);
or U2803 (N_2803,N_2769,N_2753);
nor U2804 (N_2804,N_2763,N_2755);
nor U2805 (N_2805,N_2760,N_2783);
nand U2806 (N_2806,N_2773,N_2781);
nand U2807 (N_2807,N_2759,N_2770);
nand U2808 (N_2808,N_2788,N_2791);
or U2809 (N_2809,N_2779,N_2789);
nand U2810 (N_2810,N_2777,N_2797);
or U2811 (N_2811,N_2750,N_2757);
and U2812 (N_2812,N_2758,N_2794);
nor U2813 (N_2813,N_2798,N_2766);
and U2814 (N_2814,N_2775,N_2762);
and U2815 (N_2815,N_2780,N_2795);
nand U2816 (N_2816,N_2774,N_2792);
or U2817 (N_2817,N_2771,N_2784);
nor U2818 (N_2818,N_2782,N_2761);
nor U2819 (N_2819,N_2768,N_2787);
or U2820 (N_2820,N_2765,N_2751);
nand U2821 (N_2821,N_2799,N_2764);
xor U2822 (N_2822,N_2790,N_2778);
nand U2823 (N_2823,N_2772,N_2793);
nor U2824 (N_2824,N_2796,N_2785);
or U2825 (N_2825,N_2758,N_2768);
or U2826 (N_2826,N_2789,N_2751);
or U2827 (N_2827,N_2763,N_2776);
xnor U2828 (N_2828,N_2774,N_2754);
nand U2829 (N_2829,N_2765,N_2757);
or U2830 (N_2830,N_2753,N_2752);
or U2831 (N_2831,N_2764,N_2762);
or U2832 (N_2832,N_2751,N_2759);
and U2833 (N_2833,N_2792,N_2783);
nand U2834 (N_2834,N_2763,N_2782);
or U2835 (N_2835,N_2754,N_2798);
nand U2836 (N_2836,N_2781,N_2753);
and U2837 (N_2837,N_2771,N_2762);
nand U2838 (N_2838,N_2781,N_2759);
nand U2839 (N_2839,N_2763,N_2788);
and U2840 (N_2840,N_2787,N_2784);
nand U2841 (N_2841,N_2779,N_2754);
nand U2842 (N_2842,N_2750,N_2782);
nand U2843 (N_2843,N_2788,N_2751);
nand U2844 (N_2844,N_2787,N_2771);
or U2845 (N_2845,N_2785,N_2755);
nand U2846 (N_2846,N_2768,N_2798);
and U2847 (N_2847,N_2791,N_2781);
nor U2848 (N_2848,N_2758,N_2751);
and U2849 (N_2849,N_2792,N_2766);
nor U2850 (N_2850,N_2817,N_2821);
nor U2851 (N_2851,N_2813,N_2842);
xor U2852 (N_2852,N_2811,N_2812);
or U2853 (N_2853,N_2844,N_2839);
nand U2854 (N_2854,N_2822,N_2808);
or U2855 (N_2855,N_2829,N_2832);
nand U2856 (N_2856,N_2810,N_2803);
nand U2857 (N_2857,N_2837,N_2835);
nand U2858 (N_2858,N_2845,N_2816);
nand U2859 (N_2859,N_2807,N_2833);
nand U2860 (N_2860,N_2849,N_2802);
nor U2861 (N_2861,N_2826,N_2834);
and U2862 (N_2862,N_2800,N_2801);
or U2863 (N_2863,N_2830,N_2818);
or U2864 (N_2864,N_2848,N_2824);
nand U2865 (N_2865,N_2815,N_2819);
and U2866 (N_2866,N_2846,N_2820);
nor U2867 (N_2867,N_2806,N_2804);
nor U2868 (N_2868,N_2841,N_2831);
or U2869 (N_2869,N_2847,N_2825);
or U2870 (N_2870,N_2827,N_2823);
and U2871 (N_2871,N_2805,N_2838);
or U2872 (N_2872,N_2809,N_2843);
or U2873 (N_2873,N_2828,N_2840);
nand U2874 (N_2874,N_2814,N_2836);
nor U2875 (N_2875,N_2812,N_2820);
or U2876 (N_2876,N_2834,N_2809);
nor U2877 (N_2877,N_2828,N_2837);
or U2878 (N_2878,N_2838,N_2806);
nand U2879 (N_2879,N_2826,N_2801);
or U2880 (N_2880,N_2839,N_2815);
and U2881 (N_2881,N_2828,N_2841);
and U2882 (N_2882,N_2836,N_2843);
nor U2883 (N_2883,N_2811,N_2841);
nand U2884 (N_2884,N_2848,N_2807);
and U2885 (N_2885,N_2819,N_2805);
xor U2886 (N_2886,N_2846,N_2812);
xnor U2887 (N_2887,N_2800,N_2813);
nand U2888 (N_2888,N_2805,N_2814);
xor U2889 (N_2889,N_2805,N_2845);
nand U2890 (N_2890,N_2816,N_2804);
and U2891 (N_2891,N_2801,N_2813);
and U2892 (N_2892,N_2808,N_2846);
nor U2893 (N_2893,N_2841,N_2812);
nor U2894 (N_2894,N_2803,N_2836);
nand U2895 (N_2895,N_2810,N_2844);
or U2896 (N_2896,N_2819,N_2807);
nand U2897 (N_2897,N_2814,N_2842);
nor U2898 (N_2898,N_2832,N_2816);
nand U2899 (N_2899,N_2807,N_2847);
or U2900 (N_2900,N_2856,N_2873);
nand U2901 (N_2901,N_2880,N_2864);
and U2902 (N_2902,N_2868,N_2857);
or U2903 (N_2903,N_2896,N_2859);
nor U2904 (N_2904,N_2899,N_2869);
nor U2905 (N_2905,N_2867,N_2866);
or U2906 (N_2906,N_2892,N_2854);
xor U2907 (N_2907,N_2874,N_2897);
and U2908 (N_2908,N_2883,N_2872);
and U2909 (N_2909,N_2852,N_2885);
and U2910 (N_2910,N_2895,N_2853);
and U2911 (N_2911,N_2887,N_2875);
xor U2912 (N_2912,N_2858,N_2850);
nor U2913 (N_2913,N_2893,N_2881);
or U2914 (N_2914,N_2863,N_2865);
nor U2915 (N_2915,N_2879,N_2884);
nand U2916 (N_2916,N_2861,N_2898);
nor U2917 (N_2917,N_2877,N_2878);
nor U2918 (N_2918,N_2882,N_2862);
and U2919 (N_2919,N_2860,N_2894);
nor U2920 (N_2920,N_2871,N_2851);
nand U2921 (N_2921,N_2890,N_2889);
and U2922 (N_2922,N_2886,N_2891);
or U2923 (N_2923,N_2876,N_2870);
and U2924 (N_2924,N_2888,N_2855);
or U2925 (N_2925,N_2873,N_2874);
nand U2926 (N_2926,N_2876,N_2886);
nand U2927 (N_2927,N_2877,N_2869);
nand U2928 (N_2928,N_2865,N_2889);
nor U2929 (N_2929,N_2857,N_2884);
nor U2930 (N_2930,N_2865,N_2894);
nor U2931 (N_2931,N_2869,N_2878);
and U2932 (N_2932,N_2899,N_2852);
nand U2933 (N_2933,N_2868,N_2864);
and U2934 (N_2934,N_2893,N_2872);
nor U2935 (N_2935,N_2852,N_2870);
nand U2936 (N_2936,N_2875,N_2864);
nand U2937 (N_2937,N_2858,N_2870);
and U2938 (N_2938,N_2897,N_2885);
or U2939 (N_2939,N_2885,N_2858);
nand U2940 (N_2940,N_2859,N_2885);
or U2941 (N_2941,N_2891,N_2890);
or U2942 (N_2942,N_2867,N_2881);
nor U2943 (N_2943,N_2869,N_2850);
nand U2944 (N_2944,N_2893,N_2868);
or U2945 (N_2945,N_2894,N_2886);
nand U2946 (N_2946,N_2896,N_2866);
nor U2947 (N_2947,N_2885,N_2888);
or U2948 (N_2948,N_2860,N_2880);
nor U2949 (N_2949,N_2896,N_2875);
or U2950 (N_2950,N_2919,N_2925);
nand U2951 (N_2951,N_2933,N_2935);
nand U2952 (N_2952,N_2915,N_2923);
xor U2953 (N_2953,N_2934,N_2909);
or U2954 (N_2954,N_2926,N_2922);
and U2955 (N_2955,N_2931,N_2949);
xnor U2956 (N_2956,N_2900,N_2944);
xnor U2957 (N_2957,N_2902,N_2917);
nor U2958 (N_2958,N_2906,N_2938);
and U2959 (N_2959,N_2920,N_2937);
nor U2960 (N_2960,N_2904,N_2929);
nor U2961 (N_2961,N_2908,N_2911);
or U2962 (N_2962,N_2936,N_2918);
or U2963 (N_2963,N_2942,N_2945);
xnor U2964 (N_2964,N_2905,N_2901);
or U2965 (N_2965,N_2921,N_2903);
nor U2966 (N_2966,N_2940,N_2939);
and U2967 (N_2967,N_2928,N_2941);
nand U2968 (N_2968,N_2948,N_2927);
and U2969 (N_2969,N_2946,N_2914);
or U2970 (N_2970,N_2912,N_2907);
nand U2971 (N_2971,N_2924,N_2947);
nor U2972 (N_2972,N_2932,N_2943);
or U2973 (N_2973,N_2930,N_2910);
and U2974 (N_2974,N_2916,N_2913);
or U2975 (N_2975,N_2924,N_2916);
and U2976 (N_2976,N_2903,N_2923);
and U2977 (N_2977,N_2919,N_2912);
or U2978 (N_2978,N_2914,N_2911);
and U2979 (N_2979,N_2933,N_2916);
nor U2980 (N_2980,N_2918,N_2901);
xor U2981 (N_2981,N_2912,N_2917);
nor U2982 (N_2982,N_2938,N_2903);
nand U2983 (N_2983,N_2937,N_2929);
nand U2984 (N_2984,N_2913,N_2911);
and U2985 (N_2985,N_2942,N_2941);
and U2986 (N_2986,N_2920,N_2906);
nor U2987 (N_2987,N_2907,N_2936);
or U2988 (N_2988,N_2924,N_2938);
nand U2989 (N_2989,N_2924,N_2904);
or U2990 (N_2990,N_2930,N_2926);
nand U2991 (N_2991,N_2942,N_2924);
and U2992 (N_2992,N_2908,N_2924);
nand U2993 (N_2993,N_2949,N_2900);
or U2994 (N_2994,N_2915,N_2942);
or U2995 (N_2995,N_2922,N_2902);
xnor U2996 (N_2996,N_2917,N_2921);
nor U2997 (N_2997,N_2919,N_2918);
nor U2998 (N_2998,N_2915,N_2943);
nand U2999 (N_2999,N_2914,N_2926);
or UO_0 (O_0,N_2969,N_2992);
or UO_1 (O_1,N_2984,N_2971);
or UO_2 (O_2,N_2989,N_2996);
nand UO_3 (O_3,N_2995,N_2999);
and UO_4 (O_4,N_2973,N_2993);
nand UO_5 (O_5,N_2965,N_2967);
or UO_6 (O_6,N_2958,N_2957);
nor UO_7 (O_7,N_2953,N_2951);
xor UO_8 (O_8,N_2991,N_2963);
and UO_9 (O_9,N_2961,N_2976);
nand UO_10 (O_10,N_2970,N_2974);
nand UO_11 (O_11,N_2972,N_2980);
nor UO_12 (O_12,N_2998,N_2952);
nand UO_13 (O_13,N_2985,N_2981);
nand UO_14 (O_14,N_2968,N_2954);
and UO_15 (O_15,N_2960,N_2983);
nand UO_16 (O_16,N_2986,N_2956);
nor UO_17 (O_17,N_2997,N_2979);
and UO_18 (O_18,N_2964,N_2987);
nand UO_19 (O_19,N_2994,N_2978);
and UO_20 (O_20,N_2988,N_2966);
or UO_21 (O_21,N_2959,N_2962);
nor UO_22 (O_22,N_2990,N_2975);
or UO_23 (O_23,N_2950,N_2955);
nor UO_24 (O_24,N_2977,N_2982);
and UO_25 (O_25,N_2975,N_2984);
nand UO_26 (O_26,N_2966,N_2967);
or UO_27 (O_27,N_2960,N_2972);
or UO_28 (O_28,N_2975,N_2956);
and UO_29 (O_29,N_2951,N_2961);
nand UO_30 (O_30,N_2973,N_2954);
and UO_31 (O_31,N_2966,N_2989);
nor UO_32 (O_32,N_2991,N_2956);
or UO_33 (O_33,N_2984,N_2985);
xnor UO_34 (O_34,N_2966,N_2997);
nor UO_35 (O_35,N_2950,N_2999);
and UO_36 (O_36,N_2977,N_2999);
nor UO_37 (O_37,N_2952,N_2991);
and UO_38 (O_38,N_2958,N_2974);
nand UO_39 (O_39,N_2955,N_2954);
nor UO_40 (O_40,N_2983,N_2993);
nand UO_41 (O_41,N_2961,N_2967);
nand UO_42 (O_42,N_2979,N_2967);
nor UO_43 (O_43,N_2988,N_2959);
nand UO_44 (O_44,N_2970,N_2961);
nand UO_45 (O_45,N_2962,N_2958);
nor UO_46 (O_46,N_2993,N_2978);
or UO_47 (O_47,N_2962,N_2952);
or UO_48 (O_48,N_2969,N_2999);
and UO_49 (O_49,N_2981,N_2986);
and UO_50 (O_50,N_2980,N_2971);
and UO_51 (O_51,N_2999,N_2997);
xor UO_52 (O_52,N_2976,N_2962);
or UO_53 (O_53,N_2960,N_2975);
and UO_54 (O_54,N_2972,N_2997);
and UO_55 (O_55,N_2950,N_2953);
nor UO_56 (O_56,N_2982,N_2997);
and UO_57 (O_57,N_2994,N_2983);
nand UO_58 (O_58,N_2960,N_2961);
nand UO_59 (O_59,N_2964,N_2952);
or UO_60 (O_60,N_2976,N_2968);
nor UO_61 (O_61,N_2977,N_2975);
or UO_62 (O_62,N_2983,N_2954);
nand UO_63 (O_63,N_2955,N_2982);
nand UO_64 (O_64,N_2953,N_2999);
nor UO_65 (O_65,N_2999,N_2987);
and UO_66 (O_66,N_2980,N_2984);
xnor UO_67 (O_67,N_2982,N_2973);
xor UO_68 (O_68,N_2999,N_2967);
xnor UO_69 (O_69,N_2989,N_2955);
or UO_70 (O_70,N_2977,N_2995);
nor UO_71 (O_71,N_2963,N_2952);
or UO_72 (O_72,N_2992,N_2960);
or UO_73 (O_73,N_2982,N_2994);
nand UO_74 (O_74,N_2984,N_2951);
nand UO_75 (O_75,N_2978,N_2981);
or UO_76 (O_76,N_2959,N_2980);
nor UO_77 (O_77,N_2977,N_2998);
nor UO_78 (O_78,N_2978,N_2963);
nand UO_79 (O_79,N_2998,N_2981);
nor UO_80 (O_80,N_2967,N_2983);
or UO_81 (O_81,N_2963,N_2985);
and UO_82 (O_82,N_2996,N_2969);
and UO_83 (O_83,N_2955,N_2994);
and UO_84 (O_84,N_2958,N_2986);
or UO_85 (O_85,N_2977,N_2953);
or UO_86 (O_86,N_2951,N_2956);
and UO_87 (O_87,N_2973,N_2968);
xnor UO_88 (O_88,N_2960,N_2999);
or UO_89 (O_89,N_2960,N_2980);
and UO_90 (O_90,N_2956,N_2999);
nand UO_91 (O_91,N_2955,N_2969);
xnor UO_92 (O_92,N_2993,N_2979);
nor UO_93 (O_93,N_2982,N_2974);
nand UO_94 (O_94,N_2987,N_2998);
nor UO_95 (O_95,N_2997,N_2975);
or UO_96 (O_96,N_2967,N_2985);
nand UO_97 (O_97,N_2952,N_2977);
xnor UO_98 (O_98,N_2950,N_2977);
nor UO_99 (O_99,N_2951,N_2978);
or UO_100 (O_100,N_2966,N_2985);
nand UO_101 (O_101,N_2969,N_2971);
and UO_102 (O_102,N_2995,N_2988);
nand UO_103 (O_103,N_2959,N_2969);
nor UO_104 (O_104,N_2980,N_2950);
or UO_105 (O_105,N_2987,N_2950);
nor UO_106 (O_106,N_2962,N_2960);
or UO_107 (O_107,N_2985,N_2983);
xnor UO_108 (O_108,N_2959,N_2993);
and UO_109 (O_109,N_2968,N_2959);
or UO_110 (O_110,N_2997,N_2977);
nor UO_111 (O_111,N_2960,N_2995);
or UO_112 (O_112,N_2957,N_2963);
nor UO_113 (O_113,N_2982,N_2972);
and UO_114 (O_114,N_2982,N_2967);
and UO_115 (O_115,N_2957,N_2955);
nor UO_116 (O_116,N_2994,N_2951);
and UO_117 (O_117,N_2987,N_2968);
nand UO_118 (O_118,N_2984,N_2958);
and UO_119 (O_119,N_2973,N_2964);
nand UO_120 (O_120,N_2955,N_2980);
or UO_121 (O_121,N_2978,N_2991);
or UO_122 (O_122,N_2968,N_2961);
nand UO_123 (O_123,N_2965,N_2990);
xnor UO_124 (O_124,N_2982,N_2988);
or UO_125 (O_125,N_2993,N_2989);
nor UO_126 (O_126,N_2960,N_2987);
or UO_127 (O_127,N_2988,N_2979);
and UO_128 (O_128,N_2965,N_2994);
nand UO_129 (O_129,N_2958,N_2955);
nand UO_130 (O_130,N_2957,N_2982);
nor UO_131 (O_131,N_2990,N_2968);
and UO_132 (O_132,N_2998,N_2983);
nor UO_133 (O_133,N_2980,N_2952);
xor UO_134 (O_134,N_2967,N_2980);
nand UO_135 (O_135,N_2990,N_2989);
or UO_136 (O_136,N_2958,N_2960);
nor UO_137 (O_137,N_2992,N_2952);
or UO_138 (O_138,N_2983,N_2976);
or UO_139 (O_139,N_2956,N_2993);
nand UO_140 (O_140,N_2970,N_2996);
and UO_141 (O_141,N_2958,N_2950);
and UO_142 (O_142,N_2993,N_2984);
or UO_143 (O_143,N_2966,N_2998);
and UO_144 (O_144,N_2989,N_2994);
and UO_145 (O_145,N_2989,N_2959);
xor UO_146 (O_146,N_2998,N_2993);
and UO_147 (O_147,N_2991,N_2992);
nand UO_148 (O_148,N_2985,N_2960);
nor UO_149 (O_149,N_2966,N_2960);
nor UO_150 (O_150,N_2973,N_2999);
and UO_151 (O_151,N_2961,N_2969);
or UO_152 (O_152,N_2996,N_2951);
xor UO_153 (O_153,N_2997,N_2965);
nor UO_154 (O_154,N_2992,N_2999);
and UO_155 (O_155,N_2961,N_2997);
nor UO_156 (O_156,N_2988,N_2977);
and UO_157 (O_157,N_2952,N_2969);
and UO_158 (O_158,N_2983,N_2957);
nor UO_159 (O_159,N_2977,N_2961);
nand UO_160 (O_160,N_2987,N_2953);
and UO_161 (O_161,N_2981,N_2997);
nand UO_162 (O_162,N_2957,N_2978);
nor UO_163 (O_163,N_2990,N_2977);
and UO_164 (O_164,N_2980,N_2992);
and UO_165 (O_165,N_2985,N_2995);
nor UO_166 (O_166,N_2966,N_2950);
and UO_167 (O_167,N_2956,N_2963);
and UO_168 (O_168,N_2963,N_2993);
or UO_169 (O_169,N_2983,N_2973);
nand UO_170 (O_170,N_2972,N_2966);
and UO_171 (O_171,N_2968,N_2984);
xnor UO_172 (O_172,N_2978,N_2973);
or UO_173 (O_173,N_2995,N_2974);
or UO_174 (O_174,N_2959,N_2951);
nand UO_175 (O_175,N_2997,N_2964);
or UO_176 (O_176,N_2968,N_2972);
and UO_177 (O_177,N_2965,N_2982);
or UO_178 (O_178,N_2985,N_2976);
xnor UO_179 (O_179,N_2984,N_2955);
nor UO_180 (O_180,N_2981,N_2993);
nand UO_181 (O_181,N_2964,N_2978);
nand UO_182 (O_182,N_2978,N_2965);
and UO_183 (O_183,N_2952,N_2988);
nand UO_184 (O_184,N_2994,N_2981);
or UO_185 (O_185,N_2972,N_2954);
nand UO_186 (O_186,N_2999,N_2951);
xnor UO_187 (O_187,N_2978,N_2982);
nor UO_188 (O_188,N_2957,N_2977);
and UO_189 (O_189,N_2973,N_2989);
nor UO_190 (O_190,N_2986,N_2989);
and UO_191 (O_191,N_2985,N_2951);
and UO_192 (O_192,N_2981,N_2970);
nand UO_193 (O_193,N_2964,N_2984);
or UO_194 (O_194,N_2969,N_2982);
xor UO_195 (O_195,N_2996,N_2973);
nand UO_196 (O_196,N_2961,N_2963);
or UO_197 (O_197,N_2959,N_2967);
or UO_198 (O_198,N_2976,N_2971);
xor UO_199 (O_199,N_2986,N_2967);
or UO_200 (O_200,N_2990,N_2991);
or UO_201 (O_201,N_2992,N_2975);
and UO_202 (O_202,N_2954,N_2967);
or UO_203 (O_203,N_2955,N_2973);
and UO_204 (O_204,N_2991,N_2982);
and UO_205 (O_205,N_2980,N_2961);
and UO_206 (O_206,N_2970,N_2955);
and UO_207 (O_207,N_2962,N_2969);
nand UO_208 (O_208,N_2953,N_2970);
nand UO_209 (O_209,N_2954,N_2991);
nand UO_210 (O_210,N_2967,N_2971);
xor UO_211 (O_211,N_2983,N_2974);
xor UO_212 (O_212,N_2992,N_2984);
nand UO_213 (O_213,N_2963,N_2998);
and UO_214 (O_214,N_2963,N_2992);
or UO_215 (O_215,N_2974,N_2975);
xor UO_216 (O_216,N_2979,N_2996);
nor UO_217 (O_217,N_2967,N_2972);
and UO_218 (O_218,N_2979,N_2960);
nand UO_219 (O_219,N_2979,N_2980);
nand UO_220 (O_220,N_2975,N_2998);
or UO_221 (O_221,N_2950,N_2982);
and UO_222 (O_222,N_2957,N_2990);
xor UO_223 (O_223,N_2972,N_2953);
and UO_224 (O_224,N_2985,N_2965);
nor UO_225 (O_225,N_2995,N_2956);
nor UO_226 (O_226,N_2968,N_2986);
nand UO_227 (O_227,N_2957,N_2979);
nor UO_228 (O_228,N_2981,N_2971);
or UO_229 (O_229,N_2962,N_2972);
or UO_230 (O_230,N_2974,N_2963);
or UO_231 (O_231,N_2959,N_2985);
and UO_232 (O_232,N_2964,N_2990);
or UO_233 (O_233,N_2975,N_2996);
nand UO_234 (O_234,N_2970,N_2963);
nand UO_235 (O_235,N_2969,N_2979);
nand UO_236 (O_236,N_2973,N_2974);
nor UO_237 (O_237,N_2993,N_2995);
xnor UO_238 (O_238,N_2993,N_2996);
and UO_239 (O_239,N_2976,N_2957);
xnor UO_240 (O_240,N_2987,N_2996);
and UO_241 (O_241,N_2952,N_2989);
nor UO_242 (O_242,N_2984,N_2967);
nor UO_243 (O_243,N_2991,N_2983);
and UO_244 (O_244,N_2971,N_2992);
xnor UO_245 (O_245,N_2966,N_2971);
or UO_246 (O_246,N_2955,N_2993);
nor UO_247 (O_247,N_2969,N_2953);
and UO_248 (O_248,N_2959,N_2987);
or UO_249 (O_249,N_2960,N_2991);
xnor UO_250 (O_250,N_2952,N_2970);
or UO_251 (O_251,N_2989,N_2991);
or UO_252 (O_252,N_2975,N_2967);
or UO_253 (O_253,N_2993,N_2986);
nand UO_254 (O_254,N_2980,N_2956);
and UO_255 (O_255,N_2997,N_2974);
and UO_256 (O_256,N_2986,N_2961);
and UO_257 (O_257,N_2977,N_2996);
or UO_258 (O_258,N_2952,N_2983);
nor UO_259 (O_259,N_2988,N_2987);
and UO_260 (O_260,N_2987,N_2981);
and UO_261 (O_261,N_2992,N_2966);
nand UO_262 (O_262,N_2997,N_2952);
nor UO_263 (O_263,N_2956,N_2981);
xnor UO_264 (O_264,N_2979,N_2958);
or UO_265 (O_265,N_2997,N_2962);
or UO_266 (O_266,N_2978,N_2972);
nor UO_267 (O_267,N_2962,N_2979);
or UO_268 (O_268,N_2971,N_2959);
nor UO_269 (O_269,N_2995,N_2964);
nor UO_270 (O_270,N_2958,N_2994);
and UO_271 (O_271,N_2964,N_2980);
or UO_272 (O_272,N_2968,N_2978);
nand UO_273 (O_273,N_2993,N_2988);
or UO_274 (O_274,N_2962,N_2967);
nand UO_275 (O_275,N_2985,N_2996);
xnor UO_276 (O_276,N_2988,N_2963);
or UO_277 (O_277,N_2959,N_2977);
and UO_278 (O_278,N_2963,N_2954);
nand UO_279 (O_279,N_2991,N_2967);
nor UO_280 (O_280,N_2977,N_2974);
nor UO_281 (O_281,N_2962,N_2986);
xor UO_282 (O_282,N_2952,N_2995);
or UO_283 (O_283,N_2987,N_2972);
or UO_284 (O_284,N_2981,N_2991);
nor UO_285 (O_285,N_2965,N_2954);
nand UO_286 (O_286,N_2952,N_2981);
nand UO_287 (O_287,N_2973,N_2971);
or UO_288 (O_288,N_2970,N_2976);
xor UO_289 (O_289,N_2971,N_2979);
nor UO_290 (O_290,N_2991,N_2972);
nor UO_291 (O_291,N_2988,N_2964);
and UO_292 (O_292,N_2960,N_2978);
and UO_293 (O_293,N_2975,N_2954);
and UO_294 (O_294,N_2989,N_2950);
nand UO_295 (O_295,N_2993,N_2976);
nand UO_296 (O_296,N_2965,N_2958);
nor UO_297 (O_297,N_2953,N_2961);
or UO_298 (O_298,N_2969,N_2997);
nand UO_299 (O_299,N_2968,N_2979);
nor UO_300 (O_300,N_2965,N_2959);
nand UO_301 (O_301,N_2965,N_2962);
and UO_302 (O_302,N_2968,N_2965);
and UO_303 (O_303,N_2973,N_2995);
nand UO_304 (O_304,N_2969,N_2951);
nor UO_305 (O_305,N_2986,N_2959);
xnor UO_306 (O_306,N_2978,N_2954);
nor UO_307 (O_307,N_2998,N_2980);
nor UO_308 (O_308,N_2967,N_2963);
nor UO_309 (O_309,N_2995,N_2957);
xnor UO_310 (O_310,N_2996,N_2965);
nand UO_311 (O_311,N_2990,N_2985);
nand UO_312 (O_312,N_2974,N_2955);
or UO_313 (O_313,N_2998,N_2992);
or UO_314 (O_314,N_2971,N_2987);
nor UO_315 (O_315,N_2966,N_2959);
and UO_316 (O_316,N_2970,N_2991);
nand UO_317 (O_317,N_2975,N_2986);
and UO_318 (O_318,N_2977,N_2984);
xnor UO_319 (O_319,N_2950,N_2984);
nand UO_320 (O_320,N_2987,N_2954);
and UO_321 (O_321,N_2969,N_2988);
and UO_322 (O_322,N_2956,N_2959);
and UO_323 (O_323,N_2966,N_2979);
nor UO_324 (O_324,N_2977,N_2972);
or UO_325 (O_325,N_2973,N_2986);
nand UO_326 (O_326,N_2973,N_2960);
nand UO_327 (O_327,N_2954,N_2986);
and UO_328 (O_328,N_2970,N_2971);
and UO_329 (O_329,N_2961,N_2990);
or UO_330 (O_330,N_2957,N_2992);
and UO_331 (O_331,N_2957,N_2973);
nand UO_332 (O_332,N_2956,N_2990);
nand UO_333 (O_333,N_2986,N_2979);
and UO_334 (O_334,N_2994,N_2990);
or UO_335 (O_335,N_2994,N_2988);
or UO_336 (O_336,N_2958,N_2951);
nor UO_337 (O_337,N_2991,N_2950);
nand UO_338 (O_338,N_2968,N_2981);
and UO_339 (O_339,N_2992,N_2964);
xnor UO_340 (O_340,N_2990,N_2950);
or UO_341 (O_341,N_2954,N_2984);
nand UO_342 (O_342,N_2992,N_2954);
and UO_343 (O_343,N_2976,N_2950);
and UO_344 (O_344,N_2991,N_2980);
xor UO_345 (O_345,N_2954,N_2979);
nor UO_346 (O_346,N_2981,N_2979);
and UO_347 (O_347,N_2974,N_2951);
or UO_348 (O_348,N_2984,N_2979);
nand UO_349 (O_349,N_2987,N_2952);
nor UO_350 (O_350,N_2963,N_2981);
and UO_351 (O_351,N_2998,N_2996);
and UO_352 (O_352,N_2977,N_2986);
or UO_353 (O_353,N_2996,N_2994);
nand UO_354 (O_354,N_2967,N_2976);
or UO_355 (O_355,N_2962,N_2957);
nor UO_356 (O_356,N_2999,N_2996);
or UO_357 (O_357,N_2960,N_2981);
nor UO_358 (O_358,N_2996,N_2981);
nor UO_359 (O_359,N_2975,N_2952);
nor UO_360 (O_360,N_2970,N_2993);
nor UO_361 (O_361,N_2987,N_2976);
xnor UO_362 (O_362,N_2972,N_2999);
nand UO_363 (O_363,N_2973,N_2975);
nand UO_364 (O_364,N_2964,N_2950);
nand UO_365 (O_365,N_2958,N_2996);
or UO_366 (O_366,N_2982,N_2971);
nand UO_367 (O_367,N_2985,N_2999);
and UO_368 (O_368,N_2980,N_2954);
or UO_369 (O_369,N_2964,N_2982);
nand UO_370 (O_370,N_2997,N_2987);
and UO_371 (O_371,N_2951,N_2986);
nor UO_372 (O_372,N_2987,N_2951);
xnor UO_373 (O_373,N_2976,N_2966);
nor UO_374 (O_374,N_2971,N_2951);
or UO_375 (O_375,N_2982,N_2998);
and UO_376 (O_376,N_2989,N_2961);
or UO_377 (O_377,N_2992,N_2977);
xor UO_378 (O_378,N_2978,N_2971);
nand UO_379 (O_379,N_2975,N_2983);
xor UO_380 (O_380,N_2982,N_2975);
or UO_381 (O_381,N_2965,N_2957);
xnor UO_382 (O_382,N_2982,N_2953);
nand UO_383 (O_383,N_2985,N_2980);
nand UO_384 (O_384,N_2965,N_2970);
nand UO_385 (O_385,N_2958,N_2991);
and UO_386 (O_386,N_2994,N_2987);
or UO_387 (O_387,N_2971,N_2972);
and UO_388 (O_388,N_2985,N_2987);
and UO_389 (O_389,N_2979,N_2998);
nor UO_390 (O_390,N_2997,N_2958);
nor UO_391 (O_391,N_2964,N_2959);
or UO_392 (O_392,N_2987,N_2966);
nand UO_393 (O_393,N_2997,N_2991);
nor UO_394 (O_394,N_2970,N_2973);
xnor UO_395 (O_395,N_2966,N_2958);
or UO_396 (O_396,N_2957,N_2984);
nand UO_397 (O_397,N_2964,N_2955);
or UO_398 (O_398,N_2996,N_2991);
nor UO_399 (O_399,N_2990,N_2981);
and UO_400 (O_400,N_2969,N_2967);
nor UO_401 (O_401,N_2962,N_2992);
nand UO_402 (O_402,N_2975,N_2972);
or UO_403 (O_403,N_2995,N_2959);
nor UO_404 (O_404,N_2982,N_2984);
and UO_405 (O_405,N_2955,N_2976);
nor UO_406 (O_406,N_2963,N_2969);
nand UO_407 (O_407,N_2954,N_2976);
and UO_408 (O_408,N_2968,N_2999);
nor UO_409 (O_409,N_2956,N_2997);
and UO_410 (O_410,N_2970,N_2984);
nor UO_411 (O_411,N_2989,N_2997);
xnor UO_412 (O_412,N_2971,N_2994);
and UO_413 (O_413,N_2975,N_2964);
and UO_414 (O_414,N_2977,N_2971);
nor UO_415 (O_415,N_2950,N_2959);
or UO_416 (O_416,N_2966,N_2984);
and UO_417 (O_417,N_2980,N_2983);
and UO_418 (O_418,N_2956,N_2978);
and UO_419 (O_419,N_2964,N_2951);
and UO_420 (O_420,N_2995,N_2981);
or UO_421 (O_421,N_2999,N_2962);
nand UO_422 (O_422,N_2988,N_2998);
and UO_423 (O_423,N_2978,N_2969);
and UO_424 (O_424,N_2996,N_2995);
nand UO_425 (O_425,N_2970,N_2950);
or UO_426 (O_426,N_2983,N_2978);
or UO_427 (O_427,N_2999,N_2965);
or UO_428 (O_428,N_2955,N_2952);
nand UO_429 (O_429,N_2998,N_2957);
nor UO_430 (O_430,N_2992,N_2982);
and UO_431 (O_431,N_2960,N_2963);
and UO_432 (O_432,N_2983,N_2981);
nand UO_433 (O_433,N_2997,N_2983);
nand UO_434 (O_434,N_2953,N_2989);
and UO_435 (O_435,N_2974,N_2990);
or UO_436 (O_436,N_2993,N_2999);
nor UO_437 (O_437,N_2970,N_2983);
or UO_438 (O_438,N_2979,N_2972);
and UO_439 (O_439,N_2984,N_2961);
xor UO_440 (O_440,N_2991,N_2969);
nand UO_441 (O_441,N_2972,N_2992);
nand UO_442 (O_442,N_2996,N_2961);
or UO_443 (O_443,N_2960,N_2970);
or UO_444 (O_444,N_2963,N_2995);
xor UO_445 (O_445,N_2998,N_2951);
nor UO_446 (O_446,N_2998,N_2961);
and UO_447 (O_447,N_2953,N_2975);
and UO_448 (O_448,N_2964,N_2979);
and UO_449 (O_449,N_2962,N_2995);
or UO_450 (O_450,N_2999,N_2983);
nor UO_451 (O_451,N_2977,N_2991);
or UO_452 (O_452,N_2967,N_2951);
or UO_453 (O_453,N_2973,N_2987);
nand UO_454 (O_454,N_2960,N_2968);
xor UO_455 (O_455,N_2977,N_2958);
nor UO_456 (O_456,N_2996,N_2980);
or UO_457 (O_457,N_2969,N_2958);
and UO_458 (O_458,N_2974,N_2988);
and UO_459 (O_459,N_2993,N_2982);
nand UO_460 (O_460,N_2960,N_2965);
and UO_461 (O_461,N_2951,N_2966);
nand UO_462 (O_462,N_2988,N_2990);
or UO_463 (O_463,N_2952,N_2979);
and UO_464 (O_464,N_2950,N_2978);
nor UO_465 (O_465,N_2981,N_2984);
nor UO_466 (O_466,N_2985,N_2955);
nand UO_467 (O_467,N_2967,N_2968);
nand UO_468 (O_468,N_2994,N_2991);
nor UO_469 (O_469,N_2952,N_2974);
or UO_470 (O_470,N_2970,N_2998);
and UO_471 (O_471,N_2996,N_2955);
nand UO_472 (O_472,N_2979,N_2999);
nand UO_473 (O_473,N_2972,N_2981);
and UO_474 (O_474,N_2963,N_2953);
or UO_475 (O_475,N_2967,N_2989);
nand UO_476 (O_476,N_2984,N_2960);
or UO_477 (O_477,N_2976,N_2965);
nand UO_478 (O_478,N_2998,N_2984);
and UO_479 (O_479,N_2968,N_2980);
and UO_480 (O_480,N_2979,N_2982);
or UO_481 (O_481,N_2989,N_2965);
nand UO_482 (O_482,N_2996,N_2984);
xnor UO_483 (O_483,N_2973,N_2994);
or UO_484 (O_484,N_2950,N_2954);
and UO_485 (O_485,N_2980,N_2993);
nand UO_486 (O_486,N_2964,N_2962);
nor UO_487 (O_487,N_2999,N_2971);
nand UO_488 (O_488,N_2973,N_2956);
nand UO_489 (O_489,N_2982,N_2958);
nand UO_490 (O_490,N_2968,N_2966);
or UO_491 (O_491,N_2957,N_2960);
or UO_492 (O_492,N_2972,N_2986);
nor UO_493 (O_493,N_2953,N_2995);
and UO_494 (O_494,N_2969,N_2983);
or UO_495 (O_495,N_2980,N_2962);
and UO_496 (O_496,N_2964,N_2956);
or UO_497 (O_497,N_2978,N_2999);
or UO_498 (O_498,N_2976,N_2979);
nor UO_499 (O_499,N_2952,N_2958);
endmodule