module basic_2000_20000_2500_50_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_125,In_1529);
xor U1 (N_1,In_830,In_77);
nand U2 (N_2,In_528,In_513);
or U3 (N_3,In_835,In_310);
xnor U4 (N_4,In_1572,In_283);
xor U5 (N_5,In_1696,In_906);
nand U6 (N_6,In_1632,In_1087);
nand U7 (N_7,In_1278,In_858);
and U8 (N_8,In_862,In_1579);
and U9 (N_9,In_1584,In_475);
xor U10 (N_10,In_1850,In_1937);
and U11 (N_11,In_1586,In_1780);
xnor U12 (N_12,In_198,In_1117);
nor U13 (N_13,In_326,In_1428);
nor U14 (N_14,In_437,In_892);
and U15 (N_15,In_1980,In_1309);
or U16 (N_16,In_760,In_399);
nand U17 (N_17,In_1897,In_1982);
and U18 (N_18,In_1465,In_932);
nand U19 (N_19,In_112,In_1744);
or U20 (N_20,In_1438,In_618);
and U21 (N_21,In_903,In_424);
nand U22 (N_22,In_130,In_378);
and U23 (N_23,In_246,In_1211);
and U24 (N_24,In_37,In_694);
nor U25 (N_25,In_572,In_749);
and U26 (N_26,In_1967,In_490);
xor U27 (N_27,In_361,In_1292);
nand U28 (N_28,In_1155,In_730);
xor U29 (N_29,In_1644,In_967);
xnor U30 (N_30,In_466,In_408);
or U31 (N_31,In_190,In_1437);
or U32 (N_32,In_1760,In_1506);
or U33 (N_33,In_1607,In_943);
xnor U34 (N_34,In_1197,In_1416);
and U35 (N_35,In_761,In_822);
nor U36 (N_36,In_365,In_1302);
or U37 (N_37,In_1731,In_1135);
xor U38 (N_38,In_36,In_131);
and U39 (N_39,In_956,In_1362);
nor U40 (N_40,In_1468,In_15);
or U41 (N_41,In_734,In_1993);
xor U42 (N_42,In_1386,In_1985);
and U43 (N_43,In_1119,In_419);
nand U44 (N_44,In_1355,In_260);
and U45 (N_45,In_1422,In_281);
or U46 (N_46,In_599,In_679);
xor U47 (N_47,In_1611,In_1411);
nor U48 (N_48,In_232,In_1409);
and U49 (N_49,In_1886,In_651);
nand U50 (N_50,In_442,In_1589);
xnor U51 (N_51,In_1866,In_733);
xor U52 (N_52,In_1233,In_810);
nand U53 (N_53,In_1005,In_295);
or U54 (N_54,In_1681,In_1374);
or U55 (N_55,In_499,In_481);
xor U56 (N_56,In_1766,In_1826);
nor U57 (N_57,In_1732,In_1845);
or U58 (N_58,In_1306,In_620);
and U59 (N_59,In_1481,In_495);
nand U60 (N_60,In_71,In_1380);
nor U61 (N_61,In_409,In_316);
or U62 (N_62,In_39,In_1577);
nor U63 (N_63,In_1040,In_1361);
or U64 (N_64,In_1771,In_1829);
or U65 (N_65,In_1467,In_177);
or U66 (N_66,In_1175,In_1718);
nand U67 (N_67,In_706,In_879);
nor U68 (N_68,In_1103,In_287);
nand U69 (N_69,In_160,In_547);
xnor U70 (N_70,In_24,In_1665);
and U71 (N_71,In_300,In_476);
and U72 (N_72,In_17,In_28);
xnor U73 (N_73,In_537,In_874);
and U74 (N_74,In_1132,In_55);
or U75 (N_75,In_649,In_1401);
and U76 (N_76,In_1170,In_1657);
and U77 (N_77,In_1446,In_253);
nand U78 (N_78,In_1196,In_1171);
nand U79 (N_79,In_1253,In_1252);
nor U80 (N_80,In_1613,In_109);
nand U81 (N_81,In_431,In_617);
nor U82 (N_82,In_1851,In_303);
or U83 (N_83,In_1999,In_1311);
or U84 (N_84,In_970,In_257);
and U85 (N_85,In_477,In_1041);
and U86 (N_86,In_472,In_918);
or U87 (N_87,In_1182,In_1493);
nor U88 (N_88,In_823,In_1646);
nand U89 (N_89,In_355,In_1935);
nand U90 (N_90,In_1963,In_85);
nor U91 (N_91,In_802,In_995);
nand U92 (N_92,In_1090,In_594);
nand U93 (N_93,In_697,In_615);
nor U94 (N_94,In_1367,In_1214);
nor U95 (N_95,In_610,In_1026);
and U96 (N_96,In_1046,In_924);
and U97 (N_97,In_702,In_1460);
and U98 (N_98,In_1693,In_645);
or U99 (N_99,In_541,In_1178);
xnor U100 (N_100,In_33,In_1803);
xor U101 (N_101,In_840,In_1535);
nand U102 (N_102,In_359,In_781);
nor U103 (N_103,In_348,In_1787);
nand U104 (N_104,In_1838,In_1740);
nor U105 (N_105,In_167,In_740);
nor U106 (N_106,In_330,In_13);
nand U107 (N_107,In_241,In_855);
nor U108 (N_108,In_1501,In_1141);
nand U109 (N_109,In_843,In_341);
xor U110 (N_110,In_1741,In_1686);
and U111 (N_111,In_1562,In_342);
or U112 (N_112,In_80,In_356);
nand U113 (N_113,In_363,In_1753);
or U114 (N_114,In_1847,In_1316);
xnor U115 (N_115,In_1247,In_380);
and U116 (N_116,In_1218,In_1398);
or U117 (N_117,In_1708,In_542);
nor U118 (N_118,In_1588,In_911);
or U119 (N_119,In_517,In_1350);
nand U120 (N_120,In_589,In_1720);
nand U121 (N_121,In_975,In_1615);
and U122 (N_122,In_423,In_1463);
nor U123 (N_123,In_974,In_1516);
or U124 (N_124,In_1234,In_1342);
and U125 (N_125,In_1814,In_159);
or U126 (N_126,In_169,In_1358);
nand U127 (N_127,In_62,In_1183);
nand U128 (N_128,In_1599,In_1840);
or U129 (N_129,In_165,In_1348);
or U130 (N_130,In_385,In_1415);
or U131 (N_131,In_779,In_44);
nand U132 (N_132,In_338,In_1654);
and U133 (N_133,In_1899,In_57);
nand U134 (N_134,In_444,In_1142);
and U135 (N_135,In_1507,In_1448);
nand U136 (N_136,In_1689,In_535);
nand U137 (N_137,In_1420,In_1271);
or U138 (N_138,In_1491,In_1734);
nor U139 (N_139,In_1834,In_1921);
xor U140 (N_140,In_171,In_1435);
nand U141 (N_141,In_1076,In_1541);
xor U142 (N_142,In_1106,In_878);
and U143 (N_143,In_521,In_1860);
or U144 (N_144,In_1048,In_628);
or U145 (N_145,In_1251,In_1531);
and U146 (N_146,In_433,In_392);
and U147 (N_147,In_1578,In_1620);
nand U148 (N_148,In_1407,In_581);
or U149 (N_149,In_337,In_1939);
or U150 (N_150,In_755,In_496);
nor U151 (N_151,In_1173,In_1598);
nor U152 (N_152,In_820,In_153);
or U153 (N_153,In_895,In_211);
nand U154 (N_154,In_1502,In_1757);
xnor U155 (N_155,In_681,In_1763);
and U156 (N_156,In_939,In_529);
nand U157 (N_157,In_1167,In_1496);
and U158 (N_158,In_902,In_1893);
nand U159 (N_159,In_1489,In_482);
nand U160 (N_160,In_233,In_208);
and U161 (N_161,In_884,In_1261);
xor U162 (N_162,In_1272,In_212);
xnor U163 (N_163,In_1210,In_262);
nand U164 (N_164,In_880,In_1239);
and U165 (N_165,In_61,In_1185);
xor U166 (N_166,In_391,In_514);
or U167 (N_167,In_1494,In_1205);
or U168 (N_168,In_248,In_909);
nor U169 (N_169,In_523,In_1928);
or U170 (N_170,In_657,In_888);
nand U171 (N_171,In_1984,In_844);
nand U172 (N_172,In_789,In_1610);
or U173 (N_173,In_1756,In_1244);
nor U174 (N_174,In_806,In_1277);
and U175 (N_175,In_546,In_1536);
xnor U176 (N_176,In_123,In_435);
or U177 (N_177,In_427,In_519);
nor U178 (N_178,In_1429,In_1102);
and U179 (N_179,In_1621,In_1474);
nand U180 (N_180,In_1129,In_331);
and U181 (N_181,In_1749,In_1545);
and U182 (N_182,In_564,In_1052);
and U183 (N_183,In_114,In_1458);
and U184 (N_184,In_1349,In_3);
and U185 (N_185,In_750,In_268);
nand U186 (N_186,In_440,In_1525);
or U187 (N_187,In_282,In_604);
nand U188 (N_188,In_309,In_774);
nor U189 (N_189,In_1554,In_1330);
or U190 (N_190,In_1835,In_1037);
and U191 (N_191,In_1235,In_30);
nand U192 (N_192,In_113,In_473);
xor U193 (N_193,In_415,In_711);
xor U194 (N_194,In_86,In_721);
nand U195 (N_195,In_307,In_118);
nand U196 (N_196,In_1558,In_966);
xor U197 (N_197,In_816,In_1553);
and U198 (N_198,In_221,In_983);
or U199 (N_199,In_1518,In_543);
nand U200 (N_200,In_1697,In_197);
xor U201 (N_201,In_1109,In_1294);
xor U202 (N_202,In_1034,In_782);
and U203 (N_203,In_658,In_91);
nor U204 (N_204,In_1122,In_72);
xor U205 (N_205,In_460,In_20);
xor U206 (N_206,In_1890,In_1807);
nand U207 (N_207,In_1371,In_201);
and U208 (N_208,In_454,In_1013);
xor U209 (N_209,In_596,In_797);
nor U210 (N_210,In_941,In_10);
xor U211 (N_211,In_531,In_1867);
or U212 (N_212,In_695,In_9);
nand U213 (N_213,In_381,In_92);
nand U214 (N_214,In_1637,In_1120);
and U215 (N_215,In_560,In_947);
and U216 (N_216,In_1707,In_1432);
xor U217 (N_217,In_1955,In_582);
xnor U218 (N_218,In_1878,In_1922);
nor U219 (N_219,In_478,In_1100);
nand U220 (N_220,In_1715,In_1776);
and U221 (N_221,In_11,In_120);
xor U222 (N_222,In_1476,In_162);
nand U223 (N_223,In_905,In_25);
nand U224 (N_224,In_1791,In_1022);
nor U225 (N_225,In_1816,In_1056);
or U226 (N_226,In_1759,In_677);
or U227 (N_227,In_1376,In_124);
nand U228 (N_228,In_718,In_16);
and U229 (N_229,In_961,In_1324);
xnor U230 (N_230,In_1488,In_522);
or U231 (N_231,In_642,In_981);
or U232 (N_232,In_1616,In_989);
and U233 (N_233,In_545,In_1439);
and U234 (N_234,In_1364,In_1224);
nor U235 (N_235,In_1550,In_405);
nand U236 (N_236,In_207,In_1849);
xnor U237 (N_237,In_1369,In_1169);
or U238 (N_238,In_856,In_1743);
xor U239 (N_239,In_1671,In_1390);
and U240 (N_240,In_978,In_999);
and U241 (N_241,In_1914,In_687);
and U242 (N_242,In_374,In_1569);
xnor U243 (N_243,In_51,In_1652);
nor U244 (N_244,In_673,In_1334);
nand U245 (N_245,In_728,In_402);
xnor U246 (N_246,In_353,In_1282);
nor U247 (N_247,In_461,In_705);
or U248 (N_248,In_686,In_1781);
nor U249 (N_249,In_881,In_1910);
nand U250 (N_250,In_296,In_1746);
nand U251 (N_251,In_1846,In_189);
xor U252 (N_252,In_1470,In_573);
or U253 (N_253,In_52,In_1168);
xnor U254 (N_254,In_222,In_1918);
xnor U255 (N_255,In_1130,In_867);
or U256 (N_256,In_1118,In_1951);
nor U257 (N_257,In_847,In_1965);
and U258 (N_258,In_271,In_824);
and U259 (N_259,In_1735,In_135);
or U260 (N_260,In_653,In_921);
xnor U261 (N_261,In_58,In_266);
or U262 (N_262,In_629,In_1012);
xnor U263 (N_263,In_1755,In_950);
nand U264 (N_264,In_137,In_1571);
or U265 (N_265,In_1023,In_647);
nor U266 (N_266,In_891,In_945);
or U267 (N_267,In_636,In_915);
xnor U268 (N_268,In_1357,In_1243);
xor U269 (N_269,In_1062,In_877);
and U270 (N_270,In_486,In_491);
or U271 (N_271,In_1209,In_436);
nand U272 (N_272,In_1971,In_904);
or U273 (N_273,In_870,In_1279);
xnor U274 (N_274,In_1312,In_848);
xnor U275 (N_275,In_1642,In_1523);
or U276 (N_276,In_723,In_1232);
nor U277 (N_277,In_1704,In_846);
nor U278 (N_278,In_787,In_149);
and U279 (N_279,In_247,In_1956);
or U280 (N_280,In_1412,In_1815);
nor U281 (N_281,In_1901,In_108);
and U282 (N_282,In_333,In_682);
or U283 (N_283,In_462,In_994);
nor U284 (N_284,In_41,In_621);
or U285 (N_285,In_1139,In_1112);
and U286 (N_286,In_930,In_1841);
xor U287 (N_287,In_1275,In_413);
and U288 (N_288,In_725,In_1166);
nand U289 (N_289,In_968,In_140);
nor U290 (N_290,In_1727,In_364);
nand U291 (N_291,In_641,In_231);
and U292 (N_292,In_676,In_347);
and U293 (N_293,In_731,In_116);
or U294 (N_294,In_1952,In_141);
nor U295 (N_295,In_1177,In_1811);
or U296 (N_296,In_1079,In_1363);
or U297 (N_297,In_1832,In_554);
nand U298 (N_298,In_747,In_898);
nand U299 (N_299,In_258,In_1549);
or U300 (N_300,In_14,In_1500);
nand U301 (N_301,In_1674,In_1464);
nand U302 (N_302,In_456,In_626);
xnor U303 (N_303,In_1286,In_1931);
and U304 (N_304,In_900,In_1195);
and U305 (N_305,In_1942,In_758);
and U306 (N_306,In_1709,In_1336);
nand U307 (N_307,In_1086,In_837);
and U308 (N_308,In_1146,In_259);
or U309 (N_309,In_1843,In_97);
nor U310 (N_310,In_771,In_1695);
nor U311 (N_311,In_1977,In_1888);
nor U312 (N_312,In_1938,In_325);
or U313 (N_313,In_1069,In_948);
nor U314 (N_314,In_1149,In_1246);
nand U315 (N_315,In_1020,In_783);
and U316 (N_316,In_1736,In_969);
and U317 (N_317,In_1094,In_1485);
nor U318 (N_318,In_1303,In_1359);
nor U319 (N_319,In_193,In_289);
or U320 (N_320,In_288,In_390);
and U321 (N_321,In_147,In_954);
xnor U322 (N_322,In_26,In_0);
or U323 (N_323,In_412,In_1031);
or U324 (N_324,In_1403,In_1212);
nand U325 (N_325,In_1213,In_446);
nor U326 (N_326,In_1869,In_1783);
xor U327 (N_327,In_611,In_1080);
nand U328 (N_328,In_1260,In_619);
nand U329 (N_329,In_996,In_154);
or U330 (N_330,In_622,In_1471);
or U331 (N_331,In_990,In_1307);
and U332 (N_332,In_314,In_1713);
nand U333 (N_333,In_1511,In_1539);
and U334 (N_334,In_1907,In_205);
xnor U335 (N_335,In_143,In_1961);
nand U336 (N_336,In_1388,In_1236);
and U337 (N_337,In_1634,In_1199);
or U338 (N_338,In_386,In_1091);
xnor U339 (N_339,In_766,In_850);
xnor U340 (N_340,In_865,In_1104);
nor U341 (N_341,In_1974,In_21);
and U342 (N_342,In_410,In_685);
and U343 (N_343,In_1830,In_1478);
nand U344 (N_344,In_592,In_317);
xnor U345 (N_345,In_1131,In_172);
or U346 (N_346,In_242,In_1773);
and U347 (N_347,In_194,In_1378);
xor U348 (N_348,In_261,In_196);
or U349 (N_349,In_95,In_1839);
nand U350 (N_350,In_469,In_1902);
nand U351 (N_351,In_204,In_777);
nand U352 (N_352,In_767,In_1114);
nor U353 (N_353,In_971,In_949);
xor U354 (N_354,In_45,In_1819);
nor U355 (N_355,In_1200,In_1524);
xor U356 (N_356,In_959,In_1556);
nand U357 (N_357,In_1870,In_1095);
nand U358 (N_358,In_393,In_1221);
and U359 (N_359,In_588,In_370);
and U360 (N_360,In_689,In_1084);
and U361 (N_361,In_1635,In_1134);
nand U362 (N_362,In_857,In_1987);
nor U363 (N_363,In_1580,In_1770);
xnor U364 (N_364,In_19,In_1626);
nand U365 (N_365,In_605,In_530);
xor U366 (N_366,In_576,In_1414);
nand U367 (N_367,In_265,In_1038);
or U368 (N_368,In_133,In_1677);
nand U369 (N_369,In_226,In_1053);
and U370 (N_370,In_1721,In_650);
or U371 (N_371,In_826,In_744);
and U372 (N_372,In_1190,In_866);
xnor U373 (N_373,In_1662,In_1750);
nand U374 (N_374,In_668,In_1944);
and U375 (N_375,In_1601,In_1653);
and U376 (N_376,In_276,In_1029);
or U377 (N_377,In_1399,In_1394);
nor U378 (N_378,In_1565,In_346);
or U379 (N_379,In_1219,In_34);
or U380 (N_380,In_1447,In_1220);
and U381 (N_381,In_128,In_663);
xnor U382 (N_382,In_164,In_773);
or U383 (N_383,In_1176,In_1868);
and U384 (N_384,In_1801,In_1612);
xor U385 (N_385,In_644,In_304);
nor U386 (N_386,In_591,In_285);
xor U387 (N_387,In_1490,In_748);
or U388 (N_388,In_1421,In_631);
xnor U389 (N_389,In_400,In_1875);
nand U390 (N_390,In_666,In_578);
xnor U391 (N_391,In_175,In_1010);
xor U392 (N_392,In_1527,In_1014);
or U393 (N_393,In_1650,In_1794);
nor U394 (N_394,In_1136,In_312);
nor U395 (N_395,In_1881,In_503);
nand U396 (N_396,In_1331,In_1699);
and U397 (N_397,In_1994,In_1649);
and U398 (N_398,In_6,In_506);
or U399 (N_399,In_351,In_1934);
and U400 (N_400,In_814,N_251);
or U401 (N_401,In_1949,N_204);
xnor U402 (N_402,In_349,In_1258);
nor U403 (N_403,In_1154,In_786);
xor U404 (N_404,In_1582,In_665);
nor U405 (N_405,In_1975,In_953);
xor U406 (N_406,In_237,N_49);
nand U407 (N_407,In_813,In_350);
xor U408 (N_408,In_1360,N_317);
or U409 (N_409,N_30,N_324);
nand U410 (N_410,In_1152,In_1824);
nor U411 (N_411,In_920,In_606);
nor U412 (N_412,N_391,In_321);
nor U413 (N_413,In_267,In_1655);
nand U414 (N_414,In_1692,N_91);
and U415 (N_415,In_1365,N_309);
or U416 (N_416,N_399,In_1730);
and U417 (N_417,In_507,N_283);
xnor U418 (N_418,In_827,In_1701);
or U419 (N_419,In_1528,In_1017);
or U420 (N_420,In_864,In_1647);
xnor U421 (N_421,N_54,In_195);
nor U422 (N_422,In_674,In_1594);
nor U423 (N_423,N_332,In_65);
nand U424 (N_424,In_883,In_1690);
nor U425 (N_425,N_295,In_1267);
and U426 (N_426,In_1786,In_1552);
or U427 (N_427,In_1717,In_168);
and U428 (N_428,In_73,In_639);
nor U429 (N_429,In_1186,In_1784);
nor U430 (N_430,In_940,N_296);
nor U431 (N_431,N_189,In_518);
nand U432 (N_432,In_1680,N_242);
nor U433 (N_433,In_121,N_249);
or U434 (N_434,N_174,In_717);
nor U435 (N_435,In_1051,In_1078);
and U436 (N_436,In_1187,N_207);
nand U437 (N_437,In_79,N_142);
nand U438 (N_438,In_1973,In_291);
xor U439 (N_439,In_464,N_387);
nand U440 (N_440,In_1329,In_534);
nand U441 (N_441,In_586,In_429);
nor U442 (N_442,In_1992,In_148);
nor U443 (N_443,N_282,In_151);
nand U444 (N_444,In_1706,In_1593);
nor U445 (N_445,In_1225,In_320);
and U446 (N_446,In_142,In_1273);
nor U447 (N_447,In_1544,In_1263);
xor U448 (N_448,N_2,N_308);
and U449 (N_449,In_377,In_914);
or U450 (N_450,In_700,In_957);
or U451 (N_451,In_286,N_259);
or U452 (N_452,In_1033,In_759);
nand U453 (N_453,N_240,In_245);
xor U454 (N_454,In_1248,N_335);
nor U455 (N_455,N_197,In_1011);
and U456 (N_456,In_1499,N_378);
or U457 (N_457,In_101,In_1855);
nand U458 (N_458,In_1879,In_255);
nand U459 (N_459,In_1676,N_325);
xnor U460 (N_460,In_1002,N_40);
nor U461 (N_461,In_1898,In_1284);
nand U462 (N_462,In_818,In_1018);
nand U463 (N_463,In_780,N_150);
and U464 (N_464,In_1664,In_1323);
or U465 (N_465,In_1274,In_1315);
or U466 (N_466,In_775,N_320);
or U467 (N_467,In_1895,In_1366);
xor U468 (N_468,N_24,In_812);
nand U469 (N_469,In_551,In_691);
and U470 (N_470,In_1058,N_173);
nand U471 (N_471,N_149,In_1833);
and U472 (N_472,N_247,In_512);
or U473 (N_473,In_1976,N_115);
or U474 (N_474,In_1449,N_58);
and U475 (N_475,In_1916,N_107);
or U476 (N_476,In_1920,In_178);
nor U477 (N_477,In_751,In_693);
and U478 (N_478,N_6,In_368);
nand U479 (N_479,N_17,In_982);
or U480 (N_480,In_4,In_992);
and U481 (N_481,In_188,In_1392);
or U482 (N_482,In_703,In_1148);
and U483 (N_483,In_1368,N_201);
or U484 (N_484,In_709,N_31);
or U485 (N_485,In_1405,N_342);
nor U486 (N_486,In_669,In_479);
nand U487 (N_487,In_887,In_318);
xnor U488 (N_488,In_516,In_106);
nand U489 (N_489,In_933,N_18);
nand U490 (N_490,In_185,In_269);
nand U491 (N_491,N_127,N_101);
xor U492 (N_492,In_93,N_57);
or U493 (N_493,In_707,In_483);
nand U494 (N_494,N_111,In_157);
or U495 (N_495,In_1030,In_280);
or U496 (N_496,In_1997,In_1540);
or U497 (N_497,In_1848,N_108);
xnor U498 (N_498,In_984,In_1758);
and U499 (N_499,In_1754,In_1473);
or U500 (N_500,In_161,N_228);
or U501 (N_501,In_1008,N_160);
nand U502 (N_502,In_1059,In_1061);
and U503 (N_503,In_614,In_1070);
nor U504 (N_504,In_1472,In_1687);
nor U505 (N_505,In_1877,In_593);
or U506 (N_506,N_106,In_497);
xor U507 (N_507,In_1067,In_53);
and U508 (N_508,N_53,In_1747);
nor U509 (N_509,In_1861,In_1633);
nor U510 (N_510,N_66,In_216);
or U511 (N_511,N_80,In_384);
or U512 (N_512,In_234,N_10);
or U513 (N_513,In_389,In_293);
and U514 (N_514,In_1133,In_449);
xor U515 (N_515,In_1858,In_1228);
nor U516 (N_516,In_1085,In_1081);
and U517 (N_517,N_215,N_81);
xor U518 (N_518,In_1308,In_1515);
nand U519 (N_519,In_986,In_1822);
nor U520 (N_520,In_696,In_821);
nand U521 (N_521,In_407,In_1560);
or U522 (N_522,In_1180,N_141);
or U523 (N_523,N_77,N_181);
nand U524 (N_524,In_1852,In_1291);
nand U525 (N_525,In_358,N_323);
nor U526 (N_526,In_1285,In_63);
nor U527 (N_527,N_70,In_1636);
nand U528 (N_528,In_1150,In_754);
xor U529 (N_529,N_148,In_463);
nor U530 (N_530,In_963,In_1505);
nor U531 (N_531,In_1343,In_568);
or U532 (N_532,N_370,N_95);
or U533 (N_533,N_102,In_680);
nand U534 (N_534,N_63,In_230);
nor U535 (N_535,In_166,N_263);
nor U536 (N_536,In_343,In_583);
and U537 (N_537,In_1,In_1418);
xnor U538 (N_538,In_1618,In_1156);
and U539 (N_539,In_158,In_1887);
nand U540 (N_540,In_652,N_365);
xor U541 (N_541,In_646,In_875);
nor U542 (N_542,In_1054,In_1127);
xor U543 (N_543,N_69,In_1673);
or U544 (N_544,In_319,In_1385);
or U545 (N_545,In_553,In_1947);
or U546 (N_546,In_965,In_1964);
nor U547 (N_547,In_671,In_1960);
xor U548 (N_548,N_206,In_256);
or U549 (N_549,In_1534,In_1948);
nand U550 (N_550,In_923,In_480);
nor U551 (N_551,In_1457,N_273);
xnor U552 (N_552,N_380,N_193);
xnor U553 (N_553,In_1006,N_164);
nand U554 (N_554,In_1055,In_272);
xor U555 (N_555,N_13,In_1487);
nand U556 (N_556,N_339,In_1778);
and U557 (N_557,In_438,In_1161);
nor U558 (N_558,In_603,In_1570);
or U559 (N_559,In_1445,In_1434);
nand U560 (N_560,In_49,In_1946);
xnor U561 (N_561,In_129,N_390);
and U562 (N_562,N_395,In_559);
xor U563 (N_563,N_267,In_524);
or U564 (N_564,In_727,In_1262);
and U565 (N_565,In_819,In_788);
nor U566 (N_566,In_736,In_552);
nand U567 (N_567,N_297,In_270);
or U568 (N_568,In_298,In_1503);
nor U569 (N_569,In_1452,In_1548);
xnor U570 (N_570,N_19,In_76);
or U571 (N_571,N_316,In_42);
nand U572 (N_572,In_1333,In_1806);
nand U573 (N_573,N_28,In_863);
xnor U574 (N_574,In_1559,N_129);
nand U575 (N_575,In_88,In_765);
or U576 (N_576,In_985,In_275);
nor U577 (N_577,In_1728,N_336);
nand U578 (N_578,In_1772,N_5);
or U579 (N_579,In_1854,In_1019);
nand U580 (N_580,In_624,In_1953);
xor U581 (N_581,N_147,In_470);
xor U582 (N_582,In_1889,In_322);
or U583 (N_583,In_1793,In_831);
nand U584 (N_584,In_439,N_341);
or U585 (N_585,N_137,In_1800);
and U586 (N_586,In_1640,In_916);
or U587 (N_587,In_1475,In_1479);
or U588 (N_588,In_1957,In_224);
or U589 (N_589,In_732,N_331);
or U590 (N_590,In_1925,In_1395);
or U591 (N_591,In_894,In_1779);
nor U592 (N_592,In_548,In_662);
nor U593 (N_593,In_430,In_1563);
nor U594 (N_594,In_1075,In_1016);
or U595 (N_595,In_297,In_110);
nor U596 (N_596,In_928,In_69);
and U597 (N_597,In_468,In_406);
xor U598 (N_598,In_1981,N_225);
or U599 (N_599,N_37,In_683);
or U600 (N_600,In_743,In_1923);
and U601 (N_601,N_293,In_1441);
or U602 (N_602,In_366,In_1711);
and U603 (N_603,N_105,N_198);
nand U604 (N_604,N_311,N_125);
or U605 (N_605,In_1995,In_1522);
xor U606 (N_606,In_1983,In_1325);
nand U607 (N_607,N_99,N_45);
xnor U608 (N_608,In_485,In_1733);
and U609 (N_609,In_1347,N_236);
nor U610 (N_610,N_328,In_1862);
nor U611 (N_611,In_1105,In_801);
and U612 (N_612,In_912,N_381);
nor U613 (N_613,In_1685,In_1208);
xor U614 (N_614,In_713,In_910);
or U615 (N_615,In_1609,N_188);
nor U616 (N_616,N_145,In_1188);
and U617 (N_617,In_661,In_250);
nor U618 (N_618,N_210,In_917);
xor U619 (N_619,In_770,In_89);
xnor U620 (N_620,In_1461,N_110);
nor U621 (N_621,N_165,In_1605);
xnor U622 (N_622,In_1372,In_678);
xor U623 (N_623,In_958,In_48);
nand U624 (N_624,N_185,In_1241);
xnor U625 (N_625,In_715,In_235);
nand U626 (N_626,In_763,In_973);
nand U627 (N_627,In_1227,In_1327);
or U628 (N_628,In_373,In_371);
or U629 (N_629,In_416,N_88);
nor U630 (N_630,In_1319,N_132);
nand U631 (N_631,In_1238,In_1798);
nor U632 (N_632,In_1396,N_90);
nand U633 (N_633,In_1389,N_46);
nor U634 (N_634,N_205,In_375);
nor U635 (N_635,N_123,N_42);
xor U636 (N_636,In_1073,In_869);
nor U637 (N_637,In_799,In_1165);
and U638 (N_638,N_194,In_223);
nor U639 (N_639,In_352,In_1564);
nand U640 (N_640,N_299,In_710);
xnor U641 (N_641,In_1972,In_1587);
xor U642 (N_642,N_278,In_432);
nor U643 (N_643,N_208,In_672);
xnor U644 (N_644,In_849,N_352);
xnor U645 (N_645,In_1590,N_238);
nand U646 (N_646,In_1124,In_1064);
nand U647 (N_647,In_422,In_471);
or U648 (N_648,In_511,In_1283);
xor U649 (N_649,In_1513,In_574);
nor U650 (N_650,In_238,In_396);
nor U651 (N_651,In_897,In_785);
or U652 (N_652,In_1748,In_987);
and U653 (N_653,In_1480,N_229);
or U654 (N_654,In_1945,In_808);
xnor U655 (N_655,N_61,In_1624);
nand U656 (N_656,In_94,In_842);
or U657 (N_657,In_1093,In_284);
and U658 (N_658,In_616,In_1604);
or U659 (N_659,In_335,In_183);
xnor U660 (N_660,N_287,N_271);
xor U661 (N_661,In_369,N_302);
and U662 (N_662,N_139,In_1537);
and U663 (N_663,In_99,In_218);
or U664 (N_664,N_166,In_279);
nor U665 (N_665,In_1335,N_371);
or U666 (N_666,In_453,In_122);
and U667 (N_667,In_421,In_1259);
xor U668 (N_668,In_1063,N_298);
or U669 (N_669,N_256,In_345);
nor U670 (N_670,N_74,In_931);
xnor U671 (N_671,In_181,N_182);
nand U672 (N_672,N_364,N_306);
nand U673 (N_673,N_213,In_1958);
nor U674 (N_674,N_368,N_161);
nor U675 (N_675,N_358,In_1024);
and U676 (N_676,In_569,In_1099);
xnor U677 (N_677,N_73,In_315);
or U678 (N_678,In_306,In_1509);
xor U679 (N_679,N_103,N_349);
and U680 (N_680,In_1809,In_214);
and U681 (N_681,In_70,In_1844);
and U682 (N_682,In_817,In_1096);
nand U683 (N_683,In_1250,In_1543);
or U684 (N_684,In_401,In_1116);
xnor U685 (N_685,In_1710,In_404);
xnor U686 (N_686,In_979,In_1108);
nor U687 (N_687,In_75,In_127);
nand U688 (N_688,In_332,In_1021);
nor U689 (N_689,In_502,In_1317);
xor U690 (N_690,In_550,N_214);
nor U691 (N_691,N_268,In_379);
or U692 (N_692,N_333,In_719);
nand U693 (N_693,In_1281,In_1561);
xnor U694 (N_694,In_1345,N_233);
nor U695 (N_695,In_1301,In_768);
nand U696 (N_696,N_122,N_221);
or U697 (N_697,N_398,In_239);
or U698 (N_698,N_226,In_240);
nor U699 (N_699,In_1911,In_1328);
nor U700 (N_700,N_48,In_1266);
nand U701 (N_701,In_1597,N_16);
xor U702 (N_702,In_1047,In_107);
and U703 (N_703,N_244,N_175);
xnor U704 (N_704,In_1774,N_357);
xnor U705 (N_705,In_584,In_1828);
and U706 (N_706,In_1631,In_1206);
nand U707 (N_707,In_1222,In_1813);
xor U708 (N_708,In_1163,N_265);
and U709 (N_709,In_1785,In_1913);
nand U710 (N_710,In_1310,In_493);
and U711 (N_711,In_807,In_1044);
nand U712 (N_712,In_1998,N_104);
and U713 (N_713,In_708,In_1892);
and U714 (N_714,In_510,In_329);
or U715 (N_715,In_834,In_1712);
nor U716 (N_716,In_1648,N_313);
nand U717 (N_717,In_1765,N_375);
and U718 (N_718,In_1906,N_183);
nor U719 (N_719,In_1645,In_525);
xnor U720 (N_720,In_1391,In_299);
or U721 (N_721,In_1477,In_539);
nand U722 (N_722,In_598,In_1144);
xor U723 (N_723,In_757,In_1293);
xor U724 (N_724,N_43,In_132);
xnor U725 (N_725,In_1482,N_131);
nand U726 (N_726,In_1147,N_270);
nor U727 (N_727,In_1658,In_675);
and U728 (N_728,N_116,In_1092);
and U729 (N_729,N_153,In_795);
or U730 (N_730,In_1703,In_139);
nand U731 (N_731,In_1346,In_187);
or U732 (N_732,In_1497,In_388);
nor U733 (N_733,In_145,N_345);
and U734 (N_734,In_809,In_458);
xor U735 (N_735,N_276,In_798);
nor U736 (N_736,In_796,N_144);
nand U737 (N_737,In_1143,In_1884);
nand U738 (N_738,In_173,In_1768);
or U739 (N_739,In_1450,In_467);
nand U740 (N_740,In_487,In_776);
nand U741 (N_741,In_951,In_1679);
nor U742 (N_742,In_1043,In_1304);
nand U743 (N_743,In_625,In_1700);
xnor U744 (N_744,N_84,In_35);
xnor U745 (N_745,In_1423,In_1694);
or U746 (N_746,In_1410,N_327);
or U747 (N_747,In_1436,In_587);
or U748 (N_748,N_186,In_465);
or U749 (N_749,In_1817,In_778);
xor U750 (N_750,N_72,In_1547);
nand U751 (N_751,In_1486,N_29);
nand U752 (N_752,In_1900,In_1417);
xnor U753 (N_753,In_1512,In_451);
nand U754 (N_754,In_1583,In_1035);
and U755 (N_755,N_176,In_1568);
or U756 (N_756,In_1249,N_245);
nor U757 (N_757,In_907,N_162);
or U758 (N_758,N_224,In_1926);
or U759 (N_759,In_1125,In_508);
nor U760 (N_760,N_7,In_1969);
nand U761 (N_761,In_1666,N_212);
xnor U762 (N_762,In_40,N_55);
nor U763 (N_763,In_1719,N_384);
xor U764 (N_764,In_459,In_1426);
xnor U765 (N_765,In_1160,N_138);
and U766 (N_766,In_1000,In_1408);
nand U767 (N_767,N_120,In_566);
or U768 (N_768,In_1510,In_825);
or U769 (N_769,In_203,In_1903);
nor U770 (N_770,In_1337,In_1268);
nand U771 (N_771,In_1752,In_684);
and U772 (N_772,In_2,N_171);
xnor U773 (N_773,N_82,In_793);
or U774 (N_774,In_1140,N_373);
nand U775 (N_775,N_168,In_1113);
nand U776 (N_776,In_1962,In_1651);
nor U777 (N_777,In_1625,In_1986);
nand U778 (N_778,N_359,N_156);
nand U779 (N_779,N_372,In_1404);
xor U780 (N_780,In_946,In_38);
xor U781 (N_781,In_492,In_640);
xor U782 (N_782,In_1876,In_1193);
xnor U783 (N_783,In_1353,In_998);
nor U784 (N_784,In_1818,N_12);
xnor U785 (N_785,In_890,N_353);
nand U786 (N_786,In_301,In_1827);
and U787 (N_787,In_1521,In_1678);
or U788 (N_788,N_272,N_155);
or U789 (N_789,N_258,In_745);
and U790 (N_790,In_1520,In_1789);
or U791 (N_791,In_1810,N_109);
xnor U792 (N_792,In_59,In_1455);
xnor U793 (N_793,In_138,In_22);
and U794 (N_794,In_1873,In_1991);
or U795 (N_795,In_1656,N_118);
xor U796 (N_796,In_134,In_562);
nor U797 (N_797,In_1402,N_78);
nor U798 (N_798,In_868,In_1805);
and U799 (N_799,In_845,In_83);
nand U800 (N_800,In_290,N_584);
nand U801 (N_801,N_557,N_478);
nor U802 (N_802,In_1001,N_770);
and U803 (N_803,In_1538,N_281);
or U804 (N_804,In_323,N_93);
xnor U805 (N_805,N_541,N_619);
xor U806 (N_806,N_594,N_522);
and U807 (N_807,N_179,In_1217);
nor U808 (N_808,In_1908,N_791);
nor U809 (N_809,N_498,In_1660);
or U810 (N_810,N_628,N_337);
nand U811 (N_811,N_566,In_1280);
xnor U812 (N_812,N_409,In_1387);
or U813 (N_813,In_1189,In_841);
and U814 (N_814,N_635,N_638);
or U815 (N_815,In_1111,In_254);
nand U816 (N_816,N_169,In_1406);
nand U817 (N_817,In_1683,In_1162);
xor U818 (N_818,N_616,In_278);
or U819 (N_819,In_1172,N_76);
xor U820 (N_820,In_1230,In_1608);
and U821 (N_821,N_366,In_1504);
and U822 (N_822,N_360,In_357);
nand U823 (N_823,N_27,N_152);
nand U824 (N_824,N_492,N_319);
and U825 (N_825,In_1351,N_701);
xor U826 (N_826,In_804,N_581);
nand U827 (N_827,N_751,In_854);
nand U828 (N_828,In_425,In_720);
and U829 (N_829,In_1915,N_675);
or U830 (N_830,N_307,In_1782);
nor U831 (N_831,In_1194,N_704);
and U832 (N_832,N_443,In_1705);
xor U833 (N_833,In_1585,In_146);
or U834 (N_834,In_362,In_557);
and U835 (N_835,In_1229,N_475);
and U836 (N_836,N_354,N_441);
xor U837 (N_837,N_178,N_394);
nor U838 (N_838,N_304,In_136);
nor U839 (N_839,N_468,In_500);
xor U840 (N_840,N_389,N_545);
and U841 (N_841,In_1296,N_59);
xnor U842 (N_842,In_955,In_729);
and U843 (N_843,N_697,In_98);
nor U844 (N_844,N_219,In_570);
nor U845 (N_845,N_708,N_234);
or U846 (N_846,N_568,In_1519);
xor U847 (N_847,N_779,N_669);
nor U848 (N_848,N_430,N_781);
or U849 (N_849,In_411,N_793);
nor U850 (N_850,N_393,In_251);
nor U851 (N_851,In_360,N_496);
nor U852 (N_852,N_35,In_833);
nor U853 (N_853,In_1050,In_1231);
nor U854 (N_854,In_104,In_68);
nand U855 (N_855,N_472,In_274);
nand U856 (N_856,N_577,N_491);
xnor U857 (N_857,N_694,N_501);
nor U858 (N_858,In_1567,N_44);
or U859 (N_859,N_799,N_348);
nor U860 (N_860,N_787,N_126);
nand U861 (N_861,In_1245,In_1574);
and U862 (N_862,In_634,N_464);
and U863 (N_863,In_1602,N_462);
nor U864 (N_864,N_437,In_311);
nand U865 (N_865,N_683,In_1808);
or U866 (N_866,N_290,N_343);
nand U867 (N_867,N_529,In_27);
nor U868 (N_868,In_1932,N_223);
or U869 (N_869,In_249,N_624);
or U870 (N_870,In_308,In_1725);
xnor U871 (N_871,N_218,In_612);
nand U872 (N_872,In_174,In_561);
xor U873 (N_873,In_455,N_135);
nand U874 (N_874,N_569,N_667);
xor U875 (N_875,In_398,In_1533);
nand U876 (N_876,In_1430,In_81);
xnor U877 (N_877,N_703,In_229);
nand U878 (N_878,In_1912,N_388);
xnor U879 (N_879,N_747,In_1462);
or U880 (N_880,N_143,N_253);
nand U881 (N_881,N_4,N_586);
and U882 (N_882,In_851,N_547);
nand U883 (N_883,In_1723,In_1641);
and U884 (N_884,N_36,N_642);
xor U885 (N_885,N_474,In_1060);
nor U886 (N_886,N_134,In_1517);
and U887 (N_887,In_1356,N_611);
nor U888 (N_888,N_759,N_794);
and U889 (N_889,N_419,In_1551);
or U890 (N_890,N_203,N_3);
or U891 (N_891,In_623,N_636);
nor U892 (N_892,N_62,In_936);
nor U893 (N_893,N_556,In_1077);
xor U894 (N_894,N_25,In_938);
or U895 (N_895,In_1812,In_829);
xnor U896 (N_896,N_606,N_286);
and U897 (N_897,N_698,N_749);
xor U898 (N_898,N_670,In_1684);
nand U899 (N_899,In_191,N_476);
and U900 (N_900,N_274,N_752);
and U901 (N_901,In_1305,N_97);
and U902 (N_902,In_1207,N_315);
and U903 (N_903,N_222,N_502);
xor U904 (N_904,In_1722,In_1856);
and U905 (N_905,In_1042,In_152);
nand U906 (N_906,N_617,N_291);
xnor U907 (N_907,N_653,N_163);
xnor U908 (N_908,N_482,N_459);
xor U909 (N_909,N_486,N_15);
nor U910 (N_910,In_1883,N_89);
and U911 (N_911,In_1738,N_629);
and U912 (N_912,N_657,In_1257);
or U913 (N_913,N_321,N_379);
nand U914 (N_914,In_597,In_1466);
or U915 (N_915,In_772,N_609);
or U916 (N_916,In_1629,In_515);
nand U917 (N_917,N_374,N_682);
xnor U918 (N_918,In_339,N_622);
or U919 (N_919,In_1996,In_828);
nor U920 (N_920,In_292,In_1341);
or U921 (N_921,In_1128,In_1313);
and U922 (N_922,N_621,In_724);
nor U923 (N_923,N_220,In_980);
nand U924 (N_924,In_236,N_717);
nor U925 (N_925,In_1724,N_660);
nand U926 (N_926,In_1764,N_367);
and U927 (N_927,N_158,In_742);
and U928 (N_928,In_549,N_754);
nand U929 (N_929,N_216,N_350);
or U930 (N_930,N_170,N_191);
nor U931 (N_931,N_199,In_336);
or U932 (N_932,N_177,In_1970);
and U933 (N_933,In_1943,In_885);
nor U934 (N_934,N_768,N_778);
xor U935 (N_935,In_1322,N_9);
nand U936 (N_936,In_738,N_648);
and U937 (N_937,In_1338,In_1295);
or U938 (N_938,In_434,N_85);
and U939 (N_939,N_382,In_1659);
nor U940 (N_940,In_1698,In_526);
nor U941 (N_941,N_257,In_1820);
nor U942 (N_942,In_784,N_753);
and U943 (N_943,N_405,In_1138);
or U944 (N_944,In_1400,N_429);
xnor U945 (N_945,In_1823,In_1242);
nor U946 (N_946,N_561,N_172);
xor U947 (N_947,N_260,In_1573);
nor U948 (N_948,In_952,N_266);
or U949 (N_949,N_718,N_607);
and U950 (N_950,N_157,In_180);
xnor U951 (N_951,In_452,N_356);
or U952 (N_952,N_726,N_495);
xor U953 (N_953,N_154,N_605);
nand U954 (N_954,In_838,N_524);
xor U955 (N_955,N_686,N_289);
and U956 (N_956,N_543,In_919);
nor U957 (N_957,N_292,N_542);
or U958 (N_958,N_128,In_1256);
nand U959 (N_959,In_1097,N_696);
xnor U960 (N_960,N_731,N_23);
xnor U961 (N_961,N_576,N_444);
nor U962 (N_962,In_428,N_513);
and U963 (N_963,N_285,In_354);
xnor U964 (N_964,N_544,In_753);
nand U965 (N_965,N_67,In_934);
and U966 (N_966,In_790,In_1592);
xnor U967 (N_967,N_457,N_0);
xnor U968 (N_968,In_7,N_738);
nor U969 (N_969,In_372,In_1978);
or U970 (N_970,N_668,N_420);
nand U971 (N_971,In_376,In_103);
and U972 (N_972,In_1575,N_243);
nor U973 (N_973,In_1270,In_414);
nor U974 (N_974,In_294,In_484);
and U975 (N_975,N_416,In_1115);
nand U976 (N_976,N_512,In_716);
nor U977 (N_977,N_706,In_901);
or U978 (N_978,In_1751,In_1045);
xor U979 (N_979,N_499,In_737);
xor U980 (N_980,N_615,N_386);
nor U981 (N_981,In_1373,N_618);
or U982 (N_982,In_220,In_752);
and U983 (N_983,N_663,In_213);
nand U984 (N_984,N_20,In_1179);
nand U985 (N_985,N_508,In_1297);
and U986 (N_986,N_425,In_1203);
or U987 (N_987,In_1057,N_723);
nor U988 (N_988,In_313,In_1675);
nor U989 (N_989,In_1688,N_451);
or U990 (N_990,N_180,N_22);
and U991 (N_991,N_51,In_1240);
and U992 (N_992,In_635,In_871);
nand U993 (N_993,N_526,N_275);
nand U994 (N_994,In_1905,N_737);
nor U995 (N_995,In_1742,In_443);
nor U996 (N_996,In_859,In_769);
xnor U997 (N_997,N_310,In_1300);
xor U998 (N_998,In_1137,In_893);
nand U999 (N_999,In_1595,In_227);
nor U1000 (N_1000,In_1672,N_528);
xnor U1001 (N_1001,N_52,In_1226);
and U1002 (N_1002,N_797,In_1557);
or U1003 (N_1003,N_401,In_1049);
xnor U1004 (N_1004,In_670,N_573);
or U1005 (N_1005,In_988,In_1821);
and U1006 (N_1006,N_644,N_217);
nand U1007 (N_1007,N_538,In_1526);
xor U1008 (N_1008,In_1427,N_567);
or U1009 (N_1009,N_534,In_1600);
nand U1010 (N_1010,N_509,N_432);
xnor U1011 (N_1011,N_728,N_789);
nand U1012 (N_1012,In_328,N_477);
nand U1013 (N_1013,In_1865,In_1617);
nand U1014 (N_1014,N_344,N_583);
xnor U1015 (N_1015,N_626,N_329);
nor U1016 (N_1016,In_1254,N_695);
and U1017 (N_1017,In_1714,N_469);
nor U1018 (N_1018,In_115,In_23);
xnor U1019 (N_1019,In_1158,In_1383);
nor U1020 (N_1020,N_555,N_705);
and U1021 (N_1021,In_540,N_757);
xnor U1022 (N_1022,N_133,In_1661);
xor U1023 (N_1023,N_484,N_724);
nor U1024 (N_1024,N_408,In_861);
xor U1025 (N_1025,N_200,In_1159);
nand U1026 (N_1026,N_454,In_1909);
xnor U1027 (N_1027,In_1716,N_60);
or U1028 (N_1028,In_1532,N_772);
xnor U1029 (N_1029,N_119,N_294);
or U1030 (N_1030,N_64,N_361);
or U1031 (N_1031,In_1375,In_664);
xor U1032 (N_1032,In_637,N_431);
nand U1033 (N_1033,N_614,In_155);
nand U1034 (N_1034,N_400,N_414);
or U1035 (N_1035,In_1198,In_1456);
nor U1036 (N_1036,In_590,In_1638);
xnor U1037 (N_1037,N_322,In_991);
and U1038 (N_1038,In_417,N_404);
or U1039 (N_1039,In_654,In_532);
or U1040 (N_1040,In_722,In_839);
nand U1041 (N_1041,In_1966,In_712);
and U1042 (N_1042,N_376,In_1431);
or U1043 (N_1043,In_119,N_507);
or U1044 (N_1044,In_1968,In_1089);
nor U1045 (N_1045,In_1622,In_860);
xor U1046 (N_1046,N_604,N_688);
and U1047 (N_1047,N_427,N_413);
xor U1048 (N_1048,N_550,N_687);
and U1049 (N_1049,In_630,In_50);
or U1050 (N_1050,In_1459,In_1872);
nand U1051 (N_1051,In_1988,N_318);
nor U1052 (N_1052,N_504,In_1775);
or U1053 (N_1053,N_563,N_346);
xnor U1054 (N_1054,N_458,N_756);
nand U1055 (N_1055,N_571,In_1831);
or U1056 (N_1056,In_217,N_314);
and U1057 (N_1057,N_664,N_510);
nor U1058 (N_1058,N_473,In_1804);
nand U1059 (N_1059,N_601,N_546);
nor U1060 (N_1060,In_876,In_1204);
nor U1061 (N_1061,N_767,N_575);
nand U1062 (N_1062,In_60,N_665);
nand U1063 (N_1063,In_756,In_565);
nand U1064 (N_1064,N_530,In_1340);
nor U1065 (N_1065,In_504,N_421);
or U1066 (N_1066,N_570,In_1790);
nor U1067 (N_1067,N_572,N_643);
xnor U1068 (N_1068,N_436,N_340);
or U1069 (N_1069,N_411,N_514);
nor U1070 (N_1070,N_646,N_521);
nand U1071 (N_1071,N_392,N_305);
xnor U1072 (N_1072,N_39,In_1454);
or U1073 (N_1073,In_1318,In_1663);
nor U1074 (N_1074,In_520,In_186);
xor U1075 (N_1075,N_719,In_87);
xnor U1076 (N_1076,N_250,N_86);
nor U1077 (N_1077,N_681,N_641);
nor U1078 (N_1078,N_788,In_896);
nand U1079 (N_1079,In_418,N_279);
xor U1080 (N_1080,N_746,In_872);
xor U1081 (N_1081,N_487,In_580);
and U1082 (N_1082,N_721,In_1936);
nand U1083 (N_1083,In_176,In_209);
nand U1084 (N_1084,In_1792,In_1737);
nor U1085 (N_1085,In_972,N_549);
xnor U1086 (N_1086,N_124,N_776);
and U1087 (N_1087,N_255,In_100);
nor U1088 (N_1088,N_795,In_340);
nor U1089 (N_1089,In_1904,N_418);
xor U1090 (N_1090,In_56,In_395);
xor U1091 (N_1091,In_922,In_1216);
and U1092 (N_1092,N_362,In_667);
xnor U1093 (N_1093,N_130,In_78);
and U1094 (N_1094,In_1424,N_516);
and U1095 (N_1095,N_671,N_755);
nor U1096 (N_1096,In_1379,In_387);
nor U1097 (N_1097,In_1027,In_117);
nor U1098 (N_1098,In_305,In_613);
xor U1099 (N_1099,In_764,N_722);
and U1100 (N_1100,In_714,In_1799);
xnor U1101 (N_1101,In_1453,N_523);
nand U1102 (N_1102,In_1107,In_1451);
xnor U1103 (N_1103,In_853,N_300);
and U1104 (N_1104,In_215,In_726);
nor U1105 (N_1105,In_794,N_764);
xor U1106 (N_1106,In_1891,N_634);
xor U1107 (N_1107,In_5,In_882);
nor U1108 (N_1108,N_600,In_1397);
nor U1109 (N_1109,N_32,N_613);
and U1110 (N_1110,N_693,In_899);
and U1111 (N_1111,In_1777,In_1603);
xnor U1112 (N_1112,N_50,In_367);
and U1113 (N_1113,N_403,N_602);
xor U1114 (N_1114,In_344,N_196);
or U1115 (N_1115,In_1382,N_396);
and U1116 (N_1116,In_1871,N_231);
nor U1117 (N_1117,N_515,N_599);
or U1118 (N_1118,In_12,N_654);
and U1119 (N_1119,N_729,N_485);
nand U1120 (N_1120,N_574,In_1071);
nor U1121 (N_1121,In_1036,N_301);
nand U1122 (N_1122,In_264,In_1669);
or U1123 (N_1123,N_209,N_483);
nor U1124 (N_1124,N_412,In_1927);
nand U1125 (N_1125,N_553,N_733);
nand U1126 (N_1126,In_1702,In_1853);
nor U1127 (N_1127,In_1314,N_280);
nor U1128 (N_1128,N_230,N_727);
xnor U1129 (N_1129,N_691,In_1745);
and U1130 (N_1130,N_782,In_1151);
nor U1131 (N_1131,In_1483,N_700);
nand U1132 (N_1132,In_243,N_494);
or U1133 (N_1133,N_262,N_465);
and U1134 (N_1134,N_715,N_232);
or U1135 (N_1135,In_1924,N_453);
nand U1136 (N_1136,N_237,In_1929);
nor U1137 (N_1137,In_43,N_792);
nor U1138 (N_1138,In_1223,N_732);
nor U1139 (N_1139,In_633,N_26);
nor U1140 (N_1140,In_488,In_1514);
and U1141 (N_1141,N_535,N_417);
nand U1142 (N_1142,In_1933,In_1627);
nor U1143 (N_1143,In_976,N_113);
nand U1144 (N_1144,In_219,In_1576);
or U1145 (N_1145,N_678,In_192);
and U1146 (N_1146,N_596,In_741);
or U1147 (N_1147,N_520,In_1009);
nand U1148 (N_1148,N_712,In_929);
or U1149 (N_1149,In_1896,In_1384);
and U1150 (N_1150,In_1643,N_736);
nand U1151 (N_1151,N_422,In_643);
or U1152 (N_1152,N_652,In_944);
and U1153 (N_1153,In_1320,In_800);
nand U1154 (N_1154,In_1795,N_740);
xor U1155 (N_1155,In_1344,N_117);
nor U1156 (N_1156,In_324,In_585);
nor U1157 (N_1157,In_244,N_590);
or U1158 (N_1158,In_1508,N_679);
nor U1159 (N_1159,In_1101,In_555);
xor U1160 (N_1160,In_273,In_445);
nor U1161 (N_1161,In_1442,N_455);
and U1162 (N_1162,N_235,In_474);
xnor U1163 (N_1163,N_623,N_303);
xor U1164 (N_1164,N_564,N_761);
nand U1165 (N_1165,In_1836,N_647);
xor U1166 (N_1166,In_1145,In_1072);
or U1167 (N_1167,In_836,In_803);
or U1168 (N_1168,N_745,In_46);
or U1169 (N_1169,N_725,In_156);
nand U1170 (N_1170,In_1237,In_1003);
or U1171 (N_1171,N_450,In_403);
nand U1172 (N_1172,N_780,In_200);
or U1173 (N_1173,N_610,In_1619);
nand U1174 (N_1174,N_410,In_228);
or U1175 (N_1175,N_146,N_593);
or U1176 (N_1176,In_962,N_689);
or U1177 (N_1177,In_1623,In_182);
or U1178 (N_1178,In_746,In_441);
xor U1179 (N_1179,In_1265,In_448);
nor U1180 (N_1180,N_562,N_75);
and U1181 (N_1181,N_140,N_100);
or U1182 (N_1182,N_239,In_1326);
nand U1183 (N_1183,N_588,In_54);
xnor U1184 (N_1184,In_563,In_31);
nor U1185 (N_1185,In_964,In_1894);
xnor U1186 (N_1186,N_190,N_666);
and U1187 (N_1187,In_67,In_571);
and U1188 (N_1188,In_1670,N_548);
and U1189 (N_1189,In_32,N_383);
and U1190 (N_1190,N_83,In_1546);
and U1191 (N_1191,In_8,N_461);
xor U1192 (N_1192,In_1015,In_1074);
and U1193 (N_1193,In_1191,In_1542);
nor U1194 (N_1194,N_587,In_1469);
nor U1195 (N_1195,In_144,N_603);
nand U1196 (N_1196,In_1729,N_505);
xnor U1197 (N_1197,N_14,N_87);
xor U1198 (N_1198,N_151,N_684);
or U1199 (N_1199,N_312,In_394);
or U1200 (N_1200,N_1170,N_434);
nand U1201 (N_1201,N_969,N_1085);
or U1202 (N_1202,N_597,In_960);
or U1203 (N_1203,N_407,N_1187);
nand U1204 (N_1204,In_29,In_1298);
nor U1205 (N_1205,N_1093,In_1088);
and U1206 (N_1206,N_989,N_828);
nor U1207 (N_1207,N_651,In_1419);
xnor U1208 (N_1208,N_735,N_579);
nand U1209 (N_1209,N_739,N_1135);
nor U1210 (N_1210,N_1043,In_84);
or U1211 (N_1211,N_1029,In_993);
nand U1212 (N_1212,N_1031,N_806);
xnor U1213 (N_1213,N_261,N_826);
nand U1214 (N_1214,N_1016,In_1354);
xor U1215 (N_1215,N_956,N_1126);
or U1216 (N_1216,N_907,N_862);
and U1217 (N_1217,In_1039,N_1019);
and U1218 (N_1218,In_1842,N_713);
or U1219 (N_1219,In_811,N_1109);
nand U1220 (N_1220,N_1021,In_601);
nand U1221 (N_1221,In_1950,N_880);
nor U1222 (N_1222,N_973,N_92);
nand U1223 (N_1223,N_1133,N_1049);
xor U1224 (N_1224,N_608,N_1115);
nor U1225 (N_1225,N_971,In_692);
or U1226 (N_1226,N_330,N_860);
nor U1227 (N_1227,N_1056,N_1167);
nand U1228 (N_1228,N_673,N_783);
and U1229 (N_1229,N_864,N_655);
or U1230 (N_1230,N_1188,In_1857);
nand U1231 (N_1231,N_195,N_829);
or U1232 (N_1232,In_225,N_1015);
or U1233 (N_1233,N_1018,N_1173);
nor U1234 (N_1234,In_704,N_808);
nor U1235 (N_1235,N_918,N_277);
nor U1236 (N_1236,N_992,N_1158);
nand U1237 (N_1237,N_506,N_1091);
nor U1238 (N_1238,N_537,N_997);
and U1239 (N_1239,N_625,N_519);
nand U1240 (N_1240,N_958,In_536);
xor U1241 (N_1241,N_916,N_714);
xnor U1242 (N_1242,N_1168,N_1116);
xnor U1243 (N_1243,N_929,N_982);
nor U1244 (N_1244,N_730,N_269);
xor U1245 (N_1245,N_931,N_674);
or U1246 (N_1246,N_68,N_872);
or U1247 (N_1247,N_1190,N_857);
xnor U1248 (N_1248,N_986,N_1176);
or U1249 (N_1249,N_533,N_640);
xor U1250 (N_1250,N_1137,N_1035);
nand U1251 (N_1251,N_351,N_865);
and U1252 (N_1252,In_889,N_932);
nand U1253 (N_1253,N_943,N_1055);
or U1254 (N_1254,N_922,N_467);
and U1255 (N_1255,N_838,N_1072);
xnor U1256 (N_1256,N_954,N_585);
nor U1257 (N_1257,N_1169,In_1788);
nand U1258 (N_1258,N_1193,N_1079);
nor U1259 (N_1259,N_765,N_831);
nand U1260 (N_1260,N_844,N_202);
nand U1261 (N_1261,N_843,N_627);
xor U1262 (N_1262,N_1191,In_1614);
nor U1263 (N_1263,In_1290,In_688);
nor U1264 (N_1264,N_439,In_567);
nor U1265 (N_1265,N_909,N_1014);
or U1266 (N_1266,N_639,N_460);
xnor U1267 (N_1267,N_879,N_871);
nand U1268 (N_1268,N_899,N_743);
xor U1269 (N_1269,In_1288,N_552);
nand U1270 (N_1270,N_934,N_1070);
and U1271 (N_1271,N_1113,N_869);
and U1272 (N_1272,In_1990,N_874);
or U1273 (N_1273,In_1769,N_1077);
nand U1274 (N_1274,In_18,In_327);
nand U1275 (N_1275,N_1020,In_1581);
nand U1276 (N_1276,N_136,In_1157);
nor U1277 (N_1277,N_1057,N_377);
or U1278 (N_1278,N_942,N_1051);
xor U1279 (N_1279,N_1157,N_819);
or U1280 (N_1280,In_815,N_1089);
xnor U1281 (N_1281,N_592,N_1013);
nand U1282 (N_1282,N_881,N_786);
or U1283 (N_1283,N_1117,N_518);
nor U1284 (N_1284,In_873,In_1299);
nor U1285 (N_1285,N_1151,N_580);
xnor U1286 (N_1286,N_813,N_56);
nand U1287 (N_1287,N_903,N_1112);
nand U1288 (N_1288,N_649,In_1837);
xnor U1289 (N_1289,N_1185,N_1046);
or U1290 (N_1290,N_656,N_187);
nand U1291 (N_1291,In_602,N_822);
and U1292 (N_1292,N_466,N_1102);
or U1293 (N_1293,N_1196,In_1941);
nor U1294 (N_1294,In_659,In_426);
nand U1295 (N_1295,N_995,N_525);
or U1296 (N_1296,N_1165,N_511);
nor U1297 (N_1297,In_1726,In_1321);
or U1298 (N_1298,N_910,N_167);
nor U1299 (N_1299,N_711,N_925);
or U1300 (N_1300,In_655,N_1);
xnor U1301 (N_1301,N_905,N_944);
xor U1302 (N_1302,N_870,In_163);
nor U1303 (N_1303,N_868,N_815);
xnor U1304 (N_1304,In_1885,N_896);
or U1305 (N_1305,N_661,N_633);
or U1306 (N_1306,N_863,N_1149);
nor U1307 (N_1307,N_650,N_1136);
and U1308 (N_1308,N_1146,N_1106);
or U1309 (N_1309,N_1037,In_739);
nand U1310 (N_1310,N_825,N_961);
and U1311 (N_1311,N_426,N_835);
xnor U1312 (N_1312,N_886,In_1066);
xnor U1313 (N_1313,In_1989,N_979);
nand U1314 (N_1314,In_1530,N_758);
and U1315 (N_1315,In_1184,In_1393);
xor U1316 (N_1316,N_1071,N_834);
nand U1317 (N_1317,In_977,N_121);
and U1318 (N_1318,N_1114,N_937);
and U1319 (N_1319,N_326,In_1566);
nand U1320 (N_1320,N_21,N_741);
or U1321 (N_1321,N_1162,N_1009);
nor U1322 (N_1322,N_1123,In_937);
or U1323 (N_1323,N_742,N_1027);
or U1324 (N_1324,In_263,In_494);
and U1325 (N_1325,N_1003,N_560);
nand U1326 (N_1326,N_762,In_1668);
nor U1327 (N_1327,N_1131,N_1061);
xnor U1328 (N_1328,N_1084,N_559);
nor U1329 (N_1329,In_600,N_471);
and U1330 (N_1330,N_1198,N_987);
or U1331 (N_1331,In_1153,N_338);
and U1332 (N_1332,N_488,In_1796);
nand U1333 (N_1333,N_435,N_846);
nor U1334 (N_1334,N_470,N_1033);
nor U1335 (N_1335,N_334,N_895);
or U1336 (N_1336,N_565,N_589);
xnor U1337 (N_1337,In_1596,N_824);
and U1338 (N_1338,N_1058,N_1005);
nand U1339 (N_1339,N_930,N_503);
and U1340 (N_1340,N_1095,N_1087);
or U1341 (N_1341,In_1882,N_821);
and U1342 (N_1342,In_1339,N_252);
nor U1343 (N_1343,N_710,N_591);
nor U1344 (N_1344,N_423,N_892);
nor U1345 (N_1345,N_489,N_1023);
xor U1346 (N_1346,N_1160,N_1148);
xnor U1347 (N_1347,N_65,N_852);
nand U1348 (N_1348,N_1140,N_440);
xnor U1349 (N_1349,N_919,In_627);
xnor U1350 (N_1350,N_1002,In_252);
nand U1351 (N_1351,N_960,N_915);
nor U1352 (N_1352,N_1097,N_803);
or U1353 (N_1353,In_1425,N_962);
xnor U1354 (N_1354,N_452,In_792);
and U1355 (N_1355,N_1034,In_935);
nand U1356 (N_1356,In_1591,N_784);
and U1357 (N_1357,In_1825,In_82);
or U1358 (N_1358,N_598,N_1145);
or U1359 (N_1359,N_785,N_807);
nor U1360 (N_1360,N_8,In_1352);
xor U1361 (N_1361,N_773,N_424);
nor U1362 (N_1362,N_1090,N_532);
nand U1363 (N_1363,N_71,N_842);
nor U1364 (N_1364,N_955,N_1179);
or U1365 (N_1365,In_1082,In_1940);
xor U1366 (N_1366,N_612,In_1068);
nor U1367 (N_1367,N_832,N_449);
nand U1368 (N_1368,N_1122,N_902);
or U1369 (N_1369,N_928,N_631);
nand U1370 (N_1370,N_748,N_947);
and U1371 (N_1371,In_1443,N_830);
or U1372 (N_1372,N_981,N_1088);
xnor U1373 (N_1373,N_867,N_873);
xor U1374 (N_1374,In_334,N_941);
nor U1375 (N_1375,N_1124,N_1110);
and U1376 (N_1376,N_1104,N_975);
xor U1377 (N_1377,N_1098,N_991);
or U1378 (N_1378,N_1125,N_959);
and U1379 (N_1379,N_923,In_170);
or U1380 (N_1380,In_735,N_1010);
or U1381 (N_1381,In_699,N_11);
or U1382 (N_1382,In_1930,N_889);
nand U1383 (N_1383,N_1161,N_1026);
nor U1384 (N_1384,N_1081,In_184);
or U1385 (N_1385,N_848,N_854);
or U1386 (N_1386,In_942,N_645);
xor U1387 (N_1387,N_837,N_1139);
nand U1388 (N_1388,N_978,N_112);
nor U1389 (N_1389,N_1041,N_816);
and U1390 (N_1390,In_105,In_1007);
nor U1391 (N_1391,N_804,N_578);
and U1392 (N_1392,In_66,N_481);
nor U1393 (N_1393,In_1433,N_347);
or U1394 (N_1394,N_1143,In_527);
and U1395 (N_1395,N_888,N_1052);
nand U1396 (N_1396,N_1011,In_74);
or U1397 (N_1397,N_447,N_1028);
nand U1398 (N_1398,In_1606,In_805);
xor U1399 (N_1399,N_1119,N_709);
and U1400 (N_1400,N_428,N_936);
nand U1401 (N_1401,N_893,N_288);
and U1402 (N_1402,N_406,In_1444);
nand U1403 (N_1403,In_556,In_1767);
or U1404 (N_1404,N_812,N_680);
or U1405 (N_1405,In_1484,N_802);
nor U1406 (N_1406,N_847,N_861);
nor U1407 (N_1407,N_994,In_690);
nand U1408 (N_1408,N_983,N_841);
nand U1409 (N_1409,N_1065,N_1174);
or U1410 (N_1410,N_866,N_1166);
nand U1411 (N_1411,In_1025,In_1276);
nor U1412 (N_1412,N_878,N_1008);
nor U1413 (N_1413,N_818,In_1123);
and U1414 (N_1414,In_558,N_446);
or U1415 (N_1415,N_970,N_853);
nand U1416 (N_1416,N_1080,In_1628);
xor U1417 (N_1417,In_533,N_1156);
xnor U1418 (N_1418,N_433,N_904);
nor U1419 (N_1419,In_150,N_1069);
nand U1420 (N_1420,N_385,N_1096);
or U1421 (N_1421,In_126,N_96);
nor U1422 (N_1422,N_692,N_763);
or U1423 (N_1423,N_849,N_998);
or U1424 (N_1424,In_538,N_775);
and U1425 (N_1425,N_913,N_876);
nor U1426 (N_1426,N_536,N_926);
nor U1427 (N_1427,In_47,N_1044);
nor U1428 (N_1428,N_1155,N_1000);
or U1429 (N_1429,N_456,In_1377);
xor U1430 (N_1430,N_891,In_302);
nand U1431 (N_1431,In_420,In_1289);
and U1432 (N_1432,In_908,N_1141);
xor U1433 (N_1433,N_977,N_1004);
nor U1434 (N_1434,N_953,N_796);
nor U1435 (N_1435,N_885,N_810);
or U1436 (N_1436,In_1762,N_949);
xnor U1437 (N_1437,N_1108,N_875);
and U1438 (N_1438,In_210,N_554);
xnor U1439 (N_1439,N_1182,N_699);
xor U1440 (N_1440,N_658,In_1370);
nor U1441 (N_1441,N_1107,N_927);
or U1442 (N_1442,N_790,N_445);
or U1443 (N_1443,N_939,In_1630);
or U1444 (N_1444,In_698,N_284);
nor U1445 (N_1445,In_1639,N_463);
and U1446 (N_1446,In_90,In_501);
xor U1447 (N_1447,In_701,In_1440);
xnor U1448 (N_1448,N_1045,N_1074);
nor U1449 (N_1449,N_911,N_950);
or U1450 (N_1450,N_672,In_1381);
xnor U1451 (N_1451,N_1144,N_850);
xor U1452 (N_1452,N_769,N_493);
nand U1453 (N_1453,N_1062,In_1098);
or U1454 (N_1454,N_801,N_690);
nor U1455 (N_1455,In_1028,N_1175);
nand U1456 (N_1456,N_47,N_1094);
nor U1457 (N_1457,N_1189,N_1121);
xnor U1458 (N_1458,In_206,In_64);
nand U1459 (N_1459,N_1181,N_734);
xor U1460 (N_1460,In_656,N_1138);
nor U1461 (N_1461,In_927,In_791);
and U1462 (N_1462,N_707,N_820);
or U1463 (N_1463,N_894,N_985);
and U1464 (N_1464,N_716,N_1086);
and U1465 (N_1465,N_369,N_98);
nor U1466 (N_1466,N_1197,N_490);
xnor U1467 (N_1467,N_750,N_999);
nor U1468 (N_1468,In_886,N_884);
nand U1469 (N_1469,N_227,In_1255);
or U1470 (N_1470,N_531,N_996);
xor U1471 (N_1471,In_913,N_1163);
nor U1472 (N_1472,N_777,In_489);
and U1473 (N_1473,N_851,In_579);
and U1474 (N_1474,N_34,N_1142);
nor U1475 (N_1475,N_1025,In_852);
xnor U1476 (N_1476,N_1159,N_1127);
and U1477 (N_1477,N_1194,N_952);
xnor U1478 (N_1478,N_877,N_1152);
or U1479 (N_1479,In_111,N_448);
nand U1480 (N_1480,N_964,N_1184);
or U1481 (N_1481,N_1092,In_1739);
xnor U1482 (N_1482,N_702,N_211);
and U1483 (N_1483,In_1979,N_500);
or U1484 (N_1484,N_192,N_974);
nand U1485 (N_1485,N_965,N_1134);
xor U1486 (N_1486,In_199,N_972);
nand U1487 (N_1487,N_898,In_762);
or U1488 (N_1488,In_832,N_415);
nand U1489 (N_1489,In_926,In_1032);
or U1490 (N_1490,In_660,In_382);
or U1491 (N_1491,In_505,In_1215);
nand U1492 (N_1492,In_277,N_632);
and U1493 (N_1493,In_595,N_827);
or U1494 (N_1494,N_1053,In_1181);
nor U1495 (N_1495,N_938,In_1174);
and U1496 (N_1496,N_744,N_1054);
and U1497 (N_1497,N_94,N_1047);
and U1498 (N_1498,N_1059,N_833);
xnor U1499 (N_1499,N_442,N_397);
xor U1500 (N_1500,N_1017,N_1171);
nand U1501 (N_1501,N_1120,N_840);
nor U1502 (N_1502,In_1917,In_1880);
or U1503 (N_1503,N_517,N_1068);
nor U1504 (N_1504,In_179,N_906);
nand U1505 (N_1505,N_1012,N_1164);
nand U1506 (N_1506,N_984,In_383);
nor U1507 (N_1507,N_800,N_836);
nand U1508 (N_1508,In_609,N_662);
nand U1509 (N_1509,In_509,N_1192);
xor U1510 (N_1510,In_397,N_551);
nor U1511 (N_1511,In_1269,N_1082);
and U1512 (N_1512,In_1864,N_912);
and U1513 (N_1513,N_845,N_766);
xor U1514 (N_1514,N_855,N_1183);
nand U1515 (N_1515,N_814,In_1121);
and U1516 (N_1516,N_1038,N_1180);
and U1517 (N_1517,In_1413,N_1001);
and U1518 (N_1518,N_1132,N_882);
and U1519 (N_1519,N_1100,N_1101);
or U1520 (N_1520,N_990,N_951);
or U1521 (N_1521,In_202,N_539);
xnor U1522 (N_1522,In_575,N_1039);
and U1523 (N_1523,In_1863,In_1126);
xnor U1524 (N_1524,In_1919,N_1153);
or U1525 (N_1525,In_1065,N_264);
and U1526 (N_1526,N_1022,N_620);
xor U1527 (N_1527,N_908,N_1060);
and U1528 (N_1528,N_901,N_159);
xor U1529 (N_1529,N_980,N_1105);
and U1530 (N_1530,In_1110,N_1006);
xnor U1531 (N_1531,N_1172,N_963);
nand U1532 (N_1532,N_184,N_558);
and U1533 (N_1533,In_1004,N_774);
or U1534 (N_1534,N_1036,N_1177);
nand U1535 (N_1535,N_1032,N_1064);
xnor U1536 (N_1536,In_96,N_527);
nand U1537 (N_1537,N_809,In_632);
nand U1538 (N_1538,N_859,N_1030);
and U1539 (N_1539,In_447,N_582);
nor U1540 (N_1540,N_479,In_1691);
nand U1541 (N_1541,N_1007,N_957);
nand U1542 (N_1542,N_1067,In_997);
and U1543 (N_1543,N_946,In_1264);
nand U1544 (N_1544,N_1099,N_677);
and U1545 (N_1545,N_676,In_1332);
and U1546 (N_1546,N_1147,N_595);
xor U1547 (N_1547,N_1073,N_890);
and U1548 (N_1548,N_839,In_1202);
nand U1549 (N_1549,N_856,N_1075);
xor U1550 (N_1550,N_967,In_1495);
nor U1551 (N_1551,N_114,N_1195);
nand U1552 (N_1552,N_630,N_1048);
nand U1553 (N_1553,N_246,N_968);
xnor U1554 (N_1554,N_858,N_1024);
nor U1555 (N_1555,N_935,N_1042);
or U1556 (N_1556,N_33,In_450);
nor U1557 (N_1557,In_638,N_798);
xor U1558 (N_1558,N_363,N_241);
xor U1559 (N_1559,N_1103,In_1761);
nand U1560 (N_1560,In_925,In_1874);
nor U1561 (N_1561,In_648,N_823);
nand U1562 (N_1562,N_1130,N_659);
nor U1563 (N_1563,N_637,N_41);
xor U1564 (N_1564,In_608,In_1802);
xnor U1565 (N_1565,N_1083,N_1186);
xor U1566 (N_1566,In_577,N_1129);
nand U1567 (N_1567,In_498,N_897);
or U1568 (N_1568,N_945,N_248);
nand U1569 (N_1569,In_1287,N_940);
nor U1570 (N_1570,N_760,N_720);
and U1571 (N_1571,In_544,N_497);
nor U1572 (N_1572,N_685,N_993);
or U1573 (N_1573,In_1959,N_254);
nand U1574 (N_1574,N_921,N_966);
xnor U1575 (N_1575,N_1040,N_1050);
nor U1576 (N_1576,In_1201,N_1111);
nor U1577 (N_1577,N_540,N_1150);
or U1578 (N_1578,In_1682,N_883);
and U1579 (N_1579,In_607,N_1128);
xor U1580 (N_1580,N_933,N_438);
and U1581 (N_1581,N_771,N_355);
or U1582 (N_1582,In_1492,In_1954);
nand U1583 (N_1583,N_402,N_920);
nor U1584 (N_1584,N_480,N_805);
or U1585 (N_1585,N_914,N_1078);
xnor U1586 (N_1586,In_1797,N_38);
or U1587 (N_1587,N_1063,N_1076);
nand U1588 (N_1588,N_917,N_976);
or U1589 (N_1589,N_887,In_1083);
or U1590 (N_1590,N_1118,N_1178);
xor U1591 (N_1591,N_817,In_457);
nor U1592 (N_1592,In_1192,N_811);
nor U1593 (N_1593,N_79,N_924);
and U1594 (N_1594,N_948,N_900);
nor U1595 (N_1595,In_1498,In_1859);
nor U1596 (N_1596,In_1555,In_102);
nand U1597 (N_1597,In_1164,In_1667);
nor U1598 (N_1598,N_988,N_1199);
and U1599 (N_1599,N_1066,N_1154);
nor U1600 (N_1600,N_1310,N_1219);
nor U1601 (N_1601,N_1469,N_1457);
and U1602 (N_1602,N_1546,N_1277);
xor U1603 (N_1603,N_1307,N_1321);
or U1604 (N_1604,N_1240,N_1204);
or U1605 (N_1605,N_1203,N_1570);
nor U1606 (N_1606,N_1281,N_1487);
and U1607 (N_1607,N_1211,N_1507);
xnor U1608 (N_1608,N_1360,N_1560);
nand U1609 (N_1609,N_1593,N_1244);
or U1610 (N_1610,N_1447,N_1477);
xnor U1611 (N_1611,N_1229,N_1391);
and U1612 (N_1612,N_1298,N_1557);
or U1613 (N_1613,N_1418,N_1235);
xnor U1614 (N_1614,N_1493,N_1414);
nor U1615 (N_1615,N_1522,N_1597);
xor U1616 (N_1616,N_1529,N_1440);
or U1617 (N_1617,N_1396,N_1237);
nand U1618 (N_1618,N_1508,N_1351);
nand U1619 (N_1619,N_1227,N_1231);
nor U1620 (N_1620,N_1410,N_1595);
and U1621 (N_1621,N_1500,N_1382);
nand U1622 (N_1622,N_1584,N_1363);
nand U1623 (N_1623,N_1448,N_1384);
xnor U1624 (N_1624,N_1379,N_1536);
and U1625 (N_1625,N_1545,N_1539);
nand U1626 (N_1626,N_1403,N_1358);
nor U1627 (N_1627,N_1577,N_1389);
or U1628 (N_1628,N_1398,N_1484);
or U1629 (N_1629,N_1427,N_1323);
or U1630 (N_1630,N_1230,N_1374);
nand U1631 (N_1631,N_1460,N_1376);
xnor U1632 (N_1632,N_1263,N_1491);
and U1633 (N_1633,N_1406,N_1425);
xor U1634 (N_1634,N_1302,N_1413);
or U1635 (N_1635,N_1481,N_1354);
xor U1636 (N_1636,N_1269,N_1415);
nand U1637 (N_1637,N_1588,N_1261);
nand U1638 (N_1638,N_1565,N_1473);
xnor U1639 (N_1639,N_1348,N_1258);
or U1640 (N_1640,N_1551,N_1340);
nor U1641 (N_1641,N_1483,N_1350);
and U1642 (N_1642,N_1377,N_1392);
nor U1643 (N_1643,N_1397,N_1355);
and U1644 (N_1644,N_1504,N_1375);
xor U1645 (N_1645,N_1475,N_1494);
nand U1646 (N_1646,N_1547,N_1490);
nor U1647 (N_1647,N_1503,N_1409);
nand U1648 (N_1648,N_1569,N_1554);
or U1649 (N_1649,N_1598,N_1209);
nor U1650 (N_1650,N_1515,N_1318);
or U1651 (N_1651,N_1564,N_1256);
and U1652 (N_1652,N_1214,N_1459);
or U1653 (N_1653,N_1501,N_1502);
and U1654 (N_1654,N_1516,N_1378);
or U1655 (N_1655,N_1566,N_1580);
nand U1656 (N_1656,N_1294,N_1239);
nand U1657 (N_1657,N_1257,N_1401);
xnor U1658 (N_1658,N_1583,N_1300);
nand U1659 (N_1659,N_1543,N_1246);
nor U1660 (N_1660,N_1293,N_1559);
nand U1661 (N_1661,N_1317,N_1439);
and U1662 (N_1662,N_1524,N_1304);
xnor U1663 (N_1663,N_1297,N_1313);
nand U1664 (N_1664,N_1287,N_1444);
nand U1665 (N_1665,N_1552,N_1549);
and U1666 (N_1666,N_1278,N_1544);
and U1667 (N_1667,N_1341,N_1364);
xnor U1668 (N_1668,N_1537,N_1567);
nand U1669 (N_1669,N_1387,N_1541);
nand U1670 (N_1670,N_1486,N_1513);
and U1671 (N_1671,N_1213,N_1412);
xor U1672 (N_1672,N_1563,N_1370);
nor U1673 (N_1673,N_1590,N_1324);
or U1674 (N_1674,N_1367,N_1417);
xor U1675 (N_1675,N_1451,N_1489);
nand U1676 (N_1676,N_1372,N_1200);
xor U1677 (N_1677,N_1579,N_1238);
nand U1678 (N_1678,N_1453,N_1306);
nor U1679 (N_1679,N_1356,N_1326);
xnor U1680 (N_1680,N_1201,N_1420);
nor U1681 (N_1681,N_1575,N_1366);
or U1682 (N_1682,N_1337,N_1290);
and U1683 (N_1683,N_1283,N_1435);
xnor U1684 (N_1684,N_1308,N_1437);
or U1685 (N_1685,N_1292,N_1373);
xnor U1686 (N_1686,N_1436,N_1492);
nand U1687 (N_1687,N_1215,N_1592);
nand U1688 (N_1688,N_1568,N_1434);
or U1689 (N_1689,N_1393,N_1446);
nor U1690 (N_1690,N_1480,N_1485);
xor U1691 (N_1691,N_1510,N_1234);
and U1692 (N_1692,N_1338,N_1352);
nand U1693 (N_1693,N_1582,N_1241);
or U1694 (N_1694,N_1520,N_1249);
xor U1695 (N_1695,N_1576,N_1380);
xnor U1696 (N_1696,N_1556,N_1207);
nand U1697 (N_1697,N_1443,N_1255);
xor U1698 (N_1698,N_1368,N_1478);
nor U1699 (N_1699,N_1349,N_1599);
nand U1700 (N_1700,N_1433,N_1525);
or U1701 (N_1701,N_1216,N_1466);
nor U1702 (N_1702,N_1596,N_1540);
and U1703 (N_1703,N_1571,N_1250);
or U1704 (N_1704,N_1267,N_1225);
and U1705 (N_1705,N_1528,N_1388);
or U1706 (N_1706,N_1498,N_1402);
or U1707 (N_1707,N_1431,N_1330);
nor U1708 (N_1708,N_1472,N_1311);
nor U1709 (N_1709,N_1463,N_1386);
and U1710 (N_1710,N_1328,N_1586);
nor U1711 (N_1711,N_1521,N_1438);
nand U1712 (N_1712,N_1254,N_1224);
nand U1713 (N_1713,N_1523,N_1479);
xor U1714 (N_1714,N_1221,N_1266);
nor U1715 (N_1715,N_1301,N_1344);
and U1716 (N_1716,N_1284,N_1482);
or U1717 (N_1717,N_1573,N_1468);
nand U1718 (N_1718,N_1538,N_1345);
and U1719 (N_1719,N_1456,N_1353);
nor U1720 (N_1720,N_1303,N_1419);
xor U1721 (N_1721,N_1519,N_1562);
nor U1722 (N_1722,N_1532,N_1594);
xor U1723 (N_1723,N_1408,N_1411);
or U1724 (N_1724,N_1553,N_1289);
nand U1725 (N_1725,N_1530,N_1223);
nor U1726 (N_1726,N_1424,N_1445);
or U1727 (N_1727,N_1470,N_1404);
xor U1728 (N_1728,N_1399,N_1262);
or U1729 (N_1729,N_1242,N_1359);
nand U1730 (N_1730,N_1454,N_1587);
xor U1731 (N_1731,N_1581,N_1295);
nor U1732 (N_1732,N_1394,N_1488);
nand U1733 (N_1733,N_1305,N_1282);
or U1734 (N_1734,N_1534,N_1429);
nand U1735 (N_1735,N_1461,N_1268);
nor U1736 (N_1736,N_1316,N_1251);
and U1737 (N_1737,N_1499,N_1205);
xor U1738 (N_1738,N_1511,N_1476);
or U1739 (N_1739,N_1400,N_1442);
xnor U1740 (N_1740,N_1589,N_1361);
or U1741 (N_1741,N_1464,N_1212);
nor U1742 (N_1742,N_1315,N_1346);
xor U1743 (N_1743,N_1558,N_1274);
or U1744 (N_1744,N_1407,N_1259);
and U1745 (N_1745,N_1342,N_1248);
or U1746 (N_1746,N_1329,N_1327);
xor U1747 (N_1747,N_1471,N_1578);
nor U1748 (N_1748,N_1390,N_1371);
nor U1749 (N_1749,N_1265,N_1347);
and U1750 (N_1750,N_1343,N_1217);
or U1751 (N_1751,N_1285,N_1512);
xnor U1752 (N_1752,N_1270,N_1286);
nand U1753 (N_1753,N_1572,N_1228);
nand U1754 (N_1754,N_1405,N_1369);
nor U1755 (N_1755,N_1245,N_1465);
or U1756 (N_1756,N_1220,N_1243);
and U1757 (N_1757,N_1260,N_1236);
and U1758 (N_1758,N_1331,N_1381);
or U1759 (N_1759,N_1385,N_1550);
or U1760 (N_1760,N_1322,N_1574);
nor U1761 (N_1761,N_1309,N_1526);
or U1762 (N_1762,N_1333,N_1273);
nor U1763 (N_1763,N_1296,N_1423);
and U1764 (N_1764,N_1222,N_1426);
or U1765 (N_1765,N_1202,N_1276);
and U1766 (N_1766,N_1312,N_1291);
xnor U1767 (N_1767,N_1383,N_1319);
nand U1768 (N_1768,N_1208,N_1505);
or U1769 (N_1769,N_1253,N_1288);
nand U1770 (N_1770,N_1339,N_1275);
nor U1771 (N_1771,N_1206,N_1467);
and U1772 (N_1772,N_1336,N_1226);
nand U1773 (N_1773,N_1455,N_1527);
and U1774 (N_1774,N_1535,N_1365);
xor U1775 (N_1775,N_1441,N_1450);
xor U1776 (N_1776,N_1462,N_1210);
xnor U1777 (N_1777,N_1531,N_1514);
xor U1778 (N_1778,N_1458,N_1334);
nor U1779 (N_1779,N_1591,N_1416);
or U1780 (N_1780,N_1449,N_1517);
or U1781 (N_1781,N_1422,N_1264);
nor U1782 (N_1782,N_1335,N_1279);
xor U1783 (N_1783,N_1542,N_1561);
nand U1784 (N_1784,N_1280,N_1320);
nand U1785 (N_1785,N_1474,N_1555);
and U1786 (N_1786,N_1332,N_1247);
nor U1787 (N_1787,N_1495,N_1421);
or U1788 (N_1788,N_1357,N_1509);
and U1789 (N_1789,N_1271,N_1314);
nand U1790 (N_1790,N_1218,N_1362);
and U1791 (N_1791,N_1533,N_1452);
xor U1792 (N_1792,N_1585,N_1432);
xor U1793 (N_1793,N_1496,N_1233);
nor U1794 (N_1794,N_1252,N_1325);
nand U1795 (N_1795,N_1272,N_1518);
xnor U1796 (N_1796,N_1497,N_1299);
and U1797 (N_1797,N_1548,N_1428);
nor U1798 (N_1798,N_1430,N_1232);
and U1799 (N_1799,N_1395,N_1506);
xnor U1800 (N_1800,N_1353,N_1338);
or U1801 (N_1801,N_1458,N_1398);
nor U1802 (N_1802,N_1411,N_1539);
or U1803 (N_1803,N_1320,N_1429);
nor U1804 (N_1804,N_1595,N_1533);
or U1805 (N_1805,N_1207,N_1583);
or U1806 (N_1806,N_1401,N_1318);
xor U1807 (N_1807,N_1529,N_1442);
xnor U1808 (N_1808,N_1326,N_1361);
xnor U1809 (N_1809,N_1544,N_1436);
xor U1810 (N_1810,N_1577,N_1480);
or U1811 (N_1811,N_1368,N_1446);
xor U1812 (N_1812,N_1501,N_1599);
nor U1813 (N_1813,N_1381,N_1442);
nor U1814 (N_1814,N_1476,N_1236);
or U1815 (N_1815,N_1597,N_1271);
nor U1816 (N_1816,N_1594,N_1573);
or U1817 (N_1817,N_1524,N_1402);
and U1818 (N_1818,N_1589,N_1579);
xnor U1819 (N_1819,N_1394,N_1336);
xor U1820 (N_1820,N_1364,N_1327);
nand U1821 (N_1821,N_1472,N_1346);
xnor U1822 (N_1822,N_1340,N_1520);
nand U1823 (N_1823,N_1478,N_1443);
nor U1824 (N_1824,N_1404,N_1326);
or U1825 (N_1825,N_1244,N_1317);
nor U1826 (N_1826,N_1491,N_1480);
xnor U1827 (N_1827,N_1384,N_1373);
and U1828 (N_1828,N_1289,N_1415);
nor U1829 (N_1829,N_1394,N_1541);
or U1830 (N_1830,N_1355,N_1504);
nand U1831 (N_1831,N_1431,N_1237);
and U1832 (N_1832,N_1409,N_1428);
and U1833 (N_1833,N_1595,N_1205);
xnor U1834 (N_1834,N_1278,N_1465);
or U1835 (N_1835,N_1469,N_1542);
xor U1836 (N_1836,N_1491,N_1546);
and U1837 (N_1837,N_1577,N_1278);
nor U1838 (N_1838,N_1539,N_1495);
nor U1839 (N_1839,N_1304,N_1461);
and U1840 (N_1840,N_1529,N_1315);
xnor U1841 (N_1841,N_1395,N_1419);
nor U1842 (N_1842,N_1461,N_1270);
or U1843 (N_1843,N_1532,N_1307);
and U1844 (N_1844,N_1304,N_1418);
and U1845 (N_1845,N_1220,N_1240);
or U1846 (N_1846,N_1503,N_1410);
and U1847 (N_1847,N_1455,N_1340);
nor U1848 (N_1848,N_1419,N_1537);
or U1849 (N_1849,N_1441,N_1569);
or U1850 (N_1850,N_1506,N_1575);
and U1851 (N_1851,N_1443,N_1231);
and U1852 (N_1852,N_1401,N_1408);
xor U1853 (N_1853,N_1547,N_1555);
or U1854 (N_1854,N_1485,N_1387);
or U1855 (N_1855,N_1367,N_1307);
nor U1856 (N_1856,N_1480,N_1361);
nand U1857 (N_1857,N_1598,N_1253);
xor U1858 (N_1858,N_1452,N_1246);
nor U1859 (N_1859,N_1278,N_1380);
nor U1860 (N_1860,N_1398,N_1575);
xor U1861 (N_1861,N_1505,N_1342);
xnor U1862 (N_1862,N_1488,N_1390);
nand U1863 (N_1863,N_1255,N_1599);
nor U1864 (N_1864,N_1403,N_1540);
and U1865 (N_1865,N_1414,N_1436);
xor U1866 (N_1866,N_1454,N_1461);
nor U1867 (N_1867,N_1327,N_1511);
xor U1868 (N_1868,N_1257,N_1535);
xor U1869 (N_1869,N_1366,N_1419);
nand U1870 (N_1870,N_1317,N_1574);
xor U1871 (N_1871,N_1384,N_1208);
nor U1872 (N_1872,N_1303,N_1436);
nor U1873 (N_1873,N_1210,N_1240);
nand U1874 (N_1874,N_1395,N_1307);
nor U1875 (N_1875,N_1558,N_1520);
nor U1876 (N_1876,N_1204,N_1553);
and U1877 (N_1877,N_1562,N_1551);
and U1878 (N_1878,N_1475,N_1323);
nand U1879 (N_1879,N_1340,N_1219);
xor U1880 (N_1880,N_1413,N_1529);
and U1881 (N_1881,N_1205,N_1293);
and U1882 (N_1882,N_1497,N_1538);
xor U1883 (N_1883,N_1502,N_1574);
nor U1884 (N_1884,N_1408,N_1368);
and U1885 (N_1885,N_1232,N_1380);
xnor U1886 (N_1886,N_1216,N_1274);
nor U1887 (N_1887,N_1495,N_1212);
nor U1888 (N_1888,N_1477,N_1515);
nor U1889 (N_1889,N_1214,N_1507);
or U1890 (N_1890,N_1539,N_1281);
nor U1891 (N_1891,N_1265,N_1393);
nor U1892 (N_1892,N_1460,N_1369);
xnor U1893 (N_1893,N_1482,N_1207);
and U1894 (N_1894,N_1303,N_1457);
xnor U1895 (N_1895,N_1376,N_1406);
and U1896 (N_1896,N_1333,N_1475);
or U1897 (N_1897,N_1345,N_1432);
nand U1898 (N_1898,N_1403,N_1522);
and U1899 (N_1899,N_1335,N_1526);
nor U1900 (N_1900,N_1317,N_1258);
nand U1901 (N_1901,N_1478,N_1260);
nand U1902 (N_1902,N_1599,N_1319);
xnor U1903 (N_1903,N_1304,N_1403);
nor U1904 (N_1904,N_1253,N_1512);
or U1905 (N_1905,N_1366,N_1237);
or U1906 (N_1906,N_1380,N_1570);
and U1907 (N_1907,N_1542,N_1336);
xnor U1908 (N_1908,N_1594,N_1494);
and U1909 (N_1909,N_1474,N_1224);
nand U1910 (N_1910,N_1572,N_1368);
nand U1911 (N_1911,N_1589,N_1342);
nand U1912 (N_1912,N_1552,N_1413);
xnor U1913 (N_1913,N_1592,N_1261);
or U1914 (N_1914,N_1476,N_1403);
and U1915 (N_1915,N_1353,N_1567);
xor U1916 (N_1916,N_1587,N_1402);
and U1917 (N_1917,N_1513,N_1317);
and U1918 (N_1918,N_1582,N_1230);
and U1919 (N_1919,N_1408,N_1311);
and U1920 (N_1920,N_1226,N_1529);
and U1921 (N_1921,N_1488,N_1377);
nand U1922 (N_1922,N_1354,N_1593);
or U1923 (N_1923,N_1523,N_1573);
or U1924 (N_1924,N_1447,N_1341);
nor U1925 (N_1925,N_1459,N_1418);
or U1926 (N_1926,N_1208,N_1225);
and U1927 (N_1927,N_1373,N_1216);
xnor U1928 (N_1928,N_1419,N_1432);
or U1929 (N_1929,N_1392,N_1228);
nand U1930 (N_1930,N_1329,N_1477);
or U1931 (N_1931,N_1213,N_1546);
nand U1932 (N_1932,N_1596,N_1356);
and U1933 (N_1933,N_1434,N_1425);
nor U1934 (N_1934,N_1408,N_1573);
nor U1935 (N_1935,N_1228,N_1458);
nand U1936 (N_1936,N_1360,N_1423);
nand U1937 (N_1937,N_1255,N_1408);
nand U1938 (N_1938,N_1436,N_1320);
nor U1939 (N_1939,N_1308,N_1532);
nand U1940 (N_1940,N_1561,N_1214);
nand U1941 (N_1941,N_1353,N_1439);
nor U1942 (N_1942,N_1477,N_1251);
and U1943 (N_1943,N_1299,N_1250);
nand U1944 (N_1944,N_1417,N_1203);
or U1945 (N_1945,N_1502,N_1458);
and U1946 (N_1946,N_1419,N_1494);
nand U1947 (N_1947,N_1583,N_1266);
and U1948 (N_1948,N_1356,N_1344);
xnor U1949 (N_1949,N_1315,N_1251);
nor U1950 (N_1950,N_1449,N_1446);
nand U1951 (N_1951,N_1565,N_1331);
nor U1952 (N_1952,N_1452,N_1229);
nand U1953 (N_1953,N_1446,N_1443);
xor U1954 (N_1954,N_1240,N_1308);
and U1955 (N_1955,N_1574,N_1232);
xor U1956 (N_1956,N_1544,N_1534);
or U1957 (N_1957,N_1481,N_1431);
and U1958 (N_1958,N_1450,N_1365);
nor U1959 (N_1959,N_1400,N_1300);
or U1960 (N_1960,N_1396,N_1469);
xor U1961 (N_1961,N_1200,N_1475);
xnor U1962 (N_1962,N_1503,N_1265);
nand U1963 (N_1963,N_1450,N_1206);
xor U1964 (N_1964,N_1301,N_1489);
nand U1965 (N_1965,N_1539,N_1442);
and U1966 (N_1966,N_1240,N_1371);
nor U1967 (N_1967,N_1507,N_1478);
nand U1968 (N_1968,N_1363,N_1536);
nor U1969 (N_1969,N_1348,N_1591);
xnor U1970 (N_1970,N_1471,N_1597);
nand U1971 (N_1971,N_1505,N_1504);
nand U1972 (N_1972,N_1587,N_1563);
nand U1973 (N_1973,N_1321,N_1516);
xor U1974 (N_1974,N_1567,N_1559);
or U1975 (N_1975,N_1521,N_1253);
or U1976 (N_1976,N_1468,N_1246);
nor U1977 (N_1977,N_1522,N_1586);
xnor U1978 (N_1978,N_1389,N_1512);
and U1979 (N_1979,N_1572,N_1423);
and U1980 (N_1980,N_1517,N_1356);
or U1981 (N_1981,N_1591,N_1532);
nand U1982 (N_1982,N_1264,N_1451);
xor U1983 (N_1983,N_1544,N_1530);
xor U1984 (N_1984,N_1502,N_1543);
xor U1985 (N_1985,N_1240,N_1422);
or U1986 (N_1986,N_1213,N_1507);
xor U1987 (N_1987,N_1510,N_1480);
or U1988 (N_1988,N_1293,N_1452);
xnor U1989 (N_1989,N_1387,N_1357);
nor U1990 (N_1990,N_1364,N_1569);
xnor U1991 (N_1991,N_1442,N_1369);
xor U1992 (N_1992,N_1506,N_1550);
and U1993 (N_1993,N_1320,N_1332);
nand U1994 (N_1994,N_1584,N_1440);
or U1995 (N_1995,N_1450,N_1561);
nor U1996 (N_1996,N_1491,N_1449);
nand U1997 (N_1997,N_1265,N_1326);
nand U1998 (N_1998,N_1265,N_1422);
nand U1999 (N_1999,N_1398,N_1334);
nor U2000 (N_2000,N_1918,N_1809);
and U2001 (N_2001,N_1841,N_1931);
nor U2002 (N_2002,N_1829,N_1772);
or U2003 (N_2003,N_1985,N_1638);
nand U2004 (N_2004,N_1935,N_1778);
or U2005 (N_2005,N_1796,N_1894);
xnor U2006 (N_2006,N_1752,N_1703);
or U2007 (N_2007,N_1819,N_1727);
or U2008 (N_2008,N_1782,N_1605);
and U2009 (N_2009,N_1804,N_1818);
xor U2010 (N_2010,N_1890,N_1730);
xnor U2011 (N_2011,N_1876,N_1639);
or U2012 (N_2012,N_1905,N_1929);
nand U2013 (N_2013,N_1789,N_1739);
nand U2014 (N_2014,N_1755,N_1734);
xor U2015 (N_2015,N_1705,N_1943);
nor U2016 (N_2016,N_1653,N_1736);
xnor U2017 (N_2017,N_1847,N_1883);
nand U2018 (N_2018,N_1775,N_1821);
or U2019 (N_2019,N_1997,N_1707);
xnor U2020 (N_2020,N_1628,N_1825);
or U2021 (N_2021,N_1853,N_1741);
xnor U2022 (N_2022,N_1652,N_1783);
xor U2023 (N_2023,N_1948,N_1802);
nand U2024 (N_2024,N_1683,N_1682);
xnor U2025 (N_2025,N_1871,N_1774);
or U2026 (N_2026,N_1610,N_1831);
and U2027 (N_2027,N_1770,N_1824);
nand U2028 (N_2028,N_1887,N_1793);
nor U2029 (N_2029,N_1642,N_1658);
nand U2030 (N_2030,N_1897,N_1679);
and U2031 (N_2031,N_1945,N_1711);
nor U2032 (N_2032,N_1938,N_1870);
or U2033 (N_2033,N_1696,N_1768);
nor U2034 (N_2034,N_1636,N_1827);
and U2035 (N_2035,N_1877,N_1830);
nor U2036 (N_2036,N_1650,N_1840);
nor U2037 (N_2037,N_1872,N_1822);
or U2038 (N_2038,N_1800,N_1867);
nand U2039 (N_2039,N_1915,N_1828);
or U2040 (N_2040,N_1973,N_1903);
and U2041 (N_2041,N_1603,N_1635);
xor U2042 (N_2042,N_1993,N_1919);
xor U2043 (N_2043,N_1732,N_1979);
or U2044 (N_2044,N_1851,N_1917);
or U2045 (N_2045,N_1771,N_1728);
and U2046 (N_2046,N_1712,N_1923);
or U2047 (N_2047,N_1644,N_1620);
or U2048 (N_2048,N_1602,N_1624);
xor U2049 (N_2049,N_1699,N_1992);
nand U2050 (N_2050,N_1893,N_1916);
or U2051 (N_2051,N_1842,N_1777);
xor U2052 (N_2052,N_1814,N_1799);
nand U2053 (N_2053,N_1868,N_1687);
xnor U2054 (N_2054,N_1902,N_1663);
nand U2055 (N_2055,N_1776,N_1749);
and U2056 (N_2056,N_1634,N_1823);
and U2057 (N_2057,N_1694,N_1601);
xor U2058 (N_2058,N_1714,N_1666);
and U2059 (N_2059,N_1688,N_1615);
xnor U2060 (N_2060,N_1745,N_1672);
xor U2061 (N_2061,N_1880,N_1660);
or U2062 (N_2062,N_1906,N_1989);
nor U2063 (N_2063,N_1954,N_1686);
nand U2064 (N_2064,N_1692,N_1884);
or U2065 (N_2065,N_1701,N_1691);
xnor U2066 (N_2066,N_1717,N_1813);
nor U2067 (N_2067,N_1996,N_1801);
xor U2068 (N_2068,N_1860,N_1901);
nand U2069 (N_2069,N_1669,N_1965);
and U2070 (N_2070,N_1951,N_1889);
xnor U2071 (N_2071,N_1640,N_1910);
xor U2072 (N_2072,N_1643,N_1994);
xor U2073 (N_2073,N_1864,N_1859);
nand U2074 (N_2074,N_1875,N_1963);
nor U2075 (N_2075,N_1855,N_1735);
xnor U2076 (N_2076,N_1632,N_1627);
or U2077 (N_2077,N_1836,N_1758);
xor U2078 (N_2078,N_1806,N_1773);
or U2079 (N_2079,N_1788,N_1983);
nor U2080 (N_2080,N_1879,N_1631);
nor U2081 (N_2081,N_1898,N_1764);
or U2082 (N_2082,N_1892,N_1926);
xor U2083 (N_2083,N_1927,N_1737);
xor U2084 (N_2084,N_1680,N_1724);
xnor U2085 (N_2085,N_1656,N_1961);
and U2086 (N_2086,N_1837,N_1808);
nor U2087 (N_2087,N_1698,N_1689);
and U2088 (N_2088,N_1953,N_1874);
and U2089 (N_2089,N_1922,N_1896);
nand U2090 (N_2090,N_1986,N_1817);
nand U2091 (N_2091,N_1957,N_1982);
or U2092 (N_2092,N_1629,N_1934);
xor U2093 (N_2093,N_1908,N_1664);
and U2094 (N_2094,N_1862,N_1609);
and U2095 (N_2095,N_1678,N_1803);
nand U2096 (N_2096,N_1622,N_1654);
and U2097 (N_2097,N_1975,N_1939);
or U2098 (N_2098,N_1600,N_1684);
xnor U2099 (N_2099,N_1646,N_1647);
nor U2100 (N_2100,N_1606,N_1740);
nand U2101 (N_2101,N_1865,N_1878);
xor U2102 (N_2102,N_1968,N_1978);
nand U2103 (N_2103,N_1676,N_1668);
or U2104 (N_2104,N_1759,N_1748);
nor U2105 (N_2105,N_1866,N_1671);
or U2106 (N_2106,N_1845,N_1747);
nor U2107 (N_2107,N_1838,N_1932);
or U2108 (N_2108,N_1805,N_1988);
xor U2109 (N_2109,N_1888,N_1785);
nand U2110 (N_2110,N_1667,N_1882);
nand U2111 (N_2111,N_1742,N_1611);
xnor U2112 (N_2112,N_1921,N_1861);
or U2113 (N_2113,N_1956,N_1706);
or U2114 (N_2114,N_1750,N_1990);
and U2115 (N_2115,N_1858,N_1987);
and U2116 (N_2116,N_1885,N_1835);
and U2117 (N_2117,N_1784,N_1630);
or U2118 (N_2118,N_1812,N_1940);
or U2119 (N_2119,N_1607,N_1625);
nor U2120 (N_2120,N_1746,N_1913);
or U2121 (N_2121,N_1955,N_1744);
or U2122 (N_2122,N_1947,N_1645);
xor U2123 (N_2123,N_1780,N_1604);
or U2124 (N_2124,N_1621,N_1942);
and U2125 (N_2125,N_1977,N_1949);
and U2126 (N_2126,N_1904,N_1655);
or U2127 (N_2127,N_1962,N_1966);
or U2128 (N_2128,N_1700,N_1729);
nand U2129 (N_2129,N_1924,N_1895);
or U2130 (N_2130,N_1914,N_1704);
and U2131 (N_2131,N_1786,N_1815);
nand U2132 (N_2132,N_1826,N_1713);
or U2133 (N_2133,N_1991,N_1781);
and U2134 (N_2134,N_1795,N_1753);
and U2135 (N_2135,N_1765,N_1719);
xor U2136 (N_2136,N_1976,N_1751);
nand U2137 (N_2137,N_1900,N_1899);
xnor U2138 (N_2138,N_1769,N_1834);
and U2139 (N_2139,N_1854,N_1849);
nor U2140 (N_2140,N_1807,N_1761);
nor U2141 (N_2141,N_1791,N_1970);
or U2142 (N_2142,N_1626,N_1675);
and U2143 (N_2143,N_1873,N_1708);
nor U2144 (N_2144,N_1946,N_1738);
and U2145 (N_2145,N_1941,N_1794);
nand U2146 (N_2146,N_1731,N_1810);
and U2147 (N_2147,N_1674,N_1725);
or U2148 (N_2148,N_1608,N_1722);
nand U2149 (N_2149,N_1619,N_1733);
and U2150 (N_2150,N_1633,N_1662);
xnor U2151 (N_2151,N_1648,N_1743);
nand U2152 (N_2152,N_1863,N_1756);
nand U2153 (N_2153,N_1612,N_1613);
nor U2154 (N_2154,N_1848,N_1843);
xnor U2155 (N_2155,N_1816,N_1677);
and U2156 (N_2156,N_1670,N_1617);
nor U2157 (N_2157,N_1651,N_1790);
or U2158 (N_2158,N_1980,N_1623);
and U2159 (N_2159,N_1797,N_1886);
nand U2160 (N_2160,N_1685,N_1767);
xor U2161 (N_2161,N_1762,N_1820);
nor U2162 (N_2162,N_1928,N_1937);
nor U2163 (N_2163,N_1936,N_1657);
nor U2164 (N_2164,N_1641,N_1766);
nor U2165 (N_2165,N_1850,N_1869);
nor U2166 (N_2166,N_1999,N_1757);
or U2167 (N_2167,N_1709,N_1909);
or U2168 (N_2168,N_1787,N_1984);
or U2169 (N_2169,N_1998,N_1907);
nor U2170 (N_2170,N_1839,N_1881);
nand U2171 (N_2171,N_1958,N_1856);
nand U2172 (N_2172,N_1891,N_1971);
nor U2173 (N_2173,N_1912,N_1726);
nand U2174 (N_2174,N_1779,N_1690);
and U2175 (N_2175,N_1811,N_1930);
xor U2176 (N_2176,N_1964,N_1702);
nor U2177 (N_2177,N_1754,N_1833);
nand U2178 (N_2178,N_1763,N_1697);
nand U2179 (N_2179,N_1974,N_1673);
or U2180 (N_2180,N_1723,N_1960);
and U2181 (N_2181,N_1852,N_1972);
xor U2182 (N_2182,N_1792,N_1721);
nand U2183 (N_2183,N_1959,N_1981);
or U2184 (N_2184,N_1952,N_1911);
nor U2185 (N_2185,N_1844,N_1846);
nor U2186 (N_2186,N_1720,N_1618);
and U2187 (N_2187,N_1710,N_1944);
or U2188 (N_2188,N_1693,N_1716);
xor U2189 (N_2189,N_1760,N_1995);
and U2190 (N_2190,N_1920,N_1933);
nor U2191 (N_2191,N_1718,N_1665);
xor U2192 (N_2192,N_1857,N_1614);
and U2193 (N_2193,N_1925,N_1967);
nand U2194 (N_2194,N_1649,N_1616);
nor U2195 (N_2195,N_1661,N_1798);
and U2196 (N_2196,N_1969,N_1950);
xor U2197 (N_2197,N_1659,N_1715);
nor U2198 (N_2198,N_1681,N_1832);
nor U2199 (N_2199,N_1695,N_1637);
xor U2200 (N_2200,N_1791,N_1700);
xor U2201 (N_2201,N_1978,N_1783);
or U2202 (N_2202,N_1668,N_1893);
nand U2203 (N_2203,N_1827,N_1741);
and U2204 (N_2204,N_1834,N_1785);
xor U2205 (N_2205,N_1714,N_1664);
or U2206 (N_2206,N_1987,N_1606);
nand U2207 (N_2207,N_1795,N_1683);
nand U2208 (N_2208,N_1939,N_1789);
nand U2209 (N_2209,N_1881,N_1880);
and U2210 (N_2210,N_1960,N_1780);
and U2211 (N_2211,N_1647,N_1975);
xnor U2212 (N_2212,N_1953,N_1787);
nand U2213 (N_2213,N_1730,N_1788);
xnor U2214 (N_2214,N_1895,N_1715);
or U2215 (N_2215,N_1918,N_1926);
and U2216 (N_2216,N_1714,N_1729);
nand U2217 (N_2217,N_1749,N_1815);
nand U2218 (N_2218,N_1763,N_1992);
and U2219 (N_2219,N_1708,N_1881);
and U2220 (N_2220,N_1612,N_1601);
and U2221 (N_2221,N_1688,N_1729);
nand U2222 (N_2222,N_1762,N_1833);
xor U2223 (N_2223,N_1742,N_1916);
nand U2224 (N_2224,N_1861,N_1647);
nand U2225 (N_2225,N_1852,N_1743);
xor U2226 (N_2226,N_1902,N_1765);
or U2227 (N_2227,N_1924,N_1934);
nor U2228 (N_2228,N_1970,N_1694);
or U2229 (N_2229,N_1717,N_1853);
nor U2230 (N_2230,N_1682,N_1870);
nand U2231 (N_2231,N_1991,N_1615);
or U2232 (N_2232,N_1653,N_1868);
or U2233 (N_2233,N_1717,N_1956);
nand U2234 (N_2234,N_1625,N_1753);
nand U2235 (N_2235,N_1655,N_1997);
and U2236 (N_2236,N_1661,N_1897);
and U2237 (N_2237,N_1978,N_1730);
or U2238 (N_2238,N_1631,N_1921);
nor U2239 (N_2239,N_1708,N_1717);
nand U2240 (N_2240,N_1893,N_1662);
nor U2241 (N_2241,N_1906,N_1837);
and U2242 (N_2242,N_1693,N_1930);
and U2243 (N_2243,N_1873,N_1874);
nor U2244 (N_2244,N_1849,N_1926);
and U2245 (N_2245,N_1949,N_1835);
or U2246 (N_2246,N_1669,N_1998);
or U2247 (N_2247,N_1631,N_1714);
xnor U2248 (N_2248,N_1832,N_1642);
or U2249 (N_2249,N_1742,N_1709);
nand U2250 (N_2250,N_1951,N_1931);
and U2251 (N_2251,N_1863,N_1859);
nor U2252 (N_2252,N_1917,N_1613);
and U2253 (N_2253,N_1948,N_1915);
nor U2254 (N_2254,N_1867,N_1704);
nand U2255 (N_2255,N_1830,N_1995);
or U2256 (N_2256,N_1810,N_1642);
nand U2257 (N_2257,N_1856,N_1778);
xor U2258 (N_2258,N_1625,N_1898);
and U2259 (N_2259,N_1612,N_1985);
or U2260 (N_2260,N_1816,N_1940);
nand U2261 (N_2261,N_1934,N_1965);
xor U2262 (N_2262,N_1780,N_1906);
xnor U2263 (N_2263,N_1818,N_1792);
nand U2264 (N_2264,N_1866,N_1840);
xnor U2265 (N_2265,N_1639,N_1911);
nand U2266 (N_2266,N_1921,N_1917);
or U2267 (N_2267,N_1779,N_1908);
nand U2268 (N_2268,N_1919,N_1907);
and U2269 (N_2269,N_1954,N_1703);
and U2270 (N_2270,N_1838,N_1794);
nand U2271 (N_2271,N_1973,N_1748);
nor U2272 (N_2272,N_1772,N_1712);
nand U2273 (N_2273,N_1602,N_1623);
or U2274 (N_2274,N_1904,N_1895);
and U2275 (N_2275,N_1769,N_1673);
nor U2276 (N_2276,N_1974,N_1861);
and U2277 (N_2277,N_1740,N_1961);
nand U2278 (N_2278,N_1993,N_1747);
or U2279 (N_2279,N_1952,N_1724);
nor U2280 (N_2280,N_1972,N_1749);
xor U2281 (N_2281,N_1852,N_1731);
nor U2282 (N_2282,N_1772,N_1738);
nand U2283 (N_2283,N_1920,N_1662);
and U2284 (N_2284,N_1839,N_1963);
or U2285 (N_2285,N_1829,N_1765);
and U2286 (N_2286,N_1789,N_1830);
or U2287 (N_2287,N_1994,N_1838);
or U2288 (N_2288,N_1699,N_1706);
xor U2289 (N_2289,N_1923,N_1877);
xor U2290 (N_2290,N_1807,N_1866);
nand U2291 (N_2291,N_1714,N_1771);
xnor U2292 (N_2292,N_1643,N_1766);
or U2293 (N_2293,N_1918,N_1623);
nand U2294 (N_2294,N_1653,N_1931);
nor U2295 (N_2295,N_1931,N_1801);
nand U2296 (N_2296,N_1998,N_1789);
xnor U2297 (N_2297,N_1821,N_1973);
xnor U2298 (N_2298,N_1990,N_1724);
nand U2299 (N_2299,N_1960,N_1867);
nand U2300 (N_2300,N_1967,N_1657);
xor U2301 (N_2301,N_1912,N_1975);
and U2302 (N_2302,N_1794,N_1896);
and U2303 (N_2303,N_1657,N_1933);
and U2304 (N_2304,N_1729,N_1963);
or U2305 (N_2305,N_1815,N_1927);
nor U2306 (N_2306,N_1774,N_1993);
xnor U2307 (N_2307,N_1973,N_1879);
xor U2308 (N_2308,N_1894,N_1697);
nand U2309 (N_2309,N_1859,N_1720);
and U2310 (N_2310,N_1991,N_1713);
xor U2311 (N_2311,N_1682,N_1912);
nand U2312 (N_2312,N_1649,N_1700);
or U2313 (N_2313,N_1627,N_1729);
nor U2314 (N_2314,N_1809,N_1934);
nor U2315 (N_2315,N_1899,N_1693);
or U2316 (N_2316,N_1917,N_1763);
nor U2317 (N_2317,N_1857,N_1769);
xor U2318 (N_2318,N_1974,N_1917);
or U2319 (N_2319,N_1947,N_1702);
nand U2320 (N_2320,N_1701,N_1736);
xor U2321 (N_2321,N_1769,N_1615);
nor U2322 (N_2322,N_1754,N_1912);
xnor U2323 (N_2323,N_1611,N_1797);
and U2324 (N_2324,N_1983,N_1879);
and U2325 (N_2325,N_1989,N_1965);
or U2326 (N_2326,N_1760,N_1769);
nand U2327 (N_2327,N_1748,N_1648);
nor U2328 (N_2328,N_1680,N_1811);
and U2329 (N_2329,N_1923,N_1717);
xnor U2330 (N_2330,N_1653,N_1819);
nand U2331 (N_2331,N_1630,N_1995);
xor U2332 (N_2332,N_1772,N_1677);
xor U2333 (N_2333,N_1915,N_1919);
xnor U2334 (N_2334,N_1766,N_1828);
and U2335 (N_2335,N_1867,N_1644);
and U2336 (N_2336,N_1980,N_1717);
or U2337 (N_2337,N_1828,N_1950);
xnor U2338 (N_2338,N_1754,N_1987);
nand U2339 (N_2339,N_1731,N_1798);
nor U2340 (N_2340,N_1645,N_1725);
xnor U2341 (N_2341,N_1740,N_1710);
or U2342 (N_2342,N_1957,N_1712);
or U2343 (N_2343,N_1762,N_1948);
and U2344 (N_2344,N_1828,N_1701);
and U2345 (N_2345,N_1774,N_1734);
nor U2346 (N_2346,N_1828,N_1714);
or U2347 (N_2347,N_1610,N_1666);
or U2348 (N_2348,N_1876,N_1657);
xnor U2349 (N_2349,N_1697,N_1786);
nand U2350 (N_2350,N_1780,N_1612);
nor U2351 (N_2351,N_1864,N_1619);
or U2352 (N_2352,N_1830,N_1794);
and U2353 (N_2353,N_1789,N_1619);
or U2354 (N_2354,N_1917,N_1793);
or U2355 (N_2355,N_1809,N_1853);
or U2356 (N_2356,N_1785,N_1938);
nand U2357 (N_2357,N_1694,N_1817);
nand U2358 (N_2358,N_1601,N_1992);
xnor U2359 (N_2359,N_1887,N_1705);
xnor U2360 (N_2360,N_1985,N_1649);
or U2361 (N_2361,N_1963,N_1889);
or U2362 (N_2362,N_1767,N_1970);
xnor U2363 (N_2363,N_1959,N_1777);
and U2364 (N_2364,N_1955,N_1760);
nand U2365 (N_2365,N_1755,N_1632);
xor U2366 (N_2366,N_1808,N_1771);
nor U2367 (N_2367,N_1860,N_1648);
and U2368 (N_2368,N_1750,N_1908);
nand U2369 (N_2369,N_1750,N_1807);
and U2370 (N_2370,N_1905,N_1668);
and U2371 (N_2371,N_1970,N_1677);
or U2372 (N_2372,N_1646,N_1972);
xnor U2373 (N_2373,N_1815,N_1901);
nor U2374 (N_2374,N_1697,N_1856);
nor U2375 (N_2375,N_1729,N_1657);
and U2376 (N_2376,N_1962,N_1716);
or U2377 (N_2377,N_1772,N_1732);
and U2378 (N_2378,N_1928,N_1666);
nor U2379 (N_2379,N_1658,N_1914);
nor U2380 (N_2380,N_1860,N_1836);
and U2381 (N_2381,N_1693,N_1621);
and U2382 (N_2382,N_1666,N_1806);
xnor U2383 (N_2383,N_1973,N_1883);
or U2384 (N_2384,N_1998,N_1796);
nor U2385 (N_2385,N_1761,N_1636);
xnor U2386 (N_2386,N_1678,N_1715);
and U2387 (N_2387,N_1993,N_1978);
and U2388 (N_2388,N_1707,N_1788);
or U2389 (N_2389,N_1969,N_1958);
nand U2390 (N_2390,N_1950,N_1642);
nor U2391 (N_2391,N_1854,N_1730);
and U2392 (N_2392,N_1830,N_1893);
xor U2393 (N_2393,N_1893,N_1634);
nand U2394 (N_2394,N_1853,N_1739);
nor U2395 (N_2395,N_1738,N_1871);
nor U2396 (N_2396,N_1968,N_1679);
or U2397 (N_2397,N_1942,N_1863);
or U2398 (N_2398,N_1815,N_1625);
or U2399 (N_2399,N_1951,N_1846);
nor U2400 (N_2400,N_2060,N_2368);
nand U2401 (N_2401,N_2205,N_2260);
and U2402 (N_2402,N_2176,N_2316);
nor U2403 (N_2403,N_2083,N_2197);
or U2404 (N_2404,N_2158,N_2146);
xnor U2405 (N_2405,N_2072,N_2134);
xor U2406 (N_2406,N_2399,N_2355);
or U2407 (N_2407,N_2321,N_2221);
xor U2408 (N_2408,N_2335,N_2137);
nand U2409 (N_2409,N_2129,N_2374);
and U2410 (N_2410,N_2286,N_2087);
nand U2411 (N_2411,N_2284,N_2163);
and U2412 (N_2412,N_2034,N_2073);
nand U2413 (N_2413,N_2192,N_2128);
or U2414 (N_2414,N_2104,N_2045);
nor U2415 (N_2415,N_2081,N_2040);
and U2416 (N_2416,N_2113,N_2080);
xor U2417 (N_2417,N_2255,N_2082);
nor U2418 (N_2418,N_2145,N_2002);
nand U2419 (N_2419,N_2085,N_2035);
xnor U2420 (N_2420,N_2195,N_2244);
xnor U2421 (N_2421,N_2300,N_2105);
nor U2422 (N_2422,N_2165,N_2025);
xor U2423 (N_2423,N_2102,N_2161);
and U2424 (N_2424,N_2396,N_2347);
xnor U2425 (N_2425,N_2276,N_2089);
or U2426 (N_2426,N_2175,N_2078);
nand U2427 (N_2427,N_2182,N_2301);
and U2428 (N_2428,N_2314,N_2190);
or U2429 (N_2429,N_2203,N_2055);
and U2430 (N_2430,N_2044,N_2001);
and U2431 (N_2431,N_2006,N_2220);
and U2432 (N_2432,N_2262,N_2224);
or U2433 (N_2433,N_2343,N_2223);
and U2434 (N_2434,N_2144,N_2273);
xnor U2435 (N_2435,N_2028,N_2349);
or U2436 (N_2436,N_2313,N_2373);
and U2437 (N_2437,N_2041,N_2050);
xnor U2438 (N_2438,N_2333,N_2246);
nor U2439 (N_2439,N_2193,N_2160);
or U2440 (N_2440,N_2210,N_2027);
nand U2441 (N_2441,N_2334,N_2249);
nor U2442 (N_2442,N_2005,N_2215);
xnor U2443 (N_2443,N_2311,N_2365);
nor U2444 (N_2444,N_2213,N_2381);
nor U2445 (N_2445,N_2162,N_2394);
xnor U2446 (N_2446,N_2047,N_2339);
nor U2447 (N_2447,N_2397,N_2164);
and U2448 (N_2448,N_2004,N_2065);
or U2449 (N_2449,N_2388,N_2098);
and U2450 (N_2450,N_2125,N_2283);
or U2451 (N_2451,N_2243,N_2212);
or U2452 (N_2452,N_2299,N_2180);
xnor U2453 (N_2453,N_2337,N_2013);
or U2454 (N_2454,N_2222,N_2174);
and U2455 (N_2455,N_2353,N_2076);
xnor U2456 (N_2456,N_2068,N_2110);
nor U2457 (N_2457,N_2209,N_2239);
xor U2458 (N_2458,N_2189,N_2183);
or U2459 (N_2459,N_2207,N_2282);
or U2460 (N_2460,N_2367,N_2166);
xnor U2461 (N_2461,N_2218,N_2070);
and U2462 (N_2462,N_2277,N_2188);
and U2463 (N_2463,N_2201,N_2066);
and U2464 (N_2464,N_2024,N_2122);
xor U2465 (N_2465,N_2360,N_2115);
and U2466 (N_2466,N_2154,N_2121);
nor U2467 (N_2467,N_2211,N_2395);
nand U2468 (N_2468,N_2235,N_2305);
nand U2469 (N_2469,N_2214,N_2196);
or U2470 (N_2470,N_2018,N_2118);
nand U2471 (N_2471,N_2320,N_2285);
or U2472 (N_2472,N_2170,N_2251);
nand U2473 (N_2473,N_2185,N_2023);
nand U2474 (N_2474,N_2269,N_2309);
or U2475 (N_2475,N_2229,N_2140);
xnor U2476 (N_2476,N_2017,N_2238);
or U2477 (N_2477,N_2356,N_2369);
and U2478 (N_2478,N_2342,N_2323);
nor U2479 (N_2479,N_2088,N_2053);
nor U2480 (N_2480,N_2265,N_2109);
nor U2481 (N_2481,N_2217,N_2268);
and U2482 (N_2482,N_2206,N_2131);
nor U2483 (N_2483,N_2370,N_2330);
and U2484 (N_2484,N_2363,N_2091);
xor U2485 (N_2485,N_2127,N_2296);
or U2486 (N_2486,N_2142,N_2208);
nand U2487 (N_2487,N_2227,N_2147);
nand U2488 (N_2488,N_2271,N_2107);
nand U2489 (N_2489,N_2312,N_2124);
xor U2490 (N_2490,N_2219,N_2287);
or U2491 (N_2491,N_2303,N_2346);
nor U2492 (N_2492,N_2240,N_2295);
xor U2493 (N_2493,N_2380,N_2186);
nor U2494 (N_2494,N_2059,N_2058);
or U2495 (N_2495,N_2371,N_2332);
nand U2496 (N_2496,N_2226,N_2184);
nor U2497 (N_2497,N_2338,N_2015);
xor U2498 (N_2498,N_2138,N_2084);
and U2499 (N_2499,N_2278,N_2069);
nand U2500 (N_2500,N_2362,N_2079);
xor U2501 (N_2501,N_2225,N_2272);
and U2502 (N_2502,N_2386,N_2198);
xnor U2503 (N_2503,N_2351,N_2293);
nand U2504 (N_2504,N_2061,N_2011);
and U2505 (N_2505,N_2012,N_2385);
nor U2506 (N_2506,N_2359,N_2019);
nor U2507 (N_2507,N_2191,N_2031);
or U2508 (N_2508,N_2324,N_2086);
nand U2509 (N_2509,N_2094,N_2008);
and U2510 (N_2510,N_2156,N_2052);
nand U2511 (N_2511,N_2391,N_2248);
xnor U2512 (N_2512,N_2003,N_2267);
and U2513 (N_2513,N_2171,N_2111);
xor U2514 (N_2514,N_2100,N_2384);
xor U2515 (N_2515,N_2092,N_2049);
or U2516 (N_2516,N_2114,N_2062);
and U2517 (N_2517,N_2204,N_2143);
xnor U2518 (N_2518,N_2231,N_2039);
nor U2519 (N_2519,N_2043,N_2064);
nor U2520 (N_2520,N_2292,N_2009);
and U2521 (N_2521,N_2095,N_2241);
nand U2522 (N_2522,N_2310,N_2177);
or U2523 (N_2523,N_2152,N_2390);
nor U2524 (N_2524,N_2297,N_2315);
xnor U2525 (N_2525,N_2232,N_2281);
nand U2526 (N_2526,N_2392,N_2307);
nand U2527 (N_2527,N_2126,N_2357);
nor U2528 (N_2528,N_2000,N_2033);
xor U2529 (N_2529,N_2364,N_2187);
nor U2530 (N_2530,N_2266,N_2151);
and U2531 (N_2531,N_2378,N_2074);
and U2532 (N_2532,N_2096,N_2148);
or U2533 (N_2533,N_2294,N_2398);
nor U2534 (N_2534,N_2132,N_2366);
nand U2535 (N_2535,N_2030,N_2010);
nor U2536 (N_2536,N_2067,N_2341);
or U2537 (N_2537,N_2179,N_2093);
xnor U2538 (N_2538,N_2135,N_2327);
and U2539 (N_2539,N_2375,N_2014);
nor U2540 (N_2540,N_2336,N_2358);
xor U2541 (N_2541,N_2036,N_2106);
and U2542 (N_2542,N_2288,N_2291);
nand U2543 (N_2543,N_2331,N_2150);
nand U2544 (N_2544,N_2290,N_2117);
xor U2545 (N_2545,N_2306,N_2382);
and U2546 (N_2546,N_2167,N_2236);
nand U2547 (N_2547,N_2377,N_2157);
xnor U2548 (N_2548,N_2200,N_2199);
nor U2549 (N_2549,N_2021,N_2063);
nor U2550 (N_2550,N_2259,N_2046);
nand U2551 (N_2551,N_2354,N_2141);
nand U2552 (N_2552,N_2340,N_2274);
and U2553 (N_2553,N_2181,N_2112);
xor U2554 (N_2554,N_2233,N_2298);
nor U2555 (N_2555,N_2123,N_2099);
or U2556 (N_2556,N_2302,N_2257);
or U2557 (N_2557,N_2228,N_2242);
and U2558 (N_2558,N_2376,N_2261);
nor U2559 (N_2559,N_2056,N_2350);
and U2560 (N_2560,N_2383,N_2270);
and U2561 (N_2561,N_2263,N_2130);
xor U2562 (N_2562,N_2032,N_2352);
nand U2563 (N_2563,N_2252,N_2054);
nand U2564 (N_2564,N_2318,N_2139);
nor U2565 (N_2565,N_2389,N_2256);
nand U2566 (N_2566,N_2379,N_2326);
and U2567 (N_2567,N_2254,N_2234);
or U2568 (N_2568,N_2328,N_2387);
or U2569 (N_2569,N_2230,N_2325);
nand U2570 (N_2570,N_2250,N_2022);
nor U2571 (N_2571,N_2097,N_2178);
nand U2572 (N_2572,N_2101,N_2202);
nand U2573 (N_2573,N_2247,N_2361);
and U2574 (N_2574,N_2042,N_2264);
or U2575 (N_2575,N_2169,N_2133);
nor U2576 (N_2576,N_2155,N_2304);
and U2577 (N_2577,N_2159,N_2279);
nor U2578 (N_2578,N_2194,N_2319);
nor U2579 (N_2579,N_2393,N_2016);
xnor U2580 (N_2580,N_2037,N_2172);
xor U2581 (N_2581,N_2308,N_2020);
xor U2582 (N_2582,N_2071,N_2153);
and U2583 (N_2583,N_2051,N_2322);
xor U2584 (N_2584,N_2329,N_2253);
and U2585 (N_2585,N_2372,N_2120);
or U2586 (N_2586,N_2007,N_2289);
nor U2587 (N_2587,N_2216,N_2168);
nand U2588 (N_2588,N_2245,N_2136);
nor U2589 (N_2589,N_2077,N_2344);
or U2590 (N_2590,N_2149,N_2026);
xor U2591 (N_2591,N_2090,N_2038);
nor U2592 (N_2592,N_2048,N_2057);
xnor U2593 (N_2593,N_2348,N_2103);
or U2594 (N_2594,N_2119,N_2075);
xor U2595 (N_2595,N_2108,N_2173);
or U2596 (N_2596,N_2275,N_2345);
nor U2597 (N_2597,N_2116,N_2317);
nand U2598 (N_2598,N_2258,N_2237);
nor U2599 (N_2599,N_2029,N_2280);
or U2600 (N_2600,N_2258,N_2298);
or U2601 (N_2601,N_2337,N_2226);
xnor U2602 (N_2602,N_2104,N_2375);
nand U2603 (N_2603,N_2234,N_2042);
nor U2604 (N_2604,N_2138,N_2223);
or U2605 (N_2605,N_2006,N_2157);
and U2606 (N_2606,N_2130,N_2356);
or U2607 (N_2607,N_2253,N_2062);
or U2608 (N_2608,N_2076,N_2382);
nor U2609 (N_2609,N_2144,N_2195);
nor U2610 (N_2610,N_2124,N_2355);
nand U2611 (N_2611,N_2316,N_2262);
and U2612 (N_2612,N_2301,N_2241);
and U2613 (N_2613,N_2128,N_2006);
nor U2614 (N_2614,N_2076,N_2197);
nand U2615 (N_2615,N_2396,N_2077);
and U2616 (N_2616,N_2069,N_2388);
and U2617 (N_2617,N_2028,N_2233);
xnor U2618 (N_2618,N_2164,N_2153);
nand U2619 (N_2619,N_2172,N_2114);
or U2620 (N_2620,N_2231,N_2188);
nand U2621 (N_2621,N_2334,N_2300);
nand U2622 (N_2622,N_2129,N_2130);
xnor U2623 (N_2623,N_2005,N_2127);
and U2624 (N_2624,N_2399,N_2123);
and U2625 (N_2625,N_2024,N_2219);
or U2626 (N_2626,N_2236,N_2221);
nand U2627 (N_2627,N_2346,N_2337);
xnor U2628 (N_2628,N_2175,N_2291);
nor U2629 (N_2629,N_2169,N_2342);
xor U2630 (N_2630,N_2027,N_2386);
and U2631 (N_2631,N_2201,N_2328);
nand U2632 (N_2632,N_2020,N_2162);
or U2633 (N_2633,N_2092,N_2042);
nand U2634 (N_2634,N_2129,N_2089);
or U2635 (N_2635,N_2083,N_2107);
nor U2636 (N_2636,N_2100,N_2357);
or U2637 (N_2637,N_2330,N_2087);
nand U2638 (N_2638,N_2240,N_2228);
and U2639 (N_2639,N_2399,N_2394);
or U2640 (N_2640,N_2270,N_2043);
nand U2641 (N_2641,N_2134,N_2222);
nor U2642 (N_2642,N_2323,N_2095);
and U2643 (N_2643,N_2124,N_2057);
and U2644 (N_2644,N_2241,N_2105);
xor U2645 (N_2645,N_2288,N_2340);
and U2646 (N_2646,N_2201,N_2178);
or U2647 (N_2647,N_2342,N_2043);
xnor U2648 (N_2648,N_2212,N_2204);
xor U2649 (N_2649,N_2029,N_2372);
nand U2650 (N_2650,N_2284,N_2184);
xor U2651 (N_2651,N_2053,N_2037);
or U2652 (N_2652,N_2161,N_2247);
nor U2653 (N_2653,N_2158,N_2137);
xnor U2654 (N_2654,N_2017,N_2388);
and U2655 (N_2655,N_2085,N_2362);
nor U2656 (N_2656,N_2157,N_2052);
and U2657 (N_2657,N_2249,N_2363);
xnor U2658 (N_2658,N_2120,N_2333);
or U2659 (N_2659,N_2246,N_2113);
or U2660 (N_2660,N_2176,N_2283);
and U2661 (N_2661,N_2371,N_2340);
and U2662 (N_2662,N_2091,N_2098);
xnor U2663 (N_2663,N_2085,N_2093);
nor U2664 (N_2664,N_2015,N_2373);
nand U2665 (N_2665,N_2157,N_2373);
or U2666 (N_2666,N_2001,N_2299);
nor U2667 (N_2667,N_2320,N_2101);
or U2668 (N_2668,N_2256,N_2352);
nand U2669 (N_2669,N_2109,N_2226);
nand U2670 (N_2670,N_2357,N_2293);
and U2671 (N_2671,N_2134,N_2375);
and U2672 (N_2672,N_2178,N_2253);
nand U2673 (N_2673,N_2159,N_2262);
and U2674 (N_2674,N_2168,N_2110);
and U2675 (N_2675,N_2096,N_2340);
or U2676 (N_2676,N_2095,N_2086);
or U2677 (N_2677,N_2092,N_2345);
nand U2678 (N_2678,N_2068,N_2297);
xor U2679 (N_2679,N_2177,N_2294);
nand U2680 (N_2680,N_2264,N_2113);
nor U2681 (N_2681,N_2210,N_2193);
xor U2682 (N_2682,N_2335,N_2162);
xnor U2683 (N_2683,N_2134,N_2255);
xor U2684 (N_2684,N_2213,N_2243);
nand U2685 (N_2685,N_2096,N_2198);
nor U2686 (N_2686,N_2198,N_2106);
nand U2687 (N_2687,N_2294,N_2370);
or U2688 (N_2688,N_2340,N_2225);
and U2689 (N_2689,N_2098,N_2169);
or U2690 (N_2690,N_2003,N_2157);
or U2691 (N_2691,N_2104,N_2374);
xor U2692 (N_2692,N_2170,N_2106);
nand U2693 (N_2693,N_2119,N_2224);
or U2694 (N_2694,N_2227,N_2185);
or U2695 (N_2695,N_2366,N_2099);
nor U2696 (N_2696,N_2164,N_2393);
xnor U2697 (N_2697,N_2337,N_2093);
and U2698 (N_2698,N_2209,N_2148);
or U2699 (N_2699,N_2175,N_2250);
nand U2700 (N_2700,N_2022,N_2399);
nand U2701 (N_2701,N_2039,N_2325);
xor U2702 (N_2702,N_2270,N_2164);
or U2703 (N_2703,N_2394,N_2183);
nand U2704 (N_2704,N_2314,N_2163);
or U2705 (N_2705,N_2199,N_2246);
xnor U2706 (N_2706,N_2268,N_2048);
xor U2707 (N_2707,N_2314,N_2067);
nand U2708 (N_2708,N_2175,N_2272);
nand U2709 (N_2709,N_2253,N_2338);
xnor U2710 (N_2710,N_2248,N_2079);
nor U2711 (N_2711,N_2245,N_2157);
xor U2712 (N_2712,N_2007,N_2211);
or U2713 (N_2713,N_2315,N_2249);
or U2714 (N_2714,N_2283,N_2203);
or U2715 (N_2715,N_2309,N_2004);
or U2716 (N_2716,N_2188,N_2258);
nand U2717 (N_2717,N_2257,N_2182);
and U2718 (N_2718,N_2167,N_2177);
nand U2719 (N_2719,N_2234,N_2319);
nor U2720 (N_2720,N_2345,N_2304);
and U2721 (N_2721,N_2085,N_2083);
or U2722 (N_2722,N_2211,N_2040);
nor U2723 (N_2723,N_2216,N_2229);
nor U2724 (N_2724,N_2188,N_2217);
xor U2725 (N_2725,N_2094,N_2076);
nor U2726 (N_2726,N_2305,N_2315);
and U2727 (N_2727,N_2311,N_2175);
or U2728 (N_2728,N_2100,N_2090);
and U2729 (N_2729,N_2000,N_2090);
or U2730 (N_2730,N_2190,N_2235);
nor U2731 (N_2731,N_2369,N_2348);
nor U2732 (N_2732,N_2018,N_2059);
nor U2733 (N_2733,N_2063,N_2277);
nand U2734 (N_2734,N_2261,N_2168);
or U2735 (N_2735,N_2323,N_2014);
xnor U2736 (N_2736,N_2323,N_2233);
nor U2737 (N_2737,N_2309,N_2247);
xnor U2738 (N_2738,N_2057,N_2216);
nand U2739 (N_2739,N_2124,N_2171);
nor U2740 (N_2740,N_2037,N_2397);
nor U2741 (N_2741,N_2049,N_2154);
nor U2742 (N_2742,N_2389,N_2277);
xnor U2743 (N_2743,N_2295,N_2223);
or U2744 (N_2744,N_2288,N_2182);
and U2745 (N_2745,N_2353,N_2338);
nand U2746 (N_2746,N_2292,N_2342);
xnor U2747 (N_2747,N_2239,N_2117);
or U2748 (N_2748,N_2158,N_2059);
and U2749 (N_2749,N_2161,N_2000);
and U2750 (N_2750,N_2114,N_2386);
nor U2751 (N_2751,N_2088,N_2241);
xnor U2752 (N_2752,N_2183,N_2247);
nor U2753 (N_2753,N_2223,N_2162);
xor U2754 (N_2754,N_2013,N_2331);
and U2755 (N_2755,N_2051,N_2156);
and U2756 (N_2756,N_2225,N_2309);
and U2757 (N_2757,N_2378,N_2349);
and U2758 (N_2758,N_2306,N_2002);
or U2759 (N_2759,N_2168,N_2160);
nor U2760 (N_2760,N_2278,N_2144);
xor U2761 (N_2761,N_2185,N_2396);
and U2762 (N_2762,N_2049,N_2261);
or U2763 (N_2763,N_2320,N_2124);
and U2764 (N_2764,N_2308,N_2286);
nand U2765 (N_2765,N_2111,N_2154);
or U2766 (N_2766,N_2243,N_2175);
or U2767 (N_2767,N_2315,N_2384);
nand U2768 (N_2768,N_2025,N_2111);
xor U2769 (N_2769,N_2269,N_2105);
and U2770 (N_2770,N_2196,N_2206);
nand U2771 (N_2771,N_2245,N_2142);
or U2772 (N_2772,N_2022,N_2354);
or U2773 (N_2773,N_2360,N_2342);
and U2774 (N_2774,N_2037,N_2133);
nor U2775 (N_2775,N_2136,N_2007);
nand U2776 (N_2776,N_2296,N_2300);
nor U2777 (N_2777,N_2023,N_2345);
or U2778 (N_2778,N_2315,N_2206);
nand U2779 (N_2779,N_2201,N_2089);
and U2780 (N_2780,N_2246,N_2202);
nand U2781 (N_2781,N_2012,N_2231);
or U2782 (N_2782,N_2015,N_2331);
nor U2783 (N_2783,N_2014,N_2134);
nand U2784 (N_2784,N_2037,N_2016);
nand U2785 (N_2785,N_2254,N_2390);
or U2786 (N_2786,N_2114,N_2352);
nor U2787 (N_2787,N_2278,N_2171);
nor U2788 (N_2788,N_2342,N_2023);
nor U2789 (N_2789,N_2322,N_2399);
nand U2790 (N_2790,N_2283,N_2360);
and U2791 (N_2791,N_2187,N_2198);
or U2792 (N_2792,N_2225,N_2339);
or U2793 (N_2793,N_2374,N_2353);
nor U2794 (N_2794,N_2208,N_2217);
and U2795 (N_2795,N_2148,N_2013);
nand U2796 (N_2796,N_2294,N_2328);
and U2797 (N_2797,N_2100,N_2324);
nor U2798 (N_2798,N_2005,N_2210);
and U2799 (N_2799,N_2257,N_2100);
xnor U2800 (N_2800,N_2767,N_2597);
nand U2801 (N_2801,N_2666,N_2604);
and U2802 (N_2802,N_2747,N_2710);
or U2803 (N_2803,N_2755,N_2403);
xnor U2804 (N_2804,N_2501,N_2646);
and U2805 (N_2805,N_2639,N_2749);
nor U2806 (N_2806,N_2557,N_2503);
nor U2807 (N_2807,N_2550,N_2561);
and U2808 (N_2808,N_2431,N_2434);
nor U2809 (N_2809,N_2697,N_2757);
xor U2810 (N_2810,N_2512,N_2536);
nor U2811 (N_2811,N_2762,N_2791);
xor U2812 (N_2812,N_2785,N_2740);
nand U2813 (N_2813,N_2407,N_2613);
xor U2814 (N_2814,N_2635,N_2753);
nor U2815 (N_2815,N_2717,N_2469);
nand U2816 (N_2816,N_2461,N_2544);
xor U2817 (N_2817,N_2578,N_2517);
xor U2818 (N_2818,N_2455,N_2584);
xnor U2819 (N_2819,N_2594,N_2577);
or U2820 (N_2820,N_2663,N_2445);
and U2821 (N_2821,N_2508,N_2644);
nand U2822 (N_2822,N_2502,N_2545);
xnor U2823 (N_2823,N_2532,N_2499);
and U2824 (N_2824,N_2721,N_2798);
or U2825 (N_2825,N_2625,N_2645);
or U2826 (N_2826,N_2631,N_2659);
and U2827 (N_2827,N_2700,N_2492);
nor U2828 (N_2828,N_2526,N_2795);
xor U2829 (N_2829,N_2706,N_2765);
or U2830 (N_2830,N_2680,N_2602);
xnor U2831 (N_2831,N_2539,N_2574);
xnor U2832 (N_2832,N_2596,N_2592);
and U2833 (N_2833,N_2648,N_2610);
and U2834 (N_2834,N_2588,N_2543);
and U2835 (N_2835,N_2522,N_2427);
or U2836 (N_2836,N_2519,N_2662);
and U2837 (N_2837,N_2770,N_2589);
nor U2838 (N_2838,N_2570,N_2443);
nor U2839 (N_2839,N_2579,N_2568);
nor U2840 (N_2840,N_2565,N_2473);
and U2841 (N_2841,N_2474,N_2695);
and U2842 (N_2842,N_2490,N_2690);
xnor U2843 (N_2843,N_2410,N_2673);
xor U2844 (N_2844,N_2677,N_2459);
or U2845 (N_2845,N_2601,N_2718);
xor U2846 (N_2846,N_2457,N_2513);
nor U2847 (N_2847,N_2716,N_2510);
nand U2848 (N_2848,N_2741,N_2616);
nor U2849 (N_2849,N_2612,N_2769);
or U2850 (N_2850,N_2679,N_2413);
and U2851 (N_2851,N_2701,N_2494);
nor U2852 (N_2852,N_2529,N_2754);
nand U2853 (N_2853,N_2689,N_2569);
nand U2854 (N_2854,N_2711,N_2524);
and U2855 (N_2855,N_2752,N_2630);
nand U2856 (N_2856,N_2655,N_2796);
xor U2857 (N_2857,N_2456,N_2731);
or U2858 (N_2858,N_2719,N_2500);
and U2859 (N_2859,N_2462,N_2507);
nand U2860 (N_2860,N_2555,N_2424);
xor U2861 (N_2861,N_2687,N_2436);
and U2862 (N_2862,N_2738,N_2627);
nor U2863 (N_2863,N_2575,N_2426);
nor U2864 (N_2864,N_2739,N_2748);
xnor U2865 (N_2865,N_2642,N_2771);
or U2866 (N_2866,N_2799,N_2476);
and U2867 (N_2867,N_2661,N_2651);
or U2868 (N_2868,N_2676,N_2732);
nand U2869 (N_2869,N_2538,N_2734);
nand U2870 (N_2870,N_2730,N_2636);
nor U2871 (N_2871,N_2783,N_2486);
nand U2872 (N_2872,N_2707,N_2685);
or U2873 (N_2873,N_2764,N_2566);
or U2874 (N_2874,N_2556,N_2735);
xor U2875 (N_2875,N_2599,N_2440);
and U2876 (N_2876,N_2609,N_2760);
and U2877 (N_2877,N_2743,N_2665);
xor U2878 (N_2878,N_2465,N_2514);
and U2879 (N_2879,N_2414,N_2729);
xor U2880 (N_2880,N_2678,N_2653);
and U2881 (N_2881,N_2515,N_2647);
and U2882 (N_2882,N_2422,N_2475);
or U2883 (N_2883,N_2758,N_2429);
xnor U2884 (N_2884,N_2726,N_2542);
xor U2885 (N_2885,N_2621,N_2400);
nand U2886 (N_2886,N_2571,N_2595);
nand U2887 (N_2887,N_2709,N_2782);
nand U2888 (N_2888,N_2606,N_2790);
or U2889 (N_2889,N_2691,N_2776);
nor U2890 (N_2890,N_2549,N_2447);
xnor U2891 (N_2891,N_2727,N_2547);
xor U2892 (N_2892,N_2591,N_2667);
and U2893 (N_2893,N_2437,N_2598);
nor U2894 (N_2894,N_2792,N_2686);
or U2895 (N_2895,N_2480,N_2643);
xor U2896 (N_2896,N_2699,N_2745);
nand U2897 (N_2897,N_2497,N_2696);
nor U2898 (N_2898,N_2546,N_2654);
xor U2899 (N_2899,N_2441,N_2681);
nor U2900 (N_2900,N_2506,N_2766);
or U2901 (N_2901,N_2493,N_2618);
or U2902 (N_2902,N_2423,N_2511);
nand U2903 (N_2903,N_2432,N_2778);
nor U2904 (N_2904,N_2797,N_2482);
xnor U2905 (N_2905,N_2684,N_2736);
and U2906 (N_2906,N_2786,N_2484);
and U2907 (N_2907,N_2672,N_2564);
or U2908 (N_2908,N_2585,N_2773);
nand U2909 (N_2909,N_2458,N_2603);
nor U2910 (N_2910,N_2420,N_2478);
or U2911 (N_2911,N_2438,N_2567);
xor U2912 (N_2912,N_2518,N_2664);
xor U2913 (N_2913,N_2611,N_2713);
or U2914 (N_2914,N_2638,N_2472);
and U2915 (N_2915,N_2504,N_2694);
or U2916 (N_2916,N_2608,N_2780);
or U2917 (N_2917,N_2516,N_2615);
nor U2918 (N_2918,N_2628,N_2537);
and U2919 (N_2919,N_2781,N_2406);
xnor U2920 (N_2920,N_2671,N_2471);
and U2921 (N_2921,N_2558,N_2725);
nand U2922 (N_2922,N_2415,N_2728);
and U2923 (N_2923,N_2590,N_2531);
xor U2924 (N_2924,N_2534,N_2626);
and U2925 (N_2925,N_2405,N_2450);
xnor U2926 (N_2926,N_2712,N_2614);
nand U2927 (N_2927,N_2402,N_2703);
nor U2928 (N_2928,N_2408,N_2487);
or U2929 (N_2929,N_2656,N_2620);
nor U2930 (N_2930,N_2793,N_2650);
and U2931 (N_2931,N_2768,N_2789);
nand U2932 (N_2932,N_2633,N_2533);
nor U2933 (N_2933,N_2724,N_2452);
xor U2934 (N_2934,N_2553,N_2525);
and U2935 (N_2935,N_2759,N_2756);
nand U2936 (N_2936,N_2401,N_2640);
or U2937 (N_2937,N_2583,N_2479);
xnor U2938 (N_2938,N_2698,N_2433);
or U2939 (N_2939,N_2488,N_2463);
and U2940 (N_2940,N_2714,N_2491);
and U2941 (N_2941,N_2468,N_2742);
and U2942 (N_2942,N_2586,N_2554);
or U2943 (N_2943,N_2404,N_2784);
or U2944 (N_2944,N_2419,N_2751);
nand U2945 (N_2945,N_2669,N_2541);
nand U2946 (N_2946,N_2505,N_2425);
and U2947 (N_2947,N_2788,N_2520);
and U2948 (N_2948,N_2466,N_2582);
xnor U2949 (N_2949,N_2551,N_2683);
nor U2950 (N_2950,N_2617,N_2600);
nor U2951 (N_2951,N_2411,N_2449);
and U2952 (N_2952,N_2622,N_2763);
nor U2953 (N_2953,N_2451,N_2435);
and U2954 (N_2954,N_2485,N_2715);
nor U2955 (N_2955,N_2439,N_2562);
or U2956 (N_2956,N_2668,N_2409);
xnor U2957 (N_2957,N_2623,N_2787);
nor U2958 (N_2958,N_2417,N_2708);
xnor U2959 (N_2959,N_2720,N_2675);
or U2960 (N_2960,N_2775,N_2464);
and U2961 (N_2961,N_2704,N_2552);
nor U2962 (N_2962,N_2774,N_2421);
nand U2963 (N_2963,N_2535,N_2746);
or U2964 (N_2964,N_2779,N_2495);
xnor U2965 (N_2965,N_2682,N_2772);
and U2966 (N_2966,N_2477,N_2607);
or U2967 (N_2967,N_2418,N_2528);
or U2968 (N_2968,N_2540,N_2498);
and U2969 (N_2969,N_2674,N_2560);
nand U2970 (N_2970,N_2460,N_2576);
xnor U2971 (N_2971,N_2652,N_2527);
nand U2972 (N_2972,N_2670,N_2641);
and U2973 (N_2973,N_2481,N_2572);
nand U2974 (N_2974,N_2548,N_2649);
xnor U2975 (N_2975,N_2521,N_2483);
or U2976 (N_2976,N_2777,N_2489);
nor U2977 (N_2977,N_2693,N_2761);
and U2978 (N_2978,N_2722,N_2750);
xnor U2979 (N_2979,N_2573,N_2509);
or U2980 (N_2980,N_2688,N_2737);
or U2981 (N_2981,N_2530,N_2619);
and U2982 (N_2982,N_2467,N_2453);
nor U2983 (N_2983,N_2416,N_2559);
nand U2984 (N_2984,N_2794,N_2496);
xor U2985 (N_2985,N_2657,N_2444);
nand U2986 (N_2986,N_2470,N_2587);
nor U2987 (N_2987,N_2634,N_2605);
nor U2988 (N_2988,N_2523,N_2705);
and U2989 (N_2989,N_2637,N_2448);
and U2990 (N_2990,N_2660,N_2430);
and U2991 (N_2991,N_2629,N_2692);
xor U2992 (N_2992,N_2658,N_2454);
or U2993 (N_2993,N_2580,N_2412);
xnor U2994 (N_2994,N_2428,N_2723);
or U2995 (N_2995,N_2593,N_2702);
xnor U2996 (N_2996,N_2581,N_2446);
or U2997 (N_2997,N_2563,N_2744);
xnor U2998 (N_2998,N_2442,N_2632);
nor U2999 (N_2999,N_2733,N_2624);
nand U3000 (N_3000,N_2574,N_2609);
nor U3001 (N_3001,N_2530,N_2432);
nor U3002 (N_3002,N_2492,N_2734);
nand U3003 (N_3003,N_2783,N_2628);
xnor U3004 (N_3004,N_2600,N_2412);
and U3005 (N_3005,N_2731,N_2624);
or U3006 (N_3006,N_2450,N_2556);
nand U3007 (N_3007,N_2495,N_2589);
nor U3008 (N_3008,N_2766,N_2715);
nand U3009 (N_3009,N_2592,N_2738);
or U3010 (N_3010,N_2761,N_2738);
nor U3011 (N_3011,N_2719,N_2694);
nand U3012 (N_3012,N_2477,N_2794);
xor U3013 (N_3013,N_2745,N_2654);
nor U3014 (N_3014,N_2470,N_2769);
nand U3015 (N_3015,N_2790,N_2793);
xor U3016 (N_3016,N_2430,N_2729);
nor U3017 (N_3017,N_2561,N_2725);
nor U3018 (N_3018,N_2447,N_2506);
nor U3019 (N_3019,N_2720,N_2764);
and U3020 (N_3020,N_2599,N_2505);
nor U3021 (N_3021,N_2771,N_2437);
xor U3022 (N_3022,N_2468,N_2782);
xor U3023 (N_3023,N_2774,N_2495);
or U3024 (N_3024,N_2657,N_2490);
and U3025 (N_3025,N_2763,N_2667);
nand U3026 (N_3026,N_2674,N_2581);
nor U3027 (N_3027,N_2558,N_2577);
nand U3028 (N_3028,N_2665,N_2713);
nand U3029 (N_3029,N_2582,N_2570);
xor U3030 (N_3030,N_2669,N_2726);
and U3031 (N_3031,N_2679,N_2525);
or U3032 (N_3032,N_2642,N_2457);
and U3033 (N_3033,N_2563,N_2606);
xnor U3034 (N_3034,N_2765,N_2641);
and U3035 (N_3035,N_2516,N_2746);
or U3036 (N_3036,N_2570,N_2682);
and U3037 (N_3037,N_2596,N_2411);
or U3038 (N_3038,N_2486,N_2438);
nor U3039 (N_3039,N_2432,N_2496);
xnor U3040 (N_3040,N_2786,N_2655);
nor U3041 (N_3041,N_2589,N_2528);
nor U3042 (N_3042,N_2671,N_2412);
and U3043 (N_3043,N_2781,N_2411);
nand U3044 (N_3044,N_2633,N_2607);
nor U3045 (N_3045,N_2439,N_2785);
and U3046 (N_3046,N_2774,N_2706);
nor U3047 (N_3047,N_2466,N_2699);
nand U3048 (N_3048,N_2709,N_2688);
nand U3049 (N_3049,N_2523,N_2428);
xnor U3050 (N_3050,N_2604,N_2785);
nor U3051 (N_3051,N_2456,N_2418);
nor U3052 (N_3052,N_2669,N_2435);
nor U3053 (N_3053,N_2593,N_2665);
nand U3054 (N_3054,N_2531,N_2564);
nand U3055 (N_3055,N_2550,N_2677);
and U3056 (N_3056,N_2477,N_2650);
xor U3057 (N_3057,N_2613,N_2712);
nor U3058 (N_3058,N_2589,N_2688);
xor U3059 (N_3059,N_2618,N_2467);
and U3060 (N_3060,N_2726,N_2616);
and U3061 (N_3061,N_2412,N_2733);
xor U3062 (N_3062,N_2700,N_2652);
and U3063 (N_3063,N_2608,N_2648);
and U3064 (N_3064,N_2725,N_2450);
and U3065 (N_3065,N_2418,N_2455);
xnor U3066 (N_3066,N_2699,N_2520);
nor U3067 (N_3067,N_2487,N_2591);
or U3068 (N_3068,N_2455,N_2663);
or U3069 (N_3069,N_2557,N_2480);
nand U3070 (N_3070,N_2517,N_2769);
or U3071 (N_3071,N_2784,N_2773);
or U3072 (N_3072,N_2575,N_2593);
xor U3073 (N_3073,N_2411,N_2435);
or U3074 (N_3074,N_2559,N_2670);
and U3075 (N_3075,N_2431,N_2730);
or U3076 (N_3076,N_2479,N_2631);
xor U3077 (N_3077,N_2450,N_2588);
xnor U3078 (N_3078,N_2644,N_2767);
and U3079 (N_3079,N_2573,N_2728);
or U3080 (N_3080,N_2514,N_2705);
nand U3081 (N_3081,N_2761,N_2561);
xnor U3082 (N_3082,N_2677,N_2746);
or U3083 (N_3083,N_2782,N_2424);
nor U3084 (N_3084,N_2672,N_2773);
nor U3085 (N_3085,N_2751,N_2444);
or U3086 (N_3086,N_2523,N_2623);
nor U3087 (N_3087,N_2436,N_2495);
and U3088 (N_3088,N_2560,N_2745);
or U3089 (N_3089,N_2768,N_2431);
nand U3090 (N_3090,N_2757,N_2510);
xor U3091 (N_3091,N_2765,N_2681);
or U3092 (N_3092,N_2569,N_2437);
or U3093 (N_3093,N_2494,N_2737);
or U3094 (N_3094,N_2702,N_2465);
or U3095 (N_3095,N_2471,N_2558);
and U3096 (N_3096,N_2636,N_2664);
nor U3097 (N_3097,N_2550,N_2616);
xor U3098 (N_3098,N_2477,N_2521);
or U3099 (N_3099,N_2553,N_2522);
and U3100 (N_3100,N_2757,N_2502);
or U3101 (N_3101,N_2614,N_2441);
nand U3102 (N_3102,N_2567,N_2508);
and U3103 (N_3103,N_2534,N_2459);
or U3104 (N_3104,N_2589,N_2438);
nor U3105 (N_3105,N_2703,N_2695);
or U3106 (N_3106,N_2423,N_2413);
nand U3107 (N_3107,N_2684,N_2740);
xnor U3108 (N_3108,N_2566,N_2588);
or U3109 (N_3109,N_2617,N_2721);
nand U3110 (N_3110,N_2765,N_2563);
xor U3111 (N_3111,N_2663,N_2562);
nor U3112 (N_3112,N_2684,N_2477);
and U3113 (N_3113,N_2703,N_2463);
or U3114 (N_3114,N_2491,N_2432);
and U3115 (N_3115,N_2454,N_2694);
nor U3116 (N_3116,N_2506,N_2574);
and U3117 (N_3117,N_2734,N_2750);
nand U3118 (N_3118,N_2408,N_2572);
nand U3119 (N_3119,N_2538,N_2401);
or U3120 (N_3120,N_2697,N_2526);
xor U3121 (N_3121,N_2669,N_2462);
nor U3122 (N_3122,N_2738,N_2520);
or U3123 (N_3123,N_2678,N_2513);
and U3124 (N_3124,N_2658,N_2499);
or U3125 (N_3125,N_2546,N_2562);
or U3126 (N_3126,N_2443,N_2470);
xor U3127 (N_3127,N_2439,N_2404);
and U3128 (N_3128,N_2582,N_2444);
or U3129 (N_3129,N_2775,N_2679);
xor U3130 (N_3130,N_2763,N_2635);
nor U3131 (N_3131,N_2750,N_2546);
xor U3132 (N_3132,N_2732,N_2502);
and U3133 (N_3133,N_2743,N_2462);
xor U3134 (N_3134,N_2466,N_2767);
or U3135 (N_3135,N_2796,N_2406);
or U3136 (N_3136,N_2490,N_2488);
or U3137 (N_3137,N_2590,N_2731);
xor U3138 (N_3138,N_2615,N_2582);
xnor U3139 (N_3139,N_2793,N_2713);
nor U3140 (N_3140,N_2698,N_2429);
and U3141 (N_3141,N_2635,N_2738);
or U3142 (N_3142,N_2779,N_2759);
nand U3143 (N_3143,N_2766,N_2709);
nor U3144 (N_3144,N_2706,N_2438);
nor U3145 (N_3145,N_2499,N_2475);
xnor U3146 (N_3146,N_2412,N_2744);
or U3147 (N_3147,N_2733,N_2719);
xor U3148 (N_3148,N_2717,N_2758);
nor U3149 (N_3149,N_2734,N_2733);
nand U3150 (N_3150,N_2449,N_2793);
or U3151 (N_3151,N_2715,N_2549);
and U3152 (N_3152,N_2576,N_2612);
nor U3153 (N_3153,N_2722,N_2503);
nor U3154 (N_3154,N_2793,N_2531);
xor U3155 (N_3155,N_2686,N_2712);
and U3156 (N_3156,N_2793,N_2485);
nand U3157 (N_3157,N_2763,N_2704);
or U3158 (N_3158,N_2520,N_2525);
xnor U3159 (N_3159,N_2485,N_2781);
xor U3160 (N_3160,N_2703,N_2476);
and U3161 (N_3161,N_2459,N_2641);
or U3162 (N_3162,N_2652,N_2795);
and U3163 (N_3163,N_2796,N_2413);
nor U3164 (N_3164,N_2439,N_2441);
and U3165 (N_3165,N_2667,N_2546);
or U3166 (N_3166,N_2410,N_2508);
or U3167 (N_3167,N_2782,N_2772);
nand U3168 (N_3168,N_2475,N_2511);
nand U3169 (N_3169,N_2745,N_2484);
nor U3170 (N_3170,N_2409,N_2761);
or U3171 (N_3171,N_2523,N_2493);
nor U3172 (N_3172,N_2711,N_2794);
nor U3173 (N_3173,N_2651,N_2624);
nor U3174 (N_3174,N_2778,N_2505);
or U3175 (N_3175,N_2697,N_2536);
nand U3176 (N_3176,N_2436,N_2769);
nand U3177 (N_3177,N_2603,N_2585);
nor U3178 (N_3178,N_2698,N_2599);
nand U3179 (N_3179,N_2617,N_2737);
and U3180 (N_3180,N_2747,N_2589);
nand U3181 (N_3181,N_2789,N_2723);
xnor U3182 (N_3182,N_2430,N_2531);
or U3183 (N_3183,N_2714,N_2629);
nor U3184 (N_3184,N_2704,N_2507);
or U3185 (N_3185,N_2452,N_2423);
and U3186 (N_3186,N_2660,N_2743);
and U3187 (N_3187,N_2433,N_2565);
nor U3188 (N_3188,N_2797,N_2766);
nor U3189 (N_3189,N_2578,N_2620);
xnor U3190 (N_3190,N_2563,N_2693);
xor U3191 (N_3191,N_2544,N_2536);
and U3192 (N_3192,N_2441,N_2533);
nor U3193 (N_3193,N_2598,N_2766);
or U3194 (N_3194,N_2641,N_2678);
nand U3195 (N_3195,N_2578,N_2508);
nor U3196 (N_3196,N_2497,N_2746);
xnor U3197 (N_3197,N_2639,N_2650);
and U3198 (N_3198,N_2599,N_2442);
and U3199 (N_3199,N_2763,N_2540);
nand U3200 (N_3200,N_2942,N_3081);
xnor U3201 (N_3201,N_2884,N_2814);
or U3202 (N_3202,N_2867,N_3042);
nand U3203 (N_3203,N_2940,N_3052);
or U3204 (N_3204,N_2857,N_2923);
and U3205 (N_3205,N_2980,N_3145);
and U3206 (N_3206,N_2821,N_3022);
and U3207 (N_3207,N_2965,N_3066);
nor U3208 (N_3208,N_3157,N_3027);
or U3209 (N_3209,N_2936,N_3077);
nor U3210 (N_3210,N_3071,N_2977);
xnor U3211 (N_3211,N_3011,N_2892);
nand U3212 (N_3212,N_3174,N_2924);
xnor U3213 (N_3213,N_3087,N_3195);
xnor U3214 (N_3214,N_3045,N_3028);
nor U3215 (N_3215,N_3194,N_3057);
or U3216 (N_3216,N_2916,N_3094);
nand U3217 (N_3217,N_2969,N_2907);
or U3218 (N_3218,N_3024,N_3199);
and U3219 (N_3219,N_2811,N_3059);
nor U3220 (N_3220,N_3013,N_3017);
and U3221 (N_3221,N_2870,N_3175);
nand U3222 (N_3222,N_2982,N_3067);
xor U3223 (N_3223,N_2882,N_2911);
or U3224 (N_3224,N_2993,N_3193);
nand U3225 (N_3225,N_3043,N_3047);
or U3226 (N_3226,N_3086,N_3169);
nand U3227 (N_3227,N_3030,N_2888);
and U3228 (N_3228,N_2932,N_2875);
nand U3229 (N_3229,N_3164,N_3080);
nor U3230 (N_3230,N_3056,N_2910);
nor U3231 (N_3231,N_2938,N_2822);
and U3232 (N_3232,N_3069,N_3050);
and U3233 (N_3233,N_3113,N_3105);
xnor U3234 (N_3234,N_3159,N_2863);
nor U3235 (N_3235,N_2970,N_2948);
nor U3236 (N_3236,N_2803,N_3070);
and U3237 (N_3237,N_3021,N_2869);
or U3238 (N_3238,N_3141,N_3109);
nor U3239 (N_3239,N_3123,N_2902);
and U3240 (N_3240,N_2873,N_3138);
xor U3241 (N_3241,N_2997,N_2960);
nor U3242 (N_3242,N_3114,N_3139);
nand U3243 (N_3243,N_2978,N_3039);
nand U3244 (N_3244,N_3010,N_3106);
nor U3245 (N_3245,N_2836,N_3085);
nand U3246 (N_3246,N_2835,N_3187);
and U3247 (N_3247,N_3020,N_3144);
or U3248 (N_3248,N_3023,N_2878);
nand U3249 (N_3249,N_3177,N_2930);
and U3250 (N_3250,N_3036,N_2889);
nor U3251 (N_3251,N_2823,N_2840);
and U3252 (N_3252,N_3063,N_3001);
nor U3253 (N_3253,N_3183,N_3108);
or U3254 (N_3254,N_3018,N_3092);
and U3255 (N_3255,N_2956,N_2856);
nand U3256 (N_3256,N_3046,N_3096);
or U3257 (N_3257,N_3014,N_3127);
or U3258 (N_3258,N_3053,N_3125);
nor U3259 (N_3259,N_2824,N_3034);
nand U3260 (N_3260,N_3076,N_3156);
or U3261 (N_3261,N_3009,N_2800);
or U3262 (N_3262,N_2895,N_3111);
nand U3263 (N_3263,N_3176,N_2818);
xor U3264 (N_3264,N_2917,N_2904);
nor U3265 (N_3265,N_2944,N_3132);
nand U3266 (N_3266,N_3115,N_3197);
nand U3267 (N_3267,N_2999,N_2862);
nor U3268 (N_3268,N_3015,N_2816);
and U3269 (N_3269,N_2843,N_3116);
or U3270 (N_3270,N_3110,N_2830);
xor U3271 (N_3271,N_3058,N_2897);
nor U3272 (N_3272,N_3182,N_3078);
nand U3273 (N_3273,N_3090,N_3065);
nor U3274 (N_3274,N_2927,N_2951);
xnor U3275 (N_3275,N_2920,N_3137);
nor U3276 (N_3276,N_3165,N_3075);
nand U3277 (N_3277,N_3186,N_3135);
or U3278 (N_3278,N_2988,N_3190);
xor U3279 (N_3279,N_2914,N_3072);
or U3280 (N_3280,N_3130,N_3032);
or U3281 (N_3281,N_3098,N_2883);
nor U3282 (N_3282,N_3008,N_2898);
or U3283 (N_3283,N_2935,N_3041);
nor U3284 (N_3284,N_3134,N_3097);
and U3285 (N_3285,N_3196,N_2954);
or U3286 (N_3286,N_2894,N_2903);
nand U3287 (N_3287,N_2880,N_3153);
xor U3288 (N_3288,N_2807,N_2842);
nand U3289 (N_3289,N_2934,N_3044);
xor U3290 (N_3290,N_3149,N_3026);
xnor U3291 (N_3291,N_2900,N_2893);
and U3292 (N_3292,N_2953,N_3198);
or U3293 (N_3293,N_3136,N_2804);
and U3294 (N_3294,N_2957,N_2958);
nor U3295 (N_3295,N_3162,N_3006);
xnor U3296 (N_3296,N_3124,N_2806);
nand U3297 (N_3297,N_2881,N_3131);
xor U3298 (N_3298,N_3061,N_2986);
and U3299 (N_3299,N_2974,N_2879);
nand U3300 (N_3300,N_3192,N_2901);
xnor U3301 (N_3301,N_2855,N_3184);
and U3302 (N_3302,N_3181,N_2861);
nand U3303 (N_3303,N_3016,N_2913);
xor U3304 (N_3304,N_2809,N_2967);
nand U3305 (N_3305,N_2860,N_3143);
nor U3306 (N_3306,N_3148,N_2994);
nand U3307 (N_3307,N_3003,N_2899);
or U3308 (N_3308,N_3005,N_2896);
nor U3309 (N_3309,N_2962,N_3064);
or U3310 (N_3310,N_3121,N_3188);
and U3311 (N_3311,N_2908,N_3099);
or U3312 (N_3312,N_3152,N_2819);
nor U3313 (N_3313,N_2912,N_2952);
nand U3314 (N_3314,N_3191,N_2817);
or U3315 (N_3315,N_3160,N_2925);
and U3316 (N_3316,N_2955,N_2802);
or U3317 (N_3317,N_2847,N_2837);
and U3318 (N_3318,N_2996,N_2964);
or U3319 (N_3319,N_2992,N_2987);
and U3320 (N_3320,N_2961,N_2947);
nor U3321 (N_3321,N_3107,N_2998);
xnor U3322 (N_3322,N_2846,N_2808);
nand U3323 (N_3323,N_3048,N_2946);
xor U3324 (N_3324,N_2915,N_3012);
nand U3325 (N_3325,N_2849,N_3189);
or U3326 (N_3326,N_3073,N_2963);
nor U3327 (N_3327,N_3089,N_3102);
xor U3328 (N_3328,N_2890,N_2810);
xnor U3329 (N_3329,N_2877,N_2959);
nor U3330 (N_3330,N_2852,N_2825);
nor U3331 (N_3331,N_2865,N_2926);
nor U3332 (N_3332,N_3068,N_3185);
and U3333 (N_3333,N_2829,N_2838);
and U3334 (N_3334,N_3093,N_2909);
or U3335 (N_3335,N_2981,N_2989);
nor U3336 (N_3336,N_3122,N_2858);
xor U3337 (N_3337,N_3007,N_2905);
or U3338 (N_3338,N_3154,N_3147);
xnor U3339 (N_3339,N_2941,N_3155);
or U3340 (N_3340,N_3095,N_3163);
or U3341 (N_3341,N_3171,N_2866);
and U3342 (N_3342,N_3120,N_3035);
xnor U3343 (N_3343,N_2968,N_3126);
or U3344 (N_3344,N_2885,N_2971);
nor U3345 (N_3345,N_3180,N_2859);
xnor U3346 (N_3346,N_3170,N_2972);
and U3347 (N_3347,N_3151,N_2801);
nand U3348 (N_3348,N_2945,N_2995);
nor U3349 (N_3349,N_2828,N_3040);
nand U3350 (N_3350,N_3082,N_2906);
nand U3351 (N_3351,N_3084,N_3037);
nor U3352 (N_3352,N_3103,N_3055);
nor U3353 (N_3353,N_3038,N_3173);
nor U3354 (N_3354,N_3142,N_3150);
nand U3355 (N_3355,N_3117,N_2939);
nor U3356 (N_3356,N_2990,N_2891);
or U3357 (N_3357,N_3049,N_3158);
or U3358 (N_3358,N_3079,N_2841);
nand U3359 (N_3359,N_2854,N_3074);
and U3360 (N_3360,N_2950,N_2844);
nor U3361 (N_3361,N_2929,N_3112);
nor U3362 (N_3362,N_2918,N_3168);
nand U3363 (N_3363,N_2876,N_2834);
nand U3364 (N_3364,N_2919,N_2983);
or U3365 (N_3365,N_2886,N_3029);
nor U3366 (N_3366,N_2868,N_3031);
xnor U3367 (N_3367,N_3100,N_3119);
nand U3368 (N_3368,N_3128,N_2984);
and U3369 (N_3369,N_3060,N_2813);
xor U3370 (N_3370,N_2872,N_2931);
xnor U3371 (N_3371,N_3088,N_2943);
or U3372 (N_3372,N_2985,N_3025);
or U3373 (N_3373,N_2973,N_2815);
nand U3374 (N_3374,N_2820,N_2812);
nor U3375 (N_3375,N_2949,N_2831);
xnor U3376 (N_3376,N_3172,N_2871);
nor U3377 (N_3377,N_3178,N_2933);
and U3378 (N_3378,N_3019,N_2850);
nor U3379 (N_3379,N_3062,N_3166);
nand U3380 (N_3380,N_3161,N_3054);
or U3381 (N_3381,N_3002,N_2887);
or U3382 (N_3382,N_3000,N_3133);
nor U3383 (N_3383,N_3033,N_2979);
nand U3384 (N_3384,N_2832,N_2975);
nor U3385 (N_3385,N_2921,N_2848);
or U3386 (N_3386,N_2874,N_3140);
nor U3387 (N_3387,N_3004,N_2928);
or U3388 (N_3388,N_3104,N_3091);
or U3389 (N_3389,N_2827,N_2826);
nand U3390 (N_3390,N_3146,N_3083);
nor U3391 (N_3391,N_2864,N_3179);
and U3392 (N_3392,N_2851,N_2991);
nand U3393 (N_3393,N_2966,N_2805);
nor U3394 (N_3394,N_3129,N_3101);
xnor U3395 (N_3395,N_3051,N_2976);
or U3396 (N_3396,N_2853,N_3118);
or U3397 (N_3397,N_2922,N_2839);
nand U3398 (N_3398,N_2845,N_2937);
and U3399 (N_3399,N_2833,N_3167);
nor U3400 (N_3400,N_3159,N_3021);
nor U3401 (N_3401,N_3014,N_2999);
nor U3402 (N_3402,N_2808,N_3015);
and U3403 (N_3403,N_2806,N_2944);
nand U3404 (N_3404,N_2902,N_2965);
nor U3405 (N_3405,N_2932,N_3076);
or U3406 (N_3406,N_3097,N_2881);
nand U3407 (N_3407,N_2872,N_2954);
and U3408 (N_3408,N_2819,N_3072);
xor U3409 (N_3409,N_2801,N_2951);
or U3410 (N_3410,N_3179,N_3051);
nor U3411 (N_3411,N_3055,N_2875);
xnor U3412 (N_3412,N_3145,N_3133);
xor U3413 (N_3413,N_3156,N_3132);
xnor U3414 (N_3414,N_3105,N_3161);
or U3415 (N_3415,N_3080,N_3174);
nand U3416 (N_3416,N_2803,N_2907);
nor U3417 (N_3417,N_3144,N_3101);
and U3418 (N_3418,N_3016,N_2899);
nor U3419 (N_3419,N_2877,N_3074);
nand U3420 (N_3420,N_2965,N_2803);
and U3421 (N_3421,N_2980,N_3110);
xor U3422 (N_3422,N_2868,N_2921);
xnor U3423 (N_3423,N_3050,N_2983);
nand U3424 (N_3424,N_2806,N_3052);
nand U3425 (N_3425,N_3071,N_2823);
and U3426 (N_3426,N_2885,N_3168);
and U3427 (N_3427,N_2853,N_3178);
nor U3428 (N_3428,N_2912,N_2823);
or U3429 (N_3429,N_3148,N_3019);
xor U3430 (N_3430,N_3175,N_3050);
nor U3431 (N_3431,N_3150,N_3066);
nor U3432 (N_3432,N_3006,N_2882);
nand U3433 (N_3433,N_3148,N_3184);
xnor U3434 (N_3434,N_3145,N_3158);
or U3435 (N_3435,N_3064,N_3049);
and U3436 (N_3436,N_3084,N_2985);
nor U3437 (N_3437,N_2999,N_3051);
or U3438 (N_3438,N_2924,N_2936);
and U3439 (N_3439,N_2940,N_2922);
nand U3440 (N_3440,N_3120,N_3169);
nand U3441 (N_3441,N_2845,N_2984);
xnor U3442 (N_3442,N_2996,N_3009);
nor U3443 (N_3443,N_2876,N_2950);
xnor U3444 (N_3444,N_3000,N_3059);
and U3445 (N_3445,N_2947,N_2914);
or U3446 (N_3446,N_2887,N_3052);
nand U3447 (N_3447,N_3029,N_3065);
nor U3448 (N_3448,N_3140,N_2833);
or U3449 (N_3449,N_2830,N_3020);
or U3450 (N_3450,N_3054,N_3074);
and U3451 (N_3451,N_2970,N_2810);
xnor U3452 (N_3452,N_2836,N_2967);
nor U3453 (N_3453,N_2876,N_2869);
nand U3454 (N_3454,N_2953,N_2840);
and U3455 (N_3455,N_3116,N_3189);
and U3456 (N_3456,N_3192,N_2935);
and U3457 (N_3457,N_2831,N_2993);
and U3458 (N_3458,N_3084,N_2943);
and U3459 (N_3459,N_2962,N_2952);
xnor U3460 (N_3460,N_2863,N_3088);
and U3461 (N_3461,N_2865,N_3018);
or U3462 (N_3462,N_2993,N_3148);
nor U3463 (N_3463,N_3120,N_2927);
nand U3464 (N_3464,N_2815,N_3096);
and U3465 (N_3465,N_2982,N_2811);
nand U3466 (N_3466,N_3167,N_3083);
or U3467 (N_3467,N_3091,N_3071);
nor U3468 (N_3468,N_3054,N_3105);
or U3469 (N_3469,N_2976,N_2956);
and U3470 (N_3470,N_2929,N_2892);
nor U3471 (N_3471,N_2999,N_2814);
nor U3472 (N_3472,N_3084,N_3113);
nand U3473 (N_3473,N_2824,N_2933);
and U3474 (N_3474,N_3121,N_3019);
or U3475 (N_3475,N_2883,N_3153);
nand U3476 (N_3476,N_2952,N_2876);
xnor U3477 (N_3477,N_3136,N_3127);
nor U3478 (N_3478,N_3010,N_2866);
or U3479 (N_3479,N_3127,N_3075);
and U3480 (N_3480,N_3196,N_2930);
xnor U3481 (N_3481,N_3144,N_3198);
nor U3482 (N_3482,N_2802,N_3035);
xor U3483 (N_3483,N_3081,N_3123);
nor U3484 (N_3484,N_3088,N_2868);
nand U3485 (N_3485,N_2938,N_2958);
nand U3486 (N_3486,N_3029,N_3135);
or U3487 (N_3487,N_2963,N_2808);
xor U3488 (N_3488,N_3040,N_2885);
nor U3489 (N_3489,N_2847,N_2982);
nand U3490 (N_3490,N_3192,N_3027);
xnor U3491 (N_3491,N_2925,N_3134);
nand U3492 (N_3492,N_3077,N_3083);
nor U3493 (N_3493,N_2992,N_2867);
and U3494 (N_3494,N_2837,N_3000);
nor U3495 (N_3495,N_2928,N_2858);
nand U3496 (N_3496,N_3038,N_2867);
nor U3497 (N_3497,N_3066,N_3132);
and U3498 (N_3498,N_3006,N_2926);
or U3499 (N_3499,N_3074,N_2906);
xnor U3500 (N_3500,N_3008,N_2894);
xnor U3501 (N_3501,N_3042,N_2873);
nor U3502 (N_3502,N_3158,N_3150);
xor U3503 (N_3503,N_3156,N_3073);
xor U3504 (N_3504,N_3094,N_2928);
xor U3505 (N_3505,N_2934,N_3193);
xnor U3506 (N_3506,N_2813,N_2939);
nor U3507 (N_3507,N_2892,N_2941);
xor U3508 (N_3508,N_3051,N_3030);
and U3509 (N_3509,N_2854,N_3186);
xor U3510 (N_3510,N_2988,N_2806);
nand U3511 (N_3511,N_3172,N_2843);
nand U3512 (N_3512,N_2904,N_3036);
or U3513 (N_3513,N_2809,N_2957);
xnor U3514 (N_3514,N_2807,N_2831);
and U3515 (N_3515,N_2977,N_3102);
or U3516 (N_3516,N_3119,N_2873);
and U3517 (N_3517,N_2937,N_2827);
and U3518 (N_3518,N_3122,N_2826);
or U3519 (N_3519,N_3189,N_2951);
and U3520 (N_3520,N_3046,N_2808);
nand U3521 (N_3521,N_2941,N_3171);
xor U3522 (N_3522,N_3062,N_2911);
nand U3523 (N_3523,N_3165,N_2884);
xnor U3524 (N_3524,N_3111,N_2847);
or U3525 (N_3525,N_2897,N_3090);
or U3526 (N_3526,N_2867,N_3009);
or U3527 (N_3527,N_2904,N_3015);
nor U3528 (N_3528,N_2879,N_2821);
or U3529 (N_3529,N_3065,N_2815);
xor U3530 (N_3530,N_3030,N_2882);
and U3531 (N_3531,N_2864,N_2915);
nand U3532 (N_3532,N_2929,N_2994);
and U3533 (N_3533,N_3135,N_3043);
nand U3534 (N_3534,N_2891,N_3144);
xnor U3535 (N_3535,N_3008,N_3196);
nor U3536 (N_3536,N_2854,N_2915);
and U3537 (N_3537,N_2861,N_3182);
nand U3538 (N_3538,N_3040,N_3124);
xnor U3539 (N_3539,N_2898,N_3082);
nand U3540 (N_3540,N_3096,N_3140);
or U3541 (N_3541,N_2996,N_2812);
and U3542 (N_3542,N_3130,N_2907);
xor U3543 (N_3543,N_3077,N_2972);
and U3544 (N_3544,N_3026,N_2943);
nor U3545 (N_3545,N_3186,N_3121);
nor U3546 (N_3546,N_3061,N_2856);
nor U3547 (N_3547,N_3006,N_3030);
xnor U3548 (N_3548,N_3115,N_2894);
and U3549 (N_3549,N_3187,N_2889);
and U3550 (N_3550,N_2901,N_2989);
and U3551 (N_3551,N_2824,N_2919);
xor U3552 (N_3552,N_3158,N_2928);
or U3553 (N_3553,N_3019,N_3184);
nand U3554 (N_3554,N_3032,N_3039);
xnor U3555 (N_3555,N_2889,N_3180);
nor U3556 (N_3556,N_3105,N_2968);
nor U3557 (N_3557,N_3169,N_2819);
and U3558 (N_3558,N_2835,N_3144);
and U3559 (N_3559,N_3138,N_3155);
nor U3560 (N_3560,N_2916,N_3064);
or U3561 (N_3561,N_3075,N_2897);
and U3562 (N_3562,N_3153,N_3193);
xor U3563 (N_3563,N_2867,N_3130);
nand U3564 (N_3564,N_2867,N_3167);
nor U3565 (N_3565,N_3042,N_3056);
xnor U3566 (N_3566,N_3194,N_3091);
and U3567 (N_3567,N_2974,N_3117);
nor U3568 (N_3568,N_3040,N_3071);
and U3569 (N_3569,N_2945,N_2918);
nor U3570 (N_3570,N_3024,N_3146);
and U3571 (N_3571,N_2912,N_2856);
xnor U3572 (N_3572,N_2908,N_2948);
nand U3573 (N_3573,N_2923,N_2975);
and U3574 (N_3574,N_2992,N_3161);
nand U3575 (N_3575,N_2880,N_3086);
or U3576 (N_3576,N_3094,N_2911);
or U3577 (N_3577,N_3013,N_2925);
nor U3578 (N_3578,N_2900,N_3193);
nand U3579 (N_3579,N_3051,N_3066);
and U3580 (N_3580,N_3077,N_2976);
and U3581 (N_3581,N_2892,N_2938);
or U3582 (N_3582,N_3031,N_2811);
and U3583 (N_3583,N_3106,N_3167);
nand U3584 (N_3584,N_2807,N_3073);
nand U3585 (N_3585,N_2864,N_3047);
or U3586 (N_3586,N_3109,N_2938);
xor U3587 (N_3587,N_2982,N_3196);
or U3588 (N_3588,N_3108,N_3017);
nor U3589 (N_3589,N_2801,N_2973);
nor U3590 (N_3590,N_2994,N_3184);
nor U3591 (N_3591,N_2800,N_3187);
or U3592 (N_3592,N_3018,N_2950);
nor U3593 (N_3593,N_2811,N_2979);
nor U3594 (N_3594,N_2800,N_3001);
xnor U3595 (N_3595,N_3159,N_2941);
or U3596 (N_3596,N_2918,N_2922);
xnor U3597 (N_3597,N_2930,N_3097);
nand U3598 (N_3598,N_2849,N_3040);
nor U3599 (N_3599,N_3179,N_3004);
and U3600 (N_3600,N_3397,N_3336);
xnor U3601 (N_3601,N_3437,N_3299);
nor U3602 (N_3602,N_3459,N_3369);
nor U3603 (N_3603,N_3452,N_3288);
nand U3604 (N_3604,N_3577,N_3365);
xnor U3605 (N_3605,N_3387,N_3416);
nand U3606 (N_3606,N_3325,N_3464);
xnor U3607 (N_3607,N_3465,N_3575);
and U3608 (N_3608,N_3213,N_3320);
xnor U3609 (N_3609,N_3393,N_3547);
and U3610 (N_3610,N_3311,N_3259);
and U3611 (N_3611,N_3264,N_3447);
and U3612 (N_3612,N_3216,N_3305);
xnor U3613 (N_3613,N_3364,N_3413);
or U3614 (N_3614,N_3515,N_3513);
or U3615 (N_3615,N_3519,N_3543);
xor U3616 (N_3616,N_3417,N_3301);
xor U3617 (N_3617,N_3540,N_3472);
or U3618 (N_3618,N_3240,N_3330);
and U3619 (N_3619,N_3383,N_3319);
xor U3620 (N_3620,N_3255,N_3436);
xor U3621 (N_3621,N_3410,N_3275);
nor U3622 (N_3622,N_3594,N_3475);
and U3623 (N_3623,N_3399,N_3585);
or U3624 (N_3624,N_3498,N_3244);
nor U3625 (N_3625,N_3202,N_3396);
nor U3626 (N_3626,N_3376,N_3507);
xor U3627 (N_3627,N_3555,N_3420);
and U3628 (N_3628,N_3212,N_3407);
nor U3629 (N_3629,N_3208,N_3433);
nand U3630 (N_3630,N_3250,N_3296);
nand U3631 (N_3631,N_3286,N_3551);
and U3632 (N_3632,N_3354,N_3500);
or U3633 (N_3633,N_3386,N_3548);
xor U3634 (N_3634,N_3228,N_3532);
nor U3635 (N_3635,N_3215,N_3586);
nor U3636 (N_3636,N_3245,N_3221);
and U3637 (N_3637,N_3293,N_3317);
nand U3638 (N_3638,N_3374,N_3297);
and U3639 (N_3639,N_3344,N_3243);
xor U3640 (N_3640,N_3552,N_3388);
and U3641 (N_3641,N_3321,N_3484);
nor U3642 (N_3642,N_3556,N_3518);
and U3643 (N_3643,N_3308,N_3405);
and U3644 (N_3644,N_3347,N_3313);
and U3645 (N_3645,N_3384,N_3576);
xnor U3646 (N_3646,N_3581,N_3342);
nand U3647 (N_3647,N_3415,N_3520);
and U3648 (N_3648,N_3303,N_3289);
and U3649 (N_3649,N_3522,N_3403);
or U3650 (N_3650,N_3377,N_3566);
xnor U3651 (N_3651,N_3430,N_3345);
or U3652 (N_3652,N_3537,N_3200);
xnor U3653 (N_3653,N_3477,N_3404);
and U3654 (N_3654,N_3220,N_3483);
nand U3655 (N_3655,N_3453,N_3267);
nand U3656 (N_3656,N_3573,N_3579);
or U3657 (N_3657,N_3569,N_3442);
and U3658 (N_3658,N_3290,N_3458);
or U3659 (N_3659,N_3489,N_3315);
nand U3660 (N_3660,N_3593,N_3528);
and U3661 (N_3661,N_3428,N_3438);
nor U3662 (N_3662,N_3266,N_3571);
xor U3663 (N_3663,N_3359,N_3389);
nand U3664 (N_3664,N_3524,N_3280);
nand U3665 (N_3665,N_3274,N_3260);
or U3666 (N_3666,N_3578,N_3252);
xor U3667 (N_3667,N_3281,N_3511);
or U3668 (N_3668,N_3271,N_3310);
xnor U3669 (N_3669,N_3331,N_3599);
xnor U3670 (N_3670,N_3362,N_3368);
and U3671 (N_3671,N_3559,N_3201);
and U3672 (N_3672,N_3482,N_3486);
nand U3673 (N_3673,N_3360,N_3446);
nor U3674 (N_3674,N_3381,N_3278);
and U3675 (N_3675,N_3338,N_3233);
or U3676 (N_3676,N_3277,N_3309);
nand U3677 (N_3677,N_3440,N_3523);
nor U3678 (N_3678,N_3235,N_3598);
and U3679 (N_3679,N_3203,N_3249);
xnor U3680 (N_3680,N_3525,N_3570);
nand U3681 (N_3681,N_3490,N_3287);
nand U3682 (N_3682,N_3401,N_3595);
or U3683 (N_3683,N_3535,N_3558);
nand U3684 (N_3684,N_3379,N_3390);
or U3685 (N_3685,N_3485,N_3580);
or U3686 (N_3686,N_3361,N_3402);
nand U3687 (N_3687,N_3514,N_3496);
and U3688 (N_3688,N_3352,N_3391);
and U3689 (N_3689,N_3234,N_3488);
nor U3690 (N_3690,N_3246,N_3307);
or U3691 (N_3691,N_3589,N_3517);
xnor U3692 (N_3692,N_3409,N_3539);
nand U3693 (N_3693,N_3291,N_3545);
and U3694 (N_3694,N_3263,N_3568);
nand U3695 (N_3695,N_3516,N_3242);
and U3696 (N_3696,N_3257,N_3341);
and U3697 (N_3697,N_3348,N_3258);
nor U3698 (N_3698,N_3300,N_3451);
xnor U3699 (N_3699,N_3499,N_3455);
or U3700 (N_3700,N_3592,N_3423);
nand U3701 (N_3701,N_3424,N_3512);
nor U3702 (N_3702,N_3529,N_3225);
and U3703 (N_3703,N_3449,N_3471);
nor U3704 (N_3704,N_3346,N_3501);
nor U3705 (N_3705,N_3429,N_3314);
xnor U3706 (N_3706,N_3487,N_3406);
nand U3707 (N_3707,N_3236,N_3253);
nand U3708 (N_3708,N_3448,N_3334);
xnor U3709 (N_3709,N_3494,N_3256);
or U3710 (N_3710,N_3375,N_3412);
xnor U3711 (N_3711,N_3443,N_3357);
or U3712 (N_3712,N_3505,N_3370);
or U3713 (N_3713,N_3553,N_3468);
and U3714 (N_3714,N_3339,N_3340);
and U3715 (N_3715,N_3533,N_3355);
and U3716 (N_3716,N_3343,N_3439);
nand U3717 (N_3717,N_3597,N_3276);
and U3718 (N_3718,N_3363,N_3426);
or U3719 (N_3719,N_3434,N_3408);
xnor U3720 (N_3720,N_3469,N_3265);
or U3721 (N_3721,N_3380,N_3549);
or U3722 (N_3722,N_3304,N_3544);
nor U3723 (N_3723,N_3435,N_3527);
nand U3724 (N_3724,N_3400,N_3230);
xor U3725 (N_3725,N_3226,N_3506);
xor U3726 (N_3726,N_3481,N_3584);
nand U3727 (N_3727,N_3470,N_3295);
nand U3728 (N_3728,N_3510,N_3454);
or U3729 (N_3729,N_3385,N_3419);
nand U3730 (N_3730,N_3480,N_3398);
and U3731 (N_3731,N_3542,N_3335);
or U3732 (N_3732,N_3350,N_3560);
and U3733 (N_3733,N_3241,N_3508);
nor U3734 (N_3734,N_3421,N_3588);
and U3735 (N_3735,N_3431,N_3209);
and U3736 (N_3736,N_3332,N_3318);
nor U3737 (N_3737,N_3229,N_3450);
or U3738 (N_3738,N_3298,N_3227);
and U3739 (N_3739,N_3272,N_3427);
nand U3740 (N_3740,N_3563,N_3232);
or U3741 (N_3741,N_3463,N_3503);
or U3742 (N_3742,N_3461,N_3382);
or U3743 (N_3743,N_3546,N_3590);
and U3744 (N_3744,N_3541,N_3282);
or U3745 (N_3745,N_3204,N_3474);
or U3746 (N_3746,N_3239,N_3283);
xnor U3747 (N_3747,N_3284,N_3306);
and U3748 (N_3748,N_3326,N_3333);
or U3749 (N_3749,N_3587,N_3531);
and U3750 (N_3750,N_3268,N_3536);
nand U3751 (N_3751,N_3222,N_3279);
nor U3752 (N_3752,N_3378,N_3596);
xor U3753 (N_3753,N_3583,N_3425);
or U3754 (N_3754,N_3353,N_3254);
nor U3755 (N_3755,N_3358,N_3247);
nand U3756 (N_3756,N_3562,N_3432);
or U3757 (N_3757,N_3491,N_3324);
nor U3758 (N_3758,N_3273,N_3493);
nand U3759 (N_3759,N_3561,N_3509);
nand U3760 (N_3760,N_3237,N_3591);
or U3761 (N_3761,N_3476,N_3557);
and U3762 (N_3762,N_3564,N_3554);
nand U3763 (N_3763,N_3251,N_3316);
xor U3764 (N_3764,N_3466,N_3418);
nand U3765 (N_3765,N_3462,N_3478);
nor U3766 (N_3766,N_3460,N_3223);
nor U3767 (N_3767,N_3224,N_3582);
xnor U3768 (N_3768,N_3312,N_3521);
nor U3769 (N_3769,N_3322,N_3392);
nand U3770 (N_3770,N_3444,N_3349);
xnor U3771 (N_3771,N_3248,N_3269);
and U3772 (N_3772,N_3411,N_3367);
xnor U3773 (N_3773,N_3572,N_3565);
xnor U3774 (N_3774,N_3270,N_3302);
xnor U3775 (N_3775,N_3497,N_3337);
nand U3776 (N_3776,N_3479,N_3567);
and U3777 (N_3777,N_3526,N_3414);
and U3778 (N_3778,N_3323,N_3441);
and U3779 (N_3779,N_3218,N_3504);
nand U3780 (N_3780,N_3502,N_3214);
nand U3781 (N_3781,N_3329,N_3445);
xnor U3782 (N_3782,N_3456,N_3356);
or U3783 (N_3783,N_3473,N_3327);
and U3784 (N_3784,N_3534,N_3238);
xor U3785 (N_3785,N_3292,N_3467);
xnor U3786 (N_3786,N_3394,N_3371);
or U3787 (N_3787,N_3207,N_3219);
and U3788 (N_3788,N_3262,N_3285);
nand U3789 (N_3789,N_3206,N_3495);
and U3790 (N_3790,N_3328,N_3550);
and U3791 (N_3791,N_3205,N_3574);
and U3792 (N_3792,N_3457,N_3422);
nor U3793 (N_3793,N_3492,N_3294);
nor U3794 (N_3794,N_3217,N_3538);
and U3795 (N_3795,N_3372,N_3373);
or U3796 (N_3796,N_3261,N_3231);
nor U3797 (N_3797,N_3210,N_3395);
and U3798 (N_3798,N_3211,N_3366);
nand U3799 (N_3799,N_3530,N_3351);
and U3800 (N_3800,N_3532,N_3472);
nand U3801 (N_3801,N_3203,N_3390);
xor U3802 (N_3802,N_3327,N_3446);
xnor U3803 (N_3803,N_3217,N_3238);
nor U3804 (N_3804,N_3512,N_3213);
nor U3805 (N_3805,N_3568,N_3385);
nand U3806 (N_3806,N_3576,N_3400);
xnor U3807 (N_3807,N_3233,N_3255);
xnor U3808 (N_3808,N_3487,N_3322);
and U3809 (N_3809,N_3598,N_3203);
nor U3810 (N_3810,N_3475,N_3598);
or U3811 (N_3811,N_3349,N_3490);
nand U3812 (N_3812,N_3376,N_3260);
and U3813 (N_3813,N_3463,N_3587);
nor U3814 (N_3814,N_3254,N_3330);
xnor U3815 (N_3815,N_3317,N_3330);
xnor U3816 (N_3816,N_3384,N_3457);
nand U3817 (N_3817,N_3300,N_3365);
xnor U3818 (N_3818,N_3294,N_3367);
or U3819 (N_3819,N_3219,N_3221);
nor U3820 (N_3820,N_3539,N_3435);
xor U3821 (N_3821,N_3227,N_3592);
nand U3822 (N_3822,N_3432,N_3338);
and U3823 (N_3823,N_3305,N_3319);
and U3824 (N_3824,N_3415,N_3229);
or U3825 (N_3825,N_3406,N_3204);
and U3826 (N_3826,N_3327,N_3364);
or U3827 (N_3827,N_3252,N_3276);
or U3828 (N_3828,N_3557,N_3589);
xnor U3829 (N_3829,N_3597,N_3539);
or U3830 (N_3830,N_3284,N_3428);
xnor U3831 (N_3831,N_3500,N_3320);
and U3832 (N_3832,N_3368,N_3218);
or U3833 (N_3833,N_3568,N_3411);
or U3834 (N_3834,N_3390,N_3249);
nand U3835 (N_3835,N_3436,N_3261);
nand U3836 (N_3836,N_3369,N_3411);
nand U3837 (N_3837,N_3473,N_3341);
nor U3838 (N_3838,N_3590,N_3263);
nor U3839 (N_3839,N_3583,N_3238);
or U3840 (N_3840,N_3208,N_3542);
nor U3841 (N_3841,N_3494,N_3385);
and U3842 (N_3842,N_3577,N_3255);
or U3843 (N_3843,N_3255,N_3417);
nor U3844 (N_3844,N_3378,N_3215);
nor U3845 (N_3845,N_3506,N_3316);
nand U3846 (N_3846,N_3584,N_3597);
xor U3847 (N_3847,N_3552,N_3515);
or U3848 (N_3848,N_3581,N_3533);
xor U3849 (N_3849,N_3519,N_3394);
xnor U3850 (N_3850,N_3556,N_3489);
nor U3851 (N_3851,N_3297,N_3535);
and U3852 (N_3852,N_3290,N_3494);
xnor U3853 (N_3853,N_3488,N_3244);
and U3854 (N_3854,N_3285,N_3245);
nor U3855 (N_3855,N_3350,N_3282);
or U3856 (N_3856,N_3560,N_3374);
xnor U3857 (N_3857,N_3421,N_3526);
or U3858 (N_3858,N_3209,N_3563);
xor U3859 (N_3859,N_3480,N_3494);
and U3860 (N_3860,N_3201,N_3323);
xor U3861 (N_3861,N_3435,N_3259);
xor U3862 (N_3862,N_3360,N_3491);
nor U3863 (N_3863,N_3519,N_3475);
nand U3864 (N_3864,N_3367,N_3562);
nor U3865 (N_3865,N_3266,N_3233);
nand U3866 (N_3866,N_3309,N_3215);
nor U3867 (N_3867,N_3364,N_3507);
and U3868 (N_3868,N_3593,N_3446);
xor U3869 (N_3869,N_3353,N_3208);
nor U3870 (N_3870,N_3535,N_3318);
nand U3871 (N_3871,N_3510,N_3290);
xor U3872 (N_3872,N_3208,N_3543);
and U3873 (N_3873,N_3352,N_3593);
or U3874 (N_3874,N_3394,N_3365);
nand U3875 (N_3875,N_3353,N_3379);
xnor U3876 (N_3876,N_3380,N_3452);
and U3877 (N_3877,N_3298,N_3218);
nor U3878 (N_3878,N_3248,N_3231);
xnor U3879 (N_3879,N_3274,N_3226);
and U3880 (N_3880,N_3433,N_3396);
or U3881 (N_3881,N_3569,N_3559);
and U3882 (N_3882,N_3403,N_3222);
nor U3883 (N_3883,N_3433,N_3543);
or U3884 (N_3884,N_3568,N_3426);
nand U3885 (N_3885,N_3473,N_3579);
or U3886 (N_3886,N_3253,N_3531);
xor U3887 (N_3887,N_3393,N_3317);
xnor U3888 (N_3888,N_3522,N_3348);
and U3889 (N_3889,N_3429,N_3366);
and U3890 (N_3890,N_3426,N_3536);
nand U3891 (N_3891,N_3530,N_3489);
nor U3892 (N_3892,N_3225,N_3324);
and U3893 (N_3893,N_3371,N_3575);
nand U3894 (N_3894,N_3270,N_3532);
nand U3895 (N_3895,N_3439,N_3323);
xnor U3896 (N_3896,N_3221,N_3380);
xor U3897 (N_3897,N_3498,N_3486);
nand U3898 (N_3898,N_3502,N_3542);
xnor U3899 (N_3899,N_3253,N_3289);
nand U3900 (N_3900,N_3404,N_3425);
nor U3901 (N_3901,N_3229,N_3459);
and U3902 (N_3902,N_3556,N_3483);
nor U3903 (N_3903,N_3568,N_3214);
nor U3904 (N_3904,N_3242,N_3485);
or U3905 (N_3905,N_3265,N_3275);
nand U3906 (N_3906,N_3240,N_3568);
and U3907 (N_3907,N_3435,N_3578);
and U3908 (N_3908,N_3460,N_3475);
nor U3909 (N_3909,N_3327,N_3304);
and U3910 (N_3910,N_3515,N_3204);
or U3911 (N_3911,N_3562,N_3224);
xor U3912 (N_3912,N_3289,N_3209);
and U3913 (N_3913,N_3581,N_3421);
and U3914 (N_3914,N_3544,N_3479);
or U3915 (N_3915,N_3350,N_3302);
nand U3916 (N_3916,N_3279,N_3537);
xor U3917 (N_3917,N_3321,N_3514);
and U3918 (N_3918,N_3455,N_3390);
and U3919 (N_3919,N_3371,N_3201);
or U3920 (N_3920,N_3307,N_3212);
xor U3921 (N_3921,N_3528,N_3299);
and U3922 (N_3922,N_3252,N_3386);
xor U3923 (N_3923,N_3340,N_3482);
nor U3924 (N_3924,N_3300,N_3498);
or U3925 (N_3925,N_3471,N_3543);
or U3926 (N_3926,N_3584,N_3503);
and U3927 (N_3927,N_3312,N_3490);
xnor U3928 (N_3928,N_3287,N_3473);
xor U3929 (N_3929,N_3356,N_3260);
xnor U3930 (N_3930,N_3480,N_3268);
and U3931 (N_3931,N_3573,N_3315);
nor U3932 (N_3932,N_3410,N_3404);
nand U3933 (N_3933,N_3320,N_3567);
or U3934 (N_3934,N_3591,N_3290);
and U3935 (N_3935,N_3336,N_3239);
xnor U3936 (N_3936,N_3422,N_3272);
nor U3937 (N_3937,N_3253,N_3445);
or U3938 (N_3938,N_3571,N_3203);
and U3939 (N_3939,N_3544,N_3593);
nand U3940 (N_3940,N_3298,N_3444);
or U3941 (N_3941,N_3396,N_3429);
nor U3942 (N_3942,N_3565,N_3567);
or U3943 (N_3943,N_3569,N_3303);
xnor U3944 (N_3944,N_3462,N_3236);
xor U3945 (N_3945,N_3562,N_3493);
and U3946 (N_3946,N_3261,N_3373);
and U3947 (N_3947,N_3359,N_3579);
and U3948 (N_3948,N_3325,N_3274);
nor U3949 (N_3949,N_3216,N_3412);
nor U3950 (N_3950,N_3391,N_3429);
and U3951 (N_3951,N_3517,N_3262);
xor U3952 (N_3952,N_3413,N_3273);
or U3953 (N_3953,N_3520,N_3259);
nor U3954 (N_3954,N_3520,N_3508);
nand U3955 (N_3955,N_3549,N_3303);
or U3956 (N_3956,N_3297,N_3394);
xnor U3957 (N_3957,N_3394,N_3495);
nor U3958 (N_3958,N_3420,N_3464);
and U3959 (N_3959,N_3405,N_3517);
or U3960 (N_3960,N_3427,N_3234);
or U3961 (N_3961,N_3444,N_3551);
nor U3962 (N_3962,N_3224,N_3501);
xor U3963 (N_3963,N_3414,N_3585);
and U3964 (N_3964,N_3219,N_3578);
or U3965 (N_3965,N_3592,N_3518);
nor U3966 (N_3966,N_3410,N_3469);
xnor U3967 (N_3967,N_3452,N_3572);
nor U3968 (N_3968,N_3573,N_3401);
and U3969 (N_3969,N_3271,N_3588);
xor U3970 (N_3970,N_3480,N_3208);
xnor U3971 (N_3971,N_3251,N_3284);
xnor U3972 (N_3972,N_3389,N_3262);
xor U3973 (N_3973,N_3411,N_3572);
nand U3974 (N_3974,N_3550,N_3210);
or U3975 (N_3975,N_3328,N_3370);
nor U3976 (N_3976,N_3287,N_3513);
and U3977 (N_3977,N_3302,N_3295);
xor U3978 (N_3978,N_3482,N_3323);
nor U3979 (N_3979,N_3439,N_3226);
or U3980 (N_3980,N_3482,N_3536);
or U3981 (N_3981,N_3382,N_3455);
xnor U3982 (N_3982,N_3228,N_3554);
nand U3983 (N_3983,N_3206,N_3340);
and U3984 (N_3984,N_3270,N_3254);
and U3985 (N_3985,N_3274,N_3395);
nor U3986 (N_3986,N_3548,N_3272);
nand U3987 (N_3987,N_3516,N_3533);
and U3988 (N_3988,N_3536,N_3584);
and U3989 (N_3989,N_3232,N_3356);
xnor U3990 (N_3990,N_3319,N_3294);
nand U3991 (N_3991,N_3543,N_3572);
and U3992 (N_3992,N_3328,N_3322);
nor U3993 (N_3993,N_3408,N_3583);
and U3994 (N_3994,N_3230,N_3452);
nor U3995 (N_3995,N_3310,N_3278);
xor U3996 (N_3996,N_3423,N_3324);
xnor U3997 (N_3997,N_3304,N_3595);
and U3998 (N_3998,N_3507,N_3222);
and U3999 (N_3999,N_3254,N_3382);
nand U4000 (N_4000,N_3946,N_3891);
nand U4001 (N_4001,N_3647,N_3658);
or U4002 (N_4002,N_3986,N_3970);
nand U4003 (N_4003,N_3818,N_3764);
nor U4004 (N_4004,N_3616,N_3793);
xor U4005 (N_4005,N_3928,N_3754);
nor U4006 (N_4006,N_3856,N_3614);
nand U4007 (N_4007,N_3613,N_3819);
nor U4008 (N_4008,N_3643,N_3657);
or U4009 (N_4009,N_3915,N_3994);
nor U4010 (N_4010,N_3778,N_3889);
xnor U4011 (N_4011,N_3888,N_3779);
and U4012 (N_4012,N_3997,N_3917);
and U4013 (N_4013,N_3622,N_3831);
xnor U4014 (N_4014,N_3869,N_3874);
nand U4015 (N_4015,N_3842,N_3992);
and U4016 (N_4016,N_3908,N_3863);
nor U4017 (N_4017,N_3985,N_3822);
and U4018 (N_4018,N_3799,N_3674);
or U4019 (N_4019,N_3820,N_3884);
and U4020 (N_4020,N_3980,N_3641);
nor U4021 (N_4021,N_3781,N_3835);
nor U4022 (N_4022,N_3875,N_3911);
nand U4023 (N_4023,N_3668,N_3965);
and U4024 (N_4024,N_3853,N_3769);
or U4025 (N_4025,N_3857,N_3787);
or U4026 (N_4026,N_3731,N_3852);
xor U4027 (N_4027,N_3768,N_3677);
xor U4028 (N_4028,N_3619,N_3810);
and U4029 (N_4029,N_3930,N_3605);
and U4030 (N_4030,N_3881,N_3895);
xor U4031 (N_4031,N_3757,N_3760);
xor U4032 (N_4032,N_3692,N_3618);
nand U4033 (N_4033,N_3938,N_3897);
xor U4034 (N_4034,N_3995,N_3828);
nand U4035 (N_4035,N_3709,N_3685);
or U4036 (N_4036,N_3808,N_3752);
nor U4037 (N_4037,N_3950,N_3681);
xnor U4038 (N_4038,N_3940,N_3639);
or U4039 (N_4039,N_3987,N_3607);
xnor U4040 (N_4040,N_3979,N_3748);
nor U4041 (N_4041,N_3784,N_3664);
nand U4042 (N_4042,N_3785,N_3803);
nor U4043 (N_4043,N_3601,N_3813);
xnor U4044 (N_4044,N_3976,N_3719);
nor U4045 (N_4045,N_3743,N_3916);
nand U4046 (N_4046,N_3659,N_3814);
or U4047 (N_4047,N_3633,N_3744);
and U4048 (N_4048,N_3967,N_3772);
xor U4049 (N_4049,N_3998,N_3626);
or U4050 (N_4050,N_3766,N_3996);
xnor U4051 (N_4051,N_3661,N_3735);
nor U4052 (N_4052,N_3617,N_3797);
and U4053 (N_4053,N_3937,N_3761);
or U4054 (N_4054,N_3859,N_3910);
nand U4055 (N_4055,N_3839,N_3654);
xor U4056 (N_4056,N_3829,N_3697);
xor U4057 (N_4057,N_3783,N_3836);
xnor U4058 (N_4058,N_3920,N_3759);
xor U4059 (N_4059,N_3826,N_3890);
or U4060 (N_4060,N_3963,N_3846);
nor U4061 (N_4061,N_3789,N_3882);
nand U4062 (N_4062,N_3901,N_3900);
xnor U4063 (N_4063,N_3947,N_3800);
xor U4064 (N_4064,N_3913,N_3712);
or U4065 (N_4065,N_3717,N_3838);
xnor U4066 (N_4066,N_3955,N_3790);
xnor U4067 (N_4067,N_3956,N_3713);
nand U4068 (N_4068,N_3740,N_3922);
xnor U4069 (N_4069,N_3868,N_3816);
xor U4070 (N_4070,N_3720,N_3791);
nor U4071 (N_4071,N_3912,N_3724);
nand U4072 (N_4072,N_3612,N_3929);
xnor U4073 (N_4073,N_3688,N_3861);
nor U4074 (N_4074,N_3615,N_3708);
nand U4075 (N_4075,N_3858,N_3945);
and U4076 (N_4076,N_3958,N_3939);
or U4077 (N_4077,N_3646,N_3952);
xnor U4078 (N_4078,N_3978,N_3725);
nand U4079 (N_4079,N_3966,N_3726);
nor U4080 (N_4080,N_3722,N_3974);
nor U4081 (N_4081,N_3666,N_3749);
or U4082 (N_4082,N_3732,N_3737);
and U4083 (N_4083,N_3751,N_3848);
xnor U4084 (N_4084,N_3621,N_3623);
and U4085 (N_4085,N_3756,N_3683);
nor U4086 (N_4086,N_3843,N_3642);
xor U4087 (N_4087,N_3798,N_3951);
and U4088 (N_4088,N_3933,N_3854);
nand U4089 (N_4089,N_3753,N_3672);
nor U4090 (N_4090,N_3993,N_3892);
nand U4091 (N_4091,N_3703,N_3871);
xor U4092 (N_4092,N_3801,N_3669);
nand U4093 (N_4093,N_3960,N_3921);
and U4094 (N_4094,N_3651,N_3811);
or U4095 (N_4095,N_3847,N_3765);
or U4096 (N_4096,N_3600,N_3827);
nand U4097 (N_4097,N_3638,N_3834);
nand U4098 (N_4098,N_3699,N_3809);
or U4099 (N_4099,N_3865,N_3914);
and U4100 (N_4100,N_3653,N_3776);
xnor U4101 (N_4101,N_3948,N_3625);
xnor U4102 (N_4102,N_3935,N_3794);
or U4103 (N_4103,N_3629,N_3782);
nand U4104 (N_4104,N_3775,N_3927);
and U4105 (N_4105,N_3953,N_3807);
nor U4106 (N_4106,N_3870,N_3670);
and U4107 (N_4107,N_3893,N_3802);
and U4108 (N_4108,N_3907,N_3841);
nor U4109 (N_4109,N_3705,N_3867);
nand U4110 (N_4110,N_3902,N_3806);
and U4111 (N_4111,N_3990,N_3758);
and U4112 (N_4112,N_3701,N_3873);
and U4113 (N_4113,N_3736,N_3886);
nand U4114 (N_4114,N_3649,N_3704);
nand U4115 (N_4115,N_3932,N_3747);
xor U4116 (N_4116,N_3795,N_3942);
nand U4117 (N_4117,N_3718,N_3849);
nand U4118 (N_4118,N_3792,N_3983);
xor U4119 (N_4119,N_3796,N_3606);
and U4120 (N_4120,N_3924,N_3648);
and U4121 (N_4121,N_3624,N_3608);
and U4122 (N_4122,N_3714,N_3679);
xor U4123 (N_4123,N_3943,N_3788);
nor U4124 (N_4124,N_3899,N_3830);
or U4125 (N_4125,N_3894,N_3691);
and U4126 (N_4126,N_3815,N_3962);
nand U4127 (N_4127,N_3931,N_3905);
nand U4128 (N_4128,N_3773,N_3898);
and U4129 (N_4129,N_3862,N_3663);
and U4130 (N_4130,N_3696,N_3972);
nand U4131 (N_4131,N_3655,N_3635);
nor U4132 (N_4132,N_3727,N_3650);
nand U4133 (N_4133,N_3973,N_3729);
and U4134 (N_4134,N_3968,N_3887);
and U4135 (N_4135,N_3770,N_3872);
or U4136 (N_4136,N_3684,N_3989);
nand U4137 (N_4137,N_3777,N_3825);
and U4138 (N_4138,N_3604,N_3975);
xor U4139 (N_4139,N_3711,N_3755);
nor U4140 (N_4140,N_3812,N_3961);
nor U4141 (N_4141,N_3730,N_3762);
and U4142 (N_4142,N_3750,N_3675);
nor U4143 (N_4143,N_3671,N_3738);
nor U4144 (N_4144,N_3774,N_3906);
and U4145 (N_4145,N_3926,N_3767);
or U4146 (N_4146,N_3925,N_3686);
xnor U4147 (N_4147,N_3602,N_3860);
and U4148 (N_4148,N_3630,N_3728);
xnor U4149 (N_4149,N_3878,N_3833);
nor U4150 (N_4150,N_3866,N_3662);
nand U4151 (N_4151,N_3982,N_3676);
and U4152 (N_4152,N_3876,N_3954);
or U4153 (N_4153,N_3636,N_3631);
xor U4154 (N_4154,N_3620,N_3823);
nand U4155 (N_4155,N_3851,N_3637);
nor U4156 (N_4156,N_3904,N_3941);
nand U4157 (N_4157,N_3628,N_3879);
or U4158 (N_4158,N_3690,N_3780);
or U4159 (N_4159,N_3885,N_3864);
nor U4160 (N_4160,N_3880,N_3909);
or U4161 (N_4161,N_3644,N_3923);
nand U4162 (N_4162,N_3964,N_3919);
and U4163 (N_4163,N_3999,N_3733);
xnor U4164 (N_4164,N_3610,N_3949);
or U4165 (N_4165,N_3609,N_3603);
xnor U4166 (N_4166,N_3786,N_3832);
or U4167 (N_4167,N_3734,N_3693);
nor U4168 (N_4168,N_3805,N_3840);
and U4169 (N_4169,N_3632,N_3745);
xor U4170 (N_4170,N_3821,N_3746);
xnor U4171 (N_4171,N_3845,N_3660);
or U4172 (N_4172,N_3971,N_3896);
xor U4173 (N_4173,N_3689,N_3977);
nor U4174 (N_4174,N_3640,N_3716);
xnor U4175 (N_4175,N_3883,N_3959);
xnor U4176 (N_4176,N_3824,N_3665);
xor U4177 (N_4177,N_3936,N_3877);
xnor U4178 (N_4178,N_3981,N_3715);
and U4179 (N_4179,N_3702,N_3678);
nand U4180 (N_4180,N_3627,N_3804);
xnor U4181 (N_4181,N_3850,N_3652);
nand U4182 (N_4182,N_3687,N_3721);
xnor U4183 (N_4183,N_3944,N_3742);
xnor U4184 (N_4184,N_3984,N_3969);
and U4185 (N_4185,N_3695,N_3723);
nor U4186 (N_4186,N_3634,N_3771);
and U4187 (N_4187,N_3673,N_3707);
xor U4188 (N_4188,N_3656,N_3645);
nor U4189 (N_4189,N_3855,N_3934);
nor U4190 (N_4190,N_3741,N_3694);
nor U4191 (N_4191,N_3957,N_3710);
or U4192 (N_4192,N_3837,N_3918);
nor U4193 (N_4193,N_3682,N_3739);
xnor U4194 (N_4194,N_3611,N_3817);
or U4195 (N_4195,N_3700,N_3680);
nand U4196 (N_4196,N_3844,N_3698);
and U4197 (N_4197,N_3763,N_3667);
nor U4198 (N_4198,N_3988,N_3991);
xor U4199 (N_4199,N_3903,N_3706);
xor U4200 (N_4200,N_3602,N_3894);
or U4201 (N_4201,N_3966,N_3671);
nand U4202 (N_4202,N_3863,N_3697);
or U4203 (N_4203,N_3896,N_3741);
and U4204 (N_4204,N_3662,N_3752);
and U4205 (N_4205,N_3718,N_3730);
xnor U4206 (N_4206,N_3704,N_3811);
nand U4207 (N_4207,N_3610,N_3656);
nor U4208 (N_4208,N_3845,N_3813);
nor U4209 (N_4209,N_3924,N_3914);
nor U4210 (N_4210,N_3776,N_3630);
or U4211 (N_4211,N_3630,N_3757);
or U4212 (N_4212,N_3900,N_3956);
xor U4213 (N_4213,N_3846,N_3947);
nand U4214 (N_4214,N_3938,N_3999);
nor U4215 (N_4215,N_3915,N_3613);
and U4216 (N_4216,N_3852,N_3791);
nand U4217 (N_4217,N_3739,N_3925);
xnor U4218 (N_4218,N_3855,N_3858);
nor U4219 (N_4219,N_3908,N_3836);
and U4220 (N_4220,N_3818,N_3819);
xor U4221 (N_4221,N_3813,N_3854);
nand U4222 (N_4222,N_3884,N_3868);
nor U4223 (N_4223,N_3753,N_3640);
and U4224 (N_4224,N_3824,N_3935);
xor U4225 (N_4225,N_3909,N_3853);
nand U4226 (N_4226,N_3987,N_3742);
xor U4227 (N_4227,N_3690,N_3639);
xnor U4228 (N_4228,N_3646,N_3906);
xor U4229 (N_4229,N_3767,N_3820);
or U4230 (N_4230,N_3887,N_3811);
nand U4231 (N_4231,N_3902,N_3968);
xor U4232 (N_4232,N_3706,N_3935);
xor U4233 (N_4233,N_3762,N_3720);
nor U4234 (N_4234,N_3864,N_3912);
and U4235 (N_4235,N_3961,N_3627);
nor U4236 (N_4236,N_3959,N_3984);
and U4237 (N_4237,N_3850,N_3614);
nor U4238 (N_4238,N_3858,N_3785);
or U4239 (N_4239,N_3986,N_3849);
or U4240 (N_4240,N_3880,N_3628);
xor U4241 (N_4241,N_3862,N_3738);
or U4242 (N_4242,N_3716,N_3741);
and U4243 (N_4243,N_3636,N_3614);
nor U4244 (N_4244,N_3979,N_3801);
and U4245 (N_4245,N_3662,N_3857);
nand U4246 (N_4246,N_3916,N_3682);
nand U4247 (N_4247,N_3845,N_3882);
nor U4248 (N_4248,N_3967,N_3947);
xnor U4249 (N_4249,N_3809,N_3777);
nor U4250 (N_4250,N_3783,N_3791);
nor U4251 (N_4251,N_3733,N_3700);
nor U4252 (N_4252,N_3676,N_3975);
nor U4253 (N_4253,N_3962,N_3712);
xnor U4254 (N_4254,N_3619,N_3718);
nand U4255 (N_4255,N_3714,N_3656);
xnor U4256 (N_4256,N_3764,N_3908);
xnor U4257 (N_4257,N_3982,N_3873);
nor U4258 (N_4258,N_3801,N_3792);
nor U4259 (N_4259,N_3714,N_3764);
or U4260 (N_4260,N_3885,N_3656);
and U4261 (N_4261,N_3784,N_3774);
or U4262 (N_4262,N_3878,N_3943);
nor U4263 (N_4263,N_3957,N_3908);
xor U4264 (N_4264,N_3890,N_3650);
xnor U4265 (N_4265,N_3818,N_3761);
nand U4266 (N_4266,N_3727,N_3632);
nand U4267 (N_4267,N_3679,N_3768);
and U4268 (N_4268,N_3921,N_3948);
nor U4269 (N_4269,N_3984,N_3752);
nor U4270 (N_4270,N_3866,N_3878);
and U4271 (N_4271,N_3637,N_3756);
and U4272 (N_4272,N_3982,N_3809);
or U4273 (N_4273,N_3646,N_3799);
or U4274 (N_4274,N_3659,N_3798);
nand U4275 (N_4275,N_3941,N_3713);
nor U4276 (N_4276,N_3885,N_3887);
nor U4277 (N_4277,N_3638,N_3802);
xor U4278 (N_4278,N_3848,N_3768);
nor U4279 (N_4279,N_3971,N_3618);
or U4280 (N_4280,N_3981,N_3930);
nor U4281 (N_4281,N_3935,N_3876);
or U4282 (N_4282,N_3645,N_3793);
and U4283 (N_4283,N_3694,N_3850);
nand U4284 (N_4284,N_3853,N_3885);
xor U4285 (N_4285,N_3827,N_3826);
nand U4286 (N_4286,N_3629,N_3836);
and U4287 (N_4287,N_3855,N_3971);
nor U4288 (N_4288,N_3691,N_3929);
nand U4289 (N_4289,N_3606,N_3660);
and U4290 (N_4290,N_3831,N_3821);
nand U4291 (N_4291,N_3954,N_3927);
nand U4292 (N_4292,N_3939,N_3635);
xor U4293 (N_4293,N_3957,N_3842);
nor U4294 (N_4294,N_3680,N_3862);
or U4295 (N_4295,N_3659,N_3768);
nor U4296 (N_4296,N_3677,N_3892);
and U4297 (N_4297,N_3677,N_3808);
and U4298 (N_4298,N_3941,N_3609);
and U4299 (N_4299,N_3715,N_3774);
or U4300 (N_4300,N_3799,N_3826);
nor U4301 (N_4301,N_3725,N_3643);
nor U4302 (N_4302,N_3691,N_3637);
xnor U4303 (N_4303,N_3827,N_3719);
and U4304 (N_4304,N_3709,N_3984);
and U4305 (N_4305,N_3773,N_3890);
xor U4306 (N_4306,N_3970,N_3865);
or U4307 (N_4307,N_3721,N_3816);
xor U4308 (N_4308,N_3865,N_3817);
nor U4309 (N_4309,N_3749,N_3622);
nand U4310 (N_4310,N_3926,N_3683);
xor U4311 (N_4311,N_3897,N_3691);
or U4312 (N_4312,N_3865,N_3658);
and U4313 (N_4313,N_3703,N_3769);
nor U4314 (N_4314,N_3818,N_3996);
and U4315 (N_4315,N_3780,N_3995);
or U4316 (N_4316,N_3725,N_3924);
and U4317 (N_4317,N_3877,N_3792);
xnor U4318 (N_4318,N_3814,N_3970);
xnor U4319 (N_4319,N_3695,N_3842);
nor U4320 (N_4320,N_3755,N_3953);
or U4321 (N_4321,N_3743,N_3795);
and U4322 (N_4322,N_3760,N_3910);
or U4323 (N_4323,N_3788,N_3976);
xor U4324 (N_4324,N_3728,N_3916);
xnor U4325 (N_4325,N_3862,N_3800);
nand U4326 (N_4326,N_3638,N_3659);
nand U4327 (N_4327,N_3835,N_3944);
nand U4328 (N_4328,N_3606,N_3908);
xnor U4329 (N_4329,N_3929,N_3977);
nor U4330 (N_4330,N_3751,N_3851);
nor U4331 (N_4331,N_3949,N_3953);
nor U4332 (N_4332,N_3697,N_3834);
nor U4333 (N_4333,N_3713,N_3890);
nor U4334 (N_4334,N_3759,N_3638);
nor U4335 (N_4335,N_3691,N_3923);
or U4336 (N_4336,N_3689,N_3974);
nand U4337 (N_4337,N_3884,N_3930);
xor U4338 (N_4338,N_3705,N_3731);
or U4339 (N_4339,N_3841,N_3962);
nor U4340 (N_4340,N_3733,N_3709);
or U4341 (N_4341,N_3747,N_3920);
and U4342 (N_4342,N_3849,N_3724);
nor U4343 (N_4343,N_3608,N_3983);
nor U4344 (N_4344,N_3810,N_3637);
nand U4345 (N_4345,N_3890,N_3815);
xor U4346 (N_4346,N_3666,N_3746);
xor U4347 (N_4347,N_3708,N_3736);
and U4348 (N_4348,N_3996,N_3609);
nand U4349 (N_4349,N_3914,N_3848);
nand U4350 (N_4350,N_3988,N_3604);
and U4351 (N_4351,N_3797,N_3832);
or U4352 (N_4352,N_3860,N_3940);
nand U4353 (N_4353,N_3850,N_3729);
nand U4354 (N_4354,N_3778,N_3884);
nor U4355 (N_4355,N_3695,N_3943);
or U4356 (N_4356,N_3684,N_3958);
and U4357 (N_4357,N_3988,N_3888);
xnor U4358 (N_4358,N_3931,N_3901);
and U4359 (N_4359,N_3646,N_3911);
or U4360 (N_4360,N_3743,N_3765);
nor U4361 (N_4361,N_3793,N_3831);
or U4362 (N_4362,N_3689,N_3973);
nor U4363 (N_4363,N_3889,N_3670);
and U4364 (N_4364,N_3878,N_3979);
nor U4365 (N_4365,N_3639,N_3779);
nor U4366 (N_4366,N_3635,N_3904);
xnor U4367 (N_4367,N_3653,N_3990);
and U4368 (N_4368,N_3775,N_3720);
and U4369 (N_4369,N_3725,N_3806);
nand U4370 (N_4370,N_3645,N_3842);
or U4371 (N_4371,N_3810,N_3622);
nor U4372 (N_4372,N_3958,N_3905);
nor U4373 (N_4373,N_3857,N_3648);
nand U4374 (N_4374,N_3650,N_3619);
xnor U4375 (N_4375,N_3825,N_3717);
nor U4376 (N_4376,N_3790,N_3984);
nand U4377 (N_4377,N_3681,N_3774);
nand U4378 (N_4378,N_3844,N_3633);
nor U4379 (N_4379,N_3771,N_3817);
nand U4380 (N_4380,N_3942,N_3820);
or U4381 (N_4381,N_3724,N_3968);
and U4382 (N_4382,N_3985,N_3781);
or U4383 (N_4383,N_3984,N_3928);
or U4384 (N_4384,N_3689,N_3902);
or U4385 (N_4385,N_3609,N_3806);
nand U4386 (N_4386,N_3679,N_3955);
xor U4387 (N_4387,N_3857,N_3761);
nand U4388 (N_4388,N_3807,N_3981);
nor U4389 (N_4389,N_3775,N_3897);
xor U4390 (N_4390,N_3740,N_3752);
or U4391 (N_4391,N_3987,N_3648);
nand U4392 (N_4392,N_3725,N_3894);
nor U4393 (N_4393,N_3922,N_3622);
nor U4394 (N_4394,N_3671,N_3861);
and U4395 (N_4395,N_3791,N_3665);
and U4396 (N_4396,N_3826,N_3978);
or U4397 (N_4397,N_3684,N_3817);
xor U4398 (N_4398,N_3891,N_3744);
nor U4399 (N_4399,N_3606,N_3970);
nor U4400 (N_4400,N_4235,N_4043);
nor U4401 (N_4401,N_4119,N_4292);
or U4402 (N_4402,N_4349,N_4357);
nand U4403 (N_4403,N_4014,N_4037);
nand U4404 (N_4404,N_4003,N_4098);
and U4405 (N_4405,N_4061,N_4040);
nand U4406 (N_4406,N_4064,N_4175);
nor U4407 (N_4407,N_4232,N_4179);
nor U4408 (N_4408,N_4122,N_4218);
nand U4409 (N_4409,N_4124,N_4009);
or U4410 (N_4410,N_4373,N_4036);
nor U4411 (N_4411,N_4144,N_4103);
nor U4412 (N_4412,N_4159,N_4306);
nand U4413 (N_4413,N_4033,N_4273);
and U4414 (N_4414,N_4184,N_4131);
and U4415 (N_4415,N_4091,N_4125);
nand U4416 (N_4416,N_4007,N_4332);
nor U4417 (N_4417,N_4345,N_4303);
nor U4418 (N_4418,N_4266,N_4284);
xor U4419 (N_4419,N_4379,N_4169);
nor U4420 (N_4420,N_4153,N_4154);
nor U4421 (N_4421,N_4073,N_4195);
or U4422 (N_4422,N_4164,N_4028);
xnor U4423 (N_4423,N_4324,N_4145);
or U4424 (N_4424,N_4127,N_4060);
xor U4425 (N_4425,N_4287,N_4253);
or U4426 (N_4426,N_4078,N_4305);
nor U4427 (N_4427,N_4231,N_4076);
nand U4428 (N_4428,N_4258,N_4369);
nand U4429 (N_4429,N_4215,N_4044);
nand U4430 (N_4430,N_4167,N_4304);
or U4431 (N_4431,N_4170,N_4364);
nor U4432 (N_4432,N_4294,N_4228);
nor U4433 (N_4433,N_4263,N_4210);
nand U4434 (N_4434,N_4199,N_4398);
nor U4435 (N_4435,N_4281,N_4390);
and U4436 (N_4436,N_4217,N_4270);
and U4437 (N_4437,N_4381,N_4027);
and U4438 (N_4438,N_4155,N_4185);
and U4439 (N_4439,N_4276,N_4102);
or U4440 (N_4440,N_4180,N_4008);
xnor U4441 (N_4441,N_4205,N_4326);
nor U4442 (N_4442,N_4149,N_4242);
and U4443 (N_4443,N_4069,N_4178);
or U4444 (N_4444,N_4212,N_4322);
xnor U4445 (N_4445,N_4187,N_4338);
or U4446 (N_4446,N_4116,N_4348);
nor U4447 (N_4447,N_4042,N_4307);
and U4448 (N_4448,N_4331,N_4347);
nand U4449 (N_4449,N_4298,N_4255);
xor U4450 (N_4450,N_4237,N_4090);
nand U4451 (N_4451,N_4084,N_4129);
or U4452 (N_4452,N_4196,N_4296);
nor U4453 (N_4453,N_4362,N_4146);
and U4454 (N_4454,N_4058,N_4280);
xnor U4455 (N_4455,N_4189,N_4101);
xnor U4456 (N_4456,N_4117,N_4399);
nor U4457 (N_4457,N_4262,N_4055);
nor U4458 (N_4458,N_4039,N_4285);
nor U4459 (N_4459,N_4290,N_4275);
or U4460 (N_4460,N_4063,N_4236);
and U4461 (N_4461,N_4261,N_4260);
xor U4462 (N_4462,N_4100,N_4315);
xor U4463 (N_4463,N_4227,N_4051);
and U4464 (N_4464,N_4107,N_4319);
xor U4465 (N_4465,N_4222,N_4297);
or U4466 (N_4466,N_4291,N_4377);
and U4467 (N_4467,N_4372,N_4134);
nand U4468 (N_4468,N_4375,N_4193);
and U4469 (N_4469,N_4109,N_4035);
nand U4470 (N_4470,N_4111,N_4209);
nor U4471 (N_4471,N_4163,N_4165);
nand U4472 (N_4472,N_4320,N_4392);
or U4473 (N_4473,N_4239,N_4395);
nor U4474 (N_4474,N_4360,N_4389);
nand U4475 (N_4475,N_4343,N_4085);
and U4476 (N_4476,N_4310,N_4207);
and U4477 (N_4477,N_4350,N_4341);
and U4478 (N_4478,N_4220,N_4197);
nand U4479 (N_4479,N_4191,N_4230);
nand U4480 (N_4480,N_4151,N_4378);
nor U4481 (N_4481,N_4138,N_4142);
and U4482 (N_4482,N_4206,N_4160);
or U4483 (N_4483,N_4268,N_4106);
and U4484 (N_4484,N_4264,N_4030);
xor U4485 (N_4485,N_4295,N_4046);
xnor U4486 (N_4486,N_4249,N_4173);
nand U4487 (N_4487,N_4045,N_4004);
nand U4488 (N_4488,N_4000,N_4265);
nand U4489 (N_4489,N_4067,N_4359);
nor U4490 (N_4490,N_4087,N_4133);
nand U4491 (N_4491,N_4309,N_4023);
and U4492 (N_4492,N_4182,N_4120);
nand U4493 (N_4493,N_4074,N_4204);
nand U4494 (N_4494,N_4346,N_4066);
xnor U4495 (N_4495,N_4384,N_4325);
and U4496 (N_4496,N_4137,N_4024);
nor U4497 (N_4497,N_4368,N_4128);
or U4498 (N_4498,N_4010,N_4118);
xor U4499 (N_4499,N_4140,N_4246);
and U4500 (N_4500,N_4080,N_4286);
xnor U4501 (N_4501,N_4257,N_4186);
or U4502 (N_4502,N_4011,N_4302);
nand U4503 (N_4503,N_4351,N_4086);
and U4504 (N_4504,N_4370,N_4354);
or U4505 (N_4505,N_4225,N_4130);
and U4506 (N_4506,N_4157,N_4089);
xor U4507 (N_4507,N_4203,N_4147);
nor U4508 (N_4508,N_4136,N_4070);
xnor U4509 (N_4509,N_4126,N_4022);
and U4510 (N_4510,N_4054,N_4172);
nand U4511 (N_4511,N_4282,N_4123);
or U4512 (N_4512,N_4358,N_4352);
or U4513 (N_4513,N_4079,N_4293);
or U4514 (N_4514,N_4200,N_4015);
or U4515 (N_4515,N_4355,N_4081);
nand U4516 (N_4516,N_4301,N_4314);
and U4517 (N_4517,N_4254,N_4386);
xor U4518 (N_4518,N_4077,N_4397);
or U4519 (N_4519,N_4244,N_4376);
and U4520 (N_4520,N_4267,N_4393);
and U4521 (N_4521,N_4213,N_4367);
or U4522 (N_4522,N_4248,N_4238);
nor U4523 (N_4523,N_4374,N_4323);
or U4524 (N_4524,N_4018,N_4247);
xnor U4525 (N_4525,N_4176,N_4013);
and U4526 (N_4526,N_4068,N_4313);
nor U4527 (N_4527,N_4095,N_4034);
and U4528 (N_4528,N_4016,N_4334);
nor U4529 (N_4529,N_4094,N_4216);
nor U4530 (N_4530,N_4391,N_4041);
xnor U4531 (N_4531,N_4214,N_4156);
and U4532 (N_4532,N_4245,N_4083);
and U4533 (N_4533,N_4056,N_4071);
nand U4534 (N_4534,N_4190,N_4300);
nand U4535 (N_4535,N_4366,N_4002);
and U4536 (N_4536,N_4387,N_4219);
or U4537 (N_4537,N_4113,N_4208);
nor U4538 (N_4538,N_4283,N_4330);
xnor U4539 (N_4539,N_4017,N_4318);
and U4540 (N_4540,N_4031,N_4234);
xnor U4541 (N_4541,N_4029,N_4135);
xor U4542 (N_4542,N_4168,N_4050);
nor U4543 (N_4543,N_4224,N_4032);
nor U4544 (N_4544,N_4006,N_4026);
nand U4545 (N_4545,N_4139,N_4394);
and U4546 (N_4546,N_4361,N_4177);
nand U4547 (N_4547,N_4241,N_4328);
nand U4548 (N_4548,N_4308,N_4088);
nand U4549 (N_4549,N_4166,N_4344);
xor U4550 (N_4550,N_4382,N_4271);
or U4551 (N_4551,N_4161,N_4251);
nand U4552 (N_4552,N_4108,N_4082);
xor U4553 (N_4553,N_4048,N_4380);
nand U4554 (N_4554,N_4259,N_4025);
or U4555 (N_4555,N_4223,N_4150);
and U4556 (N_4556,N_4112,N_4115);
nor U4557 (N_4557,N_4057,N_4152);
nor U4558 (N_4558,N_4385,N_4049);
xor U4559 (N_4559,N_4299,N_4202);
nand U4560 (N_4560,N_4194,N_4141);
xor U4561 (N_4561,N_4277,N_4311);
and U4562 (N_4562,N_4047,N_4226);
or U4563 (N_4563,N_4337,N_4132);
or U4564 (N_4564,N_4019,N_4038);
nand U4565 (N_4565,N_4121,N_4012);
nand U4566 (N_4566,N_4110,N_4221);
nand U4567 (N_4567,N_4105,N_4252);
nand U4568 (N_4568,N_4396,N_4339);
xor U4569 (N_4569,N_4053,N_4188);
nand U4570 (N_4570,N_4062,N_4059);
xnor U4571 (N_4571,N_4329,N_4288);
nor U4572 (N_4572,N_4274,N_4229);
and U4573 (N_4573,N_4092,N_4183);
or U4574 (N_4574,N_4336,N_4340);
or U4575 (N_4575,N_4192,N_4371);
and U4576 (N_4576,N_4356,N_4279);
nand U4577 (N_4577,N_4021,N_4335);
nand U4578 (N_4578,N_4099,N_4001);
xor U4579 (N_4579,N_4201,N_4321);
nand U4580 (N_4580,N_4233,N_4174);
nand U4581 (N_4581,N_4052,N_4316);
and U4582 (N_4582,N_4317,N_4148);
xnor U4583 (N_4583,N_4333,N_4342);
nand U4584 (N_4584,N_4289,N_4240);
or U4585 (N_4585,N_4181,N_4243);
and U4586 (N_4586,N_4093,N_4256);
nand U4587 (N_4587,N_4162,N_4272);
nand U4588 (N_4588,N_4327,N_4198);
nand U4589 (N_4589,N_4114,N_4353);
xnor U4590 (N_4590,N_4143,N_4388);
nor U4591 (N_4591,N_4075,N_4211);
and U4592 (N_4592,N_4363,N_4269);
xnor U4593 (N_4593,N_4096,N_4158);
and U4594 (N_4594,N_4104,N_4365);
xnor U4595 (N_4595,N_4065,N_4005);
xnor U4596 (N_4596,N_4250,N_4072);
or U4597 (N_4597,N_4020,N_4171);
nand U4598 (N_4598,N_4097,N_4383);
or U4599 (N_4599,N_4278,N_4312);
nand U4600 (N_4600,N_4128,N_4296);
nor U4601 (N_4601,N_4283,N_4258);
nor U4602 (N_4602,N_4220,N_4239);
xor U4603 (N_4603,N_4203,N_4370);
nand U4604 (N_4604,N_4351,N_4185);
and U4605 (N_4605,N_4350,N_4273);
xor U4606 (N_4606,N_4012,N_4094);
nor U4607 (N_4607,N_4000,N_4043);
nand U4608 (N_4608,N_4172,N_4163);
xnor U4609 (N_4609,N_4335,N_4082);
nand U4610 (N_4610,N_4093,N_4350);
and U4611 (N_4611,N_4222,N_4072);
or U4612 (N_4612,N_4213,N_4358);
xor U4613 (N_4613,N_4346,N_4017);
nand U4614 (N_4614,N_4069,N_4256);
xnor U4615 (N_4615,N_4262,N_4287);
nor U4616 (N_4616,N_4280,N_4326);
and U4617 (N_4617,N_4290,N_4211);
nor U4618 (N_4618,N_4179,N_4368);
xnor U4619 (N_4619,N_4218,N_4079);
or U4620 (N_4620,N_4248,N_4300);
nor U4621 (N_4621,N_4394,N_4145);
nor U4622 (N_4622,N_4028,N_4107);
and U4623 (N_4623,N_4149,N_4076);
or U4624 (N_4624,N_4038,N_4160);
or U4625 (N_4625,N_4012,N_4234);
or U4626 (N_4626,N_4326,N_4101);
or U4627 (N_4627,N_4198,N_4183);
or U4628 (N_4628,N_4020,N_4220);
or U4629 (N_4629,N_4086,N_4388);
or U4630 (N_4630,N_4072,N_4077);
and U4631 (N_4631,N_4069,N_4368);
or U4632 (N_4632,N_4103,N_4161);
and U4633 (N_4633,N_4177,N_4048);
and U4634 (N_4634,N_4038,N_4020);
nor U4635 (N_4635,N_4192,N_4379);
and U4636 (N_4636,N_4185,N_4132);
xor U4637 (N_4637,N_4338,N_4032);
nand U4638 (N_4638,N_4225,N_4355);
xor U4639 (N_4639,N_4198,N_4278);
nor U4640 (N_4640,N_4310,N_4231);
nand U4641 (N_4641,N_4379,N_4115);
or U4642 (N_4642,N_4278,N_4326);
nor U4643 (N_4643,N_4138,N_4080);
or U4644 (N_4644,N_4087,N_4011);
nand U4645 (N_4645,N_4243,N_4197);
or U4646 (N_4646,N_4378,N_4121);
nor U4647 (N_4647,N_4237,N_4313);
or U4648 (N_4648,N_4263,N_4204);
or U4649 (N_4649,N_4392,N_4134);
nand U4650 (N_4650,N_4252,N_4372);
and U4651 (N_4651,N_4046,N_4319);
nor U4652 (N_4652,N_4211,N_4150);
xor U4653 (N_4653,N_4014,N_4095);
nand U4654 (N_4654,N_4088,N_4144);
and U4655 (N_4655,N_4286,N_4376);
xnor U4656 (N_4656,N_4074,N_4128);
nand U4657 (N_4657,N_4075,N_4254);
xnor U4658 (N_4658,N_4057,N_4248);
nand U4659 (N_4659,N_4172,N_4217);
and U4660 (N_4660,N_4063,N_4362);
nor U4661 (N_4661,N_4129,N_4025);
nor U4662 (N_4662,N_4037,N_4032);
xor U4663 (N_4663,N_4093,N_4045);
or U4664 (N_4664,N_4121,N_4318);
and U4665 (N_4665,N_4193,N_4089);
or U4666 (N_4666,N_4181,N_4388);
and U4667 (N_4667,N_4142,N_4394);
and U4668 (N_4668,N_4242,N_4167);
xnor U4669 (N_4669,N_4351,N_4330);
xnor U4670 (N_4670,N_4152,N_4309);
nor U4671 (N_4671,N_4040,N_4372);
xor U4672 (N_4672,N_4200,N_4273);
nand U4673 (N_4673,N_4087,N_4283);
or U4674 (N_4674,N_4329,N_4388);
nand U4675 (N_4675,N_4286,N_4322);
or U4676 (N_4676,N_4209,N_4350);
xor U4677 (N_4677,N_4184,N_4067);
or U4678 (N_4678,N_4357,N_4380);
xnor U4679 (N_4679,N_4310,N_4216);
nor U4680 (N_4680,N_4376,N_4104);
nand U4681 (N_4681,N_4259,N_4122);
and U4682 (N_4682,N_4141,N_4059);
nor U4683 (N_4683,N_4316,N_4169);
nor U4684 (N_4684,N_4173,N_4103);
nand U4685 (N_4685,N_4240,N_4367);
nor U4686 (N_4686,N_4004,N_4358);
nand U4687 (N_4687,N_4073,N_4163);
or U4688 (N_4688,N_4044,N_4174);
or U4689 (N_4689,N_4374,N_4068);
and U4690 (N_4690,N_4386,N_4005);
and U4691 (N_4691,N_4330,N_4053);
xnor U4692 (N_4692,N_4081,N_4257);
nor U4693 (N_4693,N_4366,N_4145);
or U4694 (N_4694,N_4357,N_4045);
or U4695 (N_4695,N_4396,N_4088);
xnor U4696 (N_4696,N_4194,N_4188);
nor U4697 (N_4697,N_4108,N_4090);
and U4698 (N_4698,N_4092,N_4046);
nor U4699 (N_4699,N_4186,N_4298);
xnor U4700 (N_4700,N_4364,N_4128);
or U4701 (N_4701,N_4054,N_4222);
or U4702 (N_4702,N_4069,N_4191);
nor U4703 (N_4703,N_4214,N_4084);
or U4704 (N_4704,N_4335,N_4240);
and U4705 (N_4705,N_4301,N_4331);
and U4706 (N_4706,N_4103,N_4304);
xor U4707 (N_4707,N_4129,N_4028);
nand U4708 (N_4708,N_4105,N_4206);
nor U4709 (N_4709,N_4214,N_4322);
nand U4710 (N_4710,N_4307,N_4229);
nand U4711 (N_4711,N_4137,N_4211);
or U4712 (N_4712,N_4327,N_4069);
and U4713 (N_4713,N_4341,N_4326);
nor U4714 (N_4714,N_4365,N_4089);
nand U4715 (N_4715,N_4337,N_4331);
or U4716 (N_4716,N_4180,N_4207);
and U4717 (N_4717,N_4376,N_4384);
xor U4718 (N_4718,N_4106,N_4287);
or U4719 (N_4719,N_4077,N_4198);
nand U4720 (N_4720,N_4174,N_4386);
or U4721 (N_4721,N_4118,N_4368);
and U4722 (N_4722,N_4011,N_4304);
nor U4723 (N_4723,N_4029,N_4169);
nor U4724 (N_4724,N_4136,N_4280);
nor U4725 (N_4725,N_4314,N_4062);
or U4726 (N_4726,N_4351,N_4053);
and U4727 (N_4727,N_4137,N_4394);
or U4728 (N_4728,N_4136,N_4277);
or U4729 (N_4729,N_4377,N_4021);
nand U4730 (N_4730,N_4339,N_4325);
xor U4731 (N_4731,N_4023,N_4381);
xor U4732 (N_4732,N_4218,N_4113);
xnor U4733 (N_4733,N_4342,N_4123);
nand U4734 (N_4734,N_4032,N_4364);
nand U4735 (N_4735,N_4065,N_4310);
nand U4736 (N_4736,N_4069,N_4270);
and U4737 (N_4737,N_4207,N_4334);
or U4738 (N_4738,N_4389,N_4186);
or U4739 (N_4739,N_4161,N_4038);
nor U4740 (N_4740,N_4160,N_4347);
or U4741 (N_4741,N_4008,N_4366);
nor U4742 (N_4742,N_4010,N_4245);
nor U4743 (N_4743,N_4201,N_4161);
xnor U4744 (N_4744,N_4329,N_4041);
nand U4745 (N_4745,N_4314,N_4095);
and U4746 (N_4746,N_4100,N_4181);
or U4747 (N_4747,N_4306,N_4365);
nand U4748 (N_4748,N_4349,N_4026);
nor U4749 (N_4749,N_4119,N_4084);
nand U4750 (N_4750,N_4125,N_4397);
xnor U4751 (N_4751,N_4339,N_4036);
and U4752 (N_4752,N_4266,N_4208);
or U4753 (N_4753,N_4366,N_4147);
xor U4754 (N_4754,N_4199,N_4323);
and U4755 (N_4755,N_4343,N_4105);
and U4756 (N_4756,N_4371,N_4182);
or U4757 (N_4757,N_4135,N_4343);
and U4758 (N_4758,N_4179,N_4023);
nor U4759 (N_4759,N_4065,N_4316);
xnor U4760 (N_4760,N_4083,N_4133);
nor U4761 (N_4761,N_4008,N_4132);
or U4762 (N_4762,N_4181,N_4317);
xor U4763 (N_4763,N_4053,N_4077);
xor U4764 (N_4764,N_4280,N_4192);
nor U4765 (N_4765,N_4118,N_4314);
xor U4766 (N_4766,N_4398,N_4328);
nor U4767 (N_4767,N_4212,N_4233);
or U4768 (N_4768,N_4239,N_4397);
nand U4769 (N_4769,N_4201,N_4373);
and U4770 (N_4770,N_4339,N_4237);
nor U4771 (N_4771,N_4261,N_4097);
nand U4772 (N_4772,N_4121,N_4397);
and U4773 (N_4773,N_4370,N_4000);
nor U4774 (N_4774,N_4194,N_4117);
nand U4775 (N_4775,N_4394,N_4072);
or U4776 (N_4776,N_4354,N_4193);
nand U4777 (N_4777,N_4384,N_4098);
or U4778 (N_4778,N_4150,N_4329);
nor U4779 (N_4779,N_4076,N_4253);
or U4780 (N_4780,N_4070,N_4162);
and U4781 (N_4781,N_4238,N_4260);
nand U4782 (N_4782,N_4045,N_4119);
xnor U4783 (N_4783,N_4243,N_4357);
nor U4784 (N_4784,N_4368,N_4253);
or U4785 (N_4785,N_4131,N_4078);
xor U4786 (N_4786,N_4116,N_4317);
xnor U4787 (N_4787,N_4369,N_4106);
xnor U4788 (N_4788,N_4192,N_4343);
nor U4789 (N_4789,N_4196,N_4040);
and U4790 (N_4790,N_4072,N_4159);
and U4791 (N_4791,N_4302,N_4318);
xnor U4792 (N_4792,N_4172,N_4246);
xnor U4793 (N_4793,N_4124,N_4275);
xnor U4794 (N_4794,N_4089,N_4236);
and U4795 (N_4795,N_4250,N_4203);
nor U4796 (N_4796,N_4223,N_4093);
or U4797 (N_4797,N_4395,N_4055);
nor U4798 (N_4798,N_4184,N_4399);
or U4799 (N_4799,N_4194,N_4219);
nor U4800 (N_4800,N_4631,N_4736);
nor U4801 (N_4801,N_4774,N_4595);
and U4802 (N_4802,N_4478,N_4436);
nor U4803 (N_4803,N_4666,N_4675);
nand U4804 (N_4804,N_4641,N_4657);
and U4805 (N_4805,N_4614,N_4670);
nand U4806 (N_4806,N_4501,N_4743);
xor U4807 (N_4807,N_4459,N_4739);
nor U4808 (N_4808,N_4645,N_4734);
and U4809 (N_4809,N_4552,N_4699);
nand U4810 (N_4810,N_4655,N_4713);
nor U4811 (N_4811,N_4785,N_4747);
or U4812 (N_4812,N_4454,N_4742);
nor U4813 (N_4813,N_4504,N_4402);
nand U4814 (N_4814,N_4708,N_4538);
nand U4815 (N_4815,N_4542,N_4619);
or U4816 (N_4816,N_4681,N_4450);
and U4817 (N_4817,N_4517,N_4585);
xor U4818 (N_4818,N_4591,N_4669);
and U4819 (N_4819,N_4559,N_4745);
nand U4820 (N_4820,N_4607,N_4465);
xnor U4821 (N_4821,N_4626,N_4502);
xnor U4822 (N_4822,N_4579,N_4405);
xor U4823 (N_4823,N_4461,N_4409);
and U4824 (N_4824,N_4594,N_4404);
nor U4825 (N_4825,N_4612,N_4788);
xor U4826 (N_4826,N_4428,N_4432);
nor U4827 (N_4827,N_4578,N_4593);
or U4828 (N_4828,N_4440,N_4470);
nand U4829 (N_4829,N_4768,N_4627);
xor U4830 (N_4830,N_4413,N_4705);
xor U4831 (N_4831,N_4427,N_4541);
xnor U4832 (N_4832,N_4716,N_4714);
or U4833 (N_4833,N_4582,N_4475);
and U4834 (N_4834,N_4799,N_4407);
nor U4835 (N_4835,N_4639,N_4796);
xnor U4836 (N_4836,N_4483,N_4602);
or U4837 (N_4837,N_4457,N_4656);
nand U4838 (N_4838,N_4629,N_4625);
and U4839 (N_4839,N_4782,N_4507);
and U4840 (N_4840,N_4481,N_4786);
and U4841 (N_4841,N_4644,N_4773);
nand U4842 (N_4842,N_4726,N_4537);
or U4843 (N_4843,N_4671,N_4635);
xnor U4844 (N_4844,N_4509,N_4587);
nor U4845 (N_4845,N_4697,N_4623);
xnor U4846 (N_4846,N_4676,N_4425);
nand U4847 (N_4847,N_4487,N_4590);
nand U4848 (N_4848,N_4609,N_4673);
nor U4849 (N_4849,N_4679,N_4511);
nand U4850 (N_4850,N_4456,N_4685);
or U4851 (N_4851,N_4752,N_4581);
nand U4852 (N_4852,N_4599,N_4558);
nand U4853 (N_4853,N_4779,N_4632);
xnor U4854 (N_4854,N_4452,N_4760);
nor U4855 (N_4855,N_4534,N_4571);
and U4856 (N_4856,N_4680,N_4777);
and U4857 (N_4857,N_4667,N_4648);
nor U4858 (N_4858,N_4674,N_4664);
xnor U4859 (N_4859,N_4691,N_4683);
nand U4860 (N_4860,N_4439,N_4492);
nand U4861 (N_4861,N_4488,N_4567);
and U4862 (N_4862,N_4763,N_4496);
nand U4863 (N_4863,N_4493,N_4416);
nand U4864 (N_4864,N_4575,N_4446);
xor U4865 (N_4865,N_4408,N_4431);
nor U4866 (N_4866,N_4729,N_4503);
and U4867 (N_4867,N_4702,N_4566);
and U4868 (N_4868,N_4784,N_4577);
xnor U4869 (N_4869,N_4555,N_4433);
and U4870 (N_4870,N_4663,N_4758);
nand U4871 (N_4871,N_4617,N_4518);
or U4872 (N_4872,N_4410,N_4678);
nand U4873 (N_4873,N_4560,N_4471);
nand U4874 (N_4874,N_4530,N_4448);
xor U4875 (N_4875,N_4548,N_4622);
nand U4876 (N_4876,N_4480,N_4414);
nor U4877 (N_4877,N_4430,N_4766);
nor U4878 (N_4878,N_4717,N_4624);
nor U4879 (N_4879,N_4564,N_4418);
and U4880 (N_4880,N_4419,N_4565);
nand U4881 (N_4881,N_4715,N_4464);
nor U4882 (N_4882,N_4574,N_4449);
nand U4883 (N_4883,N_4740,N_4539);
nor U4884 (N_4884,N_4514,N_4444);
xor U4885 (N_4885,N_4458,N_4570);
and U4886 (N_4886,N_4651,N_4688);
and U4887 (N_4887,N_4479,N_4435);
xnor U4888 (N_4888,N_4605,N_4649);
and U4889 (N_4889,N_4469,N_4654);
xor U4890 (N_4890,N_4700,N_4429);
xnor U4891 (N_4891,N_4776,N_4755);
and U4892 (N_4892,N_4535,N_4415);
or U4893 (N_4893,N_4462,N_4672);
nand U4894 (N_4894,N_4698,N_4762);
nand U4895 (N_4895,N_4422,N_4725);
or U4896 (N_4896,N_4484,N_4721);
nand U4897 (N_4897,N_4783,N_4753);
nor U4898 (N_4898,N_4772,N_4723);
nor U4899 (N_4899,N_4746,N_4621);
or U4900 (N_4900,N_4598,N_4600);
or U4901 (N_4901,N_4618,N_4549);
xor U4902 (N_4902,N_4434,N_4490);
xnor U4903 (N_4903,N_4665,N_4642);
and U4904 (N_4904,N_4767,N_4769);
xor U4905 (N_4905,N_4401,N_4491);
nand U4906 (N_4906,N_4728,N_4573);
xnor U4907 (N_4907,N_4513,N_4426);
or U4908 (N_4908,N_4506,N_4797);
and U4909 (N_4909,N_4677,N_4524);
and U4910 (N_4910,N_4532,N_4695);
nor U4911 (N_4911,N_4443,N_4712);
nor U4912 (N_4912,N_4731,N_4580);
or U4913 (N_4913,N_4778,N_4550);
or U4914 (N_4914,N_4437,N_4525);
and U4915 (N_4915,N_4749,N_4756);
nand U4916 (N_4916,N_4790,N_4597);
xor U4917 (N_4917,N_4711,N_4730);
or U4918 (N_4918,N_4424,N_4472);
or U4919 (N_4919,N_4562,N_4720);
nand U4920 (N_4920,N_4761,N_4494);
and U4921 (N_4921,N_4604,N_4710);
nor U4922 (N_4922,N_4610,N_4466);
nand U4923 (N_4923,N_4658,N_4704);
nor U4924 (N_4924,N_4554,N_4781);
nor U4925 (N_4925,N_4596,N_4719);
nor U4926 (N_4926,N_4576,N_4601);
nor U4927 (N_4927,N_4653,N_4613);
or U4928 (N_4928,N_4727,N_4545);
or U4929 (N_4929,N_4637,N_4467);
nor U4930 (N_4930,N_4588,N_4460);
or U4931 (N_4931,N_4592,N_4792);
nor U4932 (N_4932,N_4531,N_4659);
xor U4933 (N_4933,N_4751,N_4793);
nand U4934 (N_4934,N_4724,N_4586);
nor U4935 (N_4935,N_4606,N_4476);
xnor U4936 (N_4936,N_4445,N_4505);
nand U4937 (N_4937,N_4500,N_4709);
or U4938 (N_4938,N_4744,N_4640);
or U4939 (N_4939,N_4764,N_4489);
or U4940 (N_4940,N_4696,N_4608);
nor U4941 (N_4941,N_4474,N_4741);
nor U4942 (N_4942,N_4738,N_4557);
and U4943 (N_4943,N_4718,N_4692);
nor U4944 (N_4944,N_4423,N_4633);
and U4945 (N_4945,N_4543,N_4668);
xor U4946 (N_4946,N_4643,N_4522);
or U4947 (N_4947,N_4703,N_4701);
and U4948 (N_4948,N_4690,N_4789);
nor U4949 (N_4949,N_4661,N_4498);
and U4950 (N_4950,N_4463,N_4447);
or U4951 (N_4951,N_4561,N_4516);
nand U4952 (N_4952,N_4400,N_4519);
nand U4953 (N_4953,N_4536,N_4551);
nand U4954 (N_4954,N_4750,N_4438);
nand U4955 (N_4955,N_4455,N_4453);
and U4956 (N_4956,N_4482,N_4693);
nand U4957 (N_4957,N_4497,N_4411);
nand U4958 (N_4958,N_4528,N_4611);
nand U4959 (N_4959,N_4652,N_4794);
and U4960 (N_4960,N_4647,N_4634);
xor U4961 (N_4961,N_4529,N_4508);
nand U4962 (N_4962,N_4630,N_4616);
or U4963 (N_4963,N_4737,N_4689);
nor U4964 (N_4964,N_4420,N_4795);
and U4965 (N_4965,N_4620,N_4406);
nor U4966 (N_4966,N_4775,N_4540);
or U4967 (N_4967,N_4707,N_4572);
xnor U4968 (N_4968,N_4547,N_4770);
nand U4969 (N_4969,N_4527,N_4722);
xnor U4970 (N_4970,N_4636,N_4735);
xor U4971 (N_4971,N_4510,N_4798);
and U4972 (N_4972,N_4546,N_4486);
and U4973 (N_4973,N_4477,N_4583);
xor U4974 (N_4974,N_4628,N_4417);
or U4975 (N_4975,N_4473,N_4421);
nand U4976 (N_4976,N_4733,N_4650);
nor U4977 (N_4977,N_4441,N_4694);
nor U4978 (N_4978,N_4780,N_4589);
and U4979 (N_4979,N_4638,N_4512);
xor U4980 (N_4980,N_4544,N_4660);
and U4981 (N_4981,N_4771,N_4686);
or U4982 (N_4982,N_4646,N_4748);
nor U4983 (N_4983,N_4759,N_4568);
nand U4984 (N_4984,N_4556,N_4403);
nor U4985 (N_4985,N_4451,N_4754);
or U4986 (N_4986,N_4533,N_4787);
or U4987 (N_4987,N_4682,N_4526);
or U4988 (N_4988,N_4523,N_4553);
nor U4989 (N_4989,N_4791,N_4521);
xnor U4990 (N_4990,N_4468,N_4687);
xor U4991 (N_4991,N_4615,N_4603);
nand U4992 (N_4992,N_4520,N_4584);
nor U4993 (N_4993,N_4495,N_4412);
and U4994 (N_4994,N_4757,N_4499);
or U4995 (N_4995,N_4706,N_4732);
nand U4996 (N_4996,N_4563,N_4442);
nand U4997 (N_4997,N_4515,N_4765);
nand U4998 (N_4998,N_4485,N_4684);
xor U4999 (N_4999,N_4662,N_4569);
xnor U5000 (N_5000,N_4781,N_4471);
nand U5001 (N_5001,N_4586,N_4650);
nor U5002 (N_5002,N_4571,N_4626);
nor U5003 (N_5003,N_4637,N_4619);
xor U5004 (N_5004,N_4782,N_4680);
or U5005 (N_5005,N_4544,N_4691);
xnor U5006 (N_5006,N_4555,N_4584);
or U5007 (N_5007,N_4791,N_4588);
or U5008 (N_5008,N_4554,N_4763);
nand U5009 (N_5009,N_4511,N_4519);
or U5010 (N_5010,N_4411,N_4737);
nand U5011 (N_5011,N_4515,N_4542);
xor U5012 (N_5012,N_4612,N_4697);
nor U5013 (N_5013,N_4700,N_4706);
and U5014 (N_5014,N_4781,N_4473);
nor U5015 (N_5015,N_4670,N_4718);
xor U5016 (N_5016,N_4735,N_4531);
nor U5017 (N_5017,N_4432,N_4642);
or U5018 (N_5018,N_4499,N_4416);
and U5019 (N_5019,N_4754,N_4569);
nand U5020 (N_5020,N_4513,N_4652);
xor U5021 (N_5021,N_4498,N_4753);
or U5022 (N_5022,N_4796,N_4625);
and U5023 (N_5023,N_4508,N_4428);
or U5024 (N_5024,N_4435,N_4641);
nor U5025 (N_5025,N_4696,N_4749);
nand U5026 (N_5026,N_4677,N_4583);
or U5027 (N_5027,N_4450,N_4632);
nand U5028 (N_5028,N_4771,N_4630);
nand U5029 (N_5029,N_4404,N_4615);
nand U5030 (N_5030,N_4590,N_4463);
nand U5031 (N_5031,N_4440,N_4655);
and U5032 (N_5032,N_4604,N_4590);
nand U5033 (N_5033,N_4485,N_4659);
or U5034 (N_5034,N_4493,N_4536);
and U5035 (N_5035,N_4666,N_4776);
nor U5036 (N_5036,N_4775,N_4403);
nor U5037 (N_5037,N_4464,N_4559);
and U5038 (N_5038,N_4429,N_4524);
nor U5039 (N_5039,N_4690,N_4733);
nand U5040 (N_5040,N_4761,N_4496);
nor U5041 (N_5041,N_4574,N_4707);
nand U5042 (N_5042,N_4577,N_4497);
and U5043 (N_5043,N_4697,N_4421);
xnor U5044 (N_5044,N_4670,N_4492);
xnor U5045 (N_5045,N_4706,N_4537);
xor U5046 (N_5046,N_4637,N_4772);
xor U5047 (N_5047,N_4692,N_4751);
nor U5048 (N_5048,N_4436,N_4784);
nand U5049 (N_5049,N_4590,N_4473);
xor U5050 (N_5050,N_4726,N_4588);
and U5051 (N_5051,N_4576,N_4672);
xor U5052 (N_5052,N_4666,N_4543);
or U5053 (N_5053,N_4707,N_4466);
nand U5054 (N_5054,N_4556,N_4563);
nand U5055 (N_5055,N_4739,N_4775);
and U5056 (N_5056,N_4588,N_4692);
xnor U5057 (N_5057,N_4485,N_4755);
and U5058 (N_5058,N_4702,N_4595);
nand U5059 (N_5059,N_4689,N_4463);
nor U5060 (N_5060,N_4530,N_4433);
xor U5061 (N_5061,N_4427,N_4477);
nor U5062 (N_5062,N_4783,N_4627);
nor U5063 (N_5063,N_4636,N_4633);
or U5064 (N_5064,N_4558,N_4670);
nand U5065 (N_5065,N_4692,N_4791);
xnor U5066 (N_5066,N_4613,N_4494);
nor U5067 (N_5067,N_4573,N_4766);
xor U5068 (N_5068,N_4666,N_4563);
nor U5069 (N_5069,N_4632,N_4788);
and U5070 (N_5070,N_4451,N_4529);
and U5071 (N_5071,N_4796,N_4516);
and U5072 (N_5072,N_4610,N_4413);
nand U5073 (N_5073,N_4618,N_4467);
xnor U5074 (N_5074,N_4736,N_4495);
and U5075 (N_5075,N_4602,N_4678);
and U5076 (N_5076,N_4632,N_4427);
and U5077 (N_5077,N_4759,N_4688);
nor U5078 (N_5078,N_4423,N_4694);
xor U5079 (N_5079,N_4690,N_4426);
nand U5080 (N_5080,N_4468,N_4420);
nor U5081 (N_5081,N_4457,N_4465);
nor U5082 (N_5082,N_4565,N_4469);
nand U5083 (N_5083,N_4525,N_4467);
and U5084 (N_5084,N_4712,N_4643);
or U5085 (N_5085,N_4509,N_4472);
nand U5086 (N_5086,N_4475,N_4443);
or U5087 (N_5087,N_4432,N_4544);
and U5088 (N_5088,N_4466,N_4475);
or U5089 (N_5089,N_4400,N_4451);
and U5090 (N_5090,N_4506,N_4718);
nand U5091 (N_5091,N_4415,N_4787);
or U5092 (N_5092,N_4776,N_4432);
and U5093 (N_5093,N_4578,N_4580);
or U5094 (N_5094,N_4605,N_4485);
nor U5095 (N_5095,N_4765,N_4691);
xnor U5096 (N_5096,N_4479,N_4784);
and U5097 (N_5097,N_4684,N_4720);
and U5098 (N_5098,N_4650,N_4500);
nand U5099 (N_5099,N_4494,N_4543);
nor U5100 (N_5100,N_4507,N_4656);
nor U5101 (N_5101,N_4740,N_4691);
xor U5102 (N_5102,N_4645,N_4400);
xor U5103 (N_5103,N_4662,N_4650);
nor U5104 (N_5104,N_4504,N_4526);
nand U5105 (N_5105,N_4657,N_4610);
xor U5106 (N_5106,N_4664,N_4594);
nor U5107 (N_5107,N_4731,N_4426);
xnor U5108 (N_5108,N_4776,N_4698);
or U5109 (N_5109,N_4452,N_4547);
or U5110 (N_5110,N_4724,N_4512);
nor U5111 (N_5111,N_4572,N_4657);
nand U5112 (N_5112,N_4766,N_4743);
nor U5113 (N_5113,N_4429,N_4691);
or U5114 (N_5114,N_4568,N_4463);
nand U5115 (N_5115,N_4595,N_4697);
and U5116 (N_5116,N_4529,N_4751);
or U5117 (N_5117,N_4568,N_4763);
nor U5118 (N_5118,N_4525,N_4549);
or U5119 (N_5119,N_4440,N_4554);
or U5120 (N_5120,N_4540,N_4667);
nor U5121 (N_5121,N_4599,N_4574);
nand U5122 (N_5122,N_4787,N_4783);
and U5123 (N_5123,N_4453,N_4407);
nand U5124 (N_5124,N_4716,N_4598);
or U5125 (N_5125,N_4656,N_4658);
xnor U5126 (N_5126,N_4569,N_4416);
xor U5127 (N_5127,N_4485,N_4771);
and U5128 (N_5128,N_4581,N_4600);
nor U5129 (N_5129,N_4549,N_4533);
and U5130 (N_5130,N_4747,N_4468);
nand U5131 (N_5131,N_4451,N_4602);
xnor U5132 (N_5132,N_4656,N_4722);
xnor U5133 (N_5133,N_4527,N_4550);
xnor U5134 (N_5134,N_4700,N_4760);
nand U5135 (N_5135,N_4581,N_4420);
or U5136 (N_5136,N_4465,N_4785);
xnor U5137 (N_5137,N_4543,N_4588);
nand U5138 (N_5138,N_4445,N_4430);
nand U5139 (N_5139,N_4537,N_4590);
nand U5140 (N_5140,N_4747,N_4770);
and U5141 (N_5141,N_4470,N_4786);
or U5142 (N_5142,N_4795,N_4608);
xnor U5143 (N_5143,N_4699,N_4472);
nor U5144 (N_5144,N_4688,N_4761);
nand U5145 (N_5145,N_4754,N_4418);
nand U5146 (N_5146,N_4699,N_4765);
and U5147 (N_5147,N_4593,N_4602);
or U5148 (N_5148,N_4516,N_4461);
nor U5149 (N_5149,N_4575,N_4751);
and U5150 (N_5150,N_4650,N_4744);
nor U5151 (N_5151,N_4455,N_4409);
xor U5152 (N_5152,N_4456,N_4735);
and U5153 (N_5153,N_4754,N_4555);
or U5154 (N_5154,N_4658,N_4663);
nand U5155 (N_5155,N_4665,N_4674);
nor U5156 (N_5156,N_4725,N_4652);
nor U5157 (N_5157,N_4563,N_4497);
nand U5158 (N_5158,N_4651,N_4505);
nand U5159 (N_5159,N_4446,N_4678);
and U5160 (N_5160,N_4451,N_4485);
or U5161 (N_5161,N_4719,N_4742);
or U5162 (N_5162,N_4429,N_4609);
xor U5163 (N_5163,N_4608,N_4732);
and U5164 (N_5164,N_4591,N_4798);
nor U5165 (N_5165,N_4756,N_4643);
or U5166 (N_5166,N_4739,N_4490);
and U5167 (N_5167,N_4598,N_4710);
xnor U5168 (N_5168,N_4521,N_4594);
nor U5169 (N_5169,N_4736,N_4681);
or U5170 (N_5170,N_4657,N_4745);
and U5171 (N_5171,N_4728,N_4441);
nor U5172 (N_5172,N_4421,N_4635);
nor U5173 (N_5173,N_4572,N_4633);
and U5174 (N_5174,N_4689,N_4550);
nor U5175 (N_5175,N_4673,N_4695);
xor U5176 (N_5176,N_4548,N_4455);
and U5177 (N_5177,N_4782,N_4626);
or U5178 (N_5178,N_4697,N_4683);
nor U5179 (N_5179,N_4604,N_4739);
and U5180 (N_5180,N_4646,N_4475);
xor U5181 (N_5181,N_4592,N_4474);
and U5182 (N_5182,N_4470,N_4703);
and U5183 (N_5183,N_4513,N_4681);
and U5184 (N_5184,N_4473,N_4544);
nor U5185 (N_5185,N_4792,N_4551);
xnor U5186 (N_5186,N_4529,N_4411);
or U5187 (N_5187,N_4727,N_4683);
nand U5188 (N_5188,N_4627,N_4690);
xnor U5189 (N_5189,N_4619,N_4462);
nand U5190 (N_5190,N_4678,N_4786);
nor U5191 (N_5191,N_4637,N_4402);
xor U5192 (N_5192,N_4576,N_4494);
nor U5193 (N_5193,N_4773,N_4714);
xor U5194 (N_5194,N_4516,N_4680);
or U5195 (N_5195,N_4769,N_4751);
nand U5196 (N_5196,N_4465,N_4642);
nand U5197 (N_5197,N_4406,N_4767);
or U5198 (N_5198,N_4614,N_4445);
or U5199 (N_5199,N_4638,N_4439);
nor U5200 (N_5200,N_4982,N_4901);
xor U5201 (N_5201,N_5128,N_5117);
xor U5202 (N_5202,N_4929,N_4971);
and U5203 (N_5203,N_4874,N_4962);
and U5204 (N_5204,N_4868,N_5172);
nand U5205 (N_5205,N_4927,N_4914);
nand U5206 (N_5206,N_5163,N_4871);
or U5207 (N_5207,N_4854,N_4824);
nor U5208 (N_5208,N_5045,N_5090);
nor U5209 (N_5209,N_4875,N_5111);
and U5210 (N_5210,N_5006,N_5134);
xnor U5211 (N_5211,N_4813,N_4973);
xor U5212 (N_5212,N_5061,N_4975);
and U5213 (N_5213,N_4947,N_5144);
nand U5214 (N_5214,N_4888,N_5124);
xnor U5215 (N_5215,N_5156,N_4828);
xor U5216 (N_5216,N_4839,N_4832);
xnor U5217 (N_5217,N_4864,N_4990);
xor U5218 (N_5218,N_5030,N_5119);
and U5219 (N_5219,N_4848,N_5048);
xor U5220 (N_5220,N_4918,N_4843);
or U5221 (N_5221,N_4998,N_5131);
or U5222 (N_5222,N_4847,N_5059);
xnor U5223 (N_5223,N_4806,N_4924);
or U5224 (N_5224,N_5114,N_5143);
or U5225 (N_5225,N_4899,N_5051);
or U5226 (N_5226,N_5009,N_4978);
or U5227 (N_5227,N_4861,N_5107);
xnor U5228 (N_5228,N_5181,N_4820);
nand U5229 (N_5229,N_5087,N_5094);
nand U5230 (N_5230,N_4849,N_5071);
xnor U5231 (N_5231,N_5150,N_4816);
xor U5232 (N_5232,N_4908,N_5195);
and U5233 (N_5233,N_5038,N_5164);
nand U5234 (N_5234,N_4801,N_5193);
xor U5235 (N_5235,N_4906,N_5154);
or U5236 (N_5236,N_5097,N_4993);
nor U5237 (N_5237,N_4943,N_4844);
or U5238 (N_5238,N_5069,N_4877);
and U5239 (N_5239,N_4881,N_5004);
xor U5240 (N_5240,N_5192,N_5166);
or U5241 (N_5241,N_5060,N_5028);
nor U5242 (N_5242,N_5159,N_4919);
and U5243 (N_5243,N_4822,N_5112);
nor U5244 (N_5244,N_4926,N_4841);
and U5245 (N_5245,N_5186,N_4850);
or U5246 (N_5246,N_4840,N_4934);
or U5247 (N_5247,N_5039,N_5089);
nor U5248 (N_5248,N_5176,N_4895);
nand U5249 (N_5249,N_4903,N_5135);
nand U5250 (N_5250,N_4956,N_4931);
xor U5251 (N_5251,N_5158,N_5019);
xnor U5252 (N_5252,N_5033,N_5093);
and U5253 (N_5253,N_4967,N_4838);
xor U5254 (N_5254,N_4987,N_4862);
nor U5255 (N_5255,N_5018,N_4831);
and U5256 (N_5256,N_5024,N_5070);
and U5257 (N_5257,N_4885,N_4856);
nand U5258 (N_5258,N_4916,N_5102);
or U5259 (N_5259,N_4949,N_4858);
nor U5260 (N_5260,N_4823,N_4898);
xor U5261 (N_5261,N_5005,N_4890);
and U5262 (N_5262,N_5072,N_4970);
or U5263 (N_5263,N_4827,N_4939);
xor U5264 (N_5264,N_5113,N_5196);
xnor U5265 (N_5265,N_4977,N_4857);
xor U5266 (N_5266,N_4957,N_4866);
xnor U5267 (N_5267,N_5095,N_4936);
nor U5268 (N_5268,N_4966,N_4997);
nand U5269 (N_5269,N_5189,N_5041);
nor U5270 (N_5270,N_5153,N_5013);
nand U5271 (N_5271,N_4892,N_4860);
and U5272 (N_5272,N_4963,N_5098);
and U5273 (N_5273,N_4902,N_5180);
nor U5274 (N_5274,N_5050,N_5110);
nor U5275 (N_5275,N_5141,N_5055);
nand U5276 (N_5276,N_4933,N_5105);
nor U5277 (N_5277,N_4870,N_4894);
nand U5278 (N_5278,N_4955,N_5199);
or U5279 (N_5279,N_4979,N_5000);
xnor U5280 (N_5280,N_4986,N_5007);
nor U5281 (N_5281,N_4923,N_4938);
xnor U5282 (N_5282,N_4921,N_4922);
xnor U5283 (N_5283,N_5037,N_4859);
and U5284 (N_5284,N_4964,N_5091);
and U5285 (N_5285,N_5052,N_5025);
nor U5286 (N_5286,N_5032,N_5167);
or U5287 (N_5287,N_4804,N_5122);
or U5288 (N_5288,N_5003,N_5015);
nand U5289 (N_5289,N_4985,N_4909);
xor U5290 (N_5290,N_5140,N_5026);
xor U5291 (N_5291,N_5047,N_4992);
and U5292 (N_5292,N_4837,N_4989);
nor U5293 (N_5293,N_4876,N_4833);
nor U5294 (N_5294,N_5121,N_4836);
nor U5295 (N_5295,N_4818,N_5165);
nand U5296 (N_5296,N_4910,N_5155);
or U5297 (N_5297,N_5147,N_4920);
xnor U5298 (N_5298,N_4878,N_5130);
and U5299 (N_5299,N_4995,N_4805);
or U5300 (N_5300,N_5044,N_4951);
or U5301 (N_5301,N_5099,N_4851);
xor U5302 (N_5302,N_5146,N_5109);
or U5303 (N_5303,N_4960,N_4965);
nor U5304 (N_5304,N_4981,N_4915);
and U5305 (N_5305,N_4800,N_5001);
or U5306 (N_5306,N_5085,N_4983);
nand U5307 (N_5307,N_5139,N_4814);
xnor U5308 (N_5308,N_4991,N_4867);
xnor U5309 (N_5309,N_4879,N_4897);
xnor U5310 (N_5310,N_5088,N_5101);
xnor U5311 (N_5311,N_5075,N_4980);
and U5312 (N_5312,N_5178,N_5017);
nor U5313 (N_5313,N_4807,N_5132);
nor U5314 (N_5314,N_5062,N_4930);
and U5315 (N_5315,N_5184,N_5142);
and U5316 (N_5316,N_5022,N_4900);
xnor U5317 (N_5317,N_4912,N_5068);
or U5318 (N_5318,N_4935,N_5149);
or U5319 (N_5319,N_4953,N_5057);
and U5320 (N_5320,N_4948,N_5034);
nand U5321 (N_5321,N_5125,N_5187);
and U5322 (N_5322,N_5151,N_4809);
or U5323 (N_5323,N_5067,N_5104);
nand U5324 (N_5324,N_4817,N_5073);
nand U5325 (N_5325,N_5120,N_4887);
or U5326 (N_5326,N_5191,N_4996);
and U5327 (N_5327,N_5171,N_4976);
nand U5328 (N_5328,N_4893,N_5058);
or U5329 (N_5329,N_5138,N_4937);
nand U5330 (N_5330,N_4855,N_5157);
xor U5331 (N_5331,N_4869,N_5198);
nor U5332 (N_5332,N_4826,N_4958);
xnor U5333 (N_5333,N_4944,N_4819);
nand U5334 (N_5334,N_5115,N_5152);
nand U5335 (N_5335,N_4803,N_5076);
nand U5336 (N_5336,N_4917,N_5065);
xor U5337 (N_5337,N_5148,N_4907);
and U5338 (N_5338,N_4972,N_4846);
or U5339 (N_5339,N_5096,N_5123);
and U5340 (N_5340,N_4815,N_4911);
xnor U5341 (N_5341,N_5127,N_4974);
nor U5342 (N_5342,N_4886,N_4946);
xnor U5343 (N_5343,N_5043,N_5053);
nand U5344 (N_5344,N_4942,N_4852);
nand U5345 (N_5345,N_4825,N_5197);
nor U5346 (N_5346,N_4896,N_4845);
nand U5347 (N_5347,N_4835,N_5188);
nand U5348 (N_5348,N_4940,N_5092);
nor U5349 (N_5349,N_5129,N_4821);
nor U5350 (N_5350,N_4884,N_4811);
nand U5351 (N_5351,N_4952,N_5194);
and U5352 (N_5352,N_5012,N_5086);
xor U5353 (N_5353,N_4999,N_5027);
or U5354 (N_5354,N_4810,N_5020);
xnor U5355 (N_5355,N_5066,N_4863);
or U5356 (N_5356,N_5078,N_5031);
nor U5357 (N_5357,N_5046,N_5162);
nor U5358 (N_5358,N_4968,N_5023);
xor U5359 (N_5359,N_5168,N_5080);
nand U5360 (N_5360,N_5161,N_5002);
and U5361 (N_5361,N_4988,N_4880);
and U5362 (N_5362,N_5082,N_5016);
xor U5363 (N_5363,N_4945,N_4812);
and U5364 (N_5364,N_4842,N_4872);
and U5365 (N_5365,N_4853,N_5040);
and U5366 (N_5366,N_5049,N_5064);
and U5367 (N_5367,N_5084,N_4891);
and U5368 (N_5368,N_5174,N_5083);
and U5369 (N_5369,N_5056,N_4873);
xnor U5370 (N_5370,N_5175,N_4925);
xor U5371 (N_5371,N_5035,N_5126);
and U5372 (N_5372,N_4959,N_5008);
or U5373 (N_5373,N_5042,N_4932);
or U5374 (N_5374,N_4984,N_5137);
nand U5375 (N_5375,N_5183,N_5182);
or U5376 (N_5376,N_5106,N_5173);
nor U5377 (N_5377,N_4834,N_5179);
nand U5378 (N_5378,N_4830,N_4950);
and U5379 (N_5379,N_4941,N_4969);
nor U5380 (N_5380,N_5108,N_5021);
and U5381 (N_5381,N_4802,N_4808);
nor U5382 (N_5382,N_5054,N_5074);
xor U5383 (N_5383,N_4913,N_4889);
xnor U5384 (N_5384,N_5116,N_4865);
nand U5385 (N_5385,N_4928,N_5079);
and U5386 (N_5386,N_4883,N_5118);
nor U5387 (N_5387,N_5077,N_5100);
nor U5388 (N_5388,N_5011,N_5036);
xnor U5389 (N_5389,N_5169,N_4882);
nand U5390 (N_5390,N_4954,N_5160);
xnor U5391 (N_5391,N_5136,N_5185);
nor U5392 (N_5392,N_5010,N_5081);
and U5393 (N_5393,N_4994,N_5029);
xnor U5394 (N_5394,N_4829,N_5103);
and U5395 (N_5395,N_5145,N_5190);
nor U5396 (N_5396,N_5063,N_4904);
xnor U5397 (N_5397,N_4905,N_5133);
xor U5398 (N_5398,N_5177,N_5014);
nor U5399 (N_5399,N_5170,N_4961);
nand U5400 (N_5400,N_5060,N_5168);
nand U5401 (N_5401,N_5050,N_4819);
or U5402 (N_5402,N_4874,N_5031);
nor U5403 (N_5403,N_4978,N_4852);
nand U5404 (N_5404,N_5024,N_4803);
nand U5405 (N_5405,N_5086,N_5190);
nand U5406 (N_5406,N_4804,N_4997);
nor U5407 (N_5407,N_5197,N_4861);
and U5408 (N_5408,N_4857,N_5126);
and U5409 (N_5409,N_4975,N_4928);
nor U5410 (N_5410,N_4868,N_5111);
nor U5411 (N_5411,N_5105,N_5116);
xnor U5412 (N_5412,N_5093,N_4928);
nand U5413 (N_5413,N_5085,N_5098);
xnor U5414 (N_5414,N_4853,N_5130);
nand U5415 (N_5415,N_5189,N_5128);
nor U5416 (N_5416,N_5119,N_5153);
and U5417 (N_5417,N_4858,N_4906);
and U5418 (N_5418,N_4926,N_5100);
nor U5419 (N_5419,N_4997,N_5110);
xnor U5420 (N_5420,N_5190,N_5109);
nand U5421 (N_5421,N_5100,N_4902);
or U5422 (N_5422,N_4825,N_5156);
xor U5423 (N_5423,N_4995,N_5139);
and U5424 (N_5424,N_5067,N_4819);
nand U5425 (N_5425,N_5037,N_5146);
or U5426 (N_5426,N_5046,N_5188);
xor U5427 (N_5427,N_5137,N_4817);
nand U5428 (N_5428,N_4973,N_5078);
or U5429 (N_5429,N_4820,N_5164);
nand U5430 (N_5430,N_5118,N_4901);
and U5431 (N_5431,N_4904,N_4902);
xnor U5432 (N_5432,N_4851,N_4813);
xor U5433 (N_5433,N_4922,N_4956);
and U5434 (N_5434,N_4817,N_5042);
nand U5435 (N_5435,N_4837,N_5016);
nor U5436 (N_5436,N_4920,N_5078);
xor U5437 (N_5437,N_5141,N_5020);
and U5438 (N_5438,N_4862,N_4917);
and U5439 (N_5439,N_4895,N_5084);
nand U5440 (N_5440,N_5041,N_5154);
nor U5441 (N_5441,N_4948,N_4919);
and U5442 (N_5442,N_4837,N_5098);
nor U5443 (N_5443,N_4857,N_4950);
nand U5444 (N_5444,N_4923,N_5083);
nand U5445 (N_5445,N_5026,N_5046);
and U5446 (N_5446,N_5014,N_5147);
or U5447 (N_5447,N_4813,N_4890);
and U5448 (N_5448,N_4800,N_5070);
xnor U5449 (N_5449,N_5177,N_4863);
and U5450 (N_5450,N_4986,N_5133);
nand U5451 (N_5451,N_5128,N_5154);
xnor U5452 (N_5452,N_4970,N_4816);
and U5453 (N_5453,N_5042,N_4946);
nand U5454 (N_5454,N_4832,N_5028);
nor U5455 (N_5455,N_5059,N_5013);
and U5456 (N_5456,N_4913,N_4851);
nor U5457 (N_5457,N_4995,N_4830);
and U5458 (N_5458,N_4973,N_5136);
or U5459 (N_5459,N_5005,N_4829);
and U5460 (N_5460,N_4953,N_5015);
and U5461 (N_5461,N_4838,N_4959);
and U5462 (N_5462,N_5193,N_5013);
nor U5463 (N_5463,N_5020,N_5138);
xor U5464 (N_5464,N_4849,N_4823);
or U5465 (N_5465,N_4931,N_4876);
xor U5466 (N_5466,N_4818,N_5093);
or U5467 (N_5467,N_5196,N_5002);
nand U5468 (N_5468,N_4965,N_5129);
nor U5469 (N_5469,N_4857,N_5163);
or U5470 (N_5470,N_4960,N_4968);
and U5471 (N_5471,N_4812,N_4955);
or U5472 (N_5472,N_5103,N_4877);
nor U5473 (N_5473,N_5042,N_4963);
nand U5474 (N_5474,N_5150,N_5107);
nor U5475 (N_5475,N_4964,N_4887);
or U5476 (N_5476,N_4905,N_4991);
nand U5477 (N_5477,N_4950,N_4982);
or U5478 (N_5478,N_4970,N_5116);
nor U5479 (N_5479,N_5124,N_4884);
or U5480 (N_5480,N_5145,N_5165);
or U5481 (N_5481,N_4882,N_5164);
nand U5482 (N_5482,N_4919,N_5120);
nor U5483 (N_5483,N_4917,N_4888);
nor U5484 (N_5484,N_4879,N_5157);
and U5485 (N_5485,N_5123,N_4809);
and U5486 (N_5486,N_4991,N_4955);
nand U5487 (N_5487,N_5057,N_4835);
xor U5488 (N_5488,N_4866,N_4923);
nand U5489 (N_5489,N_5160,N_4970);
and U5490 (N_5490,N_4996,N_5064);
nor U5491 (N_5491,N_5102,N_4967);
nor U5492 (N_5492,N_5011,N_4830);
nor U5493 (N_5493,N_5056,N_4900);
or U5494 (N_5494,N_4879,N_4995);
nand U5495 (N_5495,N_5082,N_5093);
nand U5496 (N_5496,N_5112,N_4947);
or U5497 (N_5497,N_5181,N_5127);
and U5498 (N_5498,N_5166,N_4958);
nand U5499 (N_5499,N_5106,N_4826);
nand U5500 (N_5500,N_4838,N_5158);
xnor U5501 (N_5501,N_5033,N_4830);
nand U5502 (N_5502,N_4989,N_5095);
and U5503 (N_5503,N_4883,N_5042);
nand U5504 (N_5504,N_5154,N_5038);
xnor U5505 (N_5505,N_4859,N_5117);
and U5506 (N_5506,N_4868,N_5048);
and U5507 (N_5507,N_4925,N_5024);
nor U5508 (N_5508,N_4884,N_5065);
nand U5509 (N_5509,N_4899,N_4985);
nor U5510 (N_5510,N_5104,N_4975);
nor U5511 (N_5511,N_5138,N_5140);
and U5512 (N_5512,N_4802,N_5011);
and U5513 (N_5513,N_5196,N_4966);
and U5514 (N_5514,N_4978,N_5015);
and U5515 (N_5515,N_4946,N_4968);
xnor U5516 (N_5516,N_5106,N_5036);
nor U5517 (N_5517,N_4841,N_5082);
nor U5518 (N_5518,N_5177,N_4817);
nand U5519 (N_5519,N_5077,N_4848);
nand U5520 (N_5520,N_4953,N_4873);
and U5521 (N_5521,N_5137,N_5149);
nor U5522 (N_5522,N_4975,N_5041);
and U5523 (N_5523,N_4913,N_5147);
xor U5524 (N_5524,N_5029,N_4821);
nor U5525 (N_5525,N_5193,N_4908);
nand U5526 (N_5526,N_4964,N_4951);
nor U5527 (N_5527,N_4938,N_4952);
nand U5528 (N_5528,N_4810,N_5098);
nor U5529 (N_5529,N_5190,N_5106);
nand U5530 (N_5530,N_4911,N_4977);
or U5531 (N_5531,N_4937,N_5128);
xor U5532 (N_5532,N_5199,N_5089);
xor U5533 (N_5533,N_4892,N_4879);
or U5534 (N_5534,N_4952,N_5186);
and U5535 (N_5535,N_4815,N_4955);
nor U5536 (N_5536,N_4978,N_4976);
nand U5537 (N_5537,N_4934,N_5134);
nand U5538 (N_5538,N_4909,N_5118);
xor U5539 (N_5539,N_5160,N_4900);
nor U5540 (N_5540,N_4847,N_5117);
nor U5541 (N_5541,N_4846,N_4931);
xor U5542 (N_5542,N_4943,N_4974);
and U5543 (N_5543,N_5137,N_5138);
xnor U5544 (N_5544,N_4833,N_5044);
xor U5545 (N_5545,N_4895,N_4851);
xnor U5546 (N_5546,N_4910,N_5125);
or U5547 (N_5547,N_4924,N_4859);
nor U5548 (N_5548,N_4838,N_5087);
xnor U5549 (N_5549,N_5047,N_4897);
or U5550 (N_5550,N_5129,N_5048);
xnor U5551 (N_5551,N_4919,N_5156);
nor U5552 (N_5552,N_4845,N_4864);
nor U5553 (N_5553,N_4991,N_5020);
or U5554 (N_5554,N_5181,N_4947);
xor U5555 (N_5555,N_4905,N_4995);
and U5556 (N_5556,N_5044,N_5062);
or U5557 (N_5557,N_4908,N_4850);
and U5558 (N_5558,N_4848,N_5126);
xnor U5559 (N_5559,N_5064,N_5081);
xnor U5560 (N_5560,N_5143,N_4827);
xor U5561 (N_5561,N_4902,N_5185);
xor U5562 (N_5562,N_4977,N_5195);
nor U5563 (N_5563,N_4936,N_5147);
and U5564 (N_5564,N_4826,N_4923);
nor U5565 (N_5565,N_5088,N_4842);
xor U5566 (N_5566,N_5035,N_5095);
xnor U5567 (N_5567,N_4873,N_5122);
or U5568 (N_5568,N_5149,N_4895);
and U5569 (N_5569,N_5060,N_4860);
nand U5570 (N_5570,N_5162,N_4944);
nand U5571 (N_5571,N_4883,N_4927);
xor U5572 (N_5572,N_4936,N_4851);
xnor U5573 (N_5573,N_5097,N_5133);
nor U5574 (N_5574,N_4846,N_5107);
nor U5575 (N_5575,N_4921,N_4882);
nor U5576 (N_5576,N_5044,N_4905);
nor U5577 (N_5577,N_4895,N_4993);
nor U5578 (N_5578,N_4916,N_4835);
xnor U5579 (N_5579,N_4978,N_4818);
xnor U5580 (N_5580,N_5178,N_5001);
nand U5581 (N_5581,N_5188,N_4923);
nand U5582 (N_5582,N_4816,N_4812);
xnor U5583 (N_5583,N_5086,N_4978);
nor U5584 (N_5584,N_4937,N_5099);
or U5585 (N_5585,N_5133,N_5101);
or U5586 (N_5586,N_4889,N_4899);
nor U5587 (N_5587,N_5107,N_5013);
xor U5588 (N_5588,N_5026,N_5011);
nor U5589 (N_5589,N_4981,N_5176);
or U5590 (N_5590,N_4924,N_5009);
nand U5591 (N_5591,N_5057,N_4954);
or U5592 (N_5592,N_5087,N_4849);
xor U5593 (N_5593,N_4801,N_4889);
xnor U5594 (N_5594,N_4867,N_4910);
nand U5595 (N_5595,N_4900,N_5018);
or U5596 (N_5596,N_4957,N_5121);
nor U5597 (N_5597,N_4987,N_5117);
or U5598 (N_5598,N_5022,N_4919);
nand U5599 (N_5599,N_4873,N_5184);
nor U5600 (N_5600,N_5343,N_5401);
and U5601 (N_5601,N_5422,N_5397);
nand U5602 (N_5602,N_5202,N_5566);
and U5603 (N_5603,N_5411,N_5584);
and U5604 (N_5604,N_5517,N_5449);
xnor U5605 (N_5605,N_5344,N_5567);
and U5606 (N_5606,N_5231,N_5406);
and U5607 (N_5607,N_5587,N_5501);
nand U5608 (N_5608,N_5282,N_5267);
nor U5609 (N_5609,N_5529,N_5573);
and U5610 (N_5610,N_5513,N_5433);
xor U5611 (N_5611,N_5580,N_5516);
nor U5612 (N_5612,N_5214,N_5360);
nand U5613 (N_5613,N_5218,N_5375);
xor U5614 (N_5614,N_5346,N_5519);
nand U5615 (N_5615,N_5296,N_5475);
nor U5616 (N_5616,N_5301,N_5207);
xnor U5617 (N_5617,N_5380,N_5465);
nor U5618 (N_5618,N_5310,N_5549);
or U5619 (N_5619,N_5277,N_5377);
nand U5620 (N_5620,N_5498,N_5261);
and U5621 (N_5621,N_5209,N_5398);
xnor U5622 (N_5622,N_5395,N_5404);
or U5623 (N_5623,N_5376,N_5252);
nor U5624 (N_5624,N_5553,N_5279);
nand U5625 (N_5625,N_5420,N_5438);
xor U5626 (N_5626,N_5414,N_5291);
nor U5627 (N_5627,N_5226,N_5505);
nand U5628 (N_5628,N_5251,N_5457);
or U5629 (N_5629,N_5281,N_5421);
or U5630 (N_5630,N_5366,N_5405);
and U5631 (N_5631,N_5307,N_5211);
nand U5632 (N_5632,N_5562,N_5456);
nor U5633 (N_5633,N_5364,N_5309);
or U5634 (N_5634,N_5381,N_5382);
or U5635 (N_5635,N_5256,N_5490);
and U5636 (N_5636,N_5290,N_5353);
or U5637 (N_5637,N_5544,N_5551);
or U5638 (N_5638,N_5329,N_5531);
and U5639 (N_5639,N_5315,N_5536);
nor U5640 (N_5640,N_5459,N_5439);
nand U5641 (N_5641,N_5356,N_5265);
nand U5642 (N_5642,N_5337,N_5451);
xnor U5643 (N_5643,N_5582,N_5471);
nor U5644 (N_5644,N_5208,N_5488);
and U5645 (N_5645,N_5571,N_5273);
and U5646 (N_5646,N_5317,N_5470);
xnor U5647 (N_5647,N_5493,N_5204);
or U5648 (N_5648,N_5468,N_5502);
and U5649 (N_5649,N_5403,N_5423);
or U5650 (N_5650,N_5259,N_5585);
nand U5651 (N_5651,N_5407,N_5312);
nor U5652 (N_5652,N_5563,N_5595);
nor U5653 (N_5653,N_5324,N_5286);
or U5654 (N_5654,N_5472,N_5320);
nor U5655 (N_5655,N_5328,N_5210);
xnor U5656 (N_5656,N_5283,N_5316);
xnor U5657 (N_5657,N_5213,N_5447);
nand U5658 (N_5658,N_5539,N_5358);
and U5659 (N_5659,N_5245,N_5576);
nor U5660 (N_5660,N_5284,N_5361);
xor U5661 (N_5661,N_5460,N_5349);
and U5662 (N_5662,N_5367,N_5327);
nor U5663 (N_5663,N_5200,N_5342);
or U5664 (N_5664,N_5441,N_5446);
nand U5665 (N_5665,N_5492,N_5295);
nand U5666 (N_5666,N_5430,N_5491);
or U5667 (N_5667,N_5368,N_5285);
xor U5668 (N_5668,N_5354,N_5436);
and U5669 (N_5669,N_5257,N_5432);
nor U5670 (N_5670,N_5485,N_5378);
and U5671 (N_5671,N_5321,N_5527);
or U5672 (N_5672,N_5541,N_5311);
nor U5673 (N_5673,N_5463,N_5201);
nand U5674 (N_5674,N_5522,N_5440);
or U5675 (N_5675,N_5340,N_5363);
nand U5676 (N_5676,N_5483,N_5511);
or U5677 (N_5677,N_5552,N_5396);
or U5678 (N_5678,N_5355,N_5258);
nor U5679 (N_5679,N_5305,N_5274);
nor U5680 (N_5680,N_5219,N_5480);
xor U5681 (N_5681,N_5287,N_5383);
and U5682 (N_5682,N_5484,N_5275);
nand U5683 (N_5683,N_5350,N_5462);
xnor U5684 (N_5684,N_5238,N_5509);
nand U5685 (N_5685,N_5525,N_5532);
nand U5686 (N_5686,N_5220,N_5297);
nand U5687 (N_5687,N_5540,N_5336);
xor U5688 (N_5688,N_5535,N_5523);
xnor U5689 (N_5689,N_5215,N_5565);
or U5690 (N_5690,N_5444,N_5384);
nand U5691 (N_5691,N_5306,N_5270);
or U5692 (N_5692,N_5599,N_5334);
and U5693 (N_5693,N_5443,N_5326);
nand U5694 (N_5694,N_5554,N_5589);
nand U5695 (N_5695,N_5391,N_5216);
nand U5696 (N_5696,N_5335,N_5507);
xor U5697 (N_5697,N_5419,N_5524);
nand U5698 (N_5698,N_5481,N_5469);
xor U5699 (N_5699,N_5276,N_5300);
nand U5700 (N_5700,N_5400,N_5445);
nand U5701 (N_5701,N_5597,N_5359);
nor U5702 (N_5702,N_5564,N_5203);
or U5703 (N_5703,N_5388,N_5427);
nand U5704 (N_5704,N_5234,N_5244);
nor U5705 (N_5705,N_5435,N_5534);
nand U5706 (N_5706,N_5303,N_5240);
nand U5707 (N_5707,N_5393,N_5345);
xor U5708 (N_5708,N_5370,N_5586);
nor U5709 (N_5709,N_5508,N_5530);
nor U5710 (N_5710,N_5572,N_5431);
xor U5711 (N_5711,N_5561,N_5548);
or U5712 (N_5712,N_5598,N_5250);
nor U5713 (N_5713,N_5387,N_5246);
and U5714 (N_5714,N_5494,N_5331);
or U5715 (N_5715,N_5547,N_5222);
nand U5716 (N_5716,N_5372,N_5302);
nand U5717 (N_5717,N_5537,N_5241);
nand U5718 (N_5718,N_5578,N_5255);
and U5719 (N_5719,N_5520,N_5409);
nand U5720 (N_5720,N_5521,N_5233);
nand U5721 (N_5721,N_5374,N_5487);
nor U5722 (N_5722,N_5596,N_5591);
nor U5723 (N_5723,N_5365,N_5289);
or U5724 (N_5724,N_5533,N_5308);
and U5725 (N_5725,N_5338,N_5394);
nand U5726 (N_5726,N_5538,N_5332);
and U5727 (N_5727,N_5357,N_5410);
nor U5728 (N_5728,N_5212,N_5236);
xnor U5729 (N_5729,N_5514,N_5559);
nor U5730 (N_5730,N_5434,N_5272);
nor U5731 (N_5731,N_5323,N_5280);
nor U5732 (N_5732,N_5504,N_5497);
or U5733 (N_5733,N_5243,N_5428);
and U5734 (N_5734,N_5228,N_5249);
nand U5735 (N_5735,N_5319,N_5474);
and U5736 (N_5736,N_5512,N_5515);
or U5737 (N_5737,N_5330,N_5489);
and U5738 (N_5738,N_5402,N_5556);
or U5739 (N_5739,N_5528,N_5299);
nor U5740 (N_5740,N_5424,N_5333);
nand U5741 (N_5741,N_5339,N_5399);
and U5742 (N_5742,N_5429,N_5466);
or U5743 (N_5743,N_5221,N_5503);
xor U5744 (N_5744,N_5313,N_5526);
nand U5745 (N_5745,N_5412,N_5304);
or U5746 (N_5746,N_5269,N_5314);
and U5747 (N_5747,N_5569,N_5351);
xor U5748 (N_5748,N_5450,N_5543);
nor U5749 (N_5749,N_5217,N_5482);
and U5750 (N_5750,N_5389,N_5206);
or U5751 (N_5751,N_5254,N_5477);
xnor U5752 (N_5752,N_5426,N_5278);
or U5753 (N_5753,N_5570,N_5479);
and U5754 (N_5754,N_5232,N_5293);
nand U5755 (N_5755,N_5464,N_5266);
or U5756 (N_5756,N_5542,N_5341);
nand U5757 (N_5757,N_5235,N_5593);
and U5758 (N_5758,N_5558,N_5292);
or U5759 (N_5759,N_5461,N_5448);
nand U5760 (N_5760,N_5557,N_5425);
nor U5761 (N_5761,N_5499,N_5574);
and U5762 (N_5762,N_5458,N_5506);
nand U5763 (N_5763,N_5486,N_5473);
nor U5764 (N_5764,N_5510,N_5237);
nand U5765 (N_5765,N_5590,N_5223);
nor U5766 (N_5766,N_5288,N_5294);
nor U5767 (N_5767,N_5348,N_5392);
xor U5768 (N_5768,N_5229,N_5362);
nand U5769 (N_5769,N_5577,N_5417);
xnor U5770 (N_5770,N_5253,N_5373);
or U5771 (N_5771,N_5416,N_5495);
and U5772 (N_5772,N_5518,N_5581);
xnor U5773 (N_5773,N_5453,N_5369);
xnor U5774 (N_5774,N_5545,N_5379);
and U5775 (N_5775,N_5476,N_5496);
or U5776 (N_5776,N_5271,N_5413);
nand U5777 (N_5777,N_5583,N_5262);
xnor U5778 (N_5778,N_5437,N_5478);
nor U5779 (N_5779,N_5371,N_5239);
nor U5780 (N_5780,N_5224,N_5352);
nand U5781 (N_5781,N_5452,N_5568);
or U5782 (N_5782,N_5268,N_5247);
and U5783 (N_5783,N_5579,N_5500);
and U5784 (N_5784,N_5594,N_5225);
xor U5785 (N_5785,N_5415,N_5325);
and U5786 (N_5786,N_5385,N_5260);
and U5787 (N_5787,N_5230,N_5546);
or U5788 (N_5788,N_5467,N_5205);
nor U5789 (N_5789,N_5386,N_5560);
xor U5790 (N_5790,N_5248,N_5347);
nand U5791 (N_5791,N_5550,N_5298);
and U5792 (N_5792,N_5454,N_5264);
nor U5793 (N_5793,N_5455,N_5418);
xor U5794 (N_5794,N_5227,N_5390);
and U5795 (N_5795,N_5442,N_5263);
nand U5796 (N_5796,N_5318,N_5322);
nor U5797 (N_5797,N_5408,N_5242);
or U5798 (N_5798,N_5575,N_5555);
nor U5799 (N_5799,N_5592,N_5588);
xnor U5800 (N_5800,N_5316,N_5229);
nor U5801 (N_5801,N_5258,N_5281);
xor U5802 (N_5802,N_5289,N_5542);
nand U5803 (N_5803,N_5460,N_5304);
nand U5804 (N_5804,N_5508,N_5262);
and U5805 (N_5805,N_5513,N_5478);
nand U5806 (N_5806,N_5330,N_5377);
nand U5807 (N_5807,N_5236,N_5537);
nand U5808 (N_5808,N_5462,N_5279);
nand U5809 (N_5809,N_5479,N_5236);
and U5810 (N_5810,N_5416,N_5286);
and U5811 (N_5811,N_5260,N_5583);
and U5812 (N_5812,N_5596,N_5561);
and U5813 (N_5813,N_5305,N_5465);
nand U5814 (N_5814,N_5253,N_5494);
xnor U5815 (N_5815,N_5328,N_5344);
xor U5816 (N_5816,N_5206,N_5486);
and U5817 (N_5817,N_5473,N_5421);
nand U5818 (N_5818,N_5377,N_5274);
nand U5819 (N_5819,N_5223,N_5243);
or U5820 (N_5820,N_5245,N_5416);
and U5821 (N_5821,N_5538,N_5284);
or U5822 (N_5822,N_5233,N_5327);
xor U5823 (N_5823,N_5543,N_5228);
nand U5824 (N_5824,N_5491,N_5493);
xor U5825 (N_5825,N_5593,N_5455);
xor U5826 (N_5826,N_5431,N_5493);
xor U5827 (N_5827,N_5256,N_5572);
or U5828 (N_5828,N_5568,N_5406);
and U5829 (N_5829,N_5229,N_5385);
and U5830 (N_5830,N_5558,N_5215);
and U5831 (N_5831,N_5314,N_5464);
nor U5832 (N_5832,N_5424,N_5204);
nand U5833 (N_5833,N_5598,N_5510);
or U5834 (N_5834,N_5523,N_5391);
or U5835 (N_5835,N_5552,N_5420);
or U5836 (N_5836,N_5477,N_5312);
nand U5837 (N_5837,N_5576,N_5300);
nand U5838 (N_5838,N_5572,N_5413);
xor U5839 (N_5839,N_5548,N_5571);
nor U5840 (N_5840,N_5235,N_5334);
nor U5841 (N_5841,N_5273,N_5378);
nor U5842 (N_5842,N_5543,N_5324);
nor U5843 (N_5843,N_5414,N_5418);
xnor U5844 (N_5844,N_5290,N_5333);
or U5845 (N_5845,N_5349,N_5207);
xnor U5846 (N_5846,N_5586,N_5469);
nor U5847 (N_5847,N_5431,N_5212);
or U5848 (N_5848,N_5506,N_5213);
nor U5849 (N_5849,N_5443,N_5421);
or U5850 (N_5850,N_5485,N_5233);
nor U5851 (N_5851,N_5335,N_5518);
xor U5852 (N_5852,N_5409,N_5427);
nand U5853 (N_5853,N_5315,N_5438);
and U5854 (N_5854,N_5476,N_5354);
nand U5855 (N_5855,N_5342,N_5337);
and U5856 (N_5856,N_5323,N_5201);
nor U5857 (N_5857,N_5420,N_5377);
or U5858 (N_5858,N_5518,N_5311);
nor U5859 (N_5859,N_5570,N_5443);
nor U5860 (N_5860,N_5287,N_5507);
nand U5861 (N_5861,N_5200,N_5313);
nor U5862 (N_5862,N_5507,N_5377);
nor U5863 (N_5863,N_5494,N_5434);
or U5864 (N_5864,N_5264,N_5361);
and U5865 (N_5865,N_5396,N_5495);
nand U5866 (N_5866,N_5508,N_5350);
and U5867 (N_5867,N_5539,N_5362);
or U5868 (N_5868,N_5362,N_5493);
nor U5869 (N_5869,N_5456,N_5275);
xnor U5870 (N_5870,N_5463,N_5518);
nor U5871 (N_5871,N_5518,N_5294);
and U5872 (N_5872,N_5316,N_5274);
and U5873 (N_5873,N_5599,N_5550);
xor U5874 (N_5874,N_5491,N_5409);
nor U5875 (N_5875,N_5284,N_5558);
xor U5876 (N_5876,N_5291,N_5440);
nand U5877 (N_5877,N_5367,N_5510);
xor U5878 (N_5878,N_5468,N_5363);
nand U5879 (N_5879,N_5326,N_5520);
and U5880 (N_5880,N_5587,N_5422);
nor U5881 (N_5881,N_5590,N_5460);
and U5882 (N_5882,N_5567,N_5495);
xnor U5883 (N_5883,N_5233,N_5205);
and U5884 (N_5884,N_5481,N_5571);
nor U5885 (N_5885,N_5399,N_5392);
xor U5886 (N_5886,N_5484,N_5466);
nor U5887 (N_5887,N_5530,N_5585);
and U5888 (N_5888,N_5291,N_5438);
nand U5889 (N_5889,N_5445,N_5462);
nor U5890 (N_5890,N_5458,N_5353);
or U5891 (N_5891,N_5326,N_5366);
xor U5892 (N_5892,N_5531,N_5369);
nor U5893 (N_5893,N_5433,N_5456);
and U5894 (N_5894,N_5408,N_5211);
nand U5895 (N_5895,N_5229,N_5205);
or U5896 (N_5896,N_5313,N_5367);
nor U5897 (N_5897,N_5504,N_5332);
nand U5898 (N_5898,N_5502,N_5312);
nor U5899 (N_5899,N_5431,N_5469);
and U5900 (N_5900,N_5461,N_5447);
xor U5901 (N_5901,N_5380,N_5508);
xnor U5902 (N_5902,N_5537,N_5237);
nand U5903 (N_5903,N_5503,N_5351);
xnor U5904 (N_5904,N_5242,N_5354);
or U5905 (N_5905,N_5405,N_5247);
xor U5906 (N_5906,N_5343,N_5248);
nor U5907 (N_5907,N_5403,N_5469);
or U5908 (N_5908,N_5512,N_5259);
nor U5909 (N_5909,N_5318,N_5543);
and U5910 (N_5910,N_5417,N_5555);
and U5911 (N_5911,N_5358,N_5232);
and U5912 (N_5912,N_5400,N_5237);
nand U5913 (N_5913,N_5583,N_5524);
and U5914 (N_5914,N_5274,N_5275);
nand U5915 (N_5915,N_5562,N_5237);
nand U5916 (N_5916,N_5392,N_5353);
nand U5917 (N_5917,N_5431,N_5583);
xor U5918 (N_5918,N_5577,N_5518);
nand U5919 (N_5919,N_5593,N_5397);
nor U5920 (N_5920,N_5490,N_5457);
xor U5921 (N_5921,N_5231,N_5599);
or U5922 (N_5922,N_5284,N_5248);
or U5923 (N_5923,N_5456,N_5450);
nand U5924 (N_5924,N_5384,N_5357);
xor U5925 (N_5925,N_5584,N_5320);
or U5926 (N_5926,N_5510,N_5503);
or U5927 (N_5927,N_5416,N_5270);
or U5928 (N_5928,N_5333,N_5543);
nor U5929 (N_5929,N_5497,N_5217);
or U5930 (N_5930,N_5443,N_5296);
nand U5931 (N_5931,N_5513,N_5423);
and U5932 (N_5932,N_5513,N_5598);
xor U5933 (N_5933,N_5331,N_5370);
and U5934 (N_5934,N_5587,N_5259);
and U5935 (N_5935,N_5213,N_5439);
xnor U5936 (N_5936,N_5396,N_5487);
nand U5937 (N_5937,N_5508,N_5295);
xor U5938 (N_5938,N_5360,N_5385);
nor U5939 (N_5939,N_5577,N_5223);
and U5940 (N_5940,N_5552,N_5324);
nor U5941 (N_5941,N_5333,N_5586);
nor U5942 (N_5942,N_5444,N_5251);
xor U5943 (N_5943,N_5210,N_5342);
nor U5944 (N_5944,N_5230,N_5237);
and U5945 (N_5945,N_5284,N_5439);
and U5946 (N_5946,N_5495,N_5393);
nor U5947 (N_5947,N_5425,N_5501);
xor U5948 (N_5948,N_5364,N_5255);
xor U5949 (N_5949,N_5265,N_5483);
and U5950 (N_5950,N_5497,N_5344);
nor U5951 (N_5951,N_5258,N_5362);
or U5952 (N_5952,N_5251,N_5337);
xor U5953 (N_5953,N_5253,N_5383);
xnor U5954 (N_5954,N_5409,N_5434);
and U5955 (N_5955,N_5506,N_5253);
nor U5956 (N_5956,N_5283,N_5497);
and U5957 (N_5957,N_5488,N_5235);
or U5958 (N_5958,N_5411,N_5536);
and U5959 (N_5959,N_5212,N_5338);
and U5960 (N_5960,N_5559,N_5208);
xor U5961 (N_5961,N_5453,N_5338);
xnor U5962 (N_5962,N_5474,N_5562);
xor U5963 (N_5963,N_5516,N_5473);
nor U5964 (N_5964,N_5521,N_5224);
nand U5965 (N_5965,N_5350,N_5355);
xnor U5966 (N_5966,N_5555,N_5271);
nor U5967 (N_5967,N_5309,N_5445);
and U5968 (N_5968,N_5532,N_5495);
and U5969 (N_5969,N_5299,N_5379);
and U5970 (N_5970,N_5307,N_5486);
xor U5971 (N_5971,N_5236,N_5372);
xnor U5972 (N_5972,N_5314,N_5466);
nand U5973 (N_5973,N_5282,N_5421);
and U5974 (N_5974,N_5259,N_5283);
or U5975 (N_5975,N_5336,N_5212);
or U5976 (N_5976,N_5560,N_5231);
and U5977 (N_5977,N_5517,N_5572);
xnor U5978 (N_5978,N_5277,N_5342);
and U5979 (N_5979,N_5554,N_5417);
and U5980 (N_5980,N_5341,N_5248);
nor U5981 (N_5981,N_5347,N_5213);
or U5982 (N_5982,N_5491,N_5466);
and U5983 (N_5983,N_5583,N_5567);
and U5984 (N_5984,N_5397,N_5549);
nor U5985 (N_5985,N_5315,N_5455);
xnor U5986 (N_5986,N_5585,N_5508);
nand U5987 (N_5987,N_5386,N_5381);
or U5988 (N_5988,N_5502,N_5226);
xor U5989 (N_5989,N_5331,N_5289);
nor U5990 (N_5990,N_5392,N_5536);
and U5991 (N_5991,N_5233,N_5559);
xor U5992 (N_5992,N_5389,N_5516);
nor U5993 (N_5993,N_5388,N_5206);
nand U5994 (N_5994,N_5234,N_5372);
or U5995 (N_5995,N_5385,N_5597);
xnor U5996 (N_5996,N_5234,N_5306);
nand U5997 (N_5997,N_5459,N_5417);
nand U5998 (N_5998,N_5484,N_5531);
nor U5999 (N_5999,N_5440,N_5537);
or U6000 (N_6000,N_5712,N_5642);
or U6001 (N_6001,N_5610,N_5802);
nor U6002 (N_6002,N_5664,N_5630);
nor U6003 (N_6003,N_5961,N_5612);
xnor U6004 (N_6004,N_5833,N_5732);
and U6005 (N_6005,N_5821,N_5853);
xnor U6006 (N_6006,N_5710,N_5753);
and U6007 (N_6007,N_5893,N_5764);
or U6008 (N_6008,N_5621,N_5625);
or U6009 (N_6009,N_5626,N_5771);
or U6010 (N_6010,N_5787,N_5840);
or U6011 (N_6011,N_5768,N_5872);
nor U6012 (N_6012,N_5613,N_5786);
or U6013 (N_6013,N_5982,N_5917);
or U6014 (N_6014,N_5865,N_5806);
nand U6015 (N_6015,N_5656,N_5719);
and U6016 (N_6016,N_5900,N_5862);
or U6017 (N_6017,N_5793,N_5720);
nor U6018 (N_6018,N_5682,N_5641);
xnor U6019 (N_6019,N_5636,N_5800);
nor U6020 (N_6020,N_5644,N_5733);
and U6021 (N_6021,N_5954,N_5678);
nand U6022 (N_6022,N_5690,N_5938);
xor U6023 (N_6023,N_5918,N_5637);
and U6024 (N_6024,N_5958,N_5974);
or U6025 (N_6025,N_5773,N_5639);
xnor U6026 (N_6026,N_5929,N_5699);
and U6027 (N_6027,N_5651,N_5850);
nor U6028 (N_6028,N_5646,N_5962);
nand U6029 (N_6029,N_5703,N_5859);
nor U6030 (N_6030,N_5640,N_5946);
nand U6031 (N_6031,N_5628,N_5908);
xor U6032 (N_6032,N_5913,N_5836);
xor U6033 (N_6033,N_5981,N_5987);
nand U6034 (N_6034,N_5686,N_5940);
and U6035 (N_6035,N_5658,N_5684);
or U6036 (N_6036,N_5835,N_5671);
and U6037 (N_6037,N_5889,N_5864);
and U6038 (N_6038,N_5968,N_5777);
and U6039 (N_6039,N_5881,N_5914);
nand U6040 (N_6040,N_5890,N_5711);
or U6041 (N_6041,N_5995,N_5925);
nand U6042 (N_6042,N_5746,N_5869);
nor U6043 (N_6043,N_5848,N_5619);
and U6044 (N_6044,N_5614,N_5805);
and U6045 (N_6045,N_5897,N_5822);
nor U6046 (N_6046,N_5886,N_5663);
and U6047 (N_6047,N_5604,N_5873);
nor U6048 (N_6048,N_5912,N_5676);
nand U6049 (N_6049,N_5696,N_5722);
xnor U6050 (N_6050,N_5863,N_5898);
or U6051 (N_6051,N_5951,N_5615);
xnor U6052 (N_6052,N_5706,N_5799);
and U6053 (N_6053,N_5718,N_5747);
nand U6054 (N_6054,N_5880,N_5724);
or U6055 (N_6055,N_5757,N_5774);
or U6056 (N_6056,N_5736,N_5755);
and U6057 (N_6057,N_5815,N_5823);
nor U6058 (N_6058,N_5643,N_5655);
or U6059 (N_6059,N_5980,N_5879);
nor U6060 (N_6060,N_5931,N_5708);
nor U6061 (N_6061,N_5989,N_5731);
or U6062 (N_6062,N_5607,N_5785);
nand U6063 (N_6063,N_5972,N_5947);
nand U6064 (N_6064,N_5854,N_5867);
and U6065 (N_6065,N_5677,N_5965);
nand U6066 (N_6066,N_5936,N_5996);
or U6067 (N_6067,N_5928,N_5804);
nand U6068 (N_6068,N_5910,N_5659);
and U6069 (N_6069,N_5971,N_5933);
and U6070 (N_6070,N_5691,N_5674);
nand U6071 (N_6071,N_5809,N_5741);
and U6072 (N_6072,N_5950,N_5838);
nor U6073 (N_6073,N_5895,N_5780);
nor U6074 (N_6074,N_5993,N_5675);
xor U6075 (N_6075,N_5909,N_5698);
nand U6076 (N_6076,N_5779,N_5681);
xor U6077 (N_6077,N_5679,N_5795);
nor U6078 (N_6078,N_5834,N_5846);
nor U6079 (N_6079,N_5858,N_5700);
or U6080 (N_6080,N_5990,N_5969);
or U6081 (N_6081,N_5784,N_5807);
or U6082 (N_6082,N_5662,N_5616);
nand U6083 (N_6083,N_5737,N_5645);
and U6084 (N_6084,N_5852,N_5666);
and U6085 (N_6085,N_5957,N_5824);
nor U6086 (N_6086,N_5670,N_5654);
nand U6087 (N_6087,N_5901,N_5716);
xnor U6088 (N_6088,N_5624,N_5728);
nor U6089 (N_6089,N_5622,N_5767);
and U6090 (N_6090,N_5752,N_5832);
and U6091 (N_6091,N_5683,N_5756);
and U6092 (N_6092,N_5647,N_5882);
xnor U6093 (N_6093,N_5668,N_5949);
nand U6094 (N_6094,N_5916,N_5794);
nor U6095 (N_6095,N_5808,N_5744);
or U6096 (N_6096,N_5892,N_5915);
and U6097 (N_6097,N_5966,N_5874);
nor U6098 (N_6098,N_5792,N_5934);
or U6099 (N_6099,N_5817,N_5932);
nor U6100 (N_6100,N_5760,N_5891);
or U6101 (N_6101,N_5870,N_5661);
nand U6102 (N_6102,N_5941,N_5725);
and U6103 (N_6103,N_5751,N_5721);
or U6104 (N_6104,N_5749,N_5829);
nand U6105 (N_6105,N_5798,N_5876);
nor U6106 (N_6106,N_5635,N_5960);
xor U6107 (N_6107,N_5772,N_5955);
nor U6108 (N_6108,N_5801,N_5887);
nand U6109 (N_6109,N_5944,N_5868);
nor U6110 (N_6110,N_5877,N_5902);
nor U6111 (N_6111,N_5937,N_5855);
nor U6112 (N_6112,N_5758,N_5715);
and U6113 (N_6113,N_5687,N_5945);
nand U6114 (N_6114,N_5992,N_5739);
and U6115 (N_6115,N_5866,N_5704);
nor U6116 (N_6116,N_5796,N_5707);
and U6117 (N_6117,N_5723,N_5906);
or U6118 (N_6118,N_5797,N_5692);
nor U6119 (N_6119,N_5790,N_5776);
or U6120 (N_6120,N_5783,N_5648);
or U6121 (N_6121,N_5841,N_5831);
nor U6122 (N_6122,N_5973,N_5611);
nand U6123 (N_6123,N_5618,N_5759);
xnor U6124 (N_6124,N_5782,N_5977);
or U6125 (N_6125,N_5942,N_5688);
nor U6126 (N_6126,N_5813,N_5921);
or U6127 (N_6127,N_5847,N_5632);
and U6128 (N_6128,N_5788,N_5979);
nor U6129 (N_6129,N_5861,N_5775);
or U6130 (N_6130,N_5726,N_5924);
xnor U6131 (N_6131,N_5789,N_5964);
xnor U6132 (N_6132,N_5629,N_5814);
or U6133 (N_6133,N_5871,N_5888);
xor U6134 (N_6134,N_5601,N_5754);
nand U6135 (N_6135,N_5602,N_5899);
and U6136 (N_6136,N_5903,N_5709);
nor U6137 (N_6137,N_5884,N_5907);
and U6138 (N_6138,N_5983,N_5763);
xor U6139 (N_6139,N_5830,N_5603);
nand U6140 (N_6140,N_5689,N_5600);
nand U6141 (N_6141,N_5702,N_5713);
nand U6142 (N_6142,N_5935,N_5761);
xor U6143 (N_6143,N_5812,N_5717);
or U6144 (N_6144,N_5894,N_5837);
and U6145 (N_6145,N_5939,N_5770);
and U6146 (N_6146,N_5740,N_5694);
and U6147 (N_6147,N_5652,N_5967);
or U6148 (N_6148,N_5672,N_5705);
xnor U6149 (N_6149,N_5693,N_5984);
nand U6150 (N_6150,N_5849,N_5927);
nor U6151 (N_6151,N_5999,N_5791);
or U6152 (N_6152,N_5742,N_5634);
and U6153 (N_6153,N_5926,N_5856);
or U6154 (N_6154,N_5669,N_5998);
or U6155 (N_6155,N_5997,N_5978);
nand U6156 (N_6156,N_5851,N_5943);
or U6157 (N_6157,N_5623,N_5839);
nand U6158 (N_6158,N_5673,N_5734);
xor U6159 (N_6159,N_5638,N_5631);
nand U6160 (N_6160,N_5762,N_5811);
nand U6161 (N_6161,N_5920,N_5714);
or U6162 (N_6162,N_5970,N_5665);
nand U6163 (N_6163,N_5956,N_5953);
nand U6164 (N_6164,N_5701,N_5653);
xnor U6165 (N_6165,N_5769,N_5857);
nand U6166 (N_6166,N_5609,N_5875);
xor U6167 (N_6167,N_5878,N_5743);
nor U6168 (N_6168,N_5991,N_5633);
nand U6169 (N_6169,N_5975,N_5826);
and U6170 (N_6170,N_5627,N_5781);
nand U6171 (N_6171,N_5766,N_5745);
and U6172 (N_6172,N_5985,N_5930);
or U6173 (N_6173,N_5994,N_5845);
nand U6174 (N_6174,N_5738,N_5919);
nand U6175 (N_6175,N_5986,N_5606);
and U6176 (N_6176,N_5843,N_5735);
and U6177 (N_6177,N_5608,N_5952);
nor U6178 (N_6178,N_5883,N_5605);
nor U6179 (N_6179,N_5765,N_5810);
and U6180 (N_6180,N_5860,N_5617);
xnor U6181 (N_6181,N_5650,N_5827);
xor U6182 (N_6182,N_5963,N_5695);
nand U6183 (N_6183,N_5828,N_5904);
nand U6184 (N_6184,N_5657,N_5685);
nand U6185 (N_6185,N_5748,N_5896);
and U6186 (N_6186,N_5727,N_5885);
nor U6187 (N_6187,N_5750,N_5842);
nand U6188 (N_6188,N_5697,N_5816);
nor U6189 (N_6189,N_5976,N_5730);
nand U6190 (N_6190,N_5778,N_5649);
or U6191 (N_6191,N_5819,N_5923);
nor U6192 (N_6192,N_5905,N_5680);
xor U6193 (N_6193,N_5667,N_5729);
nor U6194 (N_6194,N_5948,N_5660);
xnor U6195 (N_6195,N_5620,N_5820);
or U6196 (N_6196,N_5911,N_5959);
xnor U6197 (N_6197,N_5922,N_5825);
xor U6198 (N_6198,N_5818,N_5988);
nor U6199 (N_6199,N_5803,N_5844);
or U6200 (N_6200,N_5962,N_5637);
and U6201 (N_6201,N_5624,N_5631);
nand U6202 (N_6202,N_5966,N_5953);
and U6203 (N_6203,N_5676,N_5669);
nand U6204 (N_6204,N_5773,N_5720);
nor U6205 (N_6205,N_5858,N_5777);
nand U6206 (N_6206,N_5817,N_5860);
xor U6207 (N_6207,N_5793,N_5655);
or U6208 (N_6208,N_5833,N_5615);
nand U6209 (N_6209,N_5628,N_5742);
nand U6210 (N_6210,N_5924,N_5838);
xnor U6211 (N_6211,N_5814,N_5890);
nor U6212 (N_6212,N_5664,N_5657);
or U6213 (N_6213,N_5897,N_5771);
or U6214 (N_6214,N_5993,N_5861);
or U6215 (N_6215,N_5863,N_5973);
nand U6216 (N_6216,N_5837,N_5654);
and U6217 (N_6217,N_5902,N_5977);
or U6218 (N_6218,N_5897,N_5711);
nor U6219 (N_6219,N_5876,N_5834);
xor U6220 (N_6220,N_5690,N_5948);
nor U6221 (N_6221,N_5739,N_5913);
or U6222 (N_6222,N_5656,N_5677);
xor U6223 (N_6223,N_5726,N_5844);
and U6224 (N_6224,N_5663,N_5999);
xor U6225 (N_6225,N_5788,N_5775);
and U6226 (N_6226,N_5629,N_5654);
and U6227 (N_6227,N_5924,N_5600);
nor U6228 (N_6228,N_5839,N_5700);
or U6229 (N_6229,N_5983,N_5672);
xnor U6230 (N_6230,N_5722,N_5736);
xor U6231 (N_6231,N_5740,N_5853);
and U6232 (N_6232,N_5983,N_5836);
and U6233 (N_6233,N_5674,N_5938);
nand U6234 (N_6234,N_5712,N_5684);
or U6235 (N_6235,N_5933,N_5884);
nand U6236 (N_6236,N_5925,N_5764);
nand U6237 (N_6237,N_5783,N_5726);
nand U6238 (N_6238,N_5648,N_5923);
nor U6239 (N_6239,N_5860,N_5721);
or U6240 (N_6240,N_5760,N_5686);
nor U6241 (N_6241,N_5657,N_5993);
xor U6242 (N_6242,N_5799,N_5805);
xor U6243 (N_6243,N_5627,N_5977);
nor U6244 (N_6244,N_5736,N_5831);
or U6245 (N_6245,N_5835,N_5701);
nor U6246 (N_6246,N_5911,N_5746);
nand U6247 (N_6247,N_5961,N_5649);
or U6248 (N_6248,N_5818,N_5959);
and U6249 (N_6249,N_5679,N_5659);
nand U6250 (N_6250,N_5729,N_5735);
nor U6251 (N_6251,N_5851,N_5681);
or U6252 (N_6252,N_5698,N_5851);
nand U6253 (N_6253,N_5674,N_5809);
nand U6254 (N_6254,N_5809,N_5713);
and U6255 (N_6255,N_5800,N_5726);
or U6256 (N_6256,N_5880,N_5950);
nor U6257 (N_6257,N_5820,N_5931);
xnor U6258 (N_6258,N_5727,N_5636);
and U6259 (N_6259,N_5966,N_5960);
nor U6260 (N_6260,N_5697,N_5870);
or U6261 (N_6261,N_5979,N_5840);
xnor U6262 (N_6262,N_5811,N_5909);
xor U6263 (N_6263,N_5821,N_5809);
and U6264 (N_6264,N_5947,N_5671);
and U6265 (N_6265,N_5663,N_5725);
and U6266 (N_6266,N_5765,N_5661);
and U6267 (N_6267,N_5716,N_5695);
or U6268 (N_6268,N_5825,N_5772);
nand U6269 (N_6269,N_5888,N_5615);
nand U6270 (N_6270,N_5934,N_5707);
nor U6271 (N_6271,N_5874,N_5624);
nand U6272 (N_6272,N_5649,N_5973);
nor U6273 (N_6273,N_5632,N_5996);
nand U6274 (N_6274,N_5880,N_5949);
and U6275 (N_6275,N_5601,N_5996);
xnor U6276 (N_6276,N_5980,N_5974);
nand U6277 (N_6277,N_5656,N_5798);
or U6278 (N_6278,N_5665,N_5640);
nand U6279 (N_6279,N_5970,N_5827);
xor U6280 (N_6280,N_5907,N_5788);
or U6281 (N_6281,N_5843,N_5740);
or U6282 (N_6282,N_5607,N_5957);
xnor U6283 (N_6283,N_5917,N_5645);
or U6284 (N_6284,N_5879,N_5826);
nor U6285 (N_6285,N_5890,N_5654);
nand U6286 (N_6286,N_5825,N_5727);
nor U6287 (N_6287,N_5771,N_5641);
and U6288 (N_6288,N_5935,N_5815);
xor U6289 (N_6289,N_5975,N_5837);
nand U6290 (N_6290,N_5887,N_5935);
or U6291 (N_6291,N_5650,N_5966);
and U6292 (N_6292,N_5824,N_5638);
nand U6293 (N_6293,N_5853,N_5753);
or U6294 (N_6294,N_5760,N_5842);
or U6295 (N_6295,N_5852,N_5996);
or U6296 (N_6296,N_5964,N_5787);
or U6297 (N_6297,N_5982,N_5629);
or U6298 (N_6298,N_5784,N_5622);
nor U6299 (N_6299,N_5900,N_5689);
nand U6300 (N_6300,N_5925,N_5747);
nand U6301 (N_6301,N_5878,N_5943);
or U6302 (N_6302,N_5991,N_5947);
nor U6303 (N_6303,N_5654,N_5953);
and U6304 (N_6304,N_5732,N_5861);
or U6305 (N_6305,N_5927,N_5955);
and U6306 (N_6306,N_5818,N_5986);
nor U6307 (N_6307,N_5622,N_5615);
or U6308 (N_6308,N_5670,N_5617);
nand U6309 (N_6309,N_5639,N_5604);
nor U6310 (N_6310,N_5909,N_5641);
and U6311 (N_6311,N_5908,N_5636);
xnor U6312 (N_6312,N_5650,N_5805);
xor U6313 (N_6313,N_5922,N_5886);
and U6314 (N_6314,N_5916,N_5945);
xnor U6315 (N_6315,N_5744,N_5792);
xor U6316 (N_6316,N_5681,N_5796);
xnor U6317 (N_6317,N_5850,N_5868);
xor U6318 (N_6318,N_5602,N_5794);
and U6319 (N_6319,N_5758,N_5771);
nand U6320 (N_6320,N_5618,N_5608);
nand U6321 (N_6321,N_5872,N_5695);
xor U6322 (N_6322,N_5854,N_5851);
nand U6323 (N_6323,N_5973,N_5832);
or U6324 (N_6324,N_5925,N_5733);
xnor U6325 (N_6325,N_5928,N_5686);
nand U6326 (N_6326,N_5892,N_5894);
xor U6327 (N_6327,N_5691,N_5653);
nand U6328 (N_6328,N_5728,N_5606);
and U6329 (N_6329,N_5749,N_5689);
and U6330 (N_6330,N_5737,N_5646);
xor U6331 (N_6331,N_5825,N_5765);
nand U6332 (N_6332,N_5855,N_5736);
or U6333 (N_6333,N_5860,N_5877);
nor U6334 (N_6334,N_5948,N_5669);
and U6335 (N_6335,N_5765,N_5921);
nor U6336 (N_6336,N_5963,N_5730);
xor U6337 (N_6337,N_5600,N_5988);
nand U6338 (N_6338,N_5744,N_5963);
nor U6339 (N_6339,N_5768,N_5718);
and U6340 (N_6340,N_5643,N_5970);
xor U6341 (N_6341,N_5707,N_5767);
xor U6342 (N_6342,N_5919,N_5804);
nor U6343 (N_6343,N_5937,N_5971);
nor U6344 (N_6344,N_5777,N_5925);
or U6345 (N_6345,N_5783,N_5638);
or U6346 (N_6346,N_5713,N_5645);
or U6347 (N_6347,N_5692,N_5672);
and U6348 (N_6348,N_5826,N_5760);
or U6349 (N_6349,N_5698,N_5704);
and U6350 (N_6350,N_5940,N_5681);
and U6351 (N_6351,N_5869,N_5673);
nand U6352 (N_6352,N_5788,N_5616);
and U6353 (N_6353,N_5805,N_5740);
xnor U6354 (N_6354,N_5829,N_5876);
xnor U6355 (N_6355,N_5712,N_5627);
xnor U6356 (N_6356,N_5758,N_5788);
nand U6357 (N_6357,N_5787,N_5753);
xnor U6358 (N_6358,N_5666,N_5902);
nand U6359 (N_6359,N_5986,N_5854);
nand U6360 (N_6360,N_5660,N_5794);
or U6361 (N_6361,N_5869,N_5966);
nor U6362 (N_6362,N_5888,N_5889);
and U6363 (N_6363,N_5787,N_5739);
nor U6364 (N_6364,N_5646,N_5660);
or U6365 (N_6365,N_5740,N_5631);
or U6366 (N_6366,N_5742,N_5981);
and U6367 (N_6367,N_5772,N_5896);
or U6368 (N_6368,N_5805,N_5616);
and U6369 (N_6369,N_5707,N_5625);
nand U6370 (N_6370,N_5824,N_5605);
and U6371 (N_6371,N_5689,N_5848);
nand U6372 (N_6372,N_5606,N_5619);
xor U6373 (N_6373,N_5881,N_5721);
and U6374 (N_6374,N_5818,N_5797);
nor U6375 (N_6375,N_5769,N_5787);
nor U6376 (N_6376,N_5760,N_5681);
nor U6377 (N_6377,N_5972,N_5727);
or U6378 (N_6378,N_5853,N_5902);
nand U6379 (N_6379,N_5907,N_5880);
or U6380 (N_6380,N_5689,N_5966);
xor U6381 (N_6381,N_5915,N_5724);
nor U6382 (N_6382,N_5834,N_5623);
xor U6383 (N_6383,N_5848,N_5706);
or U6384 (N_6384,N_5682,N_5989);
or U6385 (N_6385,N_5897,N_5959);
and U6386 (N_6386,N_5748,N_5636);
nand U6387 (N_6387,N_5814,N_5855);
nor U6388 (N_6388,N_5885,N_5967);
xor U6389 (N_6389,N_5627,N_5973);
nand U6390 (N_6390,N_5772,N_5645);
nor U6391 (N_6391,N_5648,N_5968);
nor U6392 (N_6392,N_5670,N_5787);
nor U6393 (N_6393,N_5712,N_5934);
xnor U6394 (N_6394,N_5759,N_5797);
nor U6395 (N_6395,N_5955,N_5818);
nand U6396 (N_6396,N_5973,N_5810);
or U6397 (N_6397,N_5896,N_5875);
nor U6398 (N_6398,N_5718,N_5906);
and U6399 (N_6399,N_5915,N_5802);
nand U6400 (N_6400,N_6054,N_6387);
xor U6401 (N_6401,N_6229,N_6190);
and U6402 (N_6402,N_6294,N_6084);
nand U6403 (N_6403,N_6126,N_6311);
nand U6404 (N_6404,N_6373,N_6318);
xor U6405 (N_6405,N_6134,N_6013);
or U6406 (N_6406,N_6206,N_6297);
nor U6407 (N_6407,N_6191,N_6069);
nand U6408 (N_6408,N_6292,N_6181);
or U6409 (N_6409,N_6231,N_6299);
or U6410 (N_6410,N_6110,N_6383);
nand U6411 (N_6411,N_6379,N_6377);
or U6412 (N_6412,N_6378,N_6274);
nor U6413 (N_6413,N_6317,N_6083);
and U6414 (N_6414,N_6262,N_6359);
xnor U6415 (N_6415,N_6355,N_6173);
or U6416 (N_6416,N_6330,N_6144);
xor U6417 (N_6417,N_6205,N_6033);
or U6418 (N_6418,N_6275,N_6088);
or U6419 (N_6419,N_6321,N_6012);
xnor U6420 (N_6420,N_6128,N_6391);
xor U6421 (N_6421,N_6298,N_6167);
nand U6422 (N_6422,N_6019,N_6176);
xnor U6423 (N_6423,N_6165,N_6367);
xnor U6424 (N_6424,N_6296,N_6303);
and U6425 (N_6425,N_6150,N_6185);
nand U6426 (N_6426,N_6023,N_6301);
nand U6427 (N_6427,N_6120,N_6133);
nand U6428 (N_6428,N_6009,N_6123);
nand U6429 (N_6429,N_6241,N_6112);
and U6430 (N_6430,N_6052,N_6334);
nor U6431 (N_6431,N_6184,N_6148);
or U6432 (N_6432,N_6029,N_6001);
nor U6433 (N_6433,N_6041,N_6125);
xor U6434 (N_6434,N_6224,N_6008);
xor U6435 (N_6435,N_6356,N_6341);
nor U6436 (N_6436,N_6203,N_6364);
xnor U6437 (N_6437,N_6223,N_6073);
xor U6438 (N_6438,N_6220,N_6056);
and U6439 (N_6439,N_6360,N_6238);
and U6440 (N_6440,N_6113,N_6263);
or U6441 (N_6441,N_6328,N_6003);
xnor U6442 (N_6442,N_6159,N_6142);
or U6443 (N_6443,N_6219,N_6390);
xnor U6444 (N_6444,N_6157,N_6352);
and U6445 (N_6445,N_6246,N_6104);
nand U6446 (N_6446,N_6027,N_6258);
nand U6447 (N_6447,N_6198,N_6022);
and U6448 (N_6448,N_6040,N_6332);
and U6449 (N_6449,N_6090,N_6266);
nand U6450 (N_6450,N_6000,N_6077);
nor U6451 (N_6451,N_6339,N_6396);
or U6452 (N_6452,N_6154,N_6098);
and U6453 (N_6453,N_6018,N_6232);
or U6454 (N_6454,N_6047,N_6247);
xnor U6455 (N_6455,N_6172,N_6031);
nor U6456 (N_6456,N_6269,N_6228);
nand U6457 (N_6457,N_6058,N_6350);
nor U6458 (N_6458,N_6175,N_6323);
nor U6459 (N_6459,N_6064,N_6315);
and U6460 (N_6460,N_6314,N_6124);
or U6461 (N_6461,N_6143,N_6305);
nor U6462 (N_6462,N_6138,N_6192);
xor U6463 (N_6463,N_6014,N_6340);
and U6464 (N_6464,N_6074,N_6285);
xor U6465 (N_6465,N_6108,N_6200);
and U6466 (N_6466,N_6156,N_6271);
nand U6467 (N_6467,N_6394,N_6245);
or U6468 (N_6468,N_6240,N_6072);
xor U6469 (N_6469,N_6070,N_6049);
nand U6470 (N_6470,N_6147,N_6320);
xor U6471 (N_6471,N_6376,N_6280);
xor U6472 (N_6472,N_6213,N_6121);
xnor U6473 (N_6473,N_6208,N_6291);
and U6474 (N_6474,N_6392,N_6252);
or U6475 (N_6475,N_6371,N_6114);
xor U6476 (N_6476,N_6362,N_6264);
nand U6477 (N_6477,N_6358,N_6122);
nand U6478 (N_6478,N_6270,N_6044);
nor U6479 (N_6479,N_6107,N_6091);
and U6480 (N_6480,N_6267,N_6386);
or U6481 (N_6481,N_6046,N_6168);
nand U6482 (N_6482,N_6131,N_6368);
nor U6483 (N_6483,N_6024,N_6153);
xor U6484 (N_6484,N_6011,N_6006);
xnor U6485 (N_6485,N_6209,N_6326);
nor U6486 (N_6486,N_6227,N_6081);
nand U6487 (N_6487,N_6369,N_6366);
nand U6488 (N_6488,N_6349,N_6094);
nor U6489 (N_6489,N_6053,N_6163);
nand U6490 (N_6490,N_6319,N_6251);
and U6491 (N_6491,N_6365,N_6109);
or U6492 (N_6492,N_6076,N_6100);
and U6493 (N_6493,N_6132,N_6197);
or U6494 (N_6494,N_6034,N_6007);
xnor U6495 (N_6495,N_6374,N_6067);
or U6496 (N_6496,N_6199,N_6169);
or U6497 (N_6497,N_6370,N_6178);
and U6498 (N_6498,N_6177,N_6155);
and U6499 (N_6499,N_6233,N_6039);
nand U6500 (N_6500,N_6015,N_6017);
xnor U6501 (N_6501,N_6343,N_6038);
xnor U6502 (N_6502,N_6141,N_6093);
and U6503 (N_6503,N_6261,N_6204);
and U6504 (N_6504,N_6036,N_6244);
and U6505 (N_6505,N_6277,N_6381);
and U6506 (N_6506,N_6187,N_6331);
nand U6507 (N_6507,N_6080,N_6284);
nand U6508 (N_6508,N_6020,N_6145);
xor U6509 (N_6509,N_6353,N_6162);
nand U6510 (N_6510,N_6186,N_6062);
or U6511 (N_6511,N_6035,N_6086);
and U6512 (N_6512,N_6278,N_6057);
nor U6513 (N_6513,N_6136,N_6242);
or U6514 (N_6514,N_6119,N_6382);
and U6515 (N_6515,N_6043,N_6236);
nor U6516 (N_6516,N_6272,N_6324);
xnor U6517 (N_6517,N_6174,N_6068);
xor U6518 (N_6518,N_6243,N_6234);
nor U6519 (N_6519,N_6158,N_6268);
and U6520 (N_6520,N_6188,N_6254);
xor U6521 (N_6521,N_6050,N_6201);
nor U6522 (N_6522,N_6384,N_6361);
and U6523 (N_6523,N_6030,N_6097);
nand U6524 (N_6524,N_6065,N_6180);
nor U6525 (N_6525,N_6344,N_6265);
xnor U6526 (N_6526,N_6348,N_6214);
or U6527 (N_6527,N_6295,N_6127);
and U6528 (N_6528,N_6388,N_6004);
nand U6529 (N_6529,N_6071,N_6256);
and U6530 (N_6530,N_6286,N_6257);
or U6531 (N_6531,N_6102,N_6166);
nor U6532 (N_6532,N_6025,N_6316);
and U6533 (N_6533,N_6250,N_6021);
nand U6534 (N_6534,N_6078,N_6304);
and U6535 (N_6535,N_6363,N_6336);
or U6536 (N_6536,N_6397,N_6060);
or U6537 (N_6537,N_6276,N_6235);
and U6538 (N_6538,N_6079,N_6161);
or U6539 (N_6539,N_6273,N_6260);
xor U6540 (N_6540,N_6338,N_6389);
nand U6541 (N_6541,N_6116,N_6225);
xnor U6542 (N_6542,N_6327,N_6117);
nor U6543 (N_6543,N_6032,N_6005);
or U6544 (N_6544,N_6302,N_6310);
nor U6545 (N_6545,N_6335,N_6010);
nand U6546 (N_6546,N_6309,N_6230);
xor U6547 (N_6547,N_6095,N_6207);
and U6548 (N_6548,N_6048,N_6193);
or U6549 (N_6549,N_6002,N_6248);
nor U6550 (N_6550,N_6111,N_6026);
or U6551 (N_6551,N_6239,N_6137);
nor U6552 (N_6552,N_6259,N_6281);
or U6553 (N_6553,N_6152,N_6087);
or U6554 (N_6554,N_6151,N_6313);
and U6555 (N_6555,N_6346,N_6333);
xnor U6556 (N_6556,N_6082,N_6300);
xnor U6557 (N_6557,N_6115,N_6216);
nand U6558 (N_6558,N_6312,N_6101);
or U6559 (N_6559,N_6237,N_6255);
nand U6560 (N_6560,N_6182,N_6221);
and U6561 (N_6561,N_6282,N_6195);
nor U6562 (N_6562,N_6160,N_6249);
or U6563 (N_6563,N_6398,N_6211);
xnor U6564 (N_6564,N_6325,N_6253);
and U6565 (N_6565,N_6061,N_6194);
nor U6566 (N_6566,N_6045,N_6171);
nand U6567 (N_6567,N_6287,N_6105);
nand U6568 (N_6568,N_6329,N_6179);
nor U6569 (N_6569,N_6106,N_6308);
xor U6570 (N_6570,N_6037,N_6089);
nor U6571 (N_6571,N_6149,N_6202);
xor U6572 (N_6572,N_6393,N_6289);
xor U6573 (N_6573,N_6103,N_6075);
xnor U6574 (N_6574,N_6357,N_6130);
and U6575 (N_6575,N_6063,N_6099);
nor U6576 (N_6576,N_6354,N_6222);
or U6577 (N_6577,N_6347,N_6226);
xnor U6578 (N_6578,N_6375,N_6140);
nand U6579 (N_6579,N_6016,N_6096);
xor U6580 (N_6580,N_6399,N_6183);
nand U6581 (N_6581,N_6380,N_6042);
nand U6582 (N_6582,N_6164,N_6337);
xnor U6583 (N_6583,N_6170,N_6092);
and U6584 (N_6584,N_6215,N_6189);
nor U6585 (N_6585,N_6139,N_6293);
and U6586 (N_6586,N_6085,N_6283);
xor U6587 (N_6587,N_6051,N_6395);
or U6588 (N_6588,N_6196,N_6129);
xor U6589 (N_6589,N_6066,N_6217);
xnor U6590 (N_6590,N_6212,N_6118);
or U6591 (N_6591,N_6135,N_6385);
nor U6592 (N_6592,N_6028,N_6306);
xor U6593 (N_6593,N_6351,N_6307);
or U6594 (N_6594,N_6288,N_6342);
nor U6595 (N_6595,N_6290,N_6218);
xnor U6596 (N_6596,N_6146,N_6210);
and U6597 (N_6597,N_6322,N_6279);
or U6598 (N_6598,N_6372,N_6059);
or U6599 (N_6599,N_6055,N_6345);
and U6600 (N_6600,N_6073,N_6193);
and U6601 (N_6601,N_6053,N_6285);
nand U6602 (N_6602,N_6189,N_6168);
nor U6603 (N_6603,N_6383,N_6223);
or U6604 (N_6604,N_6142,N_6360);
and U6605 (N_6605,N_6353,N_6303);
or U6606 (N_6606,N_6245,N_6142);
xnor U6607 (N_6607,N_6101,N_6079);
and U6608 (N_6608,N_6310,N_6163);
or U6609 (N_6609,N_6073,N_6147);
and U6610 (N_6610,N_6183,N_6019);
and U6611 (N_6611,N_6144,N_6366);
xor U6612 (N_6612,N_6366,N_6345);
or U6613 (N_6613,N_6084,N_6232);
and U6614 (N_6614,N_6367,N_6029);
nand U6615 (N_6615,N_6107,N_6360);
xor U6616 (N_6616,N_6173,N_6031);
xor U6617 (N_6617,N_6043,N_6226);
or U6618 (N_6618,N_6196,N_6030);
or U6619 (N_6619,N_6232,N_6047);
or U6620 (N_6620,N_6135,N_6258);
and U6621 (N_6621,N_6065,N_6064);
xor U6622 (N_6622,N_6363,N_6394);
xor U6623 (N_6623,N_6150,N_6002);
and U6624 (N_6624,N_6302,N_6198);
nand U6625 (N_6625,N_6116,N_6089);
nand U6626 (N_6626,N_6146,N_6223);
xor U6627 (N_6627,N_6159,N_6125);
or U6628 (N_6628,N_6353,N_6193);
nand U6629 (N_6629,N_6338,N_6171);
nand U6630 (N_6630,N_6088,N_6054);
nor U6631 (N_6631,N_6133,N_6000);
and U6632 (N_6632,N_6316,N_6066);
xor U6633 (N_6633,N_6071,N_6234);
nor U6634 (N_6634,N_6169,N_6132);
nand U6635 (N_6635,N_6065,N_6043);
nand U6636 (N_6636,N_6141,N_6367);
and U6637 (N_6637,N_6277,N_6266);
xor U6638 (N_6638,N_6225,N_6242);
and U6639 (N_6639,N_6095,N_6271);
and U6640 (N_6640,N_6218,N_6269);
xnor U6641 (N_6641,N_6108,N_6182);
or U6642 (N_6642,N_6238,N_6030);
or U6643 (N_6643,N_6032,N_6378);
nor U6644 (N_6644,N_6016,N_6232);
or U6645 (N_6645,N_6351,N_6167);
and U6646 (N_6646,N_6347,N_6037);
or U6647 (N_6647,N_6104,N_6385);
nand U6648 (N_6648,N_6381,N_6121);
and U6649 (N_6649,N_6203,N_6087);
and U6650 (N_6650,N_6142,N_6391);
nor U6651 (N_6651,N_6086,N_6348);
or U6652 (N_6652,N_6027,N_6312);
and U6653 (N_6653,N_6051,N_6268);
nand U6654 (N_6654,N_6047,N_6394);
nor U6655 (N_6655,N_6190,N_6042);
and U6656 (N_6656,N_6305,N_6231);
nand U6657 (N_6657,N_6284,N_6103);
or U6658 (N_6658,N_6211,N_6103);
nand U6659 (N_6659,N_6302,N_6391);
xor U6660 (N_6660,N_6217,N_6273);
or U6661 (N_6661,N_6033,N_6000);
and U6662 (N_6662,N_6079,N_6258);
nand U6663 (N_6663,N_6377,N_6366);
nor U6664 (N_6664,N_6095,N_6074);
xor U6665 (N_6665,N_6369,N_6071);
nand U6666 (N_6666,N_6312,N_6186);
or U6667 (N_6667,N_6068,N_6026);
nor U6668 (N_6668,N_6169,N_6353);
or U6669 (N_6669,N_6257,N_6199);
nand U6670 (N_6670,N_6174,N_6078);
nand U6671 (N_6671,N_6212,N_6060);
and U6672 (N_6672,N_6056,N_6091);
nand U6673 (N_6673,N_6262,N_6092);
nand U6674 (N_6674,N_6080,N_6242);
nor U6675 (N_6675,N_6182,N_6117);
nand U6676 (N_6676,N_6357,N_6112);
or U6677 (N_6677,N_6287,N_6176);
xnor U6678 (N_6678,N_6309,N_6070);
nand U6679 (N_6679,N_6230,N_6174);
xnor U6680 (N_6680,N_6075,N_6117);
nand U6681 (N_6681,N_6088,N_6001);
nand U6682 (N_6682,N_6145,N_6382);
xnor U6683 (N_6683,N_6092,N_6344);
xnor U6684 (N_6684,N_6186,N_6046);
xnor U6685 (N_6685,N_6257,N_6177);
or U6686 (N_6686,N_6127,N_6399);
or U6687 (N_6687,N_6173,N_6121);
nand U6688 (N_6688,N_6218,N_6193);
and U6689 (N_6689,N_6373,N_6300);
and U6690 (N_6690,N_6214,N_6089);
xor U6691 (N_6691,N_6365,N_6247);
xor U6692 (N_6692,N_6372,N_6250);
or U6693 (N_6693,N_6240,N_6257);
nand U6694 (N_6694,N_6238,N_6185);
and U6695 (N_6695,N_6238,N_6394);
xor U6696 (N_6696,N_6065,N_6059);
nand U6697 (N_6697,N_6244,N_6138);
and U6698 (N_6698,N_6296,N_6207);
or U6699 (N_6699,N_6139,N_6376);
and U6700 (N_6700,N_6182,N_6009);
or U6701 (N_6701,N_6091,N_6213);
nor U6702 (N_6702,N_6388,N_6046);
or U6703 (N_6703,N_6337,N_6257);
or U6704 (N_6704,N_6169,N_6076);
nor U6705 (N_6705,N_6165,N_6112);
nand U6706 (N_6706,N_6069,N_6150);
nor U6707 (N_6707,N_6198,N_6268);
nor U6708 (N_6708,N_6183,N_6053);
nor U6709 (N_6709,N_6205,N_6053);
nand U6710 (N_6710,N_6352,N_6132);
nor U6711 (N_6711,N_6126,N_6138);
nor U6712 (N_6712,N_6263,N_6035);
or U6713 (N_6713,N_6118,N_6370);
or U6714 (N_6714,N_6373,N_6216);
nor U6715 (N_6715,N_6108,N_6294);
nor U6716 (N_6716,N_6200,N_6110);
and U6717 (N_6717,N_6269,N_6057);
xor U6718 (N_6718,N_6338,N_6059);
xor U6719 (N_6719,N_6192,N_6133);
nor U6720 (N_6720,N_6057,N_6307);
nor U6721 (N_6721,N_6155,N_6318);
nand U6722 (N_6722,N_6116,N_6113);
and U6723 (N_6723,N_6061,N_6183);
and U6724 (N_6724,N_6289,N_6145);
and U6725 (N_6725,N_6131,N_6282);
or U6726 (N_6726,N_6168,N_6362);
nand U6727 (N_6727,N_6087,N_6141);
and U6728 (N_6728,N_6115,N_6399);
nand U6729 (N_6729,N_6020,N_6050);
and U6730 (N_6730,N_6138,N_6117);
nand U6731 (N_6731,N_6263,N_6018);
and U6732 (N_6732,N_6352,N_6208);
nor U6733 (N_6733,N_6393,N_6243);
and U6734 (N_6734,N_6215,N_6115);
nand U6735 (N_6735,N_6199,N_6042);
or U6736 (N_6736,N_6005,N_6134);
nand U6737 (N_6737,N_6327,N_6119);
nand U6738 (N_6738,N_6211,N_6199);
nand U6739 (N_6739,N_6228,N_6181);
nor U6740 (N_6740,N_6344,N_6345);
nor U6741 (N_6741,N_6268,N_6063);
and U6742 (N_6742,N_6129,N_6328);
nand U6743 (N_6743,N_6365,N_6069);
nand U6744 (N_6744,N_6044,N_6006);
xnor U6745 (N_6745,N_6363,N_6152);
nand U6746 (N_6746,N_6112,N_6386);
xor U6747 (N_6747,N_6381,N_6204);
and U6748 (N_6748,N_6059,N_6331);
nand U6749 (N_6749,N_6149,N_6067);
or U6750 (N_6750,N_6196,N_6153);
nand U6751 (N_6751,N_6139,N_6340);
nor U6752 (N_6752,N_6380,N_6323);
and U6753 (N_6753,N_6330,N_6251);
or U6754 (N_6754,N_6024,N_6096);
xnor U6755 (N_6755,N_6397,N_6045);
or U6756 (N_6756,N_6348,N_6004);
or U6757 (N_6757,N_6009,N_6239);
and U6758 (N_6758,N_6071,N_6363);
nand U6759 (N_6759,N_6247,N_6224);
xnor U6760 (N_6760,N_6209,N_6020);
xor U6761 (N_6761,N_6327,N_6348);
and U6762 (N_6762,N_6236,N_6104);
xor U6763 (N_6763,N_6232,N_6389);
and U6764 (N_6764,N_6037,N_6220);
nor U6765 (N_6765,N_6392,N_6323);
and U6766 (N_6766,N_6326,N_6087);
or U6767 (N_6767,N_6332,N_6083);
and U6768 (N_6768,N_6319,N_6179);
nand U6769 (N_6769,N_6255,N_6337);
nand U6770 (N_6770,N_6352,N_6166);
xnor U6771 (N_6771,N_6188,N_6022);
xor U6772 (N_6772,N_6248,N_6217);
xor U6773 (N_6773,N_6021,N_6354);
xor U6774 (N_6774,N_6234,N_6119);
nor U6775 (N_6775,N_6076,N_6342);
and U6776 (N_6776,N_6091,N_6344);
and U6777 (N_6777,N_6195,N_6363);
nand U6778 (N_6778,N_6117,N_6163);
xor U6779 (N_6779,N_6100,N_6268);
nor U6780 (N_6780,N_6177,N_6278);
xnor U6781 (N_6781,N_6326,N_6294);
and U6782 (N_6782,N_6222,N_6339);
nor U6783 (N_6783,N_6100,N_6263);
nor U6784 (N_6784,N_6197,N_6140);
nand U6785 (N_6785,N_6237,N_6155);
xnor U6786 (N_6786,N_6197,N_6025);
xor U6787 (N_6787,N_6130,N_6163);
nor U6788 (N_6788,N_6133,N_6005);
and U6789 (N_6789,N_6130,N_6117);
xor U6790 (N_6790,N_6030,N_6394);
nand U6791 (N_6791,N_6084,N_6252);
or U6792 (N_6792,N_6140,N_6316);
xnor U6793 (N_6793,N_6323,N_6241);
xor U6794 (N_6794,N_6368,N_6183);
xnor U6795 (N_6795,N_6344,N_6070);
nor U6796 (N_6796,N_6133,N_6029);
xnor U6797 (N_6797,N_6343,N_6026);
and U6798 (N_6798,N_6222,N_6146);
or U6799 (N_6799,N_6096,N_6297);
nand U6800 (N_6800,N_6603,N_6762);
xor U6801 (N_6801,N_6612,N_6685);
or U6802 (N_6802,N_6593,N_6674);
nand U6803 (N_6803,N_6658,N_6416);
and U6804 (N_6804,N_6670,N_6592);
nor U6805 (N_6805,N_6598,N_6659);
or U6806 (N_6806,N_6536,N_6437);
xor U6807 (N_6807,N_6664,N_6627);
nor U6808 (N_6808,N_6504,N_6630);
or U6809 (N_6809,N_6464,N_6533);
xor U6810 (N_6810,N_6410,N_6678);
and U6811 (N_6811,N_6700,N_6411);
and U6812 (N_6812,N_6571,N_6525);
nand U6813 (N_6813,N_6716,N_6462);
nand U6814 (N_6814,N_6714,N_6488);
xor U6815 (N_6815,N_6693,N_6417);
and U6816 (N_6816,N_6610,N_6441);
xor U6817 (N_6817,N_6653,N_6463);
nand U6818 (N_6818,N_6643,N_6672);
and U6819 (N_6819,N_6446,N_6471);
nor U6820 (N_6820,N_6620,N_6759);
or U6821 (N_6821,N_6616,N_6505);
nand U6822 (N_6822,N_6535,N_6466);
nand U6823 (N_6823,N_6764,N_6496);
and U6824 (N_6824,N_6420,N_6461);
or U6825 (N_6825,N_6673,N_6640);
nor U6826 (N_6826,N_6622,N_6413);
nor U6827 (N_6827,N_6553,N_6769);
and U6828 (N_6828,N_6549,N_6541);
or U6829 (N_6829,N_6782,N_6711);
nor U6830 (N_6830,N_6430,N_6529);
nor U6831 (N_6831,N_6587,N_6526);
xnor U6832 (N_6832,N_6585,N_6527);
nand U6833 (N_6833,N_6478,N_6698);
nand U6834 (N_6834,N_6418,N_6723);
xnor U6835 (N_6835,N_6491,N_6498);
or U6836 (N_6836,N_6720,N_6511);
nor U6837 (N_6837,N_6677,N_6475);
and U6838 (N_6838,N_6788,N_6433);
nand U6839 (N_6839,N_6727,N_6798);
nand U6840 (N_6840,N_6792,N_6402);
nand U6841 (N_6841,N_6785,N_6794);
xnor U6842 (N_6842,N_6611,N_6739);
nand U6843 (N_6843,N_6539,N_6408);
or U6844 (N_6844,N_6775,N_6765);
nor U6845 (N_6845,N_6669,N_6754);
xnor U6846 (N_6846,N_6486,N_6558);
xnor U6847 (N_6847,N_6712,N_6545);
nand U6848 (N_6848,N_6600,N_6542);
nor U6849 (N_6849,N_6735,N_6731);
nand U6850 (N_6850,N_6540,N_6427);
nor U6851 (N_6851,N_6614,N_6582);
xnor U6852 (N_6852,N_6752,N_6688);
xor U6853 (N_6853,N_6618,N_6734);
or U6854 (N_6854,N_6523,N_6750);
nand U6855 (N_6855,N_6732,N_6569);
nand U6856 (N_6856,N_6636,N_6586);
nor U6857 (N_6857,N_6487,N_6400);
or U6858 (N_6858,N_6479,N_6634);
xor U6859 (N_6859,N_6635,N_6633);
or U6860 (N_6860,N_6607,N_6524);
nand U6861 (N_6861,N_6628,N_6438);
xor U6862 (N_6862,N_6647,N_6605);
nand U6863 (N_6863,N_6662,N_6422);
or U6864 (N_6864,N_6748,N_6546);
and U6865 (N_6865,N_6589,N_6451);
nor U6866 (N_6866,N_6690,N_6744);
or U6867 (N_6867,N_6468,N_6512);
or U6868 (N_6868,N_6440,N_6435);
or U6869 (N_6869,N_6497,N_6426);
nand U6870 (N_6870,N_6613,N_6729);
xnor U6871 (N_6871,N_6531,N_6608);
nor U6872 (N_6872,N_6706,N_6648);
and U6873 (N_6873,N_6449,N_6623);
nor U6874 (N_6874,N_6564,N_6476);
and U6875 (N_6875,N_6573,N_6642);
nor U6876 (N_6876,N_6555,N_6718);
xor U6877 (N_6877,N_6683,N_6768);
or U6878 (N_6878,N_6793,N_6431);
nor U6879 (N_6879,N_6489,N_6588);
and U6880 (N_6880,N_6641,N_6493);
nor U6881 (N_6881,N_6483,N_6518);
and U6882 (N_6882,N_6601,N_6575);
nand U6883 (N_6883,N_6760,N_6660);
xnor U6884 (N_6884,N_6691,N_6455);
xnor U6885 (N_6885,N_6557,N_6442);
or U6886 (N_6886,N_6509,N_6639);
and U6887 (N_6887,N_6652,N_6574);
nand U6888 (N_6888,N_6503,N_6580);
or U6889 (N_6889,N_6767,N_6409);
xor U6890 (N_6890,N_6522,N_6770);
xnor U6891 (N_6891,N_6681,N_6448);
nor U6892 (N_6892,N_6757,N_6758);
and U6893 (N_6893,N_6715,N_6684);
and U6894 (N_6894,N_6406,N_6661);
or U6895 (N_6895,N_6704,N_6710);
xor U6896 (N_6896,N_6457,N_6773);
nor U6897 (N_6897,N_6679,N_6705);
and U6898 (N_6898,N_6507,N_6519);
nor U6899 (N_6899,N_6741,N_6756);
or U6900 (N_6900,N_6783,N_6777);
and U6901 (N_6901,N_6746,N_6733);
nor U6902 (N_6902,N_6469,N_6763);
nor U6903 (N_6903,N_6766,N_6405);
nand U6904 (N_6904,N_6554,N_6506);
or U6905 (N_6905,N_6730,N_6687);
nand U6906 (N_6906,N_6740,N_6452);
xnor U6907 (N_6907,N_6456,N_6532);
nand U6908 (N_6908,N_6521,N_6755);
nor U6909 (N_6909,N_6439,N_6563);
xnor U6910 (N_6910,N_6692,N_6528);
nor U6911 (N_6911,N_6708,N_6599);
nor U6912 (N_6912,N_6703,N_6790);
and U6913 (N_6913,N_6444,N_6717);
nor U6914 (N_6914,N_6774,N_6595);
or U6915 (N_6915,N_6619,N_6638);
and U6916 (N_6916,N_6501,N_6725);
or U6917 (N_6917,N_6454,N_6629);
and U6918 (N_6918,N_6722,N_6772);
and U6919 (N_6919,N_6702,N_6445);
nor U6920 (N_6920,N_6728,N_6548);
nand U6921 (N_6921,N_6434,N_6707);
and U6922 (N_6922,N_6481,N_6726);
nor U6923 (N_6923,N_6631,N_6666);
and U6924 (N_6924,N_6753,N_6514);
xnor U6925 (N_6925,N_6781,N_6537);
nor U6926 (N_6926,N_6671,N_6625);
and U6927 (N_6927,N_6578,N_6577);
nor U6928 (N_6928,N_6745,N_6667);
xor U6929 (N_6929,N_6552,N_6458);
or U6930 (N_6930,N_6637,N_6499);
nand U6931 (N_6931,N_6749,N_6477);
nand U6932 (N_6932,N_6516,N_6695);
or U6933 (N_6933,N_6494,N_6530);
nand U6934 (N_6934,N_6665,N_6484);
xnor U6935 (N_6935,N_6567,N_6615);
nand U6936 (N_6936,N_6737,N_6655);
nor U6937 (N_6937,N_6594,N_6492);
and U6938 (N_6938,N_6645,N_6676);
and U6939 (N_6939,N_6778,N_6584);
and U6940 (N_6940,N_6675,N_6787);
xor U6941 (N_6941,N_6621,N_6649);
nor U6942 (N_6942,N_6550,N_6490);
xor U6943 (N_6943,N_6544,N_6459);
nor U6944 (N_6944,N_6579,N_6590);
nand U6945 (N_6945,N_6551,N_6784);
xor U6946 (N_6946,N_6689,N_6606);
nor U6947 (N_6947,N_6510,N_6414);
xor U6948 (N_6948,N_6650,N_6560);
nand U6949 (N_6949,N_6515,N_6776);
nand U6950 (N_6950,N_6421,N_6412);
xor U6951 (N_6951,N_6566,N_6470);
and U6952 (N_6952,N_6480,N_6596);
or U6953 (N_6953,N_6424,N_6565);
and U6954 (N_6954,N_6508,N_6656);
xor U6955 (N_6955,N_6404,N_6561);
and U6956 (N_6956,N_6436,N_6696);
xor U6957 (N_6957,N_6697,N_6686);
nand U6958 (N_6958,N_6626,N_6576);
and U6959 (N_6959,N_6721,N_6602);
nor U6960 (N_6960,N_6502,N_6403);
and U6961 (N_6961,N_6780,N_6419);
xor U6962 (N_6962,N_6407,N_6751);
and U6963 (N_6963,N_6568,N_6500);
nor U6964 (N_6964,N_6657,N_6791);
or U6965 (N_6965,N_6646,N_6482);
xnor U6966 (N_6966,N_6699,N_6556);
xor U6967 (N_6967,N_6543,N_6415);
or U6968 (N_6968,N_6789,N_6591);
and U6969 (N_6969,N_6654,N_6495);
and U6970 (N_6970,N_6473,N_6624);
nor U6971 (N_6971,N_6795,N_6572);
or U6972 (N_6972,N_6786,N_6538);
and U6973 (N_6973,N_6709,N_6779);
and U6974 (N_6974,N_6583,N_6632);
nor U6975 (N_6975,N_6736,N_6747);
or U6976 (N_6976,N_6663,N_6797);
or U6977 (N_6977,N_6724,N_6713);
nor U6978 (N_6978,N_6401,N_6570);
nor U6979 (N_6979,N_6513,N_6453);
or U6980 (N_6980,N_6609,N_6559);
or U6981 (N_6981,N_6534,N_6443);
and U6982 (N_6982,N_6432,N_6447);
and U6983 (N_6983,N_6581,N_6547);
xnor U6984 (N_6984,N_6742,N_6668);
and U6985 (N_6985,N_6450,N_6425);
nor U6986 (N_6986,N_6701,N_6465);
or U6987 (N_6987,N_6467,N_6719);
xnor U6988 (N_6988,N_6738,N_6796);
and U6989 (N_6989,N_6474,N_6743);
and U6990 (N_6990,N_6562,N_6651);
xnor U6991 (N_6991,N_6682,N_6597);
nand U6992 (N_6992,N_6460,N_6694);
or U6993 (N_6993,N_6429,N_6520);
nor U6994 (N_6994,N_6428,N_6423);
or U6995 (N_6995,N_6485,N_6517);
or U6996 (N_6996,N_6680,N_6771);
or U6997 (N_6997,N_6761,N_6617);
nand U6998 (N_6998,N_6604,N_6644);
nor U6999 (N_6999,N_6472,N_6799);
nor U7000 (N_7000,N_6576,N_6734);
nor U7001 (N_7001,N_6455,N_6664);
nand U7002 (N_7002,N_6486,N_6602);
or U7003 (N_7003,N_6565,N_6722);
nor U7004 (N_7004,N_6632,N_6622);
nand U7005 (N_7005,N_6591,N_6713);
xor U7006 (N_7006,N_6405,N_6606);
or U7007 (N_7007,N_6629,N_6475);
or U7008 (N_7008,N_6577,N_6477);
nor U7009 (N_7009,N_6763,N_6632);
and U7010 (N_7010,N_6499,N_6484);
and U7011 (N_7011,N_6511,N_6713);
xnor U7012 (N_7012,N_6534,N_6465);
nor U7013 (N_7013,N_6719,N_6588);
nor U7014 (N_7014,N_6623,N_6442);
nand U7015 (N_7015,N_6758,N_6796);
or U7016 (N_7016,N_6494,N_6589);
or U7017 (N_7017,N_6606,N_6537);
and U7018 (N_7018,N_6738,N_6756);
and U7019 (N_7019,N_6733,N_6580);
nor U7020 (N_7020,N_6754,N_6726);
xor U7021 (N_7021,N_6438,N_6552);
nand U7022 (N_7022,N_6555,N_6729);
xnor U7023 (N_7023,N_6769,N_6733);
nor U7024 (N_7024,N_6779,N_6481);
xor U7025 (N_7025,N_6701,N_6476);
nand U7026 (N_7026,N_6466,N_6689);
and U7027 (N_7027,N_6606,N_6573);
and U7028 (N_7028,N_6419,N_6690);
xor U7029 (N_7029,N_6664,N_6409);
or U7030 (N_7030,N_6414,N_6548);
nor U7031 (N_7031,N_6549,N_6576);
and U7032 (N_7032,N_6420,N_6536);
or U7033 (N_7033,N_6790,N_6787);
nand U7034 (N_7034,N_6542,N_6526);
nand U7035 (N_7035,N_6541,N_6693);
and U7036 (N_7036,N_6492,N_6772);
nor U7037 (N_7037,N_6730,N_6663);
xnor U7038 (N_7038,N_6464,N_6502);
xnor U7039 (N_7039,N_6711,N_6517);
nand U7040 (N_7040,N_6595,N_6413);
nor U7041 (N_7041,N_6403,N_6716);
nor U7042 (N_7042,N_6422,N_6745);
and U7043 (N_7043,N_6422,N_6695);
nand U7044 (N_7044,N_6422,N_6540);
nor U7045 (N_7045,N_6576,N_6468);
nand U7046 (N_7046,N_6469,N_6630);
and U7047 (N_7047,N_6485,N_6422);
nand U7048 (N_7048,N_6768,N_6762);
xor U7049 (N_7049,N_6459,N_6528);
xnor U7050 (N_7050,N_6634,N_6532);
and U7051 (N_7051,N_6663,N_6401);
or U7052 (N_7052,N_6603,N_6684);
nor U7053 (N_7053,N_6478,N_6435);
xor U7054 (N_7054,N_6514,N_6495);
xnor U7055 (N_7055,N_6744,N_6727);
xor U7056 (N_7056,N_6599,N_6501);
nor U7057 (N_7057,N_6593,N_6746);
or U7058 (N_7058,N_6701,N_6466);
xor U7059 (N_7059,N_6609,N_6653);
nand U7060 (N_7060,N_6433,N_6513);
and U7061 (N_7061,N_6531,N_6781);
nor U7062 (N_7062,N_6573,N_6662);
nor U7063 (N_7063,N_6550,N_6526);
xor U7064 (N_7064,N_6702,N_6762);
nor U7065 (N_7065,N_6456,N_6786);
or U7066 (N_7066,N_6728,N_6651);
and U7067 (N_7067,N_6498,N_6780);
nor U7068 (N_7068,N_6495,N_6661);
xnor U7069 (N_7069,N_6604,N_6466);
nand U7070 (N_7070,N_6502,N_6579);
nand U7071 (N_7071,N_6423,N_6679);
nor U7072 (N_7072,N_6545,N_6799);
nor U7073 (N_7073,N_6713,N_6734);
nor U7074 (N_7074,N_6580,N_6687);
and U7075 (N_7075,N_6461,N_6434);
nand U7076 (N_7076,N_6673,N_6486);
nor U7077 (N_7077,N_6672,N_6511);
and U7078 (N_7078,N_6656,N_6481);
nand U7079 (N_7079,N_6470,N_6703);
or U7080 (N_7080,N_6758,N_6548);
xor U7081 (N_7081,N_6750,N_6474);
and U7082 (N_7082,N_6763,N_6710);
or U7083 (N_7083,N_6439,N_6441);
nand U7084 (N_7084,N_6726,N_6602);
and U7085 (N_7085,N_6742,N_6424);
and U7086 (N_7086,N_6788,N_6412);
nand U7087 (N_7087,N_6796,N_6587);
xor U7088 (N_7088,N_6776,N_6590);
and U7089 (N_7089,N_6628,N_6463);
nand U7090 (N_7090,N_6416,N_6404);
nand U7091 (N_7091,N_6542,N_6778);
nor U7092 (N_7092,N_6599,N_6401);
xor U7093 (N_7093,N_6631,N_6532);
and U7094 (N_7094,N_6585,N_6551);
and U7095 (N_7095,N_6430,N_6473);
nor U7096 (N_7096,N_6614,N_6559);
nor U7097 (N_7097,N_6720,N_6531);
nand U7098 (N_7098,N_6443,N_6638);
and U7099 (N_7099,N_6541,N_6534);
nand U7100 (N_7100,N_6427,N_6634);
or U7101 (N_7101,N_6604,N_6698);
or U7102 (N_7102,N_6738,N_6637);
nor U7103 (N_7103,N_6766,N_6789);
and U7104 (N_7104,N_6618,N_6524);
and U7105 (N_7105,N_6628,N_6739);
xnor U7106 (N_7106,N_6443,N_6777);
or U7107 (N_7107,N_6614,N_6523);
and U7108 (N_7108,N_6544,N_6456);
nand U7109 (N_7109,N_6776,N_6738);
nand U7110 (N_7110,N_6528,N_6468);
or U7111 (N_7111,N_6549,N_6551);
nand U7112 (N_7112,N_6660,N_6539);
nand U7113 (N_7113,N_6428,N_6529);
nand U7114 (N_7114,N_6701,N_6580);
nand U7115 (N_7115,N_6619,N_6614);
xnor U7116 (N_7116,N_6607,N_6710);
xnor U7117 (N_7117,N_6404,N_6467);
xor U7118 (N_7118,N_6739,N_6718);
and U7119 (N_7119,N_6407,N_6410);
or U7120 (N_7120,N_6490,N_6472);
xnor U7121 (N_7121,N_6632,N_6676);
or U7122 (N_7122,N_6579,N_6678);
nand U7123 (N_7123,N_6569,N_6653);
nand U7124 (N_7124,N_6779,N_6705);
nor U7125 (N_7125,N_6404,N_6479);
nand U7126 (N_7126,N_6648,N_6523);
nor U7127 (N_7127,N_6685,N_6484);
and U7128 (N_7128,N_6508,N_6785);
nor U7129 (N_7129,N_6474,N_6620);
xnor U7130 (N_7130,N_6774,N_6561);
xor U7131 (N_7131,N_6404,N_6774);
and U7132 (N_7132,N_6551,N_6741);
nand U7133 (N_7133,N_6539,N_6457);
or U7134 (N_7134,N_6667,N_6439);
nor U7135 (N_7135,N_6789,N_6599);
nor U7136 (N_7136,N_6759,N_6730);
or U7137 (N_7137,N_6481,N_6620);
xnor U7138 (N_7138,N_6476,N_6454);
and U7139 (N_7139,N_6620,N_6510);
nor U7140 (N_7140,N_6482,N_6623);
or U7141 (N_7141,N_6408,N_6577);
xnor U7142 (N_7142,N_6752,N_6493);
and U7143 (N_7143,N_6593,N_6788);
nand U7144 (N_7144,N_6562,N_6759);
or U7145 (N_7145,N_6475,N_6796);
and U7146 (N_7146,N_6786,N_6627);
xor U7147 (N_7147,N_6724,N_6462);
nor U7148 (N_7148,N_6420,N_6404);
and U7149 (N_7149,N_6522,N_6696);
nand U7150 (N_7150,N_6449,N_6797);
or U7151 (N_7151,N_6538,N_6624);
and U7152 (N_7152,N_6621,N_6633);
xnor U7153 (N_7153,N_6544,N_6522);
and U7154 (N_7154,N_6425,N_6623);
nor U7155 (N_7155,N_6495,N_6698);
or U7156 (N_7156,N_6508,N_6527);
or U7157 (N_7157,N_6640,N_6569);
and U7158 (N_7158,N_6647,N_6514);
or U7159 (N_7159,N_6630,N_6759);
and U7160 (N_7160,N_6421,N_6785);
or U7161 (N_7161,N_6748,N_6603);
nand U7162 (N_7162,N_6711,N_6446);
nor U7163 (N_7163,N_6539,N_6495);
nand U7164 (N_7164,N_6527,N_6418);
or U7165 (N_7165,N_6788,N_6721);
nor U7166 (N_7166,N_6792,N_6662);
nand U7167 (N_7167,N_6766,N_6534);
and U7168 (N_7168,N_6633,N_6434);
nand U7169 (N_7169,N_6542,N_6653);
or U7170 (N_7170,N_6733,N_6514);
nand U7171 (N_7171,N_6532,N_6719);
nand U7172 (N_7172,N_6535,N_6658);
and U7173 (N_7173,N_6628,N_6787);
xnor U7174 (N_7174,N_6421,N_6662);
nand U7175 (N_7175,N_6516,N_6678);
nor U7176 (N_7176,N_6711,N_6575);
nor U7177 (N_7177,N_6476,N_6499);
xnor U7178 (N_7178,N_6593,N_6678);
nand U7179 (N_7179,N_6655,N_6759);
or U7180 (N_7180,N_6591,N_6672);
and U7181 (N_7181,N_6637,N_6498);
or U7182 (N_7182,N_6601,N_6592);
and U7183 (N_7183,N_6696,N_6723);
nand U7184 (N_7184,N_6640,N_6570);
nor U7185 (N_7185,N_6434,N_6605);
and U7186 (N_7186,N_6587,N_6475);
and U7187 (N_7187,N_6668,N_6473);
or U7188 (N_7188,N_6762,N_6710);
and U7189 (N_7189,N_6756,N_6425);
or U7190 (N_7190,N_6523,N_6733);
nor U7191 (N_7191,N_6639,N_6603);
nor U7192 (N_7192,N_6740,N_6723);
xnor U7193 (N_7193,N_6797,N_6668);
xor U7194 (N_7194,N_6625,N_6437);
nor U7195 (N_7195,N_6553,N_6545);
xor U7196 (N_7196,N_6401,N_6760);
nor U7197 (N_7197,N_6630,N_6711);
and U7198 (N_7198,N_6702,N_6422);
and U7199 (N_7199,N_6605,N_6444);
or U7200 (N_7200,N_7092,N_7162);
nand U7201 (N_7201,N_6840,N_7059);
nand U7202 (N_7202,N_7196,N_6937);
or U7203 (N_7203,N_7117,N_7017);
xnor U7204 (N_7204,N_6864,N_6944);
nand U7205 (N_7205,N_7172,N_6917);
xor U7206 (N_7206,N_6888,N_7097);
and U7207 (N_7207,N_6902,N_7166);
nand U7208 (N_7208,N_6988,N_6914);
or U7209 (N_7209,N_6906,N_7121);
and U7210 (N_7210,N_6996,N_6878);
or U7211 (N_7211,N_6825,N_7078);
xnor U7212 (N_7212,N_7113,N_6813);
and U7213 (N_7213,N_7047,N_7108);
nor U7214 (N_7214,N_6950,N_6828);
nor U7215 (N_7215,N_6926,N_6810);
and U7216 (N_7216,N_6838,N_7192);
nor U7217 (N_7217,N_6946,N_6871);
nor U7218 (N_7218,N_7091,N_7020);
nand U7219 (N_7219,N_6970,N_6829);
nor U7220 (N_7220,N_7007,N_7120);
nand U7221 (N_7221,N_6977,N_7013);
xor U7222 (N_7222,N_6851,N_6862);
xor U7223 (N_7223,N_7105,N_7174);
nor U7224 (N_7224,N_6932,N_7035);
and U7225 (N_7225,N_7008,N_6963);
xor U7226 (N_7226,N_7137,N_7039);
nor U7227 (N_7227,N_7000,N_7094);
and U7228 (N_7228,N_6811,N_7150);
or U7229 (N_7229,N_6887,N_6848);
and U7230 (N_7230,N_6859,N_6817);
nand U7231 (N_7231,N_6891,N_7132);
xor U7232 (N_7232,N_6989,N_7089);
nand U7233 (N_7233,N_7067,N_7096);
or U7234 (N_7234,N_7074,N_7019);
xor U7235 (N_7235,N_7180,N_7084);
nor U7236 (N_7236,N_7189,N_7048);
nor U7237 (N_7237,N_6857,N_6834);
nor U7238 (N_7238,N_7186,N_7011);
or U7239 (N_7239,N_7182,N_6923);
xor U7240 (N_7240,N_7038,N_6849);
nand U7241 (N_7241,N_7001,N_7041);
or U7242 (N_7242,N_7027,N_7109);
xnor U7243 (N_7243,N_7076,N_6876);
xor U7244 (N_7244,N_6965,N_7064);
or U7245 (N_7245,N_7088,N_6998);
or U7246 (N_7246,N_6985,N_6837);
nand U7247 (N_7247,N_7024,N_7181);
nor U7248 (N_7248,N_6841,N_6873);
nor U7249 (N_7249,N_6918,N_6905);
nand U7250 (N_7250,N_7055,N_6819);
xor U7251 (N_7251,N_6896,N_6883);
nor U7252 (N_7252,N_7145,N_6933);
nor U7253 (N_7253,N_6928,N_7036);
or U7254 (N_7254,N_7033,N_6874);
nor U7255 (N_7255,N_7177,N_6969);
and U7256 (N_7256,N_7183,N_6904);
or U7257 (N_7257,N_7133,N_6952);
and U7258 (N_7258,N_7114,N_6842);
or U7259 (N_7259,N_7191,N_7100);
nand U7260 (N_7260,N_7131,N_7073);
nand U7261 (N_7261,N_7135,N_7103);
nand U7262 (N_7262,N_7195,N_6967);
nor U7263 (N_7263,N_7151,N_6916);
nand U7264 (N_7264,N_6858,N_6850);
nor U7265 (N_7265,N_6846,N_7026);
xnor U7266 (N_7266,N_6884,N_7141);
nor U7267 (N_7267,N_6854,N_7063);
xor U7268 (N_7268,N_6939,N_6968);
nor U7269 (N_7269,N_6853,N_6861);
and U7270 (N_7270,N_7045,N_7106);
nor U7271 (N_7271,N_6881,N_7075);
nand U7272 (N_7272,N_7102,N_6991);
nand U7273 (N_7273,N_6865,N_6856);
xor U7274 (N_7274,N_7146,N_6921);
nand U7275 (N_7275,N_7030,N_6978);
xor U7276 (N_7276,N_7079,N_7126);
or U7277 (N_7277,N_7193,N_6855);
nand U7278 (N_7278,N_7168,N_7157);
nor U7279 (N_7279,N_7051,N_7171);
or U7280 (N_7280,N_6826,N_7134);
and U7281 (N_7281,N_6993,N_6957);
xnor U7282 (N_7282,N_7056,N_7003);
and U7283 (N_7283,N_7197,N_6992);
or U7284 (N_7284,N_7149,N_6909);
and U7285 (N_7285,N_6990,N_6930);
nor U7286 (N_7286,N_7163,N_6924);
or U7287 (N_7287,N_6972,N_7184);
and U7288 (N_7288,N_6955,N_6979);
or U7289 (N_7289,N_6984,N_7148);
xnor U7290 (N_7290,N_7085,N_7175);
xnor U7291 (N_7291,N_6897,N_6835);
and U7292 (N_7292,N_6942,N_7169);
or U7293 (N_7293,N_6997,N_7142);
and U7294 (N_7294,N_6925,N_7115);
xnor U7295 (N_7295,N_6959,N_7040);
nand U7296 (N_7296,N_7021,N_6886);
and U7297 (N_7297,N_6995,N_6934);
or U7298 (N_7298,N_7170,N_7116);
or U7299 (N_7299,N_6814,N_6833);
xor U7300 (N_7300,N_7068,N_6958);
or U7301 (N_7301,N_6877,N_6895);
and U7302 (N_7302,N_6976,N_6831);
xor U7303 (N_7303,N_7129,N_7049);
and U7304 (N_7304,N_6948,N_7160);
or U7305 (N_7305,N_7086,N_7031);
nand U7306 (N_7306,N_7173,N_7054);
xnor U7307 (N_7307,N_6845,N_6919);
or U7308 (N_7308,N_7152,N_6818);
or U7309 (N_7309,N_7034,N_6815);
or U7310 (N_7310,N_7093,N_6879);
and U7311 (N_7311,N_6847,N_7065);
and U7312 (N_7312,N_6824,N_7005);
and U7313 (N_7313,N_6900,N_6869);
or U7314 (N_7314,N_7104,N_7138);
nand U7315 (N_7315,N_7198,N_6938);
xnor U7316 (N_7316,N_6945,N_7111);
xor U7317 (N_7317,N_6800,N_6894);
or U7318 (N_7318,N_7187,N_6901);
or U7319 (N_7319,N_6807,N_6872);
or U7320 (N_7320,N_7053,N_6867);
nor U7321 (N_7321,N_6983,N_7128);
nor U7322 (N_7322,N_7071,N_7147);
and U7323 (N_7323,N_7122,N_6860);
xnor U7324 (N_7324,N_6999,N_7012);
and U7325 (N_7325,N_6806,N_7025);
xor U7326 (N_7326,N_7070,N_6836);
or U7327 (N_7327,N_7099,N_6920);
nor U7328 (N_7328,N_7098,N_6823);
nand U7329 (N_7329,N_7127,N_7124);
xnor U7330 (N_7330,N_6980,N_6975);
nand U7331 (N_7331,N_7123,N_7154);
nor U7332 (N_7332,N_7022,N_7110);
and U7333 (N_7333,N_7010,N_7058);
nor U7334 (N_7334,N_6922,N_7082);
or U7335 (N_7335,N_6940,N_6903);
or U7336 (N_7336,N_6947,N_6852);
or U7337 (N_7337,N_7090,N_7066);
and U7338 (N_7338,N_6843,N_7062);
nand U7339 (N_7339,N_6808,N_7188);
and U7340 (N_7340,N_7139,N_6870);
nor U7341 (N_7341,N_6885,N_6927);
or U7342 (N_7342,N_6804,N_6911);
nand U7343 (N_7343,N_6908,N_7130);
nor U7344 (N_7344,N_6892,N_7052);
nor U7345 (N_7345,N_6964,N_7028);
and U7346 (N_7346,N_7118,N_7158);
and U7347 (N_7347,N_6936,N_7143);
xnor U7348 (N_7348,N_7080,N_7057);
or U7349 (N_7349,N_6951,N_6961);
or U7350 (N_7350,N_7006,N_6986);
nand U7351 (N_7351,N_7095,N_6935);
and U7352 (N_7352,N_6889,N_6953);
and U7353 (N_7353,N_7159,N_7144);
nand U7354 (N_7354,N_7004,N_7077);
nor U7355 (N_7355,N_7190,N_7140);
nor U7356 (N_7356,N_7050,N_7199);
and U7357 (N_7357,N_7112,N_7083);
and U7358 (N_7358,N_7179,N_7023);
xor U7359 (N_7359,N_6801,N_6974);
nor U7360 (N_7360,N_7161,N_6812);
nand U7361 (N_7361,N_6816,N_6910);
nand U7362 (N_7362,N_7194,N_7125);
nor U7363 (N_7363,N_7185,N_7018);
or U7364 (N_7364,N_6821,N_6943);
and U7365 (N_7365,N_6915,N_7101);
and U7366 (N_7366,N_6931,N_7155);
and U7367 (N_7367,N_7167,N_6981);
nor U7368 (N_7368,N_6960,N_6844);
nand U7369 (N_7369,N_7016,N_7072);
nand U7370 (N_7370,N_7178,N_6898);
and U7371 (N_7371,N_7042,N_6803);
nor U7372 (N_7372,N_6987,N_7164);
xor U7373 (N_7373,N_6966,N_7014);
and U7374 (N_7374,N_7015,N_6868);
xor U7375 (N_7375,N_6954,N_7032);
and U7376 (N_7376,N_6994,N_7037);
xor U7377 (N_7377,N_6839,N_6832);
nand U7378 (N_7378,N_7153,N_7087);
xor U7379 (N_7379,N_6827,N_7060);
or U7380 (N_7380,N_6822,N_6890);
or U7381 (N_7381,N_6820,N_6866);
and U7382 (N_7382,N_6929,N_7061);
nand U7383 (N_7383,N_7107,N_6956);
or U7384 (N_7384,N_6949,N_6913);
and U7385 (N_7385,N_7119,N_7044);
nand U7386 (N_7386,N_6875,N_7043);
xor U7387 (N_7387,N_7165,N_7069);
nand U7388 (N_7388,N_6973,N_6805);
nand U7389 (N_7389,N_6912,N_6809);
xor U7390 (N_7390,N_7176,N_6971);
and U7391 (N_7391,N_6962,N_6899);
xnor U7392 (N_7392,N_6982,N_7002);
and U7393 (N_7393,N_6802,N_6893);
nand U7394 (N_7394,N_7136,N_7156);
nor U7395 (N_7395,N_7081,N_6941);
nor U7396 (N_7396,N_7046,N_6880);
nor U7397 (N_7397,N_6907,N_7029);
or U7398 (N_7398,N_6882,N_7009);
or U7399 (N_7399,N_6863,N_6830);
or U7400 (N_7400,N_6919,N_6916);
nor U7401 (N_7401,N_7077,N_6925);
xnor U7402 (N_7402,N_7014,N_6970);
and U7403 (N_7403,N_7052,N_6986);
and U7404 (N_7404,N_6944,N_6916);
xnor U7405 (N_7405,N_7044,N_7118);
or U7406 (N_7406,N_7005,N_6855);
nor U7407 (N_7407,N_6861,N_7097);
and U7408 (N_7408,N_6891,N_6886);
nand U7409 (N_7409,N_6961,N_6947);
nand U7410 (N_7410,N_6999,N_7016);
nor U7411 (N_7411,N_7071,N_7138);
and U7412 (N_7412,N_7185,N_6813);
and U7413 (N_7413,N_6907,N_7138);
nand U7414 (N_7414,N_6998,N_6839);
or U7415 (N_7415,N_6929,N_6824);
or U7416 (N_7416,N_6979,N_6843);
xnor U7417 (N_7417,N_6833,N_7164);
xor U7418 (N_7418,N_7197,N_6967);
nor U7419 (N_7419,N_6868,N_6867);
nand U7420 (N_7420,N_6919,N_7024);
and U7421 (N_7421,N_7184,N_6856);
or U7422 (N_7422,N_7115,N_7079);
xnor U7423 (N_7423,N_7066,N_7173);
nor U7424 (N_7424,N_7102,N_7028);
and U7425 (N_7425,N_6828,N_6915);
and U7426 (N_7426,N_7136,N_6850);
xor U7427 (N_7427,N_7130,N_6999);
or U7428 (N_7428,N_7031,N_6876);
nand U7429 (N_7429,N_7040,N_6851);
or U7430 (N_7430,N_6898,N_6960);
nand U7431 (N_7431,N_7169,N_7000);
xnor U7432 (N_7432,N_6837,N_7050);
nand U7433 (N_7433,N_6950,N_6998);
nand U7434 (N_7434,N_6860,N_7199);
or U7435 (N_7435,N_7168,N_7129);
nor U7436 (N_7436,N_7023,N_7191);
or U7437 (N_7437,N_6836,N_7182);
and U7438 (N_7438,N_6970,N_7104);
or U7439 (N_7439,N_7136,N_6993);
or U7440 (N_7440,N_6875,N_7199);
nand U7441 (N_7441,N_7004,N_6967);
xnor U7442 (N_7442,N_6872,N_6813);
xnor U7443 (N_7443,N_7083,N_7125);
or U7444 (N_7444,N_7075,N_7030);
nand U7445 (N_7445,N_6882,N_6827);
nand U7446 (N_7446,N_7161,N_7122);
and U7447 (N_7447,N_7133,N_7116);
and U7448 (N_7448,N_7023,N_6987);
and U7449 (N_7449,N_7176,N_7188);
or U7450 (N_7450,N_6828,N_7140);
and U7451 (N_7451,N_7045,N_6909);
nand U7452 (N_7452,N_7176,N_7136);
and U7453 (N_7453,N_7071,N_6948);
or U7454 (N_7454,N_6833,N_6940);
nor U7455 (N_7455,N_6811,N_7102);
or U7456 (N_7456,N_7109,N_6895);
nand U7457 (N_7457,N_6953,N_7101);
nand U7458 (N_7458,N_7044,N_7172);
nor U7459 (N_7459,N_7028,N_7007);
and U7460 (N_7460,N_7013,N_6901);
nor U7461 (N_7461,N_7019,N_7174);
nor U7462 (N_7462,N_6838,N_6848);
nand U7463 (N_7463,N_7149,N_6851);
or U7464 (N_7464,N_6897,N_6898);
nor U7465 (N_7465,N_6887,N_7149);
and U7466 (N_7466,N_7103,N_7192);
nor U7467 (N_7467,N_6927,N_6846);
nand U7468 (N_7468,N_7170,N_7123);
nand U7469 (N_7469,N_7074,N_7093);
xor U7470 (N_7470,N_7105,N_6904);
xnor U7471 (N_7471,N_6965,N_6959);
or U7472 (N_7472,N_7113,N_7074);
or U7473 (N_7473,N_7104,N_6826);
or U7474 (N_7474,N_7044,N_6822);
xor U7475 (N_7475,N_6846,N_6963);
nand U7476 (N_7476,N_6915,N_7003);
and U7477 (N_7477,N_6966,N_6855);
nand U7478 (N_7478,N_7083,N_6926);
or U7479 (N_7479,N_6944,N_6946);
nand U7480 (N_7480,N_6904,N_7052);
nand U7481 (N_7481,N_6927,N_7011);
nand U7482 (N_7482,N_7140,N_6905);
xor U7483 (N_7483,N_6926,N_6876);
nand U7484 (N_7484,N_7177,N_6958);
xnor U7485 (N_7485,N_7071,N_6842);
nor U7486 (N_7486,N_6821,N_6977);
or U7487 (N_7487,N_7094,N_6991);
nand U7488 (N_7488,N_7083,N_6832);
xor U7489 (N_7489,N_6957,N_7050);
and U7490 (N_7490,N_6966,N_7170);
and U7491 (N_7491,N_6998,N_7108);
or U7492 (N_7492,N_6993,N_7072);
nor U7493 (N_7493,N_7108,N_6882);
or U7494 (N_7494,N_6860,N_6910);
or U7495 (N_7495,N_6962,N_6986);
and U7496 (N_7496,N_6900,N_6838);
nor U7497 (N_7497,N_6930,N_7036);
xnor U7498 (N_7498,N_6862,N_6815);
nor U7499 (N_7499,N_6811,N_6949);
nand U7500 (N_7500,N_7188,N_6930);
and U7501 (N_7501,N_7199,N_6983);
nand U7502 (N_7502,N_6831,N_7036);
nand U7503 (N_7503,N_7111,N_6832);
nor U7504 (N_7504,N_7051,N_6935);
xor U7505 (N_7505,N_7023,N_6941);
nand U7506 (N_7506,N_7105,N_6826);
and U7507 (N_7507,N_7120,N_7192);
nand U7508 (N_7508,N_6803,N_7113);
or U7509 (N_7509,N_7170,N_6951);
and U7510 (N_7510,N_7145,N_7008);
and U7511 (N_7511,N_7060,N_7041);
nand U7512 (N_7512,N_7185,N_6987);
nand U7513 (N_7513,N_6931,N_7037);
xor U7514 (N_7514,N_7106,N_7177);
nand U7515 (N_7515,N_7194,N_7073);
nor U7516 (N_7516,N_6927,N_6947);
or U7517 (N_7517,N_7145,N_6996);
and U7518 (N_7518,N_6880,N_6978);
and U7519 (N_7519,N_6992,N_7080);
nand U7520 (N_7520,N_6858,N_7122);
nor U7521 (N_7521,N_6948,N_6803);
or U7522 (N_7522,N_6863,N_6825);
or U7523 (N_7523,N_7064,N_6843);
nor U7524 (N_7524,N_7037,N_7026);
or U7525 (N_7525,N_7112,N_6822);
xnor U7526 (N_7526,N_6895,N_7016);
nor U7527 (N_7527,N_7102,N_7093);
or U7528 (N_7528,N_7110,N_7142);
or U7529 (N_7529,N_7024,N_6879);
or U7530 (N_7530,N_6959,N_7160);
and U7531 (N_7531,N_6900,N_6862);
xnor U7532 (N_7532,N_7123,N_6911);
xor U7533 (N_7533,N_6815,N_6810);
xnor U7534 (N_7534,N_6880,N_6982);
nand U7535 (N_7535,N_7182,N_6999);
nor U7536 (N_7536,N_7162,N_6893);
nand U7537 (N_7537,N_7092,N_6886);
nand U7538 (N_7538,N_7087,N_7186);
xnor U7539 (N_7539,N_6976,N_6883);
nor U7540 (N_7540,N_7053,N_6946);
or U7541 (N_7541,N_6804,N_6950);
nor U7542 (N_7542,N_7112,N_7036);
nor U7543 (N_7543,N_6897,N_7180);
nor U7544 (N_7544,N_6917,N_6844);
xnor U7545 (N_7545,N_6802,N_7039);
nor U7546 (N_7546,N_7141,N_6817);
xor U7547 (N_7547,N_7029,N_6888);
and U7548 (N_7548,N_6998,N_6848);
nor U7549 (N_7549,N_7085,N_7112);
xor U7550 (N_7550,N_7100,N_6915);
or U7551 (N_7551,N_7016,N_6820);
nand U7552 (N_7552,N_6913,N_7197);
nor U7553 (N_7553,N_6978,N_6922);
nand U7554 (N_7554,N_7018,N_7154);
nand U7555 (N_7555,N_7160,N_6800);
xnor U7556 (N_7556,N_7130,N_7167);
nand U7557 (N_7557,N_7002,N_6988);
nor U7558 (N_7558,N_7125,N_7075);
nor U7559 (N_7559,N_7004,N_7191);
or U7560 (N_7560,N_6988,N_7184);
xnor U7561 (N_7561,N_6949,N_6908);
nand U7562 (N_7562,N_6879,N_6812);
or U7563 (N_7563,N_7061,N_7108);
and U7564 (N_7564,N_7148,N_7041);
nand U7565 (N_7565,N_6969,N_7096);
nand U7566 (N_7566,N_7055,N_7016);
nor U7567 (N_7567,N_6834,N_7089);
nand U7568 (N_7568,N_6908,N_6856);
or U7569 (N_7569,N_7172,N_7043);
nand U7570 (N_7570,N_7049,N_6816);
nor U7571 (N_7571,N_6885,N_7105);
nor U7572 (N_7572,N_7055,N_6839);
xnor U7573 (N_7573,N_7192,N_6941);
nor U7574 (N_7574,N_7126,N_6917);
xor U7575 (N_7575,N_6855,N_6943);
nor U7576 (N_7576,N_7004,N_7097);
or U7577 (N_7577,N_7149,N_6919);
nor U7578 (N_7578,N_7046,N_6820);
nor U7579 (N_7579,N_7143,N_6822);
or U7580 (N_7580,N_6933,N_7141);
or U7581 (N_7581,N_6916,N_6892);
xnor U7582 (N_7582,N_7179,N_7094);
and U7583 (N_7583,N_7098,N_7088);
xnor U7584 (N_7584,N_6997,N_7154);
xor U7585 (N_7585,N_7056,N_7113);
nand U7586 (N_7586,N_7152,N_6815);
nor U7587 (N_7587,N_6970,N_7065);
nor U7588 (N_7588,N_7180,N_7112);
nand U7589 (N_7589,N_6812,N_7175);
and U7590 (N_7590,N_6951,N_6804);
or U7591 (N_7591,N_6854,N_7022);
nand U7592 (N_7592,N_7064,N_7083);
nor U7593 (N_7593,N_6804,N_6958);
nand U7594 (N_7594,N_6839,N_6932);
nor U7595 (N_7595,N_7118,N_7086);
nand U7596 (N_7596,N_6910,N_7148);
nor U7597 (N_7597,N_6883,N_6907);
xnor U7598 (N_7598,N_6975,N_7150);
nand U7599 (N_7599,N_7010,N_6903);
or U7600 (N_7600,N_7333,N_7575);
or U7601 (N_7601,N_7336,N_7272);
nor U7602 (N_7602,N_7418,N_7407);
and U7603 (N_7603,N_7513,N_7254);
and U7604 (N_7604,N_7402,N_7275);
nor U7605 (N_7605,N_7561,N_7289);
xor U7606 (N_7606,N_7568,N_7494);
nor U7607 (N_7607,N_7586,N_7538);
nor U7608 (N_7608,N_7365,N_7565);
and U7609 (N_7609,N_7306,N_7342);
nand U7610 (N_7610,N_7371,N_7435);
or U7611 (N_7611,N_7355,N_7301);
xor U7612 (N_7612,N_7462,N_7475);
xor U7613 (N_7613,N_7588,N_7532);
or U7614 (N_7614,N_7359,N_7376);
and U7615 (N_7615,N_7375,N_7304);
xor U7616 (N_7616,N_7491,N_7528);
xor U7617 (N_7617,N_7283,N_7389);
xnor U7618 (N_7618,N_7471,N_7298);
xor U7619 (N_7619,N_7286,N_7244);
and U7620 (N_7620,N_7506,N_7378);
or U7621 (N_7621,N_7234,N_7539);
and U7622 (N_7622,N_7449,N_7458);
or U7623 (N_7623,N_7411,N_7570);
nand U7624 (N_7624,N_7233,N_7287);
and U7625 (N_7625,N_7522,N_7536);
nand U7626 (N_7626,N_7273,N_7447);
or U7627 (N_7627,N_7457,N_7578);
nor U7628 (N_7628,N_7476,N_7481);
and U7629 (N_7629,N_7503,N_7305);
or U7630 (N_7630,N_7470,N_7216);
and U7631 (N_7631,N_7324,N_7400);
and U7632 (N_7632,N_7420,N_7227);
or U7633 (N_7633,N_7360,N_7245);
xor U7634 (N_7634,N_7516,N_7382);
or U7635 (N_7635,N_7217,N_7383);
nand U7636 (N_7636,N_7307,N_7225);
and U7637 (N_7637,N_7487,N_7268);
and U7638 (N_7638,N_7599,N_7537);
nor U7639 (N_7639,N_7577,N_7525);
or U7640 (N_7640,N_7377,N_7564);
or U7641 (N_7641,N_7597,N_7498);
nand U7642 (N_7642,N_7448,N_7517);
nand U7643 (N_7643,N_7311,N_7293);
xnor U7644 (N_7644,N_7343,N_7214);
xnor U7645 (N_7645,N_7456,N_7261);
xnor U7646 (N_7646,N_7502,N_7403);
and U7647 (N_7647,N_7572,N_7240);
xnor U7648 (N_7648,N_7424,N_7406);
nand U7649 (N_7649,N_7468,N_7482);
xor U7650 (N_7650,N_7337,N_7238);
xor U7651 (N_7651,N_7381,N_7321);
nand U7652 (N_7652,N_7340,N_7461);
and U7653 (N_7653,N_7555,N_7302);
or U7654 (N_7654,N_7278,N_7541);
and U7655 (N_7655,N_7508,N_7255);
nand U7656 (N_7656,N_7290,N_7587);
nor U7657 (N_7657,N_7453,N_7292);
and U7658 (N_7658,N_7339,N_7466);
or U7659 (N_7659,N_7569,N_7348);
nor U7660 (N_7660,N_7551,N_7215);
xnor U7661 (N_7661,N_7454,N_7249);
nand U7662 (N_7662,N_7521,N_7423);
xnor U7663 (N_7663,N_7392,N_7437);
xor U7664 (N_7664,N_7559,N_7204);
nor U7665 (N_7665,N_7523,N_7446);
nand U7666 (N_7666,N_7390,N_7485);
xnor U7667 (N_7667,N_7530,N_7361);
or U7668 (N_7668,N_7414,N_7300);
xor U7669 (N_7669,N_7281,N_7344);
xnor U7670 (N_7670,N_7489,N_7288);
or U7671 (N_7671,N_7401,N_7439);
and U7672 (N_7672,N_7459,N_7318);
nor U7673 (N_7673,N_7202,N_7398);
or U7674 (N_7674,N_7419,N_7325);
nand U7675 (N_7675,N_7247,N_7547);
xor U7676 (N_7676,N_7550,N_7320);
nor U7677 (N_7677,N_7313,N_7330);
nor U7678 (N_7678,N_7442,N_7386);
or U7679 (N_7679,N_7370,N_7274);
nor U7680 (N_7680,N_7391,N_7428);
nor U7681 (N_7681,N_7529,N_7474);
xor U7682 (N_7682,N_7266,N_7396);
nand U7683 (N_7683,N_7315,N_7567);
nor U7684 (N_7684,N_7385,N_7504);
xor U7685 (N_7685,N_7409,N_7229);
and U7686 (N_7686,N_7515,N_7484);
nand U7687 (N_7687,N_7291,N_7251);
or U7688 (N_7688,N_7534,N_7262);
and U7689 (N_7689,N_7366,N_7368);
nor U7690 (N_7690,N_7440,N_7553);
nand U7691 (N_7691,N_7379,N_7560);
or U7692 (N_7692,N_7583,N_7380);
xnor U7693 (N_7693,N_7496,N_7248);
nor U7694 (N_7694,N_7510,N_7222);
nand U7695 (N_7695,N_7512,N_7542);
xnor U7696 (N_7696,N_7209,N_7477);
nor U7697 (N_7697,N_7438,N_7548);
or U7698 (N_7698,N_7455,N_7243);
nand U7699 (N_7699,N_7595,N_7239);
nor U7700 (N_7700,N_7533,N_7201);
xnor U7701 (N_7701,N_7479,N_7499);
xor U7702 (N_7702,N_7246,N_7579);
and U7703 (N_7703,N_7417,N_7354);
nand U7704 (N_7704,N_7467,N_7493);
and U7705 (N_7705,N_7465,N_7347);
nand U7706 (N_7706,N_7226,N_7444);
xor U7707 (N_7707,N_7388,N_7531);
and U7708 (N_7708,N_7208,N_7395);
nand U7709 (N_7709,N_7235,N_7205);
xor U7710 (N_7710,N_7257,N_7443);
nor U7711 (N_7711,N_7384,N_7480);
nor U7712 (N_7712,N_7303,N_7219);
and U7713 (N_7713,N_7279,N_7211);
or U7714 (N_7714,N_7509,N_7469);
nand U7715 (N_7715,N_7473,N_7236);
nor U7716 (N_7716,N_7230,N_7282);
and U7717 (N_7717,N_7349,N_7576);
nand U7718 (N_7718,N_7544,N_7332);
nand U7719 (N_7719,N_7399,N_7363);
nor U7720 (N_7720,N_7573,N_7258);
and U7721 (N_7721,N_7478,N_7408);
nor U7722 (N_7722,N_7232,N_7415);
and U7723 (N_7723,N_7492,N_7265);
xnor U7724 (N_7724,N_7260,N_7310);
and U7725 (N_7725,N_7270,N_7557);
or U7726 (N_7726,N_7322,N_7242);
nor U7727 (N_7727,N_7405,N_7367);
and U7728 (N_7728,N_7413,N_7472);
and U7729 (N_7729,N_7486,N_7341);
and U7730 (N_7730,N_7259,N_7284);
and U7731 (N_7731,N_7329,N_7346);
and U7732 (N_7732,N_7410,N_7206);
xor U7733 (N_7733,N_7210,N_7338);
nand U7734 (N_7734,N_7267,N_7511);
or U7735 (N_7735,N_7374,N_7524);
and U7736 (N_7736,N_7331,N_7237);
nand U7737 (N_7737,N_7527,N_7434);
xnor U7738 (N_7738,N_7543,N_7463);
and U7739 (N_7739,N_7327,N_7436);
and U7740 (N_7740,N_7269,N_7212);
or U7741 (N_7741,N_7221,N_7203);
and U7742 (N_7742,N_7430,N_7356);
or U7743 (N_7743,N_7596,N_7432);
or U7744 (N_7744,N_7425,N_7580);
xnor U7745 (N_7745,N_7317,N_7220);
or U7746 (N_7746,N_7200,N_7280);
and U7747 (N_7747,N_7526,N_7549);
xnor U7748 (N_7748,N_7224,N_7326);
xor U7749 (N_7749,N_7253,N_7213);
and U7750 (N_7750,N_7584,N_7421);
xor U7751 (N_7751,N_7593,N_7345);
nand U7752 (N_7752,N_7285,N_7563);
nand U7753 (N_7753,N_7540,N_7427);
nor U7754 (N_7754,N_7323,N_7252);
or U7755 (N_7755,N_7451,N_7566);
or U7756 (N_7756,N_7412,N_7264);
and U7757 (N_7757,N_7276,N_7445);
nand U7758 (N_7758,N_7362,N_7500);
xor U7759 (N_7759,N_7589,N_7207);
nor U7760 (N_7760,N_7334,N_7581);
nor U7761 (N_7761,N_7554,N_7590);
nor U7762 (N_7762,N_7433,N_7501);
nor U7763 (N_7763,N_7277,N_7299);
nor U7764 (N_7764,N_7452,N_7393);
and U7765 (N_7765,N_7256,N_7350);
and U7766 (N_7766,N_7552,N_7519);
xnor U7767 (N_7767,N_7295,N_7429);
xnor U7768 (N_7768,N_7271,N_7483);
and U7769 (N_7769,N_7556,N_7495);
nand U7770 (N_7770,N_7514,N_7546);
nand U7771 (N_7771,N_7364,N_7518);
or U7772 (N_7772,N_7294,N_7250);
nor U7773 (N_7773,N_7404,N_7372);
or U7774 (N_7774,N_7497,N_7416);
nand U7775 (N_7775,N_7488,N_7352);
and U7776 (N_7776,N_7309,N_7263);
nor U7777 (N_7777,N_7520,N_7574);
or U7778 (N_7778,N_7394,N_7335);
or U7779 (N_7779,N_7464,N_7312);
nand U7780 (N_7780,N_7422,N_7228);
xnor U7781 (N_7781,N_7571,N_7558);
nand U7782 (N_7782,N_7431,N_7353);
and U7783 (N_7783,N_7316,N_7460);
and U7784 (N_7784,N_7314,N_7357);
nor U7785 (N_7785,N_7387,N_7582);
nor U7786 (N_7786,N_7585,N_7562);
and U7787 (N_7787,N_7241,N_7358);
and U7788 (N_7788,N_7328,N_7373);
or U7789 (N_7789,N_7296,N_7591);
xnor U7790 (N_7790,N_7223,N_7505);
nor U7791 (N_7791,N_7598,N_7545);
xor U7792 (N_7792,N_7426,N_7441);
or U7793 (N_7793,N_7535,N_7490);
xnor U7794 (N_7794,N_7594,N_7319);
and U7795 (N_7795,N_7231,N_7397);
and U7796 (N_7796,N_7369,N_7507);
nor U7797 (N_7797,N_7297,N_7450);
and U7798 (N_7798,N_7308,N_7218);
nand U7799 (N_7799,N_7592,N_7351);
xor U7800 (N_7800,N_7412,N_7319);
nor U7801 (N_7801,N_7281,N_7407);
nor U7802 (N_7802,N_7384,N_7292);
nand U7803 (N_7803,N_7422,N_7262);
nand U7804 (N_7804,N_7450,N_7548);
nand U7805 (N_7805,N_7513,N_7413);
xor U7806 (N_7806,N_7335,N_7233);
nor U7807 (N_7807,N_7226,N_7377);
nor U7808 (N_7808,N_7212,N_7508);
xor U7809 (N_7809,N_7459,N_7474);
and U7810 (N_7810,N_7576,N_7244);
xnor U7811 (N_7811,N_7269,N_7348);
xor U7812 (N_7812,N_7227,N_7217);
or U7813 (N_7813,N_7306,N_7514);
and U7814 (N_7814,N_7336,N_7215);
nor U7815 (N_7815,N_7303,N_7368);
nor U7816 (N_7816,N_7442,N_7328);
and U7817 (N_7817,N_7201,N_7588);
xor U7818 (N_7818,N_7292,N_7559);
nor U7819 (N_7819,N_7527,N_7381);
or U7820 (N_7820,N_7513,N_7268);
or U7821 (N_7821,N_7305,N_7211);
and U7822 (N_7822,N_7418,N_7301);
and U7823 (N_7823,N_7302,N_7513);
and U7824 (N_7824,N_7596,N_7518);
nand U7825 (N_7825,N_7398,N_7368);
xnor U7826 (N_7826,N_7228,N_7580);
nand U7827 (N_7827,N_7366,N_7475);
or U7828 (N_7828,N_7211,N_7351);
nor U7829 (N_7829,N_7572,N_7484);
and U7830 (N_7830,N_7507,N_7477);
nand U7831 (N_7831,N_7368,N_7257);
or U7832 (N_7832,N_7524,N_7248);
or U7833 (N_7833,N_7341,N_7373);
or U7834 (N_7834,N_7470,N_7519);
xor U7835 (N_7835,N_7576,N_7491);
and U7836 (N_7836,N_7367,N_7400);
nand U7837 (N_7837,N_7476,N_7562);
nand U7838 (N_7838,N_7525,N_7252);
or U7839 (N_7839,N_7435,N_7359);
or U7840 (N_7840,N_7377,N_7473);
nand U7841 (N_7841,N_7361,N_7585);
nor U7842 (N_7842,N_7259,N_7309);
or U7843 (N_7843,N_7390,N_7303);
xor U7844 (N_7844,N_7584,N_7269);
or U7845 (N_7845,N_7563,N_7502);
and U7846 (N_7846,N_7388,N_7439);
nor U7847 (N_7847,N_7365,N_7371);
nor U7848 (N_7848,N_7589,N_7201);
nand U7849 (N_7849,N_7575,N_7290);
nor U7850 (N_7850,N_7523,N_7225);
nand U7851 (N_7851,N_7445,N_7462);
nor U7852 (N_7852,N_7216,N_7341);
or U7853 (N_7853,N_7589,N_7496);
nand U7854 (N_7854,N_7586,N_7338);
nand U7855 (N_7855,N_7293,N_7586);
xnor U7856 (N_7856,N_7467,N_7541);
nand U7857 (N_7857,N_7449,N_7582);
nor U7858 (N_7858,N_7421,N_7262);
nor U7859 (N_7859,N_7512,N_7321);
or U7860 (N_7860,N_7532,N_7581);
nand U7861 (N_7861,N_7522,N_7515);
nor U7862 (N_7862,N_7419,N_7497);
nand U7863 (N_7863,N_7497,N_7484);
xor U7864 (N_7864,N_7598,N_7215);
xnor U7865 (N_7865,N_7212,N_7330);
nor U7866 (N_7866,N_7463,N_7416);
nor U7867 (N_7867,N_7526,N_7208);
nand U7868 (N_7868,N_7477,N_7510);
nor U7869 (N_7869,N_7343,N_7312);
nand U7870 (N_7870,N_7581,N_7257);
xor U7871 (N_7871,N_7343,N_7423);
xor U7872 (N_7872,N_7375,N_7214);
xnor U7873 (N_7873,N_7247,N_7282);
or U7874 (N_7874,N_7560,N_7530);
nor U7875 (N_7875,N_7363,N_7550);
nor U7876 (N_7876,N_7368,N_7417);
xnor U7877 (N_7877,N_7556,N_7470);
xnor U7878 (N_7878,N_7235,N_7276);
xnor U7879 (N_7879,N_7472,N_7215);
and U7880 (N_7880,N_7570,N_7434);
nor U7881 (N_7881,N_7220,N_7408);
xor U7882 (N_7882,N_7292,N_7343);
nor U7883 (N_7883,N_7583,N_7540);
and U7884 (N_7884,N_7339,N_7597);
nor U7885 (N_7885,N_7524,N_7390);
and U7886 (N_7886,N_7437,N_7501);
nand U7887 (N_7887,N_7573,N_7410);
xnor U7888 (N_7888,N_7585,N_7428);
or U7889 (N_7889,N_7271,N_7396);
xnor U7890 (N_7890,N_7289,N_7383);
nand U7891 (N_7891,N_7346,N_7434);
and U7892 (N_7892,N_7546,N_7517);
and U7893 (N_7893,N_7581,N_7249);
nor U7894 (N_7894,N_7515,N_7391);
nand U7895 (N_7895,N_7534,N_7409);
and U7896 (N_7896,N_7247,N_7320);
or U7897 (N_7897,N_7277,N_7322);
or U7898 (N_7898,N_7471,N_7386);
or U7899 (N_7899,N_7411,N_7547);
and U7900 (N_7900,N_7566,N_7427);
and U7901 (N_7901,N_7504,N_7531);
xnor U7902 (N_7902,N_7306,N_7311);
xnor U7903 (N_7903,N_7458,N_7317);
nor U7904 (N_7904,N_7237,N_7383);
nor U7905 (N_7905,N_7353,N_7560);
or U7906 (N_7906,N_7245,N_7394);
or U7907 (N_7907,N_7292,N_7484);
or U7908 (N_7908,N_7292,N_7370);
xor U7909 (N_7909,N_7451,N_7580);
xnor U7910 (N_7910,N_7500,N_7332);
nor U7911 (N_7911,N_7530,N_7566);
and U7912 (N_7912,N_7409,N_7546);
xnor U7913 (N_7913,N_7203,N_7228);
nand U7914 (N_7914,N_7321,N_7561);
nor U7915 (N_7915,N_7380,N_7273);
or U7916 (N_7916,N_7303,N_7550);
xnor U7917 (N_7917,N_7339,N_7250);
xor U7918 (N_7918,N_7213,N_7228);
nand U7919 (N_7919,N_7200,N_7498);
xor U7920 (N_7920,N_7488,N_7461);
nor U7921 (N_7921,N_7595,N_7542);
nand U7922 (N_7922,N_7557,N_7418);
and U7923 (N_7923,N_7401,N_7527);
nor U7924 (N_7924,N_7359,N_7552);
and U7925 (N_7925,N_7410,N_7346);
nand U7926 (N_7926,N_7470,N_7413);
or U7927 (N_7927,N_7447,N_7231);
nand U7928 (N_7928,N_7559,N_7359);
and U7929 (N_7929,N_7311,N_7404);
xnor U7930 (N_7930,N_7350,N_7432);
nand U7931 (N_7931,N_7469,N_7236);
or U7932 (N_7932,N_7362,N_7481);
nor U7933 (N_7933,N_7376,N_7268);
nor U7934 (N_7934,N_7390,N_7405);
xnor U7935 (N_7935,N_7551,N_7311);
or U7936 (N_7936,N_7267,N_7239);
nor U7937 (N_7937,N_7238,N_7558);
xor U7938 (N_7938,N_7585,N_7528);
xor U7939 (N_7939,N_7466,N_7352);
xor U7940 (N_7940,N_7398,N_7470);
nand U7941 (N_7941,N_7417,N_7521);
and U7942 (N_7942,N_7474,N_7342);
nor U7943 (N_7943,N_7456,N_7311);
xor U7944 (N_7944,N_7575,N_7477);
or U7945 (N_7945,N_7467,N_7451);
nand U7946 (N_7946,N_7312,N_7541);
or U7947 (N_7947,N_7276,N_7588);
nand U7948 (N_7948,N_7278,N_7284);
nand U7949 (N_7949,N_7463,N_7329);
xor U7950 (N_7950,N_7589,N_7570);
and U7951 (N_7951,N_7534,N_7515);
and U7952 (N_7952,N_7212,N_7243);
nor U7953 (N_7953,N_7268,N_7385);
or U7954 (N_7954,N_7495,N_7336);
or U7955 (N_7955,N_7583,N_7582);
xnor U7956 (N_7956,N_7422,N_7536);
and U7957 (N_7957,N_7287,N_7396);
nor U7958 (N_7958,N_7368,N_7330);
or U7959 (N_7959,N_7327,N_7467);
nand U7960 (N_7960,N_7257,N_7375);
xor U7961 (N_7961,N_7310,N_7539);
nor U7962 (N_7962,N_7447,N_7576);
nor U7963 (N_7963,N_7449,N_7299);
nand U7964 (N_7964,N_7518,N_7356);
nor U7965 (N_7965,N_7566,N_7308);
and U7966 (N_7966,N_7296,N_7561);
or U7967 (N_7967,N_7205,N_7575);
xor U7968 (N_7968,N_7541,N_7508);
or U7969 (N_7969,N_7497,N_7205);
or U7970 (N_7970,N_7366,N_7293);
nor U7971 (N_7971,N_7345,N_7458);
and U7972 (N_7972,N_7377,N_7462);
nor U7973 (N_7973,N_7547,N_7264);
nand U7974 (N_7974,N_7214,N_7335);
xor U7975 (N_7975,N_7320,N_7422);
nand U7976 (N_7976,N_7316,N_7436);
and U7977 (N_7977,N_7334,N_7455);
nand U7978 (N_7978,N_7578,N_7358);
xnor U7979 (N_7979,N_7459,N_7267);
nor U7980 (N_7980,N_7432,N_7394);
nor U7981 (N_7981,N_7571,N_7280);
or U7982 (N_7982,N_7202,N_7537);
nand U7983 (N_7983,N_7208,N_7472);
nor U7984 (N_7984,N_7332,N_7412);
and U7985 (N_7985,N_7558,N_7331);
nand U7986 (N_7986,N_7507,N_7230);
and U7987 (N_7987,N_7308,N_7423);
xnor U7988 (N_7988,N_7580,N_7532);
xnor U7989 (N_7989,N_7201,N_7527);
nor U7990 (N_7990,N_7393,N_7309);
or U7991 (N_7991,N_7245,N_7500);
and U7992 (N_7992,N_7314,N_7447);
and U7993 (N_7993,N_7212,N_7325);
nand U7994 (N_7994,N_7430,N_7475);
and U7995 (N_7995,N_7246,N_7565);
and U7996 (N_7996,N_7432,N_7487);
and U7997 (N_7997,N_7203,N_7213);
nor U7998 (N_7998,N_7424,N_7582);
nand U7999 (N_7999,N_7305,N_7203);
xor U8000 (N_8000,N_7620,N_7864);
and U8001 (N_8001,N_7905,N_7872);
xnor U8002 (N_8002,N_7873,N_7849);
nor U8003 (N_8003,N_7800,N_7975);
xnor U8004 (N_8004,N_7831,N_7633);
xor U8005 (N_8005,N_7763,N_7867);
nor U8006 (N_8006,N_7928,N_7866);
and U8007 (N_8007,N_7755,N_7945);
nor U8008 (N_8008,N_7639,N_7699);
nand U8009 (N_8009,N_7923,N_7891);
or U8010 (N_8010,N_7992,N_7666);
xor U8011 (N_8011,N_7935,N_7914);
nor U8012 (N_8012,N_7931,N_7819);
and U8013 (N_8013,N_7895,N_7957);
or U8014 (N_8014,N_7762,N_7893);
xnor U8015 (N_8015,N_7690,N_7732);
nand U8016 (N_8016,N_7847,N_7616);
nor U8017 (N_8017,N_7653,N_7841);
xor U8018 (N_8018,N_7997,N_7939);
xnor U8019 (N_8019,N_7718,N_7824);
xor U8020 (N_8020,N_7792,N_7920);
or U8021 (N_8021,N_7960,N_7746);
and U8022 (N_8022,N_7742,N_7959);
and U8023 (N_8023,N_7936,N_7919);
xnor U8024 (N_8024,N_7693,N_7838);
xor U8025 (N_8025,N_7725,N_7686);
and U8026 (N_8026,N_7978,N_7877);
nor U8027 (N_8027,N_7655,N_7783);
and U8028 (N_8028,N_7603,N_7683);
or U8029 (N_8029,N_7940,N_7818);
xor U8030 (N_8030,N_7840,N_7708);
nand U8031 (N_8031,N_7759,N_7716);
nand U8032 (N_8032,N_7662,N_7853);
nor U8033 (N_8033,N_7617,N_7672);
nor U8034 (N_8034,N_7779,N_7976);
xor U8035 (N_8035,N_7932,N_7794);
nand U8036 (N_8036,N_7697,N_7613);
nor U8037 (N_8037,N_7814,N_7711);
nor U8038 (N_8038,N_7651,N_7869);
nand U8039 (N_8039,N_7785,N_7791);
nand U8040 (N_8040,N_7680,N_7937);
nor U8041 (N_8041,N_7607,N_7644);
nor U8042 (N_8042,N_7989,N_7868);
or U8043 (N_8043,N_7946,N_7861);
nand U8044 (N_8044,N_7676,N_7769);
xor U8045 (N_8045,N_7990,N_7605);
nor U8046 (N_8046,N_7634,N_7715);
nor U8047 (N_8047,N_7974,N_7828);
nand U8048 (N_8048,N_7961,N_7925);
and U8049 (N_8049,N_7646,N_7906);
nand U8050 (N_8050,N_7952,N_7878);
nor U8051 (N_8051,N_7816,N_7904);
nand U8052 (N_8052,N_7745,N_7956);
nand U8053 (N_8053,N_7773,N_7832);
nand U8054 (N_8054,N_7630,N_7740);
and U8055 (N_8055,N_7885,N_7736);
and U8056 (N_8056,N_7695,N_7691);
and U8057 (N_8057,N_7750,N_7684);
nor U8058 (N_8058,N_7770,N_7670);
and U8059 (N_8059,N_7747,N_7907);
nor U8060 (N_8060,N_7739,N_7806);
or U8061 (N_8061,N_7752,N_7979);
xnor U8062 (N_8062,N_7821,N_7850);
xor U8063 (N_8063,N_7805,N_7766);
xnor U8064 (N_8064,N_7884,N_7900);
nor U8065 (N_8065,N_7793,N_7733);
nand U8066 (N_8066,N_7823,N_7614);
xnor U8067 (N_8067,N_7727,N_7916);
xor U8068 (N_8068,N_7656,N_7689);
nand U8069 (N_8069,N_7668,N_7826);
and U8070 (N_8070,N_7704,N_7765);
nor U8071 (N_8071,N_7811,N_7846);
nand U8072 (N_8072,N_7921,N_7882);
xor U8073 (N_8073,N_7784,N_7659);
and U8074 (N_8074,N_7910,N_7848);
xor U8075 (N_8075,N_7851,N_7942);
nor U8076 (N_8076,N_7835,N_7673);
xnor U8077 (N_8077,N_7741,N_7754);
and U8078 (N_8078,N_7641,N_7774);
nand U8079 (N_8079,N_7981,N_7692);
xor U8080 (N_8080,N_7901,N_7638);
or U8081 (N_8081,N_7751,N_7610);
nor U8082 (N_8082,N_7650,N_7721);
nor U8083 (N_8083,N_7949,N_7714);
nor U8084 (N_8084,N_7637,N_7862);
xor U8085 (N_8085,N_7764,N_7631);
and U8086 (N_8086,N_7999,N_7667);
nor U8087 (N_8087,N_7609,N_7812);
and U8088 (N_8088,N_7606,N_7748);
and U8089 (N_8089,N_7898,N_7772);
nor U8090 (N_8090,N_7988,N_7758);
and U8091 (N_8091,N_7643,N_7948);
and U8092 (N_8092,N_7894,N_7665);
nor U8093 (N_8093,N_7694,N_7790);
or U8094 (N_8094,N_7788,N_7970);
nor U8095 (N_8095,N_7991,N_7971);
nand U8096 (N_8096,N_7782,N_7687);
nand U8097 (N_8097,N_7839,N_7664);
nand U8098 (N_8098,N_7701,N_7685);
or U8099 (N_8099,N_7982,N_7930);
and U8100 (N_8100,N_7833,N_7863);
nand U8101 (N_8101,N_7705,N_7911);
and U8102 (N_8102,N_7967,N_7852);
nor U8103 (N_8103,N_7780,N_7844);
or U8104 (N_8104,N_7843,N_7608);
or U8105 (N_8105,N_7632,N_7657);
or U8106 (N_8106,N_7767,N_7623);
xnor U8107 (N_8107,N_7600,N_7749);
and U8108 (N_8108,N_7830,N_7756);
xor U8109 (N_8109,N_7724,N_7677);
and U8110 (N_8110,N_7985,N_7887);
xnor U8111 (N_8111,N_7886,N_7880);
or U8112 (N_8112,N_7728,N_7778);
xor U8113 (N_8113,N_7915,N_7744);
or U8114 (N_8114,N_7965,N_7652);
and U8115 (N_8115,N_7856,N_7604);
xor U8116 (N_8116,N_7809,N_7980);
or U8117 (N_8117,N_7696,N_7753);
nor U8118 (N_8118,N_7698,N_7996);
nor U8119 (N_8119,N_7817,N_7836);
xnor U8120 (N_8120,N_7803,N_7682);
nor U8121 (N_8121,N_7934,N_7629);
nand U8122 (N_8122,N_7987,N_7660);
and U8123 (N_8123,N_7938,N_7776);
or U8124 (N_8124,N_7624,N_7781);
and U8125 (N_8125,N_7743,N_7615);
or U8126 (N_8126,N_7890,N_7902);
or U8127 (N_8127,N_7734,N_7947);
nand U8128 (N_8128,N_7892,N_7969);
xnor U8129 (N_8129,N_7963,N_7797);
nor U8130 (N_8130,N_7897,N_7717);
nor U8131 (N_8131,N_7827,N_7825);
nand U8132 (N_8132,N_7801,N_7927);
xor U8133 (N_8133,N_7888,N_7998);
nor U8134 (N_8134,N_7966,N_7729);
xnor U8135 (N_8135,N_7899,N_7913);
or U8136 (N_8136,N_7757,N_7995);
or U8137 (N_8137,N_7918,N_7889);
nand U8138 (N_8138,N_7972,N_7964);
nor U8139 (N_8139,N_7875,N_7908);
or U8140 (N_8140,N_7700,N_7955);
or U8141 (N_8141,N_7738,N_7786);
xnor U8142 (N_8142,N_7671,N_7903);
nand U8143 (N_8143,N_7645,N_7883);
or U8144 (N_8144,N_7636,N_7619);
xor U8145 (N_8145,N_7973,N_7612);
nand U8146 (N_8146,N_7787,N_7611);
or U8147 (N_8147,N_7775,N_7761);
and U8148 (N_8148,N_7760,N_7663);
nand U8149 (N_8149,N_7768,N_7720);
nor U8150 (N_8150,N_7829,N_7820);
nand U8151 (N_8151,N_7771,N_7621);
nand U8152 (N_8152,N_7986,N_7661);
nand U8153 (N_8153,N_7628,N_7926);
nand U8154 (N_8154,N_7710,N_7706);
or U8155 (N_8155,N_7702,N_7879);
nand U8156 (N_8156,N_7625,N_7719);
xor U8157 (N_8157,N_7804,N_7834);
nor U8158 (N_8158,N_7941,N_7722);
or U8159 (N_8159,N_7822,N_7648);
or U8160 (N_8160,N_7713,N_7675);
nor U8161 (N_8161,N_7924,N_7807);
and U8162 (N_8162,N_7654,N_7922);
or U8163 (N_8163,N_7601,N_7896);
xor U8164 (N_8164,N_7796,N_7627);
nor U8165 (N_8165,N_7837,N_7602);
nand U8166 (N_8166,N_7993,N_7865);
nand U8167 (N_8167,N_7789,N_7626);
or U8168 (N_8168,N_7968,N_7912);
xor U8169 (N_8169,N_7799,N_7635);
nand U8170 (N_8170,N_7953,N_7802);
and U8171 (N_8171,N_7707,N_7813);
xnor U8172 (N_8172,N_7798,N_7735);
nor U8173 (N_8173,N_7712,N_7669);
nand U8174 (N_8174,N_7723,N_7983);
xnor U8175 (N_8175,N_7870,N_7681);
nand U8176 (N_8176,N_7958,N_7854);
nor U8177 (N_8177,N_7954,N_7950);
or U8178 (N_8178,N_7703,N_7917);
xnor U8179 (N_8179,N_7929,N_7859);
xnor U8180 (N_8180,N_7709,N_7777);
and U8181 (N_8181,N_7881,N_7649);
or U8182 (N_8182,N_7808,N_7951);
or U8183 (N_8183,N_7731,N_7730);
and U8184 (N_8184,N_7857,N_7994);
xnor U8185 (N_8185,N_7944,N_7647);
xnor U8186 (N_8186,N_7876,N_7726);
nand U8187 (N_8187,N_7943,N_7984);
nor U8188 (N_8188,N_7860,N_7658);
nand U8189 (N_8189,N_7810,N_7977);
or U8190 (N_8190,N_7688,N_7842);
nand U8191 (N_8191,N_7737,N_7933);
and U8192 (N_8192,N_7845,N_7871);
nand U8193 (N_8193,N_7874,N_7622);
nor U8194 (N_8194,N_7642,N_7795);
or U8195 (N_8195,N_7855,N_7674);
nand U8196 (N_8196,N_7962,N_7679);
nor U8197 (N_8197,N_7640,N_7618);
nand U8198 (N_8198,N_7815,N_7678);
and U8199 (N_8199,N_7909,N_7858);
and U8200 (N_8200,N_7998,N_7892);
and U8201 (N_8201,N_7600,N_7674);
or U8202 (N_8202,N_7738,N_7676);
xor U8203 (N_8203,N_7663,N_7753);
nand U8204 (N_8204,N_7859,N_7987);
nand U8205 (N_8205,N_7774,N_7865);
nor U8206 (N_8206,N_7777,N_7941);
xor U8207 (N_8207,N_7716,N_7848);
or U8208 (N_8208,N_7895,N_7997);
nor U8209 (N_8209,N_7623,N_7862);
nor U8210 (N_8210,N_7946,N_7910);
or U8211 (N_8211,N_7986,N_7724);
xor U8212 (N_8212,N_7852,N_7777);
or U8213 (N_8213,N_7882,N_7812);
xor U8214 (N_8214,N_7895,N_7870);
and U8215 (N_8215,N_7880,N_7689);
xnor U8216 (N_8216,N_7673,N_7907);
nor U8217 (N_8217,N_7718,N_7807);
or U8218 (N_8218,N_7917,N_7603);
and U8219 (N_8219,N_7918,N_7969);
nand U8220 (N_8220,N_7688,N_7930);
or U8221 (N_8221,N_7669,N_7865);
nand U8222 (N_8222,N_7965,N_7877);
and U8223 (N_8223,N_7745,N_7969);
nor U8224 (N_8224,N_7607,N_7816);
nand U8225 (N_8225,N_7608,N_7756);
nor U8226 (N_8226,N_7844,N_7920);
xnor U8227 (N_8227,N_7605,N_7741);
nand U8228 (N_8228,N_7755,N_7999);
xnor U8229 (N_8229,N_7985,N_7735);
and U8230 (N_8230,N_7670,N_7769);
nand U8231 (N_8231,N_7942,N_7960);
or U8232 (N_8232,N_7824,N_7659);
and U8233 (N_8233,N_7677,N_7873);
and U8234 (N_8234,N_7826,N_7920);
or U8235 (N_8235,N_7927,N_7735);
xor U8236 (N_8236,N_7870,N_7818);
and U8237 (N_8237,N_7857,N_7730);
and U8238 (N_8238,N_7718,N_7828);
xor U8239 (N_8239,N_7777,N_7992);
xnor U8240 (N_8240,N_7887,N_7880);
nor U8241 (N_8241,N_7629,N_7794);
or U8242 (N_8242,N_7726,N_7829);
xor U8243 (N_8243,N_7652,N_7618);
and U8244 (N_8244,N_7725,N_7653);
or U8245 (N_8245,N_7743,N_7963);
nand U8246 (N_8246,N_7782,N_7749);
and U8247 (N_8247,N_7682,N_7937);
and U8248 (N_8248,N_7901,N_7775);
nor U8249 (N_8249,N_7967,N_7894);
xor U8250 (N_8250,N_7852,N_7751);
nor U8251 (N_8251,N_7676,N_7681);
nor U8252 (N_8252,N_7954,N_7766);
and U8253 (N_8253,N_7940,N_7769);
nand U8254 (N_8254,N_7729,N_7830);
xor U8255 (N_8255,N_7724,N_7977);
nand U8256 (N_8256,N_7769,N_7975);
nand U8257 (N_8257,N_7667,N_7861);
or U8258 (N_8258,N_7887,N_7834);
or U8259 (N_8259,N_7968,N_7845);
nand U8260 (N_8260,N_7996,N_7622);
or U8261 (N_8261,N_7833,N_7929);
or U8262 (N_8262,N_7704,N_7809);
or U8263 (N_8263,N_7612,N_7671);
nor U8264 (N_8264,N_7725,N_7611);
and U8265 (N_8265,N_7722,N_7886);
xor U8266 (N_8266,N_7760,N_7610);
and U8267 (N_8267,N_7634,N_7994);
or U8268 (N_8268,N_7708,N_7998);
and U8269 (N_8269,N_7612,N_7953);
nand U8270 (N_8270,N_7959,N_7769);
and U8271 (N_8271,N_7690,N_7701);
xor U8272 (N_8272,N_7932,N_7631);
nand U8273 (N_8273,N_7960,N_7766);
xor U8274 (N_8274,N_7967,N_7778);
xor U8275 (N_8275,N_7922,N_7636);
nor U8276 (N_8276,N_7979,N_7967);
xnor U8277 (N_8277,N_7635,N_7898);
nor U8278 (N_8278,N_7920,N_7655);
nand U8279 (N_8279,N_7606,N_7616);
nor U8280 (N_8280,N_7989,N_7741);
xor U8281 (N_8281,N_7944,N_7936);
nand U8282 (N_8282,N_7997,N_7662);
and U8283 (N_8283,N_7853,N_7627);
xor U8284 (N_8284,N_7936,N_7866);
nor U8285 (N_8285,N_7981,N_7887);
xor U8286 (N_8286,N_7865,N_7766);
or U8287 (N_8287,N_7808,N_7867);
xor U8288 (N_8288,N_7811,N_7701);
or U8289 (N_8289,N_7677,N_7995);
xnor U8290 (N_8290,N_7958,N_7846);
nor U8291 (N_8291,N_7867,N_7620);
nor U8292 (N_8292,N_7960,N_7721);
nand U8293 (N_8293,N_7840,N_7636);
xor U8294 (N_8294,N_7678,N_7970);
and U8295 (N_8295,N_7888,N_7742);
or U8296 (N_8296,N_7848,N_7968);
nor U8297 (N_8297,N_7903,N_7800);
and U8298 (N_8298,N_7772,N_7639);
and U8299 (N_8299,N_7929,N_7730);
or U8300 (N_8300,N_7851,N_7779);
or U8301 (N_8301,N_7703,N_7850);
nand U8302 (N_8302,N_7644,N_7770);
nand U8303 (N_8303,N_7739,N_7619);
or U8304 (N_8304,N_7674,N_7896);
nand U8305 (N_8305,N_7991,N_7849);
and U8306 (N_8306,N_7742,N_7866);
nand U8307 (N_8307,N_7602,N_7685);
nor U8308 (N_8308,N_7921,N_7672);
or U8309 (N_8309,N_7753,N_7839);
and U8310 (N_8310,N_7999,N_7728);
nand U8311 (N_8311,N_7763,N_7945);
and U8312 (N_8312,N_7961,N_7910);
xnor U8313 (N_8313,N_7865,N_7782);
xor U8314 (N_8314,N_7762,N_7998);
xnor U8315 (N_8315,N_7720,N_7845);
and U8316 (N_8316,N_7895,N_7754);
nand U8317 (N_8317,N_7645,N_7784);
or U8318 (N_8318,N_7812,N_7714);
nand U8319 (N_8319,N_7866,N_7899);
nand U8320 (N_8320,N_7833,N_7832);
nand U8321 (N_8321,N_7718,N_7744);
xor U8322 (N_8322,N_7671,N_7840);
and U8323 (N_8323,N_7695,N_7651);
nand U8324 (N_8324,N_7870,N_7893);
or U8325 (N_8325,N_7648,N_7736);
or U8326 (N_8326,N_7642,N_7961);
nand U8327 (N_8327,N_7912,N_7678);
or U8328 (N_8328,N_7823,N_7865);
nand U8329 (N_8329,N_7685,N_7615);
or U8330 (N_8330,N_7959,N_7680);
xor U8331 (N_8331,N_7790,N_7638);
nor U8332 (N_8332,N_7918,N_7956);
or U8333 (N_8333,N_7633,N_7860);
nand U8334 (N_8334,N_7965,N_7916);
nand U8335 (N_8335,N_7861,N_7819);
and U8336 (N_8336,N_7831,N_7734);
xnor U8337 (N_8337,N_7784,N_7603);
nor U8338 (N_8338,N_7788,N_7605);
and U8339 (N_8339,N_7879,N_7884);
xor U8340 (N_8340,N_7608,N_7619);
xor U8341 (N_8341,N_7988,N_7846);
nand U8342 (N_8342,N_7882,N_7850);
xor U8343 (N_8343,N_7685,N_7934);
nor U8344 (N_8344,N_7702,N_7885);
or U8345 (N_8345,N_7676,N_7987);
or U8346 (N_8346,N_7703,N_7712);
xnor U8347 (N_8347,N_7974,N_7943);
and U8348 (N_8348,N_7958,N_7730);
xnor U8349 (N_8349,N_7971,N_7734);
nand U8350 (N_8350,N_7982,N_7910);
nand U8351 (N_8351,N_7971,N_7895);
or U8352 (N_8352,N_7927,N_7781);
and U8353 (N_8353,N_7898,N_7785);
xor U8354 (N_8354,N_7750,N_7902);
and U8355 (N_8355,N_7683,N_7860);
nor U8356 (N_8356,N_7606,N_7882);
and U8357 (N_8357,N_7880,N_7996);
or U8358 (N_8358,N_7654,N_7955);
nand U8359 (N_8359,N_7826,N_7731);
nor U8360 (N_8360,N_7942,N_7679);
nor U8361 (N_8361,N_7907,N_7802);
xnor U8362 (N_8362,N_7878,N_7688);
and U8363 (N_8363,N_7823,N_7825);
and U8364 (N_8364,N_7889,N_7642);
nor U8365 (N_8365,N_7766,N_7681);
and U8366 (N_8366,N_7665,N_7664);
nand U8367 (N_8367,N_7744,N_7740);
or U8368 (N_8368,N_7780,N_7662);
and U8369 (N_8369,N_7922,N_7874);
xnor U8370 (N_8370,N_7707,N_7724);
or U8371 (N_8371,N_7982,N_7953);
nand U8372 (N_8372,N_7702,N_7716);
nand U8373 (N_8373,N_7883,N_7632);
or U8374 (N_8374,N_7814,N_7866);
and U8375 (N_8375,N_7790,N_7951);
xnor U8376 (N_8376,N_7747,N_7899);
or U8377 (N_8377,N_7602,N_7788);
and U8378 (N_8378,N_7866,N_7830);
nand U8379 (N_8379,N_7811,N_7800);
xor U8380 (N_8380,N_7909,N_7985);
or U8381 (N_8381,N_7894,N_7712);
and U8382 (N_8382,N_7812,N_7933);
xnor U8383 (N_8383,N_7769,N_7817);
xnor U8384 (N_8384,N_7892,N_7625);
nand U8385 (N_8385,N_7736,N_7618);
nand U8386 (N_8386,N_7877,N_7884);
nand U8387 (N_8387,N_7990,N_7834);
nand U8388 (N_8388,N_7820,N_7738);
or U8389 (N_8389,N_7687,N_7984);
and U8390 (N_8390,N_7612,N_7976);
nor U8391 (N_8391,N_7921,N_7910);
or U8392 (N_8392,N_7875,N_7792);
nand U8393 (N_8393,N_7693,N_7942);
nand U8394 (N_8394,N_7749,N_7890);
nand U8395 (N_8395,N_7696,N_7899);
xnor U8396 (N_8396,N_7631,N_7783);
or U8397 (N_8397,N_7877,N_7890);
or U8398 (N_8398,N_7929,N_7664);
or U8399 (N_8399,N_7895,N_7992);
xor U8400 (N_8400,N_8142,N_8305);
xor U8401 (N_8401,N_8124,N_8211);
xnor U8402 (N_8402,N_8369,N_8182);
nand U8403 (N_8403,N_8028,N_8014);
nor U8404 (N_8404,N_8339,N_8390);
xnor U8405 (N_8405,N_8396,N_8303);
and U8406 (N_8406,N_8131,N_8040);
and U8407 (N_8407,N_8372,N_8016);
nor U8408 (N_8408,N_8105,N_8132);
and U8409 (N_8409,N_8378,N_8264);
nor U8410 (N_8410,N_8302,N_8139);
or U8411 (N_8411,N_8000,N_8152);
and U8412 (N_8412,N_8329,N_8256);
xnor U8413 (N_8413,N_8135,N_8147);
nor U8414 (N_8414,N_8104,N_8384);
nand U8415 (N_8415,N_8265,N_8338);
or U8416 (N_8416,N_8349,N_8365);
nor U8417 (N_8417,N_8165,N_8312);
and U8418 (N_8418,N_8291,N_8190);
nand U8419 (N_8419,N_8207,N_8314);
nand U8420 (N_8420,N_8065,N_8119);
nor U8421 (N_8421,N_8184,N_8259);
and U8422 (N_8422,N_8111,N_8382);
xor U8423 (N_8423,N_8177,N_8084);
nor U8424 (N_8424,N_8304,N_8148);
nor U8425 (N_8425,N_8234,N_8230);
and U8426 (N_8426,N_8068,N_8006);
and U8427 (N_8427,N_8330,N_8261);
and U8428 (N_8428,N_8392,N_8081);
or U8429 (N_8429,N_8101,N_8073);
xor U8430 (N_8430,N_8140,N_8160);
or U8431 (N_8431,N_8394,N_8025);
and U8432 (N_8432,N_8150,N_8244);
and U8433 (N_8433,N_8385,N_8285);
xor U8434 (N_8434,N_8026,N_8062);
or U8435 (N_8435,N_8080,N_8018);
nor U8436 (N_8436,N_8227,N_8275);
nor U8437 (N_8437,N_8094,N_8398);
or U8438 (N_8438,N_8309,N_8192);
xnor U8439 (N_8439,N_8043,N_8120);
and U8440 (N_8440,N_8168,N_8308);
nor U8441 (N_8441,N_8173,N_8118);
nor U8442 (N_8442,N_8301,N_8255);
nor U8443 (N_8443,N_8219,N_8056);
xnor U8444 (N_8444,N_8097,N_8313);
nand U8445 (N_8445,N_8074,N_8204);
nand U8446 (N_8446,N_8045,N_8052);
or U8447 (N_8447,N_8186,N_8248);
or U8448 (N_8448,N_8343,N_8214);
nor U8449 (N_8449,N_8237,N_8373);
or U8450 (N_8450,N_8166,N_8281);
xor U8451 (N_8451,N_8138,N_8141);
xnor U8452 (N_8452,N_8159,N_8370);
and U8453 (N_8453,N_8143,N_8051);
and U8454 (N_8454,N_8079,N_8027);
or U8455 (N_8455,N_8042,N_8247);
nor U8456 (N_8456,N_8245,N_8151);
xnor U8457 (N_8457,N_8164,N_8125);
or U8458 (N_8458,N_8335,N_8321);
nor U8459 (N_8459,N_8034,N_8108);
nand U8460 (N_8460,N_8274,N_8181);
and U8461 (N_8461,N_8171,N_8146);
and U8462 (N_8462,N_8049,N_8300);
and U8463 (N_8463,N_8257,N_8235);
nor U8464 (N_8464,N_8037,N_8364);
nor U8465 (N_8465,N_8060,N_8020);
nand U8466 (N_8466,N_8379,N_8325);
nor U8467 (N_8467,N_8123,N_8047);
nor U8468 (N_8468,N_8340,N_8197);
or U8469 (N_8469,N_8239,N_8188);
nand U8470 (N_8470,N_8071,N_8169);
nor U8471 (N_8471,N_8130,N_8210);
nor U8472 (N_8472,N_8153,N_8093);
nand U8473 (N_8473,N_8011,N_8276);
xnor U8474 (N_8474,N_8337,N_8136);
and U8475 (N_8475,N_8199,N_8090);
or U8476 (N_8476,N_8009,N_8355);
xor U8477 (N_8477,N_8222,N_8183);
nand U8478 (N_8478,N_8038,N_8347);
and U8479 (N_8479,N_8307,N_8366);
or U8480 (N_8480,N_8203,N_8072);
nor U8481 (N_8481,N_8399,N_8267);
nor U8482 (N_8482,N_8358,N_8336);
nor U8483 (N_8483,N_8178,N_8023);
and U8484 (N_8484,N_8115,N_8076);
nand U8485 (N_8485,N_8029,N_8063);
and U8486 (N_8486,N_8240,N_8391);
and U8487 (N_8487,N_8376,N_8054);
nor U8488 (N_8488,N_8096,N_8272);
and U8489 (N_8489,N_8298,N_8057);
or U8490 (N_8490,N_8170,N_8311);
and U8491 (N_8491,N_8316,N_8185);
xnor U8492 (N_8492,N_8377,N_8002);
nor U8493 (N_8493,N_8342,N_8122);
nor U8494 (N_8494,N_8155,N_8362);
and U8495 (N_8495,N_8050,N_8066);
and U8496 (N_8496,N_8306,N_8196);
xor U8497 (N_8497,N_8258,N_8126);
and U8498 (N_8498,N_8251,N_8368);
or U8499 (N_8499,N_8320,N_8033);
or U8500 (N_8500,N_8083,N_8393);
xor U8501 (N_8501,N_8195,N_8024);
and U8502 (N_8502,N_8395,N_8315);
nand U8503 (N_8503,N_8112,N_8095);
nand U8504 (N_8504,N_8310,N_8087);
nand U8505 (N_8505,N_8107,N_8172);
and U8506 (N_8506,N_8254,N_8318);
and U8507 (N_8507,N_8326,N_8134);
and U8508 (N_8508,N_8133,N_8086);
or U8509 (N_8509,N_8193,N_8216);
nor U8510 (N_8510,N_8360,N_8232);
and U8511 (N_8511,N_8273,N_8397);
nor U8512 (N_8512,N_8290,N_8367);
xor U8513 (N_8513,N_8289,N_8041);
xor U8514 (N_8514,N_8046,N_8383);
or U8515 (N_8515,N_8341,N_8161);
xnor U8516 (N_8516,N_8295,N_8359);
and U8517 (N_8517,N_8200,N_8176);
xnor U8518 (N_8518,N_8128,N_8293);
nand U8519 (N_8519,N_8233,N_8187);
xor U8520 (N_8520,N_8371,N_8048);
xnor U8521 (N_8521,N_8114,N_8030);
or U8522 (N_8522,N_8327,N_8328);
nor U8523 (N_8523,N_8064,N_8053);
or U8524 (N_8524,N_8345,N_8154);
or U8525 (N_8525,N_8100,N_8005);
xnor U8526 (N_8526,N_8212,N_8278);
and U8527 (N_8527,N_8121,N_8163);
and U8528 (N_8528,N_8363,N_8058);
or U8529 (N_8529,N_8332,N_8228);
and U8530 (N_8530,N_8044,N_8061);
xor U8531 (N_8531,N_8268,N_8286);
nor U8532 (N_8532,N_8319,N_8277);
nor U8533 (N_8533,N_8157,N_8078);
or U8534 (N_8534,N_8113,N_8317);
nor U8535 (N_8535,N_8189,N_8032);
xor U8536 (N_8536,N_8287,N_8282);
nor U8537 (N_8537,N_8035,N_8089);
nor U8538 (N_8538,N_8116,N_8333);
xor U8539 (N_8539,N_8284,N_8149);
or U8540 (N_8540,N_8145,N_8271);
xnor U8541 (N_8541,N_8269,N_8106);
or U8542 (N_8542,N_8344,N_8213);
nand U8543 (N_8543,N_8229,N_8015);
nand U8544 (N_8544,N_8004,N_8354);
and U8545 (N_8545,N_8067,N_8174);
nand U8546 (N_8546,N_8322,N_8085);
or U8547 (N_8547,N_8003,N_8297);
xor U8548 (N_8548,N_8092,N_8158);
or U8549 (N_8549,N_8221,N_8088);
nand U8550 (N_8550,N_8069,N_8039);
or U8551 (N_8551,N_8102,N_8238);
or U8552 (N_8552,N_8175,N_8194);
and U8553 (N_8553,N_8215,N_8266);
nor U8554 (N_8554,N_8323,N_8129);
nor U8555 (N_8555,N_8001,N_8070);
or U8556 (N_8556,N_8013,N_8082);
nor U8557 (N_8557,N_8209,N_8208);
or U8558 (N_8558,N_8198,N_8217);
or U8559 (N_8559,N_8380,N_8324);
nor U8560 (N_8560,N_8225,N_8017);
and U8561 (N_8561,N_8262,N_8224);
or U8562 (N_8562,N_8249,N_8179);
xnor U8563 (N_8563,N_8010,N_8243);
and U8564 (N_8564,N_8299,N_8206);
xnor U8565 (N_8565,N_8205,N_8331);
and U8566 (N_8566,N_8117,N_8156);
and U8567 (N_8567,N_8007,N_8036);
nor U8568 (N_8568,N_8279,N_8231);
and U8569 (N_8569,N_8386,N_8109);
or U8570 (N_8570,N_8059,N_8356);
and U8571 (N_8571,N_8357,N_8202);
nor U8572 (N_8572,N_8241,N_8246);
or U8573 (N_8573,N_8280,N_8110);
nor U8574 (N_8574,N_8191,N_8019);
and U8575 (N_8575,N_8294,N_8218);
or U8576 (N_8576,N_8099,N_8162);
nor U8577 (N_8577,N_8283,N_8031);
nand U8578 (N_8578,N_8242,N_8353);
xor U8579 (N_8579,N_8260,N_8351);
or U8580 (N_8580,N_8021,N_8250);
or U8581 (N_8581,N_8350,N_8263);
nand U8582 (N_8582,N_8288,N_8180);
nand U8583 (N_8583,N_8008,N_8103);
xnor U8584 (N_8584,N_8223,N_8236);
or U8585 (N_8585,N_8334,N_8127);
or U8586 (N_8586,N_8381,N_8388);
or U8587 (N_8587,N_8253,N_8144);
and U8588 (N_8588,N_8075,N_8220);
nand U8589 (N_8589,N_8375,N_8292);
nor U8590 (N_8590,N_8352,N_8374);
and U8591 (N_8591,N_8137,N_8226);
or U8592 (N_8592,N_8387,N_8091);
xnor U8593 (N_8593,N_8077,N_8348);
and U8594 (N_8594,N_8270,N_8055);
nand U8595 (N_8595,N_8167,N_8201);
and U8596 (N_8596,N_8346,N_8098);
nand U8597 (N_8597,N_8012,N_8389);
xor U8598 (N_8598,N_8252,N_8022);
xnor U8599 (N_8599,N_8361,N_8296);
nand U8600 (N_8600,N_8136,N_8035);
or U8601 (N_8601,N_8274,N_8323);
and U8602 (N_8602,N_8194,N_8268);
nand U8603 (N_8603,N_8364,N_8324);
or U8604 (N_8604,N_8033,N_8012);
and U8605 (N_8605,N_8219,N_8194);
nor U8606 (N_8606,N_8141,N_8132);
xnor U8607 (N_8607,N_8034,N_8165);
xnor U8608 (N_8608,N_8138,N_8197);
xor U8609 (N_8609,N_8275,N_8079);
and U8610 (N_8610,N_8273,N_8086);
xnor U8611 (N_8611,N_8283,N_8371);
nand U8612 (N_8612,N_8120,N_8084);
or U8613 (N_8613,N_8318,N_8373);
xor U8614 (N_8614,N_8027,N_8121);
nand U8615 (N_8615,N_8227,N_8005);
xnor U8616 (N_8616,N_8069,N_8175);
or U8617 (N_8617,N_8393,N_8170);
or U8618 (N_8618,N_8362,N_8201);
nor U8619 (N_8619,N_8363,N_8190);
nand U8620 (N_8620,N_8364,N_8171);
nor U8621 (N_8621,N_8035,N_8104);
and U8622 (N_8622,N_8085,N_8032);
xor U8623 (N_8623,N_8193,N_8084);
xor U8624 (N_8624,N_8361,N_8248);
nor U8625 (N_8625,N_8213,N_8060);
and U8626 (N_8626,N_8397,N_8378);
and U8627 (N_8627,N_8236,N_8350);
nand U8628 (N_8628,N_8332,N_8065);
nand U8629 (N_8629,N_8160,N_8295);
or U8630 (N_8630,N_8220,N_8085);
nand U8631 (N_8631,N_8273,N_8317);
or U8632 (N_8632,N_8227,N_8172);
nor U8633 (N_8633,N_8163,N_8394);
and U8634 (N_8634,N_8370,N_8200);
nand U8635 (N_8635,N_8022,N_8021);
nor U8636 (N_8636,N_8194,N_8363);
or U8637 (N_8637,N_8268,N_8067);
and U8638 (N_8638,N_8357,N_8164);
and U8639 (N_8639,N_8247,N_8186);
or U8640 (N_8640,N_8026,N_8100);
nand U8641 (N_8641,N_8378,N_8222);
or U8642 (N_8642,N_8395,N_8084);
or U8643 (N_8643,N_8151,N_8057);
xor U8644 (N_8644,N_8305,N_8344);
and U8645 (N_8645,N_8324,N_8089);
and U8646 (N_8646,N_8102,N_8160);
and U8647 (N_8647,N_8265,N_8363);
and U8648 (N_8648,N_8175,N_8046);
xor U8649 (N_8649,N_8248,N_8357);
or U8650 (N_8650,N_8190,N_8054);
and U8651 (N_8651,N_8339,N_8291);
and U8652 (N_8652,N_8274,N_8231);
xor U8653 (N_8653,N_8264,N_8037);
nor U8654 (N_8654,N_8260,N_8021);
or U8655 (N_8655,N_8369,N_8002);
nor U8656 (N_8656,N_8103,N_8011);
nand U8657 (N_8657,N_8030,N_8371);
or U8658 (N_8658,N_8334,N_8244);
and U8659 (N_8659,N_8081,N_8132);
nor U8660 (N_8660,N_8388,N_8302);
nand U8661 (N_8661,N_8336,N_8343);
or U8662 (N_8662,N_8298,N_8248);
and U8663 (N_8663,N_8070,N_8262);
xnor U8664 (N_8664,N_8280,N_8179);
nand U8665 (N_8665,N_8213,N_8249);
xor U8666 (N_8666,N_8227,N_8174);
nand U8667 (N_8667,N_8349,N_8325);
or U8668 (N_8668,N_8309,N_8258);
or U8669 (N_8669,N_8151,N_8395);
and U8670 (N_8670,N_8353,N_8195);
nand U8671 (N_8671,N_8057,N_8167);
or U8672 (N_8672,N_8359,N_8173);
and U8673 (N_8673,N_8362,N_8394);
and U8674 (N_8674,N_8389,N_8016);
or U8675 (N_8675,N_8143,N_8342);
or U8676 (N_8676,N_8085,N_8014);
nand U8677 (N_8677,N_8268,N_8380);
and U8678 (N_8678,N_8366,N_8037);
nand U8679 (N_8679,N_8060,N_8395);
xnor U8680 (N_8680,N_8244,N_8300);
nand U8681 (N_8681,N_8247,N_8203);
xor U8682 (N_8682,N_8273,N_8165);
nand U8683 (N_8683,N_8370,N_8038);
xnor U8684 (N_8684,N_8064,N_8206);
xor U8685 (N_8685,N_8283,N_8228);
nand U8686 (N_8686,N_8235,N_8185);
xnor U8687 (N_8687,N_8157,N_8204);
nor U8688 (N_8688,N_8206,N_8213);
and U8689 (N_8689,N_8206,N_8391);
nor U8690 (N_8690,N_8338,N_8163);
or U8691 (N_8691,N_8194,N_8308);
or U8692 (N_8692,N_8388,N_8136);
nand U8693 (N_8693,N_8112,N_8341);
or U8694 (N_8694,N_8333,N_8169);
nand U8695 (N_8695,N_8057,N_8396);
or U8696 (N_8696,N_8287,N_8037);
nor U8697 (N_8697,N_8332,N_8092);
or U8698 (N_8698,N_8386,N_8117);
nand U8699 (N_8699,N_8076,N_8311);
or U8700 (N_8700,N_8131,N_8116);
nand U8701 (N_8701,N_8207,N_8323);
xnor U8702 (N_8702,N_8159,N_8375);
and U8703 (N_8703,N_8022,N_8036);
xnor U8704 (N_8704,N_8296,N_8008);
nor U8705 (N_8705,N_8180,N_8267);
and U8706 (N_8706,N_8237,N_8246);
and U8707 (N_8707,N_8147,N_8140);
xnor U8708 (N_8708,N_8212,N_8208);
nand U8709 (N_8709,N_8025,N_8069);
or U8710 (N_8710,N_8316,N_8229);
nand U8711 (N_8711,N_8216,N_8130);
or U8712 (N_8712,N_8118,N_8049);
xor U8713 (N_8713,N_8047,N_8009);
and U8714 (N_8714,N_8175,N_8203);
or U8715 (N_8715,N_8137,N_8122);
nand U8716 (N_8716,N_8076,N_8295);
or U8717 (N_8717,N_8302,N_8186);
or U8718 (N_8718,N_8200,N_8283);
nand U8719 (N_8719,N_8069,N_8349);
nor U8720 (N_8720,N_8376,N_8397);
or U8721 (N_8721,N_8179,N_8393);
nand U8722 (N_8722,N_8048,N_8130);
xor U8723 (N_8723,N_8101,N_8004);
or U8724 (N_8724,N_8268,N_8220);
or U8725 (N_8725,N_8066,N_8386);
nand U8726 (N_8726,N_8123,N_8206);
or U8727 (N_8727,N_8147,N_8156);
xor U8728 (N_8728,N_8213,N_8176);
xnor U8729 (N_8729,N_8242,N_8075);
or U8730 (N_8730,N_8120,N_8217);
or U8731 (N_8731,N_8068,N_8207);
nand U8732 (N_8732,N_8292,N_8061);
nand U8733 (N_8733,N_8008,N_8119);
nor U8734 (N_8734,N_8043,N_8297);
and U8735 (N_8735,N_8234,N_8302);
xnor U8736 (N_8736,N_8030,N_8352);
nor U8737 (N_8737,N_8121,N_8096);
nor U8738 (N_8738,N_8215,N_8193);
nor U8739 (N_8739,N_8327,N_8174);
nor U8740 (N_8740,N_8224,N_8038);
xor U8741 (N_8741,N_8138,N_8293);
or U8742 (N_8742,N_8037,N_8115);
xnor U8743 (N_8743,N_8192,N_8210);
nor U8744 (N_8744,N_8201,N_8072);
and U8745 (N_8745,N_8266,N_8063);
and U8746 (N_8746,N_8205,N_8337);
and U8747 (N_8747,N_8011,N_8274);
nor U8748 (N_8748,N_8060,N_8078);
xor U8749 (N_8749,N_8108,N_8217);
xor U8750 (N_8750,N_8053,N_8147);
and U8751 (N_8751,N_8149,N_8371);
nor U8752 (N_8752,N_8074,N_8213);
and U8753 (N_8753,N_8034,N_8250);
nand U8754 (N_8754,N_8299,N_8040);
or U8755 (N_8755,N_8109,N_8006);
and U8756 (N_8756,N_8185,N_8342);
nor U8757 (N_8757,N_8080,N_8360);
nor U8758 (N_8758,N_8303,N_8056);
or U8759 (N_8759,N_8362,N_8286);
or U8760 (N_8760,N_8090,N_8111);
nor U8761 (N_8761,N_8052,N_8098);
and U8762 (N_8762,N_8057,N_8270);
xor U8763 (N_8763,N_8379,N_8171);
or U8764 (N_8764,N_8127,N_8351);
and U8765 (N_8765,N_8169,N_8037);
xor U8766 (N_8766,N_8010,N_8157);
or U8767 (N_8767,N_8225,N_8333);
xnor U8768 (N_8768,N_8021,N_8382);
or U8769 (N_8769,N_8035,N_8100);
or U8770 (N_8770,N_8274,N_8073);
and U8771 (N_8771,N_8291,N_8334);
or U8772 (N_8772,N_8077,N_8357);
nand U8773 (N_8773,N_8170,N_8347);
and U8774 (N_8774,N_8268,N_8365);
or U8775 (N_8775,N_8271,N_8045);
nand U8776 (N_8776,N_8043,N_8362);
or U8777 (N_8777,N_8281,N_8078);
nor U8778 (N_8778,N_8232,N_8135);
or U8779 (N_8779,N_8258,N_8223);
and U8780 (N_8780,N_8202,N_8199);
nor U8781 (N_8781,N_8075,N_8141);
xor U8782 (N_8782,N_8358,N_8133);
nand U8783 (N_8783,N_8300,N_8325);
and U8784 (N_8784,N_8186,N_8292);
nor U8785 (N_8785,N_8351,N_8306);
nor U8786 (N_8786,N_8180,N_8214);
or U8787 (N_8787,N_8308,N_8166);
and U8788 (N_8788,N_8064,N_8393);
xnor U8789 (N_8789,N_8255,N_8306);
and U8790 (N_8790,N_8167,N_8027);
nand U8791 (N_8791,N_8251,N_8059);
xor U8792 (N_8792,N_8132,N_8274);
nand U8793 (N_8793,N_8003,N_8287);
nor U8794 (N_8794,N_8233,N_8373);
nand U8795 (N_8795,N_8209,N_8149);
or U8796 (N_8796,N_8077,N_8303);
and U8797 (N_8797,N_8344,N_8086);
or U8798 (N_8798,N_8082,N_8090);
xor U8799 (N_8799,N_8197,N_8206);
xor U8800 (N_8800,N_8434,N_8768);
or U8801 (N_8801,N_8706,N_8789);
nand U8802 (N_8802,N_8426,N_8703);
xor U8803 (N_8803,N_8428,N_8702);
xnor U8804 (N_8804,N_8613,N_8620);
and U8805 (N_8805,N_8565,N_8499);
nand U8806 (N_8806,N_8555,N_8720);
nand U8807 (N_8807,N_8781,N_8569);
xnor U8808 (N_8808,N_8770,N_8719);
nand U8809 (N_8809,N_8525,N_8616);
nor U8810 (N_8810,N_8679,N_8415);
and U8811 (N_8811,N_8503,N_8694);
or U8812 (N_8812,N_8466,N_8611);
nor U8813 (N_8813,N_8480,N_8442);
nand U8814 (N_8814,N_8539,N_8598);
nor U8815 (N_8815,N_8500,N_8519);
or U8816 (N_8816,N_8410,N_8491);
and U8817 (N_8817,N_8521,N_8628);
and U8818 (N_8818,N_8537,N_8663);
nor U8819 (N_8819,N_8402,N_8531);
xor U8820 (N_8820,N_8680,N_8448);
and U8821 (N_8821,N_8504,N_8748);
and U8822 (N_8822,N_8751,N_8455);
xnor U8823 (N_8823,N_8786,N_8414);
nor U8824 (N_8824,N_8427,N_8479);
nand U8825 (N_8825,N_8723,N_8743);
nand U8826 (N_8826,N_8665,N_8474);
xnor U8827 (N_8827,N_8785,N_8669);
nor U8828 (N_8828,N_8655,N_8450);
or U8829 (N_8829,N_8619,N_8766);
xor U8830 (N_8830,N_8754,N_8429);
nand U8831 (N_8831,N_8648,N_8696);
nand U8832 (N_8832,N_8653,N_8716);
xor U8833 (N_8833,N_8490,N_8452);
or U8834 (N_8834,N_8632,N_8642);
or U8835 (N_8835,N_8566,N_8691);
nor U8836 (N_8836,N_8712,N_8626);
and U8837 (N_8837,N_8534,N_8631);
nor U8838 (N_8838,N_8532,N_8467);
or U8839 (N_8839,N_8515,N_8562);
nor U8840 (N_8840,N_8722,N_8633);
nor U8841 (N_8841,N_8658,N_8511);
or U8842 (N_8842,N_8713,N_8798);
xor U8843 (N_8843,N_8693,N_8670);
nor U8844 (N_8844,N_8721,N_8661);
xnor U8845 (N_8845,N_8675,N_8441);
nor U8846 (N_8846,N_8522,N_8596);
nand U8847 (N_8847,N_8592,N_8641);
nand U8848 (N_8848,N_8697,N_8733);
nand U8849 (N_8849,N_8469,N_8627);
nor U8850 (N_8850,N_8530,N_8728);
nor U8851 (N_8851,N_8507,N_8541);
nand U8852 (N_8852,N_8659,N_8540);
and U8853 (N_8853,N_8704,N_8650);
nor U8854 (N_8854,N_8673,N_8690);
nor U8855 (N_8855,N_8581,N_8502);
nor U8856 (N_8856,N_8705,N_8656);
xor U8857 (N_8857,N_8423,N_8464);
and U8858 (N_8858,N_8477,N_8593);
xor U8859 (N_8859,N_8440,N_8484);
xor U8860 (N_8860,N_8692,N_8585);
xor U8861 (N_8861,N_8462,N_8666);
or U8862 (N_8862,N_8437,N_8518);
nand U8863 (N_8863,N_8422,N_8580);
nand U8864 (N_8864,N_8573,N_8418);
nor U8865 (N_8865,N_8408,N_8471);
nor U8866 (N_8866,N_8470,N_8589);
nor U8867 (N_8867,N_8501,N_8439);
and U8868 (N_8868,N_8623,N_8579);
xor U8869 (N_8869,N_8472,N_8784);
and U8870 (N_8870,N_8514,N_8535);
nor U8871 (N_8871,N_8454,N_8735);
and U8872 (N_8872,N_8796,N_8447);
nand U8873 (N_8873,N_8451,N_8523);
and U8874 (N_8874,N_8793,N_8652);
xor U8875 (N_8875,N_8568,N_8788);
and U8876 (N_8876,N_8438,N_8605);
xnor U8877 (N_8877,N_8404,N_8513);
nor U8878 (N_8878,N_8699,N_8453);
nor U8879 (N_8879,N_8756,N_8506);
or U8880 (N_8880,N_8591,N_8553);
or U8881 (N_8881,N_8604,N_8638);
or U8882 (N_8882,N_8497,N_8752);
and U8883 (N_8883,N_8446,N_8560);
and U8884 (N_8884,N_8738,N_8400);
or U8885 (N_8885,N_8558,N_8516);
and U8886 (N_8886,N_8584,N_8639);
xnor U8887 (N_8887,N_8629,N_8567);
or U8888 (N_8888,N_8533,N_8463);
nand U8889 (N_8889,N_8674,N_8622);
or U8890 (N_8890,N_8487,N_8767);
and U8891 (N_8891,N_8636,N_8577);
and U8892 (N_8892,N_8664,N_8481);
xnor U8893 (N_8893,N_8783,N_8729);
nor U8894 (N_8894,N_8420,N_8688);
and U8895 (N_8895,N_8630,N_8700);
and U8896 (N_8896,N_8774,N_8787);
nand U8897 (N_8897,N_8780,N_8777);
nor U8898 (N_8898,N_8776,N_8610);
nand U8899 (N_8899,N_8625,N_8778);
or U8900 (N_8900,N_8764,N_8475);
nor U8901 (N_8901,N_8473,N_8744);
nand U8902 (N_8902,N_8779,N_8763);
nor U8903 (N_8903,N_8709,N_8492);
xor U8904 (N_8904,N_8635,N_8430);
and U8905 (N_8905,N_8714,N_8747);
nor U8906 (N_8906,N_8557,N_8510);
nor U8907 (N_8907,N_8755,N_8436);
xnor U8908 (N_8908,N_8493,N_8496);
or U8909 (N_8909,N_8667,N_8771);
nor U8910 (N_8910,N_8782,N_8409);
nor U8911 (N_8911,N_8517,N_8606);
or U8912 (N_8912,N_8551,N_8730);
xor U8913 (N_8913,N_8791,N_8603);
nor U8914 (N_8914,N_8746,N_8654);
nand U8915 (N_8915,N_8765,N_8526);
nor U8916 (N_8916,N_8644,N_8740);
xor U8917 (N_8917,N_8405,N_8571);
nor U8918 (N_8918,N_8701,N_8576);
and U8919 (N_8919,N_8615,N_8758);
xnor U8920 (N_8920,N_8621,N_8677);
and U8921 (N_8921,N_8760,N_8542);
nand U8922 (N_8922,N_8682,N_8741);
and U8923 (N_8923,N_8456,N_8538);
or U8924 (N_8924,N_8505,N_8695);
or U8925 (N_8925,N_8545,N_8524);
or U8926 (N_8926,N_8757,N_8710);
xnor U8927 (N_8927,N_8753,N_8412);
nand U8928 (N_8928,N_8528,N_8407);
nor U8929 (N_8929,N_8489,N_8548);
and U8930 (N_8930,N_8676,N_8601);
xor U8931 (N_8931,N_8707,N_8544);
and U8932 (N_8932,N_8731,N_8687);
and U8933 (N_8933,N_8646,N_8640);
nand U8934 (N_8934,N_8583,N_8561);
xnor U8935 (N_8935,N_8761,N_8465);
nor U8936 (N_8936,N_8660,N_8403);
xor U8937 (N_8937,N_8671,N_8424);
and U8938 (N_8938,N_8468,N_8483);
nor U8939 (N_8939,N_8609,N_8549);
or U8940 (N_8940,N_8689,N_8684);
or U8941 (N_8941,N_8634,N_8509);
and U8942 (N_8942,N_8749,N_8457);
xnor U8943 (N_8943,N_8662,N_8794);
or U8944 (N_8944,N_8647,N_8546);
nand U8945 (N_8945,N_8726,N_8445);
xnor U8946 (N_8946,N_8586,N_8708);
or U8947 (N_8947,N_8797,N_8724);
nor U8948 (N_8948,N_8482,N_8431);
or U8949 (N_8949,N_8582,N_8529);
and U8950 (N_8950,N_8432,N_8624);
nor U8951 (N_8951,N_8547,N_8792);
and U8952 (N_8952,N_8718,N_8637);
and U8953 (N_8953,N_8643,N_8750);
nand U8954 (N_8954,N_8421,N_8618);
nor U8955 (N_8955,N_8590,N_8795);
nand U8956 (N_8956,N_8433,N_8488);
xnor U8957 (N_8957,N_8790,N_8681);
and U8958 (N_8958,N_8678,N_8425);
or U8959 (N_8959,N_8494,N_8737);
nand U8960 (N_8960,N_8612,N_8485);
and U8961 (N_8961,N_8554,N_8772);
nand U8962 (N_8962,N_8683,N_8587);
nand U8963 (N_8963,N_8769,N_8727);
nor U8964 (N_8964,N_8419,N_8498);
xor U8965 (N_8965,N_8645,N_8672);
and U8966 (N_8966,N_8668,N_8734);
or U8967 (N_8967,N_8685,N_8799);
or U8968 (N_8968,N_8739,N_8443);
nand U8969 (N_8969,N_8401,N_8649);
nand U8970 (N_8970,N_8572,N_8406);
and U8971 (N_8971,N_8411,N_8742);
nand U8972 (N_8972,N_8608,N_8745);
and U8973 (N_8973,N_8575,N_8449);
and U8974 (N_8974,N_8651,N_8460);
or U8975 (N_8975,N_8578,N_8588);
nor U8976 (N_8976,N_8476,N_8552);
and U8977 (N_8977,N_8413,N_8599);
nand U8978 (N_8978,N_8594,N_8527);
nand U8979 (N_8979,N_8600,N_8574);
xor U8980 (N_8980,N_8607,N_8614);
nand U8981 (N_8981,N_8512,N_8486);
nand U8982 (N_8982,N_8459,N_8461);
nor U8983 (N_8983,N_8736,N_8556);
and U8984 (N_8984,N_8550,N_8762);
nand U8985 (N_8985,N_8595,N_8711);
nor U8986 (N_8986,N_8717,N_8602);
nand U8987 (N_8987,N_8458,N_8563);
nand U8988 (N_8988,N_8759,N_8775);
and U8989 (N_8989,N_8508,N_8520);
xnor U8990 (N_8990,N_8564,N_8417);
xnor U8991 (N_8991,N_8686,N_8725);
and U8992 (N_8992,N_8657,N_8732);
nor U8993 (N_8993,N_8444,N_8559);
nor U8994 (N_8994,N_8495,N_8543);
and U8995 (N_8995,N_8617,N_8478);
xnor U8996 (N_8996,N_8536,N_8435);
or U8997 (N_8997,N_8773,N_8698);
nand U8998 (N_8998,N_8416,N_8597);
or U8999 (N_8999,N_8570,N_8715);
nand U9000 (N_9000,N_8575,N_8770);
xnor U9001 (N_9001,N_8717,N_8613);
nor U9002 (N_9002,N_8604,N_8594);
nor U9003 (N_9003,N_8727,N_8634);
nand U9004 (N_9004,N_8477,N_8664);
nand U9005 (N_9005,N_8568,N_8699);
nor U9006 (N_9006,N_8571,N_8707);
nor U9007 (N_9007,N_8597,N_8541);
or U9008 (N_9008,N_8619,N_8698);
nor U9009 (N_9009,N_8796,N_8667);
or U9010 (N_9010,N_8687,N_8441);
nand U9011 (N_9011,N_8444,N_8539);
and U9012 (N_9012,N_8782,N_8710);
nand U9013 (N_9013,N_8798,N_8501);
xnor U9014 (N_9014,N_8604,N_8602);
nand U9015 (N_9015,N_8792,N_8614);
xnor U9016 (N_9016,N_8542,N_8515);
nand U9017 (N_9017,N_8780,N_8755);
or U9018 (N_9018,N_8494,N_8550);
nor U9019 (N_9019,N_8760,N_8677);
xnor U9020 (N_9020,N_8789,N_8712);
nand U9021 (N_9021,N_8573,N_8603);
nor U9022 (N_9022,N_8503,N_8524);
and U9023 (N_9023,N_8619,N_8724);
nor U9024 (N_9024,N_8775,N_8509);
xor U9025 (N_9025,N_8511,N_8590);
and U9026 (N_9026,N_8601,N_8431);
and U9027 (N_9027,N_8468,N_8758);
nor U9028 (N_9028,N_8749,N_8555);
xnor U9029 (N_9029,N_8572,N_8410);
or U9030 (N_9030,N_8579,N_8667);
xor U9031 (N_9031,N_8536,N_8578);
nand U9032 (N_9032,N_8730,N_8449);
nor U9033 (N_9033,N_8471,N_8632);
xor U9034 (N_9034,N_8461,N_8565);
nor U9035 (N_9035,N_8460,N_8465);
and U9036 (N_9036,N_8607,N_8508);
or U9037 (N_9037,N_8738,N_8770);
xor U9038 (N_9038,N_8438,N_8563);
and U9039 (N_9039,N_8737,N_8667);
nor U9040 (N_9040,N_8621,N_8775);
and U9041 (N_9041,N_8508,N_8423);
xnor U9042 (N_9042,N_8476,N_8649);
xnor U9043 (N_9043,N_8527,N_8436);
and U9044 (N_9044,N_8522,N_8640);
nand U9045 (N_9045,N_8417,N_8435);
xor U9046 (N_9046,N_8638,N_8535);
xor U9047 (N_9047,N_8429,N_8549);
xor U9048 (N_9048,N_8588,N_8437);
and U9049 (N_9049,N_8591,N_8452);
nand U9050 (N_9050,N_8716,N_8593);
or U9051 (N_9051,N_8700,N_8792);
or U9052 (N_9052,N_8770,N_8493);
and U9053 (N_9053,N_8473,N_8435);
nor U9054 (N_9054,N_8649,N_8559);
xnor U9055 (N_9055,N_8534,N_8569);
nor U9056 (N_9056,N_8610,N_8639);
and U9057 (N_9057,N_8580,N_8760);
nand U9058 (N_9058,N_8523,N_8580);
and U9059 (N_9059,N_8628,N_8513);
xnor U9060 (N_9060,N_8651,N_8680);
xnor U9061 (N_9061,N_8489,N_8794);
nor U9062 (N_9062,N_8604,N_8415);
xnor U9063 (N_9063,N_8738,N_8737);
nand U9064 (N_9064,N_8578,N_8478);
and U9065 (N_9065,N_8518,N_8477);
or U9066 (N_9066,N_8689,N_8651);
xnor U9067 (N_9067,N_8480,N_8724);
xnor U9068 (N_9068,N_8558,N_8489);
xor U9069 (N_9069,N_8447,N_8423);
or U9070 (N_9070,N_8698,N_8718);
xnor U9071 (N_9071,N_8694,N_8495);
or U9072 (N_9072,N_8760,N_8506);
and U9073 (N_9073,N_8734,N_8755);
and U9074 (N_9074,N_8738,N_8583);
or U9075 (N_9075,N_8424,N_8486);
nor U9076 (N_9076,N_8615,N_8663);
nor U9077 (N_9077,N_8616,N_8679);
nor U9078 (N_9078,N_8662,N_8486);
xnor U9079 (N_9079,N_8515,N_8435);
nand U9080 (N_9080,N_8440,N_8428);
xnor U9081 (N_9081,N_8568,N_8795);
xnor U9082 (N_9082,N_8772,N_8657);
or U9083 (N_9083,N_8441,N_8785);
and U9084 (N_9084,N_8754,N_8770);
xor U9085 (N_9085,N_8600,N_8503);
nor U9086 (N_9086,N_8479,N_8428);
and U9087 (N_9087,N_8667,N_8466);
xnor U9088 (N_9088,N_8448,N_8548);
and U9089 (N_9089,N_8604,N_8477);
and U9090 (N_9090,N_8736,N_8758);
and U9091 (N_9091,N_8687,N_8655);
and U9092 (N_9092,N_8446,N_8566);
or U9093 (N_9093,N_8457,N_8465);
and U9094 (N_9094,N_8567,N_8528);
nand U9095 (N_9095,N_8729,N_8781);
xor U9096 (N_9096,N_8526,N_8785);
nand U9097 (N_9097,N_8431,N_8797);
or U9098 (N_9098,N_8583,N_8646);
nor U9099 (N_9099,N_8493,N_8617);
and U9100 (N_9100,N_8418,N_8667);
or U9101 (N_9101,N_8513,N_8414);
or U9102 (N_9102,N_8678,N_8448);
nand U9103 (N_9103,N_8760,N_8613);
nor U9104 (N_9104,N_8740,N_8577);
xor U9105 (N_9105,N_8758,N_8648);
nand U9106 (N_9106,N_8428,N_8658);
or U9107 (N_9107,N_8528,N_8592);
xnor U9108 (N_9108,N_8477,N_8578);
xor U9109 (N_9109,N_8569,N_8626);
nor U9110 (N_9110,N_8501,N_8787);
nor U9111 (N_9111,N_8770,N_8700);
or U9112 (N_9112,N_8573,N_8529);
nor U9113 (N_9113,N_8575,N_8772);
xnor U9114 (N_9114,N_8566,N_8438);
or U9115 (N_9115,N_8586,N_8584);
nand U9116 (N_9116,N_8522,N_8585);
or U9117 (N_9117,N_8723,N_8542);
or U9118 (N_9118,N_8402,N_8583);
xnor U9119 (N_9119,N_8438,N_8425);
nor U9120 (N_9120,N_8564,N_8679);
and U9121 (N_9121,N_8409,N_8604);
nor U9122 (N_9122,N_8468,N_8723);
or U9123 (N_9123,N_8442,N_8740);
xnor U9124 (N_9124,N_8799,N_8571);
or U9125 (N_9125,N_8711,N_8522);
and U9126 (N_9126,N_8517,N_8585);
and U9127 (N_9127,N_8759,N_8607);
xnor U9128 (N_9128,N_8713,N_8431);
and U9129 (N_9129,N_8787,N_8415);
xnor U9130 (N_9130,N_8752,N_8759);
nor U9131 (N_9131,N_8599,N_8640);
or U9132 (N_9132,N_8657,N_8609);
or U9133 (N_9133,N_8706,N_8623);
nand U9134 (N_9134,N_8690,N_8539);
and U9135 (N_9135,N_8502,N_8735);
xor U9136 (N_9136,N_8758,N_8560);
xor U9137 (N_9137,N_8793,N_8503);
and U9138 (N_9138,N_8756,N_8449);
xor U9139 (N_9139,N_8563,N_8568);
or U9140 (N_9140,N_8480,N_8513);
nand U9141 (N_9141,N_8715,N_8476);
and U9142 (N_9142,N_8775,N_8564);
nand U9143 (N_9143,N_8400,N_8688);
nor U9144 (N_9144,N_8748,N_8663);
and U9145 (N_9145,N_8665,N_8714);
nand U9146 (N_9146,N_8504,N_8419);
xor U9147 (N_9147,N_8659,N_8402);
and U9148 (N_9148,N_8543,N_8457);
or U9149 (N_9149,N_8771,N_8475);
xor U9150 (N_9150,N_8615,N_8488);
or U9151 (N_9151,N_8466,N_8632);
or U9152 (N_9152,N_8512,N_8694);
or U9153 (N_9153,N_8704,N_8766);
xnor U9154 (N_9154,N_8717,N_8783);
or U9155 (N_9155,N_8530,N_8737);
nor U9156 (N_9156,N_8753,N_8664);
xnor U9157 (N_9157,N_8691,N_8439);
and U9158 (N_9158,N_8777,N_8789);
nor U9159 (N_9159,N_8570,N_8559);
or U9160 (N_9160,N_8698,N_8767);
nand U9161 (N_9161,N_8799,N_8595);
nor U9162 (N_9162,N_8458,N_8660);
xnor U9163 (N_9163,N_8444,N_8553);
nand U9164 (N_9164,N_8674,N_8573);
and U9165 (N_9165,N_8510,N_8459);
and U9166 (N_9166,N_8463,N_8591);
nor U9167 (N_9167,N_8418,N_8798);
nand U9168 (N_9168,N_8634,N_8627);
xor U9169 (N_9169,N_8626,N_8567);
nor U9170 (N_9170,N_8720,N_8786);
or U9171 (N_9171,N_8743,N_8736);
nand U9172 (N_9172,N_8440,N_8695);
xor U9173 (N_9173,N_8623,N_8632);
and U9174 (N_9174,N_8771,N_8517);
or U9175 (N_9175,N_8438,N_8582);
nand U9176 (N_9176,N_8679,N_8498);
nor U9177 (N_9177,N_8467,N_8411);
xor U9178 (N_9178,N_8715,N_8798);
nand U9179 (N_9179,N_8637,N_8500);
nand U9180 (N_9180,N_8530,N_8750);
nor U9181 (N_9181,N_8755,N_8417);
or U9182 (N_9182,N_8576,N_8689);
xnor U9183 (N_9183,N_8761,N_8653);
nand U9184 (N_9184,N_8418,N_8409);
nor U9185 (N_9185,N_8692,N_8431);
nor U9186 (N_9186,N_8766,N_8705);
nand U9187 (N_9187,N_8483,N_8743);
xor U9188 (N_9188,N_8679,N_8789);
nor U9189 (N_9189,N_8431,N_8411);
nor U9190 (N_9190,N_8516,N_8707);
or U9191 (N_9191,N_8685,N_8405);
or U9192 (N_9192,N_8567,N_8590);
nor U9193 (N_9193,N_8707,N_8648);
and U9194 (N_9194,N_8645,N_8553);
xnor U9195 (N_9195,N_8682,N_8412);
nand U9196 (N_9196,N_8704,N_8551);
or U9197 (N_9197,N_8628,N_8626);
xnor U9198 (N_9198,N_8461,N_8732);
nor U9199 (N_9199,N_8490,N_8736);
and U9200 (N_9200,N_9109,N_8930);
and U9201 (N_9201,N_9175,N_9011);
xnor U9202 (N_9202,N_8813,N_9036);
and U9203 (N_9203,N_8875,N_9085);
nand U9204 (N_9204,N_9081,N_8853);
nand U9205 (N_9205,N_8925,N_8883);
xor U9206 (N_9206,N_8822,N_9114);
nor U9207 (N_9207,N_8997,N_9063);
nor U9208 (N_9208,N_9026,N_8965);
and U9209 (N_9209,N_8990,N_9054);
nor U9210 (N_9210,N_8985,N_9041);
and U9211 (N_9211,N_8869,N_9040);
or U9212 (N_9212,N_8898,N_8895);
xnor U9213 (N_9213,N_8958,N_8839);
nor U9214 (N_9214,N_9037,N_9009);
and U9215 (N_9215,N_8992,N_8834);
nor U9216 (N_9216,N_8846,N_8908);
xnor U9217 (N_9217,N_8996,N_8849);
and U9218 (N_9218,N_9127,N_9192);
and U9219 (N_9219,N_9100,N_8946);
nor U9220 (N_9220,N_9057,N_9065);
xnor U9221 (N_9221,N_8979,N_9033);
and U9222 (N_9222,N_9130,N_8810);
xor U9223 (N_9223,N_8874,N_9016);
and U9224 (N_9224,N_9053,N_9168);
or U9225 (N_9225,N_9073,N_8973);
nor U9226 (N_9226,N_8879,N_8949);
nor U9227 (N_9227,N_8963,N_9074);
nor U9228 (N_9228,N_9088,N_9008);
or U9229 (N_9229,N_9056,N_9162);
xor U9230 (N_9230,N_9119,N_8987);
nor U9231 (N_9231,N_8868,N_9050);
nand U9232 (N_9232,N_8820,N_9195);
or U9233 (N_9233,N_8824,N_9161);
nand U9234 (N_9234,N_8843,N_8901);
xor U9235 (N_9235,N_8931,N_9124);
nor U9236 (N_9236,N_9052,N_9149);
nor U9237 (N_9237,N_9187,N_9158);
xnor U9238 (N_9238,N_9047,N_8809);
nand U9239 (N_9239,N_8984,N_9121);
and U9240 (N_9240,N_8845,N_8871);
or U9241 (N_9241,N_9173,N_8886);
or U9242 (N_9242,N_9039,N_8876);
nor U9243 (N_9243,N_8815,N_8932);
xnor U9244 (N_9244,N_8988,N_8808);
and U9245 (N_9245,N_8904,N_9046);
nor U9246 (N_9246,N_8960,N_8903);
nand U9247 (N_9247,N_9086,N_8844);
and U9248 (N_9248,N_9079,N_9171);
and U9249 (N_9249,N_8881,N_8975);
and U9250 (N_9250,N_9004,N_9083);
or U9251 (N_9251,N_8961,N_9190);
and U9252 (N_9252,N_8819,N_8905);
or U9253 (N_9253,N_9105,N_9193);
and U9254 (N_9254,N_8827,N_9154);
xnor U9255 (N_9255,N_8801,N_9091);
nor U9256 (N_9256,N_8998,N_8938);
nand U9257 (N_9257,N_9166,N_8995);
xor U9258 (N_9258,N_9131,N_8914);
xor U9259 (N_9259,N_8966,N_9059);
nor U9260 (N_9260,N_8939,N_8842);
nor U9261 (N_9261,N_9156,N_9113);
xor U9262 (N_9262,N_8902,N_8877);
and U9263 (N_9263,N_8872,N_8974);
and U9264 (N_9264,N_8866,N_8863);
or U9265 (N_9265,N_8918,N_9188);
nor U9266 (N_9266,N_8880,N_8935);
or U9267 (N_9267,N_9032,N_9071);
or U9268 (N_9268,N_8882,N_9191);
nor U9269 (N_9269,N_9020,N_8894);
xor U9270 (N_9270,N_8805,N_9189);
or U9271 (N_9271,N_9178,N_9031);
xnor U9272 (N_9272,N_9185,N_9066);
or U9273 (N_9273,N_8867,N_8993);
nand U9274 (N_9274,N_8900,N_8972);
nor U9275 (N_9275,N_9140,N_9028);
and U9276 (N_9276,N_8826,N_9023);
xnor U9277 (N_9277,N_8971,N_8923);
nand U9278 (N_9278,N_8916,N_9038);
nor U9279 (N_9279,N_8897,N_8994);
nand U9280 (N_9280,N_9197,N_9148);
nand U9281 (N_9281,N_8864,N_9034);
nor U9282 (N_9282,N_9144,N_8964);
nand U9283 (N_9283,N_9029,N_8855);
nand U9284 (N_9284,N_9062,N_9024);
nor U9285 (N_9285,N_9129,N_9194);
and U9286 (N_9286,N_9172,N_8847);
or U9287 (N_9287,N_9112,N_9134);
and U9288 (N_9288,N_8989,N_8928);
xnor U9289 (N_9289,N_8982,N_8991);
xor U9290 (N_9290,N_8926,N_8951);
nor U9291 (N_9291,N_9097,N_8873);
xnor U9292 (N_9292,N_9183,N_8915);
nor U9293 (N_9293,N_9084,N_8832);
nand U9294 (N_9294,N_8841,N_8919);
and U9295 (N_9295,N_8850,N_8977);
nand U9296 (N_9296,N_8887,N_9153);
xor U9297 (N_9297,N_9170,N_8943);
and U9298 (N_9298,N_8806,N_9089);
or U9299 (N_9299,N_9164,N_9117);
nand U9300 (N_9300,N_9139,N_9001);
nor U9301 (N_9301,N_8944,N_9045);
nand U9302 (N_9302,N_9080,N_9179);
or U9303 (N_9303,N_9069,N_8899);
or U9304 (N_9304,N_8907,N_9196);
or U9305 (N_9305,N_8941,N_9058);
and U9306 (N_9306,N_8823,N_8959);
nor U9307 (N_9307,N_9005,N_8857);
and U9308 (N_9308,N_8924,N_9049);
xor U9309 (N_9309,N_9169,N_8955);
xnor U9310 (N_9310,N_9132,N_8962);
or U9311 (N_9311,N_9101,N_9143);
nand U9312 (N_9312,N_8929,N_9048);
and U9313 (N_9313,N_9107,N_8921);
xor U9314 (N_9314,N_8896,N_8833);
xnor U9315 (N_9315,N_8828,N_8862);
and U9316 (N_9316,N_9111,N_9075);
nor U9317 (N_9317,N_8968,N_8836);
or U9318 (N_9318,N_8840,N_8980);
and U9319 (N_9319,N_9147,N_8838);
or U9320 (N_9320,N_8969,N_8865);
nand U9321 (N_9321,N_8956,N_9019);
and U9322 (N_9322,N_9198,N_9155);
or U9323 (N_9323,N_8978,N_8825);
nand U9324 (N_9324,N_9022,N_9072);
and U9325 (N_9325,N_8811,N_9110);
and U9326 (N_9326,N_8976,N_9136);
nor U9327 (N_9327,N_8803,N_9106);
nor U9328 (N_9328,N_9115,N_9051);
or U9329 (N_9329,N_9021,N_8848);
nor U9330 (N_9330,N_8802,N_8859);
xnor U9331 (N_9331,N_8922,N_8888);
and U9332 (N_9332,N_9077,N_9012);
nor U9333 (N_9333,N_8927,N_9116);
or U9334 (N_9334,N_9151,N_9182);
xnor U9335 (N_9335,N_8878,N_8954);
nand U9336 (N_9336,N_8950,N_9096);
or U9337 (N_9337,N_8814,N_9174);
and U9338 (N_9338,N_9165,N_9099);
or U9339 (N_9339,N_8933,N_8957);
nand U9340 (N_9340,N_9068,N_9138);
nor U9341 (N_9341,N_8917,N_9142);
xor U9342 (N_9342,N_9092,N_9137);
xnor U9343 (N_9343,N_9003,N_9120);
and U9344 (N_9344,N_8893,N_9013);
nor U9345 (N_9345,N_9094,N_8970);
or U9346 (N_9346,N_9141,N_9122);
nand U9347 (N_9347,N_8817,N_9076);
or U9348 (N_9348,N_9126,N_8999);
or U9349 (N_9349,N_8856,N_8936);
and U9350 (N_9350,N_8948,N_9018);
nor U9351 (N_9351,N_8913,N_9199);
and U9352 (N_9352,N_8940,N_9135);
xnor U9353 (N_9353,N_9181,N_8800);
nor U9354 (N_9354,N_8909,N_9030);
nand U9355 (N_9355,N_8920,N_8945);
nor U9356 (N_9356,N_9103,N_9015);
and U9357 (N_9357,N_9104,N_9027);
and U9358 (N_9358,N_9098,N_8851);
xor U9359 (N_9359,N_9093,N_8934);
nand U9360 (N_9360,N_9082,N_8937);
and U9361 (N_9361,N_8830,N_9035);
nand U9362 (N_9362,N_8804,N_9159);
nand U9363 (N_9363,N_8870,N_9017);
xnor U9364 (N_9364,N_9014,N_9006);
nor U9365 (N_9365,N_9025,N_9108);
or U9366 (N_9366,N_9043,N_9184);
and U9367 (N_9367,N_9070,N_8906);
nand U9368 (N_9368,N_9180,N_9152);
and U9369 (N_9369,N_8860,N_8952);
and U9370 (N_9370,N_8816,N_8854);
nand U9371 (N_9371,N_8911,N_9010);
nand U9372 (N_9372,N_8885,N_9000);
or U9373 (N_9373,N_8837,N_8947);
or U9374 (N_9374,N_8981,N_8910);
xnor U9375 (N_9375,N_9095,N_9064);
and U9376 (N_9376,N_9067,N_9146);
nand U9377 (N_9377,N_9150,N_9157);
nor U9378 (N_9378,N_8852,N_9125);
and U9379 (N_9379,N_8821,N_8818);
nor U9380 (N_9380,N_8889,N_9186);
xnor U9381 (N_9381,N_9042,N_9160);
nand U9382 (N_9382,N_9078,N_8892);
nand U9383 (N_9383,N_8812,N_8890);
xor U9384 (N_9384,N_9118,N_9090);
nand U9385 (N_9385,N_9060,N_9055);
nor U9386 (N_9386,N_8953,N_8807);
nor U9387 (N_9387,N_9007,N_9061);
nor U9388 (N_9388,N_9145,N_9128);
xor U9389 (N_9389,N_8884,N_8891);
and U9390 (N_9390,N_9044,N_9087);
and U9391 (N_9391,N_9163,N_8831);
and U9392 (N_9392,N_9102,N_8942);
nand U9393 (N_9393,N_9002,N_8967);
or U9394 (N_9394,N_8835,N_8986);
nor U9395 (N_9395,N_8861,N_9123);
nand U9396 (N_9396,N_8983,N_9176);
xnor U9397 (N_9397,N_9167,N_8912);
nand U9398 (N_9398,N_9133,N_8829);
xnor U9399 (N_9399,N_8858,N_9177);
nor U9400 (N_9400,N_8880,N_8883);
xor U9401 (N_9401,N_9010,N_9102);
xor U9402 (N_9402,N_9055,N_8817);
or U9403 (N_9403,N_8863,N_9023);
and U9404 (N_9404,N_8857,N_8822);
xnor U9405 (N_9405,N_8998,N_9060);
nand U9406 (N_9406,N_8971,N_9031);
nor U9407 (N_9407,N_8988,N_9060);
or U9408 (N_9408,N_8867,N_8944);
or U9409 (N_9409,N_8817,N_8996);
xnor U9410 (N_9410,N_8874,N_9068);
nand U9411 (N_9411,N_9152,N_9161);
or U9412 (N_9412,N_8959,N_8957);
nor U9413 (N_9413,N_9178,N_9191);
nor U9414 (N_9414,N_9158,N_8892);
nor U9415 (N_9415,N_9051,N_8970);
nor U9416 (N_9416,N_8912,N_8992);
or U9417 (N_9417,N_9017,N_9047);
xnor U9418 (N_9418,N_8886,N_8971);
xor U9419 (N_9419,N_9141,N_9108);
or U9420 (N_9420,N_9074,N_8860);
nor U9421 (N_9421,N_8950,N_9173);
nor U9422 (N_9422,N_9040,N_8936);
and U9423 (N_9423,N_9092,N_8800);
or U9424 (N_9424,N_9040,N_8915);
xnor U9425 (N_9425,N_8818,N_9059);
nor U9426 (N_9426,N_9107,N_8843);
xor U9427 (N_9427,N_8968,N_8842);
nand U9428 (N_9428,N_8891,N_9040);
xnor U9429 (N_9429,N_9001,N_8875);
and U9430 (N_9430,N_9040,N_9033);
xnor U9431 (N_9431,N_8929,N_8916);
nand U9432 (N_9432,N_8888,N_8985);
nand U9433 (N_9433,N_9108,N_9084);
nor U9434 (N_9434,N_9042,N_8821);
nand U9435 (N_9435,N_9006,N_9196);
xnor U9436 (N_9436,N_8964,N_8921);
and U9437 (N_9437,N_8898,N_8966);
and U9438 (N_9438,N_9151,N_9070);
nor U9439 (N_9439,N_9168,N_9176);
nor U9440 (N_9440,N_9047,N_9148);
xor U9441 (N_9441,N_9074,N_8806);
xor U9442 (N_9442,N_8840,N_9005);
and U9443 (N_9443,N_9122,N_8947);
and U9444 (N_9444,N_9193,N_9037);
nor U9445 (N_9445,N_9139,N_9045);
nor U9446 (N_9446,N_8937,N_9193);
xnor U9447 (N_9447,N_9038,N_8886);
nor U9448 (N_9448,N_9093,N_8955);
or U9449 (N_9449,N_8953,N_8874);
xnor U9450 (N_9450,N_9162,N_8941);
nand U9451 (N_9451,N_8868,N_9054);
xnor U9452 (N_9452,N_8835,N_9093);
and U9453 (N_9453,N_8977,N_9019);
and U9454 (N_9454,N_9102,N_8887);
xor U9455 (N_9455,N_8902,N_8937);
xor U9456 (N_9456,N_9002,N_8846);
xor U9457 (N_9457,N_9168,N_8985);
and U9458 (N_9458,N_8965,N_9152);
or U9459 (N_9459,N_8930,N_8898);
nand U9460 (N_9460,N_9189,N_8970);
or U9461 (N_9461,N_9031,N_8903);
or U9462 (N_9462,N_9120,N_9183);
and U9463 (N_9463,N_9107,N_9070);
and U9464 (N_9464,N_9198,N_8872);
nor U9465 (N_9465,N_8832,N_9160);
or U9466 (N_9466,N_8985,N_8805);
and U9467 (N_9467,N_9036,N_9102);
nor U9468 (N_9468,N_8851,N_8988);
xnor U9469 (N_9469,N_8864,N_9159);
nand U9470 (N_9470,N_8815,N_8886);
nand U9471 (N_9471,N_9124,N_8934);
and U9472 (N_9472,N_9077,N_9173);
nor U9473 (N_9473,N_9001,N_9092);
nand U9474 (N_9474,N_8926,N_8903);
nand U9475 (N_9475,N_8920,N_9013);
or U9476 (N_9476,N_8905,N_8844);
xor U9477 (N_9477,N_9045,N_8894);
and U9478 (N_9478,N_9076,N_9081);
nand U9479 (N_9479,N_8943,N_8845);
xor U9480 (N_9480,N_8902,N_9151);
xnor U9481 (N_9481,N_9151,N_9130);
and U9482 (N_9482,N_8922,N_8940);
nor U9483 (N_9483,N_8973,N_9117);
or U9484 (N_9484,N_8917,N_8891);
nor U9485 (N_9485,N_9093,N_9000);
xnor U9486 (N_9486,N_8922,N_8929);
and U9487 (N_9487,N_8866,N_9013);
or U9488 (N_9488,N_8871,N_8996);
and U9489 (N_9489,N_9108,N_8809);
nor U9490 (N_9490,N_9155,N_9183);
nor U9491 (N_9491,N_9018,N_9140);
nor U9492 (N_9492,N_8957,N_8966);
and U9493 (N_9493,N_8867,N_8956);
and U9494 (N_9494,N_8950,N_8912);
nor U9495 (N_9495,N_9039,N_8951);
or U9496 (N_9496,N_9167,N_8999);
or U9497 (N_9497,N_8851,N_8940);
xor U9498 (N_9498,N_9117,N_8891);
xnor U9499 (N_9499,N_8834,N_9088);
xnor U9500 (N_9500,N_8888,N_9173);
or U9501 (N_9501,N_8991,N_8981);
nand U9502 (N_9502,N_8868,N_9175);
nor U9503 (N_9503,N_9135,N_8884);
and U9504 (N_9504,N_8885,N_8826);
xnor U9505 (N_9505,N_8978,N_9047);
nand U9506 (N_9506,N_9174,N_9159);
nor U9507 (N_9507,N_9043,N_9139);
or U9508 (N_9508,N_8862,N_8819);
nor U9509 (N_9509,N_8963,N_8823);
and U9510 (N_9510,N_8802,N_9035);
nor U9511 (N_9511,N_8880,N_9127);
and U9512 (N_9512,N_9067,N_9086);
and U9513 (N_9513,N_8980,N_9137);
xor U9514 (N_9514,N_8906,N_9199);
nand U9515 (N_9515,N_8938,N_9012);
or U9516 (N_9516,N_8927,N_9150);
nor U9517 (N_9517,N_9058,N_8803);
nor U9518 (N_9518,N_9150,N_8851);
nor U9519 (N_9519,N_8942,N_9143);
and U9520 (N_9520,N_8829,N_9042);
xor U9521 (N_9521,N_9140,N_8939);
xor U9522 (N_9522,N_8936,N_8863);
and U9523 (N_9523,N_8873,N_9122);
and U9524 (N_9524,N_9154,N_8979);
nand U9525 (N_9525,N_8857,N_9097);
nor U9526 (N_9526,N_9047,N_9108);
nand U9527 (N_9527,N_8924,N_8855);
xnor U9528 (N_9528,N_9118,N_8869);
and U9529 (N_9529,N_9019,N_8958);
nor U9530 (N_9530,N_8934,N_8817);
nand U9531 (N_9531,N_9092,N_8879);
nand U9532 (N_9532,N_9072,N_9074);
xnor U9533 (N_9533,N_9117,N_8818);
nand U9534 (N_9534,N_9073,N_9088);
or U9535 (N_9535,N_9049,N_8832);
nand U9536 (N_9536,N_8822,N_8853);
nand U9537 (N_9537,N_9155,N_9012);
and U9538 (N_9538,N_8803,N_9093);
nor U9539 (N_9539,N_9092,N_8843);
nor U9540 (N_9540,N_8952,N_9193);
nand U9541 (N_9541,N_9079,N_8998);
and U9542 (N_9542,N_9124,N_9156);
xor U9543 (N_9543,N_8943,N_9027);
and U9544 (N_9544,N_8966,N_8884);
or U9545 (N_9545,N_8932,N_8870);
nor U9546 (N_9546,N_9044,N_8888);
nand U9547 (N_9547,N_9142,N_9194);
nor U9548 (N_9548,N_9046,N_8858);
and U9549 (N_9549,N_9181,N_9081);
nor U9550 (N_9550,N_9055,N_8936);
or U9551 (N_9551,N_8959,N_8815);
nand U9552 (N_9552,N_9002,N_8817);
nor U9553 (N_9553,N_9133,N_8912);
nor U9554 (N_9554,N_8926,N_8992);
nor U9555 (N_9555,N_9073,N_9148);
xnor U9556 (N_9556,N_9001,N_9135);
xor U9557 (N_9557,N_9173,N_8925);
nor U9558 (N_9558,N_8856,N_8816);
xor U9559 (N_9559,N_9154,N_8941);
and U9560 (N_9560,N_9014,N_8835);
or U9561 (N_9561,N_8902,N_9065);
xor U9562 (N_9562,N_9096,N_8808);
xor U9563 (N_9563,N_8826,N_8886);
or U9564 (N_9564,N_8998,N_9121);
and U9565 (N_9565,N_8938,N_8971);
and U9566 (N_9566,N_8829,N_8991);
or U9567 (N_9567,N_8982,N_8974);
or U9568 (N_9568,N_8910,N_8855);
nor U9569 (N_9569,N_8953,N_9156);
or U9570 (N_9570,N_8925,N_9092);
nor U9571 (N_9571,N_9181,N_8979);
or U9572 (N_9572,N_9159,N_8940);
and U9573 (N_9573,N_9196,N_9121);
and U9574 (N_9574,N_9016,N_9029);
xor U9575 (N_9575,N_8837,N_9110);
nand U9576 (N_9576,N_8830,N_9020);
nor U9577 (N_9577,N_9177,N_9031);
or U9578 (N_9578,N_9129,N_8962);
nand U9579 (N_9579,N_8841,N_8920);
xnor U9580 (N_9580,N_8858,N_8808);
or U9581 (N_9581,N_9032,N_9083);
xor U9582 (N_9582,N_8959,N_8994);
nand U9583 (N_9583,N_8890,N_8901);
and U9584 (N_9584,N_9064,N_8890);
nand U9585 (N_9585,N_8873,N_8986);
nand U9586 (N_9586,N_8828,N_9061);
or U9587 (N_9587,N_9094,N_9100);
nand U9588 (N_9588,N_9085,N_8932);
nor U9589 (N_9589,N_9043,N_8982);
xor U9590 (N_9590,N_9170,N_8891);
or U9591 (N_9591,N_8942,N_8979);
nor U9592 (N_9592,N_8952,N_8949);
nand U9593 (N_9593,N_9128,N_8823);
and U9594 (N_9594,N_9013,N_9190);
nand U9595 (N_9595,N_9047,N_9130);
and U9596 (N_9596,N_9092,N_9192);
or U9597 (N_9597,N_9114,N_9105);
or U9598 (N_9598,N_9015,N_8902);
nand U9599 (N_9599,N_8990,N_9148);
or U9600 (N_9600,N_9505,N_9212);
or U9601 (N_9601,N_9421,N_9492);
nor U9602 (N_9602,N_9310,N_9217);
or U9603 (N_9603,N_9339,N_9228);
or U9604 (N_9604,N_9257,N_9457);
or U9605 (N_9605,N_9236,N_9334);
xor U9606 (N_9606,N_9405,N_9379);
nor U9607 (N_9607,N_9277,N_9521);
xor U9608 (N_9608,N_9571,N_9420);
nor U9609 (N_9609,N_9254,N_9592);
xnor U9610 (N_9610,N_9483,N_9263);
or U9611 (N_9611,N_9222,N_9253);
nor U9612 (N_9612,N_9301,N_9302);
or U9613 (N_9613,N_9518,N_9230);
nor U9614 (N_9614,N_9359,N_9364);
nor U9615 (N_9615,N_9308,N_9312);
or U9616 (N_9616,N_9495,N_9373);
nor U9617 (N_9617,N_9344,N_9535);
xor U9618 (N_9618,N_9557,N_9270);
nor U9619 (N_9619,N_9482,N_9210);
or U9620 (N_9620,N_9259,N_9260);
xnor U9621 (N_9621,N_9543,N_9423);
xnor U9622 (N_9622,N_9218,N_9320);
nand U9623 (N_9623,N_9425,N_9584);
xnor U9624 (N_9624,N_9589,N_9407);
nand U9625 (N_9625,N_9241,N_9568);
xnor U9626 (N_9626,N_9328,N_9374);
xnor U9627 (N_9627,N_9295,N_9509);
xnor U9628 (N_9628,N_9243,N_9501);
or U9629 (N_9629,N_9479,N_9352);
nor U9630 (N_9630,N_9264,N_9498);
nand U9631 (N_9631,N_9341,N_9544);
xor U9632 (N_9632,N_9316,N_9299);
nand U9633 (N_9633,N_9569,N_9473);
nor U9634 (N_9634,N_9465,N_9394);
xnor U9635 (N_9635,N_9456,N_9413);
xnor U9636 (N_9636,N_9377,N_9271);
nand U9637 (N_9637,N_9224,N_9343);
or U9638 (N_9638,N_9350,N_9239);
xor U9639 (N_9639,N_9381,N_9404);
xor U9640 (N_9640,N_9220,N_9366);
xnor U9641 (N_9641,N_9315,N_9294);
nand U9642 (N_9642,N_9219,N_9356);
nand U9643 (N_9643,N_9207,N_9494);
nand U9644 (N_9644,N_9227,N_9371);
and U9645 (N_9645,N_9208,N_9461);
nor U9646 (N_9646,N_9347,N_9558);
or U9647 (N_9647,N_9434,N_9332);
nor U9648 (N_9648,N_9386,N_9522);
nand U9649 (N_9649,N_9551,N_9281);
or U9650 (N_9650,N_9297,N_9417);
nand U9651 (N_9651,N_9506,N_9318);
xnor U9652 (N_9652,N_9231,N_9240);
nand U9653 (N_9653,N_9337,N_9256);
nor U9654 (N_9654,N_9365,N_9519);
or U9655 (N_9655,N_9470,N_9403);
and U9656 (N_9656,N_9205,N_9504);
and U9657 (N_9657,N_9431,N_9398);
and U9658 (N_9658,N_9586,N_9575);
and U9659 (N_9659,N_9293,N_9440);
or U9660 (N_9660,N_9533,N_9346);
nor U9661 (N_9661,N_9393,N_9242);
xor U9662 (N_9662,N_9562,N_9396);
and U9663 (N_9663,N_9276,N_9532);
nand U9664 (N_9664,N_9438,N_9587);
and U9665 (N_9665,N_9499,N_9285);
nand U9666 (N_9666,N_9237,N_9355);
nor U9667 (N_9667,N_9553,N_9454);
nand U9668 (N_9668,N_9211,N_9303);
nand U9669 (N_9669,N_9561,N_9530);
and U9670 (N_9670,N_9527,N_9515);
or U9671 (N_9671,N_9591,N_9500);
or U9672 (N_9672,N_9323,N_9460);
nand U9673 (N_9673,N_9367,N_9573);
and U9674 (N_9674,N_9448,N_9202);
xnor U9675 (N_9675,N_9549,N_9594);
and U9676 (N_9676,N_9471,N_9455);
nand U9677 (N_9677,N_9472,N_9552);
and U9678 (N_9678,N_9432,N_9349);
nand U9679 (N_9679,N_9399,N_9424);
nor U9680 (N_9680,N_9249,N_9574);
or U9681 (N_9681,N_9478,N_9468);
nand U9682 (N_9682,N_9266,N_9528);
or U9683 (N_9683,N_9416,N_9524);
and U9684 (N_9684,N_9255,N_9516);
xnor U9685 (N_9685,N_9542,N_9588);
xnor U9686 (N_9686,N_9261,N_9246);
nand U9687 (N_9687,N_9289,N_9306);
nor U9688 (N_9688,N_9436,N_9272);
nor U9689 (N_9689,N_9520,N_9340);
nor U9690 (N_9690,N_9229,N_9375);
nand U9691 (N_9691,N_9362,N_9363);
and U9692 (N_9692,N_9251,N_9410);
or U9693 (N_9693,N_9428,N_9313);
nand U9694 (N_9694,N_9376,N_9369);
nor U9695 (N_9695,N_9545,N_9389);
xnor U9696 (N_9696,N_9225,N_9469);
xor U9697 (N_9697,N_9579,N_9464);
and U9698 (N_9698,N_9331,N_9433);
nor U9699 (N_9699,N_9409,N_9514);
nor U9700 (N_9700,N_9226,N_9269);
nand U9701 (N_9701,N_9203,N_9564);
or U9702 (N_9702,N_9444,N_9508);
nand U9703 (N_9703,N_9353,N_9556);
xor U9704 (N_9704,N_9201,N_9493);
nor U9705 (N_9705,N_9419,N_9548);
xor U9706 (N_9706,N_9422,N_9442);
xnor U9707 (N_9707,N_9370,N_9491);
and U9708 (N_9708,N_9597,N_9248);
or U9709 (N_9709,N_9384,N_9290);
nor U9710 (N_9710,N_9372,N_9412);
and U9711 (N_9711,N_9443,N_9354);
xor U9712 (N_9712,N_9439,N_9582);
or U9713 (N_9713,N_9392,N_9283);
nor U9714 (N_9714,N_9475,N_9547);
or U9715 (N_9715,N_9590,N_9262);
xor U9716 (N_9716,N_9342,N_9247);
or U9717 (N_9717,N_9538,N_9480);
nand U9718 (N_9718,N_9467,N_9383);
or U9719 (N_9719,N_9387,N_9311);
nand U9720 (N_9720,N_9517,N_9279);
nor U9721 (N_9721,N_9487,N_9599);
xor U9722 (N_9722,N_9529,N_9450);
or U9723 (N_9723,N_9477,N_9512);
xnor U9724 (N_9724,N_9280,N_9577);
nand U9725 (N_9725,N_9485,N_9305);
nand U9726 (N_9726,N_9567,N_9572);
nand U9727 (N_9727,N_9513,N_9486);
or U9728 (N_9728,N_9348,N_9496);
nor U9729 (N_9729,N_9488,N_9463);
xnor U9730 (N_9730,N_9304,N_9510);
nor U9731 (N_9731,N_9531,N_9282);
nand U9732 (N_9732,N_9546,N_9418);
nor U9733 (N_9733,N_9447,N_9335);
nand U9734 (N_9734,N_9274,N_9278);
xnor U9735 (N_9735,N_9391,N_9245);
nor U9736 (N_9736,N_9415,N_9292);
and U9737 (N_9737,N_9361,N_9559);
xnor U9738 (N_9738,N_9451,N_9252);
and U9739 (N_9739,N_9336,N_9200);
or U9740 (N_9740,N_9214,N_9523);
and U9741 (N_9741,N_9430,N_9595);
or U9742 (N_9742,N_9581,N_9576);
and U9743 (N_9743,N_9435,N_9284);
xor U9744 (N_9744,N_9265,N_9233);
and U9745 (N_9745,N_9206,N_9325);
nand U9746 (N_9746,N_9484,N_9497);
nand U9747 (N_9747,N_9503,N_9296);
xor U9748 (N_9748,N_9400,N_9429);
nor U9749 (N_9749,N_9390,N_9322);
or U9750 (N_9750,N_9244,N_9250);
nand U9751 (N_9751,N_9388,N_9580);
or U9752 (N_9752,N_9273,N_9570);
or U9753 (N_9753,N_9402,N_9489);
and U9754 (N_9754,N_9314,N_9401);
nand U9755 (N_9755,N_9446,N_9327);
nand U9756 (N_9756,N_9540,N_9534);
xor U9757 (N_9757,N_9298,N_9525);
and U9758 (N_9758,N_9502,N_9541);
nand U9759 (N_9759,N_9406,N_9330);
nor U9760 (N_9760,N_9357,N_9449);
nor U9761 (N_9761,N_9490,N_9397);
or U9762 (N_9762,N_9324,N_9267);
and U9763 (N_9763,N_9452,N_9459);
or U9764 (N_9764,N_9286,N_9466);
xnor U9765 (N_9765,N_9596,N_9204);
and U9766 (N_9766,N_9317,N_9287);
xnor U9767 (N_9767,N_9445,N_9300);
and U9768 (N_9768,N_9382,N_9593);
or U9769 (N_9769,N_9481,N_9234);
xnor U9770 (N_9770,N_9326,N_9351);
xnor U9771 (N_9771,N_9550,N_9360);
nor U9772 (N_9772,N_9319,N_9539);
xor U9773 (N_9773,N_9345,N_9560);
and U9774 (N_9774,N_9235,N_9441);
xor U9775 (N_9775,N_9458,N_9566);
nand U9776 (N_9776,N_9338,N_9537);
nor U9777 (N_9777,N_9309,N_9291);
xor U9778 (N_9778,N_9358,N_9380);
and U9779 (N_9779,N_9507,N_9215);
xnor U9780 (N_9780,N_9526,N_9378);
and U9781 (N_9781,N_9563,N_9511);
and U9782 (N_9782,N_9275,N_9213);
nor U9783 (N_9783,N_9258,N_9209);
nand U9784 (N_9784,N_9307,N_9268);
or U9785 (N_9785,N_9321,N_9555);
or U9786 (N_9786,N_9462,N_9414);
or U9787 (N_9787,N_9411,N_9333);
nand U9788 (N_9788,N_9554,N_9221);
xnor U9789 (N_9789,N_9453,N_9474);
xor U9790 (N_9790,N_9598,N_9583);
xnor U9791 (N_9791,N_9536,N_9427);
and U9792 (N_9792,N_9585,N_9437);
nor U9793 (N_9793,N_9426,N_9565);
or U9794 (N_9794,N_9288,N_9216);
or U9795 (N_9795,N_9476,N_9578);
nand U9796 (N_9796,N_9385,N_9223);
and U9797 (N_9797,N_9368,N_9238);
nor U9798 (N_9798,N_9408,N_9232);
xor U9799 (N_9799,N_9395,N_9329);
or U9800 (N_9800,N_9344,N_9516);
or U9801 (N_9801,N_9368,N_9418);
xor U9802 (N_9802,N_9539,N_9410);
and U9803 (N_9803,N_9553,N_9219);
and U9804 (N_9804,N_9542,N_9592);
nor U9805 (N_9805,N_9250,N_9487);
and U9806 (N_9806,N_9497,N_9204);
nor U9807 (N_9807,N_9253,N_9316);
or U9808 (N_9808,N_9409,N_9414);
and U9809 (N_9809,N_9392,N_9304);
and U9810 (N_9810,N_9553,N_9319);
xnor U9811 (N_9811,N_9592,N_9429);
nor U9812 (N_9812,N_9391,N_9451);
xnor U9813 (N_9813,N_9228,N_9593);
or U9814 (N_9814,N_9352,N_9375);
and U9815 (N_9815,N_9253,N_9460);
xor U9816 (N_9816,N_9484,N_9588);
nor U9817 (N_9817,N_9480,N_9341);
xor U9818 (N_9818,N_9588,N_9270);
xor U9819 (N_9819,N_9475,N_9598);
or U9820 (N_9820,N_9200,N_9595);
xnor U9821 (N_9821,N_9346,N_9374);
nor U9822 (N_9822,N_9258,N_9560);
xor U9823 (N_9823,N_9382,N_9246);
nor U9824 (N_9824,N_9578,N_9562);
or U9825 (N_9825,N_9298,N_9570);
and U9826 (N_9826,N_9579,N_9347);
xor U9827 (N_9827,N_9584,N_9210);
xnor U9828 (N_9828,N_9367,N_9397);
nand U9829 (N_9829,N_9325,N_9505);
or U9830 (N_9830,N_9311,N_9390);
or U9831 (N_9831,N_9259,N_9343);
or U9832 (N_9832,N_9389,N_9399);
and U9833 (N_9833,N_9261,N_9317);
nand U9834 (N_9834,N_9385,N_9379);
xnor U9835 (N_9835,N_9388,N_9299);
and U9836 (N_9836,N_9306,N_9246);
nor U9837 (N_9837,N_9525,N_9505);
or U9838 (N_9838,N_9440,N_9422);
nor U9839 (N_9839,N_9594,N_9336);
or U9840 (N_9840,N_9219,N_9390);
nand U9841 (N_9841,N_9396,N_9261);
nor U9842 (N_9842,N_9273,N_9300);
and U9843 (N_9843,N_9529,N_9425);
nor U9844 (N_9844,N_9565,N_9321);
xnor U9845 (N_9845,N_9479,N_9372);
or U9846 (N_9846,N_9548,N_9476);
or U9847 (N_9847,N_9466,N_9421);
nand U9848 (N_9848,N_9396,N_9462);
and U9849 (N_9849,N_9567,N_9389);
nor U9850 (N_9850,N_9270,N_9429);
xnor U9851 (N_9851,N_9555,N_9269);
or U9852 (N_9852,N_9361,N_9374);
nor U9853 (N_9853,N_9335,N_9477);
nand U9854 (N_9854,N_9325,N_9484);
and U9855 (N_9855,N_9225,N_9213);
xnor U9856 (N_9856,N_9458,N_9348);
or U9857 (N_9857,N_9476,N_9326);
and U9858 (N_9858,N_9348,N_9277);
nor U9859 (N_9859,N_9219,N_9322);
or U9860 (N_9860,N_9332,N_9213);
xor U9861 (N_9861,N_9380,N_9405);
and U9862 (N_9862,N_9397,N_9539);
or U9863 (N_9863,N_9363,N_9293);
and U9864 (N_9864,N_9465,N_9548);
xor U9865 (N_9865,N_9339,N_9290);
nand U9866 (N_9866,N_9251,N_9498);
and U9867 (N_9867,N_9238,N_9396);
nand U9868 (N_9868,N_9493,N_9272);
nor U9869 (N_9869,N_9395,N_9401);
nand U9870 (N_9870,N_9378,N_9579);
or U9871 (N_9871,N_9277,N_9525);
nor U9872 (N_9872,N_9349,N_9287);
and U9873 (N_9873,N_9525,N_9396);
nand U9874 (N_9874,N_9399,N_9441);
or U9875 (N_9875,N_9545,N_9573);
xnor U9876 (N_9876,N_9336,N_9229);
nand U9877 (N_9877,N_9545,N_9329);
nand U9878 (N_9878,N_9585,N_9386);
xnor U9879 (N_9879,N_9556,N_9256);
nor U9880 (N_9880,N_9369,N_9268);
and U9881 (N_9881,N_9404,N_9565);
or U9882 (N_9882,N_9466,N_9461);
and U9883 (N_9883,N_9251,N_9589);
and U9884 (N_9884,N_9310,N_9200);
xnor U9885 (N_9885,N_9595,N_9286);
or U9886 (N_9886,N_9269,N_9543);
and U9887 (N_9887,N_9599,N_9581);
nor U9888 (N_9888,N_9289,N_9371);
or U9889 (N_9889,N_9471,N_9349);
and U9890 (N_9890,N_9466,N_9249);
xor U9891 (N_9891,N_9520,N_9595);
and U9892 (N_9892,N_9467,N_9244);
nand U9893 (N_9893,N_9234,N_9496);
nand U9894 (N_9894,N_9592,N_9227);
or U9895 (N_9895,N_9267,N_9226);
nor U9896 (N_9896,N_9221,N_9428);
nand U9897 (N_9897,N_9308,N_9404);
and U9898 (N_9898,N_9585,N_9380);
or U9899 (N_9899,N_9281,N_9530);
or U9900 (N_9900,N_9392,N_9558);
or U9901 (N_9901,N_9276,N_9517);
nand U9902 (N_9902,N_9520,N_9497);
nor U9903 (N_9903,N_9443,N_9205);
nand U9904 (N_9904,N_9387,N_9576);
or U9905 (N_9905,N_9570,N_9228);
nand U9906 (N_9906,N_9288,N_9268);
nor U9907 (N_9907,N_9336,N_9385);
and U9908 (N_9908,N_9354,N_9554);
and U9909 (N_9909,N_9309,N_9232);
xor U9910 (N_9910,N_9265,N_9510);
nor U9911 (N_9911,N_9344,N_9341);
and U9912 (N_9912,N_9476,N_9465);
nor U9913 (N_9913,N_9321,N_9235);
nand U9914 (N_9914,N_9471,N_9277);
nor U9915 (N_9915,N_9231,N_9511);
or U9916 (N_9916,N_9431,N_9488);
nand U9917 (N_9917,N_9374,N_9298);
or U9918 (N_9918,N_9396,N_9385);
nor U9919 (N_9919,N_9561,N_9492);
xnor U9920 (N_9920,N_9403,N_9359);
xor U9921 (N_9921,N_9563,N_9575);
or U9922 (N_9922,N_9357,N_9433);
or U9923 (N_9923,N_9473,N_9490);
or U9924 (N_9924,N_9453,N_9269);
and U9925 (N_9925,N_9316,N_9516);
nand U9926 (N_9926,N_9365,N_9317);
nor U9927 (N_9927,N_9357,N_9239);
or U9928 (N_9928,N_9595,N_9582);
nand U9929 (N_9929,N_9519,N_9439);
or U9930 (N_9930,N_9381,N_9583);
nand U9931 (N_9931,N_9371,N_9281);
nor U9932 (N_9932,N_9495,N_9542);
or U9933 (N_9933,N_9432,N_9582);
xor U9934 (N_9934,N_9324,N_9483);
xor U9935 (N_9935,N_9482,N_9545);
or U9936 (N_9936,N_9227,N_9463);
or U9937 (N_9937,N_9480,N_9254);
and U9938 (N_9938,N_9534,N_9200);
nand U9939 (N_9939,N_9372,N_9284);
or U9940 (N_9940,N_9471,N_9556);
or U9941 (N_9941,N_9495,N_9455);
nor U9942 (N_9942,N_9488,N_9272);
xnor U9943 (N_9943,N_9509,N_9330);
xor U9944 (N_9944,N_9258,N_9427);
nor U9945 (N_9945,N_9493,N_9576);
and U9946 (N_9946,N_9270,N_9345);
and U9947 (N_9947,N_9312,N_9358);
xnor U9948 (N_9948,N_9258,N_9525);
or U9949 (N_9949,N_9544,N_9371);
nor U9950 (N_9950,N_9486,N_9447);
xor U9951 (N_9951,N_9471,N_9257);
and U9952 (N_9952,N_9313,N_9420);
nand U9953 (N_9953,N_9484,N_9464);
xnor U9954 (N_9954,N_9347,N_9260);
or U9955 (N_9955,N_9502,N_9424);
and U9956 (N_9956,N_9460,N_9330);
or U9957 (N_9957,N_9404,N_9554);
xor U9958 (N_9958,N_9511,N_9557);
or U9959 (N_9959,N_9414,N_9474);
xnor U9960 (N_9960,N_9532,N_9422);
xnor U9961 (N_9961,N_9218,N_9371);
xor U9962 (N_9962,N_9264,N_9540);
nor U9963 (N_9963,N_9433,N_9439);
xnor U9964 (N_9964,N_9466,N_9487);
nand U9965 (N_9965,N_9337,N_9249);
nand U9966 (N_9966,N_9319,N_9308);
and U9967 (N_9967,N_9410,N_9519);
xor U9968 (N_9968,N_9520,N_9282);
xnor U9969 (N_9969,N_9521,N_9308);
nor U9970 (N_9970,N_9237,N_9411);
xor U9971 (N_9971,N_9562,N_9502);
xor U9972 (N_9972,N_9265,N_9406);
xor U9973 (N_9973,N_9260,N_9220);
nand U9974 (N_9974,N_9250,N_9459);
or U9975 (N_9975,N_9255,N_9213);
nand U9976 (N_9976,N_9513,N_9445);
and U9977 (N_9977,N_9351,N_9223);
xor U9978 (N_9978,N_9312,N_9594);
and U9979 (N_9979,N_9447,N_9238);
xnor U9980 (N_9980,N_9596,N_9468);
and U9981 (N_9981,N_9374,N_9318);
nor U9982 (N_9982,N_9325,N_9318);
nor U9983 (N_9983,N_9292,N_9255);
nor U9984 (N_9984,N_9245,N_9436);
and U9985 (N_9985,N_9332,N_9354);
nor U9986 (N_9986,N_9374,N_9440);
nand U9987 (N_9987,N_9211,N_9207);
or U9988 (N_9988,N_9529,N_9361);
and U9989 (N_9989,N_9395,N_9320);
and U9990 (N_9990,N_9569,N_9422);
nand U9991 (N_9991,N_9224,N_9368);
nand U9992 (N_9992,N_9207,N_9212);
xor U9993 (N_9993,N_9369,N_9347);
xnor U9994 (N_9994,N_9476,N_9482);
nand U9995 (N_9995,N_9328,N_9241);
xnor U9996 (N_9996,N_9380,N_9287);
xor U9997 (N_9997,N_9377,N_9201);
or U9998 (N_9998,N_9257,N_9588);
or U9999 (N_9999,N_9367,N_9209);
xnor U10000 (N_10000,N_9982,N_9796);
nand U10001 (N_10001,N_9923,N_9661);
xnor U10002 (N_10002,N_9724,N_9673);
nand U10003 (N_10003,N_9972,N_9660);
nor U10004 (N_10004,N_9784,N_9983);
or U10005 (N_10005,N_9817,N_9685);
or U10006 (N_10006,N_9688,N_9678);
and U10007 (N_10007,N_9895,N_9606);
nor U10008 (N_10008,N_9691,N_9966);
nor U10009 (N_10009,N_9870,N_9651);
or U10010 (N_10010,N_9931,N_9632);
nand U10011 (N_10011,N_9903,N_9755);
xor U10012 (N_10012,N_9937,N_9797);
xor U10013 (N_10013,N_9643,N_9863);
nand U10014 (N_10014,N_9674,N_9837);
nor U10015 (N_10015,N_9648,N_9749);
xnor U10016 (N_10016,N_9991,N_9615);
and U10017 (N_10017,N_9910,N_9786);
or U10018 (N_10018,N_9791,N_9682);
xor U10019 (N_10019,N_9725,N_9709);
and U10020 (N_10020,N_9919,N_9841);
xnor U10021 (N_10021,N_9741,N_9757);
nor U10022 (N_10022,N_9974,N_9962);
nand U10023 (N_10023,N_9617,N_9622);
and U10024 (N_10024,N_9888,N_9640);
or U10025 (N_10025,N_9732,N_9911);
or U10026 (N_10026,N_9917,N_9902);
or U10027 (N_10027,N_9747,N_9835);
nor U10028 (N_10028,N_9879,N_9627);
nand U10029 (N_10029,N_9806,N_9853);
nand U10030 (N_10030,N_9812,N_9948);
xnor U10031 (N_10031,N_9975,N_9956);
and U10032 (N_10032,N_9666,N_9996);
nand U10033 (N_10033,N_9920,N_9668);
xor U10034 (N_10034,N_9713,N_9623);
or U10035 (N_10035,N_9718,N_9953);
nor U10036 (N_10036,N_9838,N_9930);
nand U10037 (N_10037,N_9828,N_9631);
xnor U10038 (N_10038,N_9669,N_9932);
nand U10039 (N_10039,N_9899,N_9868);
and U10040 (N_10040,N_9612,N_9787);
or U10041 (N_10041,N_9773,N_9613);
nand U10042 (N_10042,N_9778,N_9915);
and U10043 (N_10043,N_9922,N_9820);
nor U10044 (N_10044,N_9827,N_9601);
nor U10045 (N_10045,N_9859,N_9811);
and U10046 (N_10046,N_9849,N_9637);
nand U10047 (N_10047,N_9605,N_9866);
nor U10048 (N_10048,N_9720,N_9715);
xnor U10049 (N_10049,N_9973,N_9958);
nand U10050 (N_10050,N_9881,N_9940);
nand U10051 (N_10051,N_9843,N_9743);
xnor U10052 (N_10052,N_9738,N_9967);
nand U10053 (N_10053,N_9672,N_9816);
xor U10054 (N_10054,N_9885,N_9933);
nand U10055 (N_10055,N_9663,N_9847);
nand U10056 (N_10056,N_9742,N_9705);
nand U10057 (N_10057,N_9833,N_9886);
xnor U10058 (N_10058,N_9684,N_9670);
and U10059 (N_10059,N_9675,N_9610);
nand U10060 (N_10060,N_9927,N_9768);
nand U10061 (N_10061,N_9943,N_9883);
or U10062 (N_10062,N_9830,N_9657);
nor U10063 (N_10063,N_9769,N_9760);
xnor U10064 (N_10064,N_9746,N_9620);
xnor U10065 (N_10065,N_9790,N_9862);
nand U10066 (N_10066,N_9751,N_9665);
xnor U10067 (N_10067,N_9635,N_9950);
xor U10068 (N_10068,N_9698,N_9887);
xnor U10069 (N_10069,N_9770,N_9716);
nand U10070 (N_10070,N_9604,N_9602);
xor U10071 (N_10071,N_9653,N_9714);
and U10072 (N_10072,N_9947,N_9628);
and U10073 (N_10073,N_9979,N_9845);
nor U10074 (N_10074,N_9638,N_9999);
or U10075 (N_10075,N_9865,N_9977);
nand U10076 (N_10076,N_9926,N_9782);
xor U10077 (N_10077,N_9736,N_9880);
xnor U10078 (N_10078,N_9846,N_9608);
nor U10079 (N_10079,N_9871,N_9916);
nand U10080 (N_10080,N_9856,N_9968);
or U10081 (N_10081,N_9803,N_9614);
nand U10082 (N_10082,N_9683,N_9925);
xnor U10083 (N_10083,N_9644,N_9810);
nand U10084 (N_10084,N_9619,N_9783);
xnor U10085 (N_10085,N_9831,N_9904);
nand U10086 (N_10086,N_9789,N_9763);
nand U10087 (N_10087,N_9706,N_9609);
xnor U10088 (N_10088,N_9961,N_9658);
and U10089 (N_10089,N_9794,N_9985);
nand U10090 (N_10090,N_9677,N_9681);
xor U10091 (N_10091,N_9938,N_9825);
xor U10092 (N_10092,N_9744,N_9703);
or U10093 (N_10093,N_9707,N_9824);
nor U10094 (N_10094,N_9992,N_9805);
xor U10095 (N_10095,N_9779,N_9689);
nand U10096 (N_10096,N_9995,N_9819);
nor U10097 (N_10097,N_9727,N_9872);
nand U10098 (N_10098,N_9801,N_9955);
nor U10099 (N_10099,N_9890,N_9893);
xnor U10100 (N_10100,N_9739,N_9944);
xnor U10101 (N_10101,N_9799,N_9659);
or U10102 (N_10102,N_9717,N_9735);
or U10103 (N_10103,N_9884,N_9882);
and U10104 (N_10104,N_9892,N_9981);
and U10105 (N_10105,N_9891,N_9662);
nand U10106 (N_10106,N_9873,N_9945);
or U10107 (N_10107,N_9936,N_9800);
xnor U10108 (N_10108,N_9792,N_9700);
nor U10109 (N_10109,N_9629,N_9645);
nor U10110 (N_10110,N_9696,N_9775);
or U10111 (N_10111,N_9752,N_9952);
nand U10112 (N_10112,N_9624,N_9804);
nor U10113 (N_10113,N_9699,N_9785);
and U10114 (N_10114,N_9721,N_9864);
nand U10115 (N_10115,N_9914,N_9924);
or U10116 (N_10116,N_9776,N_9711);
or U10117 (N_10117,N_9733,N_9951);
and U10118 (N_10118,N_9802,N_9878);
and U10119 (N_10119,N_9679,N_9842);
or U10120 (N_10120,N_9896,N_9836);
xor U10121 (N_10121,N_9928,N_9909);
and U10122 (N_10122,N_9877,N_9965);
xor U10123 (N_10123,N_9858,N_9946);
or U10124 (N_10124,N_9823,N_9852);
and U10125 (N_10125,N_9913,N_9647);
xnor U10126 (N_10126,N_9694,N_9772);
or U10127 (N_10127,N_9758,N_9636);
and U10128 (N_10128,N_9963,N_9834);
nand U10129 (N_10129,N_9600,N_9997);
nand U10130 (N_10130,N_9667,N_9702);
nand U10131 (N_10131,N_9633,N_9740);
and U10132 (N_10132,N_9993,N_9701);
nor U10133 (N_10133,N_9687,N_9754);
xnor U10134 (N_10134,N_9690,N_9656);
xor U10135 (N_10135,N_9867,N_9625);
xnor U10136 (N_10136,N_9756,N_9994);
xnor U10137 (N_10137,N_9618,N_9848);
nor U10138 (N_10138,N_9897,N_9611);
and U10139 (N_10139,N_9616,N_9971);
xor U10140 (N_10140,N_9861,N_9771);
nand U10141 (N_10141,N_9822,N_9730);
nor U10142 (N_10142,N_9989,N_9839);
nor U10143 (N_10143,N_9998,N_9765);
or U10144 (N_10144,N_9652,N_9813);
or U10145 (N_10145,N_9621,N_9815);
or U10146 (N_10146,N_9844,N_9649);
and U10147 (N_10147,N_9808,N_9646);
xnor U10148 (N_10148,N_9874,N_9697);
nand U10149 (N_10149,N_9764,N_9942);
nor U10150 (N_10150,N_9762,N_9704);
nor U10151 (N_10151,N_9807,N_9729);
and U10152 (N_10152,N_9726,N_9767);
or U10153 (N_10153,N_9650,N_9719);
xor U10154 (N_10154,N_9869,N_9712);
nor U10155 (N_10155,N_9990,N_9680);
nor U10156 (N_10156,N_9607,N_9960);
or U10157 (N_10157,N_9723,N_9978);
or U10158 (N_10158,N_9639,N_9686);
or U10159 (N_10159,N_9759,N_9780);
nand U10160 (N_10160,N_9954,N_9821);
nand U10161 (N_10161,N_9626,N_9798);
nand U10162 (N_10162,N_9964,N_9753);
nor U10163 (N_10163,N_9722,N_9901);
nand U10164 (N_10164,N_9850,N_9898);
xnor U10165 (N_10165,N_9832,N_9777);
and U10166 (N_10166,N_9671,N_9788);
nor U10167 (N_10167,N_9634,N_9818);
xnor U10168 (N_10168,N_9900,N_9934);
xor U10169 (N_10169,N_9854,N_9766);
nand U10170 (N_10170,N_9876,N_9957);
nand U10171 (N_10171,N_9695,N_9908);
or U10172 (N_10172,N_9949,N_9929);
and U10173 (N_10173,N_9855,N_9745);
xnor U10174 (N_10174,N_9921,N_9980);
nand U10175 (N_10175,N_9970,N_9781);
xor U10176 (N_10176,N_9814,N_9935);
nor U10177 (N_10177,N_9603,N_9986);
and U10178 (N_10178,N_9907,N_9793);
and U10179 (N_10179,N_9710,N_9976);
nor U10180 (N_10180,N_9641,N_9664);
xor U10181 (N_10181,N_9728,N_9795);
or U10182 (N_10182,N_9988,N_9959);
or U10183 (N_10183,N_9987,N_9774);
nor U10184 (N_10184,N_9889,N_9860);
xor U10185 (N_10185,N_9918,N_9693);
xor U10186 (N_10186,N_9731,N_9894);
and U10187 (N_10187,N_9761,N_9737);
nand U10188 (N_10188,N_9748,N_9750);
and U10189 (N_10189,N_9984,N_9809);
and U10190 (N_10190,N_9840,N_9829);
and U10191 (N_10191,N_9655,N_9912);
nor U10192 (N_10192,N_9939,N_9941);
or U10193 (N_10193,N_9905,N_9851);
xnor U10194 (N_10194,N_9969,N_9676);
xnor U10195 (N_10195,N_9642,N_9654);
nor U10196 (N_10196,N_9630,N_9692);
nand U10197 (N_10197,N_9875,N_9826);
or U10198 (N_10198,N_9708,N_9734);
nand U10199 (N_10199,N_9857,N_9906);
nand U10200 (N_10200,N_9830,N_9730);
or U10201 (N_10201,N_9913,N_9626);
xor U10202 (N_10202,N_9813,N_9785);
xnor U10203 (N_10203,N_9963,N_9642);
or U10204 (N_10204,N_9792,N_9644);
xnor U10205 (N_10205,N_9861,N_9921);
or U10206 (N_10206,N_9934,N_9775);
nor U10207 (N_10207,N_9957,N_9687);
nor U10208 (N_10208,N_9617,N_9763);
nor U10209 (N_10209,N_9745,N_9632);
xor U10210 (N_10210,N_9674,N_9845);
nor U10211 (N_10211,N_9797,N_9924);
nand U10212 (N_10212,N_9682,N_9619);
or U10213 (N_10213,N_9864,N_9910);
nand U10214 (N_10214,N_9991,N_9715);
nor U10215 (N_10215,N_9836,N_9785);
xor U10216 (N_10216,N_9714,N_9606);
xor U10217 (N_10217,N_9897,N_9971);
xor U10218 (N_10218,N_9822,N_9889);
and U10219 (N_10219,N_9717,N_9795);
or U10220 (N_10220,N_9836,N_9916);
xnor U10221 (N_10221,N_9769,N_9960);
and U10222 (N_10222,N_9673,N_9766);
nor U10223 (N_10223,N_9805,N_9681);
or U10224 (N_10224,N_9639,N_9723);
nand U10225 (N_10225,N_9908,N_9699);
nand U10226 (N_10226,N_9649,N_9652);
or U10227 (N_10227,N_9902,N_9633);
nand U10228 (N_10228,N_9969,N_9844);
and U10229 (N_10229,N_9682,N_9768);
xnor U10230 (N_10230,N_9910,N_9663);
and U10231 (N_10231,N_9856,N_9965);
and U10232 (N_10232,N_9763,N_9720);
or U10233 (N_10233,N_9716,N_9682);
nand U10234 (N_10234,N_9736,N_9754);
nor U10235 (N_10235,N_9963,N_9903);
nand U10236 (N_10236,N_9856,N_9916);
xnor U10237 (N_10237,N_9930,N_9976);
and U10238 (N_10238,N_9822,N_9648);
xor U10239 (N_10239,N_9681,N_9717);
and U10240 (N_10240,N_9779,N_9687);
nand U10241 (N_10241,N_9987,N_9670);
nand U10242 (N_10242,N_9782,N_9977);
or U10243 (N_10243,N_9668,N_9937);
nand U10244 (N_10244,N_9611,N_9641);
or U10245 (N_10245,N_9814,N_9739);
nor U10246 (N_10246,N_9622,N_9952);
nand U10247 (N_10247,N_9908,N_9688);
or U10248 (N_10248,N_9806,N_9914);
and U10249 (N_10249,N_9957,N_9721);
and U10250 (N_10250,N_9667,N_9615);
nor U10251 (N_10251,N_9700,N_9923);
and U10252 (N_10252,N_9909,N_9788);
xor U10253 (N_10253,N_9679,N_9992);
nand U10254 (N_10254,N_9657,N_9868);
nor U10255 (N_10255,N_9934,N_9812);
and U10256 (N_10256,N_9959,N_9723);
nand U10257 (N_10257,N_9674,N_9932);
nor U10258 (N_10258,N_9649,N_9995);
or U10259 (N_10259,N_9812,N_9884);
or U10260 (N_10260,N_9849,N_9853);
xor U10261 (N_10261,N_9871,N_9626);
nand U10262 (N_10262,N_9642,N_9652);
and U10263 (N_10263,N_9828,N_9695);
and U10264 (N_10264,N_9855,N_9784);
and U10265 (N_10265,N_9687,N_9603);
xor U10266 (N_10266,N_9957,N_9974);
nor U10267 (N_10267,N_9968,N_9975);
and U10268 (N_10268,N_9640,N_9896);
xor U10269 (N_10269,N_9921,N_9726);
nor U10270 (N_10270,N_9926,N_9670);
xor U10271 (N_10271,N_9724,N_9836);
nor U10272 (N_10272,N_9639,N_9831);
and U10273 (N_10273,N_9838,N_9947);
or U10274 (N_10274,N_9889,N_9851);
and U10275 (N_10275,N_9663,N_9928);
nor U10276 (N_10276,N_9966,N_9740);
nor U10277 (N_10277,N_9917,N_9720);
xnor U10278 (N_10278,N_9706,N_9700);
or U10279 (N_10279,N_9826,N_9786);
nor U10280 (N_10280,N_9990,N_9972);
or U10281 (N_10281,N_9628,N_9974);
and U10282 (N_10282,N_9777,N_9816);
xor U10283 (N_10283,N_9676,N_9925);
nor U10284 (N_10284,N_9941,N_9636);
nand U10285 (N_10285,N_9706,N_9936);
nor U10286 (N_10286,N_9622,N_9962);
nand U10287 (N_10287,N_9741,N_9665);
and U10288 (N_10288,N_9606,N_9791);
nand U10289 (N_10289,N_9843,N_9922);
nand U10290 (N_10290,N_9976,N_9767);
nor U10291 (N_10291,N_9667,N_9734);
or U10292 (N_10292,N_9765,N_9729);
nor U10293 (N_10293,N_9938,N_9703);
nand U10294 (N_10294,N_9868,N_9620);
nand U10295 (N_10295,N_9857,N_9636);
nor U10296 (N_10296,N_9648,N_9796);
nor U10297 (N_10297,N_9778,N_9972);
and U10298 (N_10298,N_9738,N_9952);
nor U10299 (N_10299,N_9930,N_9762);
xor U10300 (N_10300,N_9729,N_9897);
and U10301 (N_10301,N_9707,N_9857);
or U10302 (N_10302,N_9845,N_9981);
and U10303 (N_10303,N_9624,N_9766);
nand U10304 (N_10304,N_9950,N_9685);
xnor U10305 (N_10305,N_9947,N_9700);
nor U10306 (N_10306,N_9955,N_9744);
xnor U10307 (N_10307,N_9961,N_9699);
nand U10308 (N_10308,N_9734,N_9979);
nor U10309 (N_10309,N_9993,N_9726);
nand U10310 (N_10310,N_9692,N_9908);
nand U10311 (N_10311,N_9966,N_9956);
xnor U10312 (N_10312,N_9616,N_9701);
or U10313 (N_10313,N_9794,N_9708);
or U10314 (N_10314,N_9779,N_9697);
nand U10315 (N_10315,N_9723,N_9940);
nand U10316 (N_10316,N_9814,N_9988);
xnor U10317 (N_10317,N_9808,N_9834);
and U10318 (N_10318,N_9768,N_9846);
nor U10319 (N_10319,N_9977,N_9831);
nor U10320 (N_10320,N_9932,N_9816);
nor U10321 (N_10321,N_9952,N_9906);
nor U10322 (N_10322,N_9955,N_9788);
nand U10323 (N_10323,N_9982,N_9915);
and U10324 (N_10324,N_9793,N_9702);
nand U10325 (N_10325,N_9690,N_9619);
nand U10326 (N_10326,N_9887,N_9865);
nand U10327 (N_10327,N_9611,N_9960);
nand U10328 (N_10328,N_9761,N_9635);
or U10329 (N_10329,N_9751,N_9923);
nand U10330 (N_10330,N_9737,N_9910);
nand U10331 (N_10331,N_9887,N_9775);
xnor U10332 (N_10332,N_9641,N_9695);
and U10333 (N_10333,N_9629,N_9687);
xnor U10334 (N_10334,N_9964,N_9826);
or U10335 (N_10335,N_9697,N_9743);
xnor U10336 (N_10336,N_9892,N_9736);
nand U10337 (N_10337,N_9688,N_9948);
and U10338 (N_10338,N_9631,N_9622);
or U10339 (N_10339,N_9951,N_9635);
or U10340 (N_10340,N_9627,N_9652);
nand U10341 (N_10341,N_9722,N_9923);
and U10342 (N_10342,N_9715,N_9606);
nor U10343 (N_10343,N_9859,N_9623);
nor U10344 (N_10344,N_9749,N_9687);
or U10345 (N_10345,N_9981,N_9840);
and U10346 (N_10346,N_9687,N_9692);
nand U10347 (N_10347,N_9997,N_9965);
and U10348 (N_10348,N_9973,N_9813);
nand U10349 (N_10349,N_9951,N_9714);
nand U10350 (N_10350,N_9892,N_9751);
xor U10351 (N_10351,N_9985,N_9958);
nand U10352 (N_10352,N_9722,N_9793);
or U10353 (N_10353,N_9682,N_9698);
or U10354 (N_10354,N_9828,N_9747);
and U10355 (N_10355,N_9665,N_9672);
and U10356 (N_10356,N_9838,N_9611);
or U10357 (N_10357,N_9678,N_9805);
and U10358 (N_10358,N_9979,N_9668);
xor U10359 (N_10359,N_9879,N_9799);
and U10360 (N_10360,N_9602,N_9964);
and U10361 (N_10361,N_9656,N_9944);
or U10362 (N_10362,N_9683,N_9807);
xor U10363 (N_10363,N_9695,N_9933);
nand U10364 (N_10364,N_9808,N_9974);
nor U10365 (N_10365,N_9603,N_9827);
nand U10366 (N_10366,N_9814,N_9834);
or U10367 (N_10367,N_9776,N_9678);
xor U10368 (N_10368,N_9806,N_9958);
and U10369 (N_10369,N_9812,N_9964);
xor U10370 (N_10370,N_9729,N_9800);
nor U10371 (N_10371,N_9834,N_9860);
xor U10372 (N_10372,N_9935,N_9966);
xor U10373 (N_10373,N_9905,N_9983);
nand U10374 (N_10374,N_9732,N_9919);
xnor U10375 (N_10375,N_9787,N_9732);
and U10376 (N_10376,N_9781,N_9870);
nand U10377 (N_10377,N_9919,N_9693);
and U10378 (N_10378,N_9634,N_9630);
or U10379 (N_10379,N_9872,N_9888);
and U10380 (N_10380,N_9731,N_9975);
and U10381 (N_10381,N_9723,N_9677);
nor U10382 (N_10382,N_9854,N_9988);
or U10383 (N_10383,N_9726,N_9837);
and U10384 (N_10384,N_9728,N_9920);
nand U10385 (N_10385,N_9848,N_9900);
nand U10386 (N_10386,N_9941,N_9878);
and U10387 (N_10387,N_9622,N_9786);
nand U10388 (N_10388,N_9922,N_9735);
nor U10389 (N_10389,N_9659,N_9654);
nor U10390 (N_10390,N_9981,N_9705);
xor U10391 (N_10391,N_9652,N_9939);
nor U10392 (N_10392,N_9701,N_9668);
nor U10393 (N_10393,N_9793,N_9616);
or U10394 (N_10394,N_9684,N_9731);
xnor U10395 (N_10395,N_9808,N_9622);
xor U10396 (N_10396,N_9623,N_9773);
and U10397 (N_10397,N_9639,N_9847);
or U10398 (N_10398,N_9834,N_9997);
and U10399 (N_10399,N_9658,N_9731);
nand U10400 (N_10400,N_10129,N_10122);
nand U10401 (N_10401,N_10281,N_10194);
xor U10402 (N_10402,N_10394,N_10371);
xnor U10403 (N_10403,N_10310,N_10146);
xor U10404 (N_10404,N_10081,N_10313);
or U10405 (N_10405,N_10353,N_10270);
and U10406 (N_10406,N_10193,N_10362);
nor U10407 (N_10407,N_10140,N_10119);
or U10408 (N_10408,N_10118,N_10114);
nand U10409 (N_10409,N_10230,N_10351);
xnor U10410 (N_10410,N_10289,N_10249);
or U10411 (N_10411,N_10167,N_10079);
and U10412 (N_10412,N_10335,N_10328);
nor U10413 (N_10413,N_10205,N_10393);
and U10414 (N_10414,N_10097,N_10091);
xnor U10415 (N_10415,N_10089,N_10387);
xnor U10416 (N_10416,N_10008,N_10386);
nor U10417 (N_10417,N_10106,N_10136);
nor U10418 (N_10418,N_10283,N_10001);
nor U10419 (N_10419,N_10276,N_10088);
nor U10420 (N_10420,N_10164,N_10043);
nand U10421 (N_10421,N_10263,N_10067);
xor U10422 (N_10422,N_10176,N_10040);
nor U10423 (N_10423,N_10217,N_10004);
nor U10424 (N_10424,N_10064,N_10219);
or U10425 (N_10425,N_10050,N_10046);
xor U10426 (N_10426,N_10291,N_10000);
nand U10427 (N_10427,N_10323,N_10253);
nor U10428 (N_10428,N_10201,N_10228);
nor U10429 (N_10429,N_10054,N_10027);
and U10430 (N_10430,N_10261,N_10141);
xnor U10431 (N_10431,N_10121,N_10358);
nand U10432 (N_10432,N_10304,N_10266);
or U10433 (N_10433,N_10095,N_10180);
nand U10434 (N_10434,N_10189,N_10381);
nor U10435 (N_10435,N_10318,N_10350);
nor U10436 (N_10436,N_10195,N_10116);
and U10437 (N_10437,N_10055,N_10252);
xor U10438 (N_10438,N_10307,N_10117);
and U10439 (N_10439,N_10098,N_10020);
nor U10440 (N_10440,N_10213,N_10346);
nand U10441 (N_10441,N_10357,N_10123);
xnor U10442 (N_10442,N_10305,N_10312);
xor U10443 (N_10443,N_10080,N_10231);
and U10444 (N_10444,N_10314,N_10070);
nand U10445 (N_10445,N_10094,N_10356);
nand U10446 (N_10446,N_10085,N_10369);
xor U10447 (N_10447,N_10058,N_10345);
and U10448 (N_10448,N_10245,N_10324);
xor U10449 (N_10449,N_10077,N_10339);
xnor U10450 (N_10450,N_10147,N_10016);
or U10451 (N_10451,N_10221,N_10053);
xnor U10452 (N_10452,N_10032,N_10227);
nor U10453 (N_10453,N_10343,N_10109);
nand U10454 (N_10454,N_10246,N_10216);
and U10455 (N_10455,N_10236,N_10084);
nand U10456 (N_10456,N_10349,N_10330);
nand U10457 (N_10457,N_10374,N_10047);
and U10458 (N_10458,N_10038,N_10185);
or U10459 (N_10459,N_10075,N_10166);
and U10460 (N_10460,N_10366,N_10233);
nor U10461 (N_10461,N_10103,N_10062);
xnor U10462 (N_10462,N_10069,N_10391);
nor U10463 (N_10463,N_10153,N_10274);
nor U10464 (N_10464,N_10292,N_10255);
nor U10465 (N_10465,N_10206,N_10321);
and U10466 (N_10466,N_10316,N_10332);
and U10467 (N_10467,N_10096,N_10066);
nor U10468 (N_10468,N_10203,N_10152);
nand U10469 (N_10469,N_10171,N_10143);
nand U10470 (N_10470,N_10197,N_10113);
nand U10471 (N_10471,N_10010,N_10258);
nor U10472 (N_10472,N_10384,N_10028);
or U10473 (N_10473,N_10259,N_10173);
nor U10474 (N_10474,N_10380,N_10124);
and U10475 (N_10475,N_10375,N_10348);
nor U10476 (N_10476,N_10174,N_10224);
xnor U10477 (N_10477,N_10286,N_10015);
nor U10478 (N_10478,N_10037,N_10225);
xor U10479 (N_10479,N_10115,N_10215);
or U10480 (N_10480,N_10003,N_10244);
or U10481 (N_10481,N_10134,N_10005);
nor U10482 (N_10482,N_10334,N_10368);
xor U10483 (N_10483,N_10250,N_10126);
nor U10484 (N_10484,N_10239,N_10293);
and U10485 (N_10485,N_10187,N_10059);
and U10486 (N_10486,N_10365,N_10264);
or U10487 (N_10487,N_10135,N_10172);
nor U10488 (N_10488,N_10044,N_10102);
nand U10489 (N_10489,N_10306,N_10303);
xnor U10490 (N_10490,N_10284,N_10331);
nand U10491 (N_10491,N_10280,N_10052);
and U10492 (N_10492,N_10247,N_10026);
nor U10493 (N_10493,N_10051,N_10243);
nand U10494 (N_10494,N_10287,N_10290);
xnor U10495 (N_10495,N_10354,N_10169);
xnor U10496 (N_10496,N_10183,N_10395);
nand U10497 (N_10497,N_10065,N_10364);
and U10498 (N_10498,N_10029,N_10031);
nor U10499 (N_10499,N_10042,N_10120);
or U10500 (N_10500,N_10390,N_10017);
xnor U10501 (N_10501,N_10214,N_10056);
and U10502 (N_10502,N_10355,N_10397);
nor U10503 (N_10503,N_10199,N_10177);
and U10504 (N_10504,N_10072,N_10275);
nor U10505 (N_10505,N_10229,N_10154);
nand U10506 (N_10506,N_10130,N_10048);
nor U10507 (N_10507,N_10125,N_10396);
xor U10508 (N_10508,N_10226,N_10019);
or U10509 (N_10509,N_10133,N_10184);
nor U10510 (N_10510,N_10279,N_10188);
and U10511 (N_10511,N_10208,N_10383);
or U10512 (N_10512,N_10212,N_10168);
and U10513 (N_10513,N_10241,N_10338);
or U10514 (N_10514,N_10025,N_10389);
nand U10515 (N_10515,N_10398,N_10099);
nand U10516 (N_10516,N_10112,N_10342);
nor U10517 (N_10517,N_10254,N_10399);
xnor U10518 (N_10518,N_10311,N_10327);
or U10519 (N_10519,N_10308,N_10359);
and U10520 (N_10520,N_10156,N_10041);
xor U10521 (N_10521,N_10378,N_10127);
xnor U10522 (N_10522,N_10178,N_10341);
nand U10523 (N_10523,N_10108,N_10083);
nor U10524 (N_10524,N_10296,N_10373);
and U10525 (N_10525,N_10267,N_10014);
nand U10526 (N_10526,N_10009,N_10372);
or U10527 (N_10527,N_10149,N_10104);
or U10528 (N_10528,N_10300,N_10209);
or U10529 (N_10529,N_10260,N_10222);
xnor U10530 (N_10530,N_10376,N_10186);
and U10531 (N_10531,N_10068,N_10090);
and U10532 (N_10532,N_10060,N_10036);
xor U10533 (N_10533,N_10392,N_10063);
and U10534 (N_10534,N_10200,N_10298);
nor U10535 (N_10535,N_10271,N_10006);
nand U10536 (N_10536,N_10142,N_10082);
xor U10537 (N_10537,N_10137,N_10329);
nor U10538 (N_10538,N_10191,N_10190);
nand U10539 (N_10539,N_10370,N_10076);
nor U10540 (N_10540,N_10297,N_10223);
and U10541 (N_10541,N_10234,N_10179);
nor U10542 (N_10542,N_10377,N_10204);
nor U10543 (N_10543,N_10299,N_10333);
or U10544 (N_10544,N_10272,N_10071);
or U10545 (N_10545,N_10155,N_10278);
or U10546 (N_10546,N_10110,N_10035);
or U10547 (N_10547,N_10160,N_10128);
and U10548 (N_10548,N_10277,N_10024);
and U10549 (N_10549,N_10367,N_10023);
nand U10550 (N_10550,N_10061,N_10073);
nor U10551 (N_10551,N_10101,N_10211);
or U10552 (N_10552,N_10158,N_10295);
xor U10553 (N_10553,N_10319,N_10320);
and U10554 (N_10554,N_10011,N_10039);
nand U10555 (N_10555,N_10139,N_10257);
and U10556 (N_10556,N_10256,N_10078);
and U10557 (N_10557,N_10002,N_10340);
xor U10558 (N_10558,N_10049,N_10165);
or U10559 (N_10559,N_10034,N_10202);
xnor U10560 (N_10560,N_10317,N_10181);
or U10561 (N_10561,N_10132,N_10326);
or U10562 (N_10562,N_10198,N_10302);
nor U10563 (N_10563,N_10175,N_10162);
xor U10564 (N_10564,N_10057,N_10007);
and U10565 (N_10565,N_10045,N_10022);
xnor U10566 (N_10566,N_10033,N_10360);
xnor U10567 (N_10567,N_10074,N_10105);
nor U10568 (N_10568,N_10242,N_10379);
and U10569 (N_10569,N_10220,N_10170);
xor U10570 (N_10570,N_10268,N_10150);
and U10571 (N_10571,N_10107,N_10012);
nor U10572 (N_10572,N_10218,N_10361);
nand U10573 (N_10573,N_10159,N_10315);
nor U10574 (N_10574,N_10235,N_10251);
xnor U10575 (N_10575,N_10265,N_10294);
and U10576 (N_10576,N_10196,N_10388);
xor U10577 (N_10577,N_10269,N_10240);
or U10578 (N_10578,N_10111,N_10282);
and U10579 (N_10579,N_10144,N_10148);
or U10580 (N_10580,N_10325,N_10163);
and U10581 (N_10581,N_10382,N_10092);
and U10582 (N_10582,N_10309,N_10322);
and U10583 (N_10583,N_10021,N_10363);
nand U10584 (N_10584,N_10131,N_10138);
xor U10585 (N_10585,N_10288,N_10157);
nor U10586 (N_10586,N_10238,N_10161);
nor U10587 (N_10587,N_10248,N_10262);
and U10588 (N_10588,N_10273,N_10100);
nand U10589 (N_10589,N_10151,N_10086);
or U10590 (N_10590,N_10087,N_10336);
nand U10591 (N_10591,N_10192,N_10013);
xor U10592 (N_10592,N_10352,N_10030);
xnor U10593 (N_10593,N_10145,N_10285);
nand U10594 (N_10594,N_10207,N_10347);
xnor U10595 (N_10595,N_10210,N_10337);
xnor U10596 (N_10596,N_10018,N_10301);
nand U10597 (N_10597,N_10344,N_10237);
xor U10598 (N_10598,N_10232,N_10093);
xor U10599 (N_10599,N_10182,N_10385);
nor U10600 (N_10600,N_10348,N_10188);
or U10601 (N_10601,N_10149,N_10175);
or U10602 (N_10602,N_10220,N_10202);
or U10603 (N_10603,N_10260,N_10392);
nand U10604 (N_10604,N_10188,N_10077);
xor U10605 (N_10605,N_10015,N_10296);
xnor U10606 (N_10606,N_10299,N_10036);
nor U10607 (N_10607,N_10079,N_10114);
or U10608 (N_10608,N_10363,N_10328);
and U10609 (N_10609,N_10213,N_10221);
or U10610 (N_10610,N_10235,N_10001);
xor U10611 (N_10611,N_10082,N_10209);
nand U10612 (N_10612,N_10227,N_10149);
and U10613 (N_10613,N_10019,N_10120);
nand U10614 (N_10614,N_10259,N_10127);
xor U10615 (N_10615,N_10182,N_10364);
nand U10616 (N_10616,N_10099,N_10330);
nor U10617 (N_10617,N_10201,N_10161);
and U10618 (N_10618,N_10195,N_10363);
nand U10619 (N_10619,N_10083,N_10145);
and U10620 (N_10620,N_10203,N_10289);
nand U10621 (N_10621,N_10075,N_10261);
and U10622 (N_10622,N_10213,N_10198);
and U10623 (N_10623,N_10359,N_10350);
nor U10624 (N_10624,N_10010,N_10276);
and U10625 (N_10625,N_10076,N_10081);
xor U10626 (N_10626,N_10234,N_10337);
and U10627 (N_10627,N_10148,N_10351);
or U10628 (N_10628,N_10230,N_10107);
nor U10629 (N_10629,N_10337,N_10117);
or U10630 (N_10630,N_10225,N_10294);
and U10631 (N_10631,N_10169,N_10206);
xor U10632 (N_10632,N_10119,N_10157);
nor U10633 (N_10633,N_10254,N_10296);
nor U10634 (N_10634,N_10349,N_10306);
nor U10635 (N_10635,N_10157,N_10187);
nor U10636 (N_10636,N_10156,N_10273);
nor U10637 (N_10637,N_10104,N_10077);
or U10638 (N_10638,N_10100,N_10004);
nor U10639 (N_10639,N_10279,N_10014);
nand U10640 (N_10640,N_10178,N_10137);
or U10641 (N_10641,N_10262,N_10178);
or U10642 (N_10642,N_10047,N_10071);
nor U10643 (N_10643,N_10304,N_10015);
and U10644 (N_10644,N_10379,N_10198);
and U10645 (N_10645,N_10225,N_10047);
xnor U10646 (N_10646,N_10094,N_10351);
nand U10647 (N_10647,N_10398,N_10031);
xnor U10648 (N_10648,N_10264,N_10146);
nand U10649 (N_10649,N_10290,N_10393);
nand U10650 (N_10650,N_10078,N_10344);
nand U10651 (N_10651,N_10255,N_10273);
nand U10652 (N_10652,N_10390,N_10377);
nand U10653 (N_10653,N_10239,N_10057);
and U10654 (N_10654,N_10019,N_10220);
nand U10655 (N_10655,N_10024,N_10036);
or U10656 (N_10656,N_10126,N_10301);
nand U10657 (N_10657,N_10051,N_10264);
or U10658 (N_10658,N_10397,N_10064);
nand U10659 (N_10659,N_10217,N_10298);
or U10660 (N_10660,N_10186,N_10084);
nand U10661 (N_10661,N_10167,N_10289);
nor U10662 (N_10662,N_10386,N_10234);
nor U10663 (N_10663,N_10139,N_10327);
xor U10664 (N_10664,N_10279,N_10232);
nand U10665 (N_10665,N_10227,N_10262);
and U10666 (N_10666,N_10232,N_10012);
xor U10667 (N_10667,N_10248,N_10352);
xor U10668 (N_10668,N_10084,N_10388);
and U10669 (N_10669,N_10351,N_10177);
nor U10670 (N_10670,N_10081,N_10226);
nor U10671 (N_10671,N_10310,N_10267);
or U10672 (N_10672,N_10294,N_10030);
xnor U10673 (N_10673,N_10332,N_10216);
and U10674 (N_10674,N_10036,N_10265);
nor U10675 (N_10675,N_10153,N_10287);
and U10676 (N_10676,N_10051,N_10031);
or U10677 (N_10677,N_10021,N_10219);
or U10678 (N_10678,N_10118,N_10191);
nor U10679 (N_10679,N_10325,N_10372);
nand U10680 (N_10680,N_10239,N_10322);
and U10681 (N_10681,N_10301,N_10128);
xor U10682 (N_10682,N_10084,N_10399);
nor U10683 (N_10683,N_10088,N_10049);
xor U10684 (N_10684,N_10372,N_10343);
nand U10685 (N_10685,N_10219,N_10029);
or U10686 (N_10686,N_10329,N_10129);
nand U10687 (N_10687,N_10376,N_10345);
and U10688 (N_10688,N_10254,N_10383);
nor U10689 (N_10689,N_10268,N_10185);
xor U10690 (N_10690,N_10251,N_10132);
and U10691 (N_10691,N_10100,N_10169);
xnor U10692 (N_10692,N_10316,N_10129);
or U10693 (N_10693,N_10375,N_10189);
xor U10694 (N_10694,N_10001,N_10063);
nor U10695 (N_10695,N_10170,N_10057);
and U10696 (N_10696,N_10256,N_10385);
xor U10697 (N_10697,N_10102,N_10209);
or U10698 (N_10698,N_10102,N_10351);
and U10699 (N_10699,N_10069,N_10310);
xor U10700 (N_10700,N_10029,N_10203);
and U10701 (N_10701,N_10278,N_10171);
nand U10702 (N_10702,N_10018,N_10004);
or U10703 (N_10703,N_10388,N_10106);
nand U10704 (N_10704,N_10380,N_10395);
nand U10705 (N_10705,N_10143,N_10049);
xor U10706 (N_10706,N_10216,N_10282);
nor U10707 (N_10707,N_10279,N_10040);
nor U10708 (N_10708,N_10218,N_10114);
or U10709 (N_10709,N_10223,N_10260);
or U10710 (N_10710,N_10068,N_10041);
xnor U10711 (N_10711,N_10379,N_10168);
or U10712 (N_10712,N_10228,N_10277);
nand U10713 (N_10713,N_10218,N_10177);
nand U10714 (N_10714,N_10311,N_10155);
and U10715 (N_10715,N_10334,N_10030);
or U10716 (N_10716,N_10223,N_10208);
and U10717 (N_10717,N_10122,N_10071);
nand U10718 (N_10718,N_10287,N_10145);
or U10719 (N_10719,N_10376,N_10305);
and U10720 (N_10720,N_10111,N_10392);
nand U10721 (N_10721,N_10023,N_10267);
nor U10722 (N_10722,N_10116,N_10339);
nand U10723 (N_10723,N_10336,N_10195);
or U10724 (N_10724,N_10194,N_10050);
nor U10725 (N_10725,N_10105,N_10272);
nand U10726 (N_10726,N_10139,N_10159);
and U10727 (N_10727,N_10367,N_10146);
xor U10728 (N_10728,N_10079,N_10391);
xor U10729 (N_10729,N_10092,N_10054);
nand U10730 (N_10730,N_10163,N_10094);
xnor U10731 (N_10731,N_10022,N_10181);
xor U10732 (N_10732,N_10064,N_10213);
nand U10733 (N_10733,N_10232,N_10386);
xor U10734 (N_10734,N_10020,N_10277);
or U10735 (N_10735,N_10275,N_10237);
xnor U10736 (N_10736,N_10160,N_10381);
and U10737 (N_10737,N_10109,N_10263);
xnor U10738 (N_10738,N_10149,N_10116);
and U10739 (N_10739,N_10269,N_10058);
xnor U10740 (N_10740,N_10325,N_10327);
or U10741 (N_10741,N_10220,N_10328);
nor U10742 (N_10742,N_10055,N_10052);
and U10743 (N_10743,N_10168,N_10293);
and U10744 (N_10744,N_10226,N_10321);
and U10745 (N_10745,N_10030,N_10131);
or U10746 (N_10746,N_10059,N_10365);
nand U10747 (N_10747,N_10172,N_10283);
nor U10748 (N_10748,N_10148,N_10119);
and U10749 (N_10749,N_10234,N_10091);
or U10750 (N_10750,N_10101,N_10138);
and U10751 (N_10751,N_10060,N_10184);
nand U10752 (N_10752,N_10116,N_10260);
and U10753 (N_10753,N_10000,N_10022);
and U10754 (N_10754,N_10020,N_10199);
nand U10755 (N_10755,N_10027,N_10070);
nand U10756 (N_10756,N_10130,N_10344);
xor U10757 (N_10757,N_10084,N_10148);
nand U10758 (N_10758,N_10366,N_10364);
and U10759 (N_10759,N_10323,N_10220);
nor U10760 (N_10760,N_10380,N_10043);
nor U10761 (N_10761,N_10209,N_10151);
nand U10762 (N_10762,N_10003,N_10288);
nor U10763 (N_10763,N_10250,N_10317);
nand U10764 (N_10764,N_10213,N_10195);
and U10765 (N_10765,N_10386,N_10026);
xnor U10766 (N_10766,N_10072,N_10392);
xor U10767 (N_10767,N_10107,N_10397);
xnor U10768 (N_10768,N_10289,N_10038);
nor U10769 (N_10769,N_10162,N_10278);
nor U10770 (N_10770,N_10270,N_10002);
nand U10771 (N_10771,N_10136,N_10352);
xor U10772 (N_10772,N_10275,N_10043);
or U10773 (N_10773,N_10205,N_10203);
or U10774 (N_10774,N_10063,N_10105);
nor U10775 (N_10775,N_10340,N_10086);
xnor U10776 (N_10776,N_10135,N_10136);
xnor U10777 (N_10777,N_10196,N_10108);
and U10778 (N_10778,N_10026,N_10205);
or U10779 (N_10779,N_10380,N_10282);
or U10780 (N_10780,N_10086,N_10017);
nor U10781 (N_10781,N_10291,N_10194);
xnor U10782 (N_10782,N_10026,N_10089);
nor U10783 (N_10783,N_10214,N_10080);
nor U10784 (N_10784,N_10149,N_10024);
xor U10785 (N_10785,N_10292,N_10336);
nand U10786 (N_10786,N_10279,N_10129);
or U10787 (N_10787,N_10302,N_10290);
or U10788 (N_10788,N_10307,N_10124);
nor U10789 (N_10789,N_10019,N_10298);
nor U10790 (N_10790,N_10091,N_10133);
or U10791 (N_10791,N_10248,N_10043);
nor U10792 (N_10792,N_10012,N_10236);
xnor U10793 (N_10793,N_10208,N_10355);
nor U10794 (N_10794,N_10358,N_10015);
or U10795 (N_10795,N_10295,N_10355);
nand U10796 (N_10796,N_10008,N_10045);
and U10797 (N_10797,N_10099,N_10311);
nor U10798 (N_10798,N_10227,N_10228);
nand U10799 (N_10799,N_10070,N_10244);
or U10800 (N_10800,N_10453,N_10509);
or U10801 (N_10801,N_10448,N_10671);
xnor U10802 (N_10802,N_10720,N_10794);
nand U10803 (N_10803,N_10537,N_10524);
nand U10804 (N_10804,N_10480,N_10549);
xnor U10805 (N_10805,N_10722,N_10455);
nor U10806 (N_10806,N_10401,N_10791);
xnor U10807 (N_10807,N_10500,N_10797);
nand U10808 (N_10808,N_10484,N_10553);
or U10809 (N_10809,N_10701,N_10409);
and U10810 (N_10810,N_10573,N_10600);
nor U10811 (N_10811,N_10675,N_10646);
xor U10812 (N_10812,N_10420,N_10408);
xnor U10813 (N_10813,N_10633,N_10558);
xnor U10814 (N_10814,N_10707,N_10717);
nor U10815 (N_10815,N_10548,N_10451);
nand U10816 (N_10816,N_10793,N_10641);
and U10817 (N_10817,N_10556,N_10590);
nand U10818 (N_10818,N_10660,N_10735);
nand U10819 (N_10819,N_10623,N_10501);
nor U10820 (N_10820,N_10427,N_10767);
and U10821 (N_10821,N_10688,N_10596);
and U10822 (N_10822,N_10760,N_10606);
xor U10823 (N_10823,N_10419,N_10499);
nor U10824 (N_10824,N_10670,N_10697);
and U10825 (N_10825,N_10621,N_10622);
xnor U10826 (N_10826,N_10446,N_10561);
nor U10827 (N_10827,N_10785,N_10547);
or U10828 (N_10828,N_10658,N_10650);
xnor U10829 (N_10829,N_10464,N_10730);
xnor U10830 (N_10830,N_10435,N_10654);
xnor U10831 (N_10831,N_10610,N_10710);
nor U10832 (N_10832,N_10643,N_10598);
and U10833 (N_10833,N_10530,N_10749);
nand U10834 (N_10834,N_10443,N_10544);
nor U10835 (N_10835,N_10663,N_10692);
or U10836 (N_10836,N_10614,N_10611);
xor U10837 (N_10837,N_10784,N_10652);
or U10838 (N_10838,N_10655,N_10636);
xnor U10839 (N_10839,N_10452,N_10763);
nor U10840 (N_10840,N_10478,N_10515);
and U10841 (N_10841,N_10525,N_10560);
and U10842 (N_10842,N_10442,N_10753);
xor U10843 (N_10843,N_10689,N_10559);
or U10844 (N_10844,N_10513,N_10545);
nand U10845 (N_10845,N_10586,N_10750);
xnor U10846 (N_10846,N_10582,N_10583);
xor U10847 (N_10847,N_10539,N_10726);
or U10848 (N_10848,N_10532,N_10465);
nand U10849 (N_10849,N_10472,N_10694);
and U10850 (N_10850,N_10425,N_10746);
nor U10851 (N_10851,N_10713,N_10775);
nand U10852 (N_10852,N_10687,N_10494);
or U10853 (N_10853,N_10741,N_10661);
nor U10854 (N_10854,N_10593,N_10639);
xnor U10855 (N_10855,N_10533,N_10731);
and U10856 (N_10856,N_10521,N_10569);
or U10857 (N_10857,N_10647,N_10475);
or U10858 (N_10858,N_10754,N_10468);
nor U10859 (N_10859,N_10462,N_10624);
and U10860 (N_10860,N_10402,N_10570);
and U10861 (N_10861,N_10507,N_10644);
nand U10862 (N_10862,N_10686,N_10765);
xor U10863 (N_10863,N_10732,N_10492);
nor U10864 (N_10864,N_10781,N_10564);
and U10865 (N_10865,N_10659,N_10479);
nor U10866 (N_10866,N_10519,N_10777);
xnor U10867 (N_10867,N_10445,N_10461);
nand U10868 (N_10868,N_10540,N_10597);
nand U10869 (N_10869,N_10699,N_10782);
nor U10870 (N_10870,N_10703,N_10764);
nand U10871 (N_10871,N_10673,N_10463);
nor U10872 (N_10872,N_10729,N_10736);
nand U10873 (N_10873,N_10637,N_10577);
xnor U10874 (N_10874,N_10504,N_10578);
xor U10875 (N_10875,N_10742,N_10563);
or U10876 (N_10876,N_10587,N_10431);
xnor U10877 (N_10877,N_10551,N_10727);
and U10878 (N_10878,N_10604,N_10798);
xor U10879 (N_10879,N_10470,N_10592);
or U10880 (N_10880,N_10526,N_10555);
or U10881 (N_10881,N_10625,N_10721);
nand U10882 (N_10882,N_10576,N_10456);
xnor U10883 (N_10883,N_10469,N_10748);
or U10884 (N_10884,N_10580,N_10759);
and U10885 (N_10885,N_10541,N_10432);
or U10886 (N_10886,N_10552,N_10679);
nand U10887 (N_10887,N_10450,N_10487);
xor U10888 (N_10888,N_10602,N_10628);
or U10889 (N_10889,N_10744,N_10458);
or U10890 (N_10890,N_10787,N_10779);
nor U10891 (N_10891,N_10795,N_10529);
or U10892 (N_10892,N_10438,N_10546);
xor U10893 (N_10893,N_10407,N_10796);
nand U10894 (N_10894,N_10506,N_10664);
nand U10895 (N_10895,N_10538,N_10690);
xor U10896 (N_10896,N_10543,N_10416);
xor U10897 (N_10897,N_10649,N_10698);
nand U10898 (N_10898,N_10474,N_10486);
nand U10899 (N_10899,N_10756,N_10629);
nand U10900 (N_10900,N_10711,N_10572);
and U10901 (N_10901,N_10485,N_10734);
and U10902 (N_10902,N_10612,N_10620);
nor U10903 (N_10903,N_10723,N_10437);
nand U10904 (N_10904,N_10567,N_10762);
xnor U10905 (N_10905,N_10695,N_10712);
nand U10906 (N_10906,N_10706,N_10773);
xor U10907 (N_10907,N_10467,N_10557);
nand U10908 (N_10908,N_10424,N_10733);
xnor U10909 (N_10909,N_10516,N_10790);
or U10910 (N_10910,N_10489,N_10481);
nand U10911 (N_10911,N_10617,N_10768);
xor U10912 (N_10912,N_10584,N_10511);
nand U10913 (N_10913,N_10657,N_10769);
nor U10914 (N_10914,N_10404,N_10403);
nand U10915 (N_10915,N_10743,N_10589);
xnor U10916 (N_10916,N_10493,N_10682);
nand U10917 (N_10917,N_10594,N_10728);
nor U10918 (N_10918,N_10497,N_10498);
nor U10919 (N_10919,N_10651,N_10466);
and U10920 (N_10920,N_10770,N_10508);
and U10921 (N_10921,N_10766,N_10460);
xor U10922 (N_10922,N_10786,N_10550);
xnor U10923 (N_10923,N_10719,N_10585);
nand U10924 (N_10924,N_10792,N_10421);
xor U10925 (N_10925,N_10490,N_10608);
or U10926 (N_10926,N_10599,N_10491);
and U10927 (N_10927,N_10591,N_10778);
xnor U10928 (N_10928,N_10406,N_10662);
nor U10929 (N_10929,N_10751,N_10656);
xnor U10930 (N_10930,N_10588,N_10422);
and U10931 (N_10931,N_10457,N_10772);
xnor U10932 (N_10932,N_10528,N_10510);
and U10933 (N_10933,N_10426,N_10440);
nand U10934 (N_10934,N_10627,N_10642);
nand U10935 (N_10935,N_10441,N_10454);
nand U10936 (N_10936,N_10771,N_10618);
or U10937 (N_10937,N_10774,N_10579);
and U10938 (N_10938,N_10680,N_10613);
and U10939 (N_10939,N_10449,N_10428);
nor U10940 (N_10940,N_10444,N_10718);
or U10941 (N_10941,N_10562,N_10747);
xor U10942 (N_10942,N_10634,N_10715);
or U10943 (N_10943,N_10761,N_10648);
and U10944 (N_10944,N_10517,N_10684);
xor U10945 (N_10945,N_10737,N_10674);
nor U10946 (N_10946,N_10410,N_10411);
xnor U10947 (N_10947,N_10414,N_10716);
xor U10948 (N_10948,N_10757,N_10678);
nand U10949 (N_10949,N_10565,N_10638);
nor U10950 (N_10950,N_10789,N_10745);
and U10951 (N_10951,N_10512,N_10568);
nor U10952 (N_10952,N_10483,N_10405);
nand U10953 (N_10953,N_10714,N_10430);
xor U10954 (N_10954,N_10534,N_10640);
or U10955 (N_10955,N_10542,N_10667);
and U10956 (N_10956,N_10601,N_10704);
nor U10957 (N_10957,N_10632,N_10495);
xor U10958 (N_10958,N_10709,N_10434);
or U10959 (N_10959,N_10400,N_10645);
and U10960 (N_10960,N_10724,N_10518);
and U10961 (N_10961,N_10459,N_10799);
or U10962 (N_10962,N_10574,N_10418);
nand U10963 (N_10963,N_10669,N_10700);
and U10964 (N_10964,N_10677,N_10581);
and U10965 (N_10965,N_10554,N_10630);
nor U10966 (N_10966,N_10702,N_10488);
nand U10967 (N_10967,N_10752,N_10739);
nand U10968 (N_10968,N_10609,N_10619);
nor U10969 (N_10969,N_10738,N_10626);
xor U10970 (N_10970,N_10566,N_10776);
nor U10971 (N_10971,N_10417,N_10522);
or U10972 (N_10972,N_10412,N_10740);
and U10973 (N_10973,N_10436,N_10527);
nor U10974 (N_10974,N_10635,N_10605);
nand U10975 (N_10975,N_10503,N_10672);
or U10976 (N_10976,N_10482,N_10755);
xnor U10977 (N_10977,N_10476,N_10631);
xnor U10978 (N_10978,N_10653,N_10447);
nand U10979 (N_10979,N_10691,N_10616);
or U10980 (N_10980,N_10705,N_10607);
or U10981 (N_10981,N_10571,N_10413);
xnor U10982 (N_10982,N_10595,N_10535);
nor U10983 (N_10983,N_10433,N_10725);
nor U10984 (N_10984,N_10676,N_10665);
nor U10985 (N_10985,N_10758,N_10788);
or U10986 (N_10986,N_10685,N_10473);
xnor U10987 (N_10987,N_10496,N_10505);
xnor U10988 (N_10988,N_10615,N_10439);
nor U10989 (N_10989,N_10666,N_10696);
xor U10990 (N_10990,N_10693,N_10523);
xnor U10991 (N_10991,N_10681,N_10708);
nor U10992 (N_10992,N_10471,N_10514);
or U10993 (N_10993,N_10536,N_10415);
nor U10994 (N_10994,N_10502,N_10520);
nor U10995 (N_10995,N_10575,N_10429);
or U10996 (N_10996,N_10683,N_10531);
xnor U10997 (N_10997,N_10668,N_10477);
xnor U10998 (N_10998,N_10780,N_10423);
nand U10999 (N_10999,N_10783,N_10603);
nand U11000 (N_11000,N_10795,N_10527);
and U11001 (N_11001,N_10549,N_10560);
and U11002 (N_11002,N_10551,N_10549);
xor U11003 (N_11003,N_10548,N_10667);
and U11004 (N_11004,N_10661,N_10711);
xor U11005 (N_11005,N_10473,N_10463);
xnor U11006 (N_11006,N_10773,N_10693);
nor U11007 (N_11007,N_10445,N_10681);
and U11008 (N_11008,N_10706,N_10487);
and U11009 (N_11009,N_10733,N_10746);
xor U11010 (N_11010,N_10660,N_10452);
and U11011 (N_11011,N_10655,N_10504);
nor U11012 (N_11012,N_10485,N_10607);
or U11013 (N_11013,N_10777,N_10680);
and U11014 (N_11014,N_10795,N_10426);
nand U11015 (N_11015,N_10749,N_10641);
and U11016 (N_11016,N_10561,N_10694);
nor U11017 (N_11017,N_10655,N_10594);
xor U11018 (N_11018,N_10409,N_10756);
nor U11019 (N_11019,N_10472,N_10641);
or U11020 (N_11020,N_10413,N_10556);
and U11021 (N_11021,N_10539,N_10485);
nor U11022 (N_11022,N_10509,N_10468);
xor U11023 (N_11023,N_10498,N_10667);
or U11024 (N_11024,N_10530,N_10489);
and U11025 (N_11025,N_10773,N_10531);
and U11026 (N_11026,N_10789,N_10589);
xor U11027 (N_11027,N_10748,N_10650);
nor U11028 (N_11028,N_10612,N_10632);
and U11029 (N_11029,N_10756,N_10602);
or U11030 (N_11030,N_10781,N_10603);
xor U11031 (N_11031,N_10708,N_10413);
or U11032 (N_11032,N_10491,N_10515);
or U11033 (N_11033,N_10794,N_10493);
nand U11034 (N_11034,N_10653,N_10725);
and U11035 (N_11035,N_10561,N_10552);
or U11036 (N_11036,N_10676,N_10736);
and U11037 (N_11037,N_10458,N_10782);
or U11038 (N_11038,N_10414,N_10407);
and U11039 (N_11039,N_10603,N_10528);
nor U11040 (N_11040,N_10788,N_10565);
nand U11041 (N_11041,N_10715,N_10550);
xnor U11042 (N_11042,N_10745,N_10547);
xnor U11043 (N_11043,N_10513,N_10665);
nand U11044 (N_11044,N_10783,N_10745);
or U11045 (N_11045,N_10642,N_10496);
xor U11046 (N_11046,N_10480,N_10516);
or U11047 (N_11047,N_10743,N_10533);
xor U11048 (N_11048,N_10619,N_10413);
nand U11049 (N_11049,N_10403,N_10598);
or U11050 (N_11050,N_10481,N_10674);
and U11051 (N_11051,N_10782,N_10582);
xor U11052 (N_11052,N_10653,N_10405);
and U11053 (N_11053,N_10760,N_10610);
xor U11054 (N_11054,N_10603,N_10512);
nor U11055 (N_11055,N_10523,N_10793);
nand U11056 (N_11056,N_10683,N_10749);
and U11057 (N_11057,N_10440,N_10708);
xor U11058 (N_11058,N_10543,N_10438);
and U11059 (N_11059,N_10531,N_10794);
nand U11060 (N_11060,N_10627,N_10653);
and U11061 (N_11061,N_10565,N_10774);
and U11062 (N_11062,N_10526,N_10703);
nand U11063 (N_11063,N_10664,N_10701);
xnor U11064 (N_11064,N_10473,N_10547);
or U11065 (N_11065,N_10549,N_10462);
nor U11066 (N_11066,N_10676,N_10608);
nand U11067 (N_11067,N_10498,N_10489);
nand U11068 (N_11068,N_10453,N_10458);
and U11069 (N_11069,N_10658,N_10619);
or U11070 (N_11070,N_10573,N_10428);
and U11071 (N_11071,N_10415,N_10493);
or U11072 (N_11072,N_10605,N_10575);
or U11073 (N_11073,N_10742,N_10655);
and U11074 (N_11074,N_10790,N_10607);
nor U11075 (N_11075,N_10643,N_10636);
or U11076 (N_11076,N_10404,N_10755);
and U11077 (N_11077,N_10504,N_10560);
nand U11078 (N_11078,N_10568,N_10769);
or U11079 (N_11079,N_10696,N_10754);
nor U11080 (N_11080,N_10477,N_10445);
xnor U11081 (N_11081,N_10794,N_10440);
xnor U11082 (N_11082,N_10786,N_10527);
xor U11083 (N_11083,N_10566,N_10621);
nor U11084 (N_11084,N_10691,N_10710);
nand U11085 (N_11085,N_10507,N_10794);
nand U11086 (N_11086,N_10649,N_10764);
or U11087 (N_11087,N_10614,N_10637);
nand U11088 (N_11088,N_10593,N_10725);
or U11089 (N_11089,N_10510,N_10425);
and U11090 (N_11090,N_10778,N_10516);
xor U11091 (N_11091,N_10436,N_10718);
or U11092 (N_11092,N_10438,N_10555);
nand U11093 (N_11093,N_10655,N_10582);
xor U11094 (N_11094,N_10789,N_10594);
or U11095 (N_11095,N_10706,N_10476);
nor U11096 (N_11096,N_10470,N_10525);
xor U11097 (N_11097,N_10615,N_10515);
xnor U11098 (N_11098,N_10646,N_10486);
or U11099 (N_11099,N_10787,N_10401);
and U11100 (N_11100,N_10602,N_10734);
or U11101 (N_11101,N_10710,N_10491);
and U11102 (N_11102,N_10635,N_10692);
or U11103 (N_11103,N_10739,N_10452);
nand U11104 (N_11104,N_10634,N_10431);
nand U11105 (N_11105,N_10683,N_10442);
nand U11106 (N_11106,N_10671,N_10499);
xor U11107 (N_11107,N_10641,N_10478);
nand U11108 (N_11108,N_10420,N_10452);
nand U11109 (N_11109,N_10531,N_10406);
or U11110 (N_11110,N_10618,N_10464);
and U11111 (N_11111,N_10705,N_10536);
nand U11112 (N_11112,N_10634,N_10519);
or U11113 (N_11113,N_10505,N_10526);
nor U11114 (N_11114,N_10560,N_10466);
xor U11115 (N_11115,N_10481,N_10465);
xnor U11116 (N_11116,N_10536,N_10540);
and U11117 (N_11117,N_10617,N_10752);
nor U11118 (N_11118,N_10662,N_10784);
nand U11119 (N_11119,N_10645,N_10441);
nand U11120 (N_11120,N_10472,N_10748);
and U11121 (N_11121,N_10601,N_10730);
and U11122 (N_11122,N_10587,N_10592);
nand U11123 (N_11123,N_10527,N_10650);
and U11124 (N_11124,N_10715,N_10704);
nand U11125 (N_11125,N_10513,N_10695);
or U11126 (N_11126,N_10505,N_10613);
xnor U11127 (N_11127,N_10681,N_10772);
and U11128 (N_11128,N_10724,N_10741);
nor U11129 (N_11129,N_10483,N_10535);
and U11130 (N_11130,N_10747,N_10426);
xnor U11131 (N_11131,N_10648,N_10533);
or U11132 (N_11132,N_10635,N_10516);
and U11133 (N_11133,N_10494,N_10704);
xor U11134 (N_11134,N_10704,N_10478);
and U11135 (N_11135,N_10609,N_10650);
or U11136 (N_11136,N_10409,N_10713);
nand U11137 (N_11137,N_10539,N_10504);
and U11138 (N_11138,N_10789,N_10570);
nand U11139 (N_11139,N_10737,N_10570);
or U11140 (N_11140,N_10458,N_10735);
nand U11141 (N_11141,N_10628,N_10720);
or U11142 (N_11142,N_10519,N_10534);
nor U11143 (N_11143,N_10721,N_10400);
or U11144 (N_11144,N_10524,N_10789);
xnor U11145 (N_11145,N_10489,N_10663);
xnor U11146 (N_11146,N_10721,N_10594);
nor U11147 (N_11147,N_10401,N_10556);
nand U11148 (N_11148,N_10790,N_10603);
xnor U11149 (N_11149,N_10607,N_10717);
xnor U11150 (N_11150,N_10503,N_10682);
or U11151 (N_11151,N_10479,N_10511);
nand U11152 (N_11152,N_10473,N_10527);
xnor U11153 (N_11153,N_10713,N_10560);
nor U11154 (N_11154,N_10632,N_10607);
or U11155 (N_11155,N_10611,N_10425);
and U11156 (N_11156,N_10696,N_10410);
nand U11157 (N_11157,N_10702,N_10677);
nor U11158 (N_11158,N_10471,N_10509);
and U11159 (N_11159,N_10475,N_10469);
and U11160 (N_11160,N_10748,N_10647);
nor U11161 (N_11161,N_10526,N_10608);
xnor U11162 (N_11162,N_10585,N_10500);
and U11163 (N_11163,N_10701,N_10759);
xnor U11164 (N_11164,N_10485,N_10735);
and U11165 (N_11165,N_10668,N_10450);
or U11166 (N_11166,N_10575,N_10772);
xnor U11167 (N_11167,N_10613,N_10572);
and U11168 (N_11168,N_10421,N_10748);
or U11169 (N_11169,N_10466,N_10636);
nand U11170 (N_11170,N_10465,N_10692);
nor U11171 (N_11171,N_10664,N_10754);
xor U11172 (N_11172,N_10628,N_10773);
xnor U11173 (N_11173,N_10768,N_10540);
and U11174 (N_11174,N_10485,N_10580);
and U11175 (N_11175,N_10595,N_10632);
nand U11176 (N_11176,N_10457,N_10418);
nor U11177 (N_11177,N_10712,N_10638);
nor U11178 (N_11178,N_10527,N_10565);
nand U11179 (N_11179,N_10425,N_10546);
nor U11180 (N_11180,N_10741,N_10677);
and U11181 (N_11181,N_10497,N_10595);
nand U11182 (N_11182,N_10455,N_10414);
nand U11183 (N_11183,N_10536,N_10598);
and U11184 (N_11184,N_10476,N_10727);
nand U11185 (N_11185,N_10757,N_10414);
or U11186 (N_11186,N_10634,N_10630);
xnor U11187 (N_11187,N_10518,N_10573);
and U11188 (N_11188,N_10754,N_10722);
and U11189 (N_11189,N_10473,N_10605);
xor U11190 (N_11190,N_10697,N_10741);
nor U11191 (N_11191,N_10765,N_10487);
xnor U11192 (N_11192,N_10487,N_10403);
or U11193 (N_11193,N_10739,N_10698);
and U11194 (N_11194,N_10513,N_10486);
or U11195 (N_11195,N_10596,N_10464);
nand U11196 (N_11196,N_10662,N_10596);
or U11197 (N_11197,N_10538,N_10728);
xor U11198 (N_11198,N_10422,N_10780);
and U11199 (N_11199,N_10494,N_10757);
and U11200 (N_11200,N_11038,N_10821);
nand U11201 (N_11201,N_10976,N_10956);
and U11202 (N_11202,N_11117,N_10938);
or U11203 (N_11203,N_11030,N_11131);
nand U11204 (N_11204,N_10952,N_10964);
nor U11205 (N_11205,N_11014,N_10828);
or U11206 (N_11206,N_11066,N_11052);
nor U11207 (N_11207,N_11187,N_10838);
nand U11208 (N_11208,N_10989,N_10965);
nor U11209 (N_11209,N_10834,N_10948);
nand U11210 (N_11210,N_11114,N_10904);
or U11211 (N_11211,N_10873,N_11105);
and U11212 (N_11212,N_10829,N_11042);
nand U11213 (N_11213,N_11100,N_11194);
nor U11214 (N_11214,N_10924,N_10806);
and U11215 (N_11215,N_10903,N_11077);
or U11216 (N_11216,N_11084,N_11159);
nand U11217 (N_11217,N_10907,N_11026);
and U11218 (N_11218,N_11181,N_10982);
xor U11219 (N_11219,N_10943,N_10864);
and U11220 (N_11220,N_10919,N_10966);
nor U11221 (N_11221,N_11158,N_11076);
or U11222 (N_11222,N_10843,N_10868);
and U11223 (N_11223,N_10933,N_10851);
nor U11224 (N_11224,N_10879,N_10921);
or U11225 (N_11225,N_10836,N_11070);
xor U11226 (N_11226,N_10897,N_11022);
nor U11227 (N_11227,N_10839,N_11107);
nor U11228 (N_11228,N_11079,N_10803);
nor U11229 (N_11229,N_11065,N_10857);
nand U11230 (N_11230,N_11016,N_10874);
or U11231 (N_11231,N_11185,N_10810);
xnor U11232 (N_11232,N_10960,N_10809);
xnor U11233 (N_11233,N_11031,N_10882);
or U11234 (N_11234,N_10923,N_11049);
xor U11235 (N_11235,N_11018,N_11191);
xnor U11236 (N_11236,N_11075,N_11054);
nor U11237 (N_11237,N_10934,N_11027);
nand U11238 (N_11238,N_10862,N_11029);
or U11239 (N_11239,N_11017,N_11047);
nand U11240 (N_11240,N_11166,N_10899);
xnor U11241 (N_11241,N_11128,N_10962);
nand U11242 (N_11242,N_11103,N_11039);
xnor U11243 (N_11243,N_10972,N_10871);
nand U11244 (N_11244,N_11167,N_10967);
nor U11245 (N_11245,N_11001,N_11086);
xor U11246 (N_11246,N_10953,N_11134);
or U11247 (N_11247,N_11135,N_11125);
and U11248 (N_11248,N_10911,N_11062);
and U11249 (N_11249,N_10979,N_11010);
xnor U11250 (N_11250,N_10931,N_11148);
xor U11251 (N_11251,N_10833,N_10853);
nand U11252 (N_11252,N_11091,N_11182);
xor U11253 (N_11253,N_11126,N_11089);
and U11254 (N_11254,N_10885,N_11093);
nor U11255 (N_11255,N_11146,N_11032);
or U11256 (N_11256,N_11090,N_10996);
and U11257 (N_11257,N_11142,N_11132);
nand U11258 (N_11258,N_11150,N_10813);
xnor U11259 (N_11259,N_11147,N_10975);
and U11260 (N_11260,N_10957,N_10870);
nor U11261 (N_11261,N_10883,N_11102);
and U11262 (N_11262,N_11072,N_11118);
nor U11263 (N_11263,N_11112,N_10917);
xnor U11264 (N_11264,N_10999,N_10890);
and U11265 (N_11265,N_11170,N_11020);
xnor U11266 (N_11266,N_10808,N_10922);
xor U11267 (N_11267,N_11152,N_10855);
nor U11268 (N_11268,N_10822,N_11190);
or U11269 (N_11269,N_10867,N_10861);
nor U11270 (N_11270,N_11129,N_11155);
and U11271 (N_11271,N_11063,N_10825);
nor U11272 (N_11272,N_11183,N_10815);
xnor U11273 (N_11273,N_11083,N_10961);
nand U11274 (N_11274,N_10802,N_11035);
xor U11275 (N_11275,N_10887,N_10978);
nand U11276 (N_11276,N_10936,N_11163);
nand U11277 (N_11277,N_11064,N_11046);
nor U11278 (N_11278,N_10944,N_11099);
nor U11279 (N_11279,N_10908,N_11156);
nand U11280 (N_11280,N_11088,N_10849);
xnor U11281 (N_11281,N_11024,N_10969);
xnor U11282 (N_11282,N_10997,N_10848);
or U11283 (N_11283,N_10814,N_10894);
xnor U11284 (N_11284,N_11050,N_10805);
nand U11285 (N_11285,N_10832,N_11160);
nand U11286 (N_11286,N_11144,N_11055);
xor U11287 (N_11287,N_11085,N_10852);
and U11288 (N_11288,N_11034,N_10998);
nor U11289 (N_11289,N_10820,N_10925);
and U11290 (N_11290,N_11033,N_11108);
nor U11291 (N_11291,N_11074,N_11124);
or U11292 (N_11292,N_10995,N_10929);
xnor U11293 (N_11293,N_10914,N_11188);
xor U11294 (N_11294,N_11165,N_10840);
xnor U11295 (N_11295,N_10905,N_10951);
nor U11296 (N_11296,N_10988,N_10909);
nor U11297 (N_11297,N_10889,N_10983);
xnor U11298 (N_11298,N_10892,N_11019);
nand U11299 (N_11299,N_11157,N_10888);
nor U11300 (N_11300,N_11061,N_11081);
or U11301 (N_11301,N_11176,N_11044);
and U11302 (N_11302,N_11003,N_10986);
nor U11303 (N_11303,N_11168,N_10954);
xnor U11304 (N_11304,N_10918,N_10898);
nand U11305 (N_11305,N_11122,N_11172);
xor U11306 (N_11306,N_10824,N_11116);
and U11307 (N_11307,N_10854,N_11053);
and U11308 (N_11308,N_11040,N_10932);
and U11309 (N_11309,N_11060,N_11013);
nand U11310 (N_11310,N_10875,N_10955);
nand U11311 (N_11311,N_11104,N_11198);
nand U11312 (N_11312,N_10850,N_11000);
nor U11313 (N_11313,N_11197,N_11071);
and U11314 (N_11314,N_11145,N_10980);
or U11315 (N_11315,N_10963,N_11094);
or U11316 (N_11316,N_10949,N_11004);
xnor U11317 (N_11317,N_11025,N_10984);
nand U11318 (N_11318,N_11199,N_10912);
and U11319 (N_11319,N_11123,N_11008);
nand U11320 (N_11320,N_11092,N_11193);
nor U11321 (N_11321,N_11196,N_11012);
xor U11322 (N_11322,N_10878,N_10831);
or U11323 (N_11323,N_11139,N_11056);
xor U11324 (N_11324,N_11111,N_11021);
nand U11325 (N_11325,N_10844,N_10900);
or U11326 (N_11326,N_11069,N_11136);
xor U11327 (N_11327,N_11011,N_11133);
or U11328 (N_11328,N_11164,N_11045);
and U11329 (N_11329,N_10819,N_10994);
xnor U11330 (N_11330,N_11051,N_10895);
and U11331 (N_11331,N_11153,N_11080);
nor U11332 (N_11332,N_10891,N_10947);
xor U11333 (N_11333,N_11140,N_10920);
and U11334 (N_11334,N_10926,N_10880);
xor U11335 (N_11335,N_11121,N_10869);
nand U11336 (N_11336,N_11002,N_11192);
xnor U11337 (N_11337,N_11059,N_10837);
nand U11338 (N_11338,N_10801,N_10884);
nor U11339 (N_11339,N_10915,N_11154);
nor U11340 (N_11340,N_10942,N_11127);
and U11341 (N_11341,N_10872,N_11041);
nand U11342 (N_11342,N_11009,N_11137);
xor U11343 (N_11343,N_11067,N_11007);
nand U11344 (N_11344,N_10927,N_10827);
nor U11345 (N_11345,N_11106,N_11171);
and U11346 (N_11346,N_10811,N_11073);
nand U11347 (N_11347,N_10845,N_10991);
and U11348 (N_11348,N_11101,N_10987);
or U11349 (N_11349,N_11068,N_10807);
nand U11350 (N_11350,N_11037,N_10896);
and U11351 (N_11351,N_11149,N_11043);
nand U11352 (N_11352,N_10817,N_10812);
nand U11353 (N_11353,N_11151,N_10946);
and U11354 (N_11354,N_11161,N_10881);
or U11355 (N_11355,N_10804,N_11096);
or U11356 (N_11356,N_10876,N_11186);
nand U11357 (N_11357,N_10842,N_10886);
and U11358 (N_11358,N_10913,N_11162);
and U11359 (N_11359,N_11098,N_11177);
nand U11360 (N_11360,N_11023,N_11036);
or U11361 (N_11361,N_10859,N_11097);
xnor U11362 (N_11362,N_10826,N_10973);
or U11363 (N_11363,N_11169,N_10937);
nor U11364 (N_11364,N_10863,N_11184);
or U11365 (N_11365,N_11180,N_11005);
xnor U11366 (N_11366,N_10877,N_10835);
xnor U11367 (N_11367,N_11082,N_11173);
xor U11368 (N_11368,N_10858,N_10816);
and U11369 (N_11369,N_10847,N_10939);
nand U11370 (N_11370,N_10901,N_10866);
xor U11371 (N_11371,N_11130,N_10841);
nand U11372 (N_11372,N_10930,N_10935);
nor U11373 (N_11373,N_10941,N_10916);
and U11374 (N_11374,N_11087,N_11028);
xnor U11375 (N_11375,N_10959,N_10990);
and U11376 (N_11376,N_10830,N_10860);
xnor U11377 (N_11377,N_10992,N_10893);
nor U11378 (N_11378,N_10865,N_11110);
nand U11379 (N_11379,N_11109,N_11189);
and U11380 (N_11380,N_10985,N_11078);
nor U11381 (N_11381,N_10971,N_11058);
nor U11382 (N_11382,N_10970,N_10902);
nor U11383 (N_11383,N_11113,N_10818);
nand U11384 (N_11384,N_11143,N_11138);
nor U11385 (N_11385,N_11095,N_11175);
or U11386 (N_11386,N_10823,N_11174);
and U11387 (N_11387,N_10928,N_11195);
nand U11388 (N_11388,N_11178,N_10977);
nand U11389 (N_11389,N_11057,N_10968);
nor U11390 (N_11390,N_11141,N_11006);
or U11391 (N_11391,N_10950,N_10800);
xnor U11392 (N_11392,N_10940,N_11119);
nor U11393 (N_11393,N_10993,N_10906);
xnor U11394 (N_11394,N_11048,N_10958);
nor U11395 (N_11395,N_11179,N_10945);
nor U11396 (N_11396,N_10981,N_10910);
nand U11397 (N_11397,N_10846,N_11115);
nand U11398 (N_11398,N_10974,N_10856);
or U11399 (N_11399,N_11120,N_11015);
or U11400 (N_11400,N_10970,N_10947);
or U11401 (N_11401,N_10844,N_11059);
and U11402 (N_11402,N_11117,N_11111);
xnor U11403 (N_11403,N_10878,N_10874);
or U11404 (N_11404,N_11021,N_10994);
xnor U11405 (N_11405,N_10801,N_11152);
xnor U11406 (N_11406,N_11149,N_10926);
or U11407 (N_11407,N_10825,N_10881);
and U11408 (N_11408,N_10922,N_10980);
nor U11409 (N_11409,N_10865,N_10851);
or U11410 (N_11410,N_11052,N_11107);
xor U11411 (N_11411,N_11000,N_10843);
or U11412 (N_11412,N_10964,N_11012);
and U11413 (N_11413,N_10916,N_10986);
nor U11414 (N_11414,N_11193,N_11041);
and U11415 (N_11415,N_11096,N_11006);
nor U11416 (N_11416,N_11044,N_11100);
nand U11417 (N_11417,N_11088,N_10910);
xnor U11418 (N_11418,N_11194,N_11154);
or U11419 (N_11419,N_11087,N_10819);
nor U11420 (N_11420,N_11163,N_10840);
nor U11421 (N_11421,N_10803,N_10815);
nand U11422 (N_11422,N_10874,N_11036);
or U11423 (N_11423,N_11074,N_11135);
xnor U11424 (N_11424,N_10924,N_10934);
and U11425 (N_11425,N_11142,N_10861);
xnor U11426 (N_11426,N_11166,N_11026);
and U11427 (N_11427,N_11022,N_11028);
nand U11428 (N_11428,N_11033,N_11009);
xnor U11429 (N_11429,N_10830,N_11132);
nand U11430 (N_11430,N_10870,N_10930);
nand U11431 (N_11431,N_11172,N_11121);
nand U11432 (N_11432,N_10924,N_10892);
and U11433 (N_11433,N_11061,N_10859);
xor U11434 (N_11434,N_11185,N_10816);
or U11435 (N_11435,N_11068,N_11057);
xnor U11436 (N_11436,N_11034,N_10901);
xnor U11437 (N_11437,N_11135,N_10849);
nor U11438 (N_11438,N_10982,N_11064);
nand U11439 (N_11439,N_10815,N_10972);
or U11440 (N_11440,N_11093,N_11001);
or U11441 (N_11441,N_10824,N_10941);
and U11442 (N_11442,N_10969,N_10983);
xor U11443 (N_11443,N_11197,N_10952);
nand U11444 (N_11444,N_11095,N_11137);
or U11445 (N_11445,N_10961,N_10977);
and U11446 (N_11446,N_10923,N_11104);
and U11447 (N_11447,N_10971,N_11142);
nor U11448 (N_11448,N_11124,N_11046);
xor U11449 (N_11449,N_10867,N_10879);
nor U11450 (N_11450,N_10891,N_10804);
nor U11451 (N_11451,N_11025,N_10934);
nor U11452 (N_11452,N_11072,N_10985);
nand U11453 (N_11453,N_11072,N_10956);
nor U11454 (N_11454,N_11086,N_11191);
xnor U11455 (N_11455,N_10983,N_10929);
or U11456 (N_11456,N_11110,N_11126);
nor U11457 (N_11457,N_11180,N_10921);
or U11458 (N_11458,N_11079,N_10977);
and U11459 (N_11459,N_11199,N_11098);
and U11460 (N_11460,N_11045,N_11007);
or U11461 (N_11461,N_10862,N_11080);
nor U11462 (N_11462,N_10898,N_10969);
nand U11463 (N_11463,N_11124,N_11192);
or U11464 (N_11464,N_10929,N_10854);
and U11465 (N_11465,N_10963,N_10958);
or U11466 (N_11466,N_10983,N_10976);
or U11467 (N_11467,N_11085,N_11062);
or U11468 (N_11468,N_11100,N_11195);
nand U11469 (N_11469,N_11033,N_10932);
xnor U11470 (N_11470,N_10809,N_11071);
nand U11471 (N_11471,N_10878,N_11187);
nor U11472 (N_11472,N_10964,N_10947);
or U11473 (N_11473,N_10951,N_11070);
nor U11474 (N_11474,N_10997,N_10920);
or U11475 (N_11475,N_10965,N_10848);
nor U11476 (N_11476,N_11031,N_11136);
or U11477 (N_11477,N_11154,N_11042);
nand U11478 (N_11478,N_10997,N_10820);
xor U11479 (N_11479,N_11179,N_11015);
or U11480 (N_11480,N_11179,N_11108);
nor U11481 (N_11481,N_10998,N_10890);
or U11482 (N_11482,N_10985,N_10996);
and U11483 (N_11483,N_11048,N_11076);
and U11484 (N_11484,N_10963,N_11092);
or U11485 (N_11485,N_11088,N_11096);
nor U11486 (N_11486,N_11032,N_10871);
nand U11487 (N_11487,N_11092,N_11144);
and U11488 (N_11488,N_10850,N_10927);
or U11489 (N_11489,N_10968,N_11035);
nor U11490 (N_11490,N_10919,N_11147);
and U11491 (N_11491,N_11067,N_11116);
nand U11492 (N_11492,N_10894,N_11167);
xnor U11493 (N_11493,N_11047,N_10998);
nand U11494 (N_11494,N_11002,N_10984);
or U11495 (N_11495,N_10955,N_11105);
and U11496 (N_11496,N_11013,N_10990);
or U11497 (N_11497,N_11156,N_11036);
nor U11498 (N_11498,N_11130,N_11069);
and U11499 (N_11499,N_10873,N_10863);
and U11500 (N_11500,N_10909,N_11162);
and U11501 (N_11501,N_10911,N_10942);
or U11502 (N_11502,N_10916,N_10926);
and U11503 (N_11503,N_10875,N_10945);
and U11504 (N_11504,N_11195,N_10991);
nor U11505 (N_11505,N_11170,N_10993);
nand U11506 (N_11506,N_11138,N_10921);
xor U11507 (N_11507,N_11044,N_11146);
nor U11508 (N_11508,N_11122,N_10887);
nand U11509 (N_11509,N_10949,N_11181);
xor U11510 (N_11510,N_10900,N_11013);
or U11511 (N_11511,N_10852,N_10905);
or U11512 (N_11512,N_10965,N_11038);
and U11513 (N_11513,N_10925,N_11190);
nand U11514 (N_11514,N_11015,N_11069);
nand U11515 (N_11515,N_10965,N_11157);
nor U11516 (N_11516,N_11014,N_11164);
or U11517 (N_11517,N_11026,N_11097);
xnor U11518 (N_11518,N_10975,N_11002);
and U11519 (N_11519,N_10991,N_10854);
and U11520 (N_11520,N_11133,N_11199);
nand U11521 (N_11521,N_10835,N_10853);
xor U11522 (N_11522,N_10937,N_10908);
nand U11523 (N_11523,N_10837,N_10907);
nor U11524 (N_11524,N_11199,N_10921);
xnor U11525 (N_11525,N_11148,N_11070);
or U11526 (N_11526,N_11027,N_10921);
or U11527 (N_11527,N_10847,N_10952);
and U11528 (N_11528,N_11042,N_10872);
nand U11529 (N_11529,N_10955,N_11003);
or U11530 (N_11530,N_10904,N_10930);
nand U11531 (N_11531,N_11081,N_11044);
nor U11532 (N_11532,N_10960,N_10976);
xnor U11533 (N_11533,N_11066,N_11118);
nand U11534 (N_11534,N_10895,N_10820);
and U11535 (N_11535,N_11009,N_10986);
and U11536 (N_11536,N_11139,N_11194);
nor U11537 (N_11537,N_10958,N_11133);
and U11538 (N_11538,N_10832,N_11067);
nand U11539 (N_11539,N_11001,N_11113);
nand U11540 (N_11540,N_10819,N_11059);
and U11541 (N_11541,N_11093,N_10827);
or U11542 (N_11542,N_11113,N_11084);
xor U11543 (N_11543,N_10893,N_10923);
and U11544 (N_11544,N_10975,N_10850);
or U11545 (N_11545,N_11119,N_11111);
nor U11546 (N_11546,N_11016,N_10867);
nor U11547 (N_11547,N_10892,N_10931);
xnor U11548 (N_11548,N_11026,N_10937);
and U11549 (N_11549,N_11196,N_11153);
and U11550 (N_11550,N_11199,N_10871);
xor U11551 (N_11551,N_11144,N_11110);
nand U11552 (N_11552,N_10932,N_10939);
xnor U11553 (N_11553,N_11054,N_10806);
or U11554 (N_11554,N_11012,N_11047);
xnor U11555 (N_11555,N_10991,N_11112);
nand U11556 (N_11556,N_11019,N_10816);
and U11557 (N_11557,N_11179,N_10809);
nor U11558 (N_11558,N_10935,N_11189);
and U11559 (N_11559,N_10995,N_11071);
and U11560 (N_11560,N_11018,N_11188);
and U11561 (N_11561,N_10962,N_11136);
and U11562 (N_11562,N_11087,N_10887);
nor U11563 (N_11563,N_10969,N_11115);
and U11564 (N_11564,N_10994,N_10843);
and U11565 (N_11565,N_11045,N_11102);
nand U11566 (N_11566,N_10973,N_11120);
nor U11567 (N_11567,N_11047,N_11055);
nand U11568 (N_11568,N_11102,N_11103);
and U11569 (N_11569,N_11142,N_11117);
xor U11570 (N_11570,N_10867,N_11058);
nor U11571 (N_11571,N_11018,N_10952);
nor U11572 (N_11572,N_10958,N_11020);
nor U11573 (N_11573,N_10874,N_11098);
nand U11574 (N_11574,N_11123,N_11109);
nor U11575 (N_11575,N_11066,N_11108);
nor U11576 (N_11576,N_10872,N_11120);
and U11577 (N_11577,N_11168,N_11005);
nand U11578 (N_11578,N_11128,N_11031);
nor U11579 (N_11579,N_11031,N_10850);
or U11580 (N_11580,N_10896,N_10852);
or U11581 (N_11581,N_10976,N_11124);
nand U11582 (N_11582,N_10940,N_10950);
nor U11583 (N_11583,N_10974,N_10857);
nand U11584 (N_11584,N_11170,N_10851);
nand U11585 (N_11585,N_11114,N_10976);
or U11586 (N_11586,N_11100,N_10957);
and U11587 (N_11587,N_11134,N_10852);
xnor U11588 (N_11588,N_11123,N_10948);
nand U11589 (N_11589,N_11098,N_10994);
nand U11590 (N_11590,N_11053,N_11164);
and U11591 (N_11591,N_10859,N_10999);
and U11592 (N_11592,N_11185,N_10889);
xnor U11593 (N_11593,N_10833,N_10923);
nor U11594 (N_11594,N_10990,N_10961);
and U11595 (N_11595,N_11118,N_10958);
xnor U11596 (N_11596,N_11048,N_11113);
and U11597 (N_11597,N_10821,N_11067);
or U11598 (N_11598,N_10839,N_10928);
nor U11599 (N_11599,N_11081,N_10897);
xnor U11600 (N_11600,N_11255,N_11291);
xnor U11601 (N_11601,N_11273,N_11307);
nand U11602 (N_11602,N_11427,N_11577);
and U11603 (N_11603,N_11271,N_11405);
and U11604 (N_11604,N_11289,N_11333);
or U11605 (N_11605,N_11299,N_11527);
xnor U11606 (N_11606,N_11435,N_11399);
or U11607 (N_11607,N_11268,N_11410);
nor U11608 (N_11608,N_11279,N_11442);
nor U11609 (N_11609,N_11500,N_11473);
xor U11610 (N_11610,N_11301,N_11499);
and U11611 (N_11611,N_11436,N_11323);
and U11612 (N_11612,N_11402,N_11548);
nand U11613 (N_11613,N_11597,N_11367);
and U11614 (N_11614,N_11453,N_11201);
and U11615 (N_11615,N_11550,N_11566);
nand U11616 (N_11616,N_11554,N_11357);
nand U11617 (N_11617,N_11464,N_11318);
and U11618 (N_11618,N_11495,N_11214);
nor U11619 (N_11619,N_11474,N_11245);
or U11620 (N_11620,N_11277,N_11428);
nand U11621 (N_11621,N_11522,N_11362);
xor U11622 (N_11622,N_11272,N_11552);
nor U11623 (N_11623,N_11241,N_11356);
and U11624 (N_11624,N_11283,N_11525);
or U11625 (N_11625,N_11497,N_11248);
or U11626 (N_11626,N_11538,N_11328);
xnor U11627 (N_11627,N_11439,N_11267);
and U11628 (N_11628,N_11515,N_11544);
nand U11629 (N_11629,N_11297,N_11456);
or U11630 (N_11630,N_11386,N_11243);
nand U11631 (N_11631,N_11276,N_11282);
nand U11632 (N_11632,N_11385,N_11430);
xnor U11633 (N_11633,N_11454,N_11234);
nor U11634 (N_11634,N_11338,N_11535);
nand U11635 (N_11635,N_11217,N_11302);
and U11636 (N_11636,N_11284,N_11560);
nor U11637 (N_11637,N_11270,N_11429);
xnor U11638 (N_11638,N_11211,N_11303);
or U11639 (N_11639,N_11343,N_11533);
xor U11640 (N_11640,N_11233,N_11591);
xor U11641 (N_11641,N_11219,N_11387);
nor U11642 (N_11642,N_11596,N_11363);
and U11643 (N_11643,N_11457,N_11433);
or U11644 (N_11644,N_11575,N_11551);
nand U11645 (N_11645,N_11540,N_11599);
nor U11646 (N_11646,N_11471,N_11496);
or U11647 (N_11647,N_11524,N_11588);
nor U11648 (N_11648,N_11346,N_11585);
xnor U11649 (N_11649,N_11246,N_11371);
nand U11650 (N_11650,N_11407,N_11230);
and U11651 (N_11651,N_11300,N_11528);
and U11652 (N_11652,N_11375,N_11229);
nand U11653 (N_11653,N_11257,N_11409);
nand U11654 (N_11654,N_11223,N_11448);
xnor U11655 (N_11655,N_11361,N_11565);
nor U11656 (N_11656,N_11536,N_11462);
and U11657 (N_11657,N_11506,N_11364);
or U11658 (N_11658,N_11531,N_11526);
nor U11659 (N_11659,N_11422,N_11411);
or U11660 (N_11660,N_11290,N_11529);
and U11661 (N_11661,N_11351,N_11319);
nand U11662 (N_11662,N_11514,N_11379);
xor U11663 (N_11663,N_11341,N_11242);
or U11664 (N_11664,N_11553,N_11488);
nand U11665 (N_11665,N_11563,N_11532);
or U11666 (N_11666,N_11394,N_11306);
xnor U11667 (N_11667,N_11355,N_11417);
nor U11668 (N_11668,N_11449,N_11452);
xor U11669 (N_11669,N_11239,N_11415);
or U11670 (N_11670,N_11523,N_11256);
nand U11671 (N_11671,N_11482,N_11567);
nor U11672 (N_11672,N_11310,N_11240);
nor U11673 (N_11673,N_11459,N_11325);
and U11674 (N_11674,N_11383,N_11580);
and U11675 (N_11675,N_11269,N_11557);
or U11676 (N_11676,N_11477,N_11202);
or U11677 (N_11677,N_11468,N_11534);
xor U11678 (N_11678,N_11340,N_11424);
and U11679 (N_11679,N_11339,N_11398);
nand U11680 (N_11680,N_11481,N_11320);
or U11681 (N_11681,N_11460,N_11207);
xnor U11682 (N_11682,N_11562,N_11546);
nand U11683 (N_11683,N_11370,N_11589);
xor U11684 (N_11684,N_11480,N_11384);
nor U11685 (N_11685,N_11440,N_11359);
or U11686 (N_11686,N_11358,N_11388);
nand U11687 (N_11687,N_11516,N_11479);
or U11688 (N_11688,N_11518,N_11487);
nand U11689 (N_11689,N_11304,N_11380);
xnor U11690 (N_11690,N_11426,N_11425);
or U11691 (N_11691,N_11444,N_11331);
or U11692 (N_11692,N_11502,N_11296);
xnor U11693 (N_11693,N_11253,N_11220);
or U11694 (N_11694,N_11238,N_11483);
xor U11695 (N_11695,N_11542,N_11366);
nor U11696 (N_11696,N_11382,N_11437);
and U11697 (N_11697,N_11218,N_11315);
nor U11698 (N_11698,N_11461,N_11344);
and U11699 (N_11699,N_11579,N_11450);
xnor U11700 (N_11700,N_11587,N_11469);
nor U11701 (N_11701,N_11432,N_11505);
nor U11702 (N_11702,N_11247,N_11521);
nand U11703 (N_11703,N_11491,N_11251);
or U11704 (N_11704,N_11265,N_11445);
nor U11705 (N_11705,N_11235,N_11305);
xor U11706 (N_11706,N_11329,N_11369);
or U11707 (N_11707,N_11206,N_11221);
and U11708 (N_11708,N_11330,N_11517);
or U11709 (N_11709,N_11332,N_11421);
nor U11710 (N_11710,N_11391,N_11520);
nand U11711 (N_11711,N_11224,N_11262);
nor U11712 (N_11712,N_11286,N_11317);
or U11713 (N_11713,N_11475,N_11213);
nor U11714 (N_11714,N_11594,N_11200);
xnor U11715 (N_11715,N_11236,N_11212);
nor U11716 (N_11716,N_11418,N_11438);
or U11717 (N_11717,N_11208,N_11593);
nand U11718 (N_11718,N_11490,N_11549);
and U11719 (N_11719,N_11494,N_11598);
nand U11720 (N_11720,N_11447,N_11595);
xnor U11721 (N_11721,N_11259,N_11390);
or U11722 (N_11722,N_11498,N_11507);
and U11723 (N_11723,N_11582,N_11412);
xor U11724 (N_11724,N_11395,N_11294);
nand U11725 (N_11725,N_11569,N_11443);
xnor U11726 (N_11726,N_11466,N_11396);
nor U11727 (N_11727,N_11455,N_11232);
nor U11728 (N_11728,N_11572,N_11458);
nor U11729 (N_11729,N_11227,N_11210);
or U11730 (N_11730,N_11295,N_11237);
xnor U11731 (N_11731,N_11345,N_11376);
nor U11732 (N_11732,N_11215,N_11352);
and U11733 (N_11733,N_11349,N_11209);
nand U11734 (N_11734,N_11510,N_11222);
nand U11735 (N_11735,N_11354,N_11583);
or U11736 (N_11736,N_11508,N_11258);
nand U11737 (N_11737,N_11342,N_11278);
xnor U11738 (N_11738,N_11413,N_11400);
nand U11739 (N_11739,N_11465,N_11408);
or U11740 (N_11740,N_11463,N_11261);
nand U11741 (N_11741,N_11275,N_11492);
xnor U11742 (N_11742,N_11336,N_11397);
nand U11743 (N_11743,N_11308,N_11568);
nor U11744 (N_11744,N_11592,N_11360);
or U11745 (N_11745,N_11225,N_11280);
nor U11746 (N_11746,N_11470,N_11511);
or U11747 (N_11747,N_11543,N_11434);
xnor U11748 (N_11748,N_11314,N_11558);
or U11749 (N_11749,N_11441,N_11353);
xor U11750 (N_11750,N_11334,N_11377);
or U11751 (N_11751,N_11287,N_11423);
and U11752 (N_11752,N_11274,N_11584);
or U11753 (N_11753,N_11509,N_11249);
nand U11754 (N_11754,N_11578,N_11312);
nor U11755 (N_11755,N_11467,N_11493);
nor U11756 (N_11756,N_11264,N_11292);
or U11757 (N_11757,N_11327,N_11266);
or U11758 (N_11758,N_11513,N_11539);
or U11759 (N_11759,N_11216,N_11226);
or U11760 (N_11760,N_11335,N_11205);
nand U11761 (N_11761,N_11406,N_11451);
xor U11762 (N_11762,N_11501,N_11512);
nand U11763 (N_11763,N_11446,N_11486);
nor U11764 (N_11764,N_11348,N_11313);
or U11765 (N_11765,N_11285,N_11556);
nand U11766 (N_11766,N_11368,N_11321);
nor U11767 (N_11767,N_11260,N_11392);
and U11768 (N_11768,N_11231,N_11414);
nand U11769 (N_11769,N_11350,N_11203);
nand U11770 (N_11770,N_11337,N_11322);
nor U11771 (N_11771,N_11581,N_11571);
nand U11772 (N_11772,N_11401,N_11555);
and U11773 (N_11773,N_11403,N_11416);
xor U11774 (N_11774,N_11489,N_11419);
xnor U11775 (N_11775,N_11293,N_11309);
nor U11776 (N_11776,N_11263,N_11545);
nor U11777 (N_11777,N_11250,N_11316);
nand U11778 (N_11778,N_11252,N_11541);
and U11779 (N_11779,N_11372,N_11537);
xnor U11780 (N_11780,N_11393,N_11254);
nand U11781 (N_11781,N_11559,N_11420);
nand U11782 (N_11782,N_11378,N_11381);
or U11783 (N_11783,N_11431,N_11519);
and U11784 (N_11784,N_11244,N_11564);
nand U11785 (N_11785,N_11485,N_11347);
or U11786 (N_11786,N_11365,N_11288);
and U11787 (N_11787,N_11374,N_11228);
nor U11788 (N_11788,N_11311,N_11389);
xnor U11789 (N_11789,N_11472,N_11573);
nor U11790 (N_11790,N_11574,N_11561);
nor U11791 (N_11791,N_11484,N_11504);
and U11792 (N_11792,N_11324,N_11373);
xor U11793 (N_11793,N_11478,N_11281);
or U11794 (N_11794,N_11590,N_11503);
and U11795 (N_11795,N_11298,N_11326);
xor U11796 (N_11796,N_11476,N_11570);
or U11797 (N_11797,N_11404,N_11204);
nor U11798 (N_11798,N_11576,N_11586);
xnor U11799 (N_11799,N_11547,N_11530);
nor U11800 (N_11800,N_11402,N_11510);
or U11801 (N_11801,N_11208,N_11580);
nor U11802 (N_11802,N_11236,N_11216);
and U11803 (N_11803,N_11496,N_11387);
nor U11804 (N_11804,N_11351,N_11545);
nand U11805 (N_11805,N_11501,N_11544);
and U11806 (N_11806,N_11512,N_11425);
nor U11807 (N_11807,N_11554,N_11236);
xor U11808 (N_11808,N_11250,N_11540);
nand U11809 (N_11809,N_11494,N_11241);
nand U11810 (N_11810,N_11336,N_11525);
xor U11811 (N_11811,N_11274,N_11396);
or U11812 (N_11812,N_11575,N_11561);
and U11813 (N_11813,N_11253,N_11246);
nand U11814 (N_11814,N_11443,N_11339);
and U11815 (N_11815,N_11256,N_11230);
and U11816 (N_11816,N_11229,N_11332);
and U11817 (N_11817,N_11593,N_11245);
or U11818 (N_11818,N_11548,N_11411);
nand U11819 (N_11819,N_11406,N_11349);
xor U11820 (N_11820,N_11326,N_11481);
or U11821 (N_11821,N_11564,N_11204);
and U11822 (N_11822,N_11393,N_11450);
or U11823 (N_11823,N_11274,N_11416);
and U11824 (N_11824,N_11471,N_11242);
nand U11825 (N_11825,N_11359,N_11207);
nand U11826 (N_11826,N_11425,N_11422);
xor U11827 (N_11827,N_11578,N_11285);
nor U11828 (N_11828,N_11263,N_11508);
and U11829 (N_11829,N_11363,N_11421);
or U11830 (N_11830,N_11318,N_11490);
or U11831 (N_11831,N_11312,N_11386);
xnor U11832 (N_11832,N_11515,N_11438);
xor U11833 (N_11833,N_11275,N_11284);
or U11834 (N_11834,N_11313,N_11562);
or U11835 (N_11835,N_11447,N_11404);
nand U11836 (N_11836,N_11447,N_11409);
or U11837 (N_11837,N_11315,N_11409);
or U11838 (N_11838,N_11283,N_11566);
xor U11839 (N_11839,N_11243,N_11442);
or U11840 (N_11840,N_11432,N_11215);
nand U11841 (N_11841,N_11589,N_11349);
nor U11842 (N_11842,N_11241,N_11434);
and U11843 (N_11843,N_11350,N_11562);
nor U11844 (N_11844,N_11291,N_11476);
or U11845 (N_11845,N_11400,N_11577);
or U11846 (N_11846,N_11497,N_11205);
nand U11847 (N_11847,N_11353,N_11214);
xnor U11848 (N_11848,N_11247,N_11467);
nand U11849 (N_11849,N_11348,N_11536);
xor U11850 (N_11850,N_11474,N_11424);
xnor U11851 (N_11851,N_11530,N_11412);
or U11852 (N_11852,N_11576,N_11226);
and U11853 (N_11853,N_11499,N_11268);
or U11854 (N_11854,N_11549,N_11226);
xor U11855 (N_11855,N_11312,N_11271);
nand U11856 (N_11856,N_11399,N_11290);
nor U11857 (N_11857,N_11206,N_11373);
xor U11858 (N_11858,N_11478,N_11509);
nand U11859 (N_11859,N_11328,N_11425);
nand U11860 (N_11860,N_11460,N_11542);
and U11861 (N_11861,N_11392,N_11380);
nand U11862 (N_11862,N_11473,N_11564);
nand U11863 (N_11863,N_11504,N_11381);
or U11864 (N_11864,N_11207,N_11564);
xor U11865 (N_11865,N_11494,N_11364);
nand U11866 (N_11866,N_11477,N_11503);
nand U11867 (N_11867,N_11503,N_11428);
xor U11868 (N_11868,N_11374,N_11236);
or U11869 (N_11869,N_11493,N_11274);
nor U11870 (N_11870,N_11235,N_11494);
xor U11871 (N_11871,N_11210,N_11515);
xnor U11872 (N_11872,N_11411,N_11203);
or U11873 (N_11873,N_11308,N_11239);
nor U11874 (N_11874,N_11389,N_11480);
xor U11875 (N_11875,N_11481,N_11478);
xnor U11876 (N_11876,N_11233,N_11330);
and U11877 (N_11877,N_11318,N_11535);
nor U11878 (N_11878,N_11432,N_11303);
and U11879 (N_11879,N_11458,N_11398);
and U11880 (N_11880,N_11438,N_11341);
or U11881 (N_11881,N_11288,N_11424);
and U11882 (N_11882,N_11492,N_11207);
nor U11883 (N_11883,N_11336,N_11473);
xor U11884 (N_11884,N_11249,N_11490);
xnor U11885 (N_11885,N_11507,N_11311);
nor U11886 (N_11886,N_11283,N_11485);
or U11887 (N_11887,N_11435,N_11312);
and U11888 (N_11888,N_11596,N_11430);
nand U11889 (N_11889,N_11376,N_11364);
and U11890 (N_11890,N_11237,N_11253);
nand U11891 (N_11891,N_11519,N_11547);
nand U11892 (N_11892,N_11365,N_11470);
or U11893 (N_11893,N_11373,N_11552);
nand U11894 (N_11894,N_11547,N_11542);
or U11895 (N_11895,N_11566,N_11392);
nand U11896 (N_11896,N_11465,N_11475);
nand U11897 (N_11897,N_11303,N_11576);
nor U11898 (N_11898,N_11330,N_11293);
nand U11899 (N_11899,N_11503,N_11359);
nor U11900 (N_11900,N_11517,N_11460);
nor U11901 (N_11901,N_11561,N_11438);
and U11902 (N_11902,N_11298,N_11473);
or U11903 (N_11903,N_11436,N_11443);
nand U11904 (N_11904,N_11299,N_11513);
nand U11905 (N_11905,N_11339,N_11222);
or U11906 (N_11906,N_11538,N_11453);
nor U11907 (N_11907,N_11488,N_11433);
and U11908 (N_11908,N_11474,N_11508);
nor U11909 (N_11909,N_11386,N_11374);
xor U11910 (N_11910,N_11412,N_11510);
or U11911 (N_11911,N_11252,N_11491);
and U11912 (N_11912,N_11567,N_11274);
or U11913 (N_11913,N_11529,N_11402);
or U11914 (N_11914,N_11530,N_11559);
nor U11915 (N_11915,N_11343,N_11595);
nor U11916 (N_11916,N_11532,N_11473);
or U11917 (N_11917,N_11309,N_11502);
nor U11918 (N_11918,N_11354,N_11231);
xor U11919 (N_11919,N_11347,N_11282);
xnor U11920 (N_11920,N_11450,N_11594);
and U11921 (N_11921,N_11353,N_11341);
nor U11922 (N_11922,N_11263,N_11210);
nand U11923 (N_11923,N_11271,N_11396);
and U11924 (N_11924,N_11232,N_11399);
xor U11925 (N_11925,N_11381,N_11418);
nor U11926 (N_11926,N_11262,N_11275);
nand U11927 (N_11927,N_11435,N_11365);
xor U11928 (N_11928,N_11509,N_11227);
and U11929 (N_11929,N_11312,N_11224);
nand U11930 (N_11930,N_11210,N_11594);
or U11931 (N_11931,N_11329,N_11246);
xor U11932 (N_11932,N_11529,N_11296);
nand U11933 (N_11933,N_11223,N_11265);
and U11934 (N_11934,N_11586,N_11219);
or U11935 (N_11935,N_11276,N_11233);
nor U11936 (N_11936,N_11349,N_11460);
nand U11937 (N_11937,N_11313,N_11431);
nand U11938 (N_11938,N_11563,N_11362);
and U11939 (N_11939,N_11493,N_11213);
nor U11940 (N_11940,N_11520,N_11206);
or U11941 (N_11941,N_11366,N_11340);
or U11942 (N_11942,N_11215,N_11316);
nor U11943 (N_11943,N_11424,N_11485);
nor U11944 (N_11944,N_11417,N_11480);
xnor U11945 (N_11945,N_11412,N_11489);
and U11946 (N_11946,N_11549,N_11224);
and U11947 (N_11947,N_11485,N_11219);
xnor U11948 (N_11948,N_11467,N_11374);
or U11949 (N_11949,N_11430,N_11284);
nor U11950 (N_11950,N_11450,N_11368);
xor U11951 (N_11951,N_11305,N_11318);
or U11952 (N_11952,N_11274,N_11562);
and U11953 (N_11953,N_11295,N_11398);
nand U11954 (N_11954,N_11242,N_11210);
nor U11955 (N_11955,N_11310,N_11405);
nor U11956 (N_11956,N_11288,N_11380);
or U11957 (N_11957,N_11345,N_11477);
or U11958 (N_11958,N_11218,N_11219);
nand U11959 (N_11959,N_11574,N_11447);
xor U11960 (N_11960,N_11593,N_11406);
and U11961 (N_11961,N_11566,N_11299);
nand U11962 (N_11962,N_11529,N_11557);
nor U11963 (N_11963,N_11232,N_11251);
and U11964 (N_11964,N_11542,N_11543);
xor U11965 (N_11965,N_11377,N_11230);
nand U11966 (N_11966,N_11448,N_11287);
xnor U11967 (N_11967,N_11507,N_11590);
or U11968 (N_11968,N_11542,N_11258);
and U11969 (N_11969,N_11435,N_11393);
nor U11970 (N_11970,N_11281,N_11218);
xor U11971 (N_11971,N_11478,N_11233);
and U11972 (N_11972,N_11361,N_11459);
nand U11973 (N_11973,N_11554,N_11396);
nor U11974 (N_11974,N_11249,N_11376);
xnor U11975 (N_11975,N_11565,N_11324);
nor U11976 (N_11976,N_11247,N_11561);
nor U11977 (N_11977,N_11409,N_11344);
nor U11978 (N_11978,N_11309,N_11447);
and U11979 (N_11979,N_11313,N_11511);
xnor U11980 (N_11980,N_11246,N_11261);
nand U11981 (N_11981,N_11258,N_11338);
and U11982 (N_11982,N_11494,N_11596);
nor U11983 (N_11983,N_11539,N_11511);
and U11984 (N_11984,N_11207,N_11531);
xnor U11985 (N_11985,N_11415,N_11462);
nor U11986 (N_11986,N_11318,N_11567);
xor U11987 (N_11987,N_11255,N_11213);
xor U11988 (N_11988,N_11582,N_11507);
and U11989 (N_11989,N_11297,N_11556);
and U11990 (N_11990,N_11381,N_11512);
or U11991 (N_11991,N_11232,N_11368);
nor U11992 (N_11992,N_11369,N_11270);
xnor U11993 (N_11993,N_11543,N_11454);
or U11994 (N_11994,N_11419,N_11541);
xor U11995 (N_11995,N_11599,N_11546);
or U11996 (N_11996,N_11595,N_11392);
nand U11997 (N_11997,N_11286,N_11375);
nand U11998 (N_11998,N_11439,N_11212);
and U11999 (N_11999,N_11575,N_11460);
nor U12000 (N_12000,N_11992,N_11883);
nand U12001 (N_12001,N_11752,N_11764);
and U12002 (N_12002,N_11805,N_11945);
or U12003 (N_12003,N_11645,N_11792);
and U12004 (N_12004,N_11654,N_11985);
and U12005 (N_12005,N_11889,N_11675);
xor U12006 (N_12006,N_11920,N_11677);
or U12007 (N_12007,N_11924,N_11832);
nor U12008 (N_12008,N_11751,N_11952);
nand U12009 (N_12009,N_11875,N_11679);
nor U12010 (N_12010,N_11714,N_11624);
nor U12011 (N_12011,N_11600,N_11772);
xor U12012 (N_12012,N_11735,N_11803);
and U12013 (N_12013,N_11634,N_11800);
nand U12014 (N_12014,N_11930,N_11818);
nand U12015 (N_12015,N_11902,N_11630);
and U12016 (N_12016,N_11746,N_11975);
xnor U12017 (N_12017,N_11641,N_11936);
xor U12018 (N_12018,N_11928,N_11857);
and U12019 (N_12019,N_11865,N_11948);
xnor U12020 (N_12020,N_11726,N_11835);
nor U12021 (N_12021,N_11728,N_11842);
xnor U12022 (N_12022,N_11874,N_11963);
nor U12023 (N_12023,N_11947,N_11760);
xnor U12024 (N_12024,N_11774,N_11906);
or U12025 (N_12025,N_11721,N_11946);
nor U12026 (N_12026,N_11724,N_11727);
and U12027 (N_12027,N_11967,N_11779);
xnor U12028 (N_12028,N_11601,N_11744);
nor U12029 (N_12029,N_11910,N_11864);
xor U12030 (N_12030,N_11895,N_11608);
or U12031 (N_12031,N_11999,N_11637);
and U12032 (N_12032,N_11648,N_11871);
and U12033 (N_12033,N_11915,N_11885);
xnor U12034 (N_12034,N_11824,N_11662);
and U12035 (N_12035,N_11762,N_11738);
and U12036 (N_12036,N_11711,N_11768);
or U12037 (N_12037,N_11907,N_11862);
or U12038 (N_12038,N_11918,N_11944);
nand U12039 (N_12039,N_11604,N_11831);
nand U12040 (N_12040,N_11770,N_11827);
nor U12041 (N_12041,N_11949,N_11644);
nand U12042 (N_12042,N_11861,N_11696);
or U12043 (N_12043,N_11845,N_11739);
nor U12044 (N_12044,N_11681,N_11778);
and U12045 (N_12045,N_11761,N_11841);
or U12046 (N_12046,N_11625,N_11622);
xnor U12047 (N_12047,N_11937,N_11697);
xor U12048 (N_12048,N_11694,N_11893);
or U12049 (N_12049,N_11825,N_11847);
and U12050 (N_12050,N_11747,N_11629);
and U12051 (N_12051,N_11984,N_11958);
nand U12052 (N_12052,N_11880,N_11932);
nand U12053 (N_12053,N_11607,N_11969);
or U12054 (N_12054,N_11602,N_11631);
xor U12055 (N_12055,N_11713,N_11627);
or U12056 (N_12056,N_11923,N_11700);
xor U12057 (N_12057,N_11689,N_11703);
xnor U12058 (N_12058,N_11954,N_11725);
or U12059 (N_12059,N_11796,N_11849);
nand U12060 (N_12060,N_11609,N_11722);
or U12061 (N_12061,N_11891,N_11605);
nand U12062 (N_12062,N_11968,N_11823);
xor U12063 (N_12063,N_11898,N_11733);
or U12064 (N_12064,N_11717,N_11745);
nor U12065 (N_12065,N_11974,N_11633);
and U12066 (N_12066,N_11705,N_11942);
and U12067 (N_12067,N_11716,N_11894);
and U12068 (N_12068,N_11646,N_11672);
nor U12069 (N_12069,N_11990,N_11685);
nand U12070 (N_12070,N_11908,N_11757);
nor U12071 (N_12071,N_11647,N_11780);
and U12072 (N_12072,N_11776,N_11979);
nand U12073 (N_12073,N_11855,N_11632);
xor U12074 (N_12074,N_11859,N_11994);
nand U12075 (N_12075,N_11663,N_11678);
nand U12076 (N_12076,N_11931,N_11927);
and U12077 (N_12077,N_11753,N_11955);
nand U12078 (N_12078,N_11953,N_11731);
and U12079 (N_12079,N_11765,N_11635);
xor U12080 (N_12080,N_11988,N_11998);
xor U12081 (N_12081,N_11971,N_11695);
xor U12082 (N_12082,N_11686,N_11900);
or U12083 (N_12083,N_11884,N_11965);
or U12084 (N_12084,N_11702,N_11858);
or U12085 (N_12085,N_11653,N_11754);
nor U12086 (N_12086,N_11743,N_11795);
and U12087 (N_12087,N_11806,N_11950);
xnor U12088 (N_12088,N_11966,N_11655);
nor U12089 (N_12089,N_11737,N_11851);
nor U12090 (N_12090,N_11708,N_11904);
and U12091 (N_12091,N_11844,N_11781);
xnor U12092 (N_12092,N_11652,N_11877);
xnor U12093 (N_12093,N_11793,N_11804);
xnor U12094 (N_12094,N_11651,N_11667);
nor U12095 (N_12095,N_11960,N_11812);
or U12096 (N_12096,N_11987,N_11640);
nor U12097 (N_12097,N_11892,N_11623);
and U12098 (N_12098,N_11973,N_11661);
and U12099 (N_12099,N_11710,N_11976);
nor U12100 (N_12100,N_11811,N_11993);
nand U12101 (N_12101,N_11962,N_11912);
or U12102 (N_12102,N_11836,N_11938);
nor U12103 (N_12103,N_11911,N_11621);
or U12104 (N_12104,N_11665,N_11767);
nand U12105 (N_12105,N_11991,N_11863);
nand U12106 (N_12106,N_11660,N_11669);
and U12107 (N_12107,N_11801,N_11750);
or U12108 (N_12108,N_11788,N_11913);
and U12109 (N_12109,N_11852,N_11748);
or U12110 (N_12110,N_11899,N_11870);
or U12111 (N_12111,N_11682,N_11785);
nand U12112 (N_12112,N_11706,N_11939);
nand U12113 (N_12113,N_11691,N_11876);
nor U12114 (N_12114,N_11715,N_11850);
and U12115 (N_12115,N_11941,N_11828);
or U12116 (N_12116,N_11742,N_11854);
xnor U12117 (N_12117,N_11934,N_11896);
nor U12118 (N_12118,N_11964,N_11867);
nand U12119 (N_12119,N_11869,N_11612);
xnor U12120 (N_12120,N_11698,N_11814);
xor U12121 (N_12121,N_11903,N_11668);
nor U12122 (N_12122,N_11970,N_11997);
or U12123 (N_12123,N_11807,N_11839);
xor U12124 (N_12124,N_11853,N_11688);
nand U12125 (N_12125,N_11989,N_11886);
or U12126 (N_12126,N_11933,N_11618);
nand U12127 (N_12127,N_11943,N_11759);
or U12128 (N_12128,N_11773,N_11914);
and U12129 (N_12129,N_11787,N_11756);
and U12130 (N_12130,N_11916,N_11816);
nand U12131 (N_12131,N_11926,N_11643);
nor U12132 (N_12132,N_11673,N_11638);
and U12133 (N_12133,N_11956,N_11817);
or U12134 (N_12134,N_11690,N_11771);
and U12135 (N_12135,N_11840,N_11784);
xnor U12136 (N_12136,N_11866,N_11718);
xnor U12137 (N_12137,N_11878,N_11611);
xnor U12138 (N_12138,N_11704,N_11873);
nand U12139 (N_12139,N_11740,N_11656);
xnor U12140 (N_12140,N_11657,N_11977);
nand U12141 (N_12141,N_11613,N_11909);
or U12142 (N_12142,N_11868,N_11972);
nor U12143 (N_12143,N_11846,N_11603);
nor U12144 (N_12144,N_11917,N_11712);
nand U12145 (N_12145,N_11794,N_11996);
nand U12146 (N_12146,N_11775,N_11922);
xor U12147 (N_12147,N_11755,N_11766);
and U12148 (N_12148,N_11674,N_11925);
and U12149 (N_12149,N_11741,N_11616);
nor U12150 (N_12150,N_11730,N_11692);
or U12151 (N_12151,N_11838,N_11642);
or U12152 (N_12152,N_11882,N_11980);
or U12153 (N_12153,N_11986,N_11790);
and U12154 (N_12154,N_11940,N_11758);
and U12155 (N_12155,N_11670,N_11981);
xor U12156 (N_12156,N_11782,N_11821);
or U12157 (N_12157,N_11736,N_11961);
and U12158 (N_12158,N_11887,N_11606);
nor U12159 (N_12159,N_11872,N_11734);
xor U12160 (N_12160,N_11628,N_11732);
and U12161 (N_12161,N_11856,N_11783);
nor U12162 (N_12162,N_11723,N_11901);
nor U12163 (N_12163,N_11709,N_11664);
or U12164 (N_12164,N_11905,N_11881);
nand U12165 (N_12165,N_11995,N_11684);
or U12166 (N_12166,N_11819,N_11610);
xor U12167 (N_12167,N_11626,N_11890);
xor U12168 (N_12168,N_11809,N_11799);
or U12169 (N_12169,N_11769,N_11815);
xor U12170 (N_12170,N_11837,N_11888);
nor U12171 (N_12171,N_11982,N_11649);
nand U12172 (N_12172,N_11830,N_11719);
or U12173 (N_12173,N_11919,N_11834);
xor U12174 (N_12174,N_11951,N_11683);
nand U12175 (N_12175,N_11978,N_11935);
nor U12176 (N_12176,N_11879,N_11789);
or U12177 (N_12177,N_11791,N_11615);
nor U12178 (N_12178,N_11699,N_11720);
or U12179 (N_12179,N_11822,N_11810);
nor U12180 (N_12180,N_11650,N_11833);
nand U12181 (N_12181,N_11826,N_11617);
xnor U12182 (N_12182,N_11983,N_11959);
xnor U12183 (N_12183,N_11676,N_11636);
nand U12184 (N_12184,N_11666,N_11813);
and U12185 (N_12185,N_11619,N_11620);
and U12186 (N_12186,N_11749,N_11848);
nor U12187 (N_12187,N_11921,N_11701);
or U12188 (N_12188,N_11786,N_11820);
nor U12189 (N_12189,N_11860,N_11808);
nor U12190 (N_12190,N_11929,N_11763);
xor U12191 (N_12191,N_11707,N_11897);
nor U12192 (N_12192,N_11957,N_11658);
and U12193 (N_12193,N_11671,N_11829);
or U12194 (N_12194,N_11693,N_11843);
and U12195 (N_12195,N_11659,N_11797);
nand U12196 (N_12196,N_11639,N_11729);
and U12197 (N_12197,N_11680,N_11614);
and U12198 (N_12198,N_11687,N_11777);
and U12199 (N_12199,N_11802,N_11798);
xor U12200 (N_12200,N_11622,N_11786);
nor U12201 (N_12201,N_11910,N_11665);
or U12202 (N_12202,N_11826,N_11657);
or U12203 (N_12203,N_11725,N_11693);
nor U12204 (N_12204,N_11899,N_11754);
xnor U12205 (N_12205,N_11780,N_11752);
nand U12206 (N_12206,N_11825,N_11735);
xor U12207 (N_12207,N_11601,N_11847);
and U12208 (N_12208,N_11839,N_11826);
xnor U12209 (N_12209,N_11753,N_11863);
and U12210 (N_12210,N_11758,N_11864);
nand U12211 (N_12211,N_11672,N_11987);
nand U12212 (N_12212,N_11620,N_11932);
xnor U12213 (N_12213,N_11876,N_11645);
or U12214 (N_12214,N_11724,N_11995);
xnor U12215 (N_12215,N_11991,N_11708);
xnor U12216 (N_12216,N_11903,N_11651);
nor U12217 (N_12217,N_11948,N_11695);
or U12218 (N_12218,N_11776,N_11875);
and U12219 (N_12219,N_11680,N_11875);
nor U12220 (N_12220,N_11978,N_11647);
xor U12221 (N_12221,N_11757,N_11801);
xor U12222 (N_12222,N_11662,N_11925);
and U12223 (N_12223,N_11615,N_11901);
or U12224 (N_12224,N_11692,N_11617);
xnor U12225 (N_12225,N_11842,N_11931);
nand U12226 (N_12226,N_11993,N_11653);
nor U12227 (N_12227,N_11889,N_11932);
and U12228 (N_12228,N_11617,N_11767);
nand U12229 (N_12229,N_11625,N_11714);
xor U12230 (N_12230,N_11645,N_11854);
nand U12231 (N_12231,N_11988,N_11720);
or U12232 (N_12232,N_11668,N_11704);
or U12233 (N_12233,N_11655,N_11893);
nand U12234 (N_12234,N_11733,N_11676);
and U12235 (N_12235,N_11872,N_11893);
nor U12236 (N_12236,N_11906,N_11861);
nand U12237 (N_12237,N_11877,N_11799);
xor U12238 (N_12238,N_11717,N_11813);
or U12239 (N_12239,N_11899,N_11816);
nor U12240 (N_12240,N_11660,N_11628);
nand U12241 (N_12241,N_11875,N_11879);
and U12242 (N_12242,N_11646,N_11807);
nand U12243 (N_12243,N_11986,N_11601);
or U12244 (N_12244,N_11852,N_11676);
or U12245 (N_12245,N_11940,N_11822);
and U12246 (N_12246,N_11859,N_11694);
xor U12247 (N_12247,N_11885,N_11717);
xor U12248 (N_12248,N_11641,N_11604);
xor U12249 (N_12249,N_11864,N_11971);
nand U12250 (N_12250,N_11742,N_11730);
nor U12251 (N_12251,N_11744,N_11765);
and U12252 (N_12252,N_11850,N_11703);
and U12253 (N_12253,N_11669,N_11744);
and U12254 (N_12254,N_11831,N_11651);
xnor U12255 (N_12255,N_11731,N_11668);
nor U12256 (N_12256,N_11635,N_11993);
xor U12257 (N_12257,N_11947,N_11691);
and U12258 (N_12258,N_11611,N_11979);
or U12259 (N_12259,N_11652,N_11983);
and U12260 (N_12260,N_11833,N_11776);
nor U12261 (N_12261,N_11984,N_11783);
and U12262 (N_12262,N_11853,N_11858);
nand U12263 (N_12263,N_11828,N_11821);
or U12264 (N_12264,N_11852,N_11979);
nand U12265 (N_12265,N_11733,N_11665);
or U12266 (N_12266,N_11883,N_11740);
nor U12267 (N_12267,N_11651,N_11623);
xor U12268 (N_12268,N_11710,N_11643);
or U12269 (N_12269,N_11729,N_11892);
nor U12270 (N_12270,N_11805,N_11780);
or U12271 (N_12271,N_11617,N_11722);
xor U12272 (N_12272,N_11856,N_11959);
and U12273 (N_12273,N_11864,N_11600);
or U12274 (N_12274,N_11865,N_11601);
nor U12275 (N_12275,N_11733,N_11705);
and U12276 (N_12276,N_11706,N_11739);
nor U12277 (N_12277,N_11600,N_11704);
nor U12278 (N_12278,N_11660,N_11887);
nor U12279 (N_12279,N_11844,N_11717);
or U12280 (N_12280,N_11650,N_11893);
xnor U12281 (N_12281,N_11972,N_11744);
xnor U12282 (N_12282,N_11712,N_11636);
and U12283 (N_12283,N_11652,N_11709);
nand U12284 (N_12284,N_11900,N_11696);
or U12285 (N_12285,N_11999,N_11771);
xor U12286 (N_12286,N_11919,N_11741);
or U12287 (N_12287,N_11753,N_11962);
nor U12288 (N_12288,N_11983,N_11809);
nand U12289 (N_12289,N_11706,N_11900);
or U12290 (N_12290,N_11986,N_11741);
nand U12291 (N_12291,N_11795,N_11686);
and U12292 (N_12292,N_11648,N_11897);
or U12293 (N_12293,N_11769,N_11935);
and U12294 (N_12294,N_11770,N_11622);
and U12295 (N_12295,N_11684,N_11961);
nand U12296 (N_12296,N_11935,N_11726);
nor U12297 (N_12297,N_11865,N_11982);
or U12298 (N_12298,N_11813,N_11866);
xnor U12299 (N_12299,N_11767,N_11836);
nor U12300 (N_12300,N_11688,N_11812);
nand U12301 (N_12301,N_11650,N_11797);
xor U12302 (N_12302,N_11694,N_11750);
and U12303 (N_12303,N_11628,N_11751);
xor U12304 (N_12304,N_11845,N_11992);
or U12305 (N_12305,N_11732,N_11986);
nor U12306 (N_12306,N_11880,N_11728);
nand U12307 (N_12307,N_11817,N_11954);
xor U12308 (N_12308,N_11768,N_11910);
or U12309 (N_12309,N_11968,N_11677);
nand U12310 (N_12310,N_11948,N_11612);
and U12311 (N_12311,N_11829,N_11979);
nor U12312 (N_12312,N_11855,N_11962);
or U12313 (N_12313,N_11603,N_11775);
nand U12314 (N_12314,N_11879,N_11646);
xnor U12315 (N_12315,N_11685,N_11770);
and U12316 (N_12316,N_11798,N_11839);
or U12317 (N_12317,N_11981,N_11966);
xnor U12318 (N_12318,N_11781,N_11957);
xnor U12319 (N_12319,N_11945,N_11947);
or U12320 (N_12320,N_11744,N_11852);
or U12321 (N_12321,N_11633,N_11657);
or U12322 (N_12322,N_11879,N_11630);
and U12323 (N_12323,N_11862,N_11600);
and U12324 (N_12324,N_11769,N_11871);
nor U12325 (N_12325,N_11713,N_11726);
or U12326 (N_12326,N_11691,N_11692);
nand U12327 (N_12327,N_11887,N_11777);
nand U12328 (N_12328,N_11695,N_11769);
nand U12329 (N_12329,N_11610,N_11900);
nand U12330 (N_12330,N_11648,N_11793);
and U12331 (N_12331,N_11654,N_11649);
nand U12332 (N_12332,N_11723,N_11933);
and U12333 (N_12333,N_11612,N_11616);
and U12334 (N_12334,N_11956,N_11731);
and U12335 (N_12335,N_11965,N_11737);
nand U12336 (N_12336,N_11911,N_11837);
nor U12337 (N_12337,N_11860,N_11940);
and U12338 (N_12338,N_11726,N_11869);
nor U12339 (N_12339,N_11868,N_11933);
xnor U12340 (N_12340,N_11679,N_11917);
nand U12341 (N_12341,N_11664,N_11645);
xnor U12342 (N_12342,N_11795,N_11641);
or U12343 (N_12343,N_11779,N_11723);
xor U12344 (N_12344,N_11847,N_11861);
xnor U12345 (N_12345,N_11769,N_11892);
and U12346 (N_12346,N_11824,N_11822);
and U12347 (N_12347,N_11748,N_11807);
xnor U12348 (N_12348,N_11633,N_11782);
nand U12349 (N_12349,N_11737,N_11759);
nor U12350 (N_12350,N_11663,N_11856);
nand U12351 (N_12351,N_11647,N_11614);
or U12352 (N_12352,N_11664,N_11955);
nand U12353 (N_12353,N_11807,N_11886);
xor U12354 (N_12354,N_11874,N_11684);
nor U12355 (N_12355,N_11883,N_11954);
xnor U12356 (N_12356,N_11913,N_11985);
or U12357 (N_12357,N_11779,N_11905);
or U12358 (N_12358,N_11853,N_11757);
or U12359 (N_12359,N_11738,N_11855);
nor U12360 (N_12360,N_11643,N_11947);
xnor U12361 (N_12361,N_11869,N_11677);
or U12362 (N_12362,N_11650,N_11944);
nor U12363 (N_12363,N_11886,N_11823);
nor U12364 (N_12364,N_11749,N_11732);
and U12365 (N_12365,N_11695,N_11911);
nor U12366 (N_12366,N_11968,N_11804);
nand U12367 (N_12367,N_11950,N_11661);
xnor U12368 (N_12368,N_11669,N_11786);
xnor U12369 (N_12369,N_11772,N_11705);
nand U12370 (N_12370,N_11821,N_11600);
or U12371 (N_12371,N_11792,N_11853);
nor U12372 (N_12372,N_11629,N_11968);
nand U12373 (N_12373,N_11666,N_11932);
nand U12374 (N_12374,N_11902,N_11609);
and U12375 (N_12375,N_11622,N_11843);
xnor U12376 (N_12376,N_11749,N_11704);
nor U12377 (N_12377,N_11683,N_11972);
nand U12378 (N_12378,N_11668,N_11894);
xor U12379 (N_12379,N_11689,N_11686);
and U12380 (N_12380,N_11961,N_11965);
nand U12381 (N_12381,N_11735,N_11757);
xor U12382 (N_12382,N_11914,N_11719);
nand U12383 (N_12383,N_11649,N_11920);
xor U12384 (N_12384,N_11685,N_11660);
xor U12385 (N_12385,N_11765,N_11935);
and U12386 (N_12386,N_11706,N_11713);
nor U12387 (N_12387,N_11956,N_11966);
nand U12388 (N_12388,N_11713,N_11730);
xnor U12389 (N_12389,N_11671,N_11655);
or U12390 (N_12390,N_11784,N_11655);
nor U12391 (N_12391,N_11915,N_11821);
and U12392 (N_12392,N_11666,N_11790);
xnor U12393 (N_12393,N_11785,N_11676);
xor U12394 (N_12394,N_11639,N_11985);
xnor U12395 (N_12395,N_11618,N_11700);
and U12396 (N_12396,N_11868,N_11998);
nor U12397 (N_12397,N_11865,N_11835);
xor U12398 (N_12398,N_11717,N_11649);
nand U12399 (N_12399,N_11888,N_11732);
and U12400 (N_12400,N_12133,N_12252);
and U12401 (N_12401,N_12311,N_12233);
nand U12402 (N_12402,N_12157,N_12213);
and U12403 (N_12403,N_12281,N_12178);
xor U12404 (N_12404,N_12339,N_12345);
xor U12405 (N_12405,N_12117,N_12026);
xor U12406 (N_12406,N_12383,N_12371);
xnor U12407 (N_12407,N_12154,N_12153);
nand U12408 (N_12408,N_12007,N_12019);
xor U12409 (N_12409,N_12300,N_12273);
and U12410 (N_12410,N_12167,N_12090);
and U12411 (N_12411,N_12220,N_12299);
nand U12412 (N_12412,N_12104,N_12063);
and U12413 (N_12413,N_12195,N_12257);
nor U12414 (N_12414,N_12386,N_12150);
and U12415 (N_12415,N_12034,N_12155);
nand U12416 (N_12416,N_12262,N_12002);
or U12417 (N_12417,N_12319,N_12081);
xor U12418 (N_12418,N_12175,N_12358);
nor U12419 (N_12419,N_12335,N_12318);
or U12420 (N_12420,N_12087,N_12190);
nor U12421 (N_12421,N_12059,N_12096);
and U12422 (N_12422,N_12072,N_12303);
xor U12423 (N_12423,N_12160,N_12320);
nand U12424 (N_12424,N_12075,N_12332);
nor U12425 (N_12425,N_12103,N_12171);
nor U12426 (N_12426,N_12056,N_12214);
or U12427 (N_12427,N_12264,N_12395);
and U12428 (N_12428,N_12239,N_12014);
or U12429 (N_12429,N_12125,N_12306);
and U12430 (N_12430,N_12290,N_12271);
or U12431 (N_12431,N_12298,N_12192);
nand U12432 (N_12432,N_12084,N_12279);
xnor U12433 (N_12433,N_12206,N_12392);
or U12434 (N_12434,N_12200,N_12078);
xnor U12435 (N_12435,N_12127,N_12101);
nor U12436 (N_12436,N_12194,N_12069);
or U12437 (N_12437,N_12259,N_12006);
or U12438 (N_12438,N_12315,N_12212);
or U12439 (N_12439,N_12169,N_12211);
nor U12440 (N_12440,N_12140,N_12391);
xor U12441 (N_12441,N_12137,N_12004);
and U12442 (N_12442,N_12086,N_12361);
xnor U12443 (N_12443,N_12376,N_12053);
or U12444 (N_12444,N_12393,N_12149);
xnor U12445 (N_12445,N_12367,N_12107);
nand U12446 (N_12446,N_12351,N_12088);
nand U12447 (N_12447,N_12397,N_12139);
and U12448 (N_12448,N_12106,N_12246);
nor U12449 (N_12449,N_12049,N_12020);
or U12450 (N_12450,N_12256,N_12164);
or U12451 (N_12451,N_12050,N_12305);
and U12452 (N_12452,N_12394,N_12028);
nand U12453 (N_12453,N_12374,N_12205);
nor U12454 (N_12454,N_12384,N_12382);
nand U12455 (N_12455,N_12191,N_12209);
and U12456 (N_12456,N_12349,N_12046);
nand U12457 (N_12457,N_12285,N_12263);
nand U12458 (N_12458,N_12143,N_12141);
nor U12459 (N_12459,N_12027,N_12276);
nand U12460 (N_12460,N_12032,N_12301);
nor U12461 (N_12461,N_12013,N_12093);
and U12462 (N_12462,N_12022,N_12001);
and U12463 (N_12463,N_12323,N_12197);
and U12464 (N_12464,N_12180,N_12168);
nand U12465 (N_12465,N_12011,N_12296);
nand U12466 (N_12466,N_12362,N_12341);
xnor U12467 (N_12467,N_12291,N_12017);
or U12468 (N_12468,N_12328,N_12282);
and U12469 (N_12469,N_12280,N_12151);
xnor U12470 (N_12470,N_12105,N_12068);
nand U12471 (N_12471,N_12399,N_12148);
and U12472 (N_12472,N_12366,N_12166);
xor U12473 (N_12473,N_12184,N_12333);
or U12474 (N_12474,N_12009,N_12289);
xor U12475 (N_12475,N_12097,N_12207);
or U12476 (N_12476,N_12284,N_12360);
nand U12477 (N_12477,N_12120,N_12066);
and U12478 (N_12478,N_12052,N_12309);
xor U12479 (N_12479,N_12136,N_12265);
nand U12480 (N_12480,N_12181,N_12179);
xnor U12481 (N_12481,N_12045,N_12018);
nor U12482 (N_12482,N_12129,N_12238);
nor U12483 (N_12483,N_12354,N_12077);
and U12484 (N_12484,N_12132,N_12226);
nand U12485 (N_12485,N_12111,N_12249);
xor U12486 (N_12486,N_12352,N_12185);
nor U12487 (N_12487,N_12234,N_12251);
and U12488 (N_12488,N_12091,N_12230);
nand U12489 (N_12489,N_12219,N_12037);
and U12490 (N_12490,N_12198,N_12340);
nor U12491 (N_12491,N_12202,N_12152);
or U12492 (N_12492,N_12114,N_12080);
or U12493 (N_12493,N_12312,N_12172);
or U12494 (N_12494,N_12308,N_12231);
nor U12495 (N_12495,N_12310,N_12061);
nor U12496 (N_12496,N_12130,N_12193);
and U12497 (N_12497,N_12385,N_12044);
nor U12498 (N_12498,N_12070,N_12038);
nor U12499 (N_12499,N_12346,N_12287);
xnor U12500 (N_12500,N_12142,N_12307);
or U12501 (N_12501,N_12240,N_12123);
xor U12502 (N_12502,N_12261,N_12124);
nor U12503 (N_12503,N_12272,N_12359);
or U12504 (N_12504,N_12010,N_12369);
nand U12505 (N_12505,N_12253,N_12357);
xor U12506 (N_12506,N_12247,N_12083);
nor U12507 (N_12507,N_12036,N_12099);
or U12508 (N_12508,N_12344,N_12336);
or U12509 (N_12509,N_12347,N_12204);
nor U12510 (N_12510,N_12025,N_12331);
nand U12511 (N_12511,N_12322,N_12095);
or U12512 (N_12512,N_12108,N_12016);
xor U12513 (N_12513,N_12370,N_12245);
nand U12514 (N_12514,N_12023,N_12163);
or U12515 (N_12515,N_12267,N_12329);
xor U12516 (N_12516,N_12040,N_12244);
xnor U12517 (N_12517,N_12030,N_12270);
and U12518 (N_12518,N_12275,N_12057);
nor U12519 (N_12519,N_12356,N_12268);
nor U12520 (N_12520,N_12278,N_12208);
and U12521 (N_12521,N_12334,N_12031);
nand U12522 (N_12522,N_12389,N_12388);
xnor U12523 (N_12523,N_12047,N_12248);
nand U12524 (N_12524,N_12224,N_12098);
and U12525 (N_12525,N_12390,N_12314);
nor U12526 (N_12526,N_12100,N_12255);
and U12527 (N_12527,N_12012,N_12145);
nor U12528 (N_12528,N_12174,N_12073);
and U12529 (N_12529,N_12396,N_12325);
or U12530 (N_12530,N_12005,N_12398);
xnor U12531 (N_12531,N_12293,N_12225);
xnor U12532 (N_12532,N_12134,N_12156);
nand U12533 (N_12533,N_12294,N_12317);
and U12534 (N_12534,N_12277,N_12089);
nor U12535 (N_12535,N_12051,N_12092);
and U12536 (N_12536,N_12379,N_12229);
or U12537 (N_12537,N_12355,N_12378);
nand U12538 (N_12538,N_12039,N_12258);
nand U12539 (N_12539,N_12218,N_12161);
nand U12540 (N_12540,N_12158,N_12297);
and U12541 (N_12541,N_12326,N_12054);
nor U12542 (N_12542,N_12210,N_12330);
or U12543 (N_12543,N_12377,N_12135);
or U12544 (N_12544,N_12236,N_12241);
nor U12545 (N_12545,N_12033,N_12043);
xor U12546 (N_12546,N_12313,N_12327);
xor U12547 (N_12547,N_12131,N_12228);
xnor U12548 (N_12548,N_12292,N_12203);
nor U12549 (N_12549,N_12337,N_12221);
xnor U12550 (N_12550,N_12260,N_12062);
or U12551 (N_12551,N_12067,N_12222);
or U12552 (N_12552,N_12250,N_12342);
or U12553 (N_12553,N_12109,N_12015);
nor U12554 (N_12554,N_12302,N_12232);
nand U12555 (N_12555,N_12079,N_12165);
and U12556 (N_12556,N_12348,N_12350);
nand U12557 (N_12557,N_12235,N_12269);
and U12558 (N_12558,N_12021,N_12144);
and U12559 (N_12559,N_12375,N_12373);
nor U12560 (N_12560,N_12116,N_12128);
nor U12561 (N_12561,N_12368,N_12353);
and U12562 (N_12562,N_12372,N_12094);
or U12563 (N_12563,N_12159,N_12071);
nor U12564 (N_12564,N_12074,N_12058);
nor U12565 (N_12565,N_12364,N_12042);
xnor U12566 (N_12566,N_12201,N_12000);
or U12567 (N_12567,N_12189,N_12102);
and U12568 (N_12568,N_12183,N_12387);
or U12569 (N_12569,N_12216,N_12110);
xnor U12570 (N_12570,N_12065,N_12286);
nand U12571 (N_12571,N_12147,N_12024);
xor U12572 (N_12572,N_12304,N_12324);
and U12573 (N_12573,N_12186,N_12035);
xor U12574 (N_12574,N_12082,N_12177);
and U12575 (N_12575,N_12048,N_12173);
nor U12576 (N_12576,N_12085,N_12227);
nor U12577 (N_12577,N_12288,N_12343);
nand U12578 (N_12578,N_12243,N_12119);
or U12579 (N_12579,N_12196,N_12188);
and U12580 (N_12580,N_12199,N_12170);
nand U12581 (N_12581,N_12187,N_12223);
nor U12582 (N_12582,N_12113,N_12003);
nand U12583 (N_12583,N_12380,N_12055);
nor U12584 (N_12584,N_12121,N_12064);
nor U12585 (N_12585,N_12162,N_12060);
nand U12586 (N_12586,N_12321,N_12138);
nor U12587 (N_12587,N_12176,N_12381);
and U12588 (N_12588,N_12217,N_12008);
and U12589 (N_12589,N_12363,N_12316);
and U12590 (N_12590,N_12338,N_12146);
nor U12591 (N_12591,N_12122,N_12365);
nor U12592 (N_12592,N_12112,N_12126);
nand U12593 (N_12593,N_12215,N_12076);
nand U12594 (N_12594,N_12266,N_12182);
xor U12595 (N_12595,N_12295,N_12274);
and U12596 (N_12596,N_12242,N_12029);
nand U12597 (N_12597,N_12237,N_12115);
or U12598 (N_12598,N_12283,N_12041);
or U12599 (N_12599,N_12118,N_12254);
or U12600 (N_12600,N_12255,N_12054);
or U12601 (N_12601,N_12238,N_12094);
xnor U12602 (N_12602,N_12340,N_12333);
and U12603 (N_12603,N_12346,N_12003);
nand U12604 (N_12604,N_12318,N_12075);
or U12605 (N_12605,N_12384,N_12324);
or U12606 (N_12606,N_12252,N_12270);
and U12607 (N_12607,N_12330,N_12067);
and U12608 (N_12608,N_12151,N_12320);
nor U12609 (N_12609,N_12066,N_12315);
xor U12610 (N_12610,N_12376,N_12227);
xnor U12611 (N_12611,N_12102,N_12344);
or U12612 (N_12612,N_12252,N_12327);
or U12613 (N_12613,N_12088,N_12082);
and U12614 (N_12614,N_12207,N_12391);
nor U12615 (N_12615,N_12126,N_12141);
or U12616 (N_12616,N_12334,N_12160);
nand U12617 (N_12617,N_12297,N_12354);
xor U12618 (N_12618,N_12021,N_12315);
nor U12619 (N_12619,N_12171,N_12226);
nor U12620 (N_12620,N_12202,N_12174);
nand U12621 (N_12621,N_12201,N_12348);
and U12622 (N_12622,N_12238,N_12127);
and U12623 (N_12623,N_12257,N_12205);
and U12624 (N_12624,N_12064,N_12270);
nand U12625 (N_12625,N_12190,N_12134);
nand U12626 (N_12626,N_12011,N_12093);
nor U12627 (N_12627,N_12098,N_12203);
nand U12628 (N_12628,N_12210,N_12088);
nor U12629 (N_12629,N_12064,N_12198);
nor U12630 (N_12630,N_12092,N_12373);
and U12631 (N_12631,N_12354,N_12221);
nor U12632 (N_12632,N_12272,N_12389);
and U12633 (N_12633,N_12166,N_12254);
nor U12634 (N_12634,N_12146,N_12151);
nand U12635 (N_12635,N_12236,N_12196);
nor U12636 (N_12636,N_12294,N_12184);
nor U12637 (N_12637,N_12376,N_12389);
xor U12638 (N_12638,N_12196,N_12292);
xor U12639 (N_12639,N_12150,N_12398);
nor U12640 (N_12640,N_12104,N_12056);
and U12641 (N_12641,N_12299,N_12275);
xor U12642 (N_12642,N_12136,N_12227);
nor U12643 (N_12643,N_12393,N_12140);
nor U12644 (N_12644,N_12271,N_12342);
or U12645 (N_12645,N_12034,N_12066);
and U12646 (N_12646,N_12210,N_12227);
and U12647 (N_12647,N_12100,N_12080);
nand U12648 (N_12648,N_12288,N_12013);
nor U12649 (N_12649,N_12178,N_12211);
nor U12650 (N_12650,N_12237,N_12396);
and U12651 (N_12651,N_12329,N_12178);
nand U12652 (N_12652,N_12261,N_12366);
nand U12653 (N_12653,N_12384,N_12320);
xnor U12654 (N_12654,N_12038,N_12010);
and U12655 (N_12655,N_12386,N_12331);
and U12656 (N_12656,N_12133,N_12275);
nor U12657 (N_12657,N_12123,N_12211);
and U12658 (N_12658,N_12155,N_12225);
or U12659 (N_12659,N_12304,N_12157);
and U12660 (N_12660,N_12148,N_12194);
or U12661 (N_12661,N_12180,N_12177);
or U12662 (N_12662,N_12250,N_12229);
nand U12663 (N_12663,N_12165,N_12144);
nand U12664 (N_12664,N_12257,N_12334);
or U12665 (N_12665,N_12199,N_12014);
xnor U12666 (N_12666,N_12044,N_12386);
and U12667 (N_12667,N_12192,N_12134);
or U12668 (N_12668,N_12069,N_12112);
nor U12669 (N_12669,N_12278,N_12002);
xor U12670 (N_12670,N_12297,N_12194);
and U12671 (N_12671,N_12375,N_12134);
nor U12672 (N_12672,N_12372,N_12263);
or U12673 (N_12673,N_12210,N_12058);
and U12674 (N_12674,N_12004,N_12376);
nor U12675 (N_12675,N_12090,N_12282);
xor U12676 (N_12676,N_12170,N_12397);
nand U12677 (N_12677,N_12251,N_12103);
nor U12678 (N_12678,N_12059,N_12068);
or U12679 (N_12679,N_12205,N_12211);
nand U12680 (N_12680,N_12005,N_12190);
xnor U12681 (N_12681,N_12289,N_12205);
nor U12682 (N_12682,N_12224,N_12069);
nand U12683 (N_12683,N_12254,N_12072);
and U12684 (N_12684,N_12034,N_12240);
xnor U12685 (N_12685,N_12135,N_12384);
or U12686 (N_12686,N_12196,N_12087);
nor U12687 (N_12687,N_12021,N_12339);
or U12688 (N_12688,N_12398,N_12072);
and U12689 (N_12689,N_12195,N_12082);
and U12690 (N_12690,N_12209,N_12204);
or U12691 (N_12691,N_12217,N_12262);
or U12692 (N_12692,N_12039,N_12357);
or U12693 (N_12693,N_12232,N_12172);
xor U12694 (N_12694,N_12051,N_12121);
xor U12695 (N_12695,N_12139,N_12036);
xnor U12696 (N_12696,N_12330,N_12103);
xnor U12697 (N_12697,N_12375,N_12361);
and U12698 (N_12698,N_12186,N_12367);
xor U12699 (N_12699,N_12310,N_12297);
or U12700 (N_12700,N_12370,N_12082);
or U12701 (N_12701,N_12140,N_12286);
and U12702 (N_12702,N_12356,N_12172);
xor U12703 (N_12703,N_12197,N_12346);
xor U12704 (N_12704,N_12092,N_12090);
nand U12705 (N_12705,N_12160,N_12035);
xor U12706 (N_12706,N_12327,N_12259);
xor U12707 (N_12707,N_12097,N_12369);
nand U12708 (N_12708,N_12066,N_12139);
xor U12709 (N_12709,N_12012,N_12231);
nor U12710 (N_12710,N_12184,N_12292);
or U12711 (N_12711,N_12085,N_12321);
nor U12712 (N_12712,N_12288,N_12319);
and U12713 (N_12713,N_12290,N_12299);
nand U12714 (N_12714,N_12236,N_12269);
or U12715 (N_12715,N_12132,N_12094);
or U12716 (N_12716,N_12371,N_12247);
or U12717 (N_12717,N_12257,N_12232);
and U12718 (N_12718,N_12295,N_12376);
xnor U12719 (N_12719,N_12025,N_12265);
xor U12720 (N_12720,N_12347,N_12337);
nand U12721 (N_12721,N_12226,N_12054);
and U12722 (N_12722,N_12008,N_12035);
nand U12723 (N_12723,N_12359,N_12268);
and U12724 (N_12724,N_12114,N_12222);
and U12725 (N_12725,N_12106,N_12171);
and U12726 (N_12726,N_12329,N_12125);
and U12727 (N_12727,N_12107,N_12019);
nand U12728 (N_12728,N_12298,N_12082);
nor U12729 (N_12729,N_12021,N_12205);
and U12730 (N_12730,N_12005,N_12324);
nand U12731 (N_12731,N_12355,N_12319);
nor U12732 (N_12732,N_12142,N_12007);
nand U12733 (N_12733,N_12080,N_12250);
and U12734 (N_12734,N_12192,N_12093);
xor U12735 (N_12735,N_12171,N_12068);
xor U12736 (N_12736,N_12134,N_12330);
and U12737 (N_12737,N_12381,N_12345);
or U12738 (N_12738,N_12062,N_12203);
nor U12739 (N_12739,N_12015,N_12389);
xnor U12740 (N_12740,N_12346,N_12068);
and U12741 (N_12741,N_12076,N_12294);
nand U12742 (N_12742,N_12135,N_12383);
nand U12743 (N_12743,N_12265,N_12134);
or U12744 (N_12744,N_12168,N_12397);
nand U12745 (N_12745,N_12304,N_12109);
and U12746 (N_12746,N_12229,N_12274);
nor U12747 (N_12747,N_12325,N_12088);
and U12748 (N_12748,N_12049,N_12201);
nand U12749 (N_12749,N_12195,N_12066);
nand U12750 (N_12750,N_12071,N_12042);
xnor U12751 (N_12751,N_12254,N_12131);
and U12752 (N_12752,N_12304,N_12377);
nand U12753 (N_12753,N_12179,N_12256);
or U12754 (N_12754,N_12141,N_12064);
and U12755 (N_12755,N_12051,N_12351);
nand U12756 (N_12756,N_12255,N_12043);
nor U12757 (N_12757,N_12038,N_12189);
or U12758 (N_12758,N_12181,N_12389);
and U12759 (N_12759,N_12370,N_12356);
and U12760 (N_12760,N_12077,N_12264);
or U12761 (N_12761,N_12273,N_12054);
xor U12762 (N_12762,N_12388,N_12357);
nor U12763 (N_12763,N_12294,N_12052);
or U12764 (N_12764,N_12004,N_12354);
nor U12765 (N_12765,N_12258,N_12204);
nor U12766 (N_12766,N_12305,N_12073);
or U12767 (N_12767,N_12328,N_12287);
or U12768 (N_12768,N_12277,N_12265);
nor U12769 (N_12769,N_12125,N_12126);
or U12770 (N_12770,N_12028,N_12004);
nand U12771 (N_12771,N_12045,N_12256);
xnor U12772 (N_12772,N_12316,N_12214);
nor U12773 (N_12773,N_12321,N_12364);
nand U12774 (N_12774,N_12084,N_12246);
or U12775 (N_12775,N_12394,N_12051);
and U12776 (N_12776,N_12034,N_12394);
xor U12777 (N_12777,N_12361,N_12058);
xor U12778 (N_12778,N_12089,N_12081);
nor U12779 (N_12779,N_12246,N_12313);
or U12780 (N_12780,N_12259,N_12110);
nor U12781 (N_12781,N_12209,N_12053);
or U12782 (N_12782,N_12235,N_12283);
xnor U12783 (N_12783,N_12244,N_12339);
xor U12784 (N_12784,N_12355,N_12332);
xnor U12785 (N_12785,N_12366,N_12249);
nand U12786 (N_12786,N_12015,N_12128);
or U12787 (N_12787,N_12201,N_12340);
xnor U12788 (N_12788,N_12263,N_12021);
nor U12789 (N_12789,N_12011,N_12004);
nand U12790 (N_12790,N_12032,N_12147);
nor U12791 (N_12791,N_12255,N_12119);
nand U12792 (N_12792,N_12349,N_12005);
and U12793 (N_12793,N_12338,N_12093);
xnor U12794 (N_12794,N_12300,N_12033);
or U12795 (N_12795,N_12313,N_12136);
nor U12796 (N_12796,N_12299,N_12239);
nand U12797 (N_12797,N_12339,N_12202);
nand U12798 (N_12798,N_12117,N_12100);
nor U12799 (N_12799,N_12126,N_12271);
nor U12800 (N_12800,N_12629,N_12434);
and U12801 (N_12801,N_12491,N_12615);
or U12802 (N_12802,N_12633,N_12649);
xor U12803 (N_12803,N_12581,N_12521);
nor U12804 (N_12804,N_12774,N_12550);
and U12805 (N_12805,N_12788,N_12561);
and U12806 (N_12806,N_12791,N_12576);
xor U12807 (N_12807,N_12780,N_12664);
or U12808 (N_12808,N_12598,N_12738);
nand U12809 (N_12809,N_12622,N_12586);
or U12810 (N_12810,N_12772,N_12400);
xnor U12811 (N_12811,N_12642,N_12674);
xnor U12812 (N_12812,N_12530,N_12404);
nor U12813 (N_12813,N_12405,N_12556);
nor U12814 (N_12814,N_12459,N_12786);
nor U12815 (N_12815,N_12636,N_12527);
or U12816 (N_12816,N_12518,N_12720);
and U12817 (N_12817,N_12677,N_12456);
or U12818 (N_12818,N_12511,N_12490);
and U12819 (N_12819,N_12476,N_12416);
xor U12820 (N_12820,N_12452,N_12638);
xnor U12821 (N_12821,N_12525,N_12510);
or U12822 (N_12822,N_12486,N_12641);
nor U12823 (N_12823,N_12568,N_12450);
or U12824 (N_12824,N_12625,N_12709);
xor U12825 (N_12825,N_12706,N_12468);
nand U12826 (N_12826,N_12637,N_12538);
xor U12827 (N_12827,N_12604,N_12483);
nor U12828 (N_12828,N_12733,N_12719);
and U12829 (N_12829,N_12554,N_12793);
nand U12830 (N_12830,N_12451,N_12515);
and U12831 (N_12831,N_12635,N_12699);
xor U12832 (N_12832,N_12500,N_12467);
and U12833 (N_12833,N_12749,N_12696);
nor U12834 (N_12834,N_12574,N_12703);
nor U12835 (N_12835,N_12670,N_12667);
or U12836 (N_12836,N_12614,N_12705);
xor U12837 (N_12837,N_12631,N_12446);
xor U12838 (N_12838,N_12689,N_12588);
nand U12839 (N_12839,N_12746,N_12445);
nand U12840 (N_12840,N_12471,N_12630);
or U12841 (N_12841,N_12579,N_12401);
nor U12842 (N_12842,N_12756,N_12424);
or U12843 (N_12843,N_12547,N_12544);
nand U12844 (N_12844,N_12707,N_12484);
or U12845 (N_12845,N_12532,N_12799);
or U12846 (N_12846,N_12741,N_12565);
xor U12847 (N_12847,N_12708,N_12564);
nor U12848 (N_12848,N_12455,N_12443);
xor U12849 (N_12849,N_12536,N_12758);
xor U12850 (N_12850,N_12632,N_12702);
nand U12851 (N_12851,N_12448,N_12432);
and U12852 (N_12852,N_12698,N_12528);
nand U12853 (N_12853,N_12453,N_12747);
nand U12854 (N_12854,N_12652,N_12744);
nand U12855 (N_12855,N_12423,N_12678);
and U12856 (N_12856,N_12470,N_12514);
and U12857 (N_12857,N_12519,N_12558);
nor U12858 (N_12858,N_12686,N_12714);
nand U12859 (N_12859,N_12690,N_12534);
nand U12860 (N_12860,N_12684,N_12628);
nand U12861 (N_12861,N_12675,N_12792);
or U12862 (N_12862,N_12508,N_12728);
or U12863 (N_12863,N_12639,N_12506);
xor U12864 (N_12864,N_12543,N_12771);
nor U12865 (N_12865,N_12559,N_12757);
xor U12866 (N_12866,N_12605,N_12769);
nand U12867 (N_12867,N_12603,N_12753);
or U12868 (N_12868,N_12697,N_12512);
xor U12869 (N_12869,N_12711,N_12612);
and U12870 (N_12870,N_12685,N_12634);
or U12871 (N_12871,N_12415,N_12593);
xnor U12872 (N_12872,N_12402,N_12503);
and U12873 (N_12873,N_12431,N_12553);
and U12874 (N_12874,N_12575,N_12736);
nand U12875 (N_12875,N_12752,N_12537);
xnor U12876 (N_12876,N_12425,N_12761);
xor U12877 (N_12877,N_12681,N_12555);
and U12878 (N_12878,N_12712,N_12516);
or U12879 (N_12879,N_12726,N_12414);
and U12880 (N_12880,N_12762,N_12782);
and U12881 (N_12881,N_12611,N_12737);
xor U12882 (N_12882,N_12407,N_12669);
and U12883 (N_12883,N_12488,N_12481);
xnor U12884 (N_12884,N_12551,N_12716);
nor U12885 (N_12885,N_12600,N_12648);
nand U12886 (N_12886,N_12489,N_12729);
or U12887 (N_12887,N_12610,N_12499);
xor U12888 (N_12888,N_12722,N_12410);
or U12889 (N_12889,N_12591,N_12509);
nand U12890 (N_12890,N_12496,N_12766);
nand U12891 (N_12891,N_12778,N_12659);
nor U12892 (N_12892,N_12745,N_12580);
nand U12893 (N_12893,N_12645,N_12540);
or U12894 (N_12894,N_12430,N_12742);
and U12895 (N_12895,N_12570,N_12692);
xnor U12896 (N_12896,N_12563,N_12607);
nor U12897 (N_12897,N_12571,N_12683);
xnor U12898 (N_12898,N_12764,N_12535);
or U12899 (N_12899,N_12671,N_12673);
nor U12900 (N_12900,N_12640,N_12524);
and U12901 (N_12901,N_12582,N_12644);
nor U12902 (N_12902,N_12461,N_12546);
nand U12903 (N_12903,N_12545,N_12495);
xnor U12904 (N_12904,N_12734,N_12623);
and U12905 (N_12905,N_12613,N_12449);
nand U12906 (N_12906,N_12473,N_12701);
xor U12907 (N_12907,N_12679,N_12584);
and U12908 (N_12908,N_12754,N_12650);
and U12909 (N_12909,N_12501,N_12609);
nor U12910 (N_12910,N_12763,N_12447);
or U12911 (N_12911,N_12616,N_12457);
nor U12912 (N_12912,N_12784,N_12651);
xor U12913 (N_12913,N_12783,N_12666);
and U12914 (N_12914,N_12672,N_12776);
and U12915 (N_12915,N_12662,N_12731);
xnor U12916 (N_12916,N_12479,N_12743);
nor U12917 (N_12917,N_12596,N_12420);
xor U12918 (N_12918,N_12520,N_12492);
and U12919 (N_12919,N_12658,N_12715);
nor U12920 (N_12920,N_12522,N_12700);
xor U12921 (N_12921,N_12413,N_12750);
or U12922 (N_12922,N_12539,N_12748);
nor U12923 (N_12923,N_12428,N_12688);
nor U12924 (N_12924,N_12441,N_12533);
or U12925 (N_12925,N_12718,N_12621);
or U12926 (N_12926,N_12403,N_12597);
or U12927 (N_12927,N_12436,N_12665);
and U12928 (N_12928,N_12721,N_12724);
or U12929 (N_12929,N_12421,N_12668);
xnor U12930 (N_12930,N_12465,N_12437);
or U12931 (N_12931,N_12760,N_12504);
nor U12932 (N_12932,N_12606,N_12680);
nor U12933 (N_12933,N_12573,N_12713);
or U12934 (N_12934,N_12517,N_12777);
nor U12935 (N_12935,N_12795,N_12740);
nor U12936 (N_12936,N_12485,N_12735);
nand U12937 (N_12937,N_12592,N_12676);
nor U12938 (N_12938,N_12695,N_12585);
nand U12939 (N_12939,N_12482,N_12765);
and U12940 (N_12940,N_12493,N_12464);
xor U12941 (N_12941,N_12694,N_12643);
xor U12942 (N_12942,N_12458,N_12557);
xor U12943 (N_12943,N_12727,N_12566);
or U12944 (N_12944,N_12595,N_12572);
xor U12945 (N_12945,N_12656,N_12653);
or U12946 (N_12946,N_12442,N_12549);
and U12947 (N_12947,N_12438,N_12704);
xor U12948 (N_12948,N_12419,N_12460);
or U12949 (N_12949,N_12767,N_12779);
or U12950 (N_12950,N_12477,N_12626);
nand U12951 (N_12951,N_12412,N_12755);
nand U12952 (N_12952,N_12560,N_12472);
nand U12953 (N_12953,N_12406,N_12768);
and U12954 (N_12954,N_12601,N_12478);
or U12955 (N_12955,N_12682,N_12411);
or U12956 (N_12956,N_12751,N_12710);
nand U12957 (N_12957,N_12624,N_12647);
and U12958 (N_12958,N_12583,N_12787);
nand U12959 (N_12959,N_12739,N_12732);
nand U12960 (N_12960,N_12569,N_12790);
nand U12961 (N_12961,N_12440,N_12594);
xnor U12962 (N_12962,N_12589,N_12498);
or U12963 (N_12963,N_12627,N_12620);
or U12964 (N_12964,N_12418,N_12660);
or U12965 (N_12965,N_12505,N_12548);
nor U12966 (N_12966,N_12531,N_12439);
and U12967 (N_12967,N_12608,N_12454);
xnor U12968 (N_12968,N_12599,N_12789);
xnor U12969 (N_12969,N_12759,N_12513);
xor U12970 (N_12970,N_12542,N_12463);
or U12971 (N_12971,N_12427,N_12433);
and U12972 (N_12972,N_12444,N_12429);
nor U12973 (N_12973,N_12494,N_12497);
and U12974 (N_12974,N_12661,N_12435);
nor U12975 (N_12975,N_12618,N_12469);
xor U12976 (N_12976,N_12785,N_12691);
xor U12977 (N_12977,N_12693,N_12462);
nor U12978 (N_12978,N_12552,N_12480);
nand U12979 (N_12979,N_12798,N_12562);
and U12980 (N_12980,N_12602,N_12529);
nand U12981 (N_12981,N_12409,N_12663);
nand U12982 (N_12982,N_12770,N_12773);
xnor U12983 (N_12983,N_12567,N_12541);
nand U12984 (N_12984,N_12590,N_12655);
nor U12985 (N_12985,N_12723,N_12426);
nand U12986 (N_12986,N_12687,N_12408);
and U12987 (N_12987,N_12502,N_12781);
nand U12988 (N_12988,N_12794,N_12507);
xnor U12989 (N_12989,N_12466,N_12619);
or U12990 (N_12990,N_12417,N_12617);
nor U12991 (N_12991,N_12577,N_12796);
xnor U12992 (N_12992,N_12422,N_12526);
xnor U12993 (N_12993,N_12587,N_12475);
or U12994 (N_12994,N_12725,N_12657);
nand U12995 (N_12995,N_12487,N_12797);
nand U12996 (N_12996,N_12654,N_12646);
or U12997 (N_12997,N_12775,N_12578);
nor U12998 (N_12998,N_12717,N_12730);
nand U12999 (N_12999,N_12523,N_12474);
or U13000 (N_13000,N_12525,N_12504);
nand U13001 (N_13001,N_12733,N_12693);
nor U13002 (N_13002,N_12652,N_12723);
xor U13003 (N_13003,N_12468,N_12512);
xor U13004 (N_13004,N_12761,N_12430);
nand U13005 (N_13005,N_12519,N_12571);
xnor U13006 (N_13006,N_12634,N_12466);
nand U13007 (N_13007,N_12558,N_12646);
xor U13008 (N_13008,N_12654,N_12585);
nor U13009 (N_13009,N_12524,N_12680);
xor U13010 (N_13010,N_12643,N_12732);
or U13011 (N_13011,N_12425,N_12510);
nand U13012 (N_13012,N_12680,N_12684);
nor U13013 (N_13013,N_12578,N_12568);
nand U13014 (N_13014,N_12477,N_12649);
xor U13015 (N_13015,N_12588,N_12462);
nand U13016 (N_13016,N_12726,N_12710);
nor U13017 (N_13017,N_12776,N_12646);
or U13018 (N_13018,N_12582,N_12565);
xnor U13019 (N_13019,N_12696,N_12796);
and U13020 (N_13020,N_12598,N_12704);
nor U13021 (N_13021,N_12479,N_12650);
nand U13022 (N_13022,N_12556,N_12430);
nor U13023 (N_13023,N_12749,N_12572);
or U13024 (N_13024,N_12742,N_12682);
nor U13025 (N_13025,N_12649,N_12514);
nor U13026 (N_13026,N_12754,N_12452);
nand U13027 (N_13027,N_12431,N_12779);
and U13028 (N_13028,N_12496,N_12400);
xor U13029 (N_13029,N_12609,N_12446);
nand U13030 (N_13030,N_12476,N_12540);
nand U13031 (N_13031,N_12675,N_12411);
and U13032 (N_13032,N_12624,N_12606);
or U13033 (N_13033,N_12430,N_12617);
and U13034 (N_13034,N_12630,N_12611);
or U13035 (N_13035,N_12518,N_12639);
xor U13036 (N_13036,N_12469,N_12595);
nor U13037 (N_13037,N_12786,N_12522);
nand U13038 (N_13038,N_12471,N_12733);
nand U13039 (N_13039,N_12534,N_12496);
or U13040 (N_13040,N_12618,N_12626);
nor U13041 (N_13041,N_12512,N_12744);
xor U13042 (N_13042,N_12790,N_12416);
xnor U13043 (N_13043,N_12793,N_12705);
nor U13044 (N_13044,N_12401,N_12446);
xnor U13045 (N_13045,N_12758,N_12643);
and U13046 (N_13046,N_12768,N_12403);
and U13047 (N_13047,N_12447,N_12685);
or U13048 (N_13048,N_12473,N_12695);
nor U13049 (N_13049,N_12456,N_12602);
xnor U13050 (N_13050,N_12552,N_12721);
xor U13051 (N_13051,N_12442,N_12425);
xnor U13052 (N_13052,N_12796,N_12710);
or U13053 (N_13053,N_12737,N_12491);
or U13054 (N_13054,N_12643,N_12406);
xnor U13055 (N_13055,N_12720,N_12512);
xnor U13056 (N_13056,N_12656,N_12724);
and U13057 (N_13057,N_12443,N_12572);
or U13058 (N_13058,N_12611,N_12756);
xnor U13059 (N_13059,N_12543,N_12548);
xor U13060 (N_13060,N_12465,N_12752);
nor U13061 (N_13061,N_12509,N_12537);
and U13062 (N_13062,N_12655,N_12716);
and U13063 (N_13063,N_12790,N_12702);
nand U13064 (N_13064,N_12656,N_12567);
nor U13065 (N_13065,N_12737,N_12695);
nor U13066 (N_13066,N_12771,N_12718);
or U13067 (N_13067,N_12490,N_12528);
or U13068 (N_13068,N_12400,N_12553);
or U13069 (N_13069,N_12734,N_12652);
and U13070 (N_13070,N_12492,N_12793);
and U13071 (N_13071,N_12402,N_12448);
or U13072 (N_13072,N_12517,N_12533);
xnor U13073 (N_13073,N_12581,N_12441);
nand U13074 (N_13074,N_12541,N_12627);
nor U13075 (N_13075,N_12668,N_12509);
nor U13076 (N_13076,N_12721,N_12472);
nor U13077 (N_13077,N_12431,N_12767);
nor U13078 (N_13078,N_12469,N_12565);
nand U13079 (N_13079,N_12502,N_12518);
nor U13080 (N_13080,N_12613,N_12770);
nor U13081 (N_13081,N_12573,N_12492);
or U13082 (N_13082,N_12621,N_12679);
nand U13083 (N_13083,N_12575,N_12527);
and U13084 (N_13084,N_12699,N_12576);
nor U13085 (N_13085,N_12769,N_12410);
xor U13086 (N_13086,N_12433,N_12562);
nand U13087 (N_13087,N_12505,N_12588);
or U13088 (N_13088,N_12765,N_12508);
nor U13089 (N_13089,N_12591,N_12779);
nor U13090 (N_13090,N_12768,N_12611);
xor U13091 (N_13091,N_12695,N_12625);
nand U13092 (N_13092,N_12729,N_12410);
nor U13093 (N_13093,N_12465,N_12532);
nand U13094 (N_13094,N_12587,N_12787);
or U13095 (N_13095,N_12401,N_12626);
or U13096 (N_13096,N_12706,N_12429);
nand U13097 (N_13097,N_12431,N_12698);
nand U13098 (N_13098,N_12568,N_12455);
nor U13099 (N_13099,N_12567,N_12481);
xor U13100 (N_13100,N_12505,N_12457);
and U13101 (N_13101,N_12540,N_12496);
xor U13102 (N_13102,N_12472,N_12444);
and U13103 (N_13103,N_12447,N_12479);
nand U13104 (N_13104,N_12713,N_12553);
nand U13105 (N_13105,N_12550,N_12495);
xor U13106 (N_13106,N_12649,N_12493);
nand U13107 (N_13107,N_12621,N_12746);
or U13108 (N_13108,N_12627,N_12622);
nand U13109 (N_13109,N_12741,N_12633);
and U13110 (N_13110,N_12459,N_12418);
or U13111 (N_13111,N_12499,N_12734);
nand U13112 (N_13112,N_12699,N_12459);
nand U13113 (N_13113,N_12485,N_12539);
or U13114 (N_13114,N_12748,N_12426);
nor U13115 (N_13115,N_12760,N_12679);
nand U13116 (N_13116,N_12775,N_12687);
nor U13117 (N_13117,N_12544,N_12755);
or U13118 (N_13118,N_12744,N_12618);
or U13119 (N_13119,N_12445,N_12529);
xor U13120 (N_13120,N_12719,N_12670);
nand U13121 (N_13121,N_12708,N_12670);
and U13122 (N_13122,N_12640,N_12566);
or U13123 (N_13123,N_12514,N_12463);
nor U13124 (N_13124,N_12640,N_12495);
nor U13125 (N_13125,N_12601,N_12646);
and U13126 (N_13126,N_12597,N_12719);
nand U13127 (N_13127,N_12669,N_12413);
and U13128 (N_13128,N_12779,N_12651);
xnor U13129 (N_13129,N_12583,N_12509);
nand U13130 (N_13130,N_12401,N_12419);
or U13131 (N_13131,N_12576,N_12782);
nand U13132 (N_13132,N_12548,N_12704);
nand U13133 (N_13133,N_12625,N_12790);
nor U13134 (N_13134,N_12532,N_12615);
nor U13135 (N_13135,N_12466,N_12408);
nand U13136 (N_13136,N_12563,N_12455);
nor U13137 (N_13137,N_12672,N_12443);
xnor U13138 (N_13138,N_12748,N_12752);
or U13139 (N_13139,N_12470,N_12761);
and U13140 (N_13140,N_12737,N_12705);
and U13141 (N_13141,N_12682,N_12614);
nand U13142 (N_13142,N_12443,N_12775);
and U13143 (N_13143,N_12788,N_12424);
and U13144 (N_13144,N_12675,N_12666);
xor U13145 (N_13145,N_12767,N_12652);
nor U13146 (N_13146,N_12539,N_12776);
nand U13147 (N_13147,N_12514,N_12430);
and U13148 (N_13148,N_12583,N_12794);
nor U13149 (N_13149,N_12701,N_12560);
and U13150 (N_13150,N_12557,N_12463);
nand U13151 (N_13151,N_12552,N_12694);
nand U13152 (N_13152,N_12656,N_12577);
nor U13153 (N_13153,N_12401,N_12664);
or U13154 (N_13154,N_12731,N_12776);
nand U13155 (N_13155,N_12744,N_12510);
nor U13156 (N_13156,N_12793,N_12602);
nor U13157 (N_13157,N_12678,N_12644);
and U13158 (N_13158,N_12756,N_12552);
and U13159 (N_13159,N_12528,N_12630);
nand U13160 (N_13160,N_12787,N_12435);
xnor U13161 (N_13161,N_12665,N_12557);
nand U13162 (N_13162,N_12432,N_12403);
nand U13163 (N_13163,N_12557,N_12544);
nand U13164 (N_13164,N_12449,N_12707);
nand U13165 (N_13165,N_12760,N_12603);
and U13166 (N_13166,N_12476,N_12583);
nor U13167 (N_13167,N_12552,N_12453);
xor U13168 (N_13168,N_12799,N_12652);
xor U13169 (N_13169,N_12560,N_12468);
nor U13170 (N_13170,N_12491,N_12766);
and U13171 (N_13171,N_12629,N_12475);
nand U13172 (N_13172,N_12655,N_12745);
nand U13173 (N_13173,N_12743,N_12475);
nand U13174 (N_13174,N_12406,N_12458);
and U13175 (N_13175,N_12432,N_12774);
nand U13176 (N_13176,N_12707,N_12593);
or U13177 (N_13177,N_12471,N_12734);
xnor U13178 (N_13178,N_12561,N_12405);
nand U13179 (N_13179,N_12446,N_12710);
and U13180 (N_13180,N_12730,N_12562);
nand U13181 (N_13181,N_12687,N_12427);
xnor U13182 (N_13182,N_12539,N_12484);
nand U13183 (N_13183,N_12759,N_12739);
xnor U13184 (N_13184,N_12421,N_12656);
or U13185 (N_13185,N_12548,N_12754);
nor U13186 (N_13186,N_12677,N_12710);
and U13187 (N_13187,N_12674,N_12662);
and U13188 (N_13188,N_12474,N_12642);
xor U13189 (N_13189,N_12503,N_12788);
or U13190 (N_13190,N_12481,N_12441);
xor U13191 (N_13191,N_12521,N_12402);
or U13192 (N_13192,N_12712,N_12429);
nand U13193 (N_13193,N_12493,N_12754);
nand U13194 (N_13194,N_12705,N_12548);
or U13195 (N_13195,N_12521,N_12461);
or U13196 (N_13196,N_12704,N_12557);
nor U13197 (N_13197,N_12476,N_12537);
and U13198 (N_13198,N_12749,N_12774);
nand U13199 (N_13199,N_12775,N_12639);
and U13200 (N_13200,N_13049,N_13033);
nor U13201 (N_13201,N_13173,N_12991);
nand U13202 (N_13202,N_12818,N_12860);
nor U13203 (N_13203,N_13193,N_13119);
xor U13204 (N_13204,N_12809,N_12983);
nor U13205 (N_13205,N_13011,N_13022);
nor U13206 (N_13206,N_13075,N_12919);
nand U13207 (N_13207,N_12823,N_12902);
or U13208 (N_13208,N_13159,N_12834);
or U13209 (N_13209,N_12802,N_12957);
nor U13210 (N_13210,N_12942,N_13134);
or U13211 (N_13211,N_13186,N_12828);
nor U13212 (N_13212,N_12898,N_12814);
xnor U13213 (N_13213,N_12956,N_12847);
nand U13214 (N_13214,N_12853,N_12900);
and U13215 (N_13215,N_13028,N_13126);
nand U13216 (N_13216,N_12906,N_12967);
xnor U13217 (N_13217,N_13124,N_12855);
and U13218 (N_13218,N_13084,N_13066);
nand U13219 (N_13219,N_13076,N_12970);
nand U13220 (N_13220,N_13184,N_12918);
or U13221 (N_13221,N_13010,N_13194);
or U13222 (N_13222,N_12941,N_13185);
xnor U13223 (N_13223,N_13000,N_12872);
nand U13224 (N_13224,N_12854,N_12892);
nor U13225 (N_13225,N_12954,N_13002);
xor U13226 (N_13226,N_13086,N_12890);
xnor U13227 (N_13227,N_13112,N_13020);
nand U13228 (N_13228,N_12907,N_13074);
or U13229 (N_13229,N_12804,N_12827);
nand U13230 (N_13230,N_13047,N_13019);
and U13231 (N_13231,N_13101,N_12850);
xor U13232 (N_13232,N_12826,N_13069);
nand U13233 (N_13233,N_13068,N_13132);
xnor U13234 (N_13234,N_12899,N_13018);
nand U13235 (N_13235,N_13029,N_12897);
or U13236 (N_13236,N_13183,N_12914);
xnor U13237 (N_13237,N_13139,N_12801);
and U13238 (N_13238,N_12925,N_12840);
xor U13239 (N_13239,N_13156,N_13061);
nand U13240 (N_13240,N_12961,N_12841);
nor U13241 (N_13241,N_13079,N_12868);
xnor U13242 (N_13242,N_13157,N_12927);
and U13243 (N_13243,N_13090,N_12972);
nor U13244 (N_13244,N_13141,N_13099);
xor U13245 (N_13245,N_13016,N_12808);
xor U13246 (N_13246,N_13127,N_13071);
nand U13247 (N_13247,N_13097,N_13012);
or U13248 (N_13248,N_13014,N_13026);
nor U13249 (N_13249,N_12949,N_13095);
or U13250 (N_13250,N_13161,N_13191);
and U13251 (N_13251,N_12843,N_12977);
or U13252 (N_13252,N_13190,N_13067);
or U13253 (N_13253,N_12831,N_13130);
nor U13254 (N_13254,N_12904,N_12930);
and U13255 (N_13255,N_12875,N_12938);
xnor U13256 (N_13256,N_13053,N_12933);
nand U13257 (N_13257,N_13162,N_13180);
and U13258 (N_13258,N_12878,N_12842);
and U13259 (N_13259,N_12939,N_12937);
nor U13260 (N_13260,N_13146,N_13094);
nor U13261 (N_13261,N_13115,N_13058);
or U13262 (N_13262,N_12943,N_12971);
and U13263 (N_13263,N_12856,N_13078);
xnor U13264 (N_13264,N_13158,N_13006);
xnor U13265 (N_13265,N_13017,N_12876);
xor U13266 (N_13266,N_12888,N_12896);
nand U13267 (N_13267,N_12873,N_13135);
xnor U13268 (N_13268,N_12805,N_12978);
xnor U13269 (N_13269,N_13147,N_12921);
nand U13270 (N_13270,N_13103,N_13042);
nand U13271 (N_13271,N_12931,N_13040);
xnor U13272 (N_13272,N_12909,N_13059);
nor U13273 (N_13273,N_12926,N_12946);
xor U13274 (N_13274,N_13060,N_12817);
and U13275 (N_13275,N_13104,N_13154);
and U13276 (N_13276,N_13051,N_12999);
and U13277 (N_13277,N_12845,N_13107);
nor U13278 (N_13278,N_12852,N_12839);
nand U13279 (N_13279,N_12894,N_13063);
and U13280 (N_13280,N_13133,N_12981);
xnor U13281 (N_13281,N_13013,N_12965);
nor U13282 (N_13282,N_13034,N_12849);
or U13283 (N_13283,N_12960,N_12979);
xnor U13284 (N_13284,N_13118,N_13165);
or U13285 (N_13285,N_12889,N_12862);
nand U13286 (N_13286,N_13171,N_12953);
nand U13287 (N_13287,N_13131,N_12822);
and U13288 (N_13288,N_12851,N_13163);
xor U13289 (N_13289,N_12934,N_12833);
and U13290 (N_13290,N_13153,N_13009);
and U13291 (N_13291,N_13187,N_12883);
nor U13292 (N_13292,N_13092,N_12935);
or U13293 (N_13293,N_12969,N_13050);
nor U13294 (N_13294,N_13052,N_12830);
or U13295 (N_13295,N_13121,N_13057);
xor U13296 (N_13296,N_12859,N_13072);
nor U13297 (N_13297,N_13102,N_13054);
nor U13298 (N_13298,N_13081,N_12821);
nand U13299 (N_13299,N_12863,N_12996);
xor U13300 (N_13300,N_12973,N_12998);
nand U13301 (N_13301,N_12858,N_13167);
or U13302 (N_13302,N_13083,N_12824);
xnor U13303 (N_13303,N_12964,N_13148);
xnor U13304 (N_13304,N_12848,N_13164);
or U13305 (N_13305,N_13088,N_12944);
or U13306 (N_13306,N_12932,N_12910);
nand U13307 (N_13307,N_12807,N_12874);
nand U13308 (N_13308,N_13005,N_13003);
xnor U13309 (N_13309,N_13169,N_13070);
nor U13310 (N_13310,N_13176,N_12885);
and U13311 (N_13311,N_13155,N_12915);
or U13312 (N_13312,N_12846,N_12844);
and U13313 (N_13313,N_13109,N_12816);
and U13314 (N_13314,N_12905,N_13144);
or U13315 (N_13315,N_12988,N_13178);
and U13316 (N_13316,N_12908,N_12895);
nand U13317 (N_13317,N_13152,N_13170);
nand U13318 (N_13318,N_12924,N_13143);
nor U13319 (N_13319,N_13041,N_13149);
xnor U13320 (N_13320,N_13142,N_12866);
xnor U13321 (N_13321,N_12997,N_13015);
and U13322 (N_13322,N_12920,N_12810);
and U13323 (N_13323,N_13197,N_13073);
nor U13324 (N_13324,N_12962,N_13023);
and U13325 (N_13325,N_12829,N_12836);
or U13326 (N_13326,N_12832,N_12893);
or U13327 (N_13327,N_12877,N_13113);
nand U13328 (N_13328,N_13001,N_13037);
nand U13329 (N_13329,N_13129,N_13025);
nand U13330 (N_13330,N_13024,N_13048);
nor U13331 (N_13331,N_13043,N_12881);
nand U13332 (N_13332,N_13096,N_13082);
xnor U13333 (N_13333,N_13175,N_13108);
nor U13334 (N_13334,N_12880,N_12975);
xor U13335 (N_13335,N_13065,N_13136);
xor U13336 (N_13336,N_12980,N_13177);
and U13337 (N_13337,N_12948,N_13182);
nand U13338 (N_13338,N_12815,N_13106);
and U13339 (N_13339,N_12994,N_12936);
and U13340 (N_13340,N_13110,N_12985);
or U13341 (N_13341,N_12995,N_12901);
or U13342 (N_13342,N_13098,N_13085);
xor U13343 (N_13343,N_13046,N_12990);
nand U13344 (N_13344,N_12811,N_13122);
nor U13345 (N_13345,N_12928,N_12812);
nor U13346 (N_13346,N_13181,N_12968);
or U13347 (N_13347,N_12813,N_12879);
and U13348 (N_13348,N_12869,N_13140);
and U13349 (N_13349,N_13189,N_12913);
xor U13350 (N_13350,N_13087,N_12864);
xor U13351 (N_13351,N_12835,N_12993);
xnor U13352 (N_13352,N_12922,N_13004);
xnor U13353 (N_13353,N_13100,N_12916);
or U13354 (N_13354,N_12940,N_12803);
xor U13355 (N_13355,N_13116,N_13044);
nand U13356 (N_13356,N_12884,N_12903);
nor U13357 (N_13357,N_13196,N_12912);
xor U13358 (N_13358,N_13123,N_12923);
or U13359 (N_13359,N_13166,N_12992);
nor U13360 (N_13360,N_13093,N_13008);
xor U13361 (N_13361,N_13111,N_13138);
xnor U13362 (N_13362,N_12857,N_12820);
nor U13363 (N_13363,N_12945,N_13091);
nand U13364 (N_13364,N_12986,N_12947);
xor U13365 (N_13365,N_13055,N_12800);
nand U13366 (N_13366,N_13031,N_12887);
nor U13367 (N_13367,N_13195,N_13036);
nor U13368 (N_13368,N_13045,N_13128);
nor U13369 (N_13369,N_12951,N_13089);
and U13370 (N_13370,N_12837,N_12959);
nor U13371 (N_13371,N_12891,N_12952);
nand U13372 (N_13372,N_13032,N_13125);
or U13373 (N_13373,N_13077,N_12819);
nand U13374 (N_13374,N_12870,N_13150);
xor U13375 (N_13375,N_12882,N_13151);
xnor U13376 (N_13376,N_12982,N_12861);
and U13377 (N_13377,N_12871,N_13160);
or U13378 (N_13378,N_12838,N_13192);
or U13379 (N_13379,N_13021,N_12958);
and U13380 (N_13380,N_12950,N_12984);
or U13381 (N_13381,N_13114,N_13174);
nand U13382 (N_13382,N_12974,N_12929);
and U13383 (N_13383,N_13030,N_12989);
or U13384 (N_13384,N_13137,N_13038);
nand U13385 (N_13385,N_13080,N_13168);
or U13386 (N_13386,N_13198,N_13172);
nor U13387 (N_13387,N_13039,N_13035);
or U13388 (N_13388,N_12976,N_12987);
nor U13389 (N_13389,N_13145,N_12917);
and U13390 (N_13390,N_13199,N_13062);
or U13391 (N_13391,N_13105,N_12966);
nor U13392 (N_13392,N_12825,N_12806);
nand U13393 (N_13393,N_12867,N_13120);
nor U13394 (N_13394,N_13056,N_13007);
xnor U13395 (N_13395,N_13188,N_13027);
nor U13396 (N_13396,N_12963,N_13064);
or U13397 (N_13397,N_12886,N_13179);
nand U13398 (N_13398,N_12955,N_12911);
nand U13399 (N_13399,N_12865,N_13117);
nand U13400 (N_13400,N_13092,N_13066);
xnor U13401 (N_13401,N_13198,N_12806);
xnor U13402 (N_13402,N_13143,N_13039);
nor U13403 (N_13403,N_12825,N_12849);
nor U13404 (N_13404,N_12885,N_13009);
and U13405 (N_13405,N_13042,N_13140);
nand U13406 (N_13406,N_12945,N_13085);
nand U13407 (N_13407,N_13183,N_13100);
xnor U13408 (N_13408,N_12885,N_13115);
nand U13409 (N_13409,N_13151,N_13102);
nor U13410 (N_13410,N_12971,N_13091);
or U13411 (N_13411,N_13110,N_13119);
nor U13412 (N_13412,N_12962,N_12820);
and U13413 (N_13413,N_12985,N_13144);
and U13414 (N_13414,N_12910,N_12968);
or U13415 (N_13415,N_12801,N_12859);
nand U13416 (N_13416,N_13151,N_13145);
and U13417 (N_13417,N_12916,N_12927);
xnor U13418 (N_13418,N_13108,N_12955);
and U13419 (N_13419,N_13081,N_12837);
xor U13420 (N_13420,N_12874,N_13096);
and U13421 (N_13421,N_13092,N_12832);
xnor U13422 (N_13422,N_13095,N_13196);
and U13423 (N_13423,N_12820,N_12835);
xnor U13424 (N_13424,N_12972,N_13139);
or U13425 (N_13425,N_13082,N_12880);
nand U13426 (N_13426,N_12994,N_13112);
nand U13427 (N_13427,N_12901,N_12878);
xnor U13428 (N_13428,N_13140,N_12925);
or U13429 (N_13429,N_12856,N_12855);
or U13430 (N_13430,N_12874,N_13027);
xor U13431 (N_13431,N_12999,N_12993);
nand U13432 (N_13432,N_13031,N_12994);
xnor U13433 (N_13433,N_13165,N_13072);
nand U13434 (N_13434,N_13087,N_12958);
and U13435 (N_13435,N_13083,N_13173);
and U13436 (N_13436,N_12806,N_13006);
nor U13437 (N_13437,N_13146,N_13073);
nor U13438 (N_13438,N_13117,N_13173);
xor U13439 (N_13439,N_13064,N_12855);
nor U13440 (N_13440,N_12947,N_12977);
xor U13441 (N_13441,N_13124,N_12934);
nor U13442 (N_13442,N_13092,N_12955);
nor U13443 (N_13443,N_13182,N_13091);
xnor U13444 (N_13444,N_12851,N_13064);
and U13445 (N_13445,N_13187,N_13112);
xor U13446 (N_13446,N_13076,N_12941);
or U13447 (N_13447,N_13199,N_13051);
and U13448 (N_13448,N_12830,N_13175);
nand U13449 (N_13449,N_12859,N_12993);
or U13450 (N_13450,N_12945,N_13132);
and U13451 (N_13451,N_12903,N_12971);
and U13452 (N_13452,N_12888,N_13161);
nor U13453 (N_13453,N_13103,N_12981);
and U13454 (N_13454,N_12816,N_12833);
or U13455 (N_13455,N_13056,N_13175);
nand U13456 (N_13456,N_13028,N_12921);
and U13457 (N_13457,N_13175,N_13061);
nor U13458 (N_13458,N_13032,N_13027);
and U13459 (N_13459,N_13176,N_13064);
or U13460 (N_13460,N_12851,N_13179);
nand U13461 (N_13461,N_13088,N_13001);
or U13462 (N_13462,N_13158,N_12817);
or U13463 (N_13463,N_12977,N_12871);
and U13464 (N_13464,N_13168,N_12946);
nor U13465 (N_13465,N_12815,N_13060);
nor U13466 (N_13466,N_13086,N_12950);
nor U13467 (N_13467,N_12937,N_13185);
and U13468 (N_13468,N_12905,N_13043);
nor U13469 (N_13469,N_12920,N_13078);
nor U13470 (N_13470,N_13053,N_12819);
nor U13471 (N_13471,N_12806,N_13003);
nand U13472 (N_13472,N_12874,N_13076);
xnor U13473 (N_13473,N_12864,N_13094);
xor U13474 (N_13474,N_13083,N_12894);
nor U13475 (N_13475,N_13003,N_12978);
or U13476 (N_13476,N_13136,N_13103);
or U13477 (N_13477,N_13138,N_13129);
nor U13478 (N_13478,N_13178,N_12910);
or U13479 (N_13479,N_12816,N_13107);
and U13480 (N_13480,N_12980,N_12843);
nor U13481 (N_13481,N_12963,N_13071);
xor U13482 (N_13482,N_13152,N_12801);
nand U13483 (N_13483,N_12968,N_13079);
or U13484 (N_13484,N_13090,N_13164);
nor U13485 (N_13485,N_12939,N_13063);
nand U13486 (N_13486,N_13083,N_12830);
xnor U13487 (N_13487,N_12974,N_13162);
nand U13488 (N_13488,N_12880,N_12884);
xor U13489 (N_13489,N_13176,N_13050);
nand U13490 (N_13490,N_13162,N_12816);
xnor U13491 (N_13491,N_12858,N_12933);
nand U13492 (N_13492,N_12967,N_13122);
or U13493 (N_13493,N_12900,N_13072);
xor U13494 (N_13494,N_12845,N_12889);
and U13495 (N_13495,N_12905,N_12825);
nor U13496 (N_13496,N_13067,N_13134);
or U13497 (N_13497,N_12835,N_12840);
xor U13498 (N_13498,N_12827,N_12869);
and U13499 (N_13499,N_13159,N_13102);
or U13500 (N_13500,N_13152,N_12910);
and U13501 (N_13501,N_13162,N_12850);
or U13502 (N_13502,N_12807,N_13092);
nand U13503 (N_13503,N_13100,N_13097);
and U13504 (N_13504,N_13171,N_12813);
or U13505 (N_13505,N_12846,N_12861);
and U13506 (N_13506,N_12897,N_13112);
nor U13507 (N_13507,N_12990,N_13089);
nand U13508 (N_13508,N_13029,N_12863);
or U13509 (N_13509,N_13103,N_12962);
nor U13510 (N_13510,N_13052,N_12892);
nor U13511 (N_13511,N_12855,N_13043);
nor U13512 (N_13512,N_13025,N_13188);
nand U13513 (N_13513,N_12955,N_12847);
and U13514 (N_13514,N_12906,N_13007);
xnor U13515 (N_13515,N_13023,N_13115);
nand U13516 (N_13516,N_13112,N_12843);
nor U13517 (N_13517,N_12906,N_13097);
and U13518 (N_13518,N_13162,N_13131);
nor U13519 (N_13519,N_13003,N_13047);
and U13520 (N_13520,N_12890,N_13140);
nand U13521 (N_13521,N_13014,N_13037);
nor U13522 (N_13522,N_12813,N_13152);
or U13523 (N_13523,N_13104,N_12863);
xnor U13524 (N_13524,N_13111,N_12856);
nand U13525 (N_13525,N_13043,N_13153);
nand U13526 (N_13526,N_13017,N_12801);
and U13527 (N_13527,N_12807,N_13116);
nand U13528 (N_13528,N_12802,N_12926);
nor U13529 (N_13529,N_13191,N_13004);
and U13530 (N_13530,N_13187,N_12910);
or U13531 (N_13531,N_12899,N_12976);
nand U13532 (N_13532,N_12935,N_13052);
and U13533 (N_13533,N_12932,N_13039);
xnor U13534 (N_13534,N_13012,N_13089);
nand U13535 (N_13535,N_13082,N_13107);
nor U13536 (N_13536,N_13076,N_13166);
or U13537 (N_13537,N_13177,N_13016);
or U13538 (N_13538,N_13090,N_12851);
and U13539 (N_13539,N_13110,N_13038);
and U13540 (N_13540,N_12863,N_13101);
xor U13541 (N_13541,N_12913,N_13107);
nand U13542 (N_13542,N_13116,N_12950);
nand U13543 (N_13543,N_13130,N_13124);
nor U13544 (N_13544,N_12875,N_12978);
nor U13545 (N_13545,N_12909,N_13000);
or U13546 (N_13546,N_12829,N_13058);
nor U13547 (N_13547,N_12808,N_13013);
or U13548 (N_13548,N_13010,N_12915);
nor U13549 (N_13549,N_13031,N_12829);
xnor U13550 (N_13550,N_13198,N_13038);
nor U13551 (N_13551,N_12897,N_12868);
nand U13552 (N_13552,N_13169,N_12907);
nand U13553 (N_13553,N_12866,N_13069);
nand U13554 (N_13554,N_12831,N_13058);
nand U13555 (N_13555,N_12918,N_12979);
nor U13556 (N_13556,N_13052,N_13063);
or U13557 (N_13557,N_13095,N_12923);
or U13558 (N_13558,N_13174,N_12829);
xnor U13559 (N_13559,N_12805,N_12977);
nor U13560 (N_13560,N_13079,N_12893);
or U13561 (N_13561,N_12961,N_13098);
or U13562 (N_13562,N_13066,N_13088);
xnor U13563 (N_13563,N_12839,N_12948);
xor U13564 (N_13564,N_12888,N_12940);
and U13565 (N_13565,N_12823,N_12905);
nor U13566 (N_13566,N_13041,N_13076);
nand U13567 (N_13567,N_12830,N_13048);
nor U13568 (N_13568,N_13190,N_12915);
xor U13569 (N_13569,N_13031,N_12983);
nor U13570 (N_13570,N_12972,N_13133);
and U13571 (N_13571,N_13069,N_12991);
or U13572 (N_13572,N_13194,N_12994);
and U13573 (N_13573,N_12878,N_12861);
xnor U13574 (N_13574,N_13117,N_13066);
or U13575 (N_13575,N_13169,N_13158);
xor U13576 (N_13576,N_13012,N_12915);
nand U13577 (N_13577,N_13101,N_13137);
nand U13578 (N_13578,N_12875,N_12865);
nand U13579 (N_13579,N_12983,N_13117);
nor U13580 (N_13580,N_13172,N_12810);
or U13581 (N_13581,N_13111,N_12961);
xor U13582 (N_13582,N_13009,N_12908);
nand U13583 (N_13583,N_13092,N_12910);
xnor U13584 (N_13584,N_13186,N_13172);
xor U13585 (N_13585,N_13174,N_12947);
xnor U13586 (N_13586,N_12814,N_13039);
nor U13587 (N_13587,N_13011,N_13156);
nor U13588 (N_13588,N_12982,N_12851);
nand U13589 (N_13589,N_12804,N_13194);
and U13590 (N_13590,N_12992,N_12926);
xnor U13591 (N_13591,N_13134,N_12889);
and U13592 (N_13592,N_13061,N_12985);
and U13593 (N_13593,N_13053,N_12832);
nor U13594 (N_13594,N_13016,N_12831);
or U13595 (N_13595,N_13086,N_12912);
xnor U13596 (N_13596,N_13103,N_12845);
and U13597 (N_13597,N_12821,N_13024);
xnor U13598 (N_13598,N_13086,N_13144);
and U13599 (N_13599,N_13199,N_13035);
nor U13600 (N_13600,N_13559,N_13530);
xor U13601 (N_13601,N_13260,N_13282);
and U13602 (N_13602,N_13494,N_13216);
xor U13603 (N_13603,N_13259,N_13444);
nor U13604 (N_13604,N_13548,N_13541);
or U13605 (N_13605,N_13536,N_13438);
or U13606 (N_13606,N_13545,N_13320);
and U13607 (N_13607,N_13315,N_13360);
xnor U13608 (N_13608,N_13553,N_13466);
and U13609 (N_13609,N_13249,N_13254);
or U13610 (N_13610,N_13434,N_13273);
nand U13611 (N_13611,N_13465,N_13318);
nor U13612 (N_13612,N_13366,N_13329);
nor U13613 (N_13613,N_13392,N_13317);
or U13614 (N_13614,N_13592,N_13323);
xnor U13615 (N_13615,N_13587,N_13201);
xor U13616 (N_13616,N_13414,N_13303);
and U13617 (N_13617,N_13246,N_13326);
or U13618 (N_13618,N_13253,N_13525);
nor U13619 (N_13619,N_13212,N_13538);
nor U13620 (N_13620,N_13308,N_13584);
xor U13621 (N_13621,N_13402,N_13413);
xor U13622 (N_13622,N_13281,N_13341);
nand U13623 (N_13623,N_13575,N_13492);
nand U13624 (N_13624,N_13322,N_13412);
xor U13625 (N_13625,N_13440,N_13537);
nor U13626 (N_13626,N_13514,N_13516);
and U13627 (N_13627,N_13487,N_13241);
nand U13628 (N_13628,N_13390,N_13579);
or U13629 (N_13629,N_13554,N_13382);
or U13630 (N_13630,N_13550,N_13519);
nand U13631 (N_13631,N_13256,N_13279);
or U13632 (N_13632,N_13431,N_13343);
nand U13633 (N_13633,N_13503,N_13297);
nand U13634 (N_13634,N_13513,N_13217);
nor U13635 (N_13635,N_13331,N_13407);
or U13636 (N_13636,N_13262,N_13400);
nand U13637 (N_13637,N_13266,N_13333);
or U13638 (N_13638,N_13339,N_13580);
xnor U13639 (N_13639,N_13226,N_13277);
nand U13640 (N_13640,N_13533,N_13381);
and U13641 (N_13641,N_13286,N_13264);
or U13642 (N_13642,N_13300,N_13247);
xor U13643 (N_13643,N_13508,N_13376);
nand U13644 (N_13644,N_13258,N_13500);
and U13645 (N_13645,N_13478,N_13280);
nor U13646 (N_13646,N_13257,N_13418);
and U13647 (N_13647,N_13534,N_13454);
nor U13648 (N_13648,N_13370,N_13229);
nand U13649 (N_13649,N_13427,N_13419);
and U13650 (N_13650,N_13347,N_13557);
nor U13651 (N_13651,N_13213,N_13378);
or U13652 (N_13652,N_13396,N_13589);
nor U13653 (N_13653,N_13263,N_13416);
xnor U13654 (N_13654,N_13437,N_13476);
nand U13655 (N_13655,N_13345,N_13210);
or U13656 (N_13656,N_13274,N_13288);
and U13657 (N_13657,N_13380,N_13540);
and U13658 (N_13658,N_13599,N_13205);
nand U13659 (N_13659,N_13316,N_13566);
or U13660 (N_13660,N_13447,N_13523);
or U13661 (N_13661,N_13251,N_13406);
xor U13662 (N_13662,N_13549,N_13321);
or U13663 (N_13663,N_13235,N_13255);
nand U13664 (N_13664,N_13302,N_13325);
xor U13665 (N_13665,N_13219,N_13459);
or U13666 (N_13666,N_13207,N_13222);
nand U13667 (N_13667,N_13386,N_13574);
nand U13668 (N_13668,N_13420,N_13375);
or U13669 (N_13669,N_13479,N_13348);
and U13670 (N_13670,N_13598,N_13489);
nand U13671 (N_13671,N_13203,N_13501);
xnor U13672 (N_13672,N_13240,N_13410);
or U13673 (N_13673,N_13464,N_13445);
nand U13674 (N_13674,N_13441,N_13312);
and U13675 (N_13675,N_13577,N_13586);
xor U13676 (N_13676,N_13337,N_13232);
and U13677 (N_13677,N_13327,N_13383);
nand U13678 (N_13678,N_13563,N_13502);
or U13679 (N_13679,N_13363,N_13298);
nor U13680 (N_13680,N_13446,N_13453);
xnor U13681 (N_13681,N_13324,N_13568);
xnor U13682 (N_13682,N_13524,N_13299);
nand U13683 (N_13683,N_13475,N_13517);
nor U13684 (N_13684,N_13456,N_13428);
or U13685 (N_13685,N_13289,N_13417);
xor U13686 (N_13686,N_13356,N_13582);
or U13687 (N_13687,N_13421,N_13353);
nor U13688 (N_13688,N_13384,N_13368);
and U13689 (N_13689,N_13591,N_13543);
and U13690 (N_13690,N_13531,N_13439);
nand U13691 (N_13691,N_13509,N_13291);
and U13692 (N_13692,N_13265,N_13481);
and U13693 (N_13693,N_13372,N_13228);
nor U13694 (N_13694,N_13310,N_13387);
xor U13695 (N_13695,N_13371,N_13358);
nor U13696 (N_13696,N_13346,N_13527);
nand U13697 (N_13697,N_13261,N_13474);
nand U13698 (N_13698,N_13369,N_13362);
or U13699 (N_13699,N_13237,N_13547);
and U13700 (N_13700,N_13571,N_13483);
and U13701 (N_13701,N_13340,N_13471);
and U13702 (N_13702,N_13275,N_13344);
nand U13703 (N_13703,N_13485,N_13304);
and U13704 (N_13704,N_13578,N_13561);
nand U13705 (N_13705,N_13367,N_13330);
and U13706 (N_13706,N_13388,N_13399);
and U13707 (N_13707,N_13335,N_13520);
or U13708 (N_13708,N_13542,N_13511);
and U13709 (N_13709,N_13208,N_13585);
and U13710 (N_13710,N_13292,N_13238);
nand U13711 (N_13711,N_13433,N_13305);
xnor U13712 (N_13712,N_13521,N_13393);
and U13713 (N_13713,N_13473,N_13405);
and U13714 (N_13714,N_13460,N_13349);
nor U13715 (N_13715,N_13342,N_13234);
or U13716 (N_13716,N_13472,N_13595);
nor U13717 (N_13717,N_13546,N_13432);
or U13718 (N_13718,N_13252,N_13470);
or U13719 (N_13719,N_13209,N_13569);
nand U13720 (N_13720,N_13499,N_13354);
or U13721 (N_13721,N_13290,N_13597);
and U13722 (N_13722,N_13429,N_13458);
nor U13723 (N_13723,N_13204,N_13573);
and U13724 (N_13724,N_13214,N_13270);
and U13725 (N_13725,N_13355,N_13491);
xor U13726 (N_13726,N_13463,N_13236);
xnor U13727 (N_13727,N_13409,N_13581);
nor U13728 (N_13728,N_13436,N_13359);
nor U13729 (N_13729,N_13518,N_13462);
or U13730 (N_13730,N_13225,N_13495);
nand U13731 (N_13731,N_13596,N_13497);
xor U13732 (N_13732,N_13215,N_13552);
and U13733 (N_13733,N_13248,N_13334);
nand U13734 (N_13734,N_13200,N_13422);
or U13735 (N_13735,N_13389,N_13496);
or U13736 (N_13736,N_13336,N_13352);
or U13737 (N_13737,N_13361,N_13296);
nand U13738 (N_13738,N_13594,N_13461);
nor U13739 (N_13739,N_13364,N_13588);
nor U13740 (N_13740,N_13220,N_13233);
nor U13741 (N_13741,N_13398,N_13357);
nand U13742 (N_13742,N_13504,N_13539);
or U13743 (N_13743,N_13243,N_13468);
nand U13744 (N_13744,N_13283,N_13272);
nand U13745 (N_13745,N_13211,N_13245);
nand U13746 (N_13746,N_13424,N_13306);
and U13747 (N_13747,N_13206,N_13505);
nand U13748 (N_13748,N_13532,N_13576);
xor U13749 (N_13749,N_13408,N_13227);
nor U13750 (N_13750,N_13560,N_13564);
xor U13751 (N_13751,N_13425,N_13293);
and U13752 (N_13752,N_13507,N_13506);
and U13753 (N_13753,N_13309,N_13332);
or U13754 (N_13754,N_13284,N_13452);
xor U13755 (N_13755,N_13477,N_13269);
and U13756 (N_13756,N_13224,N_13484);
nor U13757 (N_13757,N_13469,N_13480);
or U13758 (N_13758,N_13457,N_13311);
xor U13759 (N_13759,N_13488,N_13328);
or U13760 (N_13760,N_13295,N_13319);
nand U13761 (N_13761,N_13450,N_13313);
xnor U13762 (N_13762,N_13583,N_13285);
xnor U13763 (N_13763,N_13239,N_13415);
xnor U13764 (N_13764,N_13526,N_13271);
or U13765 (N_13765,N_13558,N_13482);
nor U13766 (N_13766,N_13373,N_13377);
nand U13767 (N_13767,N_13572,N_13395);
xnor U13768 (N_13768,N_13567,N_13314);
nand U13769 (N_13769,N_13448,N_13231);
or U13770 (N_13770,N_13529,N_13449);
xnor U13771 (N_13771,N_13430,N_13486);
and U13772 (N_13772,N_13268,N_13307);
xor U13773 (N_13773,N_13221,N_13394);
and U13774 (N_13774,N_13365,N_13555);
and U13775 (N_13775,N_13223,N_13455);
xnor U13776 (N_13776,N_13287,N_13544);
xor U13777 (N_13777,N_13490,N_13338);
nor U13778 (N_13778,N_13385,N_13593);
xor U13779 (N_13779,N_13556,N_13351);
or U13780 (N_13780,N_13267,N_13551);
nor U13781 (N_13781,N_13512,N_13411);
and U13782 (N_13782,N_13590,N_13565);
nor U13783 (N_13783,N_13562,N_13230);
nand U13784 (N_13784,N_13244,N_13374);
nor U13785 (N_13785,N_13528,N_13442);
nand U13786 (N_13786,N_13276,N_13379);
and U13787 (N_13787,N_13202,N_13426);
or U13788 (N_13788,N_13493,N_13218);
and U13789 (N_13789,N_13467,N_13301);
xnor U13790 (N_13790,N_13242,N_13278);
and U13791 (N_13791,N_13350,N_13515);
nand U13792 (N_13792,N_13535,N_13294);
nand U13793 (N_13793,N_13397,N_13570);
nand U13794 (N_13794,N_13443,N_13522);
xor U13795 (N_13795,N_13423,N_13401);
nand U13796 (N_13796,N_13250,N_13451);
nand U13797 (N_13797,N_13391,N_13510);
or U13798 (N_13798,N_13403,N_13404);
or U13799 (N_13799,N_13435,N_13498);
xnor U13800 (N_13800,N_13335,N_13210);
and U13801 (N_13801,N_13258,N_13396);
xnor U13802 (N_13802,N_13309,N_13274);
or U13803 (N_13803,N_13461,N_13381);
nand U13804 (N_13804,N_13236,N_13505);
and U13805 (N_13805,N_13311,N_13330);
xor U13806 (N_13806,N_13508,N_13286);
or U13807 (N_13807,N_13467,N_13493);
nor U13808 (N_13808,N_13394,N_13527);
nand U13809 (N_13809,N_13252,N_13362);
nand U13810 (N_13810,N_13351,N_13445);
and U13811 (N_13811,N_13288,N_13388);
and U13812 (N_13812,N_13427,N_13282);
and U13813 (N_13813,N_13314,N_13406);
nor U13814 (N_13814,N_13325,N_13296);
nor U13815 (N_13815,N_13535,N_13378);
or U13816 (N_13816,N_13268,N_13297);
nor U13817 (N_13817,N_13326,N_13341);
nor U13818 (N_13818,N_13367,N_13260);
or U13819 (N_13819,N_13338,N_13580);
xor U13820 (N_13820,N_13480,N_13382);
nor U13821 (N_13821,N_13408,N_13474);
or U13822 (N_13822,N_13452,N_13443);
nand U13823 (N_13823,N_13500,N_13271);
nand U13824 (N_13824,N_13311,N_13427);
nor U13825 (N_13825,N_13351,N_13208);
and U13826 (N_13826,N_13563,N_13509);
and U13827 (N_13827,N_13286,N_13409);
or U13828 (N_13828,N_13332,N_13552);
xor U13829 (N_13829,N_13350,N_13227);
and U13830 (N_13830,N_13228,N_13579);
nor U13831 (N_13831,N_13321,N_13340);
or U13832 (N_13832,N_13526,N_13236);
or U13833 (N_13833,N_13552,N_13352);
nor U13834 (N_13834,N_13521,N_13422);
and U13835 (N_13835,N_13414,N_13454);
nor U13836 (N_13836,N_13329,N_13437);
and U13837 (N_13837,N_13409,N_13281);
and U13838 (N_13838,N_13334,N_13348);
and U13839 (N_13839,N_13266,N_13405);
and U13840 (N_13840,N_13439,N_13448);
nand U13841 (N_13841,N_13210,N_13521);
nand U13842 (N_13842,N_13378,N_13437);
xnor U13843 (N_13843,N_13372,N_13474);
and U13844 (N_13844,N_13440,N_13434);
xnor U13845 (N_13845,N_13481,N_13321);
and U13846 (N_13846,N_13279,N_13223);
or U13847 (N_13847,N_13444,N_13475);
xor U13848 (N_13848,N_13244,N_13390);
or U13849 (N_13849,N_13458,N_13537);
and U13850 (N_13850,N_13483,N_13596);
nor U13851 (N_13851,N_13415,N_13473);
nand U13852 (N_13852,N_13527,N_13339);
nand U13853 (N_13853,N_13260,N_13575);
xnor U13854 (N_13854,N_13446,N_13532);
nand U13855 (N_13855,N_13250,N_13417);
or U13856 (N_13856,N_13587,N_13307);
xor U13857 (N_13857,N_13281,N_13286);
and U13858 (N_13858,N_13318,N_13248);
xor U13859 (N_13859,N_13278,N_13369);
nand U13860 (N_13860,N_13521,N_13282);
nand U13861 (N_13861,N_13433,N_13493);
and U13862 (N_13862,N_13282,N_13542);
and U13863 (N_13863,N_13565,N_13598);
or U13864 (N_13864,N_13269,N_13395);
or U13865 (N_13865,N_13258,N_13531);
and U13866 (N_13866,N_13590,N_13429);
or U13867 (N_13867,N_13497,N_13495);
xor U13868 (N_13868,N_13475,N_13248);
or U13869 (N_13869,N_13369,N_13527);
nor U13870 (N_13870,N_13306,N_13361);
xnor U13871 (N_13871,N_13530,N_13456);
or U13872 (N_13872,N_13236,N_13541);
or U13873 (N_13873,N_13519,N_13399);
and U13874 (N_13874,N_13247,N_13529);
nor U13875 (N_13875,N_13597,N_13300);
or U13876 (N_13876,N_13396,N_13414);
and U13877 (N_13877,N_13212,N_13323);
and U13878 (N_13878,N_13301,N_13257);
or U13879 (N_13879,N_13337,N_13583);
nand U13880 (N_13880,N_13430,N_13471);
or U13881 (N_13881,N_13541,N_13280);
nor U13882 (N_13882,N_13445,N_13205);
or U13883 (N_13883,N_13493,N_13421);
or U13884 (N_13884,N_13217,N_13397);
xnor U13885 (N_13885,N_13431,N_13599);
and U13886 (N_13886,N_13444,N_13531);
nand U13887 (N_13887,N_13314,N_13339);
xor U13888 (N_13888,N_13493,N_13392);
nor U13889 (N_13889,N_13578,N_13242);
or U13890 (N_13890,N_13442,N_13285);
nand U13891 (N_13891,N_13317,N_13200);
and U13892 (N_13892,N_13300,N_13433);
nand U13893 (N_13893,N_13340,N_13268);
nand U13894 (N_13894,N_13307,N_13361);
and U13895 (N_13895,N_13384,N_13554);
nor U13896 (N_13896,N_13466,N_13497);
or U13897 (N_13897,N_13310,N_13440);
nand U13898 (N_13898,N_13251,N_13329);
and U13899 (N_13899,N_13426,N_13447);
nand U13900 (N_13900,N_13517,N_13553);
nand U13901 (N_13901,N_13230,N_13592);
nor U13902 (N_13902,N_13276,N_13571);
and U13903 (N_13903,N_13352,N_13200);
nand U13904 (N_13904,N_13226,N_13258);
and U13905 (N_13905,N_13556,N_13219);
xor U13906 (N_13906,N_13257,N_13296);
nor U13907 (N_13907,N_13518,N_13322);
or U13908 (N_13908,N_13441,N_13286);
xnor U13909 (N_13909,N_13438,N_13257);
xor U13910 (N_13910,N_13406,N_13413);
xor U13911 (N_13911,N_13207,N_13423);
or U13912 (N_13912,N_13324,N_13316);
nor U13913 (N_13913,N_13347,N_13407);
xor U13914 (N_13914,N_13267,N_13252);
nand U13915 (N_13915,N_13435,N_13449);
or U13916 (N_13916,N_13569,N_13498);
xnor U13917 (N_13917,N_13597,N_13491);
or U13918 (N_13918,N_13329,N_13261);
or U13919 (N_13919,N_13489,N_13437);
and U13920 (N_13920,N_13207,N_13541);
xor U13921 (N_13921,N_13569,N_13315);
or U13922 (N_13922,N_13447,N_13212);
nor U13923 (N_13923,N_13568,N_13470);
and U13924 (N_13924,N_13363,N_13583);
or U13925 (N_13925,N_13216,N_13241);
nand U13926 (N_13926,N_13323,N_13426);
nand U13927 (N_13927,N_13246,N_13257);
nand U13928 (N_13928,N_13563,N_13531);
or U13929 (N_13929,N_13374,N_13530);
nor U13930 (N_13930,N_13503,N_13341);
and U13931 (N_13931,N_13212,N_13364);
xor U13932 (N_13932,N_13408,N_13442);
nand U13933 (N_13933,N_13414,N_13480);
and U13934 (N_13934,N_13407,N_13201);
xnor U13935 (N_13935,N_13434,N_13208);
or U13936 (N_13936,N_13406,N_13419);
nand U13937 (N_13937,N_13495,N_13322);
and U13938 (N_13938,N_13235,N_13267);
or U13939 (N_13939,N_13294,N_13219);
nor U13940 (N_13940,N_13326,N_13332);
nand U13941 (N_13941,N_13431,N_13330);
nor U13942 (N_13942,N_13232,N_13367);
xor U13943 (N_13943,N_13589,N_13276);
xor U13944 (N_13944,N_13302,N_13502);
and U13945 (N_13945,N_13272,N_13248);
nand U13946 (N_13946,N_13267,N_13384);
and U13947 (N_13947,N_13288,N_13214);
nor U13948 (N_13948,N_13248,N_13461);
or U13949 (N_13949,N_13552,N_13461);
or U13950 (N_13950,N_13298,N_13327);
or U13951 (N_13951,N_13252,N_13523);
nor U13952 (N_13952,N_13373,N_13446);
nor U13953 (N_13953,N_13380,N_13240);
nand U13954 (N_13954,N_13522,N_13487);
xnor U13955 (N_13955,N_13552,N_13359);
nand U13956 (N_13956,N_13477,N_13226);
nor U13957 (N_13957,N_13498,N_13507);
nor U13958 (N_13958,N_13319,N_13387);
nor U13959 (N_13959,N_13360,N_13556);
xnor U13960 (N_13960,N_13440,N_13499);
and U13961 (N_13961,N_13395,N_13450);
nor U13962 (N_13962,N_13272,N_13348);
or U13963 (N_13963,N_13291,N_13211);
and U13964 (N_13964,N_13585,N_13548);
or U13965 (N_13965,N_13338,N_13590);
or U13966 (N_13966,N_13312,N_13305);
and U13967 (N_13967,N_13556,N_13347);
and U13968 (N_13968,N_13534,N_13588);
nor U13969 (N_13969,N_13488,N_13551);
nor U13970 (N_13970,N_13592,N_13218);
or U13971 (N_13971,N_13599,N_13548);
and U13972 (N_13972,N_13361,N_13437);
or U13973 (N_13973,N_13476,N_13441);
or U13974 (N_13974,N_13258,N_13376);
nand U13975 (N_13975,N_13455,N_13280);
xnor U13976 (N_13976,N_13418,N_13512);
nor U13977 (N_13977,N_13371,N_13594);
xnor U13978 (N_13978,N_13469,N_13483);
or U13979 (N_13979,N_13561,N_13281);
nand U13980 (N_13980,N_13540,N_13237);
or U13981 (N_13981,N_13221,N_13534);
nand U13982 (N_13982,N_13432,N_13573);
xor U13983 (N_13983,N_13237,N_13351);
nor U13984 (N_13984,N_13283,N_13407);
xnor U13985 (N_13985,N_13284,N_13542);
xnor U13986 (N_13986,N_13455,N_13307);
and U13987 (N_13987,N_13250,N_13264);
or U13988 (N_13988,N_13400,N_13209);
nor U13989 (N_13989,N_13469,N_13542);
or U13990 (N_13990,N_13310,N_13203);
or U13991 (N_13991,N_13327,N_13562);
nor U13992 (N_13992,N_13510,N_13508);
and U13993 (N_13993,N_13403,N_13300);
and U13994 (N_13994,N_13224,N_13527);
and U13995 (N_13995,N_13368,N_13296);
or U13996 (N_13996,N_13514,N_13493);
nand U13997 (N_13997,N_13307,N_13332);
and U13998 (N_13998,N_13560,N_13388);
or U13999 (N_13999,N_13515,N_13401);
or U14000 (N_14000,N_13789,N_13716);
or U14001 (N_14001,N_13765,N_13724);
nand U14002 (N_14002,N_13720,N_13824);
nand U14003 (N_14003,N_13618,N_13679);
nand U14004 (N_14004,N_13800,N_13877);
xor U14005 (N_14005,N_13680,N_13703);
nor U14006 (N_14006,N_13889,N_13657);
nor U14007 (N_14007,N_13777,N_13871);
xor U14008 (N_14008,N_13880,N_13661);
nand U14009 (N_14009,N_13715,N_13641);
or U14010 (N_14010,N_13602,N_13975);
xor U14011 (N_14011,N_13826,N_13902);
and U14012 (N_14012,N_13639,N_13979);
nand U14013 (N_14013,N_13686,N_13792);
nor U14014 (N_14014,N_13914,N_13947);
nor U14015 (N_14015,N_13912,N_13663);
and U14016 (N_14016,N_13901,N_13887);
nand U14017 (N_14017,N_13961,N_13814);
nand U14018 (N_14018,N_13713,N_13820);
nand U14019 (N_14019,N_13729,N_13926);
nand U14020 (N_14020,N_13832,N_13822);
xnor U14021 (N_14021,N_13885,N_13678);
nand U14022 (N_14022,N_13948,N_13896);
xnor U14023 (N_14023,N_13778,N_13834);
xor U14024 (N_14024,N_13699,N_13754);
nand U14025 (N_14025,N_13984,N_13675);
xor U14026 (N_14026,N_13853,N_13795);
nor U14027 (N_14027,N_13952,N_13849);
nand U14028 (N_14028,N_13764,N_13631);
or U14029 (N_14029,N_13684,N_13812);
nand U14030 (N_14030,N_13968,N_13904);
xor U14031 (N_14031,N_13927,N_13714);
xor U14032 (N_14032,N_13941,N_13828);
nand U14033 (N_14033,N_13770,N_13845);
xor U14034 (N_14034,N_13806,N_13980);
or U14035 (N_14035,N_13752,N_13868);
nor U14036 (N_14036,N_13647,N_13852);
or U14037 (N_14037,N_13673,N_13874);
xnor U14038 (N_14038,N_13674,N_13883);
nor U14039 (N_14039,N_13933,N_13935);
nand U14040 (N_14040,N_13791,N_13925);
nor U14041 (N_14041,N_13666,N_13794);
and U14042 (N_14042,N_13900,N_13707);
nor U14043 (N_14043,N_13760,N_13876);
xor U14044 (N_14044,N_13604,N_13704);
nand U14045 (N_14045,N_13739,N_13816);
xnor U14046 (N_14046,N_13932,N_13774);
xnor U14047 (N_14047,N_13632,N_13668);
or U14048 (N_14048,N_13950,N_13971);
xnor U14049 (N_14049,N_13808,N_13992);
or U14050 (N_14050,N_13998,N_13654);
and U14051 (N_14051,N_13861,N_13767);
nor U14052 (N_14052,N_13997,N_13987);
nor U14053 (N_14053,N_13700,N_13805);
nor U14054 (N_14054,N_13881,N_13905);
nand U14055 (N_14055,N_13804,N_13913);
nor U14056 (N_14056,N_13835,N_13859);
and U14057 (N_14057,N_13807,N_13610);
xor U14058 (N_14058,N_13911,N_13847);
or U14059 (N_14059,N_13642,N_13953);
xnor U14060 (N_14060,N_13685,N_13693);
xnor U14061 (N_14061,N_13648,N_13626);
or U14062 (N_14062,N_13972,N_13891);
or U14063 (N_14063,N_13895,N_13978);
and U14064 (N_14064,N_13687,N_13636);
xor U14065 (N_14065,N_13938,N_13709);
xnor U14066 (N_14066,N_13919,N_13793);
nand U14067 (N_14067,N_13732,N_13624);
nand U14068 (N_14068,N_13683,N_13983);
nand U14069 (N_14069,N_13612,N_13934);
xor U14070 (N_14070,N_13633,N_13817);
nand U14071 (N_14071,N_13823,N_13866);
and U14072 (N_14072,N_13917,N_13974);
or U14073 (N_14073,N_13784,N_13839);
or U14074 (N_14074,N_13977,N_13848);
or U14075 (N_14075,N_13909,N_13608);
nand U14076 (N_14076,N_13875,N_13613);
nor U14077 (N_14077,N_13655,N_13836);
and U14078 (N_14078,N_13882,N_13640);
xnor U14079 (N_14079,N_13991,N_13734);
or U14080 (N_14080,N_13884,N_13898);
or U14081 (N_14081,N_13727,N_13659);
xor U14082 (N_14082,N_13855,N_13989);
or U14083 (N_14083,N_13862,N_13782);
and U14084 (N_14084,N_13959,N_13737);
nand U14085 (N_14085,N_13603,N_13776);
or U14086 (N_14086,N_13712,N_13965);
and U14087 (N_14087,N_13827,N_13928);
nand U14088 (N_14088,N_13843,N_13711);
and U14089 (N_14089,N_13924,N_13643);
nand U14090 (N_14090,N_13981,N_13656);
or U14091 (N_14091,N_13753,N_13779);
xor U14092 (N_14092,N_13606,N_13821);
and U14093 (N_14093,N_13830,N_13811);
and U14094 (N_14094,N_13653,N_13878);
or U14095 (N_14095,N_13733,N_13923);
or U14096 (N_14096,N_13746,N_13689);
nor U14097 (N_14097,N_13630,N_13818);
nand U14098 (N_14098,N_13665,N_13735);
or U14099 (N_14099,N_13993,N_13797);
nand U14100 (N_14100,N_13728,N_13757);
nand U14101 (N_14101,N_13825,N_13694);
and U14102 (N_14102,N_13936,N_13681);
nor U14103 (N_14103,N_13740,N_13736);
nand U14104 (N_14104,N_13725,N_13634);
and U14105 (N_14105,N_13614,N_13801);
xor U14106 (N_14106,N_13677,N_13802);
xor U14107 (N_14107,N_13809,N_13745);
nand U14108 (N_14108,N_13646,N_13682);
nand U14109 (N_14109,N_13958,N_13966);
or U14110 (N_14110,N_13622,N_13854);
nand U14111 (N_14111,N_13619,N_13956);
nand U14112 (N_14112,N_13629,N_13705);
and U14113 (N_14113,N_13942,N_13787);
nor U14114 (N_14114,N_13692,N_13988);
xnor U14115 (N_14115,N_13831,N_13637);
xnor U14116 (N_14116,N_13710,N_13688);
and U14117 (N_14117,N_13755,N_13903);
nand U14118 (N_14118,N_13708,N_13899);
and U14119 (N_14119,N_13644,N_13783);
nor U14120 (N_14120,N_13892,N_13940);
nor U14121 (N_14121,N_13717,N_13813);
xor U14122 (N_14122,N_13960,N_13731);
nand U14123 (N_14123,N_13951,N_13841);
nand U14124 (N_14124,N_13999,N_13970);
or U14125 (N_14125,N_13930,N_13962);
xnor U14126 (N_14126,N_13916,N_13869);
and U14127 (N_14127,N_13769,N_13922);
and U14128 (N_14128,N_13929,N_13638);
xor U14129 (N_14129,N_13945,N_13621);
nor U14130 (N_14130,N_13844,N_13890);
and U14131 (N_14131,N_13623,N_13718);
nand U14132 (N_14132,N_13773,N_13920);
nor U14133 (N_14133,N_13837,N_13766);
nor U14134 (N_14134,N_13963,N_13625);
nor U14135 (N_14135,N_13601,N_13662);
nor U14136 (N_14136,N_13751,N_13628);
and U14137 (N_14137,N_13756,N_13994);
nor U14138 (N_14138,N_13937,N_13780);
nor U14139 (N_14139,N_13915,N_13650);
and U14140 (N_14140,N_13873,N_13858);
and U14141 (N_14141,N_13719,N_13796);
xnor U14142 (N_14142,N_13605,N_13886);
xnor U14143 (N_14143,N_13609,N_13698);
nor U14144 (N_14144,N_13872,N_13652);
and U14145 (N_14145,N_13939,N_13833);
and U14146 (N_14146,N_13671,N_13726);
or U14147 (N_14147,N_13888,N_13943);
or U14148 (N_14148,N_13747,N_13730);
nor U14149 (N_14149,N_13600,N_13645);
nand U14150 (N_14150,N_13672,N_13676);
nor U14151 (N_14151,N_13664,N_13907);
and U14152 (N_14152,N_13721,N_13857);
and U14153 (N_14153,N_13893,N_13949);
and U14154 (N_14154,N_13864,N_13722);
nor U14155 (N_14155,N_13658,N_13781);
and U14156 (N_14156,N_13763,N_13759);
nand U14157 (N_14157,N_13667,N_13616);
xnor U14158 (N_14158,N_13607,N_13840);
or U14159 (N_14159,N_13856,N_13867);
nor U14160 (N_14160,N_13790,N_13696);
and U14161 (N_14161,N_13748,N_13846);
or U14162 (N_14162,N_13660,N_13870);
and U14163 (N_14163,N_13738,N_13771);
or U14164 (N_14164,N_13620,N_13908);
nor U14165 (N_14165,N_13964,N_13986);
nand U14166 (N_14166,N_13851,N_13955);
nor U14167 (N_14167,N_13611,N_13810);
xor U14168 (N_14168,N_13985,N_13695);
nor U14169 (N_14169,N_13976,N_13615);
xnor U14170 (N_14170,N_13897,N_13838);
or U14171 (N_14171,N_13921,N_13918);
and U14172 (N_14172,N_13967,N_13750);
and U14173 (N_14173,N_13649,N_13995);
and U14174 (N_14174,N_13706,N_13946);
and U14175 (N_14175,N_13651,N_13617);
nand U14176 (N_14176,N_13842,N_13957);
xnor U14177 (N_14177,N_13786,N_13973);
and U14178 (N_14178,N_13775,N_13762);
xnor U14179 (N_14179,N_13996,N_13879);
or U14180 (N_14180,N_13969,N_13744);
and U14181 (N_14181,N_13669,N_13785);
or U14182 (N_14182,N_13627,N_13691);
and U14183 (N_14183,N_13954,N_13788);
xor U14184 (N_14184,N_13906,N_13865);
or U14185 (N_14185,N_13863,N_13742);
nor U14186 (N_14186,N_13743,N_13768);
or U14187 (N_14187,N_13635,N_13829);
and U14188 (N_14188,N_13799,N_13741);
nand U14189 (N_14189,N_13910,N_13670);
nand U14190 (N_14190,N_13819,N_13815);
nor U14191 (N_14191,N_13944,N_13749);
nand U14192 (N_14192,N_13982,N_13702);
nand U14193 (N_14193,N_13850,N_13761);
nand U14194 (N_14194,N_13931,N_13758);
nand U14195 (N_14195,N_13860,N_13803);
xnor U14196 (N_14196,N_13990,N_13701);
xor U14197 (N_14197,N_13690,N_13772);
or U14198 (N_14198,N_13798,N_13723);
or U14199 (N_14199,N_13697,N_13894);
xnor U14200 (N_14200,N_13686,N_13927);
or U14201 (N_14201,N_13682,N_13659);
or U14202 (N_14202,N_13769,N_13936);
xor U14203 (N_14203,N_13979,N_13821);
and U14204 (N_14204,N_13825,N_13926);
xor U14205 (N_14205,N_13673,N_13804);
nor U14206 (N_14206,N_13965,N_13647);
and U14207 (N_14207,N_13681,N_13635);
nand U14208 (N_14208,N_13975,N_13776);
nor U14209 (N_14209,N_13707,N_13901);
nor U14210 (N_14210,N_13938,N_13690);
or U14211 (N_14211,N_13944,N_13763);
xor U14212 (N_14212,N_13679,N_13629);
or U14213 (N_14213,N_13771,N_13917);
nand U14214 (N_14214,N_13894,N_13992);
nand U14215 (N_14215,N_13798,N_13679);
nor U14216 (N_14216,N_13744,N_13963);
nand U14217 (N_14217,N_13705,N_13767);
xnor U14218 (N_14218,N_13757,N_13831);
nand U14219 (N_14219,N_13816,N_13603);
nor U14220 (N_14220,N_13754,N_13923);
xnor U14221 (N_14221,N_13902,N_13806);
and U14222 (N_14222,N_13987,N_13649);
and U14223 (N_14223,N_13640,N_13977);
or U14224 (N_14224,N_13879,N_13777);
or U14225 (N_14225,N_13885,N_13747);
nor U14226 (N_14226,N_13940,N_13879);
nor U14227 (N_14227,N_13969,N_13860);
nand U14228 (N_14228,N_13679,N_13640);
nand U14229 (N_14229,N_13906,N_13629);
nand U14230 (N_14230,N_13700,N_13989);
or U14231 (N_14231,N_13845,N_13695);
xnor U14232 (N_14232,N_13691,N_13762);
or U14233 (N_14233,N_13655,N_13909);
or U14234 (N_14234,N_13932,N_13843);
nand U14235 (N_14235,N_13875,N_13956);
nor U14236 (N_14236,N_13666,N_13737);
nor U14237 (N_14237,N_13946,N_13649);
nand U14238 (N_14238,N_13876,N_13752);
nand U14239 (N_14239,N_13987,N_13711);
nand U14240 (N_14240,N_13980,N_13917);
or U14241 (N_14241,N_13615,N_13681);
and U14242 (N_14242,N_13632,N_13677);
nor U14243 (N_14243,N_13665,N_13756);
or U14244 (N_14244,N_13964,N_13767);
or U14245 (N_14245,N_13715,N_13854);
nor U14246 (N_14246,N_13882,N_13862);
nor U14247 (N_14247,N_13771,N_13969);
nor U14248 (N_14248,N_13801,N_13927);
nor U14249 (N_14249,N_13835,N_13967);
nand U14250 (N_14250,N_13979,N_13773);
nand U14251 (N_14251,N_13901,N_13957);
or U14252 (N_14252,N_13904,N_13609);
nor U14253 (N_14253,N_13985,N_13861);
nor U14254 (N_14254,N_13657,N_13785);
or U14255 (N_14255,N_13800,N_13949);
nor U14256 (N_14256,N_13621,N_13607);
nor U14257 (N_14257,N_13618,N_13968);
and U14258 (N_14258,N_13787,N_13759);
or U14259 (N_14259,N_13616,N_13714);
xor U14260 (N_14260,N_13860,N_13852);
nand U14261 (N_14261,N_13904,N_13885);
or U14262 (N_14262,N_13785,N_13927);
xor U14263 (N_14263,N_13663,N_13668);
and U14264 (N_14264,N_13694,N_13726);
xor U14265 (N_14265,N_13672,N_13916);
or U14266 (N_14266,N_13943,N_13636);
or U14267 (N_14267,N_13852,N_13979);
xnor U14268 (N_14268,N_13869,N_13814);
or U14269 (N_14269,N_13828,N_13902);
or U14270 (N_14270,N_13823,N_13942);
and U14271 (N_14271,N_13787,N_13782);
nand U14272 (N_14272,N_13915,N_13700);
nand U14273 (N_14273,N_13682,N_13940);
nor U14274 (N_14274,N_13983,N_13790);
and U14275 (N_14275,N_13640,N_13723);
nand U14276 (N_14276,N_13616,N_13951);
nand U14277 (N_14277,N_13928,N_13629);
nor U14278 (N_14278,N_13635,N_13872);
and U14279 (N_14279,N_13979,N_13606);
nand U14280 (N_14280,N_13623,N_13897);
nand U14281 (N_14281,N_13851,N_13727);
nor U14282 (N_14282,N_13940,N_13854);
nand U14283 (N_14283,N_13638,N_13625);
and U14284 (N_14284,N_13697,N_13617);
or U14285 (N_14285,N_13888,N_13835);
nor U14286 (N_14286,N_13647,N_13683);
or U14287 (N_14287,N_13787,N_13801);
xnor U14288 (N_14288,N_13846,N_13937);
and U14289 (N_14289,N_13926,N_13883);
nand U14290 (N_14290,N_13826,N_13832);
xnor U14291 (N_14291,N_13725,N_13894);
or U14292 (N_14292,N_13971,N_13748);
or U14293 (N_14293,N_13649,N_13613);
and U14294 (N_14294,N_13905,N_13913);
nand U14295 (N_14295,N_13753,N_13878);
nand U14296 (N_14296,N_13788,N_13621);
or U14297 (N_14297,N_13741,N_13896);
xnor U14298 (N_14298,N_13762,N_13688);
nand U14299 (N_14299,N_13975,N_13971);
or U14300 (N_14300,N_13740,N_13675);
nor U14301 (N_14301,N_13704,N_13966);
nand U14302 (N_14302,N_13688,N_13657);
xnor U14303 (N_14303,N_13669,N_13821);
nor U14304 (N_14304,N_13866,N_13613);
nand U14305 (N_14305,N_13801,N_13793);
and U14306 (N_14306,N_13692,N_13729);
nor U14307 (N_14307,N_13745,N_13779);
nand U14308 (N_14308,N_13691,N_13707);
xor U14309 (N_14309,N_13834,N_13881);
xnor U14310 (N_14310,N_13681,N_13852);
nand U14311 (N_14311,N_13922,N_13693);
and U14312 (N_14312,N_13947,N_13808);
or U14313 (N_14313,N_13750,N_13819);
or U14314 (N_14314,N_13776,N_13858);
nor U14315 (N_14315,N_13814,N_13772);
nor U14316 (N_14316,N_13721,N_13692);
and U14317 (N_14317,N_13746,N_13802);
nor U14318 (N_14318,N_13670,N_13847);
nand U14319 (N_14319,N_13852,N_13842);
xnor U14320 (N_14320,N_13739,N_13864);
nand U14321 (N_14321,N_13665,N_13993);
nor U14322 (N_14322,N_13914,N_13822);
nor U14323 (N_14323,N_13621,N_13918);
or U14324 (N_14324,N_13760,N_13959);
and U14325 (N_14325,N_13789,N_13920);
nand U14326 (N_14326,N_13630,N_13924);
nor U14327 (N_14327,N_13626,N_13628);
xnor U14328 (N_14328,N_13867,N_13775);
xor U14329 (N_14329,N_13960,N_13995);
nand U14330 (N_14330,N_13792,N_13947);
or U14331 (N_14331,N_13739,N_13860);
nand U14332 (N_14332,N_13801,N_13707);
xnor U14333 (N_14333,N_13847,N_13995);
nand U14334 (N_14334,N_13923,N_13727);
or U14335 (N_14335,N_13688,N_13783);
or U14336 (N_14336,N_13754,N_13926);
xnor U14337 (N_14337,N_13688,N_13950);
nand U14338 (N_14338,N_13999,N_13930);
nand U14339 (N_14339,N_13941,N_13889);
nand U14340 (N_14340,N_13777,N_13632);
xor U14341 (N_14341,N_13957,N_13948);
nor U14342 (N_14342,N_13993,N_13764);
and U14343 (N_14343,N_13976,N_13843);
or U14344 (N_14344,N_13988,N_13920);
xnor U14345 (N_14345,N_13884,N_13922);
and U14346 (N_14346,N_13809,N_13700);
or U14347 (N_14347,N_13969,N_13974);
or U14348 (N_14348,N_13737,N_13916);
nand U14349 (N_14349,N_13681,N_13994);
or U14350 (N_14350,N_13895,N_13932);
nor U14351 (N_14351,N_13923,N_13793);
and U14352 (N_14352,N_13682,N_13653);
nand U14353 (N_14353,N_13840,N_13657);
or U14354 (N_14354,N_13619,N_13897);
xnor U14355 (N_14355,N_13745,N_13957);
nand U14356 (N_14356,N_13892,N_13968);
nor U14357 (N_14357,N_13993,N_13728);
and U14358 (N_14358,N_13636,N_13965);
nand U14359 (N_14359,N_13865,N_13903);
nand U14360 (N_14360,N_13742,N_13711);
and U14361 (N_14361,N_13822,N_13694);
and U14362 (N_14362,N_13682,N_13660);
or U14363 (N_14363,N_13857,N_13979);
nand U14364 (N_14364,N_13629,N_13953);
and U14365 (N_14365,N_13636,N_13877);
or U14366 (N_14366,N_13717,N_13734);
nor U14367 (N_14367,N_13671,N_13753);
and U14368 (N_14368,N_13681,N_13803);
and U14369 (N_14369,N_13786,N_13777);
nand U14370 (N_14370,N_13606,N_13641);
nor U14371 (N_14371,N_13909,N_13830);
or U14372 (N_14372,N_13992,N_13939);
or U14373 (N_14373,N_13947,N_13801);
xnor U14374 (N_14374,N_13729,N_13795);
and U14375 (N_14375,N_13806,N_13636);
and U14376 (N_14376,N_13895,N_13751);
nor U14377 (N_14377,N_13768,N_13749);
nor U14378 (N_14378,N_13990,N_13751);
xor U14379 (N_14379,N_13611,N_13635);
nor U14380 (N_14380,N_13982,N_13932);
or U14381 (N_14381,N_13794,N_13603);
xnor U14382 (N_14382,N_13731,N_13744);
nand U14383 (N_14383,N_13719,N_13721);
or U14384 (N_14384,N_13842,N_13779);
and U14385 (N_14385,N_13938,N_13722);
or U14386 (N_14386,N_13850,N_13627);
nor U14387 (N_14387,N_13841,N_13706);
or U14388 (N_14388,N_13757,N_13741);
nand U14389 (N_14389,N_13667,N_13860);
nand U14390 (N_14390,N_13616,N_13970);
and U14391 (N_14391,N_13937,N_13638);
xor U14392 (N_14392,N_13718,N_13852);
or U14393 (N_14393,N_13970,N_13830);
nand U14394 (N_14394,N_13826,N_13771);
nor U14395 (N_14395,N_13992,N_13869);
nor U14396 (N_14396,N_13795,N_13871);
nand U14397 (N_14397,N_13741,N_13930);
or U14398 (N_14398,N_13852,N_13618);
or U14399 (N_14399,N_13649,N_13627);
xor U14400 (N_14400,N_14289,N_14095);
and U14401 (N_14401,N_14012,N_14317);
nor U14402 (N_14402,N_14043,N_14158);
xnor U14403 (N_14403,N_14050,N_14321);
nor U14404 (N_14404,N_14135,N_14282);
xnor U14405 (N_14405,N_14151,N_14361);
xor U14406 (N_14406,N_14199,N_14328);
and U14407 (N_14407,N_14075,N_14174);
and U14408 (N_14408,N_14014,N_14244);
nor U14409 (N_14409,N_14362,N_14077);
nand U14410 (N_14410,N_14190,N_14278);
and U14411 (N_14411,N_14291,N_14106);
nor U14412 (N_14412,N_14103,N_14006);
xnor U14413 (N_14413,N_14170,N_14379);
nor U14414 (N_14414,N_14316,N_14257);
or U14415 (N_14415,N_14118,N_14082);
or U14416 (N_14416,N_14159,N_14131);
nor U14417 (N_14417,N_14013,N_14210);
nand U14418 (N_14418,N_14280,N_14035);
nand U14419 (N_14419,N_14290,N_14065);
or U14420 (N_14420,N_14320,N_14089);
and U14421 (N_14421,N_14234,N_14222);
and U14422 (N_14422,N_14051,N_14236);
nand U14423 (N_14423,N_14059,N_14139);
nor U14424 (N_14424,N_14128,N_14143);
xnor U14425 (N_14425,N_14045,N_14134);
nor U14426 (N_14426,N_14125,N_14355);
or U14427 (N_14427,N_14345,N_14020);
xnor U14428 (N_14428,N_14096,N_14391);
or U14429 (N_14429,N_14097,N_14010);
and U14430 (N_14430,N_14274,N_14252);
and U14431 (N_14431,N_14153,N_14197);
nor U14432 (N_14432,N_14281,N_14196);
or U14433 (N_14433,N_14249,N_14230);
or U14434 (N_14434,N_14287,N_14394);
or U14435 (N_14435,N_14092,N_14276);
xor U14436 (N_14436,N_14209,N_14144);
and U14437 (N_14437,N_14195,N_14137);
and U14438 (N_14438,N_14397,N_14114);
nor U14439 (N_14439,N_14046,N_14069);
nand U14440 (N_14440,N_14398,N_14079);
or U14441 (N_14441,N_14288,N_14017);
nand U14442 (N_14442,N_14007,N_14327);
or U14443 (N_14443,N_14387,N_14066);
nand U14444 (N_14444,N_14176,N_14030);
or U14445 (N_14445,N_14200,N_14325);
xor U14446 (N_14446,N_14295,N_14009);
and U14447 (N_14447,N_14213,N_14123);
xor U14448 (N_14448,N_14293,N_14299);
and U14449 (N_14449,N_14229,N_14392);
and U14450 (N_14450,N_14330,N_14247);
nand U14451 (N_14451,N_14270,N_14022);
xnor U14452 (N_14452,N_14036,N_14313);
nor U14453 (N_14453,N_14306,N_14120);
and U14454 (N_14454,N_14370,N_14347);
nor U14455 (N_14455,N_14127,N_14116);
or U14456 (N_14456,N_14322,N_14083);
xor U14457 (N_14457,N_14262,N_14148);
xor U14458 (N_14458,N_14207,N_14349);
or U14459 (N_14459,N_14285,N_14292);
nor U14460 (N_14460,N_14179,N_14169);
nor U14461 (N_14461,N_14150,N_14231);
nand U14462 (N_14462,N_14084,N_14253);
or U14463 (N_14463,N_14216,N_14039);
nand U14464 (N_14464,N_14351,N_14189);
xnor U14465 (N_14465,N_14356,N_14042);
or U14466 (N_14466,N_14315,N_14178);
nand U14467 (N_14467,N_14377,N_14246);
nor U14468 (N_14468,N_14220,N_14121);
and U14469 (N_14469,N_14133,N_14076);
nand U14470 (N_14470,N_14323,N_14165);
and U14471 (N_14471,N_14388,N_14164);
nor U14472 (N_14472,N_14071,N_14254);
and U14473 (N_14473,N_14367,N_14272);
and U14474 (N_14474,N_14354,N_14044);
or U14475 (N_14475,N_14261,N_14058);
and U14476 (N_14476,N_14368,N_14091);
xnor U14477 (N_14477,N_14300,N_14359);
xnor U14478 (N_14478,N_14141,N_14226);
and U14479 (N_14479,N_14168,N_14228);
xor U14480 (N_14480,N_14334,N_14348);
or U14481 (N_14481,N_14344,N_14205);
nand U14482 (N_14482,N_14073,N_14049);
nor U14483 (N_14483,N_14310,N_14237);
and U14484 (N_14484,N_14111,N_14286);
or U14485 (N_14485,N_14372,N_14341);
and U14486 (N_14486,N_14033,N_14256);
nand U14487 (N_14487,N_14284,N_14031);
or U14488 (N_14488,N_14000,N_14395);
or U14489 (N_14489,N_14233,N_14085);
or U14490 (N_14490,N_14019,N_14221);
xor U14491 (N_14491,N_14166,N_14072);
xnor U14492 (N_14492,N_14070,N_14094);
or U14493 (N_14493,N_14005,N_14309);
nor U14494 (N_14494,N_14206,N_14181);
or U14495 (N_14495,N_14198,N_14382);
xor U14496 (N_14496,N_14204,N_14396);
nand U14497 (N_14497,N_14177,N_14308);
nand U14498 (N_14498,N_14173,N_14245);
nand U14499 (N_14499,N_14260,N_14343);
nor U14500 (N_14500,N_14023,N_14279);
and U14501 (N_14501,N_14264,N_14093);
or U14502 (N_14502,N_14182,N_14312);
nor U14503 (N_14503,N_14275,N_14336);
nand U14504 (N_14504,N_14203,N_14018);
xor U14505 (N_14505,N_14329,N_14064);
or U14506 (N_14506,N_14365,N_14025);
and U14507 (N_14507,N_14194,N_14269);
and U14508 (N_14508,N_14294,N_14202);
nand U14509 (N_14509,N_14184,N_14188);
or U14510 (N_14510,N_14183,N_14218);
xnor U14511 (N_14511,N_14004,N_14326);
and U14512 (N_14512,N_14371,N_14048);
or U14513 (N_14513,N_14376,N_14227);
nor U14514 (N_14514,N_14386,N_14378);
xor U14515 (N_14515,N_14283,N_14113);
nand U14516 (N_14516,N_14138,N_14307);
nor U14517 (N_14517,N_14258,N_14167);
and U14518 (N_14518,N_14298,N_14238);
nand U14519 (N_14519,N_14201,N_14160);
nor U14520 (N_14520,N_14185,N_14350);
or U14521 (N_14521,N_14132,N_14303);
and U14522 (N_14522,N_14055,N_14029);
xnor U14523 (N_14523,N_14024,N_14215);
nor U14524 (N_14524,N_14339,N_14399);
nand U14525 (N_14525,N_14109,N_14380);
xor U14526 (N_14526,N_14053,N_14068);
xor U14527 (N_14527,N_14224,N_14175);
nand U14528 (N_14528,N_14149,N_14157);
xnor U14529 (N_14529,N_14302,N_14373);
nand U14530 (N_14530,N_14074,N_14105);
xor U14531 (N_14531,N_14232,N_14266);
nor U14532 (N_14532,N_14271,N_14001);
and U14533 (N_14533,N_14104,N_14235);
nor U14534 (N_14534,N_14110,N_14061);
xor U14535 (N_14535,N_14021,N_14156);
nand U14536 (N_14536,N_14129,N_14027);
and U14537 (N_14537,N_14364,N_14219);
xnor U14538 (N_14538,N_14180,N_14047);
xnor U14539 (N_14539,N_14062,N_14360);
nor U14540 (N_14540,N_14263,N_14154);
nor U14541 (N_14541,N_14273,N_14214);
or U14542 (N_14542,N_14028,N_14060);
and U14543 (N_14543,N_14080,N_14057);
nand U14544 (N_14544,N_14117,N_14081);
and U14545 (N_14545,N_14342,N_14225);
xor U14546 (N_14546,N_14037,N_14155);
nor U14547 (N_14547,N_14086,N_14034);
nor U14548 (N_14548,N_14337,N_14305);
xnor U14549 (N_14549,N_14171,N_14340);
nor U14550 (N_14550,N_14357,N_14338);
and U14551 (N_14551,N_14374,N_14248);
or U14552 (N_14552,N_14239,N_14078);
nor U14553 (N_14553,N_14040,N_14332);
nand U14554 (N_14554,N_14100,N_14217);
nand U14555 (N_14555,N_14318,N_14152);
nor U14556 (N_14556,N_14384,N_14162);
and U14557 (N_14557,N_14041,N_14242);
and U14558 (N_14558,N_14375,N_14311);
xor U14559 (N_14559,N_14383,N_14146);
nor U14560 (N_14560,N_14193,N_14032);
and U14561 (N_14561,N_14268,N_14314);
or U14562 (N_14562,N_14277,N_14352);
xor U14563 (N_14563,N_14102,N_14296);
nand U14564 (N_14564,N_14147,N_14163);
nor U14565 (N_14565,N_14124,N_14107);
nand U14566 (N_14566,N_14385,N_14015);
or U14567 (N_14567,N_14122,N_14267);
xor U14568 (N_14568,N_14016,N_14088);
nor U14569 (N_14569,N_14297,N_14063);
nand U14570 (N_14570,N_14067,N_14301);
and U14571 (N_14571,N_14389,N_14208);
and U14572 (N_14572,N_14191,N_14363);
nor U14573 (N_14573,N_14393,N_14142);
xnor U14574 (N_14574,N_14026,N_14108);
or U14575 (N_14575,N_14240,N_14319);
xnor U14576 (N_14576,N_14101,N_14335);
nor U14577 (N_14577,N_14098,N_14366);
nand U14578 (N_14578,N_14243,N_14038);
xor U14579 (N_14579,N_14251,N_14003);
and U14580 (N_14580,N_14390,N_14172);
or U14581 (N_14581,N_14353,N_14346);
and U14582 (N_14582,N_14056,N_14119);
and U14583 (N_14583,N_14186,N_14008);
xor U14584 (N_14584,N_14331,N_14011);
and U14585 (N_14585,N_14324,N_14161);
xnor U14586 (N_14586,N_14136,N_14304);
nor U14587 (N_14587,N_14212,N_14087);
nor U14588 (N_14588,N_14187,N_14192);
xor U14589 (N_14589,N_14250,N_14145);
nor U14590 (N_14590,N_14223,N_14259);
xnor U14591 (N_14591,N_14211,N_14140);
nor U14592 (N_14592,N_14265,N_14002);
and U14593 (N_14593,N_14130,N_14255);
xnor U14594 (N_14594,N_14333,N_14090);
xnor U14595 (N_14595,N_14112,N_14099);
nor U14596 (N_14596,N_14241,N_14358);
xor U14597 (N_14597,N_14054,N_14126);
xor U14598 (N_14598,N_14052,N_14381);
or U14599 (N_14599,N_14369,N_14115);
or U14600 (N_14600,N_14143,N_14239);
xor U14601 (N_14601,N_14351,N_14285);
or U14602 (N_14602,N_14138,N_14257);
xor U14603 (N_14603,N_14164,N_14303);
or U14604 (N_14604,N_14021,N_14328);
xnor U14605 (N_14605,N_14248,N_14086);
or U14606 (N_14606,N_14346,N_14108);
nor U14607 (N_14607,N_14050,N_14054);
and U14608 (N_14608,N_14100,N_14320);
xor U14609 (N_14609,N_14115,N_14291);
nor U14610 (N_14610,N_14046,N_14250);
nor U14611 (N_14611,N_14050,N_14193);
xnor U14612 (N_14612,N_14072,N_14057);
or U14613 (N_14613,N_14158,N_14076);
or U14614 (N_14614,N_14397,N_14337);
xor U14615 (N_14615,N_14061,N_14187);
and U14616 (N_14616,N_14383,N_14283);
nor U14617 (N_14617,N_14320,N_14362);
xor U14618 (N_14618,N_14362,N_14248);
xor U14619 (N_14619,N_14390,N_14211);
and U14620 (N_14620,N_14157,N_14095);
or U14621 (N_14621,N_14036,N_14255);
nor U14622 (N_14622,N_14114,N_14169);
nor U14623 (N_14623,N_14009,N_14185);
nand U14624 (N_14624,N_14235,N_14345);
or U14625 (N_14625,N_14295,N_14003);
and U14626 (N_14626,N_14247,N_14015);
and U14627 (N_14627,N_14332,N_14150);
nor U14628 (N_14628,N_14183,N_14307);
or U14629 (N_14629,N_14109,N_14087);
nor U14630 (N_14630,N_14380,N_14300);
xor U14631 (N_14631,N_14058,N_14299);
xor U14632 (N_14632,N_14139,N_14132);
or U14633 (N_14633,N_14040,N_14165);
or U14634 (N_14634,N_14002,N_14309);
xor U14635 (N_14635,N_14204,N_14186);
nor U14636 (N_14636,N_14173,N_14263);
nand U14637 (N_14637,N_14115,N_14322);
nor U14638 (N_14638,N_14179,N_14062);
nand U14639 (N_14639,N_14162,N_14108);
nor U14640 (N_14640,N_14156,N_14295);
nand U14641 (N_14641,N_14098,N_14190);
or U14642 (N_14642,N_14092,N_14148);
or U14643 (N_14643,N_14349,N_14223);
and U14644 (N_14644,N_14005,N_14064);
or U14645 (N_14645,N_14177,N_14038);
nand U14646 (N_14646,N_14038,N_14189);
xor U14647 (N_14647,N_14170,N_14237);
nor U14648 (N_14648,N_14135,N_14189);
or U14649 (N_14649,N_14053,N_14285);
or U14650 (N_14650,N_14309,N_14111);
and U14651 (N_14651,N_14227,N_14208);
nor U14652 (N_14652,N_14260,N_14232);
nand U14653 (N_14653,N_14095,N_14306);
nand U14654 (N_14654,N_14128,N_14346);
nor U14655 (N_14655,N_14159,N_14230);
nand U14656 (N_14656,N_14128,N_14259);
and U14657 (N_14657,N_14012,N_14360);
and U14658 (N_14658,N_14324,N_14000);
nand U14659 (N_14659,N_14142,N_14119);
xor U14660 (N_14660,N_14291,N_14135);
nand U14661 (N_14661,N_14365,N_14238);
xor U14662 (N_14662,N_14367,N_14109);
nand U14663 (N_14663,N_14266,N_14234);
nand U14664 (N_14664,N_14142,N_14383);
xor U14665 (N_14665,N_14143,N_14338);
and U14666 (N_14666,N_14170,N_14279);
and U14667 (N_14667,N_14010,N_14150);
nor U14668 (N_14668,N_14274,N_14061);
and U14669 (N_14669,N_14281,N_14060);
nand U14670 (N_14670,N_14343,N_14327);
and U14671 (N_14671,N_14057,N_14083);
xnor U14672 (N_14672,N_14336,N_14089);
xnor U14673 (N_14673,N_14077,N_14225);
or U14674 (N_14674,N_14380,N_14085);
xnor U14675 (N_14675,N_14350,N_14307);
nand U14676 (N_14676,N_14315,N_14074);
and U14677 (N_14677,N_14198,N_14304);
xor U14678 (N_14678,N_14369,N_14227);
nor U14679 (N_14679,N_14066,N_14296);
or U14680 (N_14680,N_14353,N_14236);
and U14681 (N_14681,N_14079,N_14051);
and U14682 (N_14682,N_14250,N_14298);
or U14683 (N_14683,N_14321,N_14240);
and U14684 (N_14684,N_14379,N_14083);
and U14685 (N_14685,N_14123,N_14291);
and U14686 (N_14686,N_14015,N_14226);
nand U14687 (N_14687,N_14180,N_14386);
nand U14688 (N_14688,N_14342,N_14223);
and U14689 (N_14689,N_14312,N_14393);
xor U14690 (N_14690,N_14287,N_14064);
nand U14691 (N_14691,N_14289,N_14246);
or U14692 (N_14692,N_14104,N_14383);
or U14693 (N_14693,N_14136,N_14143);
nand U14694 (N_14694,N_14225,N_14296);
xnor U14695 (N_14695,N_14329,N_14028);
or U14696 (N_14696,N_14321,N_14332);
or U14697 (N_14697,N_14148,N_14337);
nor U14698 (N_14698,N_14216,N_14241);
nor U14699 (N_14699,N_14241,N_14302);
or U14700 (N_14700,N_14291,N_14124);
xor U14701 (N_14701,N_14393,N_14395);
nand U14702 (N_14702,N_14166,N_14113);
or U14703 (N_14703,N_14268,N_14169);
nand U14704 (N_14704,N_14110,N_14240);
xnor U14705 (N_14705,N_14032,N_14094);
nand U14706 (N_14706,N_14233,N_14198);
nand U14707 (N_14707,N_14266,N_14386);
nand U14708 (N_14708,N_14115,N_14071);
nand U14709 (N_14709,N_14038,N_14320);
xnor U14710 (N_14710,N_14034,N_14205);
nor U14711 (N_14711,N_14211,N_14350);
and U14712 (N_14712,N_14195,N_14053);
and U14713 (N_14713,N_14246,N_14112);
and U14714 (N_14714,N_14134,N_14310);
nor U14715 (N_14715,N_14180,N_14286);
and U14716 (N_14716,N_14075,N_14100);
or U14717 (N_14717,N_14173,N_14382);
xnor U14718 (N_14718,N_14394,N_14220);
or U14719 (N_14719,N_14129,N_14118);
or U14720 (N_14720,N_14392,N_14239);
xnor U14721 (N_14721,N_14376,N_14213);
or U14722 (N_14722,N_14075,N_14161);
xor U14723 (N_14723,N_14330,N_14097);
nand U14724 (N_14724,N_14036,N_14035);
xnor U14725 (N_14725,N_14329,N_14274);
nand U14726 (N_14726,N_14211,N_14356);
or U14727 (N_14727,N_14345,N_14388);
xnor U14728 (N_14728,N_14073,N_14364);
xor U14729 (N_14729,N_14303,N_14208);
xor U14730 (N_14730,N_14082,N_14077);
nor U14731 (N_14731,N_14294,N_14049);
nand U14732 (N_14732,N_14341,N_14220);
xnor U14733 (N_14733,N_14079,N_14028);
and U14734 (N_14734,N_14273,N_14349);
xor U14735 (N_14735,N_14055,N_14298);
xor U14736 (N_14736,N_14169,N_14304);
and U14737 (N_14737,N_14296,N_14270);
or U14738 (N_14738,N_14210,N_14002);
xnor U14739 (N_14739,N_14201,N_14333);
nand U14740 (N_14740,N_14050,N_14060);
or U14741 (N_14741,N_14375,N_14396);
nand U14742 (N_14742,N_14336,N_14375);
nand U14743 (N_14743,N_14054,N_14063);
nor U14744 (N_14744,N_14138,N_14070);
xnor U14745 (N_14745,N_14324,N_14373);
or U14746 (N_14746,N_14062,N_14030);
xnor U14747 (N_14747,N_14189,N_14268);
and U14748 (N_14748,N_14206,N_14159);
nor U14749 (N_14749,N_14200,N_14105);
nor U14750 (N_14750,N_14131,N_14196);
or U14751 (N_14751,N_14305,N_14037);
and U14752 (N_14752,N_14151,N_14039);
or U14753 (N_14753,N_14061,N_14004);
nand U14754 (N_14754,N_14165,N_14186);
nor U14755 (N_14755,N_14284,N_14329);
or U14756 (N_14756,N_14214,N_14364);
nand U14757 (N_14757,N_14188,N_14309);
and U14758 (N_14758,N_14305,N_14359);
and U14759 (N_14759,N_14073,N_14230);
nand U14760 (N_14760,N_14354,N_14142);
and U14761 (N_14761,N_14115,N_14143);
or U14762 (N_14762,N_14266,N_14230);
xor U14763 (N_14763,N_14294,N_14066);
or U14764 (N_14764,N_14151,N_14154);
nor U14765 (N_14765,N_14220,N_14325);
and U14766 (N_14766,N_14354,N_14371);
or U14767 (N_14767,N_14309,N_14169);
nand U14768 (N_14768,N_14093,N_14087);
nor U14769 (N_14769,N_14296,N_14261);
and U14770 (N_14770,N_14016,N_14290);
nand U14771 (N_14771,N_14049,N_14332);
xnor U14772 (N_14772,N_14156,N_14002);
nor U14773 (N_14773,N_14374,N_14123);
and U14774 (N_14774,N_14032,N_14188);
or U14775 (N_14775,N_14361,N_14137);
nor U14776 (N_14776,N_14092,N_14081);
xnor U14777 (N_14777,N_14296,N_14344);
xor U14778 (N_14778,N_14304,N_14178);
nand U14779 (N_14779,N_14182,N_14052);
and U14780 (N_14780,N_14272,N_14390);
and U14781 (N_14781,N_14308,N_14321);
nand U14782 (N_14782,N_14195,N_14083);
xnor U14783 (N_14783,N_14034,N_14074);
or U14784 (N_14784,N_14156,N_14214);
and U14785 (N_14785,N_14186,N_14223);
nor U14786 (N_14786,N_14053,N_14352);
nor U14787 (N_14787,N_14163,N_14082);
or U14788 (N_14788,N_14097,N_14326);
nor U14789 (N_14789,N_14199,N_14039);
nand U14790 (N_14790,N_14289,N_14082);
nand U14791 (N_14791,N_14134,N_14118);
nor U14792 (N_14792,N_14001,N_14197);
or U14793 (N_14793,N_14263,N_14157);
xor U14794 (N_14794,N_14050,N_14077);
xor U14795 (N_14795,N_14295,N_14292);
xor U14796 (N_14796,N_14368,N_14363);
and U14797 (N_14797,N_14344,N_14081);
nand U14798 (N_14798,N_14387,N_14215);
and U14799 (N_14799,N_14309,N_14319);
and U14800 (N_14800,N_14680,N_14675);
xor U14801 (N_14801,N_14782,N_14747);
nand U14802 (N_14802,N_14623,N_14505);
or U14803 (N_14803,N_14535,N_14524);
or U14804 (N_14804,N_14727,N_14784);
nor U14805 (N_14805,N_14530,N_14723);
nor U14806 (N_14806,N_14604,N_14654);
nor U14807 (N_14807,N_14421,N_14649);
nor U14808 (N_14808,N_14774,N_14650);
or U14809 (N_14809,N_14423,N_14753);
xor U14810 (N_14810,N_14508,N_14708);
and U14811 (N_14811,N_14757,N_14667);
nor U14812 (N_14812,N_14547,N_14633);
nand U14813 (N_14813,N_14588,N_14732);
and U14814 (N_14814,N_14744,N_14652);
nor U14815 (N_14815,N_14595,N_14714);
nand U14816 (N_14816,N_14578,N_14412);
nand U14817 (N_14817,N_14789,N_14448);
nor U14818 (N_14818,N_14711,N_14529);
nor U14819 (N_14819,N_14596,N_14730);
nand U14820 (N_14820,N_14587,N_14481);
nor U14821 (N_14821,N_14562,N_14779);
nor U14822 (N_14822,N_14632,N_14441);
xor U14823 (N_14823,N_14405,N_14646);
nor U14824 (N_14824,N_14540,N_14717);
nor U14825 (N_14825,N_14798,N_14579);
nand U14826 (N_14826,N_14741,N_14748);
xor U14827 (N_14827,N_14743,N_14444);
nand U14828 (N_14828,N_14491,N_14778);
or U14829 (N_14829,N_14581,N_14611);
xnor U14830 (N_14830,N_14486,N_14790);
xnor U14831 (N_14831,N_14400,N_14706);
or U14832 (N_14832,N_14752,N_14435);
or U14833 (N_14833,N_14443,N_14552);
nor U14834 (N_14834,N_14635,N_14746);
and U14835 (N_14835,N_14673,N_14734);
and U14836 (N_14836,N_14644,N_14493);
nand U14837 (N_14837,N_14773,N_14715);
nor U14838 (N_14838,N_14454,N_14565);
nand U14839 (N_14839,N_14541,N_14630);
or U14840 (N_14840,N_14425,N_14519);
or U14841 (N_14841,N_14620,N_14522);
and U14842 (N_14842,N_14659,N_14781);
and U14843 (N_14843,N_14553,N_14771);
xor U14844 (N_14844,N_14763,N_14525);
nand U14845 (N_14845,N_14564,N_14655);
or U14846 (N_14846,N_14556,N_14629);
and U14847 (N_14847,N_14512,N_14648);
or U14848 (N_14848,N_14584,N_14707);
xor U14849 (N_14849,N_14709,N_14472);
nor U14850 (N_14850,N_14726,N_14488);
nor U14851 (N_14851,N_14554,N_14456);
nor U14852 (N_14852,N_14517,N_14690);
nand U14853 (N_14853,N_14770,N_14483);
xor U14854 (N_14854,N_14526,N_14582);
or U14855 (N_14855,N_14450,N_14637);
nor U14856 (N_14856,N_14634,N_14506);
nand U14857 (N_14857,N_14721,N_14767);
or U14858 (N_14858,N_14704,N_14686);
and U14859 (N_14859,N_14432,N_14700);
nor U14860 (N_14860,N_14499,N_14760);
nand U14861 (N_14861,N_14406,N_14437);
and U14862 (N_14862,N_14403,N_14674);
xnor U14863 (N_14863,N_14568,N_14736);
or U14864 (N_14864,N_14557,N_14431);
or U14865 (N_14865,N_14788,N_14698);
nand U14866 (N_14866,N_14719,N_14785);
xnor U14867 (N_14867,N_14533,N_14549);
xor U14868 (N_14868,N_14497,N_14621);
nor U14869 (N_14869,N_14551,N_14609);
nand U14870 (N_14870,N_14641,N_14509);
and U14871 (N_14871,N_14795,N_14538);
and U14872 (N_14872,N_14695,N_14591);
or U14873 (N_14873,N_14636,N_14484);
and U14874 (N_14874,N_14415,N_14543);
nor U14875 (N_14875,N_14597,N_14567);
nor U14876 (N_14876,N_14663,N_14521);
or U14877 (N_14877,N_14451,N_14678);
nand U14878 (N_14878,N_14643,N_14657);
nand U14879 (N_14879,N_14610,N_14729);
nand U14880 (N_14880,N_14718,N_14534);
nor U14881 (N_14881,N_14761,N_14469);
nor U14882 (N_14882,N_14487,N_14658);
xor U14883 (N_14883,N_14485,N_14642);
nand U14884 (N_14884,N_14656,N_14703);
or U14885 (N_14885,N_14520,N_14699);
nand U14886 (N_14886,N_14601,N_14464);
nor U14887 (N_14887,N_14647,N_14513);
and U14888 (N_14888,N_14424,N_14574);
nand U14889 (N_14889,N_14527,N_14426);
and U14890 (N_14890,N_14797,N_14740);
and U14891 (N_14891,N_14720,N_14571);
and U14892 (N_14892,N_14780,N_14676);
nor U14893 (N_14893,N_14461,N_14672);
or U14894 (N_14894,N_14697,N_14766);
xnor U14895 (N_14895,N_14532,N_14544);
xor U14896 (N_14896,N_14615,N_14606);
nor U14897 (N_14897,N_14799,N_14762);
nand U14898 (N_14898,N_14572,N_14457);
nand U14899 (N_14899,N_14558,N_14434);
or U14900 (N_14900,N_14671,N_14537);
or U14901 (N_14901,N_14739,N_14787);
or U14902 (N_14902,N_14738,N_14545);
or U14903 (N_14903,N_14745,N_14477);
nor U14904 (N_14904,N_14542,N_14468);
nor U14905 (N_14905,N_14459,N_14617);
nand U14906 (N_14906,N_14580,N_14496);
and U14907 (N_14907,N_14705,N_14447);
or U14908 (N_14908,N_14577,N_14583);
xor U14909 (N_14909,N_14471,N_14589);
nor U14910 (N_14910,N_14414,N_14502);
or U14911 (N_14911,N_14613,N_14430);
nand U14912 (N_14912,N_14772,N_14474);
nand U14913 (N_14913,N_14501,N_14677);
and U14914 (N_14914,N_14482,N_14599);
or U14915 (N_14915,N_14751,N_14573);
nor U14916 (N_14916,N_14455,N_14476);
nor U14917 (N_14917,N_14440,N_14465);
and U14918 (N_14918,N_14687,N_14725);
xnor U14919 (N_14919,N_14645,N_14401);
and U14920 (N_14920,N_14664,N_14728);
nand U14921 (N_14921,N_14666,N_14764);
nor U14922 (N_14922,N_14592,N_14560);
and U14923 (N_14923,N_14724,N_14794);
nor U14924 (N_14924,N_14511,N_14570);
and U14925 (N_14925,N_14640,N_14460);
nor U14926 (N_14926,N_14416,N_14624);
and U14927 (N_14927,N_14507,N_14452);
nand U14928 (N_14928,N_14407,N_14593);
and U14929 (N_14929,N_14692,N_14576);
xnor U14930 (N_14930,N_14598,N_14514);
nor U14931 (N_14931,N_14463,N_14684);
nand U14932 (N_14932,N_14754,N_14622);
and U14933 (N_14933,N_14662,N_14608);
xnor U14934 (N_14934,N_14516,N_14660);
and U14935 (N_14935,N_14607,N_14548);
and U14936 (N_14936,N_14683,N_14427);
xor U14937 (N_14937,N_14561,N_14626);
or U14938 (N_14938,N_14433,N_14638);
nor U14939 (N_14939,N_14539,N_14759);
nor U14940 (N_14940,N_14470,N_14602);
nand U14941 (N_14941,N_14546,N_14563);
nor U14942 (N_14942,N_14689,N_14758);
nand U14943 (N_14943,N_14691,N_14682);
or U14944 (N_14944,N_14616,N_14793);
xor U14945 (N_14945,N_14438,N_14550);
xor U14946 (N_14946,N_14668,N_14419);
xor U14947 (N_14947,N_14429,N_14458);
and U14948 (N_14948,N_14742,N_14479);
and U14949 (N_14949,N_14409,N_14410);
and U14950 (N_14950,N_14504,N_14422);
or U14951 (N_14951,N_14614,N_14418);
nand U14952 (N_14952,N_14495,N_14478);
or U14953 (N_14953,N_14627,N_14590);
xnor U14954 (N_14954,N_14618,N_14518);
and U14955 (N_14955,N_14453,N_14737);
and U14956 (N_14956,N_14685,N_14777);
xnor U14957 (N_14957,N_14408,N_14681);
nor U14958 (N_14958,N_14467,N_14586);
nand U14959 (N_14959,N_14651,N_14769);
xor U14960 (N_14960,N_14569,N_14665);
or U14961 (N_14961,N_14442,N_14600);
nor U14962 (N_14962,N_14490,N_14439);
nand U14963 (N_14963,N_14765,N_14566);
and U14964 (N_14964,N_14515,N_14523);
xor U14965 (N_14965,N_14475,N_14555);
and U14966 (N_14966,N_14605,N_14559);
or U14967 (N_14967,N_14735,N_14701);
xnor U14968 (N_14968,N_14612,N_14411);
or U14969 (N_14969,N_14750,N_14449);
and U14970 (N_14970,N_14733,N_14404);
or U14971 (N_14971,N_14594,N_14628);
or U14972 (N_14972,N_14796,N_14462);
nand U14973 (N_14973,N_14653,N_14749);
nand U14974 (N_14974,N_14710,N_14669);
or U14975 (N_14975,N_14510,N_14436);
nor U14976 (N_14976,N_14473,N_14731);
and U14977 (N_14977,N_14791,N_14446);
xnor U14978 (N_14978,N_14445,N_14466);
nand U14979 (N_14979,N_14783,N_14402);
or U14980 (N_14980,N_14528,N_14531);
xor U14981 (N_14981,N_14498,N_14661);
and U14982 (N_14982,N_14755,N_14670);
xor U14983 (N_14983,N_14722,N_14756);
xor U14984 (N_14984,N_14679,N_14696);
nor U14985 (N_14985,N_14693,N_14702);
or U14986 (N_14986,N_14494,N_14536);
nor U14987 (N_14987,N_14713,N_14428);
xnor U14988 (N_14988,N_14503,N_14417);
xor U14989 (N_14989,N_14585,N_14768);
xnor U14990 (N_14990,N_14631,N_14625);
xnor U14991 (N_14991,N_14492,N_14480);
and U14992 (N_14992,N_14775,N_14489);
nand U14993 (N_14993,N_14694,N_14712);
xnor U14994 (N_14994,N_14716,N_14688);
and U14995 (N_14995,N_14792,N_14420);
nor U14996 (N_14996,N_14776,N_14786);
and U14997 (N_14997,N_14500,N_14575);
nand U14998 (N_14998,N_14603,N_14639);
nand U14999 (N_14999,N_14413,N_14619);
xnor U15000 (N_15000,N_14443,N_14660);
and U15001 (N_15001,N_14509,N_14720);
nand U15002 (N_15002,N_14632,N_14567);
xnor U15003 (N_15003,N_14783,N_14526);
nand U15004 (N_15004,N_14703,N_14546);
and U15005 (N_15005,N_14750,N_14719);
and U15006 (N_15006,N_14764,N_14563);
nand U15007 (N_15007,N_14587,N_14727);
nor U15008 (N_15008,N_14752,N_14671);
and U15009 (N_15009,N_14408,N_14634);
xor U15010 (N_15010,N_14781,N_14447);
or U15011 (N_15011,N_14618,N_14406);
xnor U15012 (N_15012,N_14708,N_14757);
xnor U15013 (N_15013,N_14506,N_14605);
nor U15014 (N_15014,N_14518,N_14776);
nor U15015 (N_15015,N_14593,N_14524);
and U15016 (N_15016,N_14776,N_14525);
nand U15017 (N_15017,N_14676,N_14788);
and U15018 (N_15018,N_14626,N_14598);
xor U15019 (N_15019,N_14658,N_14572);
nor U15020 (N_15020,N_14749,N_14608);
and U15021 (N_15021,N_14703,N_14615);
and U15022 (N_15022,N_14699,N_14457);
xor U15023 (N_15023,N_14530,N_14482);
nand U15024 (N_15024,N_14694,N_14622);
nor U15025 (N_15025,N_14756,N_14491);
or U15026 (N_15026,N_14567,N_14436);
xor U15027 (N_15027,N_14670,N_14400);
and U15028 (N_15028,N_14721,N_14567);
or U15029 (N_15029,N_14464,N_14439);
and U15030 (N_15030,N_14592,N_14435);
nor U15031 (N_15031,N_14426,N_14554);
nand U15032 (N_15032,N_14501,N_14675);
nor U15033 (N_15033,N_14717,N_14526);
nand U15034 (N_15034,N_14787,N_14696);
and U15035 (N_15035,N_14482,N_14650);
or U15036 (N_15036,N_14450,N_14788);
and U15037 (N_15037,N_14516,N_14571);
or U15038 (N_15038,N_14783,N_14652);
nor U15039 (N_15039,N_14646,N_14748);
xnor U15040 (N_15040,N_14467,N_14551);
or U15041 (N_15041,N_14570,N_14681);
or U15042 (N_15042,N_14524,N_14448);
nor U15043 (N_15043,N_14705,N_14763);
nor U15044 (N_15044,N_14759,N_14564);
and U15045 (N_15045,N_14787,N_14677);
and U15046 (N_15046,N_14460,N_14493);
or U15047 (N_15047,N_14677,N_14468);
nor U15048 (N_15048,N_14565,N_14668);
nand U15049 (N_15049,N_14532,N_14577);
xnor U15050 (N_15050,N_14486,N_14756);
nor U15051 (N_15051,N_14473,N_14522);
or U15052 (N_15052,N_14650,N_14434);
xor U15053 (N_15053,N_14625,N_14580);
nand U15054 (N_15054,N_14739,N_14558);
nor U15055 (N_15055,N_14774,N_14735);
or U15056 (N_15056,N_14463,N_14683);
nor U15057 (N_15057,N_14745,N_14535);
nor U15058 (N_15058,N_14748,N_14595);
or U15059 (N_15059,N_14617,N_14413);
nor U15060 (N_15060,N_14490,N_14524);
and U15061 (N_15061,N_14540,N_14406);
xnor U15062 (N_15062,N_14429,N_14685);
or U15063 (N_15063,N_14614,N_14667);
nor U15064 (N_15064,N_14508,N_14413);
or U15065 (N_15065,N_14581,N_14641);
nand U15066 (N_15066,N_14726,N_14463);
and U15067 (N_15067,N_14530,N_14545);
xor U15068 (N_15068,N_14661,N_14583);
nor U15069 (N_15069,N_14481,N_14443);
or U15070 (N_15070,N_14418,N_14452);
nand U15071 (N_15071,N_14408,N_14499);
nand U15072 (N_15072,N_14727,N_14480);
xnor U15073 (N_15073,N_14589,N_14568);
and U15074 (N_15074,N_14761,N_14684);
or U15075 (N_15075,N_14507,N_14656);
xnor U15076 (N_15076,N_14656,N_14486);
or U15077 (N_15077,N_14611,N_14707);
nand U15078 (N_15078,N_14406,N_14627);
or U15079 (N_15079,N_14662,N_14425);
xnor U15080 (N_15080,N_14480,N_14451);
nand U15081 (N_15081,N_14795,N_14649);
xor U15082 (N_15082,N_14478,N_14542);
nor U15083 (N_15083,N_14529,N_14612);
nor U15084 (N_15084,N_14706,N_14683);
nand U15085 (N_15085,N_14571,N_14760);
nor U15086 (N_15086,N_14719,N_14403);
nand U15087 (N_15087,N_14538,N_14652);
nand U15088 (N_15088,N_14705,N_14487);
nand U15089 (N_15089,N_14631,N_14533);
xnor U15090 (N_15090,N_14617,N_14411);
xor U15091 (N_15091,N_14595,N_14709);
or U15092 (N_15092,N_14504,N_14527);
xor U15093 (N_15093,N_14495,N_14628);
xor U15094 (N_15094,N_14716,N_14615);
xnor U15095 (N_15095,N_14619,N_14546);
nor U15096 (N_15096,N_14452,N_14406);
or U15097 (N_15097,N_14643,N_14519);
xnor U15098 (N_15098,N_14557,N_14476);
xnor U15099 (N_15099,N_14570,N_14638);
xor U15100 (N_15100,N_14473,N_14615);
and U15101 (N_15101,N_14497,N_14503);
or U15102 (N_15102,N_14486,N_14427);
or U15103 (N_15103,N_14612,N_14629);
xnor U15104 (N_15104,N_14491,N_14623);
nand U15105 (N_15105,N_14482,N_14654);
nand U15106 (N_15106,N_14480,N_14464);
xnor U15107 (N_15107,N_14606,N_14582);
and U15108 (N_15108,N_14439,N_14692);
nand U15109 (N_15109,N_14471,N_14675);
or U15110 (N_15110,N_14570,N_14515);
or U15111 (N_15111,N_14458,N_14754);
xnor U15112 (N_15112,N_14574,N_14784);
xnor U15113 (N_15113,N_14752,N_14615);
nand U15114 (N_15114,N_14414,N_14489);
and U15115 (N_15115,N_14684,N_14681);
or U15116 (N_15116,N_14438,N_14492);
or U15117 (N_15117,N_14689,N_14544);
nand U15118 (N_15118,N_14583,N_14598);
and U15119 (N_15119,N_14518,N_14778);
or U15120 (N_15120,N_14690,N_14402);
xor U15121 (N_15121,N_14428,N_14579);
nor U15122 (N_15122,N_14414,N_14572);
nand U15123 (N_15123,N_14581,N_14639);
or U15124 (N_15124,N_14661,N_14605);
xnor U15125 (N_15125,N_14707,N_14682);
and U15126 (N_15126,N_14407,N_14753);
nand U15127 (N_15127,N_14655,N_14635);
nand U15128 (N_15128,N_14647,N_14478);
and U15129 (N_15129,N_14571,N_14707);
nand U15130 (N_15130,N_14566,N_14486);
nor U15131 (N_15131,N_14629,N_14720);
xor U15132 (N_15132,N_14695,N_14594);
nand U15133 (N_15133,N_14751,N_14532);
or U15134 (N_15134,N_14492,N_14518);
or U15135 (N_15135,N_14487,N_14688);
or U15136 (N_15136,N_14708,N_14526);
nor U15137 (N_15137,N_14574,N_14514);
nor U15138 (N_15138,N_14607,N_14474);
nor U15139 (N_15139,N_14689,N_14561);
nor U15140 (N_15140,N_14528,N_14717);
and U15141 (N_15141,N_14573,N_14659);
nand U15142 (N_15142,N_14790,N_14574);
and U15143 (N_15143,N_14571,N_14415);
nand U15144 (N_15144,N_14462,N_14463);
and U15145 (N_15145,N_14600,N_14460);
nor U15146 (N_15146,N_14714,N_14572);
or U15147 (N_15147,N_14503,N_14594);
xor U15148 (N_15148,N_14453,N_14414);
nor U15149 (N_15149,N_14695,N_14546);
nor U15150 (N_15150,N_14624,N_14635);
nor U15151 (N_15151,N_14797,N_14656);
and U15152 (N_15152,N_14711,N_14412);
nand U15153 (N_15153,N_14471,N_14409);
or U15154 (N_15154,N_14662,N_14402);
xnor U15155 (N_15155,N_14609,N_14723);
xor U15156 (N_15156,N_14784,N_14549);
and U15157 (N_15157,N_14695,N_14525);
nor U15158 (N_15158,N_14534,N_14755);
and U15159 (N_15159,N_14416,N_14467);
nor U15160 (N_15160,N_14714,N_14503);
nand U15161 (N_15161,N_14688,N_14401);
nand U15162 (N_15162,N_14419,N_14463);
nand U15163 (N_15163,N_14739,N_14618);
nor U15164 (N_15164,N_14477,N_14635);
or U15165 (N_15165,N_14632,N_14443);
nor U15166 (N_15166,N_14692,N_14724);
xor U15167 (N_15167,N_14656,N_14669);
nand U15168 (N_15168,N_14493,N_14465);
and U15169 (N_15169,N_14528,N_14643);
and U15170 (N_15170,N_14585,N_14783);
nor U15171 (N_15171,N_14751,N_14567);
xor U15172 (N_15172,N_14521,N_14715);
xor U15173 (N_15173,N_14556,N_14765);
xor U15174 (N_15174,N_14793,N_14482);
and U15175 (N_15175,N_14582,N_14439);
xnor U15176 (N_15176,N_14524,N_14564);
and U15177 (N_15177,N_14484,N_14762);
xnor U15178 (N_15178,N_14758,N_14643);
and U15179 (N_15179,N_14677,N_14593);
and U15180 (N_15180,N_14602,N_14444);
nor U15181 (N_15181,N_14505,N_14636);
or U15182 (N_15182,N_14476,N_14678);
or U15183 (N_15183,N_14573,N_14417);
nand U15184 (N_15184,N_14739,N_14553);
xor U15185 (N_15185,N_14626,N_14771);
or U15186 (N_15186,N_14582,N_14406);
nor U15187 (N_15187,N_14746,N_14723);
xnor U15188 (N_15188,N_14401,N_14578);
xnor U15189 (N_15189,N_14682,N_14649);
xor U15190 (N_15190,N_14621,N_14564);
and U15191 (N_15191,N_14758,N_14570);
xor U15192 (N_15192,N_14717,N_14715);
nor U15193 (N_15193,N_14549,N_14610);
xnor U15194 (N_15194,N_14637,N_14569);
and U15195 (N_15195,N_14735,N_14667);
and U15196 (N_15196,N_14708,N_14619);
xor U15197 (N_15197,N_14734,N_14672);
nand U15198 (N_15198,N_14768,N_14493);
and U15199 (N_15199,N_14670,N_14727);
and U15200 (N_15200,N_15079,N_14853);
or U15201 (N_15201,N_14863,N_14934);
or U15202 (N_15202,N_14993,N_14809);
nor U15203 (N_15203,N_14962,N_14850);
and U15204 (N_15204,N_15185,N_15042);
or U15205 (N_15205,N_15061,N_15035);
nor U15206 (N_15206,N_14926,N_14901);
nor U15207 (N_15207,N_14970,N_15055);
and U15208 (N_15208,N_14900,N_14956);
xor U15209 (N_15209,N_14969,N_14996);
nor U15210 (N_15210,N_14922,N_15078);
xor U15211 (N_15211,N_14876,N_14932);
and U15212 (N_15212,N_15149,N_14843);
and U15213 (N_15213,N_15016,N_15024);
nand U15214 (N_15214,N_15182,N_14987);
or U15215 (N_15215,N_15073,N_15062);
or U15216 (N_15216,N_15069,N_15065);
or U15217 (N_15217,N_14842,N_15136);
nand U15218 (N_15218,N_15137,N_14965);
xor U15219 (N_15219,N_14930,N_14891);
nor U15220 (N_15220,N_15105,N_15031);
xnor U15221 (N_15221,N_15179,N_15199);
xnor U15222 (N_15222,N_14848,N_14890);
or U15223 (N_15223,N_15122,N_14874);
and U15224 (N_15224,N_15186,N_15006);
nor U15225 (N_15225,N_14919,N_15003);
and U15226 (N_15226,N_14920,N_14892);
xor U15227 (N_15227,N_15195,N_14946);
nor U15228 (N_15228,N_14935,N_15098);
xor U15229 (N_15229,N_15032,N_14894);
and U15230 (N_15230,N_14865,N_15094);
and U15231 (N_15231,N_15008,N_14802);
or U15232 (N_15232,N_14947,N_15027);
xor U15233 (N_15233,N_15036,N_15086);
or U15234 (N_15234,N_14806,N_14923);
or U15235 (N_15235,N_15070,N_15112);
nor U15236 (N_15236,N_14948,N_14999);
nand U15237 (N_15237,N_14974,N_15033);
xor U15238 (N_15238,N_15085,N_14955);
nand U15239 (N_15239,N_15047,N_15190);
nand U15240 (N_15240,N_14883,N_15020);
xnor U15241 (N_15241,N_14971,N_15180);
and U15242 (N_15242,N_15075,N_14852);
xnor U15243 (N_15243,N_15111,N_14849);
nor U15244 (N_15244,N_14844,N_14983);
nor U15245 (N_15245,N_15004,N_15191);
nand U15246 (N_15246,N_14985,N_15144);
nor U15247 (N_15247,N_15162,N_14879);
nor U15248 (N_15248,N_15177,N_15058);
nand U15249 (N_15249,N_14816,N_15128);
nor U15250 (N_15250,N_14885,N_14949);
or U15251 (N_15251,N_14944,N_15022);
or U15252 (N_15252,N_15138,N_14824);
and U15253 (N_15253,N_15151,N_14907);
and U15254 (N_15254,N_14941,N_15071);
nand U15255 (N_15255,N_14973,N_15146);
or U15256 (N_15256,N_15171,N_14942);
xor U15257 (N_15257,N_14927,N_15118);
nand U15258 (N_15258,N_15018,N_14821);
nand U15259 (N_15259,N_15198,N_14812);
and U15260 (N_15260,N_15045,N_15007);
xnor U15261 (N_15261,N_14937,N_15187);
nand U15262 (N_15262,N_14815,N_14840);
xor U15263 (N_15263,N_14978,N_14981);
xor U15264 (N_15264,N_14851,N_14810);
and U15265 (N_15265,N_14909,N_14915);
nand U15266 (N_15266,N_15117,N_14940);
and U15267 (N_15267,N_14833,N_14903);
xnor U15268 (N_15268,N_14868,N_15044);
xnor U15269 (N_15269,N_14838,N_15113);
xnor U15270 (N_15270,N_15120,N_14954);
xor U15271 (N_15271,N_14822,N_14814);
nor U15272 (N_15272,N_14959,N_14982);
and U15273 (N_15273,N_14857,N_14910);
nand U15274 (N_15274,N_14804,N_14882);
nand U15275 (N_15275,N_14813,N_15050);
or U15276 (N_15276,N_15013,N_15043);
nand U15277 (N_15277,N_15064,N_14984);
xnor U15278 (N_15278,N_14800,N_15099);
nor U15279 (N_15279,N_14823,N_14832);
and U15280 (N_15280,N_14951,N_15102);
or U15281 (N_15281,N_14958,N_14896);
nor U15282 (N_15282,N_15103,N_15145);
or U15283 (N_15283,N_15134,N_15131);
and U15284 (N_15284,N_15037,N_14887);
nor U15285 (N_15285,N_15126,N_15110);
nor U15286 (N_15286,N_14990,N_15125);
xnor U15287 (N_15287,N_15143,N_14827);
or U15288 (N_15288,N_15107,N_15160);
or U15289 (N_15289,N_15106,N_15097);
or U15290 (N_15290,N_15157,N_14889);
nand U15291 (N_15291,N_15021,N_14841);
or U15292 (N_15292,N_14898,N_14967);
and U15293 (N_15293,N_14914,N_15194);
nand U15294 (N_15294,N_14830,N_15000);
xnor U15295 (N_15295,N_15133,N_15141);
xnor U15296 (N_15296,N_15088,N_15012);
nand U15297 (N_15297,N_15038,N_14862);
and U15298 (N_15298,N_15135,N_15054);
or U15299 (N_15299,N_15080,N_15026);
xor U15300 (N_15300,N_14972,N_15166);
or U15301 (N_15301,N_15053,N_14859);
nor U15302 (N_15302,N_14867,N_15052);
xnor U15303 (N_15303,N_15041,N_15057);
nor U15304 (N_15304,N_14918,N_14871);
xor U15305 (N_15305,N_14906,N_14908);
nor U15306 (N_15306,N_14801,N_14864);
or U15307 (N_15307,N_14881,N_15139);
nand U15308 (N_15308,N_15193,N_14895);
nor U15309 (N_15309,N_15181,N_15176);
or U15310 (N_15310,N_15074,N_14888);
and U15311 (N_15311,N_15030,N_15002);
or U15312 (N_15312,N_14953,N_14899);
xnor U15313 (N_15313,N_15189,N_14945);
nor U15314 (N_15314,N_15156,N_15115);
xnor U15315 (N_15315,N_14831,N_14991);
xor U15316 (N_15316,N_15001,N_15108);
xnor U15317 (N_15317,N_14878,N_14839);
nor U15318 (N_15318,N_15028,N_14977);
nand U15319 (N_15319,N_15192,N_14807);
and U15320 (N_15320,N_15096,N_14911);
or U15321 (N_15321,N_14825,N_15029);
and U15322 (N_15322,N_15165,N_15060);
nor U15323 (N_15323,N_14998,N_15197);
xor U15324 (N_15324,N_15005,N_15017);
or U15325 (N_15325,N_15083,N_15158);
nor U15326 (N_15326,N_14836,N_15196);
and U15327 (N_15327,N_14936,N_14952);
or U15328 (N_15328,N_14826,N_14916);
nand U15329 (N_15329,N_15140,N_15084);
xnor U15330 (N_15330,N_14964,N_15059);
or U15331 (N_15331,N_14893,N_15172);
or U15332 (N_15332,N_15188,N_14884);
nand U15333 (N_15333,N_14873,N_15019);
nand U15334 (N_15334,N_14856,N_14811);
or U15335 (N_15335,N_14924,N_14870);
xor U15336 (N_15336,N_14980,N_14861);
nor U15337 (N_15337,N_15068,N_15147);
or U15338 (N_15338,N_14869,N_14933);
and U15339 (N_15339,N_14880,N_15169);
or U15340 (N_15340,N_14917,N_14819);
or U15341 (N_15341,N_14988,N_14854);
xor U15342 (N_15342,N_15170,N_14989);
and U15343 (N_15343,N_14928,N_15077);
nand U15344 (N_15344,N_14961,N_14829);
nand U15345 (N_15345,N_15116,N_14912);
nand U15346 (N_15346,N_14960,N_15164);
or U15347 (N_15347,N_14921,N_14803);
or U15348 (N_15348,N_14994,N_14931);
and U15349 (N_15349,N_14818,N_15150);
or U15350 (N_15350,N_15023,N_15034);
nand U15351 (N_15351,N_14995,N_15148);
and U15352 (N_15352,N_15104,N_15152);
and U15353 (N_15353,N_15114,N_15092);
nor U15354 (N_15354,N_15178,N_15100);
nand U15355 (N_15355,N_14897,N_15183);
xor U15356 (N_15356,N_15168,N_14957);
nor U15357 (N_15357,N_15048,N_14966);
nand U15358 (N_15358,N_15155,N_15067);
xnor U15359 (N_15359,N_15101,N_15076);
xnor U15360 (N_15360,N_15132,N_15130);
nor U15361 (N_15361,N_14820,N_15124);
nand U15362 (N_15362,N_15015,N_14968);
or U15363 (N_15363,N_14986,N_14808);
or U15364 (N_15364,N_15014,N_15127);
nand U15365 (N_15365,N_15142,N_15184);
nor U15366 (N_15366,N_14805,N_14963);
or U15367 (N_15367,N_15095,N_15081);
or U15368 (N_15368,N_14975,N_14858);
or U15369 (N_15369,N_14902,N_14845);
or U15370 (N_15370,N_14925,N_14834);
nor U15371 (N_15371,N_15040,N_15175);
xor U15372 (N_15372,N_15049,N_14929);
xnor U15373 (N_15373,N_15153,N_14950);
xnor U15374 (N_15374,N_15089,N_15087);
nand U15375 (N_15375,N_15163,N_15109);
nand U15376 (N_15376,N_14979,N_14939);
xor U15377 (N_15377,N_15090,N_15039);
xor U15378 (N_15378,N_15010,N_15173);
or U15379 (N_15379,N_15121,N_15161);
and U15380 (N_15380,N_15063,N_14846);
and U15381 (N_15381,N_15154,N_14943);
or U15382 (N_15382,N_15046,N_15072);
xor U15383 (N_15383,N_15167,N_15123);
nand U15384 (N_15384,N_15174,N_14872);
and U15385 (N_15385,N_15082,N_14877);
and U15386 (N_15386,N_14860,N_15011);
and U15387 (N_15387,N_14837,N_14997);
and U15388 (N_15388,N_14855,N_15056);
nor U15389 (N_15389,N_15025,N_15129);
nand U15390 (N_15390,N_14866,N_15009);
or U15391 (N_15391,N_15066,N_14847);
nor U15392 (N_15392,N_14976,N_15093);
nor U15393 (N_15393,N_15091,N_15119);
and U15394 (N_15394,N_14992,N_14913);
nor U15395 (N_15395,N_15051,N_14905);
nor U15396 (N_15396,N_14835,N_15159);
nor U15397 (N_15397,N_14886,N_14904);
or U15398 (N_15398,N_14875,N_14817);
or U15399 (N_15399,N_14938,N_14828);
or U15400 (N_15400,N_15188,N_15056);
and U15401 (N_15401,N_14998,N_14830);
nand U15402 (N_15402,N_15135,N_14838);
or U15403 (N_15403,N_14910,N_15006);
nand U15404 (N_15404,N_15182,N_15144);
and U15405 (N_15405,N_14858,N_15116);
or U15406 (N_15406,N_15090,N_14941);
or U15407 (N_15407,N_14910,N_14891);
nor U15408 (N_15408,N_14873,N_15051);
xnor U15409 (N_15409,N_15039,N_14917);
xnor U15410 (N_15410,N_14827,N_15043);
or U15411 (N_15411,N_14874,N_15063);
nand U15412 (N_15412,N_14846,N_14862);
nand U15413 (N_15413,N_15148,N_15059);
xnor U15414 (N_15414,N_15085,N_14844);
or U15415 (N_15415,N_14878,N_14931);
xnor U15416 (N_15416,N_15082,N_15125);
xnor U15417 (N_15417,N_15190,N_14879);
nand U15418 (N_15418,N_14871,N_14994);
nand U15419 (N_15419,N_14945,N_15159);
xor U15420 (N_15420,N_15039,N_14850);
and U15421 (N_15421,N_15116,N_15179);
xor U15422 (N_15422,N_14831,N_15091);
nand U15423 (N_15423,N_15149,N_15193);
nor U15424 (N_15424,N_14931,N_15183);
xor U15425 (N_15425,N_15148,N_15161);
nand U15426 (N_15426,N_14977,N_15085);
nor U15427 (N_15427,N_15146,N_15007);
nor U15428 (N_15428,N_14893,N_14995);
nor U15429 (N_15429,N_14842,N_15016);
or U15430 (N_15430,N_14824,N_14837);
nand U15431 (N_15431,N_15006,N_15029);
nor U15432 (N_15432,N_14880,N_14890);
nor U15433 (N_15433,N_14840,N_15190);
or U15434 (N_15434,N_15025,N_15021);
or U15435 (N_15435,N_15071,N_15131);
xor U15436 (N_15436,N_14854,N_15019);
xnor U15437 (N_15437,N_15082,N_15036);
xor U15438 (N_15438,N_14952,N_14803);
nor U15439 (N_15439,N_15012,N_15046);
or U15440 (N_15440,N_14883,N_15046);
or U15441 (N_15441,N_15107,N_14890);
xnor U15442 (N_15442,N_14990,N_14817);
xnor U15443 (N_15443,N_14928,N_15065);
or U15444 (N_15444,N_15075,N_14936);
and U15445 (N_15445,N_15186,N_15057);
xnor U15446 (N_15446,N_15145,N_14824);
or U15447 (N_15447,N_15020,N_14982);
and U15448 (N_15448,N_15118,N_14832);
or U15449 (N_15449,N_14905,N_14847);
xor U15450 (N_15450,N_14818,N_14898);
nand U15451 (N_15451,N_15129,N_14800);
xor U15452 (N_15452,N_14941,N_14906);
or U15453 (N_15453,N_15183,N_15063);
xor U15454 (N_15454,N_15015,N_15080);
nor U15455 (N_15455,N_15097,N_15099);
and U15456 (N_15456,N_14878,N_14829);
xnor U15457 (N_15457,N_14956,N_15172);
and U15458 (N_15458,N_15165,N_14951);
and U15459 (N_15459,N_15001,N_15112);
nand U15460 (N_15460,N_14872,N_15125);
nand U15461 (N_15461,N_14930,N_15103);
nor U15462 (N_15462,N_14967,N_14888);
nor U15463 (N_15463,N_14821,N_15060);
xnor U15464 (N_15464,N_14906,N_14867);
xnor U15465 (N_15465,N_15091,N_15017);
nor U15466 (N_15466,N_14866,N_15128);
and U15467 (N_15467,N_14955,N_14812);
nor U15468 (N_15468,N_15133,N_14867);
nor U15469 (N_15469,N_14824,N_15160);
nor U15470 (N_15470,N_15106,N_14973);
xor U15471 (N_15471,N_14992,N_14856);
nand U15472 (N_15472,N_15185,N_14857);
xnor U15473 (N_15473,N_15016,N_14895);
nand U15474 (N_15474,N_15115,N_15140);
and U15475 (N_15475,N_15059,N_14850);
nand U15476 (N_15476,N_15122,N_14845);
or U15477 (N_15477,N_14977,N_15194);
nand U15478 (N_15478,N_14997,N_14972);
or U15479 (N_15479,N_15023,N_15018);
xnor U15480 (N_15480,N_14925,N_14935);
or U15481 (N_15481,N_14833,N_14911);
xnor U15482 (N_15482,N_14848,N_15027);
and U15483 (N_15483,N_14936,N_14901);
and U15484 (N_15484,N_15068,N_15146);
nand U15485 (N_15485,N_14841,N_14880);
nand U15486 (N_15486,N_14949,N_15066);
or U15487 (N_15487,N_14996,N_15132);
nor U15488 (N_15488,N_15010,N_14870);
or U15489 (N_15489,N_14895,N_14922);
nor U15490 (N_15490,N_15118,N_14917);
xnor U15491 (N_15491,N_15036,N_14992);
xnor U15492 (N_15492,N_15126,N_14990);
nor U15493 (N_15493,N_14954,N_15081);
nor U15494 (N_15494,N_14849,N_14901);
nor U15495 (N_15495,N_15127,N_14819);
and U15496 (N_15496,N_15021,N_14825);
xor U15497 (N_15497,N_14899,N_14823);
xor U15498 (N_15498,N_14997,N_14978);
xnor U15499 (N_15499,N_15101,N_14844);
or U15500 (N_15500,N_14842,N_14863);
xor U15501 (N_15501,N_15027,N_15091);
nor U15502 (N_15502,N_14841,N_14973);
nor U15503 (N_15503,N_14880,N_14854);
nand U15504 (N_15504,N_14919,N_15164);
nor U15505 (N_15505,N_15090,N_14910);
nand U15506 (N_15506,N_15070,N_14820);
nand U15507 (N_15507,N_15076,N_14922);
nand U15508 (N_15508,N_15116,N_14901);
and U15509 (N_15509,N_15143,N_14837);
and U15510 (N_15510,N_14965,N_14844);
and U15511 (N_15511,N_15014,N_14987);
or U15512 (N_15512,N_14863,N_15002);
or U15513 (N_15513,N_14884,N_14976);
and U15514 (N_15514,N_14975,N_14894);
and U15515 (N_15515,N_15183,N_14810);
nor U15516 (N_15516,N_14860,N_14889);
nand U15517 (N_15517,N_14985,N_14815);
and U15518 (N_15518,N_14913,N_15182);
xnor U15519 (N_15519,N_14985,N_14974);
and U15520 (N_15520,N_14879,N_14918);
and U15521 (N_15521,N_15190,N_15134);
and U15522 (N_15522,N_15041,N_14992);
or U15523 (N_15523,N_14868,N_15113);
and U15524 (N_15524,N_14864,N_14820);
and U15525 (N_15525,N_15199,N_15177);
nand U15526 (N_15526,N_15155,N_15104);
nand U15527 (N_15527,N_14969,N_14934);
and U15528 (N_15528,N_14895,N_14956);
nand U15529 (N_15529,N_15160,N_14954);
xor U15530 (N_15530,N_15092,N_14966);
xnor U15531 (N_15531,N_14977,N_15114);
or U15532 (N_15532,N_15025,N_14843);
nand U15533 (N_15533,N_14872,N_15183);
nor U15534 (N_15534,N_14848,N_14821);
nor U15535 (N_15535,N_15067,N_15056);
xor U15536 (N_15536,N_15153,N_15190);
nor U15537 (N_15537,N_15023,N_14950);
nor U15538 (N_15538,N_14948,N_14804);
nand U15539 (N_15539,N_14962,N_14978);
and U15540 (N_15540,N_15054,N_14919);
or U15541 (N_15541,N_14905,N_15040);
nand U15542 (N_15542,N_15155,N_14815);
nor U15543 (N_15543,N_15063,N_15024);
or U15544 (N_15544,N_14809,N_14920);
nor U15545 (N_15545,N_15047,N_14915);
nor U15546 (N_15546,N_14834,N_14906);
xor U15547 (N_15547,N_15159,N_15075);
nand U15548 (N_15548,N_14907,N_14836);
nand U15549 (N_15549,N_14825,N_14981);
and U15550 (N_15550,N_15138,N_14853);
nand U15551 (N_15551,N_15024,N_15035);
xor U15552 (N_15552,N_14993,N_14939);
and U15553 (N_15553,N_14834,N_14950);
nor U15554 (N_15554,N_14931,N_15089);
nor U15555 (N_15555,N_14959,N_15190);
nor U15556 (N_15556,N_15053,N_15170);
nand U15557 (N_15557,N_14942,N_15134);
or U15558 (N_15558,N_14923,N_14926);
nor U15559 (N_15559,N_15109,N_14940);
nor U15560 (N_15560,N_15084,N_15175);
or U15561 (N_15561,N_14961,N_15116);
xor U15562 (N_15562,N_15161,N_14962);
nor U15563 (N_15563,N_14876,N_14977);
nor U15564 (N_15564,N_14800,N_15033);
xor U15565 (N_15565,N_15120,N_15196);
nor U15566 (N_15566,N_14849,N_15024);
nor U15567 (N_15567,N_14979,N_14867);
or U15568 (N_15568,N_15187,N_15154);
nand U15569 (N_15569,N_15137,N_14805);
nor U15570 (N_15570,N_14921,N_14812);
nand U15571 (N_15571,N_15199,N_15039);
or U15572 (N_15572,N_15169,N_15060);
and U15573 (N_15573,N_14904,N_15087);
xnor U15574 (N_15574,N_15147,N_15062);
xor U15575 (N_15575,N_14948,N_14900);
or U15576 (N_15576,N_14975,N_15198);
and U15577 (N_15577,N_14869,N_14997);
and U15578 (N_15578,N_14909,N_15044);
xnor U15579 (N_15579,N_15096,N_14962);
and U15580 (N_15580,N_15156,N_14866);
nor U15581 (N_15581,N_14906,N_15006);
nand U15582 (N_15582,N_15037,N_14937);
and U15583 (N_15583,N_14803,N_15151);
nor U15584 (N_15584,N_14913,N_14873);
and U15585 (N_15585,N_14999,N_15182);
or U15586 (N_15586,N_15171,N_14803);
nor U15587 (N_15587,N_15099,N_14810);
nor U15588 (N_15588,N_15020,N_14837);
or U15589 (N_15589,N_15180,N_14940);
nand U15590 (N_15590,N_14873,N_14947);
and U15591 (N_15591,N_14910,N_14907);
or U15592 (N_15592,N_14855,N_14854);
xnor U15593 (N_15593,N_15135,N_14830);
or U15594 (N_15594,N_15105,N_15034);
xnor U15595 (N_15595,N_14975,N_15185);
nor U15596 (N_15596,N_14887,N_14998);
or U15597 (N_15597,N_15061,N_14829);
nor U15598 (N_15598,N_15172,N_15040);
or U15599 (N_15599,N_15117,N_15031);
or U15600 (N_15600,N_15493,N_15304);
nor U15601 (N_15601,N_15378,N_15280);
nor U15602 (N_15602,N_15374,N_15536);
or U15603 (N_15603,N_15287,N_15202);
nand U15604 (N_15604,N_15276,N_15322);
nor U15605 (N_15605,N_15337,N_15343);
and U15606 (N_15606,N_15209,N_15362);
or U15607 (N_15607,N_15558,N_15239);
xnor U15608 (N_15608,N_15452,N_15565);
nor U15609 (N_15609,N_15501,N_15526);
xnor U15610 (N_15610,N_15246,N_15572);
xor U15611 (N_15611,N_15420,N_15363);
and U15612 (N_15612,N_15537,N_15282);
and U15613 (N_15613,N_15475,N_15563);
nor U15614 (N_15614,N_15308,N_15217);
and U15615 (N_15615,N_15271,N_15321);
and U15616 (N_15616,N_15522,N_15523);
and U15617 (N_15617,N_15547,N_15305);
or U15618 (N_15618,N_15402,N_15429);
xnor U15619 (N_15619,N_15510,N_15497);
nand U15620 (N_15620,N_15345,N_15208);
nand U15621 (N_15621,N_15361,N_15520);
nor U15622 (N_15622,N_15390,N_15592);
or U15623 (N_15623,N_15430,N_15240);
nand U15624 (N_15624,N_15210,N_15569);
and U15625 (N_15625,N_15479,N_15557);
and U15626 (N_15626,N_15231,N_15300);
xnor U15627 (N_15627,N_15439,N_15525);
or U15628 (N_15628,N_15260,N_15538);
or U15629 (N_15629,N_15410,N_15299);
or U15630 (N_15630,N_15443,N_15413);
xnor U15631 (N_15631,N_15532,N_15238);
and U15632 (N_15632,N_15294,N_15318);
xnor U15633 (N_15633,N_15415,N_15257);
nor U15634 (N_15634,N_15518,N_15561);
or U15635 (N_15635,N_15451,N_15460);
nor U15636 (N_15636,N_15233,N_15393);
xor U15637 (N_15637,N_15491,N_15350);
nor U15638 (N_15638,N_15423,N_15455);
or U15639 (N_15639,N_15488,N_15359);
and U15640 (N_15640,N_15505,N_15339);
nor U15641 (N_15641,N_15274,N_15449);
or U15642 (N_15642,N_15474,N_15458);
xnor U15643 (N_15643,N_15340,N_15407);
or U15644 (N_15644,N_15411,N_15293);
or U15645 (N_15645,N_15595,N_15216);
nand U15646 (N_15646,N_15213,N_15377);
nor U15647 (N_15647,N_15574,N_15462);
nand U15648 (N_15648,N_15498,N_15396);
and U15649 (N_15649,N_15492,N_15328);
or U15650 (N_15650,N_15485,N_15571);
nor U15651 (N_15651,N_15590,N_15327);
xnor U15652 (N_15652,N_15507,N_15244);
xor U15653 (N_15653,N_15292,N_15504);
xor U15654 (N_15654,N_15540,N_15567);
nand U15655 (N_15655,N_15234,N_15542);
xor U15656 (N_15656,N_15593,N_15579);
nand U15657 (N_15657,N_15319,N_15372);
and U15658 (N_15658,N_15387,N_15379);
nand U15659 (N_15659,N_15482,N_15478);
or U15660 (N_15660,N_15395,N_15367);
nand U15661 (N_15661,N_15370,N_15434);
nand U15662 (N_15662,N_15487,N_15466);
nand U15663 (N_15663,N_15323,N_15265);
nand U15664 (N_15664,N_15357,N_15316);
or U15665 (N_15665,N_15472,N_15219);
nor U15666 (N_15666,N_15235,N_15386);
and U15667 (N_15667,N_15530,N_15467);
nor U15668 (N_15668,N_15251,N_15576);
and U15669 (N_15669,N_15355,N_15405);
nand U15670 (N_15670,N_15222,N_15289);
nor U15671 (N_15671,N_15546,N_15366);
xor U15672 (N_15672,N_15469,N_15573);
nand U15673 (N_15673,N_15297,N_15221);
nor U15674 (N_15674,N_15228,N_15272);
xnor U15675 (N_15675,N_15404,N_15325);
xnor U15676 (N_15676,N_15264,N_15461);
or U15677 (N_15677,N_15566,N_15432);
nand U15678 (N_15678,N_15484,N_15514);
nor U15679 (N_15679,N_15227,N_15421);
or U15680 (N_15680,N_15438,N_15346);
or U15681 (N_15681,N_15380,N_15496);
or U15682 (N_15682,N_15495,N_15385);
nor U15683 (N_15683,N_15224,N_15425);
xor U15684 (N_15684,N_15597,N_15277);
nand U15685 (N_15685,N_15335,N_15200);
and U15686 (N_15686,N_15206,N_15435);
and U15687 (N_15687,N_15521,N_15334);
and U15688 (N_15688,N_15225,N_15422);
nor U15689 (N_15689,N_15317,N_15483);
xnor U15690 (N_15690,N_15281,N_15424);
xor U15691 (N_15691,N_15348,N_15591);
and U15692 (N_15692,N_15448,N_15551);
xnor U15693 (N_15693,N_15229,N_15416);
nor U15694 (N_15694,N_15347,N_15489);
or U15695 (N_15695,N_15583,N_15513);
nor U15696 (N_15696,N_15214,N_15440);
xnor U15697 (N_15697,N_15275,N_15531);
xnor U15698 (N_15698,N_15560,N_15311);
nor U15699 (N_15699,N_15494,N_15284);
xor U15700 (N_15700,N_15553,N_15550);
nor U15701 (N_15701,N_15204,N_15291);
xnor U15702 (N_15702,N_15476,N_15575);
nand U15703 (N_15703,N_15383,N_15309);
nand U15704 (N_15704,N_15242,N_15454);
or U15705 (N_15705,N_15330,N_15529);
and U15706 (N_15706,N_15249,N_15570);
nor U15707 (N_15707,N_15453,N_15252);
nor U15708 (N_15708,N_15268,N_15349);
nor U15709 (N_15709,N_15596,N_15427);
xor U15710 (N_15710,N_15490,N_15552);
or U15711 (N_15711,N_15486,N_15508);
and U15712 (N_15712,N_15578,N_15568);
nand U15713 (N_15713,N_15243,N_15392);
nand U15714 (N_15714,N_15223,N_15586);
xor U15715 (N_15715,N_15211,N_15302);
or U15716 (N_15716,N_15273,N_15545);
and U15717 (N_15717,N_15360,N_15266);
xnor U15718 (N_15718,N_15371,N_15356);
nor U15719 (N_15719,N_15290,N_15406);
or U15720 (N_15720,N_15418,N_15585);
nand U15721 (N_15721,N_15517,N_15519);
nor U15722 (N_15722,N_15205,N_15331);
nor U15723 (N_15723,N_15247,N_15320);
nand U15724 (N_15724,N_15237,N_15436);
and U15725 (N_15725,N_15263,N_15397);
and U15726 (N_15726,N_15506,N_15351);
xor U15727 (N_15727,N_15381,N_15500);
and U15728 (N_15728,N_15516,N_15559);
or U15729 (N_15729,N_15324,N_15384);
xnor U15730 (N_15730,N_15278,N_15203);
nand U15731 (N_15731,N_15388,N_15419);
nor U15732 (N_15732,N_15473,N_15408);
nor U15733 (N_15733,N_15218,N_15373);
nor U15734 (N_15734,N_15599,N_15255);
nand U15735 (N_15735,N_15256,N_15267);
xnor U15736 (N_15736,N_15564,N_15236);
and U15737 (N_15737,N_15344,N_15414);
nand U15738 (N_15738,N_15375,N_15212);
nand U15739 (N_15739,N_15463,N_15220);
nand U15740 (N_15740,N_15515,N_15254);
nand U15741 (N_15741,N_15301,N_15524);
or U15742 (N_15742,N_15261,N_15459);
xnor U15743 (N_15743,N_15534,N_15456);
nand U15744 (N_15744,N_15587,N_15365);
xor U15745 (N_15745,N_15303,N_15285);
xnor U15746 (N_15746,N_15446,N_15389);
or U15747 (N_15747,N_15230,N_15226);
and U15748 (N_15748,N_15241,N_15358);
xnor U15749 (N_15749,N_15465,N_15464);
nand U15750 (N_15750,N_15412,N_15588);
nor U15751 (N_15751,N_15433,N_15342);
nor U15752 (N_15752,N_15298,N_15582);
nor U15753 (N_15753,N_15376,N_15279);
and U15754 (N_15754,N_15270,N_15201);
nor U15755 (N_15755,N_15403,N_15437);
and U15756 (N_15756,N_15581,N_15354);
nor U15757 (N_15757,N_15580,N_15594);
nand U15758 (N_15758,N_15368,N_15539);
nor U15759 (N_15759,N_15250,N_15549);
xnor U15760 (N_15760,N_15283,N_15307);
and U15761 (N_15761,N_15296,N_15527);
nor U15762 (N_15762,N_15417,N_15450);
or U15763 (N_15763,N_15262,N_15533);
nand U15764 (N_15764,N_15584,N_15428);
or U15765 (N_15765,N_15258,N_15535);
nor U15766 (N_15766,N_15269,N_15468);
nand U15767 (N_15767,N_15431,N_15544);
nor U15768 (N_15768,N_15245,N_15295);
or U15769 (N_15769,N_15509,N_15471);
nor U15770 (N_15770,N_15502,N_15336);
nor U15771 (N_15771,N_15577,N_15333);
nor U15772 (N_15772,N_15444,N_15382);
or U15773 (N_15773,N_15477,N_15353);
and U15774 (N_15774,N_15480,N_15288);
nor U15775 (N_15775,N_15426,N_15554);
and U15776 (N_15776,N_15391,N_15409);
nor U15777 (N_15777,N_15400,N_15338);
and U15778 (N_15778,N_15589,N_15457);
xor U15779 (N_15779,N_15329,N_15207);
xnor U15780 (N_15780,N_15364,N_15286);
xor U15781 (N_15781,N_15442,N_15332);
nand U15782 (N_15782,N_15313,N_15511);
xnor U15783 (N_15783,N_15306,N_15555);
and U15784 (N_15784,N_15562,N_15352);
nand U15785 (N_15785,N_15556,N_15394);
xnor U15786 (N_15786,N_15598,N_15470);
nor U15787 (N_15787,N_15512,N_15541);
nor U15788 (N_15788,N_15232,N_15310);
and U15789 (N_15789,N_15499,N_15543);
or U15790 (N_15790,N_15369,N_15253);
xnor U15791 (N_15791,N_15315,N_15341);
nand U15792 (N_15792,N_15398,N_15447);
or U15793 (N_15793,N_15481,N_15259);
and U15794 (N_15794,N_15326,N_15312);
or U15795 (N_15795,N_15528,N_15445);
and U15796 (N_15796,N_15548,N_15503);
nand U15797 (N_15797,N_15248,N_15401);
nor U15798 (N_15798,N_15441,N_15314);
and U15799 (N_15799,N_15215,N_15399);
nor U15800 (N_15800,N_15466,N_15343);
nor U15801 (N_15801,N_15486,N_15549);
nor U15802 (N_15802,N_15510,N_15247);
nor U15803 (N_15803,N_15236,N_15455);
nor U15804 (N_15804,N_15211,N_15524);
xor U15805 (N_15805,N_15482,N_15205);
and U15806 (N_15806,N_15307,N_15242);
nor U15807 (N_15807,N_15253,N_15343);
nor U15808 (N_15808,N_15293,N_15309);
nand U15809 (N_15809,N_15512,N_15211);
and U15810 (N_15810,N_15555,N_15308);
xor U15811 (N_15811,N_15564,N_15444);
and U15812 (N_15812,N_15483,N_15408);
nand U15813 (N_15813,N_15355,N_15279);
and U15814 (N_15814,N_15368,N_15589);
nor U15815 (N_15815,N_15319,N_15485);
or U15816 (N_15816,N_15259,N_15292);
xnor U15817 (N_15817,N_15278,N_15491);
nor U15818 (N_15818,N_15482,N_15399);
and U15819 (N_15819,N_15493,N_15298);
or U15820 (N_15820,N_15238,N_15384);
nor U15821 (N_15821,N_15535,N_15454);
xnor U15822 (N_15822,N_15508,N_15364);
or U15823 (N_15823,N_15306,N_15312);
nand U15824 (N_15824,N_15271,N_15439);
nor U15825 (N_15825,N_15391,N_15535);
nor U15826 (N_15826,N_15597,N_15558);
or U15827 (N_15827,N_15253,N_15510);
and U15828 (N_15828,N_15384,N_15549);
or U15829 (N_15829,N_15546,N_15236);
xor U15830 (N_15830,N_15238,N_15369);
xnor U15831 (N_15831,N_15506,N_15249);
or U15832 (N_15832,N_15314,N_15586);
nor U15833 (N_15833,N_15435,N_15509);
nand U15834 (N_15834,N_15477,N_15484);
nor U15835 (N_15835,N_15546,N_15299);
nor U15836 (N_15836,N_15567,N_15283);
nor U15837 (N_15837,N_15389,N_15452);
nor U15838 (N_15838,N_15215,N_15525);
nor U15839 (N_15839,N_15233,N_15368);
and U15840 (N_15840,N_15504,N_15234);
nor U15841 (N_15841,N_15591,N_15403);
xnor U15842 (N_15842,N_15322,N_15218);
nand U15843 (N_15843,N_15500,N_15549);
xnor U15844 (N_15844,N_15451,N_15259);
xnor U15845 (N_15845,N_15460,N_15238);
nor U15846 (N_15846,N_15400,N_15462);
xnor U15847 (N_15847,N_15234,N_15259);
or U15848 (N_15848,N_15596,N_15229);
xnor U15849 (N_15849,N_15380,N_15291);
or U15850 (N_15850,N_15486,N_15533);
nand U15851 (N_15851,N_15294,N_15588);
nor U15852 (N_15852,N_15488,N_15459);
or U15853 (N_15853,N_15520,N_15433);
nand U15854 (N_15854,N_15538,N_15206);
nand U15855 (N_15855,N_15253,N_15222);
xor U15856 (N_15856,N_15358,N_15417);
and U15857 (N_15857,N_15432,N_15357);
and U15858 (N_15858,N_15432,N_15322);
xnor U15859 (N_15859,N_15549,N_15413);
or U15860 (N_15860,N_15533,N_15394);
xnor U15861 (N_15861,N_15308,N_15279);
nand U15862 (N_15862,N_15541,N_15367);
and U15863 (N_15863,N_15432,N_15427);
nor U15864 (N_15864,N_15568,N_15486);
xnor U15865 (N_15865,N_15337,N_15355);
xnor U15866 (N_15866,N_15240,N_15589);
nor U15867 (N_15867,N_15233,N_15509);
xor U15868 (N_15868,N_15336,N_15312);
xnor U15869 (N_15869,N_15460,N_15383);
and U15870 (N_15870,N_15311,N_15316);
nand U15871 (N_15871,N_15578,N_15307);
xnor U15872 (N_15872,N_15533,N_15296);
nor U15873 (N_15873,N_15514,N_15333);
nor U15874 (N_15874,N_15596,N_15230);
nand U15875 (N_15875,N_15321,N_15436);
and U15876 (N_15876,N_15463,N_15570);
or U15877 (N_15877,N_15540,N_15499);
and U15878 (N_15878,N_15469,N_15406);
and U15879 (N_15879,N_15214,N_15227);
or U15880 (N_15880,N_15323,N_15591);
and U15881 (N_15881,N_15210,N_15252);
nand U15882 (N_15882,N_15504,N_15517);
nor U15883 (N_15883,N_15577,N_15388);
or U15884 (N_15884,N_15456,N_15312);
xnor U15885 (N_15885,N_15232,N_15252);
and U15886 (N_15886,N_15396,N_15387);
nor U15887 (N_15887,N_15268,N_15383);
and U15888 (N_15888,N_15375,N_15221);
or U15889 (N_15889,N_15373,N_15284);
nand U15890 (N_15890,N_15217,N_15405);
and U15891 (N_15891,N_15495,N_15346);
nand U15892 (N_15892,N_15457,N_15428);
nand U15893 (N_15893,N_15509,N_15324);
nor U15894 (N_15894,N_15203,N_15466);
and U15895 (N_15895,N_15292,N_15430);
nand U15896 (N_15896,N_15389,N_15297);
or U15897 (N_15897,N_15549,N_15310);
or U15898 (N_15898,N_15240,N_15335);
nor U15899 (N_15899,N_15332,N_15395);
and U15900 (N_15900,N_15355,N_15588);
nand U15901 (N_15901,N_15563,N_15562);
nor U15902 (N_15902,N_15337,N_15478);
and U15903 (N_15903,N_15225,N_15357);
nand U15904 (N_15904,N_15412,N_15477);
xnor U15905 (N_15905,N_15225,N_15252);
and U15906 (N_15906,N_15555,N_15340);
nor U15907 (N_15907,N_15554,N_15254);
or U15908 (N_15908,N_15529,N_15561);
and U15909 (N_15909,N_15447,N_15588);
nor U15910 (N_15910,N_15322,N_15309);
and U15911 (N_15911,N_15232,N_15417);
nor U15912 (N_15912,N_15252,N_15238);
and U15913 (N_15913,N_15447,N_15325);
nand U15914 (N_15914,N_15374,N_15499);
and U15915 (N_15915,N_15217,N_15293);
and U15916 (N_15916,N_15465,N_15586);
nand U15917 (N_15917,N_15355,N_15502);
nand U15918 (N_15918,N_15349,N_15248);
and U15919 (N_15919,N_15304,N_15262);
xnor U15920 (N_15920,N_15417,N_15483);
or U15921 (N_15921,N_15351,N_15584);
xnor U15922 (N_15922,N_15353,N_15230);
or U15923 (N_15923,N_15352,N_15319);
or U15924 (N_15924,N_15457,N_15342);
xnor U15925 (N_15925,N_15429,N_15338);
and U15926 (N_15926,N_15255,N_15262);
nand U15927 (N_15927,N_15596,N_15424);
xnor U15928 (N_15928,N_15372,N_15526);
nor U15929 (N_15929,N_15431,N_15458);
nand U15930 (N_15930,N_15465,N_15492);
xnor U15931 (N_15931,N_15485,N_15254);
and U15932 (N_15932,N_15427,N_15236);
xnor U15933 (N_15933,N_15349,N_15208);
xor U15934 (N_15934,N_15523,N_15387);
or U15935 (N_15935,N_15539,N_15397);
xnor U15936 (N_15936,N_15447,N_15424);
nand U15937 (N_15937,N_15398,N_15298);
nand U15938 (N_15938,N_15217,N_15401);
nor U15939 (N_15939,N_15520,N_15239);
xor U15940 (N_15940,N_15397,N_15595);
and U15941 (N_15941,N_15221,N_15311);
xor U15942 (N_15942,N_15574,N_15406);
and U15943 (N_15943,N_15388,N_15548);
and U15944 (N_15944,N_15561,N_15267);
xnor U15945 (N_15945,N_15287,N_15219);
or U15946 (N_15946,N_15370,N_15365);
and U15947 (N_15947,N_15415,N_15434);
or U15948 (N_15948,N_15266,N_15364);
xor U15949 (N_15949,N_15439,N_15299);
and U15950 (N_15950,N_15441,N_15439);
xor U15951 (N_15951,N_15515,N_15566);
nor U15952 (N_15952,N_15585,N_15338);
xor U15953 (N_15953,N_15405,N_15302);
xnor U15954 (N_15954,N_15580,N_15219);
and U15955 (N_15955,N_15340,N_15439);
nand U15956 (N_15956,N_15421,N_15509);
nand U15957 (N_15957,N_15493,N_15581);
xnor U15958 (N_15958,N_15309,N_15295);
and U15959 (N_15959,N_15575,N_15408);
xnor U15960 (N_15960,N_15578,N_15324);
and U15961 (N_15961,N_15446,N_15233);
or U15962 (N_15962,N_15469,N_15431);
nor U15963 (N_15963,N_15572,N_15535);
nand U15964 (N_15964,N_15516,N_15310);
nand U15965 (N_15965,N_15438,N_15393);
xor U15966 (N_15966,N_15259,N_15503);
or U15967 (N_15967,N_15518,N_15558);
nor U15968 (N_15968,N_15262,N_15210);
nand U15969 (N_15969,N_15312,N_15441);
xnor U15970 (N_15970,N_15214,N_15572);
nand U15971 (N_15971,N_15530,N_15367);
nor U15972 (N_15972,N_15411,N_15275);
xnor U15973 (N_15973,N_15207,N_15317);
nand U15974 (N_15974,N_15221,N_15419);
and U15975 (N_15975,N_15234,N_15242);
xnor U15976 (N_15976,N_15385,N_15318);
nand U15977 (N_15977,N_15213,N_15286);
nand U15978 (N_15978,N_15200,N_15415);
nand U15979 (N_15979,N_15407,N_15274);
or U15980 (N_15980,N_15254,N_15427);
nor U15981 (N_15981,N_15598,N_15270);
and U15982 (N_15982,N_15535,N_15366);
nor U15983 (N_15983,N_15262,N_15385);
nand U15984 (N_15984,N_15491,N_15560);
or U15985 (N_15985,N_15568,N_15521);
and U15986 (N_15986,N_15440,N_15207);
nor U15987 (N_15987,N_15294,N_15495);
or U15988 (N_15988,N_15397,N_15316);
and U15989 (N_15989,N_15304,N_15249);
nand U15990 (N_15990,N_15441,N_15326);
xnor U15991 (N_15991,N_15376,N_15594);
nor U15992 (N_15992,N_15435,N_15458);
nor U15993 (N_15993,N_15548,N_15268);
nand U15994 (N_15994,N_15224,N_15362);
nand U15995 (N_15995,N_15537,N_15203);
nor U15996 (N_15996,N_15504,N_15246);
nand U15997 (N_15997,N_15389,N_15242);
xor U15998 (N_15998,N_15478,N_15531);
xor U15999 (N_15999,N_15281,N_15336);
and U16000 (N_16000,N_15947,N_15838);
nand U16001 (N_16001,N_15997,N_15792);
nor U16002 (N_16002,N_15676,N_15952);
or U16003 (N_16003,N_15945,N_15764);
and U16004 (N_16004,N_15881,N_15647);
and U16005 (N_16005,N_15907,N_15756);
and U16006 (N_16006,N_15710,N_15773);
or U16007 (N_16007,N_15995,N_15903);
xor U16008 (N_16008,N_15631,N_15716);
and U16009 (N_16009,N_15790,N_15815);
and U16010 (N_16010,N_15731,N_15877);
or U16011 (N_16011,N_15612,N_15748);
xor U16012 (N_16012,N_15973,N_15974);
and U16013 (N_16013,N_15924,N_15704);
xnor U16014 (N_16014,N_15772,N_15854);
or U16015 (N_16015,N_15806,N_15776);
xnor U16016 (N_16016,N_15630,N_15617);
or U16017 (N_16017,N_15698,N_15934);
or U16018 (N_16018,N_15921,N_15694);
nand U16019 (N_16019,N_15981,N_15692);
or U16020 (N_16020,N_15942,N_15960);
or U16021 (N_16021,N_15844,N_15887);
or U16022 (N_16022,N_15732,N_15988);
nand U16023 (N_16023,N_15965,N_15917);
nand U16024 (N_16024,N_15697,N_15798);
nand U16025 (N_16025,N_15848,N_15778);
nor U16026 (N_16026,N_15791,N_15898);
nand U16027 (N_16027,N_15992,N_15849);
xor U16028 (N_16028,N_15669,N_15739);
or U16029 (N_16029,N_15846,N_15714);
nor U16030 (N_16030,N_15969,N_15991);
and U16031 (N_16031,N_15803,N_15950);
or U16032 (N_16032,N_15636,N_15883);
or U16033 (N_16033,N_15938,N_15637);
and U16034 (N_16034,N_15724,N_15823);
nand U16035 (N_16035,N_15619,N_15789);
nand U16036 (N_16036,N_15999,N_15605);
and U16037 (N_16037,N_15654,N_15985);
or U16038 (N_16038,N_15680,N_15616);
and U16039 (N_16039,N_15750,N_15648);
nor U16040 (N_16040,N_15868,N_15735);
xnor U16041 (N_16041,N_15864,N_15674);
nand U16042 (N_16042,N_15953,N_15665);
xor U16043 (N_16043,N_15876,N_15920);
and U16044 (N_16044,N_15830,N_15662);
or U16045 (N_16045,N_15640,N_15705);
nor U16046 (N_16046,N_15908,N_15769);
or U16047 (N_16047,N_15979,N_15645);
or U16048 (N_16048,N_15891,N_15747);
nand U16049 (N_16049,N_15786,N_15930);
nor U16050 (N_16050,N_15976,N_15726);
or U16051 (N_16051,N_15784,N_15866);
nand U16052 (N_16052,N_15805,N_15851);
xnor U16053 (N_16053,N_15712,N_15836);
and U16054 (N_16054,N_15743,N_15807);
nand U16055 (N_16055,N_15730,N_15780);
and U16056 (N_16056,N_15656,N_15810);
or U16057 (N_16057,N_15996,N_15925);
or U16058 (N_16058,N_15941,N_15812);
or U16059 (N_16059,N_15837,N_15801);
or U16060 (N_16060,N_15886,N_15847);
nand U16061 (N_16061,N_15659,N_15781);
nand U16062 (N_16062,N_15977,N_15707);
or U16063 (N_16063,N_15723,N_15777);
or U16064 (N_16064,N_15989,N_15690);
or U16065 (N_16065,N_15679,N_15763);
and U16066 (N_16066,N_15774,N_15623);
xnor U16067 (N_16067,N_15821,N_15949);
and U16068 (N_16068,N_15978,N_15632);
and U16069 (N_16069,N_15845,N_15758);
or U16070 (N_16070,N_15668,N_15695);
nor U16071 (N_16071,N_15913,N_15613);
and U16072 (N_16072,N_15653,N_15975);
nand U16073 (N_16073,N_15892,N_15775);
xnor U16074 (N_16074,N_15703,N_15923);
and U16075 (N_16075,N_15682,N_15956);
xor U16076 (N_16076,N_15737,N_15753);
xor U16077 (N_16077,N_15993,N_15618);
and U16078 (N_16078,N_15893,N_15918);
nor U16079 (N_16079,N_15661,N_15833);
nor U16080 (N_16080,N_15650,N_15929);
xnor U16081 (N_16081,N_15606,N_15888);
nand U16082 (N_16082,N_15853,N_15633);
xnor U16083 (N_16083,N_15880,N_15926);
nor U16084 (N_16084,N_15608,N_15788);
xnor U16085 (N_16085,N_15994,N_15813);
nor U16086 (N_16086,N_15700,N_15809);
or U16087 (N_16087,N_15715,N_15691);
nand U16088 (N_16088,N_15787,N_15986);
nor U16089 (N_16089,N_15900,N_15884);
xnor U16090 (N_16090,N_15827,N_15754);
and U16091 (N_16091,N_15879,N_15804);
xnor U16092 (N_16092,N_15889,N_15733);
xor U16093 (N_16093,N_15600,N_15839);
xor U16094 (N_16094,N_15914,N_15931);
xor U16095 (N_16095,N_15624,N_15980);
xnor U16096 (N_16096,N_15762,N_15987);
and U16097 (N_16097,N_15760,N_15629);
or U16098 (N_16098,N_15818,N_15873);
xnor U16099 (N_16099,N_15751,N_15664);
and U16100 (N_16100,N_15615,N_15948);
xor U16101 (N_16101,N_15741,N_15660);
or U16102 (N_16102,N_15872,N_15785);
nor U16103 (N_16103,N_15939,N_15765);
nor U16104 (N_16104,N_15603,N_15708);
or U16105 (N_16105,N_15675,N_15718);
nand U16106 (N_16106,N_15983,N_15646);
or U16107 (N_16107,N_15711,N_15706);
nor U16108 (N_16108,N_15610,N_15857);
or U16109 (N_16109,N_15912,N_15782);
or U16110 (N_16110,N_15614,N_15819);
nor U16111 (N_16111,N_15644,N_15828);
nor U16112 (N_16112,N_15916,N_15936);
nand U16113 (N_16113,N_15673,N_15869);
nor U16114 (N_16114,N_15964,N_15767);
nand U16115 (N_16115,N_15797,N_15970);
nor U16116 (N_16116,N_15933,N_15688);
nand U16117 (N_16117,N_15841,N_15746);
xnor U16118 (N_16118,N_15658,N_15728);
or U16119 (N_16119,N_15943,N_15744);
and U16120 (N_16120,N_15915,N_15859);
nand U16121 (N_16121,N_15909,N_15865);
nor U16122 (N_16122,N_15685,N_15814);
and U16123 (N_16123,N_15713,N_15681);
nand U16124 (N_16124,N_15684,N_15878);
xor U16125 (N_16125,N_15897,N_15642);
xnor U16126 (N_16126,N_15800,N_15861);
xor U16127 (N_16127,N_15829,N_15719);
nor U16128 (N_16128,N_15874,N_15628);
nand U16129 (N_16129,N_15899,N_15609);
xor U16130 (N_16130,N_15602,N_15852);
xnor U16131 (N_16131,N_15755,N_15966);
or U16132 (N_16132,N_15902,N_15770);
or U16133 (N_16133,N_15689,N_15842);
xor U16134 (N_16134,N_15655,N_15875);
xnor U16135 (N_16135,N_15699,N_15937);
and U16136 (N_16136,N_15639,N_15687);
and U16137 (N_16137,N_15727,N_15783);
nand U16138 (N_16138,N_15935,N_15822);
nand U16139 (N_16139,N_15843,N_15972);
or U16140 (N_16140,N_15802,N_15749);
nor U16141 (N_16141,N_15638,N_15820);
or U16142 (N_16142,N_15811,N_15955);
nand U16143 (N_16143,N_15627,N_15862);
nor U16144 (N_16144,N_15634,N_15611);
xor U16145 (N_16145,N_15982,N_15670);
nand U16146 (N_16146,N_15890,N_15796);
xor U16147 (N_16147,N_15834,N_15896);
nor U16148 (N_16148,N_15667,N_15626);
and U16149 (N_16149,N_15677,N_15971);
nor U16150 (N_16150,N_15816,N_15725);
xnor U16151 (N_16151,N_15946,N_15871);
nor U16152 (N_16152,N_15652,N_15824);
nor U16153 (N_16153,N_15779,N_15919);
and U16154 (N_16154,N_15702,N_15906);
nor U16155 (N_16155,N_15958,N_15604);
or U16156 (N_16156,N_15709,N_15601);
xor U16157 (N_16157,N_15922,N_15752);
or U16158 (N_16158,N_15683,N_15808);
or U16159 (N_16159,N_15635,N_15940);
nand U16160 (N_16160,N_15759,N_15738);
and U16161 (N_16161,N_15729,N_15771);
or U16162 (N_16162,N_15740,N_15793);
and U16163 (N_16163,N_15734,N_15693);
xnor U16164 (N_16164,N_15858,N_15825);
xor U16165 (N_16165,N_15951,N_15643);
nor U16166 (N_16166,N_15686,N_15666);
nand U16167 (N_16167,N_15968,N_15717);
nand U16168 (N_16168,N_15696,N_15722);
nand U16169 (N_16169,N_15867,N_15651);
or U16170 (N_16170,N_15959,N_15885);
nand U16171 (N_16171,N_15721,N_15850);
or U16172 (N_16172,N_15990,N_15928);
or U16173 (N_16173,N_15720,N_15742);
nand U16174 (N_16174,N_15641,N_15962);
nand U16175 (N_16175,N_15954,N_15963);
or U16176 (N_16176,N_15984,N_15998);
nor U16177 (N_16177,N_15766,N_15607);
nand U16178 (N_16178,N_15625,N_15961);
xor U16179 (N_16179,N_15910,N_15894);
nand U16180 (N_16180,N_15761,N_15768);
and U16181 (N_16181,N_15826,N_15856);
xor U16182 (N_16182,N_15831,N_15932);
xnor U16183 (N_16183,N_15882,N_15663);
nand U16184 (N_16184,N_15832,N_15895);
nand U16185 (N_16185,N_15620,N_15794);
and U16186 (N_16186,N_15799,N_15745);
nor U16187 (N_16187,N_15657,N_15860);
or U16188 (N_16188,N_15621,N_15957);
nor U16189 (N_16189,N_15870,N_15905);
and U16190 (N_16190,N_15757,N_15863);
xor U16191 (N_16191,N_15817,N_15927);
and U16192 (N_16192,N_15840,N_15736);
nand U16193 (N_16193,N_15622,N_15901);
or U16194 (N_16194,N_15904,N_15795);
or U16195 (N_16195,N_15649,N_15855);
or U16196 (N_16196,N_15672,N_15701);
xor U16197 (N_16197,N_15678,N_15944);
nor U16198 (N_16198,N_15911,N_15671);
nor U16199 (N_16199,N_15835,N_15967);
or U16200 (N_16200,N_15938,N_15970);
or U16201 (N_16201,N_15831,N_15981);
or U16202 (N_16202,N_15637,N_15815);
nand U16203 (N_16203,N_15681,N_15702);
or U16204 (N_16204,N_15724,N_15921);
or U16205 (N_16205,N_15619,N_15959);
nor U16206 (N_16206,N_15649,N_15646);
and U16207 (N_16207,N_15697,N_15761);
or U16208 (N_16208,N_15690,N_15683);
and U16209 (N_16209,N_15605,N_15601);
nor U16210 (N_16210,N_15736,N_15654);
xnor U16211 (N_16211,N_15705,N_15749);
nand U16212 (N_16212,N_15925,N_15701);
xnor U16213 (N_16213,N_15708,N_15634);
and U16214 (N_16214,N_15679,N_15889);
nor U16215 (N_16215,N_15763,N_15962);
or U16216 (N_16216,N_15967,N_15777);
or U16217 (N_16217,N_15609,N_15706);
and U16218 (N_16218,N_15601,N_15898);
xor U16219 (N_16219,N_15804,N_15813);
and U16220 (N_16220,N_15693,N_15847);
nand U16221 (N_16221,N_15827,N_15942);
nor U16222 (N_16222,N_15813,N_15634);
and U16223 (N_16223,N_15830,N_15809);
nand U16224 (N_16224,N_15843,N_15740);
and U16225 (N_16225,N_15673,N_15659);
nand U16226 (N_16226,N_15980,N_15970);
xnor U16227 (N_16227,N_15883,N_15813);
nor U16228 (N_16228,N_15621,N_15913);
nand U16229 (N_16229,N_15680,N_15689);
or U16230 (N_16230,N_15857,N_15780);
nor U16231 (N_16231,N_15640,N_15684);
nor U16232 (N_16232,N_15805,N_15600);
or U16233 (N_16233,N_15719,N_15928);
or U16234 (N_16234,N_15993,N_15915);
nor U16235 (N_16235,N_15923,N_15608);
nand U16236 (N_16236,N_15816,N_15760);
xor U16237 (N_16237,N_15855,N_15950);
nand U16238 (N_16238,N_15953,N_15765);
nand U16239 (N_16239,N_15926,N_15843);
or U16240 (N_16240,N_15650,N_15977);
and U16241 (N_16241,N_15797,N_15677);
xor U16242 (N_16242,N_15833,N_15827);
nand U16243 (N_16243,N_15708,N_15810);
nand U16244 (N_16244,N_15794,N_15612);
xnor U16245 (N_16245,N_15689,N_15942);
and U16246 (N_16246,N_15859,N_15934);
nor U16247 (N_16247,N_15964,N_15924);
and U16248 (N_16248,N_15839,N_15669);
nand U16249 (N_16249,N_15660,N_15752);
or U16250 (N_16250,N_15659,N_15827);
nand U16251 (N_16251,N_15883,N_15845);
nand U16252 (N_16252,N_15750,N_15748);
nand U16253 (N_16253,N_15982,N_15876);
or U16254 (N_16254,N_15981,N_15899);
nand U16255 (N_16255,N_15621,N_15756);
nor U16256 (N_16256,N_15759,N_15920);
nand U16257 (N_16257,N_15749,N_15960);
nand U16258 (N_16258,N_15963,N_15695);
nor U16259 (N_16259,N_15841,N_15813);
nand U16260 (N_16260,N_15944,N_15739);
and U16261 (N_16261,N_15886,N_15942);
and U16262 (N_16262,N_15656,N_15730);
xnor U16263 (N_16263,N_15780,N_15639);
or U16264 (N_16264,N_15897,N_15656);
nor U16265 (N_16265,N_15940,N_15726);
and U16266 (N_16266,N_15842,N_15901);
or U16267 (N_16267,N_15841,N_15764);
or U16268 (N_16268,N_15784,N_15620);
xnor U16269 (N_16269,N_15644,N_15876);
and U16270 (N_16270,N_15682,N_15701);
nand U16271 (N_16271,N_15918,N_15663);
nor U16272 (N_16272,N_15867,N_15659);
or U16273 (N_16273,N_15696,N_15944);
or U16274 (N_16274,N_15935,N_15996);
and U16275 (N_16275,N_15809,N_15608);
or U16276 (N_16276,N_15841,N_15710);
nand U16277 (N_16277,N_15813,N_15801);
or U16278 (N_16278,N_15937,N_15637);
xnor U16279 (N_16279,N_15849,N_15999);
nor U16280 (N_16280,N_15721,N_15651);
and U16281 (N_16281,N_15937,N_15963);
and U16282 (N_16282,N_15639,N_15779);
xor U16283 (N_16283,N_15865,N_15699);
nand U16284 (N_16284,N_15966,N_15975);
and U16285 (N_16285,N_15735,N_15833);
or U16286 (N_16286,N_15600,N_15855);
xnor U16287 (N_16287,N_15987,N_15884);
xor U16288 (N_16288,N_15671,N_15692);
and U16289 (N_16289,N_15996,N_15922);
and U16290 (N_16290,N_15880,N_15762);
nor U16291 (N_16291,N_15739,N_15625);
xnor U16292 (N_16292,N_15827,N_15625);
and U16293 (N_16293,N_15817,N_15828);
nor U16294 (N_16294,N_15973,N_15942);
and U16295 (N_16295,N_15754,N_15851);
nand U16296 (N_16296,N_15727,N_15674);
xnor U16297 (N_16297,N_15869,N_15734);
or U16298 (N_16298,N_15717,N_15858);
nand U16299 (N_16299,N_15686,N_15669);
xor U16300 (N_16300,N_15822,N_15651);
and U16301 (N_16301,N_15865,N_15771);
nor U16302 (N_16302,N_15688,N_15995);
xor U16303 (N_16303,N_15810,N_15722);
xor U16304 (N_16304,N_15886,N_15839);
or U16305 (N_16305,N_15780,N_15901);
nand U16306 (N_16306,N_15832,N_15931);
xor U16307 (N_16307,N_15884,N_15907);
nand U16308 (N_16308,N_15921,N_15805);
nand U16309 (N_16309,N_15811,N_15791);
or U16310 (N_16310,N_15789,N_15930);
or U16311 (N_16311,N_15901,N_15854);
nor U16312 (N_16312,N_15882,N_15948);
and U16313 (N_16313,N_15895,N_15771);
nand U16314 (N_16314,N_15871,N_15776);
nand U16315 (N_16315,N_15929,N_15739);
or U16316 (N_16316,N_15770,N_15631);
nand U16317 (N_16317,N_15946,N_15668);
xor U16318 (N_16318,N_15911,N_15926);
nor U16319 (N_16319,N_15790,N_15983);
nor U16320 (N_16320,N_15793,N_15722);
nor U16321 (N_16321,N_15762,N_15738);
nor U16322 (N_16322,N_15877,N_15990);
or U16323 (N_16323,N_15878,N_15628);
nor U16324 (N_16324,N_15788,N_15665);
xnor U16325 (N_16325,N_15921,N_15750);
nand U16326 (N_16326,N_15669,N_15959);
or U16327 (N_16327,N_15874,N_15745);
nor U16328 (N_16328,N_15643,N_15981);
nor U16329 (N_16329,N_15891,N_15644);
and U16330 (N_16330,N_15812,N_15640);
or U16331 (N_16331,N_15711,N_15984);
and U16332 (N_16332,N_15771,N_15693);
xor U16333 (N_16333,N_15664,N_15978);
nand U16334 (N_16334,N_15706,N_15972);
nor U16335 (N_16335,N_15603,N_15883);
nand U16336 (N_16336,N_15772,N_15630);
or U16337 (N_16337,N_15716,N_15824);
nor U16338 (N_16338,N_15834,N_15827);
or U16339 (N_16339,N_15880,N_15999);
and U16340 (N_16340,N_15617,N_15710);
nor U16341 (N_16341,N_15959,N_15860);
nor U16342 (N_16342,N_15949,N_15869);
or U16343 (N_16343,N_15846,N_15729);
and U16344 (N_16344,N_15942,N_15816);
nand U16345 (N_16345,N_15740,N_15687);
and U16346 (N_16346,N_15924,N_15756);
nor U16347 (N_16347,N_15648,N_15726);
and U16348 (N_16348,N_15770,N_15648);
nor U16349 (N_16349,N_15607,N_15700);
nand U16350 (N_16350,N_15847,N_15936);
xor U16351 (N_16351,N_15730,N_15915);
nor U16352 (N_16352,N_15966,N_15899);
nor U16353 (N_16353,N_15874,N_15893);
xnor U16354 (N_16354,N_15808,N_15758);
nand U16355 (N_16355,N_15847,N_15751);
and U16356 (N_16356,N_15885,N_15881);
or U16357 (N_16357,N_15774,N_15798);
xnor U16358 (N_16358,N_15602,N_15902);
or U16359 (N_16359,N_15836,N_15799);
or U16360 (N_16360,N_15768,N_15884);
xnor U16361 (N_16361,N_15985,N_15931);
nor U16362 (N_16362,N_15770,N_15796);
and U16363 (N_16363,N_15862,N_15727);
nand U16364 (N_16364,N_15806,N_15904);
or U16365 (N_16365,N_15792,N_15733);
or U16366 (N_16366,N_15971,N_15914);
and U16367 (N_16367,N_15848,N_15780);
nand U16368 (N_16368,N_15693,N_15647);
nand U16369 (N_16369,N_15939,N_15903);
nand U16370 (N_16370,N_15769,N_15655);
xnor U16371 (N_16371,N_15659,N_15679);
xor U16372 (N_16372,N_15955,N_15847);
nand U16373 (N_16373,N_15994,N_15961);
xor U16374 (N_16374,N_15684,N_15766);
xnor U16375 (N_16375,N_15670,N_15972);
xor U16376 (N_16376,N_15916,N_15872);
or U16377 (N_16377,N_15875,N_15734);
xor U16378 (N_16378,N_15827,N_15817);
nor U16379 (N_16379,N_15963,N_15947);
nor U16380 (N_16380,N_15988,N_15879);
nor U16381 (N_16381,N_15998,N_15759);
nor U16382 (N_16382,N_15654,N_15953);
or U16383 (N_16383,N_15730,N_15974);
and U16384 (N_16384,N_15773,N_15658);
nand U16385 (N_16385,N_15996,N_15917);
or U16386 (N_16386,N_15946,N_15964);
nor U16387 (N_16387,N_15735,N_15949);
nor U16388 (N_16388,N_15900,N_15901);
and U16389 (N_16389,N_15872,N_15748);
xnor U16390 (N_16390,N_15624,N_15600);
and U16391 (N_16391,N_15869,N_15821);
xor U16392 (N_16392,N_15753,N_15653);
or U16393 (N_16393,N_15900,N_15841);
nor U16394 (N_16394,N_15796,N_15637);
and U16395 (N_16395,N_15661,N_15800);
and U16396 (N_16396,N_15840,N_15703);
or U16397 (N_16397,N_15898,N_15631);
and U16398 (N_16398,N_15937,N_15907);
nand U16399 (N_16399,N_15911,N_15630);
nor U16400 (N_16400,N_16247,N_16240);
or U16401 (N_16401,N_16371,N_16110);
or U16402 (N_16402,N_16094,N_16327);
and U16403 (N_16403,N_16287,N_16102);
xor U16404 (N_16404,N_16289,N_16333);
xor U16405 (N_16405,N_16085,N_16058);
xnor U16406 (N_16406,N_16356,N_16395);
or U16407 (N_16407,N_16210,N_16391);
and U16408 (N_16408,N_16388,N_16338);
nor U16409 (N_16409,N_16393,N_16115);
nor U16410 (N_16410,N_16186,N_16031);
xor U16411 (N_16411,N_16138,N_16100);
nor U16412 (N_16412,N_16321,N_16153);
and U16413 (N_16413,N_16343,N_16350);
nor U16414 (N_16414,N_16398,N_16000);
or U16415 (N_16415,N_16184,N_16368);
xor U16416 (N_16416,N_16317,N_16179);
nor U16417 (N_16417,N_16378,N_16218);
and U16418 (N_16418,N_16029,N_16018);
nand U16419 (N_16419,N_16112,N_16224);
or U16420 (N_16420,N_16047,N_16020);
nor U16421 (N_16421,N_16380,N_16004);
nor U16422 (N_16422,N_16107,N_16349);
xnor U16423 (N_16423,N_16335,N_16003);
nor U16424 (N_16424,N_16387,N_16297);
or U16425 (N_16425,N_16011,N_16290);
xnor U16426 (N_16426,N_16012,N_16131);
and U16427 (N_16427,N_16352,N_16062);
and U16428 (N_16428,N_16304,N_16291);
xnor U16429 (N_16429,N_16078,N_16330);
nor U16430 (N_16430,N_16353,N_16175);
nand U16431 (N_16431,N_16119,N_16363);
nor U16432 (N_16432,N_16268,N_16019);
nand U16433 (N_16433,N_16250,N_16208);
or U16434 (N_16434,N_16374,N_16169);
and U16435 (N_16435,N_16162,N_16278);
xnor U16436 (N_16436,N_16201,N_16167);
nand U16437 (N_16437,N_16384,N_16063);
or U16438 (N_16438,N_16230,N_16339);
or U16439 (N_16439,N_16344,N_16254);
or U16440 (N_16440,N_16303,N_16067);
xnor U16441 (N_16441,N_16358,N_16193);
or U16442 (N_16442,N_16015,N_16150);
or U16443 (N_16443,N_16315,N_16068);
or U16444 (N_16444,N_16377,N_16347);
nor U16445 (N_16445,N_16281,N_16166);
nor U16446 (N_16446,N_16164,N_16301);
and U16447 (N_16447,N_16209,N_16027);
nand U16448 (N_16448,N_16087,N_16360);
nand U16449 (N_16449,N_16362,N_16014);
nand U16450 (N_16450,N_16312,N_16373);
and U16451 (N_16451,N_16043,N_16271);
nor U16452 (N_16452,N_16065,N_16354);
nand U16453 (N_16453,N_16196,N_16013);
nor U16454 (N_16454,N_16030,N_16361);
nand U16455 (N_16455,N_16021,N_16390);
or U16456 (N_16456,N_16285,N_16049);
and U16457 (N_16457,N_16288,N_16205);
nand U16458 (N_16458,N_16274,N_16308);
nand U16459 (N_16459,N_16194,N_16149);
nand U16460 (N_16460,N_16079,N_16109);
and U16461 (N_16461,N_16171,N_16341);
or U16462 (N_16462,N_16096,N_16222);
or U16463 (N_16463,N_16090,N_16324);
nor U16464 (N_16464,N_16123,N_16242);
xnor U16465 (N_16465,N_16156,N_16044);
xnor U16466 (N_16466,N_16351,N_16323);
or U16467 (N_16467,N_16147,N_16348);
nor U16468 (N_16468,N_16234,N_16200);
or U16469 (N_16469,N_16113,N_16296);
nor U16470 (N_16470,N_16061,N_16280);
or U16471 (N_16471,N_16367,N_16117);
nor U16472 (N_16472,N_16128,N_16039);
nor U16473 (N_16473,N_16105,N_16266);
and U16474 (N_16474,N_16091,N_16257);
xnor U16475 (N_16475,N_16041,N_16237);
xnor U16476 (N_16476,N_16163,N_16177);
xor U16477 (N_16477,N_16264,N_16006);
xor U16478 (N_16478,N_16051,N_16155);
and U16479 (N_16479,N_16040,N_16217);
or U16480 (N_16480,N_16396,N_16046);
or U16481 (N_16481,N_16111,N_16122);
nand U16482 (N_16482,N_16220,N_16305);
nor U16483 (N_16483,N_16260,N_16229);
nor U16484 (N_16484,N_16146,N_16001);
nand U16485 (N_16485,N_16081,N_16397);
nor U16486 (N_16486,N_16252,N_16121);
and U16487 (N_16487,N_16139,N_16136);
xor U16488 (N_16488,N_16202,N_16060);
xnor U16489 (N_16489,N_16097,N_16292);
or U16490 (N_16490,N_16174,N_16140);
nor U16491 (N_16491,N_16022,N_16314);
or U16492 (N_16492,N_16069,N_16256);
xnor U16493 (N_16493,N_16231,N_16355);
nand U16494 (N_16494,N_16190,N_16227);
nand U16495 (N_16495,N_16346,N_16244);
or U16496 (N_16496,N_16099,N_16007);
and U16497 (N_16497,N_16212,N_16269);
nand U16498 (N_16498,N_16050,N_16165);
and U16499 (N_16499,N_16072,N_16307);
nand U16500 (N_16500,N_16214,N_16086);
nor U16501 (N_16501,N_16036,N_16197);
or U16502 (N_16502,N_16232,N_16326);
nand U16503 (N_16503,N_16071,N_16319);
nor U16504 (N_16504,N_16009,N_16249);
and U16505 (N_16505,N_16127,N_16313);
nand U16506 (N_16506,N_16369,N_16033);
and U16507 (N_16507,N_16238,N_16318);
and U16508 (N_16508,N_16026,N_16191);
xnor U16509 (N_16509,N_16253,N_16074);
xor U16510 (N_16510,N_16261,N_16028);
nor U16511 (N_16511,N_16137,N_16016);
nand U16512 (N_16512,N_16059,N_16302);
nand U16513 (N_16513,N_16080,N_16057);
xor U16514 (N_16514,N_16056,N_16328);
nand U16515 (N_16515,N_16219,N_16221);
or U16516 (N_16516,N_16160,N_16322);
xnor U16517 (N_16517,N_16054,N_16106);
xor U16518 (N_16518,N_16394,N_16329);
or U16519 (N_16519,N_16134,N_16337);
nor U16520 (N_16520,N_16265,N_16332);
xnor U16521 (N_16521,N_16089,N_16216);
nor U16522 (N_16522,N_16204,N_16181);
and U16523 (N_16523,N_16273,N_16005);
or U16524 (N_16524,N_16215,N_16255);
nand U16525 (N_16525,N_16392,N_16295);
xor U16526 (N_16526,N_16226,N_16277);
xnor U16527 (N_16527,N_16262,N_16206);
and U16528 (N_16528,N_16211,N_16176);
xnor U16529 (N_16529,N_16294,N_16172);
nor U16530 (N_16530,N_16104,N_16383);
xor U16531 (N_16531,N_16083,N_16189);
nor U16532 (N_16532,N_16108,N_16084);
or U16533 (N_16533,N_16236,N_16093);
or U16534 (N_16534,N_16366,N_16299);
nand U16535 (N_16535,N_16185,N_16331);
nor U16536 (N_16536,N_16142,N_16251);
and U16537 (N_16537,N_16235,N_16376);
or U16538 (N_16538,N_16372,N_16188);
or U16539 (N_16539,N_16073,N_16263);
nand U16540 (N_16540,N_16259,N_16114);
and U16541 (N_16541,N_16125,N_16141);
nand U16542 (N_16542,N_16055,N_16035);
nor U16543 (N_16543,N_16316,N_16286);
nand U16544 (N_16544,N_16239,N_16311);
nor U16545 (N_16545,N_16048,N_16038);
nand U16546 (N_16546,N_16382,N_16066);
nor U16547 (N_16547,N_16270,N_16075);
xor U16548 (N_16548,N_16379,N_16053);
and U16549 (N_16549,N_16023,N_16245);
or U16550 (N_16550,N_16248,N_16076);
xor U16551 (N_16551,N_16070,N_16325);
nand U16552 (N_16552,N_16152,N_16300);
and U16553 (N_16553,N_16157,N_16017);
and U16554 (N_16554,N_16203,N_16275);
nand U16555 (N_16555,N_16276,N_16381);
nand U16556 (N_16556,N_16283,N_16385);
xnor U16557 (N_16557,N_16243,N_16340);
or U16558 (N_16558,N_16133,N_16187);
xor U16559 (N_16559,N_16144,N_16306);
or U16560 (N_16560,N_16183,N_16130);
nor U16561 (N_16561,N_16182,N_16207);
nand U16562 (N_16562,N_16399,N_16284);
xnor U16563 (N_16563,N_16225,N_16077);
nand U16564 (N_16564,N_16132,N_16034);
xor U16565 (N_16565,N_16145,N_16195);
nor U16566 (N_16566,N_16135,N_16389);
nand U16567 (N_16567,N_16101,N_16334);
xnor U16568 (N_16568,N_16088,N_16223);
xor U16569 (N_16569,N_16052,N_16143);
nand U16570 (N_16570,N_16320,N_16258);
nor U16571 (N_16571,N_16116,N_16168);
xnor U16572 (N_16572,N_16279,N_16199);
nand U16573 (N_16573,N_16233,N_16148);
nand U16574 (N_16574,N_16129,N_16310);
and U16575 (N_16575,N_16092,N_16364);
nor U16576 (N_16576,N_16386,N_16158);
nand U16577 (N_16577,N_16154,N_16282);
and U16578 (N_16578,N_16098,N_16151);
xnor U16579 (N_16579,N_16298,N_16359);
nor U16580 (N_16580,N_16042,N_16025);
or U16581 (N_16581,N_16002,N_16008);
nand U16582 (N_16582,N_16213,N_16010);
and U16583 (N_16583,N_16082,N_16118);
and U16584 (N_16584,N_16064,N_16045);
nand U16585 (N_16585,N_16120,N_16095);
nor U16586 (N_16586,N_16267,N_16032);
and U16587 (N_16587,N_16309,N_16024);
nand U16588 (N_16588,N_16037,N_16180);
nand U16589 (N_16589,N_16103,N_16246);
or U16590 (N_16590,N_16272,N_16198);
nor U16591 (N_16591,N_16124,N_16241);
nand U16592 (N_16592,N_16178,N_16161);
nand U16593 (N_16593,N_16192,N_16159);
xnor U16594 (N_16594,N_16342,N_16126);
and U16595 (N_16595,N_16357,N_16170);
nand U16596 (N_16596,N_16336,N_16375);
xor U16597 (N_16597,N_16293,N_16173);
nand U16598 (N_16598,N_16365,N_16370);
nor U16599 (N_16599,N_16228,N_16345);
or U16600 (N_16600,N_16006,N_16266);
nand U16601 (N_16601,N_16206,N_16325);
xnor U16602 (N_16602,N_16188,N_16338);
and U16603 (N_16603,N_16349,N_16261);
nand U16604 (N_16604,N_16360,N_16238);
and U16605 (N_16605,N_16342,N_16176);
nor U16606 (N_16606,N_16306,N_16210);
nand U16607 (N_16607,N_16152,N_16328);
and U16608 (N_16608,N_16304,N_16294);
nor U16609 (N_16609,N_16071,N_16031);
or U16610 (N_16610,N_16168,N_16350);
or U16611 (N_16611,N_16247,N_16368);
nor U16612 (N_16612,N_16385,N_16220);
xnor U16613 (N_16613,N_16265,N_16015);
or U16614 (N_16614,N_16395,N_16010);
xnor U16615 (N_16615,N_16010,N_16044);
nand U16616 (N_16616,N_16181,N_16103);
nand U16617 (N_16617,N_16264,N_16300);
and U16618 (N_16618,N_16293,N_16214);
xnor U16619 (N_16619,N_16257,N_16258);
nand U16620 (N_16620,N_16371,N_16002);
nor U16621 (N_16621,N_16234,N_16000);
or U16622 (N_16622,N_16051,N_16276);
nand U16623 (N_16623,N_16168,N_16134);
or U16624 (N_16624,N_16341,N_16245);
or U16625 (N_16625,N_16070,N_16209);
nand U16626 (N_16626,N_16302,N_16005);
xnor U16627 (N_16627,N_16111,N_16117);
nor U16628 (N_16628,N_16105,N_16385);
nor U16629 (N_16629,N_16297,N_16356);
nor U16630 (N_16630,N_16358,N_16277);
nor U16631 (N_16631,N_16027,N_16112);
xnor U16632 (N_16632,N_16030,N_16273);
and U16633 (N_16633,N_16106,N_16376);
xnor U16634 (N_16634,N_16144,N_16237);
and U16635 (N_16635,N_16176,N_16399);
and U16636 (N_16636,N_16158,N_16243);
nor U16637 (N_16637,N_16282,N_16142);
and U16638 (N_16638,N_16330,N_16344);
nor U16639 (N_16639,N_16233,N_16311);
nor U16640 (N_16640,N_16377,N_16397);
and U16641 (N_16641,N_16031,N_16118);
nand U16642 (N_16642,N_16069,N_16138);
nand U16643 (N_16643,N_16347,N_16152);
nor U16644 (N_16644,N_16297,N_16197);
xnor U16645 (N_16645,N_16185,N_16089);
xor U16646 (N_16646,N_16094,N_16247);
xnor U16647 (N_16647,N_16157,N_16243);
nand U16648 (N_16648,N_16200,N_16184);
nand U16649 (N_16649,N_16332,N_16045);
and U16650 (N_16650,N_16164,N_16195);
and U16651 (N_16651,N_16286,N_16372);
and U16652 (N_16652,N_16142,N_16101);
xnor U16653 (N_16653,N_16039,N_16158);
and U16654 (N_16654,N_16093,N_16044);
or U16655 (N_16655,N_16028,N_16385);
and U16656 (N_16656,N_16340,N_16038);
or U16657 (N_16657,N_16298,N_16120);
or U16658 (N_16658,N_16282,N_16106);
or U16659 (N_16659,N_16088,N_16310);
and U16660 (N_16660,N_16191,N_16174);
xor U16661 (N_16661,N_16209,N_16061);
or U16662 (N_16662,N_16120,N_16371);
and U16663 (N_16663,N_16014,N_16000);
nor U16664 (N_16664,N_16232,N_16317);
nand U16665 (N_16665,N_16036,N_16364);
or U16666 (N_16666,N_16291,N_16068);
nor U16667 (N_16667,N_16257,N_16127);
or U16668 (N_16668,N_16318,N_16202);
xnor U16669 (N_16669,N_16094,N_16240);
xnor U16670 (N_16670,N_16320,N_16218);
or U16671 (N_16671,N_16287,N_16004);
or U16672 (N_16672,N_16117,N_16182);
nor U16673 (N_16673,N_16153,N_16083);
or U16674 (N_16674,N_16205,N_16043);
and U16675 (N_16675,N_16021,N_16357);
nand U16676 (N_16676,N_16315,N_16059);
and U16677 (N_16677,N_16128,N_16200);
or U16678 (N_16678,N_16263,N_16074);
and U16679 (N_16679,N_16157,N_16046);
nand U16680 (N_16680,N_16204,N_16293);
or U16681 (N_16681,N_16249,N_16064);
nand U16682 (N_16682,N_16338,N_16098);
or U16683 (N_16683,N_16092,N_16130);
nor U16684 (N_16684,N_16116,N_16157);
and U16685 (N_16685,N_16287,N_16054);
and U16686 (N_16686,N_16073,N_16146);
and U16687 (N_16687,N_16221,N_16332);
nand U16688 (N_16688,N_16326,N_16112);
xor U16689 (N_16689,N_16025,N_16113);
xor U16690 (N_16690,N_16344,N_16122);
or U16691 (N_16691,N_16312,N_16126);
or U16692 (N_16692,N_16257,N_16042);
and U16693 (N_16693,N_16283,N_16367);
and U16694 (N_16694,N_16386,N_16077);
and U16695 (N_16695,N_16083,N_16166);
and U16696 (N_16696,N_16378,N_16177);
nor U16697 (N_16697,N_16180,N_16292);
or U16698 (N_16698,N_16185,N_16018);
xnor U16699 (N_16699,N_16236,N_16152);
nand U16700 (N_16700,N_16317,N_16160);
nor U16701 (N_16701,N_16124,N_16187);
nand U16702 (N_16702,N_16188,N_16370);
xnor U16703 (N_16703,N_16110,N_16216);
or U16704 (N_16704,N_16340,N_16275);
and U16705 (N_16705,N_16391,N_16191);
nand U16706 (N_16706,N_16067,N_16129);
and U16707 (N_16707,N_16311,N_16279);
and U16708 (N_16708,N_16220,N_16214);
or U16709 (N_16709,N_16235,N_16140);
nor U16710 (N_16710,N_16166,N_16204);
nand U16711 (N_16711,N_16128,N_16028);
nand U16712 (N_16712,N_16213,N_16078);
nor U16713 (N_16713,N_16282,N_16152);
nor U16714 (N_16714,N_16366,N_16342);
and U16715 (N_16715,N_16231,N_16317);
and U16716 (N_16716,N_16247,N_16325);
or U16717 (N_16717,N_16104,N_16243);
nor U16718 (N_16718,N_16167,N_16398);
xnor U16719 (N_16719,N_16051,N_16345);
nand U16720 (N_16720,N_16360,N_16279);
xnor U16721 (N_16721,N_16278,N_16135);
or U16722 (N_16722,N_16326,N_16340);
nor U16723 (N_16723,N_16353,N_16284);
or U16724 (N_16724,N_16188,N_16388);
nor U16725 (N_16725,N_16325,N_16382);
xnor U16726 (N_16726,N_16353,N_16339);
and U16727 (N_16727,N_16277,N_16334);
xnor U16728 (N_16728,N_16064,N_16305);
and U16729 (N_16729,N_16078,N_16297);
or U16730 (N_16730,N_16084,N_16013);
and U16731 (N_16731,N_16350,N_16371);
nand U16732 (N_16732,N_16007,N_16329);
nand U16733 (N_16733,N_16075,N_16353);
xor U16734 (N_16734,N_16204,N_16147);
nand U16735 (N_16735,N_16136,N_16120);
nor U16736 (N_16736,N_16022,N_16180);
or U16737 (N_16737,N_16128,N_16060);
and U16738 (N_16738,N_16324,N_16061);
or U16739 (N_16739,N_16377,N_16369);
and U16740 (N_16740,N_16066,N_16079);
and U16741 (N_16741,N_16212,N_16103);
and U16742 (N_16742,N_16174,N_16329);
nand U16743 (N_16743,N_16375,N_16305);
and U16744 (N_16744,N_16375,N_16123);
nor U16745 (N_16745,N_16315,N_16169);
xor U16746 (N_16746,N_16141,N_16360);
or U16747 (N_16747,N_16313,N_16159);
or U16748 (N_16748,N_16012,N_16169);
nor U16749 (N_16749,N_16172,N_16292);
nand U16750 (N_16750,N_16202,N_16191);
xnor U16751 (N_16751,N_16341,N_16152);
and U16752 (N_16752,N_16182,N_16258);
and U16753 (N_16753,N_16037,N_16090);
or U16754 (N_16754,N_16100,N_16363);
or U16755 (N_16755,N_16327,N_16266);
nand U16756 (N_16756,N_16084,N_16080);
or U16757 (N_16757,N_16088,N_16172);
nand U16758 (N_16758,N_16249,N_16087);
xor U16759 (N_16759,N_16016,N_16091);
and U16760 (N_16760,N_16153,N_16110);
and U16761 (N_16761,N_16130,N_16246);
or U16762 (N_16762,N_16156,N_16329);
and U16763 (N_16763,N_16156,N_16047);
nor U16764 (N_16764,N_16125,N_16014);
xor U16765 (N_16765,N_16199,N_16287);
nor U16766 (N_16766,N_16307,N_16101);
nand U16767 (N_16767,N_16116,N_16127);
or U16768 (N_16768,N_16089,N_16301);
or U16769 (N_16769,N_16172,N_16052);
and U16770 (N_16770,N_16281,N_16025);
or U16771 (N_16771,N_16082,N_16023);
xnor U16772 (N_16772,N_16268,N_16112);
nand U16773 (N_16773,N_16144,N_16198);
nor U16774 (N_16774,N_16267,N_16155);
or U16775 (N_16775,N_16001,N_16174);
xnor U16776 (N_16776,N_16396,N_16197);
nand U16777 (N_16777,N_16170,N_16217);
nor U16778 (N_16778,N_16108,N_16080);
xor U16779 (N_16779,N_16310,N_16261);
nand U16780 (N_16780,N_16109,N_16389);
xor U16781 (N_16781,N_16147,N_16167);
nor U16782 (N_16782,N_16153,N_16105);
nor U16783 (N_16783,N_16325,N_16024);
or U16784 (N_16784,N_16060,N_16045);
or U16785 (N_16785,N_16383,N_16177);
xor U16786 (N_16786,N_16298,N_16178);
nor U16787 (N_16787,N_16391,N_16144);
nand U16788 (N_16788,N_16084,N_16229);
nand U16789 (N_16789,N_16381,N_16246);
or U16790 (N_16790,N_16353,N_16357);
and U16791 (N_16791,N_16288,N_16067);
nand U16792 (N_16792,N_16222,N_16048);
and U16793 (N_16793,N_16255,N_16052);
nor U16794 (N_16794,N_16357,N_16129);
nor U16795 (N_16795,N_16346,N_16386);
nor U16796 (N_16796,N_16145,N_16082);
nand U16797 (N_16797,N_16230,N_16301);
nand U16798 (N_16798,N_16352,N_16094);
nand U16799 (N_16799,N_16367,N_16159);
xnor U16800 (N_16800,N_16482,N_16608);
xnor U16801 (N_16801,N_16424,N_16712);
and U16802 (N_16802,N_16682,N_16427);
nor U16803 (N_16803,N_16791,N_16683);
or U16804 (N_16804,N_16741,N_16774);
xor U16805 (N_16805,N_16465,N_16722);
nor U16806 (N_16806,N_16744,N_16525);
xor U16807 (N_16807,N_16733,N_16616);
nor U16808 (N_16808,N_16438,N_16689);
nand U16809 (N_16809,N_16555,N_16495);
nor U16810 (N_16810,N_16662,N_16658);
nand U16811 (N_16811,N_16526,N_16640);
nand U16812 (N_16812,N_16556,N_16634);
or U16813 (N_16813,N_16789,N_16700);
or U16814 (N_16814,N_16579,N_16701);
and U16815 (N_16815,N_16422,N_16594);
nor U16816 (N_16816,N_16708,N_16740);
and U16817 (N_16817,N_16448,N_16778);
and U16818 (N_16818,N_16549,N_16463);
or U16819 (N_16819,N_16528,N_16641);
nor U16820 (N_16820,N_16583,N_16726);
nor U16821 (N_16821,N_16721,N_16564);
xnor U16822 (N_16822,N_16685,N_16665);
nand U16823 (N_16823,N_16512,N_16677);
or U16824 (N_16824,N_16418,N_16739);
nor U16825 (N_16825,N_16439,N_16420);
nand U16826 (N_16826,N_16470,N_16704);
nand U16827 (N_16827,N_16590,N_16647);
nor U16828 (N_16828,N_16478,N_16612);
and U16829 (N_16829,N_16725,N_16419);
nand U16830 (N_16830,N_16757,N_16500);
and U16831 (N_16831,N_16593,N_16676);
nand U16832 (N_16832,N_16591,N_16751);
nor U16833 (N_16833,N_16796,N_16713);
or U16834 (N_16834,N_16553,N_16717);
or U16835 (N_16835,N_16409,N_16541);
xor U16836 (N_16836,N_16576,N_16562);
and U16837 (N_16837,N_16643,N_16496);
nor U16838 (N_16838,N_16492,N_16669);
nand U16839 (N_16839,N_16567,N_16674);
or U16840 (N_16840,N_16570,N_16639);
xnor U16841 (N_16841,N_16601,N_16698);
or U16842 (N_16842,N_16693,N_16606);
xnor U16843 (N_16843,N_16732,N_16724);
nor U16844 (N_16844,N_16780,N_16628);
and U16845 (N_16845,N_16573,N_16670);
nand U16846 (N_16846,N_16637,N_16715);
nand U16847 (N_16847,N_16550,N_16679);
nor U16848 (N_16848,N_16401,N_16776);
or U16849 (N_16849,N_16750,N_16431);
nor U16850 (N_16850,N_16460,N_16652);
and U16851 (N_16851,N_16527,N_16445);
or U16852 (N_16852,N_16477,N_16772);
nor U16853 (N_16853,N_16582,N_16481);
or U16854 (N_16854,N_16441,N_16755);
nor U16855 (N_16855,N_16430,N_16655);
nor U16856 (N_16856,N_16544,N_16629);
nand U16857 (N_16857,N_16417,N_16534);
nor U16858 (N_16858,N_16517,N_16554);
nand U16859 (N_16859,N_16644,N_16506);
nand U16860 (N_16860,N_16766,N_16488);
nand U16861 (N_16861,N_16660,N_16692);
xnor U16862 (N_16862,N_16585,N_16672);
xnor U16863 (N_16863,N_16485,N_16603);
or U16864 (N_16864,N_16552,N_16691);
or U16865 (N_16865,N_16648,N_16519);
or U16866 (N_16866,N_16649,N_16656);
nand U16867 (N_16867,N_16786,N_16416);
or U16868 (N_16868,N_16747,N_16636);
nor U16869 (N_16869,N_16650,N_16461);
nand U16870 (N_16870,N_16530,N_16421);
and U16871 (N_16871,N_16560,N_16535);
nor U16872 (N_16872,N_16408,N_16444);
and U16873 (N_16873,N_16613,N_16602);
xnor U16874 (N_16874,N_16735,N_16542);
nand U16875 (N_16875,N_16671,N_16632);
xor U16876 (N_16876,N_16615,N_16547);
nand U16877 (N_16877,N_16497,N_16673);
and U16878 (N_16878,N_16773,N_16799);
or U16879 (N_16879,N_16754,N_16523);
nand U16880 (N_16880,N_16437,N_16659);
or U16881 (N_16881,N_16472,N_16710);
or U16882 (N_16882,N_16756,N_16548);
or U16883 (N_16883,N_16475,N_16667);
nor U16884 (N_16884,N_16759,N_16455);
xor U16885 (N_16885,N_16546,N_16447);
and U16886 (N_16886,N_16404,N_16785);
or U16887 (N_16887,N_16425,N_16462);
nor U16888 (N_16888,N_16574,N_16716);
or U16889 (N_16889,N_16738,N_16620);
nor U16890 (N_16890,N_16473,N_16469);
and U16891 (N_16891,N_16454,N_16787);
and U16892 (N_16892,N_16737,N_16749);
or U16893 (N_16893,N_16723,N_16531);
and U16894 (N_16894,N_16705,N_16697);
or U16895 (N_16895,N_16588,N_16743);
or U16896 (N_16896,N_16630,N_16798);
and U16897 (N_16897,N_16764,N_16696);
nor U16898 (N_16898,N_16433,N_16503);
xor U16899 (N_16899,N_16436,N_16578);
and U16900 (N_16900,N_16719,N_16633);
xor U16901 (N_16901,N_16501,N_16742);
and U16902 (N_16902,N_16451,N_16728);
nor U16903 (N_16903,N_16779,N_16680);
nor U16904 (N_16904,N_16790,N_16551);
nor U16905 (N_16905,N_16611,N_16638);
nand U16906 (N_16906,N_16592,N_16782);
nor U16907 (N_16907,N_16626,N_16442);
nand U16908 (N_16908,N_16484,N_16609);
nor U16909 (N_16909,N_16440,N_16498);
xnor U16910 (N_16910,N_16642,N_16449);
nor U16911 (N_16911,N_16577,N_16489);
nor U16912 (N_16912,N_16605,N_16734);
and U16913 (N_16913,N_16699,N_16758);
nor U16914 (N_16914,N_16761,N_16543);
xnor U16915 (N_16915,N_16707,N_16456);
nor U16916 (N_16916,N_16794,N_16529);
nor U16917 (N_16917,N_16486,N_16405);
and U16918 (N_16918,N_16645,N_16411);
nand U16919 (N_16919,N_16703,N_16494);
nor U16920 (N_16920,N_16664,N_16539);
or U16921 (N_16921,N_16748,N_16533);
and U16922 (N_16922,N_16797,N_16596);
xor U16923 (N_16923,N_16599,N_16627);
nand U16924 (N_16924,N_16619,N_16770);
nor U16925 (N_16925,N_16793,N_16572);
or U16926 (N_16926,N_16480,N_16400);
nor U16927 (N_16927,N_16631,N_16635);
nand U16928 (N_16928,N_16537,N_16413);
nor U16929 (N_16929,N_16769,N_16536);
or U16930 (N_16930,N_16580,N_16792);
xor U16931 (N_16931,N_16760,N_16557);
or U16932 (N_16932,N_16458,N_16471);
nand U16933 (N_16933,N_16520,N_16403);
and U16934 (N_16934,N_16688,N_16625);
and U16935 (N_16935,N_16654,N_16502);
nor U16936 (N_16936,N_16614,N_16563);
xor U16937 (N_16937,N_16663,N_16435);
or U16938 (N_16938,N_16777,N_16452);
and U16939 (N_16939,N_16571,N_16684);
nor U16940 (N_16940,N_16414,N_16622);
nor U16941 (N_16941,N_16657,N_16511);
xor U16942 (N_16942,N_16651,N_16666);
xnor U16943 (N_16943,N_16595,N_16788);
and U16944 (N_16944,N_16407,N_16402);
or U16945 (N_16945,N_16604,N_16711);
nand U16946 (N_16946,N_16493,N_16607);
or U16947 (N_16947,N_16709,N_16457);
nor U16948 (N_16948,N_16781,N_16767);
nand U16949 (N_16949,N_16623,N_16597);
or U16950 (N_16950,N_16569,N_16505);
and U16951 (N_16951,N_16428,N_16730);
nor U16952 (N_16952,N_16443,N_16516);
or U16953 (N_16953,N_16775,N_16762);
or U16954 (N_16954,N_16474,N_16745);
nand U16955 (N_16955,N_16598,N_16540);
xor U16956 (N_16956,N_16765,N_16575);
and U16957 (N_16957,N_16624,N_16718);
xnor U16958 (N_16958,N_16499,N_16412);
nand U16959 (N_16959,N_16784,N_16459);
and U16960 (N_16960,N_16686,N_16600);
and U16961 (N_16961,N_16490,N_16771);
and U16962 (N_16962,N_16695,N_16694);
nand U16963 (N_16963,N_16690,N_16746);
or U16964 (N_16964,N_16464,N_16558);
nand U16965 (N_16965,N_16432,N_16565);
nor U16966 (N_16966,N_16518,N_16584);
xnor U16967 (N_16967,N_16727,N_16508);
nand U16968 (N_16968,N_16736,N_16678);
nand U16969 (N_16969,N_16661,N_16668);
or U16970 (N_16970,N_16752,N_16687);
xnor U16971 (N_16971,N_16426,N_16646);
xnor U16972 (N_16972,N_16423,N_16681);
nand U16973 (N_16973,N_16446,N_16406);
nand U16974 (N_16974,N_16453,N_16434);
xnor U16975 (N_16975,N_16783,N_16504);
nand U16976 (N_16976,N_16618,N_16429);
nand U16977 (N_16977,N_16491,N_16487);
or U16978 (N_16978,N_16653,N_16510);
nand U16979 (N_16979,N_16410,N_16522);
nor U16980 (N_16980,N_16706,N_16476);
xnor U16981 (N_16981,N_16768,N_16514);
nor U16982 (N_16982,N_16589,N_16513);
nand U16983 (N_16983,N_16532,N_16763);
and U16984 (N_16984,N_16515,N_16720);
xor U16985 (N_16985,N_16509,N_16731);
nand U16986 (N_16986,N_16617,N_16507);
nor U16987 (N_16987,N_16729,N_16415);
nor U16988 (N_16988,N_16559,N_16714);
nand U16989 (N_16989,N_16675,N_16621);
or U16990 (N_16990,N_16479,N_16524);
xnor U16991 (N_16991,N_16753,N_16795);
nand U16992 (N_16992,N_16587,N_16545);
nor U16993 (N_16993,N_16467,N_16521);
nor U16994 (N_16994,N_16566,N_16466);
nand U16995 (N_16995,N_16538,N_16581);
or U16996 (N_16996,N_16610,N_16468);
nor U16997 (N_16997,N_16450,N_16702);
xor U16998 (N_16998,N_16483,N_16568);
and U16999 (N_16999,N_16586,N_16561);
xnor U17000 (N_17000,N_16593,N_16477);
nor U17001 (N_17001,N_16534,N_16433);
nand U17002 (N_17002,N_16428,N_16536);
and U17003 (N_17003,N_16532,N_16639);
nand U17004 (N_17004,N_16401,N_16732);
or U17005 (N_17005,N_16714,N_16639);
nor U17006 (N_17006,N_16692,N_16791);
xor U17007 (N_17007,N_16498,N_16721);
and U17008 (N_17008,N_16606,N_16481);
or U17009 (N_17009,N_16718,N_16584);
xnor U17010 (N_17010,N_16595,N_16460);
and U17011 (N_17011,N_16761,N_16601);
or U17012 (N_17012,N_16596,N_16529);
nor U17013 (N_17013,N_16443,N_16686);
or U17014 (N_17014,N_16434,N_16538);
xor U17015 (N_17015,N_16555,N_16715);
nor U17016 (N_17016,N_16777,N_16559);
nand U17017 (N_17017,N_16476,N_16664);
or U17018 (N_17018,N_16742,N_16488);
or U17019 (N_17019,N_16730,N_16522);
and U17020 (N_17020,N_16489,N_16782);
or U17021 (N_17021,N_16740,N_16761);
nor U17022 (N_17022,N_16569,N_16422);
nor U17023 (N_17023,N_16641,N_16755);
and U17024 (N_17024,N_16492,N_16755);
xor U17025 (N_17025,N_16700,N_16777);
and U17026 (N_17026,N_16513,N_16568);
and U17027 (N_17027,N_16500,N_16592);
and U17028 (N_17028,N_16738,N_16570);
nand U17029 (N_17029,N_16753,N_16636);
xnor U17030 (N_17030,N_16787,N_16580);
or U17031 (N_17031,N_16593,N_16720);
xnor U17032 (N_17032,N_16480,N_16634);
or U17033 (N_17033,N_16767,N_16423);
nand U17034 (N_17034,N_16488,N_16422);
or U17035 (N_17035,N_16501,N_16657);
or U17036 (N_17036,N_16749,N_16540);
or U17037 (N_17037,N_16445,N_16555);
nand U17038 (N_17038,N_16414,N_16600);
or U17039 (N_17039,N_16724,N_16787);
and U17040 (N_17040,N_16773,N_16449);
xor U17041 (N_17041,N_16515,N_16776);
or U17042 (N_17042,N_16676,N_16751);
and U17043 (N_17043,N_16759,N_16543);
or U17044 (N_17044,N_16572,N_16555);
nand U17045 (N_17045,N_16523,N_16675);
nand U17046 (N_17046,N_16580,N_16570);
and U17047 (N_17047,N_16536,N_16623);
nor U17048 (N_17048,N_16599,N_16411);
nor U17049 (N_17049,N_16769,N_16785);
nor U17050 (N_17050,N_16748,N_16506);
or U17051 (N_17051,N_16436,N_16765);
and U17052 (N_17052,N_16571,N_16762);
and U17053 (N_17053,N_16705,N_16673);
xor U17054 (N_17054,N_16787,N_16681);
and U17055 (N_17055,N_16455,N_16789);
xor U17056 (N_17056,N_16428,N_16676);
and U17057 (N_17057,N_16666,N_16787);
or U17058 (N_17058,N_16722,N_16695);
nand U17059 (N_17059,N_16698,N_16700);
nand U17060 (N_17060,N_16713,N_16778);
and U17061 (N_17061,N_16617,N_16575);
or U17062 (N_17062,N_16682,N_16669);
or U17063 (N_17063,N_16639,N_16410);
or U17064 (N_17064,N_16679,N_16496);
xnor U17065 (N_17065,N_16752,N_16447);
and U17066 (N_17066,N_16576,N_16627);
or U17067 (N_17067,N_16572,N_16615);
and U17068 (N_17068,N_16433,N_16527);
nor U17069 (N_17069,N_16657,N_16678);
nor U17070 (N_17070,N_16634,N_16639);
nand U17071 (N_17071,N_16758,N_16551);
or U17072 (N_17072,N_16664,N_16509);
xnor U17073 (N_17073,N_16529,N_16555);
xnor U17074 (N_17074,N_16506,N_16780);
and U17075 (N_17075,N_16618,N_16688);
and U17076 (N_17076,N_16707,N_16538);
or U17077 (N_17077,N_16707,N_16665);
nand U17078 (N_17078,N_16735,N_16685);
xor U17079 (N_17079,N_16608,N_16648);
nand U17080 (N_17080,N_16467,N_16590);
nor U17081 (N_17081,N_16544,N_16771);
xnor U17082 (N_17082,N_16595,N_16486);
xnor U17083 (N_17083,N_16503,N_16418);
xor U17084 (N_17084,N_16474,N_16643);
nand U17085 (N_17085,N_16476,N_16403);
nor U17086 (N_17086,N_16467,N_16473);
or U17087 (N_17087,N_16745,N_16432);
nor U17088 (N_17088,N_16480,N_16711);
xnor U17089 (N_17089,N_16764,N_16742);
nand U17090 (N_17090,N_16483,N_16663);
and U17091 (N_17091,N_16798,N_16581);
xor U17092 (N_17092,N_16638,N_16551);
and U17093 (N_17093,N_16774,N_16700);
xnor U17094 (N_17094,N_16538,N_16478);
xnor U17095 (N_17095,N_16563,N_16537);
or U17096 (N_17096,N_16758,N_16455);
nor U17097 (N_17097,N_16740,N_16799);
and U17098 (N_17098,N_16708,N_16620);
and U17099 (N_17099,N_16713,N_16435);
or U17100 (N_17100,N_16606,N_16684);
nand U17101 (N_17101,N_16796,N_16471);
or U17102 (N_17102,N_16777,N_16662);
and U17103 (N_17103,N_16597,N_16765);
nand U17104 (N_17104,N_16442,N_16565);
or U17105 (N_17105,N_16508,N_16409);
or U17106 (N_17106,N_16591,N_16635);
nor U17107 (N_17107,N_16775,N_16651);
xnor U17108 (N_17108,N_16426,N_16670);
nor U17109 (N_17109,N_16505,N_16665);
and U17110 (N_17110,N_16786,N_16696);
nor U17111 (N_17111,N_16666,N_16684);
or U17112 (N_17112,N_16442,N_16747);
and U17113 (N_17113,N_16754,N_16716);
nor U17114 (N_17114,N_16561,N_16506);
xor U17115 (N_17115,N_16722,N_16528);
and U17116 (N_17116,N_16730,N_16503);
nor U17117 (N_17117,N_16665,N_16491);
nand U17118 (N_17118,N_16538,N_16769);
nand U17119 (N_17119,N_16681,N_16401);
xnor U17120 (N_17120,N_16537,N_16784);
xnor U17121 (N_17121,N_16789,N_16758);
nor U17122 (N_17122,N_16720,N_16584);
and U17123 (N_17123,N_16765,N_16756);
nor U17124 (N_17124,N_16492,N_16532);
or U17125 (N_17125,N_16655,N_16463);
and U17126 (N_17126,N_16418,N_16621);
or U17127 (N_17127,N_16571,N_16782);
nand U17128 (N_17128,N_16421,N_16491);
and U17129 (N_17129,N_16537,N_16607);
xor U17130 (N_17130,N_16587,N_16670);
xnor U17131 (N_17131,N_16693,N_16563);
xor U17132 (N_17132,N_16581,N_16675);
xor U17133 (N_17133,N_16551,N_16411);
nand U17134 (N_17134,N_16783,N_16573);
nor U17135 (N_17135,N_16420,N_16438);
and U17136 (N_17136,N_16453,N_16527);
nand U17137 (N_17137,N_16409,N_16601);
or U17138 (N_17138,N_16676,N_16687);
nand U17139 (N_17139,N_16454,N_16483);
nor U17140 (N_17140,N_16753,N_16649);
nand U17141 (N_17141,N_16609,N_16527);
xnor U17142 (N_17142,N_16526,N_16537);
xor U17143 (N_17143,N_16477,N_16686);
nor U17144 (N_17144,N_16504,N_16594);
nand U17145 (N_17145,N_16592,N_16415);
nor U17146 (N_17146,N_16523,N_16645);
nand U17147 (N_17147,N_16493,N_16772);
nand U17148 (N_17148,N_16456,N_16710);
and U17149 (N_17149,N_16516,N_16734);
xnor U17150 (N_17150,N_16530,N_16528);
and U17151 (N_17151,N_16751,N_16479);
or U17152 (N_17152,N_16424,N_16777);
nand U17153 (N_17153,N_16716,N_16429);
nand U17154 (N_17154,N_16459,N_16748);
or U17155 (N_17155,N_16584,N_16716);
xnor U17156 (N_17156,N_16522,N_16525);
nor U17157 (N_17157,N_16786,N_16606);
xor U17158 (N_17158,N_16514,N_16544);
or U17159 (N_17159,N_16444,N_16616);
or U17160 (N_17160,N_16733,N_16627);
and U17161 (N_17161,N_16416,N_16788);
nand U17162 (N_17162,N_16450,N_16609);
nand U17163 (N_17163,N_16698,N_16598);
nand U17164 (N_17164,N_16741,N_16467);
nand U17165 (N_17165,N_16620,N_16411);
nand U17166 (N_17166,N_16455,N_16749);
or U17167 (N_17167,N_16605,N_16630);
xor U17168 (N_17168,N_16668,N_16541);
or U17169 (N_17169,N_16592,N_16700);
nor U17170 (N_17170,N_16540,N_16596);
nand U17171 (N_17171,N_16634,N_16630);
nor U17172 (N_17172,N_16756,N_16536);
xnor U17173 (N_17173,N_16516,N_16621);
xor U17174 (N_17174,N_16797,N_16796);
or U17175 (N_17175,N_16536,N_16689);
or U17176 (N_17176,N_16426,N_16776);
xnor U17177 (N_17177,N_16571,N_16577);
nor U17178 (N_17178,N_16441,N_16622);
or U17179 (N_17179,N_16609,N_16797);
xnor U17180 (N_17180,N_16610,N_16605);
nand U17181 (N_17181,N_16686,N_16524);
xor U17182 (N_17182,N_16705,N_16529);
xnor U17183 (N_17183,N_16696,N_16583);
nand U17184 (N_17184,N_16670,N_16636);
nand U17185 (N_17185,N_16519,N_16624);
xor U17186 (N_17186,N_16550,N_16749);
and U17187 (N_17187,N_16469,N_16509);
and U17188 (N_17188,N_16426,N_16459);
nand U17189 (N_17189,N_16416,N_16768);
or U17190 (N_17190,N_16533,N_16660);
nor U17191 (N_17191,N_16785,N_16723);
xor U17192 (N_17192,N_16412,N_16419);
nand U17193 (N_17193,N_16565,N_16609);
and U17194 (N_17194,N_16714,N_16424);
xor U17195 (N_17195,N_16614,N_16776);
nand U17196 (N_17196,N_16738,N_16401);
or U17197 (N_17197,N_16792,N_16786);
nor U17198 (N_17198,N_16527,N_16766);
nor U17199 (N_17199,N_16639,N_16513);
xnor U17200 (N_17200,N_16920,N_16934);
and U17201 (N_17201,N_16928,N_16831);
nor U17202 (N_17202,N_17114,N_17173);
or U17203 (N_17203,N_17030,N_16885);
or U17204 (N_17204,N_16911,N_16905);
nor U17205 (N_17205,N_16816,N_16962);
and U17206 (N_17206,N_16851,N_17043);
and U17207 (N_17207,N_16985,N_17163);
nand U17208 (N_17208,N_17158,N_16890);
xor U17209 (N_17209,N_16809,N_16881);
nand U17210 (N_17210,N_17012,N_17147);
nor U17211 (N_17211,N_17088,N_17174);
nor U17212 (N_17212,N_16825,N_17191);
or U17213 (N_17213,N_16827,N_17121);
and U17214 (N_17214,N_17092,N_17045);
or U17215 (N_17215,N_16992,N_17162);
and U17216 (N_17216,N_16950,N_16823);
xor U17217 (N_17217,N_17195,N_17122);
xor U17218 (N_17218,N_16848,N_17168);
and U17219 (N_17219,N_17032,N_17148);
nand U17220 (N_17220,N_17075,N_17153);
nand U17221 (N_17221,N_16941,N_17118);
or U17222 (N_17222,N_16926,N_16804);
or U17223 (N_17223,N_16971,N_16927);
nor U17224 (N_17224,N_17181,N_16899);
nand U17225 (N_17225,N_17006,N_17116);
nand U17226 (N_17226,N_17103,N_16995);
or U17227 (N_17227,N_16967,N_16955);
nand U17228 (N_17228,N_17120,N_16930);
or U17229 (N_17229,N_17136,N_16947);
nand U17230 (N_17230,N_16964,N_17176);
nand U17231 (N_17231,N_16873,N_16918);
nor U17232 (N_17232,N_17087,N_16807);
or U17233 (N_17233,N_16843,N_17070);
nor U17234 (N_17234,N_16894,N_17094);
nor U17235 (N_17235,N_17007,N_17194);
or U17236 (N_17236,N_16876,N_17129);
and U17237 (N_17237,N_16933,N_17090);
or U17238 (N_17238,N_17076,N_17101);
nor U17239 (N_17239,N_16856,N_16915);
nand U17240 (N_17240,N_16811,N_17139);
and U17241 (N_17241,N_16853,N_16986);
or U17242 (N_17242,N_17038,N_17111);
and U17243 (N_17243,N_16813,N_17019);
and U17244 (N_17244,N_16887,N_16983);
and U17245 (N_17245,N_16994,N_16949);
nand U17246 (N_17246,N_17134,N_16979);
or U17247 (N_17247,N_16892,N_17130);
and U17248 (N_17248,N_17119,N_17140);
xnor U17249 (N_17249,N_17014,N_17155);
nor U17250 (N_17250,N_16803,N_17074);
and U17251 (N_17251,N_16862,N_16879);
nor U17252 (N_17252,N_16802,N_16923);
or U17253 (N_17253,N_17033,N_17016);
nand U17254 (N_17254,N_17052,N_17110);
nor U17255 (N_17255,N_16943,N_16839);
and U17256 (N_17256,N_17026,N_17077);
nor U17257 (N_17257,N_16857,N_17082);
xor U17258 (N_17258,N_17001,N_16865);
and U17259 (N_17259,N_17131,N_17091);
and U17260 (N_17260,N_17156,N_16895);
or U17261 (N_17261,N_17000,N_17127);
or U17262 (N_17262,N_16902,N_17171);
or U17263 (N_17263,N_17172,N_17065);
nand U17264 (N_17264,N_16951,N_16925);
nand U17265 (N_17265,N_17011,N_17138);
or U17266 (N_17266,N_16996,N_17189);
xor U17267 (N_17267,N_17042,N_16860);
or U17268 (N_17268,N_17166,N_16913);
xnor U17269 (N_17269,N_17112,N_16845);
nor U17270 (N_17270,N_17058,N_17161);
nand U17271 (N_17271,N_17063,N_17080);
nand U17272 (N_17272,N_17036,N_17098);
or U17273 (N_17273,N_17044,N_16884);
or U17274 (N_17274,N_16852,N_16922);
xor U17275 (N_17275,N_16842,N_17144);
nor U17276 (N_17276,N_17193,N_16874);
and U17277 (N_17277,N_16940,N_16972);
xnor U17278 (N_17278,N_16973,N_16832);
nor U17279 (N_17279,N_16891,N_17084);
nand U17280 (N_17280,N_16869,N_16942);
or U17281 (N_17281,N_17149,N_16929);
nor U17282 (N_17282,N_17185,N_16999);
xnor U17283 (N_17283,N_17180,N_17068);
or U17284 (N_17284,N_16956,N_16976);
or U17285 (N_17285,N_17034,N_16903);
nor U17286 (N_17286,N_17023,N_17017);
nor U17287 (N_17287,N_16821,N_16919);
xor U17288 (N_17288,N_16875,N_16864);
xor U17289 (N_17289,N_17099,N_17133);
xor U17290 (N_17290,N_17165,N_16909);
xnor U17291 (N_17291,N_16838,N_17095);
nand U17292 (N_17292,N_17039,N_16847);
nor U17293 (N_17293,N_16946,N_16984);
and U17294 (N_17294,N_16906,N_16901);
nor U17295 (N_17295,N_16991,N_16914);
nand U17296 (N_17296,N_17081,N_16945);
nand U17297 (N_17297,N_16815,N_17083);
nand U17298 (N_17298,N_17051,N_17021);
nand U17299 (N_17299,N_17106,N_17196);
xor U17300 (N_17300,N_17151,N_17108);
xnor U17301 (N_17301,N_17132,N_16800);
nand U17302 (N_17302,N_16910,N_17069);
or U17303 (N_17303,N_16954,N_16829);
nor U17304 (N_17304,N_16966,N_16975);
xor U17305 (N_17305,N_17107,N_17029);
or U17306 (N_17306,N_17086,N_16896);
or U17307 (N_17307,N_16849,N_17047);
nand U17308 (N_17308,N_17024,N_16935);
nand U17309 (N_17309,N_16810,N_17157);
xnor U17310 (N_17310,N_16893,N_16826);
nand U17311 (N_17311,N_16958,N_16866);
or U17312 (N_17312,N_16888,N_17100);
or U17313 (N_17313,N_17037,N_17175);
and U17314 (N_17314,N_17072,N_16836);
or U17315 (N_17315,N_17192,N_16953);
xnor U17316 (N_17316,N_16904,N_17003);
nand U17317 (N_17317,N_16872,N_17085);
nor U17318 (N_17318,N_16814,N_16969);
xor U17319 (N_17319,N_17109,N_16963);
nor U17320 (N_17320,N_16854,N_16939);
nor U17321 (N_17321,N_16898,N_17079);
nand U17322 (N_17322,N_17137,N_16931);
or U17323 (N_17323,N_16916,N_16830);
nand U17324 (N_17324,N_16841,N_16981);
nor U17325 (N_17325,N_17146,N_17004);
or U17326 (N_17326,N_17050,N_16878);
and U17327 (N_17327,N_17197,N_17164);
and U17328 (N_17328,N_16882,N_17057);
nor U17329 (N_17329,N_17167,N_17048);
nand U17330 (N_17330,N_16880,N_16877);
nand U17331 (N_17331,N_16897,N_16801);
or U17332 (N_17332,N_16861,N_17002);
nor U17333 (N_17333,N_17169,N_16871);
xnor U17334 (N_17334,N_17053,N_16858);
nand U17335 (N_17335,N_17078,N_17059);
nor U17336 (N_17336,N_16868,N_17188);
nor U17337 (N_17337,N_17184,N_16820);
nand U17338 (N_17338,N_16908,N_16886);
nand U17339 (N_17339,N_17183,N_17198);
and U17340 (N_17340,N_17010,N_17013);
or U17341 (N_17341,N_17199,N_17005);
nor U17342 (N_17342,N_16978,N_16944);
nor U17343 (N_17343,N_17027,N_17159);
and U17344 (N_17344,N_17046,N_17123);
nor U17345 (N_17345,N_17097,N_17096);
xor U17346 (N_17346,N_17170,N_17062);
and U17347 (N_17347,N_17008,N_17143);
nand U17348 (N_17348,N_17041,N_17066);
nand U17349 (N_17349,N_17031,N_16817);
or U17350 (N_17350,N_17177,N_17152);
or U17351 (N_17351,N_17015,N_16863);
and U17352 (N_17352,N_17182,N_17154);
and U17353 (N_17353,N_17035,N_17102);
nor U17354 (N_17354,N_16980,N_17128);
xor U17355 (N_17355,N_17093,N_17104);
and U17356 (N_17356,N_16835,N_16937);
or U17357 (N_17357,N_16936,N_17142);
xnor U17358 (N_17358,N_16982,N_16957);
or U17359 (N_17359,N_16998,N_17061);
xnor U17360 (N_17360,N_17178,N_16974);
and U17361 (N_17361,N_16912,N_16824);
nor U17362 (N_17362,N_17125,N_16932);
xor U17363 (N_17363,N_17150,N_17145);
or U17364 (N_17364,N_17040,N_16805);
nor U17365 (N_17365,N_16870,N_17054);
or U17366 (N_17366,N_16965,N_17018);
nand U17367 (N_17367,N_16822,N_17186);
and U17368 (N_17368,N_17060,N_17056);
nor U17369 (N_17369,N_17179,N_16988);
nor U17370 (N_17370,N_16846,N_16917);
xor U17371 (N_17371,N_16993,N_17126);
nor U17372 (N_17372,N_17022,N_17064);
xnor U17373 (N_17373,N_16989,N_17113);
xor U17374 (N_17374,N_17187,N_16889);
or U17375 (N_17375,N_16819,N_16990);
and U17376 (N_17376,N_17105,N_16837);
nand U17377 (N_17377,N_16921,N_16970);
xnor U17378 (N_17378,N_16997,N_16948);
nor U17379 (N_17379,N_16855,N_16900);
xnor U17380 (N_17380,N_17124,N_16952);
and U17381 (N_17381,N_17160,N_16987);
or U17382 (N_17382,N_16883,N_17025);
nand U17383 (N_17383,N_16961,N_16840);
and U17384 (N_17384,N_16812,N_17089);
nand U17385 (N_17385,N_17049,N_16844);
xor U17386 (N_17386,N_16968,N_17067);
or U17387 (N_17387,N_16959,N_17028);
xor U17388 (N_17388,N_16924,N_17190);
and U17389 (N_17389,N_16907,N_16808);
and U17390 (N_17390,N_17020,N_17055);
nor U17391 (N_17391,N_17071,N_17117);
xor U17392 (N_17392,N_16806,N_17009);
nand U17393 (N_17393,N_17115,N_16938);
nor U17394 (N_17394,N_16977,N_16859);
nand U17395 (N_17395,N_16850,N_17135);
or U17396 (N_17396,N_17141,N_16818);
nand U17397 (N_17397,N_16867,N_17073);
or U17398 (N_17398,N_16960,N_16828);
and U17399 (N_17399,N_16833,N_16834);
xor U17400 (N_17400,N_17086,N_17058);
nand U17401 (N_17401,N_17111,N_17015);
xor U17402 (N_17402,N_16882,N_17170);
and U17403 (N_17403,N_16851,N_16925);
or U17404 (N_17404,N_17194,N_16992);
nor U17405 (N_17405,N_17149,N_17019);
or U17406 (N_17406,N_16949,N_16868);
or U17407 (N_17407,N_17196,N_16837);
and U17408 (N_17408,N_17002,N_16949);
xnor U17409 (N_17409,N_16894,N_17036);
and U17410 (N_17410,N_16939,N_17172);
nor U17411 (N_17411,N_17104,N_16929);
or U17412 (N_17412,N_17187,N_17000);
or U17413 (N_17413,N_16873,N_16876);
nand U17414 (N_17414,N_16984,N_16970);
and U17415 (N_17415,N_17103,N_17086);
xor U17416 (N_17416,N_16962,N_17032);
nand U17417 (N_17417,N_17105,N_16969);
xor U17418 (N_17418,N_16899,N_17052);
xor U17419 (N_17419,N_17107,N_16804);
xnor U17420 (N_17420,N_17126,N_17059);
xnor U17421 (N_17421,N_17158,N_17004);
and U17422 (N_17422,N_17034,N_17058);
nor U17423 (N_17423,N_16859,N_16988);
nor U17424 (N_17424,N_16815,N_17112);
nor U17425 (N_17425,N_17030,N_17026);
nand U17426 (N_17426,N_16905,N_16858);
or U17427 (N_17427,N_17166,N_17025);
nor U17428 (N_17428,N_16843,N_16886);
nand U17429 (N_17429,N_17157,N_17187);
nor U17430 (N_17430,N_17195,N_17071);
nand U17431 (N_17431,N_16956,N_16821);
nor U17432 (N_17432,N_16802,N_16970);
or U17433 (N_17433,N_17128,N_17005);
and U17434 (N_17434,N_17139,N_17102);
nor U17435 (N_17435,N_16985,N_16863);
and U17436 (N_17436,N_17009,N_17037);
or U17437 (N_17437,N_17116,N_17117);
xnor U17438 (N_17438,N_16993,N_17027);
nand U17439 (N_17439,N_16837,N_16929);
or U17440 (N_17440,N_16856,N_16966);
nor U17441 (N_17441,N_16815,N_16944);
or U17442 (N_17442,N_16836,N_16989);
or U17443 (N_17443,N_17157,N_17062);
or U17444 (N_17444,N_16921,N_17000);
xnor U17445 (N_17445,N_17156,N_17179);
or U17446 (N_17446,N_16857,N_17195);
or U17447 (N_17447,N_17096,N_17100);
xnor U17448 (N_17448,N_16801,N_16982);
or U17449 (N_17449,N_17010,N_17144);
or U17450 (N_17450,N_17186,N_17059);
nand U17451 (N_17451,N_17197,N_17004);
xnor U17452 (N_17452,N_17082,N_17020);
nor U17453 (N_17453,N_16949,N_17016);
nand U17454 (N_17454,N_17125,N_17001);
nand U17455 (N_17455,N_16832,N_16829);
and U17456 (N_17456,N_17123,N_17008);
xnor U17457 (N_17457,N_16990,N_16947);
xnor U17458 (N_17458,N_16942,N_17199);
or U17459 (N_17459,N_16928,N_17077);
nor U17460 (N_17460,N_16810,N_17120);
xnor U17461 (N_17461,N_17171,N_16970);
nor U17462 (N_17462,N_17135,N_17132);
xnor U17463 (N_17463,N_16883,N_16887);
or U17464 (N_17464,N_17078,N_17124);
nand U17465 (N_17465,N_17001,N_17191);
or U17466 (N_17466,N_16909,N_16871);
or U17467 (N_17467,N_16858,N_16915);
xnor U17468 (N_17468,N_16828,N_16932);
xor U17469 (N_17469,N_16847,N_17182);
nand U17470 (N_17470,N_17148,N_16922);
or U17471 (N_17471,N_16993,N_17045);
or U17472 (N_17472,N_16860,N_17087);
nor U17473 (N_17473,N_17012,N_16843);
nor U17474 (N_17474,N_17011,N_16868);
or U17475 (N_17475,N_17023,N_16873);
nand U17476 (N_17476,N_17041,N_17199);
nand U17477 (N_17477,N_17001,N_16894);
xor U17478 (N_17478,N_16845,N_17071);
xor U17479 (N_17479,N_17037,N_17091);
nor U17480 (N_17480,N_17159,N_16844);
and U17481 (N_17481,N_16867,N_16950);
and U17482 (N_17482,N_16810,N_17164);
or U17483 (N_17483,N_17167,N_17146);
xnor U17484 (N_17484,N_16832,N_17025);
nor U17485 (N_17485,N_16942,N_17042);
nor U17486 (N_17486,N_16975,N_16995);
nand U17487 (N_17487,N_17063,N_16901);
nor U17488 (N_17488,N_16902,N_17005);
or U17489 (N_17489,N_17136,N_17121);
nor U17490 (N_17490,N_16878,N_17074);
nand U17491 (N_17491,N_17010,N_16800);
and U17492 (N_17492,N_17132,N_17083);
or U17493 (N_17493,N_16922,N_16935);
or U17494 (N_17494,N_16982,N_17064);
nand U17495 (N_17495,N_16894,N_17068);
xor U17496 (N_17496,N_16853,N_17019);
and U17497 (N_17497,N_16855,N_16882);
nand U17498 (N_17498,N_17048,N_16888);
nor U17499 (N_17499,N_16912,N_16829);
xnor U17500 (N_17500,N_16874,N_17199);
xnor U17501 (N_17501,N_16932,N_17198);
nand U17502 (N_17502,N_17095,N_16957);
nand U17503 (N_17503,N_16846,N_16922);
nor U17504 (N_17504,N_16824,N_17177);
nor U17505 (N_17505,N_17017,N_17035);
nand U17506 (N_17506,N_17051,N_17056);
and U17507 (N_17507,N_16989,N_17108);
and U17508 (N_17508,N_17175,N_16853);
nand U17509 (N_17509,N_17009,N_17007);
nand U17510 (N_17510,N_17031,N_16949);
and U17511 (N_17511,N_16956,N_17101);
xor U17512 (N_17512,N_16977,N_16913);
nand U17513 (N_17513,N_17113,N_17020);
or U17514 (N_17514,N_17051,N_16805);
nand U17515 (N_17515,N_17019,N_17123);
xor U17516 (N_17516,N_17121,N_17147);
nand U17517 (N_17517,N_17004,N_16863);
or U17518 (N_17518,N_16885,N_17072);
and U17519 (N_17519,N_17123,N_17110);
xnor U17520 (N_17520,N_17152,N_17111);
nor U17521 (N_17521,N_17096,N_17140);
and U17522 (N_17522,N_17109,N_16910);
and U17523 (N_17523,N_17028,N_16849);
xor U17524 (N_17524,N_16844,N_17149);
or U17525 (N_17525,N_17194,N_17157);
nor U17526 (N_17526,N_17098,N_16856);
nand U17527 (N_17527,N_17038,N_17108);
or U17528 (N_17528,N_16962,N_17153);
nor U17529 (N_17529,N_16964,N_16842);
or U17530 (N_17530,N_16857,N_16961);
and U17531 (N_17531,N_16810,N_17078);
nand U17532 (N_17532,N_17045,N_17102);
xor U17533 (N_17533,N_17081,N_17105);
or U17534 (N_17534,N_17145,N_16968);
and U17535 (N_17535,N_16814,N_16927);
or U17536 (N_17536,N_16851,N_17087);
or U17537 (N_17537,N_16836,N_17137);
nand U17538 (N_17538,N_17042,N_16828);
or U17539 (N_17539,N_17192,N_17141);
or U17540 (N_17540,N_17100,N_16998);
and U17541 (N_17541,N_17023,N_17046);
or U17542 (N_17542,N_17125,N_16861);
or U17543 (N_17543,N_17166,N_16802);
and U17544 (N_17544,N_16942,N_16915);
and U17545 (N_17545,N_17189,N_17076);
or U17546 (N_17546,N_16973,N_16855);
and U17547 (N_17547,N_16966,N_17163);
or U17548 (N_17548,N_16809,N_17009);
and U17549 (N_17549,N_16845,N_17161);
xor U17550 (N_17550,N_17121,N_16910);
xnor U17551 (N_17551,N_17044,N_16923);
xor U17552 (N_17552,N_17177,N_16837);
or U17553 (N_17553,N_16922,N_16897);
xor U17554 (N_17554,N_17043,N_17198);
or U17555 (N_17555,N_17140,N_16944);
nand U17556 (N_17556,N_17079,N_16993);
xor U17557 (N_17557,N_16806,N_17060);
nand U17558 (N_17558,N_16994,N_16841);
and U17559 (N_17559,N_16997,N_16833);
xor U17560 (N_17560,N_16944,N_16980);
and U17561 (N_17561,N_17185,N_16814);
and U17562 (N_17562,N_17098,N_16941);
nand U17563 (N_17563,N_16945,N_16878);
nand U17564 (N_17564,N_17093,N_17067);
nand U17565 (N_17565,N_16878,N_16844);
nor U17566 (N_17566,N_16899,N_17174);
and U17567 (N_17567,N_16878,N_16958);
nor U17568 (N_17568,N_16872,N_16956);
nor U17569 (N_17569,N_17164,N_16955);
xor U17570 (N_17570,N_17090,N_16999);
nor U17571 (N_17571,N_17073,N_17165);
and U17572 (N_17572,N_17076,N_16936);
nor U17573 (N_17573,N_16890,N_17108);
or U17574 (N_17574,N_16948,N_16961);
or U17575 (N_17575,N_17074,N_16977);
or U17576 (N_17576,N_17019,N_17114);
nor U17577 (N_17577,N_17137,N_16886);
xor U17578 (N_17578,N_16919,N_16957);
or U17579 (N_17579,N_17007,N_17072);
nand U17580 (N_17580,N_17028,N_16908);
xnor U17581 (N_17581,N_17015,N_16990);
nor U17582 (N_17582,N_17146,N_17086);
nand U17583 (N_17583,N_16957,N_16887);
nor U17584 (N_17584,N_16872,N_17144);
nor U17585 (N_17585,N_16841,N_17093);
and U17586 (N_17586,N_16930,N_16804);
nor U17587 (N_17587,N_16881,N_16933);
nand U17588 (N_17588,N_16829,N_17178);
and U17589 (N_17589,N_16964,N_16953);
xnor U17590 (N_17590,N_17064,N_17104);
or U17591 (N_17591,N_17002,N_17198);
nor U17592 (N_17592,N_17071,N_17001);
or U17593 (N_17593,N_17078,N_16890);
and U17594 (N_17594,N_16836,N_17058);
and U17595 (N_17595,N_17157,N_16990);
or U17596 (N_17596,N_16864,N_17181);
nand U17597 (N_17597,N_16955,N_17114);
nor U17598 (N_17598,N_17073,N_17111);
and U17599 (N_17599,N_16970,N_16849);
and U17600 (N_17600,N_17268,N_17544);
xnor U17601 (N_17601,N_17237,N_17321);
and U17602 (N_17602,N_17390,N_17512);
nor U17603 (N_17603,N_17259,N_17476);
nor U17604 (N_17604,N_17251,N_17352);
xnor U17605 (N_17605,N_17555,N_17309);
nand U17606 (N_17606,N_17404,N_17402);
nor U17607 (N_17607,N_17599,N_17386);
nand U17608 (N_17608,N_17380,N_17280);
nand U17609 (N_17609,N_17568,N_17382);
nand U17610 (N_17610,N_17471,N_17297);
xor U17611 (N_17611,N_17523,N_17254);
nand U17612 (N_17612,N_17407,N_17423);
and U17613 (N_17613,N_17509,N_17565);
xnor U17614 (N_17614,N_17261,N_17405);
and U17615 (N_17615,N_17572,N_17442);
nor U17616 (N_17616,N_17361,N_17594);
and U17617 (N_17617,N_17463,N_17436);
nand U17618 (N_17618,N_17569,N_17547);
nand U17619 (N_17619,N_17444,N_17369);
xor U17620 (N_17620,N_17570,N_17359);
or U17621 (N_17621,N_17536,N_17593);
and U17622 (N_17622,N_17290,N_17368);
xor U17623 (N_17623,N_17560,N_17461);
xor U17624 (N_17624,N_17454,N_17406);
or U17625 (N_17625,N_17395,N_17477);
nor U17626 (N_17626,N_17500,N_17584);
xor U17627 (N_17627,N_17396,N_17457);
xnor U17628 (N_17628,N_17527,N_17265);
nor U17629 (N_17629,N_17249,N_17333);
nand U17630 (N_17630,N_17400,N_17300);
xor U17631 (N_17631,N_17514,N_17358);
xor U17632 (N_17632,N_17578,N_17281);
xor U17633 (N_17633,N_17334,N_17401);
nand U17634 (N_17634,N_17347,N_17262);
nand U17635 (N_17635,N_17235,N_17546);
or U17636 (N_17636,N_17314,N_17526);
and U17637 (N_17637,N_17545,N_17580);
or U17638 (N_17638,N_17506,N_17273);
or U17639 (N_17639,N_17350,N_17284);
or U17640 (N_17640,N_17264,N_17575);
xor U17641 (N_17641,N_17357,N_17481);
nor U17642 (N_17642,N_17286,N_17223);
nand U17643 (N_17643,N_17226,N_17256);
and U17644 (N_17644,N_17597,N_17435);
nor U17645 (N_17645,N_17559,N_17550);
or U17646 (N_17646,N_17561,N_17231);
xor U17647 (N_17647,N_17282,N_17204);
nor U17648 (N_17648,N_17270,N_17453);
or U17649 (N_17649,N_17339,N_17344);
and U17650 (N_17650,N_17552,N_17483);
or U17651 (N_17651,N_17258,N_17474);
and U17652 (N_17652,N_17385,N_17291);
and U17653 (N_17653,N_17409,N_17447);
nor U17654 (N_17654,N_17302,N_17246);
xnor U17655 (N_17655,N_17562,N_17384);
nand U17656 (N_17656,N_17459,N_17203);
and U17657 (N_17657,N_17267,N_17322);
nand U17658 (N_17658,N_17581,N_17305);
nand U17659 (N_17659,N_17387,N_17306);
and U17660 (N_17660,N_17208,N_17535);
nand U17661 (N_17661,N_17301,N_17529);
or U17662 (N_17662,N_17220,N_17504);
nor U17663 (N_17663,N_17394,N_17591);
or U17664 (N_17664,N_17521,N_17374);
nand U17665 (N_17665,N_17553,N_17293);
xor U17666 (N_17666,N_17543,N_17383);
and U17667 (N_17667,N_17243,N_17428);
nand U17668 (N_17668,N_17224,N_17424);
and U17669 (N_17669,N_17338,N_17455);
nor U17670 (N_17670,N_17485,N_17507);
nand U17671 (N_17671,N_17554,N_17213);
or U17672 (N_17672,N_17372,N_17433);
or U17673 (N_17673,N_17397,N_17482);
xor U17674 (N_17674,N_17236,N_17266);
nor U17675 (N_17675,N_17541,N_17351);
nand U17676 (N_17676,N_17327,N_17429);
and U17677 (N_17677,N_17269,N_17532);
nand U17678 (N_17678,N_17377,N_17418);
xor U17679 (N_17679,N_17313,N_17522);
xnor U17680 (N_17680,N_17375,N_17279);
or U17681 (N_17681,N_17200,N_17449);
or U17682 (N_17682,N_17381,N_17276);
or U17683 (N_17683,N_17346,N_17440);
and U17684 (N_17684,N_17530,N_17478);
or U17685 (N_17685,N_17228,N_17229);
nor U17686 (N_17686,N_17318,N_17484);
xnor U17687 (N_17687,N_17480,N_17427);
nand U17688 (N_17688,N_17439,N_17255);
nand U17689 (N_17689,N_17430,N_17233);
xor U17690 (N_17690,N_17287,N_17263);
and U17691 (N_17691,N_17363,N_17525);
and U17692 (N_17692,N_17431,N_17516);
or U17693 (N_17693,N_17391,N_17328);
nor U17694 (N_17694,N_17212,N_17242);
or U17695 (N_17695,N_17247,N_17408);
nor U17696 (N_17696,N_17425,N_17588);
or U17697 (N_17697,N_17469,N_17336);
nor U17698 (N_17698,N_17232,N_17563);
xor U17699 (N_17699,N_17348,N_17412);
and U17700 (N_17700,N_17214,N_17250);
or U17701 (N_17701,N_17470,N_17458);
and U17702 (N_17702,N_17240,N_17537);
and U17703 (N_17703,N_17283,N_17456);
and U17704 (N_17704,N_17451,N_17316);
or U17705 (N_17705,N_17586,N_17558);
nand U17706 (N_17706,N_17495,N_17294);
xor U17707 (N_17707,N_17464,N_17360);
nor U17708 (N_17708,N_17488,N_17210);
nor U17709 (N_17709,N_17211,N_17257);
xor U17710 (N_17710,N_17364,N_17467);
or U17711 (N_17711,N_17499,N_17342);
xnor U17712 (N_17712,N_17551,N_17538);
xnor U17713 (N_17713,N_17515,N_17399);
nand U17714 (N_17714,N_17271,N_17415);
and U17715 (N_17715,N_17493,N_17362);
nor U17716 (N_17716,N_17222,N_17215);
nand U17717 (N_17717,N_17345,N_17410);
nor U17718 (N_17718,N_17592,N_17533);
nor U17719 (N_17719,N_17460,N_17331);
nor U17720 (N_17720,N_17274,N_17421);
or U17721 (N_17721,N_17420,N_17355);
nand U17722 (N_17722,N_17487,N_17413);
nand U17723 (N_17723,N_17508,N_17432);
nand U17724 (N_17724,N_17341,N_17472);
nand U17725 (N_17725,N_17491,N_17520);
nand U17726 (N_17726,N_17548,N_17379);
nor U17727 (N_17727,N_17298,N_17452);
and U17728 (N_17728,N_17244,N_17389);
nand U17729 (N_17729,N_17330,N_17517);
or U17730 (N_17730,N_17426,N_17490);
nor U17731 (N_17731,N_17557,N_17317);
nand U17732 (N_17732,N_17366,N_17496);
and U17733 (N_17733,N_17388,N_17465);
nand U17734 (N_17734,N_17307,N_17354);
xnor U17735 (N_17735,N_17511,N_17275);
nor U17736 (N_17736,N_17245,N_17227);
xor U17737 (N_17737,N_17567,N_17248);
nand U17738 (N_17738,N_17335,N_17489);
or U17739 (N_17739,N_17398,N_17462);
and U17740 (N_17740,N_17519,N_17598);
nor U17741 (N_17741,N_17540,N_17238);
nand U17742 (N_17742,N_17492,N_17542);
xnor U17743 (N_17743,N_17579,N_17445);
and U17744 (N_17744,N_17253,N_17510);
nand U17745 (N_17745,N_17443,N_17218);
nand U17746 (N_17746,N_17310,N_17272);
nand U17747 (N_17747,N_17320,N_17446);
nor U17748 (N_17748,N_17539,N_17353);
or U17749 (N_17749,N_17468,N_17308);
xor U17750 (N_17750,N_17329,N_17367);
nor U17751 (N_17751,N_17583,N_17494);
and U17752 (N_17752,N_17201,N_17531);
xnor U17753 (N_17753,N_17296,N_17577);
nor U17754 (N_17754,N_17441,N_17376);
and U17755 (N_17755,N_17349,N_17566);
or U17756 (N_17756,N_17587,N_17217);
or U17757 (N_17757,N_17356,N_17524);
nor U17758 (N_17758,N_17571,N_17595);
and U17759 (N_17759,N_17403,N_17315);
or U17760 (N_17760,N_17277,N_17325);
xor U17761 (N_17761,N_17241,N_17252);
and U17762 (N_17762,N_17304,N_17589);
nand U17763 (N_17763,N_17299,N_17371);
and U17764 (N_17764,N_17378,N_17518);
or U17765 (N_17765,N_17332,N_17392);
or U17766 (N_17766,N_17323,N_17234);
nor U17767 (N_17767,N_17528,N_17411);
xnor U17768 (N_17768,N_17202,N_17502);
nand U17769 (N_17769,N_17574,N_17260);
or U17770 (N_17770,N_17343,N_17422);
or U17771 (N_17771,N_17370,N_17582);
and U17772 (N_17772,N_17479,N_17288);
xnor U17773 (N_17773,N_17311,N_17225);
xnor U17774 (N_17774,N_17576,N_17466);
xnor U17775 (N_17775,N_17417,N_17497);
nand U17776 (N_17776,N_17205,N_17501);
and U17777 (N_17777,N_17340,N_17312);
and U17778 (N_17778,N_17437,N_17585);
nand U17779 (N_17779,N_17285,N_17207);
and U17780 (N_17780,N_17505,N_17419);
xor U17781 (N_17781,N_17230,N_17292);
xnor U17782 (N_17782,N_17473,N_17486);
and U17783 (N_17783,N_17416,N_17319);
and U17784 (N_17784,N_17373,N_17450);
and U17785 (N_17785,N_17216,N_17503);
or U17786 (N_17786,N_17448,N_17573);
nor U17787 (N_17787,N_17549,N_17303);
nand U17788 (N_17788,N_17513,N_17365);
xor U17789 (N_17789,N_17393,N_17556);
xor U17790 (N_17790,N_17337,N_17295);
and U17791 (N_17791,N_17278,N_17564);
nor U17792 (N_17792,N_17475,N_17590);
nand U17793 (N_17793,N_17239,N_17596);
xnor U17794 (N_17794,N_17534,N_17219);
and U17795 (N_17795,N_17221,N_17206);
or U17796 (N_17796,N_17438,N_17324);
xor U17797 (N_17797,N_17434,N_17209);
nor U17798 (N_17798,N_17326,N_17498);
nand U17799 (N_17799,N_17289,N_17414);
or U17800 (N_17800,N_17538,N_17309);
nand U17801 (N_17801,N_17218,N_17549);
and U17802 (N_17802,N_17383,N_17286);
nand U17803 (N_17803,N_17310,N_17515);
xor U17804 (N_17804,N_17340,N_17459);
and U17805 (N_17805,N_17212,N_17459);
nand U17806 (N_17806,N_17393,N_17508);
or U17807 (N_17807,N_17398,N_17201);
or U17808 (N_17808,N_17244,N_17423);
nand U17809 (N_17809,N_17496,N_17441);
and U17810 (N_17810,N_17271,N_17295);
nand U17811 (N_17811,N_17443,N_17382);
and U17812 (N_17812,N_17386,N_17260);
and U17813 (N_17813,N_17335,N_17435);
xnor U17814 (N_17814,N_17363,N_17546);
and U17815 (N_17815,N_17468,N_17366);
nor U17816 (N_17816,N_17285,N_17436);
or U17817 (N_17817,N_17570,N_17473);
and U17818 (N_17818,N_17257,N_17331);
nand U17819 (N_17819,N_17269,N_17207);
xor U17820 (N_17820,N_17305,N_17290);
nand U17821 (N_17821,N_17427,N_17438);
nand U17822 (N_17822,N_17431,N_17432);
and U17823 (N_17823,N_17491,N_17474);
xor U17824 (N_17824,N_17398,N_17429);
and U17825 (N_17825,N_17416,N_17492);
nand U17826 (N_17826,N_17481,N_17557);
nand U17827 (N_17827,N_17346,N_17577);
nor U17828 (N_17828,N_17396,N_17285);
nand U17829 (N_17829,N_17242,N_17556);
nand U17830 (N_17830,N_17290,N_17258);
xor U17831 (N_17831,N_17330,N_17434);
or U17832 (N_17832,N_17482,N_17539);
xor U17833 (N_17833,N_17203,N_17492);
nor U17834 (N_17834,N_17530,N_17285);
and U17835 (N_17835,N_17407,N_17321);
and U17836 (N_17836,N_17538,N_17354);
or U17837 (N_17837,N_17307,N_17564);
or U17838 (N_17838,N_17468,N_17470);
nor U17839 (N_17839,N_17526,N_17341);
xnor U17840 (N_17840,N_17493,N_17394);
nor U17841 (N_17841,N_17388,N_17504);
and U17842 (N_17842,N_17235,N_17500);
xor U17843 (N_17843,N_17493,N_17318);
xor U17844 (N_17844,N_17307,N_17340);
nor U17845 (N_17845,N_17438,N_17463);
nor U17846 (N_17846,N_17527,N_17408);
nor U17847 (N_17847,N_17270,N_17544);
nand U17848 (N_17848,N_17311,N_17256);
or U17849 (N_17849,N_17406,N_17324);
xnor U17850 (N_17850,N_17244,N_17210);
nand U17851 (N_17851,N_17339,N_17547);
and U17852 (N_17852,N_17358,N_17335);
and U17853 (N_17853,N_17570,N_17509);
or U17854 (N_17854,N_17509,N_17243);
or U17855 (N_17855,N_17505,N_17519);
or U17856 (N_17856,N_17592,N_17256);
or U17857 (N_17857,N_17548,N_17258);
nand U17858 (N_17858,N_17510,N_17370);
nand U17859 (N_17859,N_17362,N_17271);
or U17860 (N_17860,N_17445,N_17433);
nor U17861 (N_17861,N_17339,N_17533);
or U17862 (N_17862,N_17346,N_17292);
or U17863 (N_17863,N_17428,N_17399);
and U17864 (N_17864,N_17328,N_17527);
or U17865 (N_17865,N_17518,N_17413);
nand U17866 (N_17866,N_17317,N_17427);
nand U17867 (N_17867,N_17212,N_17215);
or U17868 (N_17868,N_17585,N_17415);
nand U17869 (N_17869,N_17305,N_17521);
and U17870 (N_17870,N_17235,N_17292);
xnor U17871 (N_17871,N_17438,N_17588);
and U17872 (N_17872,N_17498,N_17569);
nor U17873 (N_17873,N_17212,N_17498);
xnor U17874 (N_17874,N_17421,N_17438);
and U17875 (N_17875,N_17318,N_17221);
xor U17876 (N_17876,N_17340,N_17517);
nand U17877 (N_17877,N_17370,N_17583);
nor U17878 (N_17878,N_17524,N_17504);
nand U17879 (N_17879,N_17524,N_17208);
nand U17880 (N_17880,N_17405,N_17453);
or U17881 (N_17881,N_17231,N_17315);
or U17882 (N_17882,N_17295,N_17428);
or U17883 (N_17883,N_17572,N_17578);
nor U17884 (N_17884,N_17513,N_17352);
xor U17885 (N_17885,N_17545,N_17365);
nand U17886 (N_17886,N_17430,N_17560);
nor U17887 (N_17887,N_17434,N_17531);
nor U17888 (N_17888,N_17373,N_17353);
nand U17889 (N_17889,N_17399,N_17488);
nor U17890 (N_17890,N_17350,N_17514);
and U17891 (N_17891,N_17293,N_17462);
nand U17892 (N_17892,N_17586,N_17458);
or U17893 (N_17893,N_17215,N_17443);
and U17894 (N_17894,N_17254,N_17371);
xor U17895 (N_17895,N_17281,N_17324);
nand U17896 (N_17896,N_17254,N_17395);
nand U17897 (N_17897,N_17462,N_17285);
nor U17898 (N_17898,N_17547,N_17515);
nand U17899 (N_17899,N_17307,N_17504);
nand U17900 (N_17900,N_17301,N_17395);
nand U17901 (N_17901,N_17452,N_17273);
nor U17902 (N_17902,N_17269,N_17219);
nand U17903 (N_17903,N_17476,N_17202);
and U17904 (N_17904,N_17393,N_17343);
or U17905 (N_17905,N_17595,N_17551);
nor U17906 (N_17906,N_17533,N_17579);
or U17907 (N_17907,N_17248,N_17215);
nand U17908 (N_17908,N_17456,N_17232);
xnor U17909 (N_17909,N_17577,N_17386);
or U17910 (N_17910,N_17463,N_17407);
nand U17911 (N_17911,N_17497,N_17573);
or U17912 (N_17912,N_17293,N_17220);
or U17913 (N_17913,N_17419,N_17412);
nor U17914 (N_17914,N_17315,N_17558);
nand U17915 (N_17915,N_17272,N_17538);
xnor U17916 (N_17916,N_17529,N_17587);
and U17917 (N_17917,N_17314,N_17478);
xnor U17918 (N_17918,N_17434,N_17224);
nor U17919 (N_17919,N_17350,N_17370);
nor U17920 (N_17920,N_17202,N_17489);
and U17921 (N_17921,N_17325,N_17214);
and U17922 (N_17922,N_17348,N_17410);
xor U17923 (N_17923,N_17340,N_17306);
nor U17924 (N_17924,N_17534,N_17452);
nand U17925 (N_17925,N_17591,N_17493);
nor U17926 (N_17926,N_17384,N_17534);
nor U17927 (N_17927,N_17471,N_17285);
nor U17928 (N_17928,N_17248,N_17228);
xor U17929 (N_17929,N_17549,N_17275);
nand U17930 (N_17930,N_17218,N_17420);
xor U17931 (N_17931,N_17279,N_17264);
and U17932 (N_17932,N_17269,N_17358);
nor U17933 (N_17933,N_17502,N_17541);
nor U17934 (N_17934,N_17530,N_17552);
nor U17935 (N_17935,N_17325,N_17217);
nand U17936 (N_17936,N_17374,N_17540);
or U17937 (N_17937,N_17267,N_17466);
nor U17938 (N_17938,N_17377,N_17320);
xnor U17939 (N_17939,N_17293,N_17394);
nand U17940 (N_17940,N_17275,N_17539);
and U17941 (N_17941,N_17254,N_17351);
or U17942 (N_17942,N_17218,N_17516);
or U17943 (N_17943,N_17536,N_17583);
xnor U17944 (N_17944,N_17542,N_17459);
xor U17945 (N_17945,N_17585,N_17298);
or U17946 (N_17946,N_17340,N_17275);
and U17947 (N_17947,N_17217,N_17509);
nor U17948 (N_17948,N_17269,N_17464);
nand U17949 (N_17949,N_17201,N_17396);
and U17950 (N_17950,N_17385,N_17450);
and U17951 (N_17951,N_17346,N_17251);
nand U17952 (N_17952,N_17357,N_17525);
or U17953 (N_17953,N_17527,N_17275);
xor U17954 (N_17954,N_17508,N_17299);
nor U17955 (N_17955,N_17442,N_17201);
nand U17956 (N_17956,N_17373,N_17587);
nand U17957 (N_17957,N_17275,N_17479);
nor U17958 (N_17958,N_17575,N_17426);
nor U17959 (N_17959,N_17221,N_17509);
and U17960 (N_17960,N_17351,N_17241);
nand U17961 (N_17961,N_17519,N_17344);
nor U17962 (N_17962,N_17473,N_17399);
xnor U17963 (N_17963,N_17216,N_17228);
nand U17964 (N_17964,N_17426,N_17249);
nor U17965 (N_17965,N_17421,N_17363);
xor U17966 (N_17966,N_17292,N_17514);
or U17967 (N_17967,N_17339,N_17364);
nand U17968 (N_17968,N_17450,N_17460);
nand U17969 (N_17969,N_17364,N_17427);
nand U17970 (N_17970,N_17203,N_17490);
and U17971 (N_17971,N_17368,N_17478);
or U17972 (N_17972,N_17225,N_17470);
and U17973 (N_17973,N_17580,N_17361);
or U17974 (N_17974,N_17308,N_17340);
nor U17975 (N_17975,N_17484,N_17419);
or U17976 (N_17976,N_17453,N_17501);
or U17977 (N_17977,N_17474,N_17394);
and U17978 (N_17978,N_17438,N_17319);
xnor U17979 (N_17979,N_17557,N_17364);
nand U17980 (N_17980,N_17312,N_17438);
nand U17981 (N_17981,N_17421,N_17314);
and U17982 (N_17982,N_17486,N_17390);
and U17983 (N_17983,N_17251,N_17471);
or U17984 (N_17984,N_17305,N_17356);
and U17985 (N_17985,N_17454,N_17209);
or U17986 (N_17986,N_17377,N_17428);
and U17987 (N_17987,N_17232,N_17487);
xor U17988 (N_17988,N_17384,N_17339);
or U17989 (N_17989,N_17585,N_17248);
nand U17990 (N_17990,N_17394,N_17489);
or U17991 (N_17991,N_17599,N_17282);
nand U17992 (N_17992,N_17524,N_17329);
or U17993 (N_17993,N_17333,N_17559);
nand U17994 (N_17994,N_17416,N_17570);
and U17995 (N_17995,N_17211,N_17372);
nand U17996 (N_17996,N_17201,N_17542);
nor U17997 (N_17997,N_17257,N_17474);
nor U17998 (N_17998,N_17413,N_17211);
or U17999 (N_17999,N_17374,N_17250);
and U18000 (N_18000,N_17938,N_17909);
or U18001 (N_18001,N_17645,N_17758);
or U18002 (N_18002,N_17607,N_17854);
xor U18003 (N_18003,N_17953,N_17745);
nor U18004 (N_18004,N_17624,N_17792);
nand U18005 (N_18005,N_17799,N_17676);
nand U18006 (N_18006,N_17895,N_17871);
nand U18007 (N_18007,N_17947,N_17958);
and U18008 (N_18008,N_17765,N_17775);
xor U18009 (N_18009,N_17813,N_17702);
xor U18010 (N_18010,N_17687,N_17888);
or U18011 (N_18011,N_17935,N_17724);
xor U18012 (N_18012,N_17675,N_17707);
nand U18013 (N_18013,N_17731,N_17678);
nand U18014 (N_18014,N_17749,N_17984);
xor U18015 (N_18015,N_17954,N_17756);
nand U18016 (N_18016,N_17891,N_17714);
nand U18017 (N_18017,N_17788,N_17606);
or U18018 (N_18018,N_17898,N_17801);
or U18019 (N_18019,N_17705,N_17603);
xor U18020 (N_18020,N_17650,N_17734);
and U18021 (N_18021,N_17991,N_17785);
xnor U18022 (N_18022,N_17688,N_17715);
and U18023 (N_18023,N_17965,N_17769);
and U18024 (N_18024,N_17655,N_17861);
nand U18025 (N_18025,N_17759,N_17746);
and U18026 (N_18026,N_17826,N_17730);
and U18027 (N_18027,N_17630,N_17722);
xnor U18028 (N_18028,N_17720,N_17973);
and U18029 (N_18029,N_17865,N_17784);
nand U18030 (N_18030,N_17999,N_17776);
nor U18031 (N_18031,N_17666,N_17629);
xnor U18032 (N_18032,N_17656,N_17903);
nand U18033 (N_18033,N_17740,N_17620);
nand U18034 (N_18034,N_17889,N_17639);
nor U18035 (N_18035,N_17631,N_17995);
nor U18036 (N_18036,N_17835,N_17635);
nand U18037 (N_18037,N_17673,N_17783);
nor U18038 (N_18038,N_17950,N_17608);
xor U18039 (N_18039,N_17648,N_17793);
nand U18040 (N_18040,N_17974,N_17894);
and U18041 (N_18041,N_17866,N_17695);
nand U18042 (N_18042,N_17917,N_17971);
or U18043 (N_18043,N_17632,N_17721);
xnor U18044 (N_18044,N_17770,N_17726);
or U18045 (N_18045,N_17751,N_17841);
nor U18046 (N_18046,N_17918,N_17843);
or U18047 (N_18047,N_17627,N_17636);
nand U18048 (N_18048,N_17833,N_17653);
and U18049 (N_18049,N_17619,N_17717);
nand U18050 (N_18050,N_17680,N_17920);
nor U18051 (N_18051,N_17677,N_17628);
xnor U18052 (N_18052,N_17960,N_17962);
nand U18053 (N_18053,N_17934,N_17690);
and U18054 (N_18054,N_17940,N_17786);
nor U18055 (N_18055,N_17992,N_17760);
xor U18056 (N_18056,N_17987,N_17941);
nor U18057 (N_18057,N_17613,N_17621);
and U18058 (N_18058,N_17684,N_17864);
nand U18059 (N_18059,N_17882,N_17729);
nand U18060 (N_18060,N_17994,N_17665);
nand U18061 (N_18061,N_17808,N_17807);
and U18062 (N_18062,N_17768,N_17661);
or U18063 (N_18063,N_17689,N_17615);
or U18064 (N_18064,N_17649,N_17694);
xor U18065 (N_18065,N_17744,N_17618);
nand U18066 (N_18066,N_17872,N_17989);
and U18067 (N_18067,N_17704,N_17990);
xnor U18068 (N_18068,N_17623,N_17979);
and U18069 (N_18069,N_17912,N_17884);
and U18070 (N_18070,N_17778,N_17959);
nand U18071 (N_18071,N_17916,N_17844);
xor U18072 (N_18072,N_17794,N_17646);
and U18073 (N_18073,N_17725,N_17743);
or U18074 (N_18074,N_17975,N_17928);
nor U18075 (N_18075,N_17774,N_17824);
or U18076 (N_18076,N_17637,N_17834);
or U18077 (N_18077,N_17863,N_17955);
nand U18078 (N_18078,N_17762,N_17876);
and U18079 (N_18079,N_17795,N_17828);
xnor U18080 (N_18080,N_17658,N_17977);
and U18081 (N_18081,N_17696,N_17816);
xnor U18082 (N_18082,N_17814,N_17800);
xnor U18083 (N_18083,N_17777,N_17803);
nand U18084 (N_18084,N_17733,N_17933);
xor U18085 (N_18085,N_17670,N_17811);
nor U18086 (N_18086,N_17657,N_17612);
and U18087 (N_18087,N_17883,N_17901);
xnor U18088 (N_18088,N_17877,N_17602);
and U18089 (N_18089,N_17604,N_17647);
nand U18090 (N_18090,N_17617,N_17970);
and U18091 (N_18091,N_17963,N_17858);
or U18092 (N_18092,N_17875,N_17986);
xnor U18093 (N_18093,N_17948,N_17838);
xor U18094 (N_18094,N_17719,N_17845);
nand U18095 (N_18095,N_17949,N_17790);
xnor U18096 (N_18096,N_17741,N_17908);
and U18097 (N_18097,N_17691,N_17881);
or U18098 (N_18098,N_17739,N_17944);
nand U18099 (N_18099,N_17796,N_17832);
nor U18100 (N_18100,N_17643,N_17964);
nand U18101 (N_18101,N_17701,N_17716);
xnor U18102 (N_18102,N_17867,N_17750);
and U18103 (N_18103,N_17817,N_17685);
xor U18104 (N_18104,N_17728,N_17780);
nor U18105 (N_18105,N_17668,N_17825);
or U18106 (N_18106,N_17823,N_17836);
nand U18107 (N_18107,N_17939,N_17634);
or U18108 (N_18108,N_17980,N_17752);
and U18109 (N_18109,N_17600,N_17925);
nor U18110 (N_18110,N_17831,N_17782);
or U18111 (N_18111,N_17850,N_17761);
or U18112 (N_18112,N_17922,N_17943);
nor U18113 (N_18113,N_17764,N_17905);
xnor U18114 (N_18114,N_17654,N_17878);
nor U18115 (N_18115,N_17966,N_17609);
xnor U18116 (N_18116,N_17910,N_17930);
xor U18117 (N_18117,N_17968,N_17855);
xor U18118 (N_18118,N_17893,N_17667);
nor U18119 (N_18119,N_17806,N_17737);
nand U18120 (N_18120,N_17892,N_17913);
nand U18121 (N_18121,N_17902,N_17787);
xor U18122 (N_18122,N_17779,N_17873);
nor U18123 (N_18123,N_17622,N_17683);
or U18124 (N_18124,N_17755,N_17805);
nor U18125 (N_18125,N_17983,N_17981);
nand U18126 (N_18126,N_17932,N_17697);
or U18127 (N_18127,N_17748,N_17601);
nand U18128 (N_18128,N_17846,N_17789);
nor U18129 (N_18129,N_17710,N_17699);
and U18130 (N_18130,N_17614,N_17951);
xnor U18131 (N_18131,N_17812,N_17927);
and U18132 (N_18132,N_17616,N_17810);
nand U18133 (N_18133,N_17961,N_17633);
nand U18134 (N_18134,N_17763,N_17887);
and U18135 (N_18135,N_17742,N_17923);
nand U18136 (N_18136,N_17754,N_17839);
nor U18137 (N_18137,N_17942,N_17727);
nor U18138 (N_18138,N_17899,N_17937);
nor U18139 (N_18139,N_17662,N_17626);
nand U18140 (N_18140,N_17914,N_17840);
or U18141 (N_18141,N_17957,N_17848);
nor U18142 (N_18142,N_17732,N_17856);
or U18143 (N_18143,N_17797,N_17849);
nor U18144 (N_18144,N_17982,N_17659);
and U18145 (N_18145,N_17988,N_17985);
or U18146 (N_18146,N_17712,N_17818);
nor U18147 (N_18147,N_17993,N_17804);
nand U18148 (N_18148,N_17672,N_17641);
or U18149 (N_18149,N_17897,N_17771);
nand U18150 (N_18150,N_17868,N_17837);
and U18151 (N_18151,N_17791,N_17686);
nor U18152 (N_18152,N_17640,N_17669);
and U18153 (N_18153,N_17664,N_17952);
and U18154 (N_18154,N_17660,N_17967);
xor U18155 (N_18155,N_17880,N_17700);
nand U18156 (N_18156,N_17798,N_17651);
nor U18157 (N_18157,N_17605,N_17766);
nand U18158 (N_18158,N_17642,N_17847);
xnor U18159 (N_18159,N_17679,N_17862);
nor U18160 (N_18160,N_17842,N_17767);
xor U18161 (N_18161,N_17886,N_17900);
and U18162 (N_18162,N_17708,N_17709);
nor U18163 (N_18163,N_17674,N_17706);
xor U18164 (N_18164,N_17698,N_17921);
nor U18165 (N_18165,N_17829,N_17692);
nand U18166 (N_18166,N_17747,N_17693);
nand U18167 (N_18167,N_17852,N_17815);
or U18168 (N_18168,N_17926,N_17820);
or U18169 (N_18169,N_17652,N_17997);
xnor U18170 (N_18170,N_17915,N_17819);
or U18171 (N_18171,N_17644,N_17735);
and U18172 (N_18172,N_17772,N_17956);
xnor U18173 (N_18173,N_17802,N_17869);
nand U18174 (N_18174,N_17738,N_17753);
xnor U18175 (N_18175,N_17822,N_17830);
xor U18176 (N_18176,N_17969,N_17919);
nor U18177 (N_18177,N_17809,N_17853);
nand U18178 (N_18178,N_17929,N_17870);
or U18179 (N_18179,N_17625,N_17821);
nor U18180 (N_18180,N_17945,N_17859);
nor U18181 (N_18181,N_17904,N_17860);
xnor U18182 (N_18182,N_17610,N_17703);
or U18183 (N_18183,N_17885,N_17911);
or U18184 (N_18184,N_17757,N_17936);
nor U18185 (N_18185,N_17611,N_17671);
or U18186 (N_18186,N_17998,N_17976);
nor U18187 (N_18187,N_17851,N_17736);
or U18188 (N_18188,N_17896,N_17879);
nand U18189 (N_18189,N_17663,N_17682);
xor U18190 (N_18190,N_17978,N_17946);
nand U18191 (N_18191,N_17931,N_17827);
nor U18192 (N_18192,N_17996,N_17781);
nand U18193 (N_18193,N_17713,N_17681);
nor U18194 (N_18194,N_17924,N_17773);
nand U18195 (N_18195,N_17638,N_17711);
nand U18196 (N_18196,N_17906,N_17857);
xor U18197 (N_18197,N_17718,N_17972);
or U18198 (N_18198,N_17723,N_17890);
or U18199 (N_18199,N_17874,N_17907);
nand U18200 (N_18200,N_17677,N_17815);
and U18201 (N_18201,N_17681,N_17849);
xor U18202 (N_18202,N_17859,N_17719);
xnor U18203 (N_18203,N_17818,N_17719);
xnor U18204 (N_18204,N_17850,N_17823);
and U18205 (N_18205,N_17745,N_17940);
nand U18206 (N_18206,N_17825,N_17796);
nor U18207 (N_18207,N_17635,N_17638);
nand U18208 (N_18208,N_17956,N_17938);
and U18209 (N_18209,N_17925,N_17652);
nor U18210 (N_18210,N_17931,N_17917);
and U18211 (N_18211,N_17893,N_17642);
xor U18212 (N_18212,N_17901,N_17777);
nand U18213 (N_18213,N_17974,N_17941);
and U18214 (N_18214,N_17771,N_17964);
nor U18215 (N_18215,N_17878,N_17643);
nor U18216 (N_18216,N_17939,N_17696);
nand U18217 (N_18217,N_17685,N_17710);
or U18218 (N_18218,N_17768,N_17971);
xor U18219 (N_18219,N_17785,N_17756);
nor U18220 (N_18220,N_17833,N_17947);
xnor U18221 (N_18221,N_17709,N_17657);
and U18222 (N_18222,N_17802,N_17989);
nand U18223 (N_18223,N_17965,N_17879);
or U18224 (N_18224,N_17618,N_17890);
xnor U18225 (N_18225,N_17941,N_17944);
nor U18226 (N_18226,N_17947,N_17786);
nand U18227 (N_18227,N_17718,N_17979);
and U18228 (N_18228,N_17849,N_17757);
and U18229 (N_18229,N_17738,N_17695);
or U18230 (N_18230,N_17996,N_17691);
nand U18231 (N_18231,N_17772,N_17670);
or U18232 (N_18232,N_17886,N_17705);
or U18233 (N_18233,N_17796,N_17785);
and U18234 (N_18234,N_17875,N_17624);
or U18235 (N_18235,N_17605,N_17613);
or U18236 (N_18236,N_17671,N_17943);
nor U18237 (N_18237,N_17674,N_17688);
nor U18238 (N_18238,N_17690,N_17811);
nand U18239 (N_18239,N_17897,N_17839);
and U18240 (N_18240,N_17869,N_17841);
or U18241 (N_18241,N_17936,N_17705);
or U18242 (N_18242,N_17718,N_17757);
and U18243 (N_18243,N_17944,N_17708);
and U18244 (N_18244,N_17736,N_17965);
or U18245 (N_18245,N_17809,N_17918);
xnor U18246 (N_18246,N_17943,N_17917);
xnor U18247 (N_18247,N_17910,N_17691);
and U18248 (N_18248,N_17899,N_17605);
nand U18249 (N_18249,N_17836,N_17704);
nand U18250 (N_18250,N_17977,N_17753);
xnor U18251 (N_18251,N_17803,N_17787);
nor U18252 (N_18252,N_17941,N_17965);
nand U18253 (N_18253,N_17779,N_17657);
and U18254 (N_18254,N_17843,N_17802);
xnor U18255 (N_18255,N_17697,N_17718);
or U18256 (N_18256,N_17915,N_17880);
xnor U18257 (N_18257,N_17806,N_17880);
nand U18258 (N_18258,N_17658,N_17730);
nand U18259 (N_18259,N_17778,N_17846);
xor U18260 (N_18260,N_17804,N_17856);
nor U18261 (N_18261,N_17736,N_17659);
nand U18262 (N_18262,N_17626,N_17694);
or U18263 (N_18263,N_17875,N_17772);
nor U18264 (N_18264,N_17821,N_17762);
or U18265 (N_18265,N_17661,N_17796);
nand U18266 (N_18266,N_17602,N_17854);
and U18267 (N_18267,N_17851,N_17968);
or U18268 (N_18268,N_17763,N_17643);
and U18269 (N_18269,N_17811,N_17793);
and U18270 (N_18270,N_17876,N_17775);
and U18271 (N_18271,N_17980,N_17923);
nor U18272 (N_18272,N_17861,N_17712);
or U18273 (N_18273,N_17859,N_17989);
nor U18274 (N_18274,N_17803,N_17685);
and U18275 (N_18275,N_17798,N_17990);
nor U18276 (N_18276,N_17727,N_17959);
or U18277 (N_18277,N_17986,N_17678);
nand U18278 (N_18278,N_17697,N_17976);
and U18279 (N_18279,N_17874,N_17626);
xnor U18280 (N_18280,N_17763,N_17824);
nor U18281 (N_18281,N_17816,N_17887);
nor U18282 (N_18282,N_17770,N_17832);
and U18283 (N_18283,N_17650,N_17793);
xnor U18284 (N_18284,N_17764,N_17828);
xor U18285 (N_18285,N_17775,N_17969);
nor U18286 (N_18286,N_17727,N_17632);
nand U18287 (N_18287,N_17850,N_17867);
nand U18288 (N_18288,N_17712,N_17941);
nand U18289 (N_18289,N_17659,N_17876);
nor U18290 (N_18290,N_17887,N_17631);
or U18291 (N_18291,N_17960,N_17742);
nand U18292 (N_18292,N_17961,N_17824);
nor U18293 (N_18293,N_17680,N_17850);
and U18294 (N_18294,N_17771,N_17934);
xnor U18295 (N_18295,N_17999,N_17833);
or U18296 (N_18296,N_17600,N_17876);
nand U18297 (N_18297,N_17764,N_17936);
and U18298 (N_18298,N_17941,N_17772);
nor U18299 (N_18299,N_17821,N_17774);
nand U18300 (N_18300,N_17887,N_17836);
or U18301 (N_18301,N_17948,N_17763);
or U18302 (N_18302,N_17800,N_17606);
and U18303 (N_18303,N_17938,N_17648);
nand U18304 (N_18304,N_17908,N_17792);
and U18305 (N_18305,N_17858,N_17662);
xor U18306 (N_18306,N_17747,N_17944);
nor U18307 (N_18307,N_17801,N_17837);
nand U18308 (N_18308,N_17673,N_17625);
xnor U18309 (N_18309,N_17779,N_17841);
nor U18310 (N_18310,N_17892,N_17731);
nor U18311 (N_18311,N_17820,N_17984);
or U18312 (N_18312,N_17673,N_17780);
nor U18313 (N_18313,N_17728,N_17731);
and U18314 (N_18314,N_17635,N_17836);
or U18315 (N_18315,N_17617,N_17933);
or U18316 (N_18316,N_17725,N_17818);
and U18317 (N_18317,N_17638,N_17873);
nor U18318 (N_18318,N_17936,N_17931);
xnor U18319 (N_18319,N_17959,N_17937);
nor U18320 (N_18320,N_17697,N_17619);
or U18321 (N_18321,N_17863,N_17810);
and U18322 (N_18322,N_17813,N_17724);
xor U18323 (N_18323,N_17794,N_17811);
nor U18324 (N_18324,N_17967,N_17885);
nand U18325 (N_18325,N_17995,N_17855);
or U18326 (N_18326,N_17782,N_17995);
nor U18327 (N_18327,N_17813,N_17844);
and U18328 (N_18328,N_17772,N_17688);
nand U18329 (N_18329,N_17843,N_17998);
nand U18330 (N_18330,N_17839,N_17627);
nand U18331 (N_18331,N_17670,N_17882);
xnor U18332 (N_18332,N_17829,N_17934);
nor U18333 (N_18333,N_17863,N_17936);
nand U18334 (N_18334,N_17822,N_17952);
and U18335 (N_18335,N_17996,N_17957);
or U18336 (N_18336,N_17812,N_17670);
nand U18337 (N_18337,N_17956,N_17677);
nor U18338 (N_18338,N_17801,N_17756);
nor U18339 (N_18339,N_17780,N_17719);
nor U18340 (N_18340,N_17709,N_17744);
nor U18341 (N_18341,N_17786,N_17798);
xor U18342 (N_18342,N_17932,N_17651);
xnor U18343 (N_18343,N_17993,N_17819);
xnor U18344 (N_18344,N_17907,N_17846);
nand U18345 (N_18345,N_17744,N_17785);
and U18346 (N_18346,N_17961,N_17631);
nand U18347 (N_18347,N_17932,N_17784);
nand U18348 (N_18348,N_17911,N_17638);
nand U18349 (N_18349,N_17810,N_17675);
nor U18350 (N_18350,N_17661,N_17717);
nand U18351 (N_18351,N_17947,N_17616);
nor U18352 (N_18352,N_17673,N_17828);
xnor U18353 (N_18353,N_17698,N_17884);
nor U18354 (N_18354,N_17629,N_17851);
and U18355 (N_18355,N_17985,N_17635);
nor U18356 (N_18356,N_17746,N_17891);
nand U18357 (N_18357,N_17846,N_17934);
nand U18358 (N_18358,N_17779,N_17946);
or U18359 (N_18359,N_17792,N_17847);
nor U18360 (N_18360,N_17951,N_17770);
or U18361 (N_18361,N_17878,N_17668);
or U18362 (N_18362,N_17933,N_17659);
nand U18363 (N_18363,N_17924,N_17922);
xnor U18364 (N_18364,N_17778,N_17761);
and U18365 (N_18365,N_17724,N_17956);
nand U18366 (N_18366,N_17837,N_17926);
or U18367 (N_18367,N_17868,N_17624);
or U18368 (N_18368,N_17955,N_17986);
or U18369 (N_18369,N_17894,N_17973);
and U18370 (N_18370,N_17626,N_17774);
nand U18371 (N_18371,N_17981,N_17849);
nor U18372 (N_18372,N_17831,N_17898);
nor U18373 (N_18373,N_17632,N_17677);
or U18374 (N_18374,N_17993,N_17777);
or U18375 (N_18375,N_17692,N_17911);
xor U18376 (N_18376,N_17844,N_17704);
nand U18377 (N_18377,N_17607,N_17814);
nand U18378 (N_18378,N_17920,N_17755);
nand U18379 (N_18379,N_17882,N_17955);
and U18380 (N_18380,N_17959,N_17624);
and U18381 (N_18381,N_17803,N_17766);
and U18382 (N_18382,N_17601,N_17794);
or U18383 (N_18383,N_17909,N_17686);
and U18384 (N_18384,N_17948,N_17802);
xor U18385 (N_18385,N_17811,N_17693);
or U18386 (N_18386,N_17615,N_17663);
nor U18387 (N_18387,N_17975,N_17677);
and U18388 (N_18388,N_17767,N_17947);
nor U18389 (N_18389,N_17976,N_17876);
xor U18390 (N_18390,N_17872,N_17776);
or U18391 (N_18391,N_17782,N_17983);
nor U18392 (N_18392,N_17622,N_17636);
and U18393 (N_18393,N_17970,N_17728);
xnor U18394 (N_18394,N_17630,N_17690);
nand U18395 (N_18395,N_17907,N_17935);
xor U18396 (N_18396,N_17696,N_17690);
or U18397 (N_18397,N_17686,N_17694);
nor U18398 (N_18398,N_17693,N_17784);
or U18399 (N_18399,N_17913,N_17780);
xor U18400 (N_18400,N_18132,N_18173);
nor U18401 (N_18401,N_18210,N_18373);
xnor U18402 (N_18402,N_18184,N_18007);
and U18403 (N_18403,N_18045,N_18397);
xnor U18404 (N_18404,N_18094,N_18070);
or U18405 (N_18405,N_18042,N_18179);
and U18406 (N_18406,N_18315,N_18321);
and U18407 (N_18407,N_18174,N_18113);
and U18408 (N_18408,N_18017,N_18091);
nor U18409 (N_18409,N_18016,N_18052);
or U18410 (N_18410,N_18147,N_18381);
nor U18411 (N_18411,N_18103,N_18044);
nand U18412 (N_18412,N_18061,N_18340);
nor U18413 (N_18413,N_18213,N_18365);
and U18414 (N_18414,N_18319,N_18242);
nand U18415 (N_18415,N_18396,N_18353);
and U18416 (N_18416,N_18192,N_18398);
xor U18417 (N_18417,N_18019,N_18256);
xor U18418 (N_18418,N_18366,N_18266);
nand U18419 (N_18419,N_18342,N_18236);
nor U18420 (N_18420,N_18259,N_18162);
xnor U18421 (N_18421,N_18232,N_18293);
or U18422 (N_18422,N_18200,N_18098);
nand U18423 (N_18423,N_18193,N_18287);
xnor U18424 (N_18424,N_18394,N_18360);
xnor U18425 (N_18425,N_18382,N_18385);
or U18426 (N_18426,N_18051,N_18399);
nor U18427 (N_18427,N_18300,N_18283);
nand U18428 (N_18428,N_18130,N_18237);
or U18429 (N_18429,N_18138,N_18067);
and U18430 (N_18430,N_18069,N_18082);
nand U18431 (N_18431,N_18141,N_18218);
or U18432 (N_18432,N_18101,N_18288);
xnor U18433 (N_18433,N_18367,N_18080);
or U18434 (N_18434,N_18114,N_18296);
nand U18435 (N_18435,N_18038,N_18290);
nand U18436 (N_18436,N_18043,N_18126);
nor U18437 (N_18437,N_18209,N_18206);
and U18438 (N_18438,N_18280,N_18352);
xnor U18439 (N_18439,N_18265,N_18374);
xnor U18440 (N_18440,N_18102,N_18059);
nand U18441 (N_18441,N_18207,N_18303);
nor U18442 (N_18442,N_18109,N_18166);
and U18443 (N_18443,N_18309,N_18384);
and U18444 (N_18444,N_18369,N_18092);
nor U18445 (N_18445,N_18331,N_18351);
or U18446 (N_18446,N_18375,N_18202);
nand U18447 (N_18447,N_18362,N_18063);
xor U18448 (N_18448,N_18194,N_18023);
nand U18449 (N_18449,N_18133,N_18341);
or U18450 (N_18450,N_18175,N_18234);
nand U18451 (N_18451,N_18073,N_18364);
or U18452 (N_18452,N_18235,N_18215);
nor U18453 (N_18453,N_18329,N_18274);
xor U18454 (N_18454,N_18191,N_18081);
and U18455 (N_18455,N_18269,N_18370);
nor U18456 (N_18456,N_18318,N_18273);
or U18457 (N_18457,N_18332,N_18077);
nor U18458 (N_18458,N_18157,N_18330);
and U18459 (N_18459,N_18361,N_18222);
xor U18460 (N_18460,N_18107,N_18185);
nor U18461 (N_18461,N_18262,N_18316);
nor U18462 (N_18462,N_18379,N_18134);
xor U18463 (N_18463,N_18176,N_18271);
and U18464 (N_18464,N_18211,N_18058);
or U18465 (N_18465,N_18305,N_18110);
or U18466 (N_18466,N_18050,N_18297);
xnor U18467 (N_18467,N_18068,N_18323);
xnor U18468 (N_18468,N_18100,N_18254);
xor U18469 (N_18469,N_18251,N_18257);
and U18470 (N_18470,N_18143,N_18186);
nor U18471 (N_18471,N_18203,N_18078);
and U18472 (N_18472,N_18181,N_18326);
nor U18473 (N_18473,N_18260,N_18046);
or U18474 (N_18474,N_18199,N_18311);
and U18475 (N_18475,N_18377,N_18281);
or U18476 (N_18476,N_18093,N_18011);
xor U18477 (N_18477,N_18231,N_18088);
or U18478 (N_18478,N_18247,N_18029);
and U18479 (N_18479,N_18378,N_18244);
and U18480 (N_18480,N_18097,N_18233);
xor U18481 (N_18481,N_18112,N_18263);
nand U18482 (N_18482,N_18392,N_18118);
xnor U18483 (N_18483,N_18064,N_18386);
nor U18484 (N_18484,N_18189,N_18308);
nor U18485 (N_18485,N_18208,N_18182);
xor U18486 (N_18486,N_18284,N_18136);
or U18487 (N_18487,N_18302,N_18124);
and U18488 (N_18488,N_18368,N_18275);
nand U18489 (N_18489,N_18187,N_18227);
nor U18490 (N_18490,N_18336,N_18286);
and U18491 (N_18491,N_18252,N_18239);
and U18492 (N_18492,N_18393,N_18153);
nand U18493 (N_18493,N_18060,N_18380);
and U18494 (N_18494,N_18028,N_18055);
nor U18495 (N_18495,N_18267,N_18021);
nor U18496 (N_18496,N_18142,N_18115);
and U18497 (N_18497,N_18196,N_18178);
nand U18498 (N_18498,N_18217,N_18371);
or U18499 (N_18499,N_18125,N_18165);
xor U18500 (N_18500,N_18041,N_18131);
xnor U18501 (N_18501,N_18272,N_18146);
xor U18502 (N_18502,N_18121,N_18278);
nor U18503 (N_18503,N_18020,N_18197);
nand U18504 (N_18504,N_18348,N_18212);
xnor U18505 (N_18505,N_18156,N_18040);
nor U18506 (N_18506,N_18018,N_18317);
nand U18507 (N_18507,N_18116,N_18145);
xnor U18508 (N_18508,N_18292,N_18195);
xnor U18509 (N_18509,N_18201,N_18129);
xnor U18510 (N_18510,N_18033,N_18072);
or U18511 (N_18511,N_18356,N_18172);
xor U18512 (N_18512,N_18282,N_18246);
nor U18513 (N_18513,N_18291,N_18188);
or U18514 (N_18514,N_18035,N_18279);
or U18515 (N_18515,N_18024,N_18148);
or U18516 (N_18516,N_18390,N_18026);
nor U18517 (N_18517,N_18013,N_18095);
and U18518 (N_18518,N_18241,N_18090);
or U18519 (N_18519,N_18104,N_18128);
xnor U18520 (N_18520,N_18037,N_18000);
and U18521 (N_18521,N_18027,N_18289);
and U18522 (N_18522,N_18214,N_18048);
nor U18523 (N_18523,N_18245,N_18074);
xnor U18524 (N_18524,N_18032,N_18248);
nor U18525 (N_18525,N_18306,N_18025);
nand U18526 (N_18526,N_18036,N_18395);
nand U18527 (N_18527,N_18159,N_18139);
xor U18528 (N_18528,N_18001,N_18158);
and U18529 (N_18529,N_18312,N_18304);
or U18530 (N_18530,N_18294,N_18261);
xor U18531 (N_18531,N_18137,N_18180);
xor U18532 (N_18532,N_18062,N_18216);
and U18533 (N_18533,N_18358,N_18120);
nand U18534 (N_18534,N_18183,N_18372);
and U18535 (N_18535,N_18085,N_18150);
or U18536 (N_18536,N_18350,N_18003);
nor U18537 (N_18537,N_18354,N_18117);
or U18538 (N_18538,N_18086,N_18253);
xnor U18539 (N_18539,N_18359,N_18135);
nor U18540 (N_18540,N_18111,N_18015);
and U18541 (N_18541,N_18004,N_18299);
nand U18542 (N_18542,N_18084,N_18338);
nand U18543 (N_18543,N_18391,N_18270);
or U18544 (N_18544,N_18079,N_18066);
or U18545 (N_18545,N_18089,N_18205);
xnor U18546 (N_18546,N_18099,N_18225);
xnor U18547 (N_18547,N_18164,N_18012);
and U18548 (N_18548,N_18031,N_18339);
nand U18549 (N_18549,N_18349,N_18123);
nor U18550 (N_18550,N_18005,N_18076);
or U18551 (N_18551,N_18238,N_18152);
xor U18552 (N_18552,N_18065,N_18119);
and U18553 (N_18553,N_18295,N_18009);
nor U18554 (N_18554,N_18389,N_18334);
xnor U18555 (N_18555,N_18335,N_18388);
or U18556 (N_18556,N_18325,N_18328);
or U18557 (N_18557,N_18298,N_18387);
and U18558 (N_18558,N_18160,N_18240);
nor U18559 (N_18559,N_18149,N_18177);
or U18560 (N_18560,N_18106,N_18264);
or U18561 (N_18561,N_18301,N_18355);
nand U18562 (N_18562,N_18258,N_18320);
nor U18563 (N_18563,N_18167,N_18346);
nor U18564 (N_18564,N_18171,N_18376);
xnor U18565 (N_18565,N_18357,N_18219);
xor U18566 (N_18566,N_18002,N_18006);
nand U18567 (N_18567,N_18049,N_18198);
xnor U18568 (N_18568,N_18307,N_18345);
and U18569 (N_18569,N_18034,N_18333);
nand U18570 (N_18570,N_18056,N_18170);
xnor U18571 (N_18571,N_18285,N_18083);
and U18572 (N_18572,N_18140,N_18008);
and U18573 (N_18573,N_18268,N_18204);
nand U18574 (N_18574,N_18108,N_18276);
and U18575 (N_18575,N_18223,N_18224);
or U18576 (N_18576,N_18010,N_18226);
nor U18577 (N_18577,N_18039,N_18383);
nand U18578 (N_18578,N_18047,N_18337);
xor U18579 (N_18579,N_18169,N_18277);
and U18580 (N_18580,N_18190,N_18313);
or U18581 (N_18581,N_18087,N_18363);
nand U18582 (N_18582,N_18057,N_18220);
xnor U18583 (N_18583,N_18255,N_18163);
xnor U18584 (N_18584,N_18310,N_18053);
nor U18585 (N_18585,N_18347,N_18221);
nand U18586 (N_18586,N_18151,N_18324);
nand U18587 (N_18587,N_18343,N_18071);
and U18588 (N_18588,N_18144,N_18250);
nor U18589 (N_18589,N_18344,N_18030);
nor U18590 (N_18590,N_18105,N_18122);
and U18591 (N_18591,N_18155,N_18229);
nor U18592 (N_18592,N_18322,N_18314);
nand U18593 (N_18593,N_18243,N_18075);
and U18594 (N_18594,N_18096,N_18127);
nand U18595 (N_18595,N_18154,N_18161);
or U18596 (N_18596,N_18168,N_18022);
and U18597 (N_18597,N_18230,N_18014);
nand U18598 (N_18598,N_18054,N_18249);
or U18599 (N_18599,N_18327,N_18228);
and U18600 (N_18600,N_18199,N_18359);
or U18601 (N_18601,N_18354,N_18118);
nand U18602 (N_18602,N_18070,N_18187);
nand U18603 (N_18603,N_18257,N_18023);
and U18604 (N_18604,N_18136,N_18012);
and U18605 (N_18605,N_18367,N_18138);
nor U18606 (N_18606,N_18070,N_18202);
nand U18607 (N_18607,N_18042,N_18394);
xnor U18608 (N_18608,N_18106,N_18379);
nand U18609 (N_18609,N_18015,N_18313);
xor U18610 (N_18610,N_18368,N_18220);
or U18611 (N_18611,N_18302,N_18269);
nand U18612 (N_18612,N_18281,N_18130);
xor U18613 (N_18613,N_18308,N_18051);
and U18614 (N_18614,N_18274,N_18075);
and U18615 (N_18615,N_18269,N_18140);
nand U18616 (N_18616,N_18276,N_18265);
or U18617 (N_18617,N_18058,N_18303);
or U18618 (N_18618,N_18220,N_18226);
nor U18619 (N_18619,N_18158,N_18356);
xnor U18620 (N_18620,N_18036,N_18259);
or U18621 (N_18621,N_18023,N_18396);
nor U18622 (N_18622,N_18075,N_18110);
xor U18623 (N_18623,N_18143,N_18086);
nand U18624 (N_18624,N_18116,N_18243);
nor U18625 (N_18625,N_18036,N_18134);
and U18626 (N_18626,N_18291,N_18156);
and U18627 (N_18627,N_18078,N_18034);
and U18628 (N_18628,N_18304,N_18282);
nor U18629 (N_18629,N_18069,N_18121);
nor U18630 (N_18630,N_18146,N_18083);
or U18631 (N_18631,N_18298,N_18395);
or U18632 (N_18632,N_18095,N_18162);
xnor U18633 (N_18633,N_18289,N_18137);
and U18634 (N_18634,N_18059,N_18205);
and U18635 (N_18635,N_18076,N_18255);
xnor U18636 (N_18636,N_18299,N_18203);
nand U18637 (N_18637,N_18138,N_18072);
nor U18638 (N_18638,N_18200,N_18011);
and U18639 (N_18639,N_18230,N_18140);
or U18640 (N_18640,N_18117,N_18229);
nand U18641 (N_18641,N_18308,N_18227);
nor U18642 (N_18642,N_18067,N_18108);
xnor U18643 (N_18643,N_18133,N_18040);
nor U18644 (N_18644,N_18247,N_18113);
or U18645 (N_18645,N_18370,N_18333);
or U18646 (N_18646,N_18332,N_18106);
xor U18647 (N_18647,N_18101,N_18385);
nor U18648 (N_18648,N_18237,N_18148);
nor U18649 (N_18649,N_18088,N_18017);
or U18650 (N_18650,N_18247,N_18015);
nand U18651 (N_18651,N_18163,N_18066);
or U18652 (N_18652,N_18014,N_18192);
nand U18653 (N_18653,N_18265,N_18269);
nor U18654 (N_18654,N_18373,N_18207);
xor U18655 (N_18655,N_18127,N_18004);
xnor U18656 (N_18656,N_18102,N_18321);
or U18657 (N_18657,N_18263,N_18054);
or U18658 (N_18658,N_18086,N_18241);
nor U18659 (N_18659,N_18131,N_18336);
and U18660 (N_18660,N_18025,N_18249);
nand U18661 (N_18661,N_18094,N_18385);
xnor U18662 (N_18662,N_18007,N_18386);
nand U18663 (N_18663,N_18018,N_18238);
and U18664 (N_18664,N_18354,N_18019);
nor U18665 (N_18665,N_18311,N_18376);
nand U18666 (N_18666,N_18344,N_18192);
or U18667 (N_18667,N_18055,N_18038);
xor U18668 (N_18668,N_18222,N_18217);
or U18669 (N_18669,N_18155,N_18153);
or U18670 (N_18670,N_18237,N_18263);
and U18671 (N_18671,N_18259,N_18192);
xor U18672 (N_18672,N_18007,N_18119);
xor U18673 (N_18673,N_18299,N_18073);
and U18674 (N_18674,N_18101,N_18129);
or U18675 (N_18675,N_18339,N_18171);
or U18676 (N_18676,N_18240,N_18311);
and U18677 (N_18677,N_18177,N_18295);
and U18678 (N_18678,N_18158,N_18333);
nor U18679 (N_18679,N_18243,N_18176);
xnor U18680 (N_18680,N_18257,N_18349);
xor U18681 (N_18681,N_18016,N_18017);
nor U18682 (N_18682,N_18332,N_18307);
nor U18683 (N_18683,N_18167,N_18061);
and U18684 (N_18684,N_18313,N_18321);
xnor U18685 (N_18685,N_18201,N_18172);
and U18686 (N_18686,N_18016,N_18364);
and U18687 (N_18687,N_18017,N_18399);
or U18688 (N_18688,N_18147,N_18056);
nor U18689 (N_18689,N_18141,N_18397);
nor U18690 (N_18690,N_18200,N_18180);
nand U18691 (N_18691,N_18297,N_18166);
or U18692 (N_18692,N_18380,N_18343);
nand U18693 (N_18693,N_18223,N_18316);
or U18694 (N_18694,N_18116,N_18041);
or U18695 (N_18695,N_18349,N_18167);
nor U18696 (N_18696,N_18320,N_18149);
or U18697 (N_18697,N_18221,N_18284);
xor U18698 (N_18698,N_18090,N_18215);
and U18699 (N_18699,N_18077,N_18219);
xnor U18700 (N_18700,N_18050,N_18192);
nand U18701 (N_18701,N_18224,N_18343);
and U18702 (N_18702,N_18128,N_18281);
xor U18703 (N_18703,N_18236,N_18245);
xor U18704 (N_18704,N_18238,N_18121);
or U18705 (N_18705,N_18052,N_18062);
xnor U18706 (N_18706,N_18058,N_18069);
xnor U18707 (N_18707,N_18141,N_18318);
or U18708 (N_18708,N_18386,N_18246);
or U18709 (N_18709,N_18131,N_18155);
nor U18710 (N_18710,N_18153,N_18189);
nor U18711 (N_18711,N_18119,N_18034);
nor U18712 (N_18712,N_18136,N_18339);
nand U18713 (N_18713,N_18119,N_18262);
and U18714 (N_18714,N_18257,N_18394);
nand U18715 (N_18715,N_18394,N_18078);
and U18716 (N_18716,N_18185,N_18366);
and U18717 (N_18717,N_18123,N_18391);
xor U18718 (N_18718,N_18102,N_18132);
xnor U18719 (N_18719,N_18210,N_18189);
xor U18720 (N_18720,N_18244,N_18175);
xnor U18721 (N_18721,N_18059,N_18098);
nand U18722 (N_18722,N_18363,N_18142);
xnor U18723 (N_18723,N_18246,N_18121);
or U18724 (N_18724,N_18125,N_18031);
nand U18725 (N_18725,N_18101,N_18270);
nand U18726 (N_18726,N_18035,N_18198);
or U18727 (N_18727,N_18152,N_18037);
nor U18728 (N_18728,N_18102,N_18032);
or U18729 (N_18729,N_18284,N_18114);
xnor U18730 (N_18730,N_18274,N_18134);
nand U18731 (N_18731,N_18294,N_18080);
nor U18732 (N_18732,N_18141,N_18375);
nor U18733 (N_18733,N_18270,N_18192);
xnor U18734 (N_18734,N_18054,N_18235);
and U18735 (N_18735,N_18222,N_18038);
xor U18736 (N_18736,N_18078,N_18019);
or U18737 (N_18737,N_18385,N_18245);
and U18738 (N_18738,N_18386,N_18354);
nor U18739 (N_18739,N_18357,N_18282);
nand U18740 (N_18740,N_18237,N_18151);
nand U18741 (N_18741,N_18081,N_18189);
nor U18742 (N_18742,N_18160,N_18304);
nand U18743 (N_18743,N_18077,N_18173);
nand U18744 (N_18744,N_18003,N_18112);
xor U18745 (N_18745,N_18324,N_18203);
xor U18746 (N_18746,N_18036,N_18155);
nand U18747 (N_18747,N_18372,N_18304);
xnor U18748 (N_18748,N_18279,N_18322);
or U18749 (N_18749,N_18198,N_18216);
nand U18750 (N_18750,N_18394,N_18236);
nand U18751 (N_18751,N_18329,N_18009);
and U18752 (N_18752,N_18389,N_18397);
nand U18753 (N_18753,N_18368,N_18316);
xor U18754 (N_18754,N_18337,N_18215);
and U18755 (N_18755,N_18392,N_18329);
and U18756 (N_18756,N_18258,N_18117);
nand U18757 (N_18757,N_18384,N_18004);
and U18758 (N_18758,N_18167,N_18390);
and U18759 (N_18759,N_18024,N_18145);
xor U18760 (N_18760,N_18225,N_18271);
nand U18761 (N_18761,N_18079,N_18072);
or U18762 (N_18762,N_18330,N_18220);
or U18763 (N_18763,N_18234,N_18161);
xor U18764 (N_18764,N_18131,N_18213);
nand U18765 (N_18765,N_18289,N_18159);
nand U18766 (N_18766,N_18249,N_18152);
or U18767 (N_18767,N_18099,N_18169);
or U18768 (N_18768,N_18019,N_18337);
nand U18769 (N_18769,N_18391,N_18383);
nor U18770 (N_18770,N_18094,N_18302);
and U18771 (N_18771,N_18354,N_18204);
xnor U18772 (N_18772,N_18016,N_18373);
nand U18773 (N_18773,N_18053,N_18302);
nor U18774 (N_18774,N_18030,N_18293);
xnor U18775 (N_18775,N_18253,N_18097);
and U18776 (N_18776,N_18278,N_18050);
nor U18777 (N_18777,N_18061,N_18385);
or U18778 (N_18778,N_18365,N_18353);
or U18779 (N_18779,N_18278,N_18021);
xnor U18780 (N_18780,N_18368,N_18052);
nor U18781 (N_18781,N_18213,N_18174);
xnor U18782 (N_18782,N_18380,N_18321);
nor U18783 (N_18783,N_18050,N_18032);
nand U18784 (N_18784,N_18172,N_18076);
nand U18785 (N_18785,N_18024,N_18048);
nor U18786 (N_18786,N_18175,N_18060);
nor U18787 (N_18787,N_18180,N_18121);
nor U18788 (N_18788,N_18358,N_18179);
xor U18789 (N_18789,N_18276,N_18012);
and U18790 (N_18790,N_18085,N_18284);
xnor U18791 (N_18791,N_18130,N_18095);
nor U18792 (N_18792,N_18277,N_18224);
nor U18793 (N_18793,N_18175,N_18126);
and U18794 (N_18794,N_18215,N_18219);
nor U18795 (N_18795,N_18200,N_18066);
and U18796 (N_18796,N_18005,N_18081);
nand U18797 (N_18797,N_18394,N_18135);
nand U18798 (N_18798,N_18287,N_18243);
or U18799 (N_18799,N_18171,N_18127);
xnor U18800 (N_18800,N_18676,N_18452);
and U18801 (N_18801,N_18558,N_18471);
xnor U18802 (N_18802,N_18474,N_18571);
nor U18803 (N_18803,N_18419,N_18788);
and U18804 (N_18804,N_18654,N_18731);
and U18805 (N_18805,N_18407,N_18600);
nand U18806 (N_18806,N_18410,N_18749);
nand U18807 (N_18807,N_18429,N_18628);
nand U18808 (N_18808,N_18768,N_18551);
xnor U18809 (N_18809,N_18621,N_18648);
or U18810 (N_18810,N_18555,N_18505);
nand U18811 (N_18811,N_18739,N_18553);
or U18812 (N_18812,N_18696,N_18502);
nor U18813 (N_18813,N_18678,N_18736);
nand U18814 (N_18814,N_18478,N_18629);
and U18815 (N_18815,N_18680,N_18713);
nor U18816 (N_18816,N_18504,N_18693);
nand U18817 (N_18817,N_18528,N_18671);
nor U18818 (N_18818,N_18790,N_18742);
nor U18819 (N_18819,N_18565,N_18549);
or U18820 (N_18820,N_18639,N_18583);
xnor U18821 (N_18821,N_18616,N_18506);
nor U18822 (N_18822,N_18559,N_18759);
nor U18823 (N_18823,N_18546,N_18579);
xor U18824 (N_18824,N_18699,N_18651);
and U18825 (N_18825,N_18473,N_18743);
nand U18826 (N_18826,N_18606,N_18657);
and U18827 (N_18827,N_18487,N_18434);
xor U18828 (N_18828,N_18796,N_18760);
or U18829 (N_18829,N_18577,N_18499);
xor U18830 (N_18830,N_18735,N_18544);
and U18831 (N_18831,N_18402,N_18691);
nor U18832 (N_18832,N_18681,N_18593);
nor U18833 (N_18833,N_18780,N_18554);
or U18834 (N_18834,N_18436,N_18441);
nand U18835 (N_18835,N_18787,N_18795);
or U18836 (N_18836,N_18424,N_18647);
and U18837 (N_18837,N_18650,N_18469);
or U18838 (N_18838,N_18534,N_18516);
xnor U18839 (N_18839,N_18518,N_18725);
nor U18840 (N_18840,N_18723,N_18755);
nand U18841 (N_18841,N_18415,N_18463);
nand U18842 (N_18842,N_18674,N_18754);
and U18843 (N_18843,N_18520,N_18531);
xnor U18844 (N_18844,N_18479,N_18637);
or U18845 (N_18845,N_18669,N_18776);
nor U18846 (N_18846,N_18706,N_18617);
xnor U18847 (N_18847,N_18625,N_18602);
and U18848 (N_18848,N_18576,N_18682);
or U18849 (N_18849,N_18685,N_18451);
nor U18850 (N_18850,N_18718,N_18468);
xor U18851 (N_18851,N_18717,N_18714);
or U18852 (N_18852,N_18409,N_18622);
xnor U18853 (N_18853,N_18430,N_18751);
xor U18854 (N_18854,N_18443,N_18595);
and U18855 (N_18855,N_18707,N_18454);
nand U18856 (N_18856,N_18708,N_18514);
nor U18857 (N_18857,N_18786,N_18586);
nor U18858 (N_18858,N_18476,N_18758);
xor U18859 (N_18859,N_18422,N_18644);
nand U18860 (N_18860,N_18753,N_18513);
or U18861 (N_18861,N_18575,N_18719);
nand U18862 (N_18862,N_18635,N_18726);
xor U18863 (N_18863,N_18491,N_18605);
nand U18864 (N_18864,N_18728,N_18722);
and U18865 (N_18865,N_18445,N_18435);
and U18866 (N_18866,N_18529,N_18601);
nor U18867 (N_18867,N_18568,N_18641);
xor U18868 (N_18868,N_18604,N_18455);
nor U18869 (N_18869,N_18590,N_18427);
nor U18870 (N_18870,N_18659,N_18677);
and U18871 (N_18871,N_18495,N_18794);
nor U18872 (N_18872,N_18462,N_18715);
nor U18873 (N_18873,N_18411,N_18697);
nand U18874 (N_18874,N_18401,N_18609);
or U18875 (N_18875,N_18762,N_18489);
nor U18876 (N_18876,N_18668,N_18772);
or U18877 (N_18877,N_18431,N_18740);
nor U18878 (N_18878,N_18724,N_18587);
nand U18879 (N_18879,N_18798,N_18472);
nor U18880 (N_18880,N_18596,N_18665);
nand U18881 (N_18881,N_18423,N_18750);
and U18882 (N_18882,N_18771,N_18570);
or U18883 (N_18883,N_18783,N_18704);
nand U18884 (N_18884,N_18792,N_18515);
xnor U18885 (N_18885,N_18695,N_18716);
nor U18886 (N_18886,N_18569,N_18661);
nand U18887 (N_18887,N_18556,N_18477);
nand U18888 (N_18888,N_18510,N_18607);
nand U18889 (N_18889,N_18667,N_18573);
xnor U18890 (N_18890,N_18541,N_18797);
or U18891 (N_18891,N_18611,N_18673);
or U18892 (N_18892,N_18733,N_18413);
or U18893 (N_18893,N_18535,N_18561);
xnor U18894 (N_18894,N_18785,N_18746);
nor U18895 (N_18895,N_18433,N_18727);
nor U18896 (N_18896,N_18705,N_18597);
nand U18897 (N_18897,N_18679,N_18645);
and U18898 (N_18898,N_18627,N_18711);
nor U18899 (N_18899,N_18488,N_18757);
or U18900 (N_18900,N_18581,N_18603);
and U18901 (N_18901,N_18527,N_18480);
and U18902 (N_18902,N_18594,N_18501);
or U18903 (N_18903,N_18539,N_18598);
nor U18904 (N_18904,N_18475,N_18636);
or U18905 (N_18905,N_18664,N_18763);
nand U18906 (N_18906,N_18767,N_18779);
xnor U18907 (N_18907,N_18582,N_18523);
nor U18908 (N_18908,N_18689,N_18540);
and U18909 (N_18909,N_18522,N_18512);
xor U18910 (N_18910,N_18417,N_18624);
nor U18911 (N_18911,N_18438,N_18508);
nor U18912 (N_18912,N_18702,N_18683);
nor U18913 (N_18913,N_18420,N_18765);
and U18914 (N_18914,N_18511,N_18775);
or U18915 (N_18915,N_18756,N_18626);
or U18916 (N_18916,N_18698,N_18741);
nor U18917 (N_18917,N_18703,N_18460);
xor U18918 (N_18918,N_18619,N_18405);
or U18919 (N_18919,N_18672,N_18525);
xnor U18920 (N_18920,N_18562,N_18418);
or U18921 (N_18921,N_18729,N_18481);
nand U18922 (N_18922,N_18747,N_18543);
nand U18923 (N_18923,N_18670,N_18638);
nand U18924 (N_18924,N_18620,N_18777);
nor U18925 (N_18925,N_18764,N_18578);
xor U18926 (N_18926,N_18745,N_18737);
and U18927 (N_18927,N_18646,N_18536);
and U18928 (N_18928,N_18781,N_18591);
or U18929 (N_18929,N_18769,N_18700);
nand U18930 (N_18930,N_18485,N_18614);
or U18931 (N_18931,N_18461,N_18694);
nor U18932 (N_18932,N_18428,N_18730);
or U18933 (N_18933,N_18631,N_18721);
and U18934 (N_18934,N_18437,N_18766);
nor U18935 (N_18935,N_18537,N_18521);
nand U18936 (N_18936,N_18509,N_18439);
or U18937 (N_18937,N_18748,N_18450);
or U18938 (N_18938,N_18563,N_18545);
nor U18939 (N_18939,N_18592,N_18432);
or U18940 (N_18940,N_18675,N_18538);
nor U18941 (N_18941,N_18684,N_18406);
nand U18942 (N_18942,N_18449,N_18530);
xor U18943 (N_18943,N_18687,N_18421);
and U18944 (N_18944,N_18533,N_18503);
nand U18945 (N_18945,N_18613,N_18612);
or U18946 (N_18946,N_18574,N_18466);
nor U18947 (N_18947,N_18492,N_18440);
xor U18948 (N_18948,N_18793,N_18519);
nand U18949 (N_18949,N_18608,N_18453);
or U18950 (N_18950,N_18566,N_18632);
xor U18951 (N_18951,N_18400,N_18630);
or U18952 (N_18952,N_18560,N_18618);
or U18953 (N_18953,N_18653,N_18799);
nand U18954 (N_18954,N_18580,N_18738);
nor U18955 (N_18955,N_18649,N_18784);
xnor U18956 (N_18956,N_18442,N_18734);
or U18957 (N_18957,N_18589,N_18493);
and U18958 (N_18958,N_18557,N_18752);
nor U18959 (N_18959,N_18643,N_18652);
nor U18960 (N_18960,N_18791,N_18599);
xor U18961 (N_18961,N_18459,N_18774);
and U18962 (N_18962,N_18465,N_18494);
or U18963 (N_18963,N_18482,N_18709);
nor U18964 (N_18964,N_18623,N_18500);
and U18965 (N_18965,N_18416,N_18688);
and U18966 (N_18966,N_18660,N_18634);
xnor U18967 (N_18967,N_18444,N_18662);
nor U18968 (N_18968,N_18712,N_18701);
xnor U18969 (N_18969,N_18610,N_18532);
nor U18970 (N_18970,N_18426,N_18486);
xnor U18971 (N_18971,N_18484,N_18483);
and U18972 (N_18972,N_18567,N_18448);
nand U18973 (N_18973,N_18496,N_18447);
nand U18974 (N_18974,N_18770,N_18456);
nor U18975 (N_18975,N_18732,N_18666);
and U18976 (N_18976,N_18548,N_18403);
nand U18977 (N_18977,N_18564,N_18458);
and U18978 (N_18978,N_18425,N_18552);
and U18979 (N_18979,N_18773,N_18761);
xor U18980 (N_18980,N_18585,N_18692);
and U18981 (N_18981,N_18550,N_18467);
or U18982 (N_18982,N_18457,N_18517);
nand U18983 (N_18983,N_18720,N_18526);
and U18984 (N_18984,N_18408,N_18663);
nand U18985 (N_18985,N_18497,N_18640);
and U18986 (N_18986,N_18464,N_18656);
xor U18987 (N_18987,N_18524,N_18778);
nand U18988 (N_18988,N_18412,N_18414);
xnor U18989 (N_18989,N_18507,N_18498);
or U18990 (N_18990,N_18572,N_18404);
xor U18991 (N_18991,N_18686,N_18633);
nor U18992 (N_18992,N_18584,N_18588);
xor U18993 (N_18993,N_18615,N_18658);
or U18994 (N_18994,N_18446,N_18547);
or U18995 (N_18995,N_18782,N_18642);
xnor U18996 (N_18996,N_18470,N_18690);
and U18997 (N_18997,N_18655,N_18710);
nand U18998 (N_18998,N_18542,N_18744);
nand U18999 (N_18999,N_18789,N_18490);
and U19000 (N_19000,N_18787,N_18446);
xnor U19001 (N_19001,N_18748,N_18444);
and U19002 (N_19002,N_18535,N_18719);
nand U19003 (N_19003,N_18400,N_18591);
xor U19004 (N_19004,N_18714,N_18504);
xnor U19005 (N_19005,N_18447,N_18758);
xor U19006 (N_19006,N_18628,N_18658);
nor U19007 (N_19007,N_18457,N_18786);
xor U19008 (N_19008,N_18571,N_18640);
nor U19009 (N_19009,N_18635,N_18776);
xnor U19010 (N_19010,N_18609,N_18417);
xor U19011 (N_19011,N_18508,N_18709);
nand U19012 (N_19012,N_18625,N_18617);
nand U19013 (N_19013,N_18670,N_18464);
nor U19014 (N_19014,N_18625,N_18587);
or U19015 (N_19015,N_18550,N_18526);
xor U19016 (N_19016,N_18433,N_18462);
xnor U19017 (N_19017,N_18560,N_18473);
xor U19018 (N_19018,N_18567,N_18605);
nand U19019 (N_19019,N_18732,N_18482);
xnor U19020 (N_19020,N_18748,N_18696);
or U19021 (N_19021,N_18636,N_18614);
nand U19022 (N_19022,N_18422,N_18734);
nand U19023 (N_19023,N_18411,N_18628);
nor U19024 (N_19024,N_18452,N_18510);
and U19025 (N_19025,N_18663,N_18737);
nor U19026 (N_19026,N_18610,N_18706);
nor U19027 (N_19027,N_18462,N_18689);
nand U19028 (N_19028,N_18623,N_18734);
xor U19029 (N_19029,N_18495,N_18436);
xor U19030 (N_19030,N_18752,N_18496);
and U19031 (N_19031,N_18575,N_18469);
or U19032 (N_19032,N_18464,N_18570);
and U19033 (N_19033,N_18760,N_18564);
nor U19034 (N_19034,N_18469,N_18731);
xor U19035 (N_19035,N_18634,N_18468);
nand U19036 (N_19036,N_18711,N_18471);
nor U19037 (N_19037,N_18400,N_18695);
nand U19038 (N_19038,N_18484,N_18497);
and U19039 (N_19039,N_18658,N_18694);
or U19040 (N_19040,N_18542,N_18620);
nor U19041 (N_19041,N_18460,N_18475);
xnor U19042 (N_19042,N_18536,N_18592);
or U19043 (N_19043,N_18437,N_18716);
xnor U19044 (N_19044,N_18665,N_18650);
nor U19045 (N_19045,N_18595,N_18663);
nand U19046 (N_19046,N_18568,N_18410);
nor U19047 (N_19047,N_18704,N_18575);
xnor U19048 (N_19048,N_18576,N_18772);
nor U19049 (N_19049,N_18798,N_18562);
nand U19050 (N_19050,N_18451,N_18443);
nand U19051 (N_19051,N_18708,N_18417);
and U19052 (N_19052,N_18627,N_18794);
xnor U19053 (N_19053,N_18454,N_18461);
xnor U19054 (N_19054,N_18647,N_18670);
or U19055 (N_19055,N_18734,N_18676);
xor U19056 (N_19056,N_18405,N_18589);
and U19057 (N_19057,N_18454,N_18629);
nand U19058 (N_19058,N_18624,N_18666);
nand U19059 (N_19059,N_18759,N_18710);
nor U19060 (N_19060,N_18479,N_18711);
or U19061 (N_19061,N_18699,N_18649);
xnor U19062 (N_19062,N_18452,N_18569);
or U19063 (N_19063,N_18704,N_18619);
xor U19064 (N_19064,N_18761,N_18413);
nand U19065 (N_19065,N_18588,N_18605);
nand U19066 (N_19066,N_18593,N_18620);
or U19067 (N_19067,N_18582,N_18756);
nand U19068 (N_19068,N_18502,N_18660);
or U19069 (N_19069,N_18767,N_18621);
nand U19070 (N_19070,N_18504,N_18559);
and U19071 (N_19071,N_18613,N_18718);
nor U19072 (N_19072,N_18618,N_18719);
nor U19073 (N_19073,N_18559,N_18449);
or U19074 (N_19074,N_18657,N_18563);
nand U19075 (N_19075,N_18436,N_18427);
or U19076 (N_19076,N_18744,N_18705);
or U19077 (N_19077,N_18455,N_18556);
and U19078 (N_19078,N_18405,N_18511);
xnor U19079 (N_19079,N_18454,N_18686);
or U19080 (N_19080,N_18435,N_18523);
nand U19081 (N_19081,N_18587,N_18679);
or U19082 (N_19082,N_18700,N_18521);
nand U19083 (N_19083,N_18789,N_18502);
nor U19084 (N_19084,N_18743,N_18699);
and U19085 (N_19085,N_18718,N_18768);
or U19086 (N_19086,N_18666,N_18526);
xor U19087 (N_19087,N_18474,N_18725);
nor U19088 (N_19088,N_18404,N_18405);
xor U19089 (N_19089,N_18690,N_18538);
nor U19090 (N_19090,N_18704,N_18555);
nand U19091 (N_19091,N_18751,N_18776);
or U19092 (N_19092,N_18693,N_18556);
xnor U19093 (N_19093,N_18415,N_18498);
or U19094 (N_19094,N_18685,N_18712);
nor U19095 (N_19095,N_18765,N_18497);
nand U19096 (N_19096,N_18700,N_18788);
xnor U19097 (N_19097,N_18772,N_18740);
nor U19098 (N_19098,N_18633,N_18703);
and U19099 (N_19099,N_18429,N_18695);
and U19100 (N_19100,N_18771,N_18408);
and U19101 (N_19101,N_18736,N_18471);
and U19102 (N_19102,N_18527,N_18660);
and U19103 (N_19103,N_18660,N_18632);
xnor U19104 (N_19104,N_18782,N_18407);
xor U19105 (N_19105,N_18792,N_18544);
xnor U19106 (N_19106,N_18559,N_18684);
or U19107 (N_19107,N_18799,N_18684);
nor U19108 (N_19108,N_18580,N_18756);
nand U19109 (N_19109,N_18470,N_18656);
nand U19110 (N_19110,N_18749,N_18518);
or U19111 (N_19111,N_18677,N_18490);
xor U19112 (N_19112,N_18759,N_18596);
nand U19113 (N_19113,N_18609,N_18793);
nor U19114 (N_19114,N_18763,N_18461);
xnor U19115 (N_19115,N_18725,N_18554);
nor U19116 (N_19116,N_18404,N_18760);
xnor U19117 (N_19117,N_18408,N_18425);
and U19118 (N_19118,N_18528,N_18653);
or U19119 (N_19119,N_18657,N_18498);
xnor U19120 (N_19120,N_18774,N_18749);
nand U19121 (N_19121,N_18494,N_18431);
nor U19122 (N_19122,N_18777,N_18442);
or U19123 (N_19123,N_18546,N_18656);
or U19124 (N_19124,N_18455,N_18679);
nand U19125 (N_19125,N_18550,N_18560);
nor U19126 (N_19126,N_18510,N_18716);
nor U19127 (N_19127,N_18411,N_18516);
xnor U19128 (N_19128,N_18749,N_18506);
and U19129 (N_19129,N_18611,N_18754);
and U19130 (N_19130,N_18512,N_18590);
xnor U19131 (N_19131,N_18746,N_18742);
and U19132 (N_19132,N_18543,N_18426);
nand U19133 (N_19133,N_18485,N_18665);
nor U19134 (N_19134,N_18723,N_18504);
nand U19135 (N_19135,N_18767,N_18492);
or U19136 (N_19136,N_18711,N_18556);
nor U19137 (N_19137,N_18432,N_18442);
nand U19138 (N_19138,N_18751,N_18610);
nand U19139 (N_19139,N_18733,N_18680);
and U19140 (N_19140,N_18528,N_18743);
nor U19141 (N_19141,N_18589,N_18447);
xor U19142 (N_19142,N_18778,N_18717);
and U19143 (N_19143,N_18735,N_18725);
and U19144 (N_19144,N_18446,N_18496);
nand U19145 (N_19145,N_18589,N_18776);
xnor U19146 (N_19146,N_18421,N_18492);
and U19147 (N_19147,N_18533,N_18747);
or U19148 (N_19148,N_18495,N_18760);
or U19149 (N_19149,N_18526,N_18479);
nand U19150 (N_19150,N_18447,N_18666);
nor U19151 (N_19151,N_18469,N_18714);
or U19152 (N_19152,N_18516,N_18623);
nor U19153 (N_19153,N_18493,N_18573);
and U19154 (N_19154,N_18505,N_18459);
or U19155 (N_19155,N_18610,N_18663);
xnor U19156 (N_19156,N_18605,N_18541);
xor U19157 (N_19157,N_18453,N_18754);
nand U19158 (N_19158,N_18488,N_18529);
or U19159 (N_19159,N_18608,N_18546);
nand U19160 (N_19160,N_18578,N_18439);
nor U19161 (N_19161,N_18553,N_18507);
and U19162 (N_19162,N_18729,N_18529);
and U19163 (N_19163,N_18616,N_18795);
nor U19164 (N_19164,N_18557,N_18622);
and U19165 (N_19165,N_18673,N_18782);
nand U19166 (N_19166,N_18617,N_18585);
and U19167 (N_19167,N_18425,N_18529);
nor U19168 (N_19168,N_18604,N_18759);
xor U19169 (N_19169,N_18490,N_18661);
or U19170 (N_19170,N_18478,N_18595);
xnor U19171 (N_19171,N_18659,N_18586);
xor U19172 (N_19172,N_18535,N_18773);
nand U19173 (N_19173,N_18783,N_18520);
nand U19174 (N_19174,N_18460,N_18797);
or U19175 (N_19175,N_18544,N_18601);
xor U19176 (N_19176,N_18767,N_18450);
and U19177 (N_19177,N_18759,N_18574);
or U19178 (N_19178,N_18540,N_18433);
or U19179 (N_19179,N_18772,N_18593);
or U19180 (N_19180,N_18499,N_18771);
and U19181 (N_19181,N_18435,N_18687);
or U19182 (N_19182,N_18569,N_18451);
or U19183 (N_19183,N_18424,N_18725);
nor U19184 (N_19184,N_18563,N_18625);
and U19185 (N_19185,N_18484,N_18664);
xor U19186 (N_19186,N_18508,N_18417);
xor U19187 (N_19187,N_18799,N_18579);
and U19188 (N_19188,N_18428,N_18786);
xnor U19189 (N_19189,N_18638,N_18562);
or U19190 (N_19190,N_18705,N_18688);
nor U19191 (N_19191,N_18611,N_18563);
nor U19192 (N_19192,N_18704,N_18732);
nand U19193 (N_19193,N_18783,N_18718);
nand U19194 (N_19194,N_18655,N_18402);
nor U19195 (N_19195,N_18746,N_18612);
and U19196 (N_19196,N_18539,N_18739);
xor U19197 (N_19197,N_18406,N_18607);
and U19198 (N_19198,N_18684,N_18439);
nand U19199 (N_19199,N_18629,N_18679);
or U19200 (N_19200,N_18968,N_18959);
or U19201 (N_19201,N_18976,N_18996);
or U19202 (N_19202,N_19041,N_18994);
xnor U19203 (N_19203,N_18887,N_18836);
xor U19204 (N_19204,N_19155,N_18950);
xnor U19205 (N_19205,N_19007,N_18980);
nand U19206 (N_19206,N_18992,N_18974);
and U19207 (N_19207,N_18859,N_19073);
or U19208 (N_19208,N_18800,N_18873);
xor U19209 (N_19209,N_19069,N_18977);
nand U19210 (N_19210,N_18872,N_18855);
xor U19211 (N_19211,N_19181,N_19004);
nor U19212 (N_19212,N_19123,N_19122);
nand U19213 (N_19213,N_18809,N_18816);
nand U19214 (N_19214,N_19028,N_18991);
or U19215 (N_19215,N_18814,N_19154);
xor U19216 (N_19216,N_19054,N_18903);
nor U19217 (N_19217,N_19182,N_18849);
and U19218 (N_19218,N_19140,N_18829);
or U19219 (N_19219,N_18900,N_18811);
nor U19220 (N_19220,N_18971,N_18961);
or U19221 (N_19221,N_18823,N_18820);
and U19222 (N_19222,N_18978,N_19190);
xor U19223 (N_19223,N_19177,N_19021);
and U19224 (N_19224,N_18913,N_19098);
and U19225 (N_19225,N_19114,N_19086);
nor U19226 (N_19226,N_18840,N_18926);
nand U19227 (N_19227,N_18963,N_18924);
xnor U19228 (N_19228,N_19164,N_19188);
or U19229 (N_19229,N_19023,N_18826);
and U19230 (N_19230,N_18979,N_18885);
or U19231 (N_19231,N_19011,N_18888);
or U19232 (N_19232,N_18934,N_19075);
or U19233 (N_19233,N_18905,N_19172);
nand U19234 (N_19234,N_19166,N_19153);
xor U19235 (N_19235,N_19091,N_19199);
or U19236 (N_19236,N_19040,N_19070);
or U19237 (N_19237,N_18834,N_19010);
xnor U19238 (N_19238,N_18975,N_19189);
nand U19239 (N_19239,N_19051,N_18807);
xor U19240 (N_19240,N_19198,N_18901);
nand U19241 (N_19241,N_19101,N_18935);
and U19242 (N_19242,N_18912,N_18880);
nand U19243 (N_19243,N_18874,N_18870);
and U19244 (N_19244,N_19145,N_19178);
xnor U19245 (N_19245,N_19163,N_18856);
xnor U19246 (N_19246,N_19100,N_18825);
and U19247 (N_19247,N_19032,N_18947);
nand U19248 (N_19248,N_18998,N_18857);
nand U19249 (N_19249,N_19144,N_19055);
nor U19250 (N_19250,N_19033,N_18933);
or U19251 (N_19251,N_18920,N_18884);
or U19252 (N_19252,N_18893,N_19194);
and U19253 (N_19253,N_18862,N_19096);
nor U19254 (N_19254,N_18940,N_19106);
or U19255 (N_19255,N_19186,N_18848);
nor U19256 (N_19256,N_19120,N_18812);
nor U19257 (N_19257,N_19111,N_19082);
and U19258 (N_19258,N_18941,N_18931);
nor U19259 (N_19259,N_19005,N_19142);
nand U19260 (N_19260,N_19135,N_18995);
or U19261 (N_19261,N_19170,N_19036);
nor U19262 (N_19262,N_18803,N_18891);
or U19263 (N_19263,N_18984,N_19148);
and U19264 (N_19264,N_18846,N_18938);
nor U19265 (N_19265,N_19080,N_19035);
nor U19266 (N_19266,N_19057,N_18943);
nor U19267 (N_19267,N_19015,N_19087);
and U19268 (N_19268,N_19146,N_18879);
and U19269 (N_19269,N_19008,N_19104);
nor U19270 (N_19270,N_18886,N_18923);
nor U19271 (N_19271,N_18889,N_19195);
or U19272 (N_19272,N_19134,N_19088);
or U19273 (N_19273,N_18904,N_19058);
or U19274 (N_19274,N_19171,N_19084);
nand U19275 (N_19275,N_19071,N_19185);
xor U19276 (N_19276,N_18817,N_18921);
xor U19277 (N_19277,N_18983,N_19151);
nand U19278 (N_19278,N_19090,N_19184);
or U19279 (N_19279,N_18850,N_19117);
nand U19280 (N_19280,N_18827,N_19093);
nor U19281 (N_19281,N_18922,N_19168);
nand U19282 (N_19282,N_18973,N_18802);
or U19283 (N_19283,N_18982,N_18909);
or U19284 (N_19284,N_19063,N_19147);
nand U19285 (N_19285,N_18867,N_18815);
nor U19286 (N_19286,N_19115,N_18910);
nor U19287 (N_19287,N_19026,N_18833);
nor U19288 (N_19288,N_18896,N_19017);
xor U19289 (N_19289,N_19183,N_18837);
nand U19290 (N_19290,N_19012,N_19074);
or U19291 (N_19291,N_19043,N_19160);
nand U19292 (N_19292,N_19022,N_18878);
nand U19293 (N_19293,N_19137,N_18871);
nor U19294 (N_19294,N_18967,N_18892);
or U19295 (N_19295,N_18860,N_19150);
and U19296 (N_19296,N_19009,N_19077);
xor U19297 (N_19297,N_19130,N_18813);
nand U19298 (N_19298,N_19131,N_19020);
and U19299 (N_19299,N_18927,N_18832);
xor U19300 (N_19300,N_18839,N_19099);
nand U19301 (N_19301,N_18960,N_18942);
or U19302 (N_19302,N_18883,N_18853);
xnor U19303 (N_19303,N_18985,N_19060);
xor U19304 (N_19304,N_19105,N_18894);
and U19305 (N_19305,N_19103,N_18919);
xnor U19306 (N_19306,N_19068,N_19013);
or U19307 (N_19307,N_19129,N_19102);
nand U19308 (N_19308,N_19125,N_18951);
xnor U19309 (N_19309,N_19174,N_19045);
and U19310 (N_19310,N_19061,N_18822);
or U19311 (N_19311,N_18851,N_18954);
nor U19312 (N_19312,N_19175,N_19113);
xor U19313 (N_19313,N_18882,N_19108);
nor U19314 (N_19314,N_19167,N_19132);
and U19315 (N_19315,N_19001,N_18944);
nor U19316 (N_19316,N_18830,N_19094);
xor U19317 (N_19317,N_19107,N_19046);
nand U19318 (N_19318,N_19024,N_18930);
nor U19319 (N_19319,N_19152,N_18847);
or U19320 (N_19320,N_19027,N_18808);
nand U19321 (N_19321,N_18801,N_19124);
nor U19322 (N_19322,N_18906,N_19158);
and U19323 (N_19323,N_18895,N_19079);
nor U19324 (N_19324,N_18866,N_19149);
xnor U19325 (N_19325,N_19048,N_18841);
nand U19326 (N_19326,N_19014,N_19029);
nor U19327 (N_19327,N_18831,N_18928);
or U19328 (N_19328,N_19109,N_19089);
and U19329 (N_19329,N_18865,N_19197);
nor U19330 (N_19330,N_19176,N_19025);
or U19331 (N_19331,N_18902,N_18881);
nor U19332 (N_19332,N_18890,N_19083);
and U19333 (N_19333,N_19118,N_19031);
or U19334 (N_19334,N_18949,N_19138);
or U19335 (N_19335,N_19116,N_19157);
and U19336 (N_19336,N_18806,N_18988);
nor U19337 (N_19337,N_19092,N_19064);
and U19338 (N_19338,N_19065,N_18969);
and U19339 (N_19339,N_18845,N_18824);
or U19340 (N_19340,N_19030,N_18970);
or U19341 (N_19341,N_19059,N_19072);
xor U19342 (N_19342,N_18908,N_19136);
xnor U19343 (N_19343,N_18986,N_19085);
xnor U19344 (N_19344,N_19042,N_18805);
nor U19345 (N_19345,N_18804,N_19127);
nand U19346 (N_19346,N_19034,N_18861);
and U19347 (N_19347,N_18907,N_19126);
nand U19348 (N_19348,N_19067,N_19056);
or U19349 (N_19349,N_18993,N_18911);
xnor U19350 (N_19350,N_19097,N_18828);
and U19351 (N_19351,N_19196,N_19156);
nand U19352 (N_19352,N_18946,N_19192);
xnor U19353 (N_19353,N_19191,N_19037);
xor U19354 (N_19354,N_18835,N_18843);
xnor U19355 (N_19355,N_18864,N_18869);
xnor U19356 (N_19356,N_18948,N_18972);
or U19357 (N_19357,N_19016,N_18877);
nor U19358 (N_19358,N_19180,N_19052);
nand U19359 (N_19359,N_18964,N_18981);
or U19360 (N_19360,N_18918,N_19169);
and U19361 (N_19361,N_19112,N_18987);
nor U19362 (N_19362,N_18962,N_19081);
nor U19363 (N_19363,N_18875,N_18925);
nand U19364 (N_19364,N_19002,N_19050);
nand U19365 (N_19365,N_19128,N_19187);
or U19366 (N_19366,N_19165,N_19110);
and U19367 (N_19367,N_19018,N_19139);
or U19368 (N_19368,N_18952,N_18936);
nor U19369 (N_19369,N_18965,N_19076);
or U19370 (N_19370,N_18955,N_19078);
xnor U19371 (N_19371,N_19039,N_18915);
and U19372 (N_19372,N_18821,N_18957);
and U19373 (N_19373,N_19161,N_19044);
nor U19374 (N_19374,N_18990,N_18844);
or U19375 (N_19375,N_19062,N_18818);
xor U19376 (N_19376,N_18897,N_19159);
and U19377 (N_19377,N_18854,N_19141);
nand U19378 (N_19378,N_18989,N_19193);
nand U19379 (N_19379,N_18917,N_18916);
xnor U19380 (N_19380,N_19049,N_19053);
and U19381 (N_19381,N_18858,N_18868);
nand U19382 (N_19382,N_19038,N_18953);
and U19383 (N_19383,N_19162,N_19173);
and U19384 (N_19384,N_19066,N_19179);
and U19385 (N_19385,N_18876,N_18945);
and U19386 (N_19386,N_19006,N_18810);
xor U19387 (N_19387,N_18863,N_18842);
xor U19388 (N_19388,N_19121,N_18956);
xnor U19389 (N_19389,N_18937,N_19119);
nand U19390 (N_19390,N_18898,N_18999);
and U19391 (N_19391,N_19095,N_19003);
nand U19392 (N_19392,N_18929,N_18914);
xor U19393 (N_19393,N_18966,N_18819);
xor U19394 (N_19394,N_19143,N_19047);
nand U19395 (N_19395,N_19000,N_18939);
or U19396 (N_19396,N_19133,N_18932);
nand U19397 (N_19397,N_18899,N_18838);
or U19398 (N_19398,N_18958,N_18852);
and U19399 (N_19399,N_19019,N_18997);
nor U19400 (N_19400,N_19101,N_19173);
and U19401 (N_19401,N_18941,N_19189);
and U19402 (N_19402,N_18897,N_18991);
nor U19403 (N_19403,N_19058,N_18903);
and U19404 (N_19404,N_19023,N_18845);
nand U19405 (N_19405,N_19088,N_18905);
or U19406 (N_19406,N_19114,N_19154);
nand U19407 (N_19407,N_18826,N_18861);
xnor U19408 (N_19408,N_19158,N_19090);
and U19409 (N_19409,N_19000,N_18906);
xor U19410 (N_19410,N_18943,N_19166);
or U19411 (N_19411,N_18887,N_19031);
nand U19412 (N_19412,N_18886,N_19050);
or U19413 (N_19413,N_19065,N_18973);
nor U19414 (N_19414,N_19157,N_19114);
nor U19415 (N_19415,N_19110,N_19070);
and U19416 (N_19416,N_19013,N_18921);
or U19417 (N_19417,N_19012,N_19177);
nor U19418 (N_19418,N_19159,N_18840);
nand U19419 (N_19419,N_19090,N_19087);
or U19420 (N_19420,N_19049,N_19021);
nand U19421 (N_19421,N_18808,N_18890);
and U19422 (N_19422,N_18881,N_19066);
and U19423 (N_19423,N_18809,N_18897);
and U19424 (N_19424,N_19078,N_19053);
xor U19425 (N_19425,N_19044,N_19068);
or U19426 (N_19426,N_19165,N_18879);
or U19427 (N_19427,N_19102,N_18862);
xor U19428 (N_19428,N_19160,N_18917);
nand U19429 (N_19429,N_19046,N_18993);
and U19430 (N_19430,N_18944,N_18867);
or U19431 (N_19431,N_19145,N_19049);
or U19432 (N_19432,N_19189,N_18959);
xor U19433 (N_19433,N_18972,N_19169);
nor U19434 (N_19434,N_19162,N_18825);
xor U19435 (N_19435,N_18980,N_19151);
xnor U19436 (N_19436,N_18903,N_19057);
nor U19437 (N_19437,N_19197,N_19100);
or U19438 (N_19438,N_18815,N_19177);
and U19439 (N_19439,N_19093,N_19019);
and U19440 (N_19440,N_18833,N_18857);
or U19441 (N_19441,N_18944,N_19157);
or U19442 (N_19442,N_19151,N_18855);
xnor U19443 (N_19443,N_19086,N_18858);
and U19444 (N_19444,N_19104,N_18928);
and U19445 (N_19445,N_19052,N_19145);
nor U19446 (N_19446,N_18911,N_18848);
xnor U19447 (N_19447,N_18902,N_18943);
nand U19448 (N_19448,N_19096,N_19097);
or U19449 (N_19449,N_18875,N_19196);
nand U19450 (N_19450,N_19139,N_18994);
nand U19451 (N_19451,N_19023,N_18932);
nand U19452 (N_19452,N_18954,N_19024);
nor U19453 (N_19453,N_18875,N_18989);
and U19454 (N_19454,N_19148,N_19014);
xor U19455 (N_19455,N_18835,N_18993);
xnor U19456 (N_19456,N_18885,N_19006);
nor U19457 (N_19457,N_18818,N_18861);
nand U19458 (N_19458,N_18937,N_19127);
nor U19459 (N_19459,N_19020,N_18971);
nand U19460 (N_19460,N_19011,N_18938);
and U19461 (N_19461,N_18873,N_18821);
or U19462 (N_19462,N_18841,N_19112);
nand U19463 (N_19463,N_18841,N_19148);
or U19464 (N_19464,N_19170,N_18927);
or U19465 (N_19465,N_19199,N_18953);
nand U19466 (N_19466,N_19134,N_19071);
xnor U19467 (N_19467,N_19085,N_18808);
xor U19468 (N_19468,N_19097,N_18831);
and U19469 (N_19469,N_18903,N_19082);
nand U19470 (N_19470,N_19027,N_18988);
nand U19471 (N_19471,N_18917,N_18833);
xnor U19472 (N_19472,N_19168,N_19160);
and U19473 (N_19473,N_19036,N_19150);
or U19474 (N_19474,N_18858,N_18940);
and U19475 (N_19475,N_19037,N_18837);
or U19476 (N_19476,N_18971,N_18936);
nor U19477 (N_19477,N_18892,N_18807);
nand U19478 (N_19478,N_18970,N_18889);
nor U19479 (N_19479,N_18870,N_18845);
nand U19480 (N_19480,N_19048,N_19039);
nor U19481 (N_19481,N_19184,N_18930);
and U19482 (N_19482,N_19136,N_19045);
xnor U19483 (N_19483,N_19095,N_19007);
nor U19484 (N_19484,N_19198,N_19159);
and U19485 (N_19485,N_19111,N_19005);
or U19486 (N_19486,N_19012,N_19144);
xor U19487 (N_19487,N_18939,N_18817);
nand U19488 (N_19488,N_19036,N_19177);
or U19489 (N_19489,N_19171,N_18960);
nor U19490 (N_19490,N_19057,N_18869);
nor U19491 (N_19491,N_18896,N_19196);
nand U19492 (N_19492,N_18825,N_19184);
nor U19493 (N_19493,N_19136,N_19075);
nand U19494 (N_19494,N_19055,N_19027);
xor U19495 (N_19495,N_19092,N_18943);
nand U19496 (N_19496,N_19056,N_18831);
xor U19497 (N_19497,N_18994,N_18820);
or U19498 (N_19498,N_19163,N_18956);
xor U19499 (N_19499,N_18811,N_18995);
nand U19500 (N_19500,N_19066,N_19014);
and U19501 (N_19501,N_18933,N_19100);
xnor U19502 (N_19502,N_18995,N_19123);
nor U19503 (N_19503,N_19099,N_18836);
or U19504 (N_19504,N_19141,N_18853);
or U19505 (N_19505,N_19032,N_18801);
xnor U19506 (N_19506,N_19039,N_18952);
and U19507 (N_19507,N_18831,N_19167);
nand U19508 (N_19508,N_19013,N_19006);
xor U19509 (N_19509,N_19141,N_18831);
xnor U19510 (N_19510,N_19198,N_19113);
and U19511 (N_19511,N_18830,N_18984);
nand U19512 (N_19512,N_18888,N_18884);
nor U19513 (N_19513,N_19077,N_19037);
and U19514 (N_19514,N_18940,N_18854);
nand U19515 (N_19515,N_19026,N_18999);
or U19516 (N_19516,N_19072,N_19027);
and U19517 (N_19517,N_19065,N_18870);
nand U19518 (N_19518,N_19021,N_18803);
or U19519 (N_19519,N_18934,N_19146);
or U19520 (N_19520,N_18862,N_19187);
xor U19521 (N_19521,N_18927,N_18894);
nor U19522 (N_19522,N_19013,N_18811);
or U19523 (N_19523,N_19124,N_18912);
nor U19524 (N_19524,N_18981,N_18892);
nand U19525 (N_19525,N_18867,N_18932);
and U19526 (N_19526,N_18819,N_18869);
nand U19527 (N_19527,N_19016,N_18971);
and U19528 (N_19528,N_19124,N_19105);
or U19529 (N_19529,N_19034,N_18894);
nand U19530 (N_19530,N_19179,N_18801);
and U19531 (N_19531,N_19114,N_18979);
nor U19532 (N_19532,N_18969,N_18864);
and U19533 (N_19533,N_18830,N_19079);
nand U19534 (N_19534,N_18891,N_18807);
xor U19535 (N_19535,N_18973,N_18934);
nand U19536 (N_19536,N_18810,N_18999);
nor U19537 (N_19537,N_19168,N_19051);
or U19538 (N_19538,N_18989,N_19064);
and U19539 (N_19539,N_18899,N_19172);
nor U19540 (N_19540,N_19052,N_18881);
nor U19541 (N_19541,N_19076,N_19118);
nor U19542 (N_19542,N_19119,N_19014);
xnor U19543 (N_19543,N_19183,N_18856);
nand U19544 (N_19544,N_18960,N_18842);
and U19545 (N_19545,N_19187,N_19004);
nor U19546 (N_19546,N_18955,N_18887);
nor U19547 (N_19547,N_18888,N_18807);
nor U19548 (N_19548,N_18827,N_19025);
nand U19549 (N_19549,N_18843,N_18967);
nor U19550 (N_19550,N_18919,N_18925);
nand U19551 (N_19551,N_19091,N_18921);
nand U19552 (N_19552,N_19155,N_19083);
and U19553 (N_19553,N_18876,N_19182);
nand U19554 (N_19554,N_19038,N_18919);
nor U19555 (N_19555,N_18945,N_18901);
and U19556 (N_19556,N_19159,N_18890);
and U19557 (N_19557,N_19107,N_19159);
or U19558 (N_19558,N_19013,N_19039);
nand U19559 (N_19559,N_19152,N_19143);
nand U19560 (N_19560,N_18948,N_18999);
nand U19561 (N_19561,N_18824,N_19038);
or U19562 (N_19562,N_19143,N_18837);
or U19563 (N_19563,N_18906,N_19192);
xor U19564 (N_19564,N_18994,N_18878);
or U19565 (N_19565,N_19121,N_18909);
and U19566 (N_19566,N_18844,N_19035);
nand U19567 (N_19567,N_18900,N_18846);
or U19568 (N_19568,N_19064,N_19159);
nand U19569 (N_19569,N_18902,N_19076);
nor U19570 (N_19570,N_19134,N_19131);
nand U19571 (N_19571,N_19178,N_18908);
xnor U19572 (N_19572,N_18884,N_18816);
nand U19573 (N_19573,N_18967,N_19001);
and U19574 (N_19574,N_18806,N_18923);
and U19575 (N_19575,N_19151,N_19149);
nor U19576 (N_19576,N_19159,N_19146);
xnor U19577 (N_19577,N_19055,N_18968);
and U19578 (N_19578,N_19082,N_19159);
xnor U19579 (N_19579,N_19070,N_19080);
xor U19580 (N_19580,N_19038,N_19056);
and U19581 (N_19581,N_18865,N_19159);
and U19582 (N_19582,N_18923,N_18945);
and U19583 (N_19583,N_19173,N_18924);
xor U19584 (N_19584,N_19143,N_19111);
or U19585 (N_19585,N_18882,N_19172);
or U19586 (N_19586,N_19010,N_18852);
or U19587 (N_19587,N_18857,N_18924);
and U19588 (N_19588,N_19103,N_18898);
nand U19589 (N_19589,N_18807,N_18806);
xnor U19590 (N_19590,N_18830,N_19111);
or U19591 (N_19591,N_18830,N_18895);
xor U19592 (N_19592,N_19140,N_18886);
xor U19593 (N_19593,N_19152,N_19134);
xnor U19594 (N_19594,N_18884,N_18991);
nand U19595 (N_19595,N_19081,N_19083);
and U19596 (N_19596,N_18991,N_18970);
nor U19597 (N_19597,N_18829,N_18956);
and U19598 (N_19598,N_18974,N_19071);
nand U19599 (N_19599,N_19012,N_18880);
xor U19600 (N_19600,N_19249,N_19520);
nand U19601 (N_19601,N_19587,N_19532);
xnor U19602 (N_19602,N_19325,N_19416);
nand U19603 (N_19603,N_19438,N_19549);
and U19604 (N_19604,N_19221,N_19248);
nand U19605 (N_19605,N_19254,N_19452);
or U19606 (N_19606,N_19323,N_19319);
nand U19607 (N_19607,N_19541,N_19295);
xor U19608 (N_19608,N_19457,N_19242);
xnor U19609 (N_19609,N_19312,N_19442);
nand U19610 (N_19610,N_19341,N_19332);
xor U19611 (N_19611,N_19214,N_19412);
nor U19612 (N_19612,N_19326,N_19367);
xor U19613 (N_19613,N_19203,N_19529);
and U19614 (N_19614,N_19553,N_19223);
nand U19615 (N_19615,N_19384,N_19536);
or U19616 (N_19616,N_19405,N_19200);
nor U19617 (N_19617,N_19329,N_19277);
or U19618 (N_19618,N_19379,N_19475);
or U19619 (N_19619,N_19579,N_19521);
nand U19620 (N_19620,N_19216,N_19498);
nor U19621 (N_19621,N_19358,N_19508);
and U19622 (N_19622,N_19361,N_19382);
nor U19623 (N_19623,N_19463,N_19309);
nand U19624 (N_19624,N_19310,N_19528);
nand U19625 (N_19625,N_19511,N_19399);
or U19626 (N_19626,N_19201,N_19461);
xnor U19627 (N_19627,N_19506,N_19206);
and U19628 (N_19628,N_19282,N_19568);
or U19629 (N_19629,N_19264,N_19444);
or U19630 (N_19630,N_19229,N_19231);
nor U19631 (N_19631,N_19265,N_19349);
or U19632 (N_19632,N_19253,N_19403);
and U19633 (N_19633,N_19293,N_19434);
and U19634 (N_19634,N_19429,N_19230);
nor U19635 (N_19635,N_19456,N_19345);
xnor U19636 (N_19636,N_19267,N_19268);
and U19637 (N_19637,N_19394,N_19202);
nand U19638 (N_19638,N_19303,N_19500);
or U19639 (N_19639,N_19531,N_19400);
and U19640 (N_19640,N_19540,N_19241);
nand U19641 (N_19641,N_19365,N_19467);
xnor U19642 (N_19642,N_19523,N_19575);
nor U19643 (N_19643,N_19516,N_19543);
nor U19644 (N_19644,N_19599,N_19330);
nand U19645 (N_19645,N_19313,N_19441);
and U19646 (N_19646,N_19501,N_19559);
and U19647 (N_19647,N_19235,N_19584);
and U19648 (N_19648,N_19477,N_19470);
nand U19649 (N_19649,N_19530,N_19213);
or U19650 (N_19650,N_19443,N_19421);
nand U19651 (N_19651,N_19261,N_19572);
and U19652 (N_19652,N_19390,N_19369);
nor U19653 (N_19653,N_19585,N_19449);
nor U19654 (N_19654,N_19563,N_19574);
or U19655 (N_19655,N_19460,N_19485);
nand U19656 (N_19656,N_19591,N_19245);
nor U19657 (N_19657,N_19354,N_19281);
nor U19658 (N_19658,N_19497,N_19331);
nor U19659 (N_19659,N_19351,N_19492);
or U19660 (N_19660,N_19522,N_19431);
and U19661 (N_19661,N_19411,N_19578);
xnor U19662 (N_19662,N_19550,N_19389);
xor U19663 (N_19663,N_19346,N_19424);
xnor U19664 (N_19664,N_19212,N_19571);
and U19665 (N_19665,N_19385,N_19560);
and U19666 (N_19666,N_19287,N_19474);
and U19667 (N_19667,N_19495,N_19428);
nand U19668 (N_19668,N_19391,N_19592);
nand U19669 (N_19669,N_19573,N_19483);
nand U19670 (N_19670,N_19342,N_19558);
xnor U19671 (N_19671,N_19276,N_19364);
nand U19672 (N_19672,N_19462,N_19238);
xor U19673 (N_19673,N_19533,N_19566);
xnor U19674 (N_19674,N_19598,N_19577);
xor U19675 (N_19675,N_19222,N_19311);
nand U19676 (N_19676,N_19299,N_19482);
and U19677 (N_19677,N_19557,N_19373);
nand U19678 (N_19678,N_19292,N_19469);
and U19679 (N_19679,N_19583,N_19263);
and U19680 (N_19680,N_19564,N_19551);
and U19681 (N_19681,N_19419,N_19445);
and U19682 (N_19682,N_19234,N_19348);
xor U19683 (N_19683,N_19270,N_19320);
and U19684 (N_19684,N_19576,N_19420);
xor U19685 (N_19685,N_19527,N_19339);
nor U19686 (N_19686,N_19322,N_19455);
nor U19687 (N_19687,N_19300,N_19548);
or U19688 (N_19688,N_19464,N_19552);
and U19689 (N_19689,N_19570,N_19340);
or U19690 (N_19690,N_19357,N_19496);
and U19691 (N_19691,N_19526,N_19377);
xnor U19692 (N_19692,N_19204,N_19236);
nand U19693 (N_19693,N_19225,N_19397);
and U19694 (N_19694,N_19362,N_19355);
nand U19695 (N_19695,N_19402,N_19493);
or U19696 (N_19696,N_19279,N_19308);
and U19697 (N_19697,N_19593,N_19374);
nor U19698 (N_19698,N_19580,N_19376);
or U19699 (N_19699,N_19581,N_19209);
or U19700 (N_19700,N_19366,N_19594);
nor U19701 (N_19701,N_19537,N_19383);
nand U19702 (N_19702,N_19510,N_19337);
or U19703 (N_19703,N_19415,N_19343);
or U19704 (N_19704,N_19450,N_19595);
nand U19705 (N_19705,N_19504,N_19274);
nand U19706 (N_19706,N_19418,N_19556);
nand U19707 (N_19707,N_19439,N_19258);
or U19708 (N_19708,N_19318,N_19289);
or U19709 (N_19709,N_19448,N_19280);
and U19710 (N_19710,N_19513,N_19283);
or U19711 (N_19711,N_19459,N_19275);
and U19712 (N_19712,N_19278,N_19215);
or U19713 (N_19713,N_19208,N_19271);
xor U19714 (N_19714,N_19335,N_19233);
nand U19715 (N_19715,N_19368,N_19386);
xnor U19716 (N_19716,N_19205,N_19328);
nand U19717 (N_19717,N_19512,N_19398);
nand U19718 (N_19718,N_19272,N_19306);
nor U19719 (N_19719,N_19453,N_19220);
xor U19720 (N_19720,N_19239,N_19427);
and U19721 (N_19721,N_19244,N_19321);
xnor U19722 (N_19722,N_19250,N_19596);
nand U19723 (N_19723,N_19333,N_19297);
nand U19724 (N_19724,N_19296,N_19435);
and U19725 (N_19725,N_19224,N_19381);
nor U19726 (N_19726,N_19586,N_19471);
nand U19727 (N_19727,N_19494,N_19555);
and U19728 (N_19728,N_19338,N_19324);
and U19729 (N_19729,N_19554,N_19425);
nor U19730 (N_19730,N_19465,N_19207);
or U19731 (N_19731,N_19468,N_19401);
or U19732 (N_19732,N_19519,N_19304);
nor U19733 (N_19733,N_19371,N_19378);
and U19734 (N_19734,N_19505,N_19251);
or U19735 (N_19735,N_19356,N_19436);
xor U19736 (N_19736,N_19247,N_19240);
or U19737 (N_19737,N_19488,N_19350);
and U19738 (N_19738,N_19480,N_19387);
nor U19739 (N_19739,N_19487,N_19478);
or U19740 (N_19740,N_19410,N_19307);
or U19741 (N_19741,N_19298,N_19344);
or U19742 (N_19742,N_19227,N_19433);
or U19743 (N_19743,N_19363,N_19237);
nor U19744 (N_19744,N_19597,N_19290);
nor U19745 (N_19745,N_19243,N_19408);
xnor U19746 (N_19746,N_19285,N_19524);
xor U19747 (N_19747,N_19302,N_19481);
nand U19748 (N_19748,N_19518,N_19490);
xnor U19749 (N_19749,N_19336,N_19316);
nand U19750 (N_19750,N_19525,N_19545);
nor U19751 (N_19751,N_19499,N_19502);
xor U19752 (N_19752,N_19546,N_19538);
nand U19753 (N_19753,N_19269,N_19517);
and U19754 (N_19754,N_19432,N_19217);
and U19755 (N_19755,N_19562,N_19291);
nand U19756 (N_19756,N_19370,N_19347);
and U19757 (N_19757,N_19360,N_19473);
xnor U19758 (N_19758,N_19417,N_19375);
or U19759 (N_19759,N_19305,N_19542);
nor U19760 (N_19760,N_19301,N_19422);
nor U19761 (N_19761,N_19256,N_19388);
or U19762 (N_19762,N_19228,N_19359);
or U19763 (N_19763,N_19476,N_19569);
nor U19764 (N_19764,N_19589,N_19509);
xor U19765 (N_19765,N_19334,N_19380);
and U19766 (N_19766,N_19262,N_19447);
nor U19767 (N_19767,N_19353,N_19582);
and U19768 (N_19768,N_19232,N_19284);
or U19769 (N_19769,N_19454,N_19514);
and U19770 (N_19770,N_19406,N_19539);
nand U19771 (N_19771,N_19315,N_19226);
nand U19772 (N_19772,N_19472,N_19507);
nand U19773 (N_19773,N_19423,N_19260);
or U19774 (N_19774,N_19590,N_19414);
nor U19775 (N_19775,N_19489,N_19491);
nor U19776 (N_19776,N_19430,N_19255);
and U19777 (N_19777,N_19446,N_19479);
xor U19778 (N_19778,N_19396,N_19219);
nor U19779 (N_19779,N_19451,N_19218);
or U19780 (N_19780,N_19286,N_19327);
or U19781 (N_19781,N_19515,N_19404);
nor U19782 (N_19782,N_19588,N_19544);
nor U19783 (N_19783,N_19484,N_19503);
nand U19784 (N_19784,N_19458,N_19565);
nand U19785 (N_19785,N_19395,N_19288);
and U19786 (N_19786,N_19210,N_19211);
nor U19787 (N_19787,N_19393,N_19266);
nand U19788 (N_19788,N_19409,N_19440);
nor U19789 (N_19789,N_19535,N_19413);
or U19790 (N_19790,N_19486,N_19392);
and U19791 (N_19791,N_19466,N_19294);
nor U19792 (N_19792,N_19547,N_19317);
or U19793 (N_19793,N_19561,N_19257);
nand U19794 (N_19794,N_19437,N_19426);
xnor U19795 (N_19795,N_19246,N_19567);
nor U19796 (N_19796,N_19352,N_19314);
or U19797 (N_19797,N_19259,N_19407);
xor U19798 (N_19798,N_19372,N_19252);
and U19799 (N_19799,N_19273,N_19534);
nor U19800 (N_19800,N_19230,N_19263);
and U19801 (N_19801,N_19232,N_19324);
and U19802 (N_19802,N_19239,N_19470);
xor U19803 (N_19803,N_19536,N_19506);
nor U19804 (N_19804,N_19261,N_19369);
nor U19805 (N_19805,N_19264,N_19307);
nor U19806 (N_19806,N_19315,N_19490);
and U19807 (N_19807,N_19462,N_19439);
nor U19808 (N_19808,N_19380,N_19500);
or U19809 (N_19809,N_19379,N_19543);
nand U19810 (N_19810,N_19483,N_19510);
xor U19811 (N_19811,N_19482,N_19315);
xnor U19812 (N_19812,N_19242,N_19576);
and U19813 (N_19813,N_19561,N_19500);
nand U19814 (N_19814,N_19201,N_19510);
nand U19815 (N_19815,N_19367,N_19553);
nor U19816 (N_19816,N_19230,N_19207);
or U19817 (N_19817,N_19358,N_19308);
and U19818 (N_19818,N_19354,N_19522);
nand U19819 (N_19819,N_19485,N_19591);
and U19820 (N_19820,N_19342,N_19482);
nor U19821 (N_19821,N_19329,N_19586);
nor U19822 (N_19822,N_19354,N_19371);
and U19823 (N_19823,N_19292,N_19358);
nand U19824 (N_19824,N_19553,N_19469);
xnor U19825 (N_19825,N_19200,N_19326);
nand U19826 (N_19826,N_19262,N_19464);
and U19827 (N_19827,N_19252,N_19268);
and U19828 (N_19828,N_19465,N_19552);
or U19829 (N_19829,N_19274,N_19320);
nand U19830 (N_19830,N_19267,N_19385);
nand U19831 (N_19831,N_19266,N_19582);
or U19832 (N_19832,N_19259,N_19519);
nand U19833 (N_19833,N_19569,N_19548);
and U19834 (N_19834,N_19241,N_19449);
nand U19835 (N_19835,N_19409,N_19523);
xnor U19836 (N_19836,N_19240,N_19597);
xnor U19837 (N_19837,N_19484,N_19343);
or U19838 (N_19838,N_19258,N_19541);
nor U19839 (N_19839,N_19370,N_19563);
nand U19840 (N_19840,N_19449,N_19309);
and U19841 (N_19841,N_19323,N_19353);
or U19842 (N_19842,N_19583,N_19452);
nor U19843 (N_19843,N_19231,N_19349);
xnor U19844 (N_19844,N_19486,N_19526);
and U19845 (N_19845,N_19452,N_19329);
nor U19846 (N_19846,N_19500,N_19573);
or U19847 (N_19847,N_19399,N_19351);
or U19848 (N_19848,N_19464,N_19400);
or U19849 (N_19849,N_19463,N_19573);
nor U19850 (N_19850,N_19519,N_19209);
nand U19851 (N_19851,N_19389,N_19318);
xor U19852 (N_19852,N_19556,N_19348);
xor U19853 (N_19853,N_19545,N_19420);
and U19854 (N_19854,N_19305,N_19363);
or U19855 (N_19855,N_19420,N_19465);
nand U19856 (N_19856,N_19294,N_19351);
and U19857 (N_19857,N_19512,N_19260);
nand U19858 (N_19858,N_19576,N_19339);
nand U19859 (N_19859,N_19380,N_19235);
nand U19860 (N_19860,N_19380,N_19520);
and U19861 (N_19861,N_19435,N_19324);
and U19862 (N_19862,N_19351,N_19481);
nor U19863 (N_19863,N_19469,N_19360);
nand U19864 (N_19864,N_19343,N_19589);
nor U19865 (N_19865,N_19295,N_19453);
nor U19866 (N_19866,N_19592,N_19236);
xor U19867 (N_19867,N_19201,N_19470);
or U19868 (N_19868,N_19373,N_19597);
or U19869 (N_19869,N_19590,N_19326);
or U19870 (N_19870,N_19309,N_19325);
nor U19871 (N_19871,N_19292,N_19241);
or U19872 (N_19872,N_19202,N_19568);
or U19873 (N_19873,N_19395,N_19460);
nand U19874 (N_19874,N_19512,N_19464);
xor U19875 (N_19875,N_19376,N_19260);
xnor U19876 (N_19876,N_19251,N_19553);
nand U19877 (N_19877,N_19495,N_19443);
nand U19878 (N_19878,N_19595,N_19473);
xnor U19879 (N_19879,N_19256,N_19236);
nor U19880 (N_19880,N_19245,N_19385);
and U19881 (N_19881,N_19278,N_19591);
xor U19882 (N_19882,N_19475,N_19363);
xnor U19883 (N_19883,N_19226,N_19494);
xor U19884 (N_19884,N_19495,N_19503);
and U19885 (N_19885,N_19229,N_19227);
nor U19886 (N_19886,N_19304,N_19593);
nand U19887 (N_19887,N_19353,N_19510);
and U19888 (N_19888,N_19273,N_19590);
and U19889 (N_19889,N_19300,N_19490);
xor U19890 (N_19890,N_19444,N_19206);
or U19891 (N_19891,N_19241,N_19333);
xor U19892 (N_19892,N_19474,N_19412);
nand U19893 (N_19893,N_19349,N_19388);
or U19894 (N_19894,N_19436,N_19532);
xor U19895 (N_19895,N_19419,N_19296);
nor U19896 (N_19896,N_19401,N_19247);
nor U19897 (N_19897,N_19402,N_19551);
nor U19898 (N_19898,N_19399,N_19589);
and U19899 (N_19899,N_19360,N_19272);
nor U19900 (N_19900,N_19444,N_19455);
nand U19901 (N_19901,N_19211,N_19576);
and U19902 (N_19902,N_19284,N_19293);
xnor U19903 (N_19903,N_19443,N_19335);
and U19904 (N_19904,N_19438,N_19526);
and U19905 (N_19905,N_19354,N_19221);
xor U19906 (N_19906,N_19451,N_19334);
nand U19907 (N_19907,N_19273,N_19333);
and U19908 (N_19908,N_19426,N_19214);
and U19909 (N_19909,N_19372,N_19342);
nor U19910 (N_19910,N_19319,N_19232);
nor U19911 (N_19911,N_19206,N_19280);
nor U19912 (N_19912,N_19544,N_19270);
nand U19913 (N_19913,N_19514,N_19329);
nand U19914 (N_19914,N_19337,N_19374);
and U19915 (N_19915,N_19432,N_19357);
and U19916 (N_19916,N_19444,N_19538);
or U19917 (N_19917,N_19539,N_19412);
xnor U19918 (N_19918,N_19478,N_19565);
nor U19919 (N_19919,N_19272,N_19216);
nor U19920 (N_19920,N_19535,N_19534);
xor U19921 (N_19921,N_19563,N_19403);
nor U19922 (N_19922,N_19390,N_19442);
nor U19923 (N_19923,N_19555,N_19565);
nand U19924 (N_19924,N_19205,N_19309);
nor U19925 (N_19925,N_19229,N_19336);
nor U19926 (N_19926,N_19321,N_19254);
nand U19927 (N_19927,N_19365,N_19442);
nand U19928 (N_19928,N_19413,N_19551);
nand U19929 (N_19929,N_19557,N_19448);
nor U19930 (N_19930,N_19454,N_19543);
or U19931 (N_19931,N_19376,N_19545);
and U19932 (N_19932,N_19385,N_19409);
and U19933 (N_19933,N_19317,N_19484);
and U19934 (N_19934,N_19394,N_19459);
xnor U19935 (N_19935,N_19533,N_19364);
nor U19936 (N_19936,N_19485,N_19411);
or U19937 (N_19937,N_19266,N_19512);
nand U19938 (N_19938,N_19541,N_19259);
nand U19939 (N_19939,N_19517,N_19218);
or U19940 (N_19940,N_19205,N_19448);
nor U19941 (N_19941,N_19321,N_19361);
and U19942 (N_19942,N_19546,N_19331);
and U19943 (N_19943,N_19392,N_19442);
nor U19944 (N_19944,N_19373,N_19256);
nor U19945 (N_19945,N_19222,N_19246);
xor U19946 (N_19946,N_19571,N_19406);
xor U19947 (N_19947,N_19284,N_19427);
and U19948 (N_19948,N_19534,N_19395);
nor U19949 (N_19949,N_19274,N_19458);
or U19950 (N_19950,N_19556,N_19562);
nand U19951 (N_19951,N_19243,N_19238);
nand U19952 (N_19952,N_19302,N_19303);
xor U19953 (N_19953,N_19304,N_19227);
nor U19954 (N_19954,N_19337,N_19343);
nand U19955 (N_19955,N_19509,N_19382);
nand U19956 (N_19956,N_19298,N_19569);
nor U19957 (N_19957,N_19513,N_19510);
and U19958 (N_19958,N_19337,N_19350);
nor U19959 (N_19959,N_19283,N_19447);
nand U19960 (N_19960,N_19418,N_19307);
or U19961 (N_19961,N_19501,N_19447);
nor U19962 (N_19962,N_19588,N_19258);
nor U19963 (N_19963,N_19547,N_19509);
nand U19964 (N_19964,N_19473,N_19554);
xnor U19965 (N_19965,N_19350,N_19514);
nor U19966 (N_19966,N_19254,N_19305);
and U19967 (N_19967,N_19469,N_19376);
nand U19968 (N_19968,N_19548,N_19257);
nand U19969 (N_19969,N_19362,N_19352);
nor U19970 (N_19970,N_19400,N_19450);
or U19971 (N_19971,N_19252,N_19216);
nor U19972 (N_19972,N_19505,N_19547);
or U19973 (N_19973,N_19569,N_19340);
nor U19974 (N_19974,N_19334,N_19247);
and U19975 (N_19975,N_19321,N_19595);
and U19976 (N_19976,N_19245,N_19390);
nor U19977 (N_19977,N_19456,N_19263);
xnor U19978 (N_19978,N_19365,N_19385);
xor U19979 (N_19979,N_19430,N_19564);
nand U19980 (N_19980,N_19480,N_19529);
and U19981 (N_19981,N_19517,N_19253);
and U19982 (N_19982,N_19500,N_19599);
xor U19983 (N_19983,N_19216,N_19499);
xor U19984 (N_19984,N_19292,N_19456);
nand U19985 (N_19985,N_19333,N_19319);
nor U19986 (N_19986,N_19272,N_19339);
or U19987 (N_19987,N_19272,N_19343);
nand U19988 (N_19988,N_19459,N_19341);
nand U19989 (N_19989,N_19249,N_19400);
or U19990 (N_19990,N_19466,N_19408);
nor U19991 (N_19991,N_19277,N_19506);
and U19992 (N_19992,N_19496,N_19209);
nor U19993 (N_19993,N_19591,N_19450);
nand U19994 (N_19994,N_19343,N_19308);
nand U19995 (N_19995,N_19524,N_19279);
nand U19996 (N_19996,N_19330,N_19523);
nand U19997 (N_19997,N_19407,N_19548);
xnor U19998 (N_19998,N_19497,N_19486);
nor U19999 (N_19999,N_19382,N_19577);
nand UO_0 (O_0,N_19852,N_19660);
and UO_1 (O_1,N_19871,N_19834);
nand UO_2 (O_2,N_19885,N_19684);
and UO_3 (O_3,N_19945,N_19744);
nor UO_4 (O_4,N_19876,N_19793);
and UO_5 (O_5,N_19908,N_19877);
and UO_6 (O_6,N_19629,N_19889);
and UO_7 (O_7,N_19829,N_19758);
and UO_8 (O_8,N_19708,N_19838);
and UO_9 (O_9,N_19978,N_19714);
and UO_10 (O_10,N_19833,N_19869);
xnor UO_11 (O_11,N_19973,N_19861);
nor UO_12 (O_12,N_19722,N_19902);
nor UO_13 (O_13,N_19711,N_19648);
xnor UO_14 (O_14,N_19915,N_19639);
and UO_15 (O_15,N_19953,N_19907);
and UO_16 (O_16,N_19718,N_19690);
nor UO_17 (O_17,N_19957,N_19811);
xor UO_18 (O_18,N_19842,N_19936);
nand UO_19 (O_19,N_19895,N_19602);
nor UO_20 (O_20,N_19865,N_19770);
nand UO_21 (O_21,N_19797,N_19789);
nand UO_22 (O_22,N_19952,N_19777);
or UO_23 (O_23,N_19712,N_19623);
or UO_24 (O_24,N_19686,N_19783);
nor UO_25 (O_25,N_19649,N_19863);
nand UO_26 (O_26,N_19759,N_19661);
nor UO_27 (O_27,N_19642,N_19761);
nand UO_28 (O_28,N_19676,N_19886);
xnor UO_29 (O_29,N_19940,N_19738);
and UO_30 (O_30,N_19810,N_19665);
xnor UO_31 (O_31,N_19928,N_19728);
xnor UO_32 (O_32,N_19867,N_19643);
nor UO_33 (O_33,N_19990,N_19647);
or UO_34 (O_34,N_19698,N_19827);
nor UO_35 (O_35,N_19788,N_19618);
and UO_36 (O_36,N_19925,N_19949);
nand UO_37 (O_37,N_19839,N_19848);
xor UO_38 (O_38,N_19802,N_19631);
or UO_39 (O_39,N_19812,N_19715);
nor UO_40 (O_40,N_19927,N_19751);
xor UO_41 (O_41,N_19819,N_19970);
and UO_42 (O_42,N_19866,N_19732);
nor UO_43 (O_43,N_19626,N_19693);
and UO_44 (O_44,N_19669,N_19826);
nor UO_45 (O_45,N_19746,N_19946);
nand UO_46 (O_46,N_19769,N_19939);
nand UO_47 (O_47,N_19906,N_19841);
nor UO_48 (O_48,N_19985,N_19914);
and UO_49 (O_49,N_19696,N_19781);
nor UO_50 (O_50,N_19612,N_19960);
and UO_51 (O_51,N_19792,N_19786);
nor UO_52 (O_52,N_19633,N_19723);
nor UO_53 (O_53,N_19646,N_19717);
or UO_54 (O_54,N_19737,N_19736);
or UO_55 (O_55,N_19606,N_19836);
and UO_56 (O_56,N_19859,N_19846);
and UO_57 (O_57,N_19894,N_19893);
and UO_58 (O_58,N_19987,N_19778);
or UO_59 (O_59,N_19713,N_19622);
and UO_60 (O_60,N_19685,N_19765);
nor UO_61 (O_61,N_19641,N_19683);
nand UO_62 (O_62,N_19998,N_19849);
nand UO_63 (O_63,N_19828,N_19733);
nand UO_64 (O_64,N_19837,N_19983);
and UO_65 (O_65,N_19745,N_19860);
nor UO_66 (O_66,N_19697,N_19678);
nor UO_67 (O_67,N_19701,N_19719);
and UO_68 (O_68,N_19899,N_19820);
xor UO_69 (O_69,N_19710,N_19721);
nand UO_70 (O_70,N_19659,N_19991);
or UO_71 (O_71,N_19616,N_19760);
nor UO_72 (O_72,N_19966,N_19785);
nand UO_73 (O_73,N_19607,N_19821);
nor UO_74 (O_74,N_19667,N_19743);
or UO_75 (O_75,N_19795,N_19909);
nor UO_76 (O_76,N_19615,N_19774);
and UO_77 (O_77,N_19924,N_19912);
or UO_78 (O_78,N_19932,N_19603);
xor UO_79 (O_79,N_19694,N_19611);
nor UO_80 (O_80,N_19757,N_19729);
xnor UO_81 (O_81,N_19855,N_19742);
xor UO_82 (O_82,N_19654,N_19823);
or UO_83 (O_83,N_19813,N_19725);
or UO_84 (O_84,N_19720,N_19857);
nor UO_85 (O_85,N_19816,N_19994);
nand UO_86 (O_86,N_19739,N_19993);
nand UO_87 (O_87,N_19609,N_19680);
xnor UO_88 (O_88,N_19879,N_19617);
or UO_89 (O_89,N_19668,N_19806);
nor UO_90 (O_90,N_19943,N_19628);
nor UO_91 (O_91,N_19868,N_19687);
xnor UO_92 (O_92,N_19600,N_19691);
or UO_93 (O_93,N_19805,N_19705);
xnor UO_94 (O_94,N_19692,N_19688);
nor UO_95 (O_95,N_19961,N_19716);
nor UO_96 (O_96,N_19988,N_19755);
nor UO_97 (O_97,N_19898,N_19923);
nor UO_98 (O_98,N_19790,N_19764);
and UO_99 (O_99,N_19968,N_19963);
nand UO_100 (O_100,N_19847,N_19699);
and UO_101 (O_101,N_19964,N_19864);
xor UO_102 (O_102,N_19635,N_19874);
nor UO_103 (O_103,N_19884,N_19619);
or UO_104 (O_104,N_19851,N_19657);
nand UO_105 (O_105,N_19873,N_19824);
nor UO_106 (O_106,N_19891,N_19782);
or UO_107 (O_107,N_19772,N_19892);
xor UO_108 (O_108,N_19844,N_19679);
nand UO_109 (O_109,N_19748,N_19636);
nand UO_110 (O_110,N_19870,N_19858);
nor UO_111 (O_111,N_19651,N_19630);
xor UO_112 (O_112,N_19610,N_19681);
nor UO_113 (O_113,N_19845,N_19637);
and UO_114 (O_114,N_19935,N_19766);
nor UO_115 (O_115,N_19808,N_19703);
nand UO_116 (O_116,N_19883,N_19741);
xor UO_117 (O_117,N_19972,N_19965);
xnor UO_118 (O_118,N_19640,N_19735);
nand UO_119 (O_119,N_19878,N_19904);
xor UO_120 (O_120,N_19601,N_19982);
nand UO_121 (O_121,N_19980,N_19747);
nand UO_122 (O_122,N_19677,N_19780);
and UO_123 (O_123,N_19706,N_19664);
or UO_124 (O_124,N_19627,N_19817);
xnor UO_125 (O_125,N_19634,N_19666);
and UO_126 (O_126,N_19799,N_19913);
nor UO_127 (O_127,N_19605,N_19903);
and UO_128 (O_128,N_19655,N_19709);
nand UO_129 (O_129,N_19776,N_19989);
xnor UO_130 (O_130,N_19768,N_19967);
xnor UO_131 (O_131,N_19673,N_19675);
xor UO_132 (O_132,N_19942,N_19882);
and UO_133 (O_133,N_19814,N_19702);
or UO_134 (O_134,N_19948,N_19791);
nor UO_135 (O_135,N_19921,N_19905);
xor UO_136 (O_136,N_19959,N_19815);
nand UO_137 (O_137,N_19971,N_19663);
xnor UO_138 (O_138,N_19887,N_19888);
or UO_139 (O_139,N_19650,N_19614);
and UO_140 (O_140,N_19807,N_19897);
nor UO_141 (O_141,N_19771,N_19796);
xnor UO_142 (O_142,N_19818,N_19930);
xor UO_143 (O_143,N_19682,N_19944);
nor UO_144 (O_144,N_19929,N_19901);
xor UO_145 (O_145,N_19645,N_19652);
nand UO_146 (O_146,N_19974,N_19608);
xnor UO_147 (O_147,N_19822,N_19934);
and UO_148 (O_148,N_19975,N_19794);
xor UO_149 (O_149,N_19773,N_19954);
nand UO_150 (O_150,N_19997,N_19862);
xor UO_151 (O_151,N_19853,N_19835);
or UO_152 (O_152,N_19996,N_19604);
xor UO_153 (O_153,N_19762,N_19670);
and UO_154 (O_154,N_19933,N_19767);
nor UO_155 (O_155,N_19962,N_19910);
xor UO_156 (O_156,N_19804,N_19749);
and UO_157 (O_157,N_19700,N_19941);
xor UO_158 (O_158,N_19955,N_19724);
and UO_159 (O_159,N_19775,N_19896);
xnor UO_160 (O_160,N_19801,N_19752);
xnor UO_161 (O_161,N_19832,N_19984);
or UO_162 (O_162,N_19632,N_19653);
xor UO_163 (O_163,N_19734,N_19995);
xor UO_164 (O_164,N_19707,N_19638);
xnor UO_165 (O_165,N_19726,N_19875);
nand UO_166 (O_166,N_19992,N_19809);
nor UO_167 (O_167,N_19850,N_19981);
nand UO_168 (O_168,N_19880,N_19872);
xor UO_169 (O_169,N_19856,N_19754);
xor UO_170 (O_170,N_19730,N_19621);
xor UO_171 (O_171,N_19976,N_19854);
nor UO_172 (O_172,N_19740,N_19919);
nor UO_173 (O_173,N_19951,N_19727);
and UO_174 (O_174,N_19979,N_19831);
xnor UO_175 (O_175,N_19999,N_19843);
nor UO_176 (O_176,N_19900,N_19920);
nor UO_177 (O_177,N_19986,N_19958);
xor UO_178 (O_178,N_19763,N_19779);
nor UO_179 (O_179,N_19620,N_19840);
and UO_180 (O_180,N_19644,N_19658);
nor UO_181 (O_181,N_19937,N_19938);
xor UO_182 (O_182,N_19625,N_19784);
nand UO_183 (O_183,N_19956,N_19704);
nand UO_184 (O_184,N_19787,N_19753);
nand UO_185 (O_185,N_19969,N_19931);
or UO_186 (O_186,N_19830,N_19881);
nor UO_187 (O_187,N_19656,N_19918);
nand UO_188 (O_188,N_19798,N_19800);
and UO_189 (O_189,N_19731,N_19689);
nand UO_190 (O_190,N_19671,N_19624);
nand UO_191 (O_191,N_19917,N_19890);
nor UO_192 (O_192,N_19756,N_19926);
nand UO_193 (O_193,N_19916,N_19911);
and UO_194 (O_194,N_19674,N_19695);
nor UO_195 (O_195,N_19947,N_19825);
and UO_196 (O_196,N_19662,N_19950);
or UO_197 (O_197,N_19750,N_19977);
or UO_198 (O_198,N_19613,N_19803);
nand UO_199 (O_199,N_19672,N_19922);
and UO_200 (O_200,N_19900,N_19723);
xnor UO_201 (O_201,N_19658,N_19811);
xor UO_202 (O_202,N_19989,N_19928);
xnor UO_203 (O_203,N_19930,N_19616);
nor UO_204 (O_204,N_19701,N_19793);
and UO_205 (O_205,N_19834,N_19708);
xnor UO_206 (O_206,N_19868,N_19684);
and UO_207 (O_207,N_19916,N_19675);
or UO_208 (O_208,N_19937,N_19611);
and UO_209 (O_209,N_19740,N_19934);
and UO_210 (O_210,N_19794,N_19804);
and UO_211 (O_211,N_19981,N_19980);
or UO_212 (O_212,N_19834,N_19807);
and UO_213 (O_213,N_19700,N_19635);
nor UO_214 (O_214,N_19649,N_19867);
nand UO_215 (O_215,N_19644,N_19848);
nand UO_216 (O_216,N_19834,N_19885);
xnor UO_217 (O_217,N_19654,N_19961);
and UO_218 (O_218,N_19736,N_19919);
nand UO_219 (O_219,N_19685,N_19823);
nand UO_220 (O_220,N_19702,N_19673);
nand UO_221 (O_221,N_19852,N_19903);
xor UO_222 (O_222,N_19752,N_19945);
and UO_223 (O_223,N_19771,N_19963);
nor UO_224 (O_224,N_19981,N_19642);
xor UO_225 (O_225,N_19878,N_19921);
and UO_226 (O_226,N_19709,N_19928);
nor UO_227 (O_227,N_19840,N_19784);
xor UO_228 (O_228,N_19752,N_19759);
and UO_229 (O_229,N_19986,N_19750);
and UO_230 (O_230,N_19873,N_19687);
xnor UO_231 (O_231,N_19852,N_19968);
nand UO_232 (O_232,N_19642,N_19658);
xor UO_233 (O_233,N_19986,N_19851);
or UO_234 (O_234,N_19809,N_19702);
nand UO_235 (O_235,N_19827,N_19636);
xnor UO_236 (O_236,N_19894,N_19927);
xnor UO_237 (O_237,N_19921,N_19936);
or UO_238 (O_238,N_19841,N_19673);
nand UO_239 (O_239,N_19870,N_19766);
or UO_240 (O_240,N_19619,N_19708);
nor UO_241 (O_241,N_19882,N_19900);
xor UO_242 (O_242,N_19980,N_19802);
or UO_243 (O_243,N_19950,N_19686);
or UO_244 (O_244,N_19954,N_19649);
and UO_245 (O_245,N_19907,N_19908);
nand UO_246 (O_246,N_19898,N_19688);
and UO_247 (O_247,N_19891,N_19739);
or UO_248 (O_248,N_19921,N_19799);
or UO_249 (O_249,N_19908,N_19715);
nor UO_250 (O_250,N_19831,N_19721);
or UO_251 (O_251,N_19631,N_19751);
nand UO_252 (O_252,N_19784,N_19604);
xnor UO_253 (O_253,N_19725,N_19731);
nor UO_254 (O_254,N_19817,N_19798);
and UO_255 (O_255,N_19715,N_19965);
or UO_256 (O_256,N_19699,N_19777);
nor UO_257 (O_257,N_19713,N_19797);
and UO_258 (O_258,N_19787,N_19912);
and UO_259 (O_259,N_19750,N_19700);
and UO_260 (O_260,N_19611,N_19926);
nand UO_261 (O_261,N_19770,N_19759);
xor UO_262 (O_262,N_19854,N_19659);
nor UO_263 (O_263,N_19961,N_19816);
and UO_264 (O_264,N_19656,N_19894);
nor UO_265 (O_265,N_19889,N_19930);
and UO_266 (O_266,N_19727,N_19831);
and UO_267 (O_267,N_19656,N_19998);
nand UO_268 (O_268,N_19611,N_19917);
nand UO_269 (O_269,N_19626,N_19639);
nand UO_270 (O_270,N_19827,N_19630);
and UO_271 (O_271,N_19990,N_19854);
nand UO_272 (O_272,N_19779,N_19685);
xor UO_273 (O_273,N_19775,N_19690);
nand UO_274 (O_274,N_19914,N_19668);
xor UO_275 (O_275,N_19733,N_19993);
nand UO_276 (O_276,N_19768,N_19723);
and UO_277 (O_277,N_19646,N_19604);
xor UO_278 (O_278,N_19873,N_19659);
xnor UO_279 (O_279,N_19835,N_19916);
or UO_280 (O_280,N_19980,N_19619);
and UO_281 (O_281,N_19806,N_19988);
and UO_282 (O_282,N_19619,N_19935);
xor UO_283 (O_283,N_19855,N_19789);
and UO_284 (O_284,N_19694,N_19731);
or UO_285 (O_285,N_19857,N_19887);
xnor UO_286 (O_286,N_19889,N_19686);
or UO_287 (O_287,N_19601,N_19964);
or UO_288 (O_288,N_19986,N_19869);
and UO_289 (O_289,N_19730,N_19846);
nand UO_290 (O_290,N_19750,N_19840);
nor UO_291 (O_291,N_19815,N_19798);
and UO_292 (O_292,N_19773,N_19725);
or UO_293 (O_293,N_19675,N_19791);
nand UO_294 (O_294,N_19959,N_19978);
or UO_295 (O_295,N_19917,N_19610);
nor UO_296 (O_296,N_19779,N_19997);
and UO_297 (O_297,N_19754,N_19877);
nor UO_298 (O_298,N_19956,N_19998);
xnor UO_299 (O_299,N_19804,N_19972);
nand UO_300 (O_300,N_19736,N_19861);
and UO_301 (O_301,N_19850,N_19608);
xnor UO_302 (O_302,N_19954,N_19681);
and UO_303 (O_303,N_19950,N_19891);
and UO_304 (O_304,N_19794,N_19714);
xnor UO_305 (O_305,N_19937,N_19701);
or UO_306 (O_306,N_19624,N_19799);
and UO_307 (O_307,N_19739,N_19655);
or UO_308 (O_308,N_19900,N_19883);
nand UO_309 (O_309,N_19677,N_19681);
nand UO_310 (O_310,N_19942,N_19968);
xnor UO_311 (O_311,N_19663,N_19660);
nand UO_312 (O_312,N_19901,N_19634);
or UO_313 (O_313,N_19997,N_19878);
xnor UO_314 (O_314,N_19852,N_19961);
or UO_315 (O_315,N_19721,N_19613);
and UO_316 (O_316,N_19994,N_19743);
and UO_317 (O_317,N_19826,N_19853);
and UO_318 (O_318,N_19676,N_19736);
or UO_319 (O_319,N_19742,N_19850);
or UO_320 (O_320,N_19857,N_19808);
or UO_321 (O_321,N_19956,N_19944);
nor UO_322 (O_322,N_19814,N_19642);
nand UO_323 (O_323,N_19953,N_19731);
and UO_324 (O_324,N_19640,N_19806);
xor UO_325 (O_325,N_19647,N_19909);
nand UO_326 (O_326,N_19638,N_19898);
nand UO_327 (O_327,N_19646,N_19833);
xor UO_328 (O_328,N_19974,N_19644);
or UO_329 (O_329,N_19624,N_19887);
xnor UO_330 (O_330,N_19828,N_19672);
or UO_331 (O_331,N_19845,N_19999);
nor UO_332 (O_332,N_19610,N_19726);
or UO_333 (O_333,N_19904,N_19976);
or UO_334 (O_334,N_19654,N_19872);
xnor UO_335 (O_335,N_19965,N_19758);
xnor UO_336 (O_336,N_19752,N_19828);
nand UO_337 (O_337,N_19745,N_19962);
and UO_338 (O_338,N_19623,N_19803);
or UO_339 (O_339,N_19999,N_19907);
nand UO_340 (O_340,N_19882,N_19994);
nor UO_341 (O_341,N_19699,N_19791);
or UO_342 (O_342,N_19610,N_19974);
or UO_343 (O_343,N_19762,N_19652);
or UO_344 (O_344,N_19746,N_19606);
nand UO_345 (O_345,N_19786,N_19753);
xnor UO_346 (O_346,N_19850,N_19888);
or UO_347 (O_347,N_19900,N_19648);
nor UO_348 (O_348,N_19658,N_19624);
or UO_349 (O_349,N_19686,N_19661);
nor UO_350 (O_350,N_19649,N_19763);
and UO_351 (O_351,N_19680,N_19847);
xnor UO_352 (O_352,N_19879,N_19823);
xnor UO_353 (O_353,N_19976,N_19627);
xnor UO_354 (O_354,N_19617,N_19962);
or UO_355 (O_355,N_19642,N_19785);
and UO_356 (O_356,N_19950,N_19756);
and UO_357 (O_357,N_19771,N_19843);
and UO_358 (O_358,N_19867,N_19918);
and UO_359 (O_359,N_19990,N_19788);
nand UO_360 (O_360,N_19806,N_19603);
xor UO_361 (O_361,N_19655,N_19877);
nand UO_362 (O_362,N_19644,N_19801);
or UO_363 (O_363,N_19610,N_19833);
nor UO_364 (O_364,N_19952,N_19787);
nand UO_365 (O_365,N_19826,N_19774);
and UO_366 (O_366,N_19970,N_19624);
and UO_367 (O_367,N_19669,N_19798);
or UO_368 (O_368,N_19911,N_19904);
or UO_369 (O_369,N_19848,N_19896);
nor UO_370 (O_370,N_19857,N_19981);
and UO_371 (O_371,N_19856,N_19850);
nor UO_372 (O_372,N_19630,N_19745);
nor UO_373 (O_373,N_19896,N_19664);
nor UO_374 (O_374,N_19648,N_19755);
nor UO_375 (O_375,N_19627,N_19631);
xnor UO_376 (O_376,N_19744,N_19788);
and UO_377 (O_377,N_19853,N_19804);
xnor UO_378 (O_378,N_19693,N_19976);
or UO_379 (O_379,N_19891,N_19788);
or UO_380 (O_380,N_19780,N_19983);
and UO_381 (O_381,N_19610,N_19772);
or UO_382 (O_382,N_19709,N_19604);
nor UO_383 (O_383,N_19845,N_19657);
nor UO_384 (O_384,N_19721,N_19770);
or UO_385 (O_385,N_19675,N_19635);
and UO_386 (O_386,N_19833,N_19785);
nor UO_387 (O_387,N_19883,N_19847);
and UO_388 (O_388,N_19960,N_19642);
xor UO_389 (O_389,N_19700,N_19638);
nor UO_390 (O_390,N_19723,N_19881);
and UO_391 (O_391,N_19608,N_19682);
nor UO_392 (O_392,N_19721,N_19793);
and UO_393 (O_393,N_19733,N_19660);
xnor UO_394 (O_394,N_19645,N_19601);
or UO_395 (O_395,N_19786,N_19907);
xnor UO_396 (O_396,N_19908,N_19619);
nor UO_397 (O_397,N_19972,N_19656);
and UO_398 (O_398,N_19847,N_19695);
nor UO_399 (O_399,N_19802,N_19775);
or UO_400 (O_400,N_19748,N_19669);
nand UO_401 (O_401,N_19655,N_19932);
nor UO_402 (O_402,N_19925,N_19860);
or UO_403 (O_403,N_19969,N_19698);
xor UO_404 (O_404,N_19880,N_19956);
xor UO_405 (O_405,N_19923,N_19878);
xnor UO_406 (O_406,N_19919,N_19896);
xor UO_407 (O_407,N_19832,N_19869);
and UO_408 (O_408,N_19935,N_19888);
nor UO_409 (O_409,N_19986,N_19948);
nor UO_410 (O_410,N_19620,N_19930);
or UO_411 (O_411,N_19791,N_19603);
or UO_412 (O_412,N_19970,N_19891);
xor UO_413 (O_413,N_19862,N_19955);
or UO_414 (O_414,N_19629,N_19760);
or UO_415 (O_415,N_19691,N_19668);
xnor UO_416 (O_416,N_19717,N_19643);
xor UO_417 (O_417,N_19795,N_19788);
or UO_418 (O_418,N_19649,N_19718);
and UO_419 (O_419,N_19918,N_19772);
nand UO_420 (O_420,N_19655,N_19957);
nor UO_421 (O_421,N_19985,N_19733);
nor UO_422 (O_422,N_19929,N_19928);
nor UO_423 (O_423,N_19932,N_19980);
xnor UO_424 (O_424,N_19757,N_19933);
nor UO_425 (O_425,N_19754,N_19612);
nand UO_426 (O_426,N_19720,N_19891);
nand UO_427 (O_427,N_19797,N_19770);
xor UO_428 (O_428,N_19627,N_19666);
and UO_429 (O_429,N_19755,N_19857);
nand UO_430 (O_430,N_19893,N_19886);
and UO_431 (O_431,N_19855,N_19749);
xor UO_432 (O_432,N_19814,N_19638);
and UO_433 (O_433,N_19767,N_19943);
xnor UO_434 (O_434,N_19754,N_19783);
or UO_435 (O_435,N_19739,N_19667);
xnor UO_436 (O_436,N_19933,N_19760);
or UO_437 (O_437,N_19661,N_19971);
nor UO_438 (O_438,N_19643,N_19721);
or UO_439 (O_439,N_19772,N_19723);
or UO_440 (O_440,N_19612,N_19924);
nand UO_441 (O_441,N_19850,N_19741);
nor UO_442 (O_442,N_19618,N_19701);
xnor UO_443 (O_443,N_19836,N_19947);
nor UO_444 (O_444,N_19611,N_19727);
and UO_445 (O_445,N_19826,N_19640);
nand UO_446 (O_446,N_19880,N_19909);
xnor UO_447 (O_447,N_19993,N_19671);
or UO_448 (O_448,N_19779,N_19666);
nor UO_449 (O_449,N_19749,N_19666);
and UO_450 (O_450,N_19966,N_19993);
and UO_451 (O_451,N_19711,N_19955);
and UO_452 (O_452,N_19854,N_19892);
xnor UO_453 (O_453,N_19937,N_19879);
nor UO_454 (O_454,N_19935,N_19644);
xnor UO_455 (O_455,N_19917,N_19993);
xnor UO_456 (O_456,N_19840,N_19926);
nand UO_457 (O_457,N_19758,N_19873);
or UO_458 (O_458,N_19669,N_19783);
xnor UO_459 (O_459,N_19717,N_19861);
nor UO_460 (O_460,N_19629,N_19989);
or UO_461 (O_461,N_19728,N_19893);
nor UO_462 (O_462,N_19826,N_19648);
nor UO_463 (O_463,N_19709,N_19874);
or UO_464 (O_464,N_19931,N_19790);
nor UO_465 (O_465,N_19926,N_19641);
xnor UO_466 (O_466,N_19742,N_19754);
or UO_467 (O_467,N_19948,N_19604);
nand UO_468 (O_468,N_19957,N_19642);
nor UO_469 (O_469,N_19770,N_19884);
or UO_470 (O_470,N_19951,N_19651);
and UO_471 (O_471,N_19993,N_19902);
xor UO_472 (O_472,N_19798,N_19911);
or UO_473 (O_473,N_19639,N_19939);
or UO_474 (O_474,N_19732,N_19979);
xnor UO_475 (O_475,N_19744,N_19702);
xor UO_476 (O_476,N_19759,N_19911);
or UO_477 (O_477,N_19818,N_19869);
and UO_478 (O_478,N_19672,N_19671);
nor UO_479 (O_479,N_19875,N_19971);
nand UO_480 (O_480,N_19916,N_19889);
nand UO_481 (O_481,N_19839,N_19624);
nand UO_482 (O_482,N_19840,N_19906);
or UO_483 (O_483,N_19864,N_19941);
nor UO_484 (O_484,N_19768,N_19675);
or UO_485 (O_485,N_19625,N_19637);
or UO_486 (O_486,N_19843,N_19750);
or UO_487 (O_487,N_19704,N_19733);
or UO_488 (O_488,N_19953,N_19630);
or UO_489 (O_489,N_19982,N_19908);
and UO_490 (O_490,N_19632,N_19626);
nor UO_491 (O_491,N_19899,N_19792);
nand UO_492 (O_492,N_19676,N_19940);
or UO_493 (O_493,N_19836,N_19946);
or UO_494 (O_494,N_19772,N_19766);
nor UO_495 (O_495,N_19870,N_19968);
xnor UO_496 (O_496,N_19743,N_19856);
nand UO_497 (O_497,N_19639,N_19970);
nor UO_498 (O_498,N_19795,N_19719);
xnor UO_499 (O_499,N_19644,N_19942);
xnor UO_500 (O_500,N_19628,N_19726);
or UO_501 (O_501,N_19877,N_19802);
or UO_502 (O_502,N_19703,N_19640);
xnor UO_503 (O_503,N_19863,N_19731);
nor UO_504 (O_504,N_19692,N_19739);
and UO_505 (O_505,N_19915,N_19994);
nand UO_506 (O_506,N_19892,N_19858);
and UO_507 (O_507,N_19825,N_19871);
or UO_508 (O_508,N_19684,N_19901);
xnor UO_509 (O_509,N_19930,N_19819);
and UO_510 (O_510,N_19945,N_19911);
and UO_511 (O_511,N_19951,N_19995);
nor UO_512 (O_512,N_19847,N_19838);
nand UO_513 (O_513,N_19783,N_19921);
or UO_514 (O_514,N_19778,N_19762);
nand UO_515 (O_515,N_19912,N_19921);
nor UO_516 (O_516,N_19706,N_19876);
xor UO_517 (O_517,N_19882,N_19659);
nor UO_518 (O_518,N_19725,N_19876);
and UO_519 (O_519,N_19731,N_19926);
or UO_520 (O_520,N_19679,N_19939);
and UO_521 (O_521,N_19856,N_19775);
and UO_522 (O_522,N_19655,N_19865);
xor UO_523 (O_523,N_19921,N_19677);
nand UO_524 (O_524,N_19735,N_19728);
nor UO_525 (O_525,N_19831,N_19665);
xor UO_526 (O_526,N_19701,N_19843);
and UO_527 (O_527,N_19608,N_19646);
nor UO_528 (O_528,N_19680,N_19978);
or UO_529 (O_529,N_19990,N_19725);
nor UO_530 (O_530,N_19727,N_19783);
nand UO_531 (O_531,N_19830,N_19853);
nand UO_532 (O_532,N_19951,N_19759);
and UO_533 (O_533,N_19672,N_19915);
nor UO_534 (O_534,N_19793,N_19851);
nor UO_535 (O_535,N_19683,N_19792);
nor UO_536 (O_536,N_19890,N_19816);
nand UO_537 (O_537,N_19980,N_19786);
xor UO_538 (O_538,N_19877,N_19671);
and UO_539 (O_539,N_19805,N_19821);
and UO_540 (O_540,N_19606,N_19967);
nor UO_541 (O_541,N_19779,N_19602);
or UO_542 (O_542,N_19663,N_19800);
nand UO_543 (O_543,N_19684,N_19879);
nor UO_544 (O_544,N_19605,N_19830);
or UO_545 (O_545,N_19748,N_19611);
xor UO_546 (O_546,N_19714,N_19964);
and UO_547 (O_547,N_19734,N_19897);
nor UO_548 (O_548,N_19803,N_19951);
nand UO_549 (O_549,N_19762,N_19968);
xnor UO_550 (O_550,N_19987,N_19958);
or UO_551 (O_551,N_19899,N_19654);
nor UO_552 (O_552,N_19980,N_19938);
or UO_553 (O_553,N_19861,N_19804);
and UO_554 (O_554,N_19941,N_19940);
or UO_555 (O_555,N_19674,N_19837);
and UO_556 (O_556,N_19900,N_19949);
nor UO_557 (O_557,N_19775,N_19698);
nand UO_558 (O_558,N_19992,N_19910);
xnor UO_559 (O_559,N_19987,N_19898);
xor UO_560 (O_560,N_19910,N_19757);
xor UO_561 (O_561,N_19625,N_19860);
and UO_562 (O_562,N_19973,N_19655);
or UO_563 (O_563,N_19906,N_19652);
or UO_564 (O_564,N_19678,N_19634);
and UO_565 (O_565,N_19621,N_19802);
nand UO_566 (O_566,N_19829,N_19812);
nand UO_567 (O_567,N_19790,N_19611);
nor UO_568 (O_568,N_19737,N_19982);
and UO_569 (O_569,N_19917,N_19775);
nand UO_570 (O_570,N_19762,N_19841);
xor UO_571 (O_571,N_19759,N_19780);
nand UO_572 (O_572,N_19866,N_19714);
xnor UO_573 (O_573,N_19843,N_19986);
xor UO_574 (O_574,N_19723,N_19735);
nand UO_575 (O_575,N_19818,N_19934);
nand UO_576 (O_576,N_19826,N_19773);
nor UO_577 (O_577,N_19653,N_19984);
and UO_578 (O_578,N_19979,N_19699);
nand UO_579 (O_579,N_19749,N_19791);
nor UO_580 (O_580,N_19605,N_19700);
nor UO_581 (O_581,N_19886,N_19706);
or UO_582 (O_582,N_19951,N_19755);
and UO_583 (O_583,N_19777,N_19600);
or UO_584 (O_584,N_19720,N_19814);
nand UO_585 (O_585,N_19808,N_19907);
nor UO_586 (O_586,N_19789,N_19957);
xor UO_587 (O_587,N_19822,N_19678);
nand UO_588 (O_588,N_19758,N_19619);
nand UO_589 (O_589,N_19900,N_19916);
nand UO_590 (O_590,N_19864,N_19629);
nor UO_591 (O_591,N_19637,N_19721);
and UO_592 (O_592,N_19902,N_19739);
nand UO_593 (O_593,N_19950,N_19835);
xnor UO_594 (O_594,N_19885,N_19621);
or UO_595 (O_595,N_19981,N_19828);
or UO_596 (O_596,N_19824,N_19916);
xor UO_597 (O_597,N_19617,N_19742);
xor UO_598 (O_598,N_19643,N_19669);
nor UO_599 (O_599,N_19661,N_19924);
nand UO_600 (O_600,N_19686,N_19943);
nor UO_601 (O_601,N_19860,N_19845);
or UO_602 (O_602,N_19953,N_19896);
or UO_603 (O_603,N_19963,N_19978);
nand UO_604 (O_604,N_19648,N_19707);
nand UO_605 (O_605,N_19969,N_19879);
nand UO_606 (O_606,N_19900,N_19687);
and UO_607 (O_607,N_19993,N_19992);
nor UO_608 (O_608,N_19971,N_19617);
and UO_609 (O_609,N_19736,N_19937);
and UO_610 (O_610,N_19842,N_19872);
nor UO_611 (O_611,N_19625,N_19968);
nor UO_612 (O_612,N_19883,N_19749);
and UO_613 (O_613,N_19871,N_19660);
nand UO_614 (O_614,N_19665,N_19984);
nand UO_615 (O_615,N_19941,N_19727);
and UO_616 (O_616,N_19851,N_19669);
xnor UO_617 (O_617,N_19981,N_19889);
or UO_618 (O_618,N_19664,N_19695);
and UO_619 (O_619,N_19871,N_19939);
nor UO_620 (O_620,N_19949,N_19858);
xor UO_621 (O_621,N_19965,N_19947);
nand UO_622 (O_622,N_19753,N_19618);
nand UO_623 (O_623,N_19670,N_19770);
xnor UO_624 (O_624,N_19695,N_19920);
xnor UO_625 (O_625,N_19870,N_19686);
nand UO_626 (O_626,N_19773,N_19976);
xnor UO_627 (O_627,N_19799,N_19648);
nor UO_628 (O_628,N_19699,N_19614);
xor UO_629 (O_629,N_19712,N_19707);
or UO_630 (O_630,N_19888,N_19740);
or UO_631 (O_631,N_19753,N_19850);
or UO_632 (O_632,N_19642,N_19813);
or UO_633 (O_633,N_19942,N_19751);
nand UO_634 (O_634,N_19684,N_19889);
nor UO_635 (O_635,N_19922,N_19667);
xnor UO_636 (O_636,N_19956,N_19783);
nand UO_637 (O_637,N_19961,N_19731);
and UO_638 (O_638,N_19668,N_19809);
or UO_639 (O_639,N_19972,N_19989);
nor UO_640 (O_640,N_19884,N_19962);
nor UO_641 (O_641,N_19600,N_19694);
and UO_642 (O_642,N_19785,N_19982);
nor UO_643 (O_643,N_19887,N_19720);
and UO_644 (O_644,N_19658,N_19680);
nor UO_645 (O_645,N_19893,N_19904);
or UO_646 (O_646,N_19995,N_19652);
xor UO_647 (O_647,N_19789,N_19922);
and UO_648 (O_648,N_19832,N_19938);
nor UO_649 (O_649,N_19638,N_19803);
nand UO_650 (O_650,N_19633,N_19836);
nor UO_651 (O_651,N_19884,N_19926);
xor UO_652 (O_652,N_19911,N_19615);
nor UO_653 (O_653,N_19844,N_19849);
and UO_654 (O_654,N_19701,N_19988);
nor UO_655 (O_655,N_19979,N_19736);
or UO_656 (O_656,N_19921,N_19622);
xor UO_657 (O_657,N_19915,N_19615);
and UO_658 (O_658,N_19633,N_19913);
and UO_659 (O_659,N_19935,N_19667);
xnor UO_660 (O_660,N_19788,N_19917);
nor UO_661 (O_661,N_19670,N_19726);
nand UO_662 (O_662,N_19815,N_19699);
nand UO_663 (O_663,N_19829,N_19872);
nor UO_664 (O_664,N_19705,N_19718);
nor UO_665 (O_665,N_19897,N_19708);
and UO_666 (O_666,N_19612,N_19658);
and UO_667 (O_667,N_19853,N_19669);
xor UO_668 (O_668,N_19649,N_19603);
xnor UO_669 (O_669,N_19891,N_19875);
nand UO_670 (O_670,N_19866,N_19615);
and UO_671 (O_671,N_19715,N_19929);
xor UO_672 (O_672,N_19867,N_19866);
nand UO_673 (O_673,N_19981,N_19968);
nor UO_674 (O_674,N_19975,N_19801);
nand UO_675 (O_675,N_19862,N_19734);
or UO_676 (O_676,N_19820,N_19729);
xor UO_677 (O_677,N_19639,N_19685);
and UO_678 (O_678,N_19758,N_19629);
nor UO_679 (O_679,N_19933,N_19755);
xor UO_680 (O_680,N_19603,N_19767);
nor UO_681 (O_681,N_19600,N_19955);
nor UO_682 (O_682,N_19951,N_19931);
nand UO_683 (O_683,N_19648,N_19836);
and UO_684 (O_684,N_19616,N_19904);
and UO_685 (O_685,N_19993,N_19764);
nor UO_686 (O_686,N_19660,N_19611);
nor UO_687 (O_687,N_19680,N_19834);
and UO_688 (O_688,N_19610,N_19765);
and UO_689 (O_689,N_19973,N_19794);
nand UO_690 (O_690,N_19774,N_19744);
and UO_691 (O_691,N_19698,N_19687);
and UO_692 (O_692,N_19634,N_19684);
and UO_693 (O_693,N_19782,N_19745);
or UO_694 (O_694,N_19784,N_19964);
and UO_695 (O_695,N_19605,N_19652);
nor UO_696 (O_696,N_19629,N_19706);
xor UO_697 (O_697,N_19731,N_19859);
or UO_698 (O_698,N_19605,N_19975);
or UO_699 (O_699,N_19647,N_19784);
nand UO_700 (O_700,N_19780,N_19721);
or UO_701 (O_701,N_19841,N_19810);
xnor UO_702 (O_702,N_19873,N_19814);
nor UO_703 (O_703,N_19680,N_19831);
nor UO_704 (O_704,N_19813,N_19659);
xor UO_705 (O_705,N_19939,N_19971);
nor UO_706 (O_706,N_19649,N_19788);
and UO_707 (O_707,N_19818,N_19797);
xor UO_708 (O_708,N_19824,N_19729);
xnor UO_709 (O_709,N_19974,N_19808);
or UO_710 (O_710,N_19879,N_19725);
nand UO_711 (O_711,N_19907,N_19602);
xnor UO_712 (O_712,N_19778,N_19837);
and UO_713 (O_713,N_19789,N_19683);
nand UO_714 (O_714,N_19845,N_19629);
or UO_715 (O_715,N_19985,N_19603);
xnor UO_716 (O_716,N_19632,N_19962);
nor UO_717 (O_717,N_19644,N_19998);
nor UO_718 (O_718,N_19914,N_19844);
nor UO_719 (O_719,N_19947,N_19708);
xor UO_720 (O_720,N_19744,N_19840);
and UO_721 (O_721,N_19628,N_19693);
and UO_722 (O_722,N_19800,N_19847);
nor UO_723 (O_723,N_19750,N_19627);
xor UO_724 (O_724,N_19643,N_19980);
nor UO_725 (O_725,N_19849,N_19805);
nand UO_726 (O_726,N_19602,N_19684);
or UO_727 (O_727,N_19613,N_19875);
nor UO_728 (O_728,N_19800,N_19680);
and UO_729 (O_729,N_19790,N_19886);
nor UO_730 (O_730,N_19974,N_19823);
nand UO_731 (O_731,N_19985,N_19918);
nand UO_732 (O_732,N_19682,N_19885);
or UO_733 (O_733,N_19649,N_19919);
nor UO_734 (O_734,N_19905,N_19943);
xor UO_735 (O_735,N_19902,N_19693);
and UO_736 (O_736,N_19764,N_19752);
nand UO_737 (O_737,N_19653,N_19779);
and UO_738 (O_738,N_19609,N_19630);
or UO_739 (O_739,N_19773,N_19623);
xnor UO_740 (O_740,N_19952,N_19846);
nor UO_741 (O_741,N_19896,N_19842);
nand UO_742 (O_742,N_19652,N_19763);
xor UO_743 (O_743,N_19741,N_19628);
xnor UO_744 (O_744,N_19708,N_19638);
xnor UO_745 (O_745,N_19769,N_19787);
or UO_746 (O_746,N_19917,N_19689);
nand UO_747 (O_747,N_19998,N_19650);
nand UO_748 (O_748,N_19826,N_19636);
xor UO_749 (O_749,N_19752,N_19710);
nor UO_750 (O_750,N_19758,N_19946);
and UO_751 (O_751,N_19669,N_19817);
nand UO_752 (O_752,N_19841,N_19931);
xor UO_753 (O_753,N_19703,N_19990);
and UO_754 (O_754,N_19764,N_19953);
or UO_755 (O_755,N_19923,N_19696);
and UO_756 (O_756,N_19657,N_19613);
nor UO_757 (O_757,N_19665,N_19630);
nor UO_758 (O_758,N_19814,N_19620);
or UO_759 (O_759,N_19662,N_19913);
or UO_760 (O_760,N_19857,N_19798);
nand UO_761 (O_761,N_19660,N_19908);
and UO_762 (O_762,N_19606,N_19638);
xor UO_763 (O_763,N_19850,N_19796);
xor UO_764 (O_764,N_19731,N_19804);
or UO_765 (O_765,N_19879,N_19890);
or UO_766 (O_766,N_19675,N_19842);
nor UO_767 (O_767,N_19907,N_19679);
nor UO_768 (O_768,N_19977,N_19734);
and UO_769 (O_769,N_19708,N_19731);
nand UO_770 (O_770,N_19772,N_19900);
nor UO_771 (O_771,N_19742,N_19625);
nand UO_772 (O_772,N_19662,N_19784);
xor UO_773 (O_773,N_19761,N_19889);
and UO_774 (O_774,N_19950,N_19700);
or UO_775 (O_775,N_19846,N_19937);
and UO_776 (O_776,N_19621,N_19780);
and UO_777 (O_777,N_19621,N_19663);
and UO_778 (O_778,N_19651,N_19803);
or UO_779 (O_779,N_19962,N_19947);
or UO_780 (O_780,N_19796,N_19725);
nand UO_781 (O_781,N_19826,N_19935);
nor UO_782 (O_782,N_19903,N_19846);
nand UO_783 (O_783,N_19706,N_19771);
xor UO_784 (O_784,N_19665,N_19913);
and UO_785 (O_785,N_19931,N_19755);
xnor UO_786 (O_786,N_19761,N_19890);
or UO_787 (O_787,N_19635,N_19843);
xnor UO_788 (O_788,N_19756,N_19602);
nand UO_789 (O_789,N_19960,N_19998);
and UO_790 (O_790,N_19643,N_19660);
and UO_791 (O_791,N_19783,N_19657);
and UO_792 (O_792,N_19928,N_19692);
nor UO_793 (O_793,N_19851,N_19693);
or UO_794 (O_794,N_19954,N_19980);
or UO_795 (O_795,N_19949,N_19708);
xor UO_796 (O_796,N_19716,N_19676);
and UO_797 (O_797,N_19753,N_19926);
xnor UO_798 (O_798,N_19971,N_19766);
nor UO_799 (O_799,N_19698,N_19889);
or UO_800 (O_800,N_19929,N_19788);
or UO_801 (O_801,N_19668,N_19943);
nand UO_802 (O_802,N_19973,N_19709);
nand UO_803 (O_803,N_19986,N_19810);
or UO_804 (O_804,N_19875,N_19696);
xor UO_805 (O_805,N_19834,N_19826);
and UO_806 (O_806,N_19690,N_19858);
nor UO_807 (O_807,N_19948,N_19688);
nor UO_808 (O_808,N_19656,N_19963);
nor UO_809 (O_809,N_19611,N_19997);
nand UO_810 (O_810,N_19617,N_19814);
or UO_811 (O_811,N_19755,N_19787);
nand UO_812 (O_812,N_19889,N_19729);
or UO_813 (O_813,N_19664,N_19925);
nor UO_814 (O_814,N_19792,N_19722);
nand UO_815 (O_815,N_19768,N_19991);
nor UO_816 (O_816,N_19618,N_19857);
nand UO_817 (O_817,N_19853,N_19642);
nor UO_818 (O_818,N_19705,N_19916);
nand UO_819 (O_819,N_19806,N_19723);
xor UO_820 (O_820,N_19650,N_19685);
nor UO_821 (O_821,N_19863,N_19762);
nand UO_822 (O_822,N_19794,N_19743);
and UO_823 (O_823,N_19613,N_19952);
nor UO_824 (O_824,N_19924,N_19963);
nor UO_825 (O_825,N_19955,N_19657);
nor UO_826 (O_826,N_19718,N_19614);
xnor UO_827 (O_827,N_19972,N_19822);
nand UO_828 (O_828,N_19867,N_19870);
nand UO_829 (O_829,N_19660,N_19861);
nand UO_830 (O_830,N_19653,N_19791);
nor UO_831 (O_831,N_19883,N_19895);
and UO_832 (O_832,N_19875,N_19777);
or UO_833 (O_833,N_19755,N_19656);
nand UO_834 (O_834,N_19736,N_19721);
xor UO_835 (O_835,N_19958,N_19748);
nor UO_836 (O_836,N_19689,N_19846);
and UO_837 (O_837,N_19991,N_19940);
and UO_838 (O_838,N_19797,N_19924);
nor UO_839 (O_839,N_19882,N_19961);
nor UO_840 (O_840,N_19805,N_19752);
nand UO_841 (O_841,N_19977,N_19966);
or UO_842 (O_842,N_19684,N_19658);
xnor UO_843 (O_843,N_19716,N_19991);
nand UO_844 (O_844,N_19935,N_19761);
nand UO_845 (O_845,N_19644,N_19676);
or UO_846 (O_846,N_19828,N_19820);
nand UO_847 (O_847,N_19960,N_19817);
and UO_848 (O_848,N_19682,N_19881);
xor UO_849 (O_849,N_19694,N_19890);
and UO_850 (O_850,N_19716,N_19835);
xnor UO_851 (O_851,N_19867,N_19837);
and UO_852 (O_852,N_19639,N_19833);
or UO_853 (O_853,N_19666,N_19795);
or UO_854 (O_854,N_19840,N_19934);
nand UO_855 (O_855,N_19728,N_19714);
nand UO_856 (O_856,N_19745,N_19672);
nand UO_857 (O_857,N_19629,N_19670);
nor UO_858 (O_858,N_19637,N_19811);
xor UO_859 (O_859,N_19678,N_19936);
nand UO_860 (O_860,N_19708,N_19682);
or UO_861 (O_861,N_19949,N_19606);
or UO_862 (O_862,N_19647,N_19739);
nor UO_863 (O_863,N_19959,N_19896);
nand UO_864 (O_864,N_19837,N_19759);
xnor UO_865 (O_865,N_19825,N_19951);
and UO_866 (O_866,N_19890,N_19825);
or UO_867 (O_867,N_19629,N_19902);
xor UO_868 (O_868,N_19629,N_19615);
or UO_869 (O_869,N_19953,N_19785);
nand UO_870 (O_870,N_19692,N_19911);
nor UO_871 (O_871,N_19861,N_19990);
and UO_872 (O_872,N_19907,N_19816);
xnor UO_873 (O_873,N_19960,N_19964);
or UO_874 (O_874,N_19988,N_19946);
or UO_875 (O_875,N_19666,N_19807);
or UO_876 (O_876,N_19805,N_19846);
and UO_877 (O_877,N_19911,N_19603);
nand UO_878 (O_878,N_19674,N_19883);
nand UO_879 (O_879,N_19966,N_19629);
and UO_880 (O_880,N_19934,N_19781);
or UO_881 (O_881,N_19712,N_19902);
or UO_882 (O_882,N_19786,N_19951);
nor UO_883 (O_883,N_19873,N_19629);
and UO_884 (O_884,N_19854,N_19741);
nand UO_885 (O_885,N_19991,N_19889);
and UO_886 (O_886,N_19995,N_19694);
nand UO_887 (O_887,N_19828,N_19744);
and UO_888 (O_888,N_19782,N_19953);
or UO_889 (O_889,N_19873,N_19608);
xnor UO_890 (O_890,N_19993,N_19895);
and UO_891 (O_891,N_19900,N_19635);
xnor UO_892 (O_892,N_19768,N_19746);
or UO_893 (O_893,N_19632,N_19751);
xnor UO_894 (O_894,N_19823,N_19799);
and UO_895 (O_895,N_19657,N_19651);
or UO_896 (O_896,N_19893,N_19837);
nor UO_897 (O_897,N_19921,N_19938);
nor UO_898 (O_898,N_19738,N_19843);
and UO_899 (O_899,N_19670,N_19808);
nand UO_900 (O_900,N_19781,N_19673);
and UO_901 (O_901,N_19898,N_19751);
and UO_902 (O_902,N_19862,N_19626);
nand UO_903 (O_903,N_19755,N_19942);
or UO_904 (O_904,N_19728,N_19640);
and UO_905 (O_905,N_19700,N_19782);
nand UO_906 (O_906,N_19800,N_19648);
xnor UO_907 (O_907,N_19941,N_19990);
nor UO_908 (O_908,N_19838,N_19639);
nor UO_909 (O_909,N_19688,N_19908);
and UO_910 (O_910,N_19964,N_19678);
nand UO_911 (O_911,N_19866,N_19833);
nor UO_912 (O_912,N_19674,N_19876);
and UO_913 (O_913,N_19803,N_19754);
nor UO_914 (O_914,N_19616,N_19773);
nand UO_915 (O_915,N_19739,N_19967);
nor UO_916 (O_916,N_19990,N_19922);
xnor UO_917 (O_917,N_19775,N_19921);
nor UO_918 (O_918,N_19977,N_19723);
nor UO_919 (O_919,N_19678,N_19843);
or UO_920 (O_920,N_19863,N_19916);
xnor UO_921 (O_921,N_19621,N_19814);
nand UO_922 (O_922,N_19936,N_19915);
nand UO_923 (O_923,N_19607,N_19986);
or UO_924 (O_924,N_19890,N_19787);
and UO_925 (O_925,N_19661,N_19735);
or UO_926 (O_926,N_19745,N_19960);
nand UO_927 (O_927,N_19650,N_19996);
nor UO_928 (O_928,N_19937,N_19862);
or UO_929 (O_929,N_19933,N_19706);
nor UO_930 (O_930,N_19941,N_19859);
nand UO_931 (O_931,N_19671,N_19828);
nor UO_932 (O_932,N_19614,N_19957);
nand UO_933 (O_933,N_19827,N_19619);
nor UO_934 (O_934,N_19794,N_19669);
and UO_935 (O_935,N_19679,N_19800);
nand UO_936 (O_936,N_19706,N_19602);
nand UO_937 (O_937,N_19751,N_19998);
xnor UO_938 (O_938,N_19649,N_19772);
nor UO_939 (O_939,N_19812,N_19937);
xor UO_940 (O_940,N_19673,N_19975);
and UO_941 (O_941,N_19943,N_19619);
nor UO_942 (O_942,N_19757,N_19951);
and UO_943 (O_943,N_19921,N_19741);
or UO_944 (O_944,N_19798,N_19673);
or UO_945 (O_945,N_19795,N_19783);
nor UO_946 (O_946,N_19725,N_19870);
nand UO_947 (O_947,N_19837,N_19820);
xor UO_948 (O_948,N_19744,N_19896);
xor UO_949 (O_949,N_19789,N_19981);
or UO_950 (O_950,N_19716,N_19600);
or UO_951 (O_951,N_19808,N_19692);
and UO_952 (O_952,N_19762,N_19934);
or UO_953 (O_953,N_19656,N_19934);
nor UO_954 (O_954,N_19831,N_19815);
xnor UO_955 (O_955,N_19632,N_19645);
xnor UO_956 (O_956,N_19979,N_19708);
or UO_957 (O_957,N_19854,N_19941);
and UO_958 (O_958,N_19666,N_19793);
and UO_959 (O_959,N_19822,N_19913);
or UO_960 (O_960,N_19614,N_19706);
xor UO_961 (O_961,N_19931,N_19997);
nand UO_962 (O_962,N_19887,N_19794);
xnor UO_963 (O_963,N_19880,N_19858);
xor UO_964 (O_964,N_19841,N_19600);
nand UO_965 (O_965,N_19926,N_19726);
nand UO_966 (O_966,N_19999,N_19731);
nor UO_967 (O_967,N_19979,N_19888);
and UO_968 (O_968,N_19962,N_19867);
and UO_969 (O_969,N_19709,N_19896);
nand UO_970 (O_970,N_19720,N_19740);
or UO_971 (O_971,N_19705,N_19895);
nand UO_972 (O_972,N_19838,N_19783);
and UO_973 (O_973,N_19893,N_19827);
nand UO_974 (O_974,N_19893,N_19800);
or UO_975 (O_975,N_19803,N_19626);
nand UO_976 (O_976,N_19807,N_19755);
xor UO_977 (O_977,N_19925,N_19873);
nor UO_978 (O_978,N_19982,N_19645);
or UO_979 (O_979,N_19944,N_19955);
nor UO_980 (O_980,N_19710,N_19793);
nor UO_981 (O_981,N_19671,N_19835);
and UO_982 (O_982,N_19810,N_19864);
nand UO_983 (O_983,N_19676,N_19650);
nand UO_984 (O_984,N_19702,N_19821);
and UO_985 (O_985,N_19877,N_19634);
or UO_986 (O_986,N_19836,N_19865);
xor UO_987 (O_987,N_19843,N_19962);
xor UO_988 (O_988,N_19617,N_19835);
and UO_989 (O_989,N_19625,N_19839);
xor UO_990 (O_990,N_19902,N_19974);
or UO_991 (O_991,N_19948,N_19606);
nand UO_992 (O_992,N_19791,N_19866);
and UO_993 (O_993,N_19903,N_19892);
xnor UO_994 (O_994,N_19990,N_19837);
nor UO_995 (O_995,N_19907,N_19832);
and UO_996 (O_996,N_19661,N_19786);
nor UO_997 (O_997,N_19931,N_19856);
xnor UO_998 (O_998,N_19895,N_19871);
and UO_999 (O_999,N_19894,N_19985);
and UO_1000 (O_1000,N_19919,N_19601);
nor UO_1001 (O_1001,N_19690,N_19602);
xnor UO_1002 (O_1002,N_19911,N_19972);
xor UO_1003 (O_1003,N_19852,N_19768);
nor UO_1004 (O_1004,N_19705,N_19719);
nor UO_1005 (O_1005,N_19721,N_19855);
and UO_1006 (O_1006,N_19874,N_19968);
or UO_1007 (O_1007,N_19820,N_19687);
xor UO_1008 (O_1008,N_19664,N_19862);
nor UO_1009 (O_1009,N_19928,N_19882);
and UO_1010 (O_1010,N_19723,N_19915);
and UO_1011 (O_1011,N_19677,N_19663);
xnor UO_1012 (O_1012,N_19637,N_19932);
nand UO_1013 (O_1013,N_19610,N_19936);
and UO_1014 (O_1014,N_19633,N_19830);
nand UO_1015 (O_1015,N_19843,N_19951);
or UO_1016 (O_1016,N_19639,N_19758);
or UO_1017 (O_1017,N_19707,N_19930);
xnor UO_1018 (O_1018,N_19652,N_19620);
nand UO_1019 (O_1019,N_19863,N_19833);
and UO_1020 (O_1020,N_19651,N_19721);
xnor UO_1021 (O_1021,N_19916,N_19937);
and UO_1022 (O_1022,N_19838,N_19739);
xor UO_1023 (O_1023,N_19992,N_19907);
nand UO_1024 (O_1024,N_19680,N_19659);
nor UO_1025 (O_1025,N_19819,N_19824);
or UO_1026 (O_1026,N_19757,N_19939);
nand UO_1027 (O_1027,N_19771,N_19863);
nand UO_1028 (O_1028,N_19640,N_19910);
and UO_1029 (O_1029,N_19608,N_19691);
nor UO_1030 (O_1030,N_19876,N_19610);
nand UO_1031 (O_1031,N_19719,N_19839);
and UO_1032 (O_1032,N_19748,N_19656);
nor UO_1033 (O_1033,N_19650,N_19704);
nand UO_1034 (O_1034,N_19801,N_19831);
nor UO_1035 (O_1035,N_19822,N_19995);
xor UO_1036 (O_1036,N_19949,N_19898);
nand UO_1037 (O_1037,N_19981,N_19761);
nand UO_1038 (O_1038,N_19696,N_19939);
xnor UO_1039 (O_1039,N_19753,N_19740);
xnor UO_1040 (O_1040,N_19612,N_19619);
nand UO_1041 (O_1041,N_19610,N_19608);
nor UO_1042 (O_1042,N_19780,N_19662);
nor UO_1043 (O_1043,N_19966,N_19673);
and UO_1044 (O_1044,N_19970,N_19905);
and UO_1045 (O_1045,N_19910,N_19877);
and UO_1046 (O_1046,N_19853,N_19653);
nand UO_1047 (O_1047,N_19970,N_19974);
nor UO_1048 (O_1048,N_19639,N_19829);
and UO_1049 (O_1049,N_19724,N_19883);
and UO_1050 (O_1050,N_19733,N_19830);
nand UO_1051 (O_1051,N_19921,N_19664);
or UO_1052 (O_1052,N_19718,N_19941);
nor UO_1053 (O_1053,N_19686,N_19633);
xnor UO_1054 (O_1054,N_19728,N_19804);
and UO_1055 (O_1055,N_19648,N_19634);
and UO_1056 (O_1056,N_19616,N_19666);
nand UO_1057 (O_1057,N_19776,N_19789);
and UO_1058 (O_1058,N_19677,N_19748);
nand UO_1059 (O_1059,N_19833,N_19874);
nand UO_1060 (O_1060,N_19989,N_19663);
or UO_1061 (O_1061,N_19722,N_19732);
or UO_1062 (O_1062,N_19784,N_19806);
and UO_1063 (O_1063,N_19947,N_19990);
nand UO_1064 (O_1064,N_19863,N_19700);
nor UO_1065 (O_1065,N_19838,N_19911);
nand UO_1066 (O_1066,N_19778,N_19865);
nor UO_1067 (O_1067,N_19614,N_19944);
and UO_1068 (O_1068,N_19614,N_19949);
xnor UO_1069 (O_1069,N_19818,N_19854);
nor UO_1070 (O_1070,N_19776,N_19699);
and UO_1071 (O_1071,N_19878,N_19939);
xnor UO_1072 (O_1072,N_19997,N_19943);
nor UO_1073 (O_1073,N_19996,N_19691);
nor UO_1074 (O_1074,N_19889,N_19748);
nand UO_1075 (O_1075,N_19994,N_19615);
or UO_1076 (O_1076,N_19864,N_19607);
nand UO_1077 (O_1077,N_19941,N_19934);
nand UO_1078 (O_1078,N_19628,N_19944);
or UO_1079 (O_1079,N_19808,N_19992);
xor UO_1080 (O_1080,N_19636,N_19649);
xnor UO_1081 (O_1081,N_19664,N_19837);
nor UO_1082 (O_1082,N_19878,N_19632);
xor UO_1083 (O_1083,N_19949,N_19695);
xnor UO_1084 (O_1084,N_19781,N_19870);
nand UO_1085 (O_1085,N_19616,N_19813);
nor UO_1086 (O_1086,N_19821,N_19996);
nor UO_1087 (O_1087,N_19698,N_19677);
nor UO_1088 (O_1088,N_19915,N_19706);
xor UO_1089 (O_1089,N_19638,N_19794);
or UO_1090 (O_1090,N_19941,N_19855);
and UO_1091 (O_1091,N_19693,N_19846);
nand UO_1092 (O_1092,N_19722,N_19949);
xnor UO_1093 (O_1093,N_19889,N_19728);
xor UO_1094 (O_1094,N_19694,N_19779);
nand UO_1095 (O_1095,N_19836,N_19771);
xor UO_1096 (O_1096,N_19957,N_19833);
nand UO_1097 (O_1097,N_19953,N_19857);
nor UO_1098 (O_1098,N_19962,N_19848);
and UO_1099 (O_1099,N_19807,N_19905);
nand UO_1100 (O_1100,N_19633,N_19770);
or UO_1101 (O_1101,N_19665,N_19945);
nor UO_1102 (O_1102,N_19784,N_19745);
and UO_1103 (O_1103,N_19682,N_19621);
nand UO_1104 (O_1104,N_19835,N_19654);
nand UO_1105 (O_1105,N_19671,N_19767);
nor UO_1106 (O_1106,N_19806,N_19665);
and UO_1107 (O_1107,N_19786,N_19889);
xnor UO_1108 (O_1108,N_19911,N_19999);
and UO_1109 (O_1109,N_19942,N_19938);
or UO_1110 (O_1110,N_19901,N_19706);
and UO_1111 (O_1111,N_19773,N_19990);
nand UO_1112 (O_1112,N_19958,N_19979);
nor UO_1113 (O_1113,N_19842,N_19912);
xor UO_1114 (O_1114,N_19794,N_19666);
and UO_1115 (O_1115,N_19869,N_19924);
xor UO_1116 (O_1116,N_19955,N_19732);
or UO_1117 (O_1117,N_19728,N_19680);
or UO_1118 (O_1118,N_19890,N_19755);
nand UO_1119 (O_1119,N_19933,N_19707);
xnor UO_1120 (O_1120,N_19755,N_19615);
and UO_1121 (O_1121,N_19756,N_19852);
xnor UO_1122 (O_1122,N_19935,N_19626);
and UO_1123 (O_1123,N_19868,N_19990);
nand UO_1124 (O_1124,N_19854,N_19942);
xnor UO_1125 (O_1125,N_19623,N_19823);
or UO_1126 (O_1126,N_19776,N_19769);
or UO_1127 (O_1127,N_19867,N_19701);
or UO_1128 (O_1128,N_19864,N_19619);
xor UO_1129 (O_1129,N_19712,N_19916);
xnor UO_1130 (O_1130,N_19836,N_19692);
or UO_1131 (O_1131,N_19901,N_19793);
or UO_1132 (O_1132,N_19949,N_19800);
xnor UO_1133 (O_1133,N_19809,N_19923);
nor UO_1134 (O_1134,N_19713,N_19781);
or UO_1135 (O_1135,N_19792,N_19600);
nor UO_1136 (O_1136,N_19956,N_19632);
and UO_1137 (O_1137,N_19672,N_19603);
nor UO_1138 (O_1138,N_19755,N_19719);
nor UO_1139 (O_1139,N_19834,N_19636);
xor UO_1140 (O_1140,N_19758,N_19881);
xor UO_1141 (O_1141,N_19780,N_19783);
nand UO_1142 (O_1142,N_19816,N_19949);
nor UO_1143 (O_1143,N_19773,N_19818);
xnor UO_1144 (O_1144,N_19690,N_19748);
nand UO_1145 (O_1145,N_19724,N_19923);
or UO_1146 (O_1146,N_19767,N_19678);
nand UO_1147 (O_1147,N_19799,N_19953);
nand UO_1148 (O_1148,N_19691,N_19894);
and UO_1149 (O_1149,N_19833,N_19934);
xnor UO_1150 (O_1150,N_19631,N_19628);
nand UO_1151 (O_1151,N_19726,N_19889);
xor UO_1152 (O_1152,N_19606,N_19852);
nor UO_1153 (O_1153,N_19851,N_19941);
and UO_1154 (O_1154,N_19829,N_19790);
xor UO_1155 (O_1155,N_19967,N_19969);
xor UO_1156 (O_1156,N_19693,N_19768);
and UO_1157 (O_1157,N_19689,N_19812);
nor UO_1158 (O_1158,N_19818,N_19748);
nor UO_1159 (O_1159,N_19753,N_19663);
or UO_1160 (O_1160,N_19755,N_19913);
and UO_1161 (O_1161,N_19647,N_19915);
or UO_1162 (O_1162,N_19789,N_19982);
xor UO_1163 (O_1163,N_19672,N_19664);
or UO_1164 (O_1164,N_19911,N_19987);
nor UO_1165 (O_1165,N_19975,N_19631);
nor UO_1166 (O_1166,N_19753,N_19944);
and UO_1167 (O_1167,N_19800,N_19677);
nor UO_1168 (O_1168,N_19862,N_19728);
nor UO_1169 (O_1169,N_19933,N_19616);
or UO_1170 (O_1170,N_19871,N_19958);
nand UO_1171 (O_1171,N_19899,N_19867);
nor UO_1172 (O_1172,N_19858,N_19721);
nor UO_1173 (O_1173,N_19904,N_19619);
nor UO_1174 (O_1174,N_19600,N_19820);
nand UO_1175 (O_1175,N_19913,N_19657);
xnor UO_1176 (O_1176,N_19980,N_19870);
nand UO_1177 (O_1177,N_19762,N_19604);
or UO_1178 (O_1178,N_19701,N_19769);
or UO_1179 (O_1179,N_19741,N_19759);
nor UO_1180 (O_1180,N_19631,N_19853);
or UO_1181 (O_1181,N_19953,N_19716);
nor UO_1182 (O_1182,N_19997,N_19667);
and UO_1183 (O_1183,N_19807,N_19835);
nand UO_1184 (O_1184,N_19771,N_19839);
and UO_1185 (O_1185,N_19955,N_19835);
xor UO_1186 (O_1186,N_19994,N_19973);
nand UO_1187 (O_1187,N_19781,N_19922);
nor UO_1188 (O_1188,N_19810,N_19894);
and UO_1189 (O_1189,N_19827,N_19778);
xor UO_1190 (O_1190,N_19932,N_19922);
and UO_1191 (O_1191,N_19838,N_19649);
nor UO_1192 (O_1192,N_19674,N_19832);
xor UO_1193 (O_1193,N_19791,N_19608);
and UO_1194 (O_1194,N_19740,N_19653);
xor UO_1195 (O_1195,N_19881,N_19715);
nor UO_1196 (O_1196,N_19628,N_19766);
xor UO_1197 (O_1197,N_19960,N_19851);
and UO_1198 (O_1198,N_19874,N_19919);
and UO_1199 (O_1199,N_19872,N_19741);
xor UO_1200 (O_1200,N_19808,N_19634);
nand UO_1201 (O_1201,N_19993,N_19719);
or UO_1202 (O_1202,N_19717,N_19662);
and UO_1203 (O_1203,N_19929,N_19734);
nor UO_1204 (O_1204,N_19779,N_19648);
or UO_1205 (O_1205,N_19943,N_19766);
xor UO_1206 (O_1206,N_19980,N_19726);
or UO_1207 (O_1207,N_19870,N_19878);
nor UO_1208 (O_1208,N_19881,N_19660);
nand UO_1209 (O_1209,N_19661,N_19692);
or UO_1210 (O_1210,N_19854,N_19654);
nand UO_1211 (O_1211,N_19861,N_19686);
nor UO_1212 (O_1212,N_19765,N_19741);
or UO_1213 (O_1213,N_19796,N_19789);
and UO_1214 (O_1214,N_19699,N_19677);
xor UO_1215 (O_1215,N_19684,N_19722);
nand UO_1216 (O_1216,N_19939,N_19958);
nand UO_1217 (O_1217,N_19997,N_19916);
nor UO_1218 (O_1218,N_19879,N_19967);
nand UO_1219 (O_1219,N_19615,N_19988);
xor UO_1220 (O_1220,N_19831,N_19764);
or UO_1221 (O_1221,N_19795,N_19733);
nor UO_1222 (O_1222,N_19801,N_19849);
nand UO_1223 (O_1223,N_19774,N_19743);
or UO_1224 (O_1224,N_19639,N_19720);
and UO_1225 (O_1225,N_19772,N_19894);
and UO_1226 (O_1226,N_19603,N_19635);
or UO_1227 (O_1227,N_19859,N_19895);
or UO_1228 (O_1228,N_19920,N_19763);
and UO_1229 (O_1229,N_19786,N_19944);
xor UO_1230 (O_1230,N_19916,N_19606);
nor UO_1231 (O_1231,N_19605,N_19751);
nand UO_1232 (O_1232,N_19986,N_19703);
nand UO_1233 (O_1233,N_19703,N_19952);
nor UO_1234 (O_1234,N_19914,N_19735);
xor UO_1235 (O_1235,N_19645,N_19644);
and UO_1236 (O_1236,N_19920,N_19903);
or UO_1237 (O_1237,N_19806,N_19953);
and UO_1238 (O_1238,N_19729,N_19988);
or UO_1239 (O_1239,N_19948,N_19682);
xor UO_1240 (O_1240,N_19996,N_19870);
xor UO_1241 (O_1241,N_19908,N_19898);
nor UO_1242 (O_1242,N_19905,N_19986);
nor UO_1243 (O_1243,N_19636,N_19959);
xor UO_1244 (O_1244,N_19728,N_19771);
and UO_1245 (O_1245,N_19633,N_19970);
nor UO_1246 (O_1246,N_19668,N_19810);
nand UO_1247 (O_1247,N_19681,N_19866);
nand UO_1248 (O_1248,N_19961,N_19743);
or UO_1249 (O_1249,N_19738,N_19628);
nor UO_1250 (O_1250,N_19864,N_19645);
xor UO_1251 (O_1251,N_19960,N_19988);
or UO_1252 (O_1252,N_19982,N_19654);
nor UO_1253 (O_1253,N_19733,N_19820);
or UO_1254 (O_1254,N_19729,N_19761);
xnor UO_1255 (O_1255,N_19894,N_19632);
nor UO_1256 (O_1256,N_19664,N_19914);
xnor UO_1257 (O_1257,N_19795,N_19707);
and UO_1258 (O_1258,N_19727,N_19895);
xor UO_1259 (O_1259,N_19821,N_19689);
xor UO_1260 (O_1260,N_19902,N_19975);
nor UO_1261 (O_1261,N_19857,N_19943);
and UO_1262 (O_1262,N_19722,N_19822);
nor UO_1263 (O_1263,N_19654,N_19740);
nor UO_1264 (O_1264,N_19859,N_19877);
xnor UO_1265 (O_1265,N_19848,N_19738);
and UO_1266 (O_1266,N_19907,N_19711);
and UO_1267 (O_1267,N_19833,N_19670);
xnor UO_1268 (O_1268,N_19728,N_19886);
nand UO_1269 (O_1269,N_19851,N_19895);
and UO_1270 (O_1270,N_19767,N_19605);
nand UO_1271 (O_1271,N_19864,N_19776);
or UO_1272 (O_1272,N_19741,N_19774);
nand UO_1273 (O_1273,N_19849,N_19653);
and UO_1274 (O_1274,N_19625,N_19849);
or UO_1275 (O_1275,N_19605,N_19713);
or UO_1276 (O_1276,N_19812,N_19982);
xnor UO_1277 (O_1277,N_19608,N_19827);
xnor UO_1278 (O_1278,N_19769,N_19936);
and UO_1279 (O_1279,N_19615,N_19834);
xor UO_1280 (O_1280,N_19754,N_19893);
nand UO_1281 (O_1281,N_19995,N_19702);
or UO_1282 (O_1282,N_19823,N_19889);
nor UO_1283 (O_1283,N_19771,N_19740);
xnor UO_1284 (O_1284,N_19899,N_19883);
and UO_1285 (O_1285,N_19898,N_19800);
or UO_1286 (O_1286,N_19828,N_19803);
nor UO_1287 (O_1287,N_19790,N_19635);
nand UO_1288 (O_1288,N_19638,N_19745);
and UO_1289 (O_1289,N_19600,N_19917);
nor UO_1290 (O_1290,N_19607,N_19869);
xor UO_1291 (O_1291,N_19731,N_19646);
xnor UO_1292 (O_1292,N_19769,N_19850);
or UO_1293 (O_1293,N_19796,N_19998);
nand UO_1294 (O_1294,N_19992,N_19918);
nand UO_1295 (O_1295,N_19821,N_19822);
or UO_1296 (O_1296,N_19662,N_19644);
xnor UO_1297 (O_1297,N_19951,N_19731);
or UO_1298 (O_1298,N_19715,N_19856);
and UO_1299 (O_1299,N_19872,N_19702);
and UO_1300 (O_1300,N_19657,N_19655);
nand UO_1301 (O_1301,N_19672,N_19678);
nand UO_1302 (O_1302,N_19954,N_19616);
nand UO_1303 (O_1303,N_19978,N_19991);
or UO_1304 (O_1304,N_19826,N_19663);
and UO_1305 (O_1305,N_19622,N_19666);
or UO_1306 (O_1306,N_19830,N_19625);
or UO_1307 (O_1307,N_19691,N_19727);
xnor UO_1308 (O_1308,N_19888,N_19700);
nor UO_1309 (O_1309,N_19774,N_19786);
nor UO_1310 (O_1310,N_19609,N_19818);
or UO_1311 (O_1311,N_19968,N_19683);
nand UO_1312 (O_1312,N_19950,N_19711);
nor UO_1313 (O_1313,N_19789,N_19605);
and UO_1314 (O_1314,N_19626,N_19899);
nand UO_1315 (O_1315,N_19790,N_19672);
xnor UO_1316 (O_1316,N_19600,N_19913);
xnor UO_1317 (O_1317,N_19750,N_19886);
or UO_1318 (O_1318,N_19837,N_19941);
and UO_1319 (O_1319,N_19952,N_19990);
or UO_1320 (O_1320,N_19886,N_19704);
and UO_1321 (O_1321,N_19717,N_19972);
nand UO_1322 (O_1322,N_19742,N_19944);
or UO_1323 (O_1323,N_19647,N_19948);
nor UO_1324 (O_1324,N_19745,N_19631);
nor UO_1325 (O_1325,N_19775,N_19668);
and UO_1326 (O_1326,N_19838,N_19721);
nand UO_1327 (O_1327,N_19683,N_19828);
and UO_1328 (O_1328,N_19854,N_19618);
xnor UO_1329 (O_1329,N_19732,N_19945);
and UO_1330 (O_1330,N_19681,N_19751);
nor UO_1331 (O_1331,N_19908,N_19737);
and UO_1332 (O_1332,N_19778,N_19714);
or UO_1333 (O_1333,N_19943,N_19659);
or UO_1334 (O_1334,N_19659,N_19636);
nor UO_1335 (O_1335,N_19907,N_19959);
xor UO_1336 (O_1336,N_19894,N_19788);
nand UO_1337 (O_1337,N_19663,N_19911);
nand UO_1338 (O_1338,N_19690,N_19993);
and UO_1339 (O_1339,N_19997,N_19879);
and UO_1340 (O_1340,N_19978,N_19807);
nand UO_1341 (O_1341,N_19848,N_19970);
xor UO_1342 (O_1342,N_19763,N_19801);
nor UO_1343 (O_1343,N_19919,N_19643);
xnor UO_1344 (O_1344,N_19739,N_19778);
nor UO_1345 (O_1345,N_19730,N_19999);
and UO_1346 (O_1346,N_19931,N_19754);
and UO_1347 (O_1347,N_19784,N_19630);
nor UO_1348 (O_1348,N_19657,N_19642);
or UO_1349 (O_1349,N_19807,N_19632);
xor UO_1350 (O_1350,N_19810,N_19853);
nor UO_1351 (O_1351,N_19887,N_19650);
xnor UO_1352 (O_1352,N_19635,N_19916);
and UO_1353 (O_1353,N_19689,N_19770);
nor UO_1354 (O_1354,N_19855,N_19853);
or UO_1355 (O_1355,N_19672,N_19792);
or UO_1356 (O_1356,N_19900,N_19984);
or UO_1357 (O_1357,N_19769,N_19851);
xor UO_1358 (O_1358,N_19645,N_19921);
xor UO_1359 (O_1359,N_19871,N_19733);
nor UO_1360 (O_1360,N_19694,N_19868);
nor UO_1361 (O_1361,N_19956,N_19729);
xnor UO_1362 (O_1362,N_19828,N_19869);
and UO_1363 (O_1363,N_19917,N_19976);
nor UO_1364 (O_1364,N_19725,N_19747);
xnor UO_1365 (O_1365,N_19627,N_19704);
and UO_1366 (O_1366,N_19974,N_19773);
nor UO_1367 (O_1367,N_19811,N_19975);
or UO_1368 (O_1368,N_19857,N_19913);
nand UO_1369 (O_1369,N_19698,N_19636);
nor UO_1370 (O_1370,N_19962,N_19839);
or UO_1371 (O_1371,N_19600,N_19784);
nor UO_1372 (O_1372,N_19680,N_19891);
nand UO_1373 (O_1373,N_19959,N_19951);
xor UO_1374 (O_1374,N_19968,N_19777);
xor UO_1375 (O_1375,N_19938,N_19712);
or UO_1376 (O_1376,N_19602,N_19996);
and UO_1377 (O_1377,N_19811,N_19735);
or UO_1378 (O_1378,N_19833,N_19826);
and UO_1379 (O_1379,N_19700,N_19832);
and UO_1380 (O_1380,N_19934,N_19987);
and UO_1381 (O_1381,N_19849,N_19924);
xor UO_1382 (O_1382,N_19899,N_19737);
nor UO_1383 (O_1383,N_19752,N_19628);
nand UO_1384 (O_1384,N_19676,N_19704);
and UO_1385 (O_1385,N_19638,N_19836);
and UO_1386 (O_1386,N_19760,N_19997);
xnor UO_1387 (O_1387,N_19662,N_19692);
nor UO_1388 (O_1388,N_19712,N_19785);
nor UO_1389 (O_1389,N_19777,N_19770);
xnor UO_1390 (O_1390,N_19916,N_19836);
nand UO_1391 (O_1391,N_19695,N_19809);
and UO_1392 (O_1392,N_19956,N_19761);
or UO_1393 (O_1393,N_19896,N_19979);
or UO_1394 (O_1394,N_19776,N_19615);
nor UO_1395 (O_1395,N_19690,N_19983);
nor UO_1396 (O_1396,N_19864,N_19838);
xnor UO_1397 (O_1397,N_19971,N_19817);
and UO_1398 (O_1398,N_19880,N_19840);
xor UO_1399 (O_1399,N_19775,N_19875);
nor UO_1400 (O_1400,N_19786,N_19658);
nand UO_1401 (O_1401,N_19888,N_19886);
xnor UO_1402 (O_1402,N_19825,N_19678);
and UO_1403 (O_1403,N_19922,N_19903);
nand UO_1404 (O_1404,N_19786,N_19645);
or UO_1405 (O_1405,N_19941,N_19888);
or UO_1406 (O_1406,N_19695,N_19703);
nor UO_1407 (O_1407,N_19773,N_19902);
nor UO_1408 (O_1408,N_19782,N_19875);
xor UO_1409 (O_1409,N_19992,N_19908);
nand UO_1410 (O_1410,N_19863,N_19819);
and UO_1411 (O_1411,N_19627,N_19675);
xor UO_1412 (O_1412,N_19768,N_19774);
nand UO_1413 (O_1413,N_19623,N_19994);
or UO_1414 (O_1414,N_19671,N_19928);
xnor UO_1415 (O_1415,N_19995,N_19893);
nand UO_1416 (O_1416,N_19895,N_19932);
nor UO_1417 (O_1417,N_19721,N_19674);
nand UO_1418 (O_1418,N_19988,N_19694);
nor UO_1419 (O_1419,N_19829,N_19826);
nor UO_1420 (O_1420,N_19904,N_19901);
xor UO_1421 (O_1421,N_19720,N_19653);
nor UO_1422 (O_1422,N_19988,N_19897);
nand UO_1423 (O_1423,N_19941,N_19639);
and UO_1424 (O_1424,N_19665,N_19990);
nand UO_1425 (O_1425,N_19718,N_19909);
xnor UO_1426 (O_1426,N_19844,N_19686);
nand UO_1427 (O_1427,N_19916,N_19760);
nand UO_1428 (O_1428,N_19836,N_19768);
xor UO_1429 (O_1429,N_19640,N_19922);
or UO_1430 (O_1430,N_19980,N_19806);
nand UO_1431 (O_1431,N_19856,N_19843);
nor UO_1432 (O_1432,N_19628,N_19984);
and UO_1433 (O_1433,N_19754,N_19825);
nand UO_1434 (O_1434,N_19863,N_19942);
nor UO_1435 (O_1435,N_19648,N_19871);
and UO_1436 (O_1436,N_19890,N_19956);
xnor UO_1437 (O_1437,N_19827,N_19888);
xor UO_1438 (O_1438,N_19737,N_19617);
nand UO_1439 (O_1439,N_19618,N_19966);
or UO_1440 (O_1440,N_19670,N_19718);
or UO_1441 (O_1441,N_19614,N_19714);
and UO_1442 (O_1442,N_19859,N_19834);
nand UO_1443 (O_1443,N_19642,N_19622);
nand UO_1444 (O_1444,N_19980,N_19993);
xnor UO_1445 (O_1445,N_19893,N_19808);
and UO_1446 (O_1446,N_19660,N_19888);
nor UO_1447 (O_1447,N_19705,N_19875);
and UO_1448 (O_1448,N_19936,N_19889);
or UO_1449 (O_1449,N_19693,N_19964);
xnor UO_1450 (O_1450,N_19845,N_19806);
and UO_1451 (O_1451,N_19690,N_19873);
xnor UO_1452 (O_1452,N_19904,N_19918);
xnor UO_1453 (O_1453,N_19649,N_19617);
xor UO_1454 (O_1454,N_19929,N_19922);
xor UO_1455 (O_1455,N_19731,N_19958);
nor UO_1456 (O_1456,N_19678,N_19792);
and UO_1457 (O_1457,N_19706,N_19696);
or UO_1458 (O_1458,N_19976,N_19652);
or UO_1459 (O_1459,N_19823,N_19982);
or UO_1460 (O_1460,N_19927,N_19786);
nand UO_1461 (O_1461,N_19768,N_19665);
xor UO_1462 (O_1462,N_19923,N_19818);
or UO_1463 (O_1463,N_19881,N_19651);
xnor UO_1464 (O_1464,N_19842,N_19604);
xor UO_1465 (O_1465,N_19653,N_19631);
or UO_1466 (O_1466,N_19885,N_19695);
nand UO_1467 (O_1467,N_19985,N_19729);
nand UO_1468 (O_1468,N_19859,N_19646);
or UO_1469 (O_1469,N_19799,N_19846);
or UO_1470 (O_1470,N_19818,N_19741);
nand UO_1471 (O_1471,N_19649,N_19885);
nor UO_1472 (O_1472,N_19869,N_19695);
nor UO_1473 (O_1473,N_19633,N_19881);
and UO_1474 (O_1474,N_19862,N_19676);
nand UO_1475 (O_1475,N_19759,N_19896);
xor UO_1476 (O_1476,N_19922,N_19780);
nor UO_1477 (O_1477,N_19853,N_19658);
nand UO_1478 (O_1478,N_19924,N_19743);
xnor UO_1479 (O_1479,N_19918,N_19702);
or UO_1480 (O_1480,N_19821,N_19927);
or UO_1481 (O_1481,N_19728,N_19846);
nor UO_1482 (O_1482,N_19819,N_19993);
or UO_1483 (O_1483,N_19914,N_19953);
nor UO_1484 (O_1484,N_19869,N_19839);
and UO_1485 (O_1485,N_19764,N_19887);
and UO_1486 (O_1486,N_19744,N_19873);
or UO_1487 (O_1487,N_19745,N_19924);
and UO_1488 (O_1488,N_19678,N_19699);
nand UO_1489 (O_1489,N_19926,N_19972);
and UO_1490 (O_1490,N_19858,N_19661);
xnor UO_1491 (O_1491,N_19905,N_19922);
or UO_1492 (O_1492,N_19625,N_19806);
or UO_1493 (O_1493,N_19784,N_19826);
nand UO_1494 (O_1494,N_19919,N_19636);
and UO_1495 (O_1495,N_19899,N_19768);
nand UO_1496 (O_1496,N_19605,N_19775);
nand UO_1497 (O_1497,N_19628,N_19662);
xnor UO_1498 (O_1498,N_19830,N_19642);
or UO_1499 (O_1499,N_19700,N_19601);
nand UO_1500 (O_1500,N_19669,N_19833);
nand UO_1501 (O_1501,N_19677,N_19916);
xnor UO_1502 (O_1502,N_19630,N_19899);
and UO_1503 (O_1503,N_19994,N_19838);
xnor UO_1504 (O_1504,N_19827,N_19649);
nor UO_1505 (O_1505,N_19779,N_19924);
nor UO_1506 (O_1506,N_19695,N_19828);
and UO_1507 (O_1507,N_19612,N_19667);
or UO_1508 (O_1508,N_19801,N_19663);
xnor UO_1509 (O_1509,N_19692,N_19801);
or UO_1510 (O_1510,N_19674,N_19850);
and UO_1511 (O_1511,N_19786,N_19699);
nor UO_1512 (O_1512,N_19755,N_19982);
nor UO_1513 (O_1513,N_19794,N_19832);
and UO_1514 (O_1514,N_19831,N_19716);
nand UO_1515 (O_1515,N_19994,N_19813);
or UO_1516 (O_1516,N_19700,N_19689);
xor UO_1517 (O_1517,N_19706,N_19946);
or UO_1518 (O_1518,N_19719,N_19669);
nand UO_1519 (O_1519,N_19619,N_19837);
nand UO_1520 (O_1520,N_19741,N_19981);
and UO_1521 (O_1521,N_19811,N_19956);
and UO_1522 (O_1522,N_19672,N_19674);
xnor UO_1523 (O_1523,N_19826,N_19848);
xor UO_1524 (O_1524,N_19763,N_19653);
and UO_1525 (O_1525,N_19633,N_19853);
nor UO_1526 (O_1526,N_19694,N_19792);
xor UO_1527 (O_1527,N_19966,N_19693);
or UO_1528 (O_1528,N_19798,N_19893);
nor UO_1529 (O_1529,N_19807,N_19684);
nand UO_1530 (O_1530,N_19992,N_19626);
nor UO_1531 (O_1531,N_19812,N_19833);
nor UO_1532 (O_1532,N_19890,N_19911);
or UO_1533 (O_1533,N_19986,N_19741);
and UO_1534 (O_1534,N_19934,N_19684);
xor UO_1535 (O_1535,N_19689,N_19681);
nor UO_1536 (O_1536,N_19689,N_19711);
xnor UO_1537 (O_1537,N_19706,N_19966);
nand UO_1538 (O_1538,N_19658,N_19690);
nand UO_1539 (O_1539,N_19629,N_19996);
or UO_1540 (O_1540,N_19785,N_19949);
xor UO_1541 (O_1541,N_19623,N_19657);
or UO_1542 (O_1542,N_19906,N_19979);
or UO_1543 (O_1543,N_19627,N_19736);
nand UO_1544 (O_1544,N_19945,N_19798);
nand UO_1545 (O_1545,N_19880,N_19680);
or UO_1546 (O_1546,N_19892,N_19810);
nand UO_1547 (O_1547,N_19745,N_19618);
or UO_1548 (O_1548,N_19623,N_19744);
xnor UO_1549 (O_1549,N_19866,N_19836);
xor UO_1550 (O_1550,N_19890,N_19865);
and UO_1551 (O_1551,N_19781,N_19815);
nand UO_1552 (O_1552,N_19841,N_19656);
nand UO_1553 (O_1553,N_19608,N_19881);
nand UO_1554 (O_1554,N_19697,N_19868);
nor UO_1555 (O_1555,N_19735,N_19803);
nand UO_1556 (O_1556,N_19758,N_19682);
and UO_1557 (O_1557,N_19891,N_19931);
and UO_1558 (O_1558,N_19962,N_19943);
or UO_1559 (O_1559,N_19752,N_19806);
nand UO_1560 (O_1560,N_19629,N_19690);
or UO_1561 (O_1561,N_19787,N_19875);
or UO_1562 (O_1562,N_19838,N_19922);
or UO_1563 (O_1563,N_19714,N_19634);
nor UO_1564 (O_1564,N_19824,N_19710);
or UO_1565 (O_1565,N_19976,N_19947);
nand UO_1566 (O_1566,N_19663,N_19942);
and UO_1567 (O_1567,N_19734,N_19825);
nor UO_1568 (O_1568,N_19820,N_19860);
and UO_1569 (O_1569,N_19857,N_19640);
xnor UO_1570 (O_1570,N_19672,N_19904);
and UO_1571 (O_1571,N_19608,N_19990);
and UO_1572 (O_1572,N_19929,N_19964);
nor UO_1573 (O_1573,N_19793,N_19997);
and UO_1574 (O_1574,N_19635,N_19690);
and UO_1575 (O_1575,N_19672,N_19673);
xnor UO_1576 (O_1576,N_19894,N_19908);
nand UO_1577 (O_1577,N_19718,N_19729);
and UO_1578 (O_1578,N_19942,N_19643);
nand UO_1579 (O_1579,N_19918,N_19920);
nor UO_1580 (O_1580,N_19867,N_19691);
or UO_1581 (O_1581,N_19886,N_19967);
and UO_1582 (O_1582,N_19814,N_19907);
and UO_1583 (O_1583,N_19906,N_19722);
and UO_1584 (O_1584,N_19785,N_19834);
nand UO_1585 (O_1585,N_19907,N_19831);
or UO_1586 (O_1586,N_19951,N_19619);
nor UO_1587 (O_1587,N_19929,N_19888);
nand UO_1588 (O_1588,N_19748,N_19793);
nand UO_1589 (O_1589,N_19608,N_19675);
nand UO_1590 (O_1590,N_19624,N_19950);
nor UO_1591 (O_1591,N_19898,N_19940);
and UO_1592 (O_1592,N_19864,N_19769);
nor UO_1593 (O_1593,N_19731,N_19667);
xor UO_1594 (O_1594,N_19652,N_19777);
xor UO_1595 (O_1595,N_19647,N_19691);
nor UO_1596 (O_1596,N_19818,N_19866);
nand UO_1597 (O_1597,N_19601,N_19782);
nand UO_1598 (O_1598,N_19857,N_19926);
nor UO_1599 (O_1599,N_19727,N_19613);
and UO_1600 (O_1600,N_19652,N_19647);
or UO_1601 (O_1601,N_19826,N_19684);
nand UO_1602 (O_1602,N_19859,N_19891);
or UO_1603 (O_1603,N_19808,N_19745);
nand UO_1604 (O_1604,N_19862,N_19706);
nand UO_1605 (O_1605,N_19755,N_19920);
nand UO_1606 (O_1606,N_19836,N_19917);
or UO_1607 (O_1607,N_19706,N_19923);
or UO_1608 (O_1608,N_19757,N_19821);
xnor UO_1609 (O_1609,N_19782,N_19872);
xor UO_1610 (O_1610,N_19816,N_19715);
xnor UO_1611 (O_1611,N_19745,N_19763);
nor UO_1612 (O_1612,N_19778,N_19684);
and UO_1613 (O_1613,N_19896,N_19892);
or UO_1614 (O_1614,N_19640,N_19931);
or UO_1615 (O_1615,N_19761,N_19893);
and UO_1616 (O_1616,N_19655,N_19790);
nand UO_1617 (O_1617,N_19888,N_19920);
nor UO_1618 (O_1618,N_19886,N_19995);
nand UO_1619 (O_1619,N_19888,N_19862);
xor UO_1620 (O_1620,N_19710,N_19860);
or UO_1621 (O_1621,N_19633,N_19672);
nor UO_1622 (O_1622,N_19762,N_19643);
xor UO_1623 (O_1623,N_19786,N_19798);
xnor UO_1624 (O_1624,N_19849,N_19812);
xnor UO_1625 (O_1625,N_19831,N_19982);
or UO_1626 (O_1626,N_19849,N_19629);
nand UO_1627 (O_1627,N_19990,N_19739);
or UO_1628 (O_1628,N_19604,N_19642);
nand UO_1629 (O_1629,N_19675,N_19720);
and UO_1630 (O_1630,N_19705,N_19884);
nand UO_1631 (O_1631,N_19685,N_19680);
nand UO_1632 (O_1632,N_19730,N_19918);
nor UO_1633 (O_1633,N_19889,N_19617);
xnor UO_1634 (O_1634,N_19809,N_19788);
or UO_1635 (O_1635,N_19609,N_19995);
nor UO_1636 (O_1636,N_19947,N_19847);
nor UO_1637 (O_1637,N_19742,N_19799);
and UO_1638 (O_1638,N_19701,N_19610);
xor UO_1639 (O_1639,N_19640,N_19984);
or UO_1640 (O_1640,N_19844,N_19850);
or UO_1641 (O_1641,N_19976,N_19770);
or UO_1642 (O_1642,N_19864,N_19835);
nor UO_1643 (O_1643,N_19806,N_19991);
xor UO_1644 (O_1644,N_19680,N_19960);
nand UO_1645 (O_1645,N_19883,N_19882);
xor UO_1646 (O_1646,N_19651,N_19772);
and UO_1647 (O_1647,N_19703,N_19957);
nand UO_1648 (O_1648,N_19731,N_19712);
or UO_1649 (O_1649,N_19742,N_19621);
and UO_1650 (O_1650,N_19775,N_19617);
xor UO_1651 (O_1651,N_19935,N_19733);
and UO_1652 (O_1652,N_19703,N_19837);
or UO_1653 (O_1653,N_19900,N_19889);
nand UO_1654 (O_1654,N_19711,N_19660);
or UO_1655 (O_1655,N_19617,N_19877);
xnor UO_1656 (O_1656,N_19818,N_19674);
and UO_1657 (O_1657,N_19971,N_19750);
and UO_1658 (O_1658,N_19903,N_19857);
or UO_1659 (O_1659,N_19707,N_19663);
or UO_1660 (O_1660,N_19679,N_19752);
nand UO_1661 (O_1661,N_19607,N_19712);
xor UO_1662 (O_1662,N_19912,N_19784);
or UO_1663 (O_1663,N_19933,N_19612);
or UO_1664 (O_1664,N_19806,N_19786);
xor UO_1665 (O_1665,N_19609,N_19972);
and UO_1666 (O_1666,N_19875,N_19716);
nor UO_1667 (O_1667,N_19940,N_19684);
xor UO_1668 (O_1668,N_19979,N_19678);
and UO_1669 (O_1669,N_19861,N_19747);
and UO_1670 (O_1670,N_19872,N_19960);
nor UO_1671 (O_1671,N_19827,N_19845);
and UO_1672 (O_1672,N_19621,N_19734);
nor UO_1673 (O_1673,N_19861,N_19875);
xor UO_1674 (O_1674,N_19831,N_19798);
nor UO_1675 (O_1675,N_19733,N_19875);
nor UO_1676 (O_1676,N_19728,N_19832);
nand UO_1677 (O_1677,N_19870,N_19967);
nand UO_1678 (O_1678,N_19601,N_19958);
and UO_1679 (O_1679,N_19941,N_19606);
nand UO_1680 (O_1680,N_19743,N_19725);
nand UO_1681 (O_1681,N_19783,N_19901);
nand UO_1682 (O_1682,N_19990,N_19644);
nand UO_1683 (O_1683,N_19819,N_19611);
or UO_1684 (O_1684,N_19624,N_19662);
or UO_1685 (O_1685,N_19783,N_19961);
and UO_1686 (O_1686,N_19807,N_19890);
and UO_1687 (O_1687,N_19788,N_19738);
or UO_1688 (O_1688,N_19977,N_19749);
nand UO_1689 (O_1689,N_19648,N_19920);
or UO_1690 (O_1690,N_19913,N_19872);
nand UO_1691 (O_1691,N_19791,N_19955);
xnor UO_1692 (O_1692,N_19891,N_19771);
xor UO_1693 (O_1693,N_19814,N_19605);
xnor UO_1694 (O_1694,N_19641,N_19674);
xor UO_1695 (O_1695,N_19604,N_19831);
nor UO_1696 (O_1696,N_19890,N_19626);
nand UO_1697 (O_1697,N_19854,N_19645);
or UO_1698 (O_1698,N_19834,N_19750);
and UO_1699 (O_1699,N_19685,N_19658);
xor UO_1700 (O_1700,N_19649,N_19888);
or UO_1701 (O_1701,N_19923,N_19689);
nand UO_1702 (O_1702,N_19995,N_19654);
nand UO_1703 (O_1703,N_19841,N_19982);
nand UO_1704 (O_1704,N_19786,N_19612);
and UO_1705 (O_1705,N_19789,N_19859);
or UO_1706 (O_1706,N_19881,N_19729);
or UO_1707 (O_1707,N_19959,N_19722);
nand UO_1708 (O_1708,N_19758,N_19731);
xor UO_1709 (O_1709,N_19706,N_19949);
or UO_1710 (O_1710,N_19842,N_19982);
xnor UO_1711 (O_1711,N_19779,N_19626);
or UO_1712 (O_1712,N_19625,N_19678);
xor UO_1713 (O_1713,N_19889,N_19841);
and UO_1714 (O_1714,N_19955,N_19995);
xnor UO_1715 (O_1715,N_19631,N_19944);
or UO_1716 (O_1716,N_19939,N_19765);
nand UO_1717 (O_1717,N_19803,N_19826);
nor UO_1718 (O_1718,N_19872,N_19718);
or UO_1719 (O_1719,N_19993,N_19698);
and UO_1720 (O_1720,N_19956,N_19636);
nand UO_1721 (O_1721,N_19751,N_19742);
xor UO_1722 (O_1722,N_19925,N_19724);
nor UO_1723 (O_1723,N_19825,N_19673);
xor UO_1724 (O_1724,N_19674,N_19753);
xnor UO_1725 (O_1725,N_19669,N_19909);
xor UO_1726 (O_1726,N_19948,N_19737);
and UO_1727 (O_1727,N_19741,N_19791);
or UO_1728 (O_1728,N_19762,N_19801);
or UO_1729 (O_1729,N_19881,N_19670);
nand UO_1730 (O_1730,N_19611,N_19698);
nand UO_1731 (O_1731,N_19636,N_19969);
xnor UO_1732 (O_1732,N_19994,N_19736);
xnor UO_1733 (O_1733,N_19855,N_19890);
nor UO_1734 (O_1734,N_19746,N_19702);
nand UO_1735 (O_1735,N_19629,N_19600);
or UO_1736 (O_1736,N_19754,N_19832);
nor UO_1737 (O_1737,N_19908,N_19983);
nor UO_1738 (O_1738,N_19941,N_19714);
xnor UO_1739 (O_1739,N_19795,N_19676);
and UO_1740 (O_1740,N_19708,N_19609);
nand UO_1741 (O_1741,N_19634,N_19692);
and UO_1742 (O_1742,N_19892,N_19660);
and UO_1743 (O_1743,N_19899,N_19669);
xor UO_1744 (O_1744,N_19960,N_19866);
nand UO_1745 (O_1745,N_19725,N_19756);
nor UO_1746 (O_1746,N_19944,N_19812);
xnor UO_1747 (O_1747,N_19970,N_19890);
xnor UO_1748 (O_1748,N_19609,N_19667);
and UO_1749 (O_1749,N_19988,N_19977);
nand UO_1750 (O_1750,N_19970,N_19753);
xor UO_1751 (O_1751,N_19927,N_19806);
xnor UO_1752 (O_1752,N_19688,N_19917);
xor UO_1753 (O_1753,N_19810,N_19764);
nor UO_1754 (O_1754,N_19825,N_19848);
and UO_1755 (O_1755,N_19735,N_19891);
nor UO_1756 (O_1756,N_19877,N_19879);
and UO_1757 (O_1757,N_19844,N_19760);
or UO_1758 (O_1758,N_19882,N_19778);
nand UO_1759 (O_1759,N_19622,N_19650);
or UO_1760 (O_1760,N_19849,N_19823);
nand UO_1761 (O_1761,N_19753,N_19773);
and UO_1762 (O_1762,N_19952,N_19890);
nor UO_1763 (O_1763,N_19618,N_19747);
and UO_1764 (O_1764,N_19687,N_19748);
or UO_1765 (O_1765,N_19745,N_19636);
and UO_1766 (O_1766,N_19957,N_19944);
or UO_1767 (O_1767,N_19601,N_19632);
nand UO_1768 (O_1768,N_19640,N_19882);
or UO_1769 (O_1769,N_19775,N_19770);
and UO_1770 (O_1770,N_19613,N_19934);
nand UO_1771 (O_1771,N_19909,N_19836);
nor UO_1772 (O_1772,N_19912,N_19768);
nor UO_1773 (O_1773,N_19846,N_19801);
nand UO_1774 (O_1774,N_19648,N_19745);
nor UO_1775 (O_1775,N_19922,N_19636);
or UO_1776 (O_1776,N_19773,N_19857);
xnor UO_1777 (O_1777,N_19725,N_19804);
nor UO_1778 (O_1778,N_19664,N_19895);
nand UO_1779 (O_1779,N_19915,N_19747);
nand UO_1780 (O_1780,N_19799,N_19726);
nand UO_1781 (O_1781,N_19785,N_19793);
and UO_1782 (O_1782,N_19849,N_19767);
xor UO_1783 (O_1783,N_19951,N_19898);
nand UO_1784 (O_1784,N_19704,N_19799);
nor UO_1785 (O_1785,N_19939,N_19933);
and UO_1786 (O_1786,N_19628,N_19671);
or UO_1787 (O_1787,N_19813,N_19850);
and UO_1788 (O_1788,N_19946,N_19803);
or UO_1789 (O_1789,N_19796,N_19619);
and UO_1790 (O_1790,N_19766,N_19665);
xnor UO_1791 (O_1791,N_19678,N_19804);
and UO_1792 (O_1792,N_19685,N_19710);
nand UO_1793 (O_1793,N_19867,N_19622);
nor UO_1794 (O_1794,N_19813,N_19749);
nand UO_1795 (O_1795,N_19988,N_19685);
nand UO_1796 (O_1796,N_19617,N_19654);
or UO_1797 (O_1797,N_19903,N_19921);
xor UO_1798 (O_1798,N_19950,N_19754);
nor UO_1799 (O_1799,N_19795,N_19608);
xor UO_1800 (O_1800,N_19912,N_19619);
and UO_1801 (O_1801,N_19877,N_19944);
and UO_1802 (O_1802,N_19709,N_19815);
nand UO_1803 (O_1803,N_19654,N_19661);
and UO_1804 (O_1804,N_19653,N_19834);
xor UO_1805 (O_1805,N_19688,N_19840);
xnor UO_1806 (O_1806,N_19874,N_19831);
xnor UO_1807 (O_1807,N_19731,N_19724);
xnor UO_1808 (O_1808,N_19882,N_19727);
and UO_1809 (O_1809,N_19651,N_19607);
nand UO_1810 (O_1810,N_19679,N_19737);
nor UO_1811 (O_1811,N_19882,N_19677);
or UO_1812 (O_1812,N_19891,N_19641);
or UO_1813 (O_1813,N_19794,N_19840);
nor UO_1814 (O_1814,N_19858,N_19604);
and UO_1815 (O_1815,N_19951,N_19932);
and UO_1816 (O_1816,N_19878,N_19969);
nand UO_1817 (O_1817,N_19634,N_19749);
xor UO_1818 (O_1818,N_19798,N_19738);
nor UO_1819 (O_1819,N_19938,N_19775);
nor UO_1820 (O_1820,N_19681,N_19818);
nand UO_1821 (O_1821,N_19831,N_19856);
or UO_1822 (O_1822,N_19716,N_19901);
nor UO_1823 (O_1823,N_19990,N_19920);
and UO_1824 (O_1824,N_19714,N_19753);
and UO_1825 (O_1825,N_19637,N_19975);
nand UO_1826 (O_1826,N_19836,N_19778);
or UO_1827 (O_1827,N_19967,N_19652);
nand UO_1828 (O_1828,N_19988,N_19676);
xor UO_1829 (O_1829,N_19761,N_19738);
or UO_1830 (O_1830,N_19810,N_19971);
and UO_1831 (O_1831,N_19853,N_19620);
xnor UO_1832 (O_1832,N_19699,N_19668);
or UO_1833 (O_1833,N_19981,N_19962);
or UO_1834 (O_1834,N_19952,N_19652);
or UO_1835 (O_1835,N_19943,N_19634);
and UO_1836 (O_1836,N_19796,N_19928);
nor UO_1837 (O_1837,N_19602,N_19649);
nor UO_1838 (O_1838,N_19786,N_19981);
or UO_1839 (O_1839,N_19973,N_19822);
or UO_1840 (O_1840,N_19984,N_19921);
or UO_1841 (O_1841,N_19840,N_19937);
nor UO_1842 (O_1842,N_19986,N_19701);
xnor UO_1843 (O_1843,N_19786,N_19977);
xor UO_1844 (O_1844,N_19710,N_19887);
or UO_1845 (O_1845,N_19943,N_19925);
or UO_1846 (O_1846,N_19669,N_19975);
and UO_1847 (O_1847,N_19841,N_19672);
xnor UO_1848 (O_1848,N_19653,N_19954);
nand UO_1849 (O_1849,N_19882,N_19668);
or UO_1850 (O_1850,N_19798,N_19610);
xnor UO_1851 (O_1851,N_19746,N_19745);
xor UO_1852 (O_1852,N_19727,N_19662);
xnor UO_1853 (O_1853,N_19832,N_19871);
nor UO_1854 (O_1854,N_19626,N_19644);
xor UO_1855 (O_1855,N_19931,N_19960);
or UO_1856 (O_1856,N_19705,N_19785);
and UO_1857 (O_1857,N_19881,N_19714);
nand UO_1858 (O_1858,N_19799,N_19974);
nor UO_1859 (O_1859,N_19608,N_19626);
nor UO_1860 (O_1860,N_19693,N_19823);
or UO_1861 (O_1861,N_19640,N_19681);
xor UO_1862 (O_1862,N_19769,N_19606);
and UO_1863 (O_1863,N_19938,N_19626);
or UO_1864 (O_1864,N_19954,N_19850);
nand UO_1865 (O_1865,N_19661,N_19666);
and UO_1866 (O_1866,N_19856,N_19803);
and UO_1867 (O_1867,N_19999,N_19833);
nand UO_1868 (O_1868,N_19805,N_19980);
or UO_1869 (O_1869,N_19625,N_19712);
or UO_1870 (O_1870,N_19792,N_19895);
nand UO_1871 (O_1871,N_19657,N_19690);
xor UO_1872 (O_1872,N_19728,N_19864);
xor UO_1873 (O_1873,N_19766,N_19724);
xor UO_1874 (O_1874,N_19851,N_19831);
or UO_1875 (O_1875,N_19910,N_19726);
nor UO_1876 (O_1876,N_19712,N_19927);
and UO_1877 (O_1877,N_19752,N_19896);
nand UO_1878 (O_1878,N_19777,N_19723);
and UO_1879 (O_1879,N_19930,N_19898);
nor UO_1880 (O_1880,N_19912,N_19841);
nor UO_1881 (O_1881,N_19787,N_19869);
xor UO_1882 (O_1882,N_19766,N_19756);
and UO_1883 (O_1883,N_19993,N_19797);
and UO_1884 (O_1884,N_19964,N_19640);
nand UO_1885 (O_1885,N_19916,N_19898);
xor UO_1886 (O_1886,N_19784,N_19728);
or UO_1887 (O_1887,N_19816,N_19695);
or UO_1888 (O_1888,N_19819,N_19673);
or UO_1889 (O_1889,N_19816,N_19746);
xor UO_1890 (O_1890,N_19652,N_19614);
nand UO_1891 (O_1891,N_19756,N_19616);
or UO_1892 (O_1892,N_19823,N_19947);
and UO_1893 (O_1893,N_19833,N_19880);
and UO_1894 (O_1894,N_19972,N_19857);
xor UO_1895 (O_1895,N_19622,N_19850);
or UO_1896 (O_1896,N_19601,N_19938);
and UO_1897 (O_1897,N_19797,N_19748);
and UO_1898 (O_1898,N_19925,N_19770);
or UO_1899 (O_1899,N_19797,N_19641);
and UO_1900 (O_1900,N_19941,N_19731);
xor UO_1901 (O_1901,N_19666,N_19837);
nor UO_1902 (O_1902,N_19710,N_19953);
nor UO_1903 (O_1903,N_19913,N_19999);
or UO_1904 (O_1904,N_19766,N_19604);
and UO_1905 (O_1905,N_19982,N_19678);
xnor UO_1906 (O_1906,N_19622,N_19643);
xor UO_1907 (O_1907,N_19770,N_19821);
xor UO_1908 (O_1908,N_19984,N_19771);
and UO_1909 (O_1909,N_19943,N_19977);
nor UO_1910 (O_1910,N_19743,N_19895);
xnor UO_1911 (O_1911,N_19945,N_19632);
nor UO_1912 (O_1912,N_19815,N_19887);
or UO_1913 (O_1913,N_19739,N_19737);
nor UO_1914 (O_1914,N_19740,N_19977);
nand UO_1915 (O_1915,N_19902,N_19748);
or UO_1916 (O_1916,N_19912,N_19838);
and UO_1917 (O_1917,N_19782,N_19659);
xnor UO_1918 (O_1918,N_19649,N_19766);
and UO_1919 (O_1919,N_19609,N_19870);
nor UO_1920 (O_1920,N_19924,N_19972);
and UO_1921 (O_1921,N_19952,N_19991);
xor UO_1922 (O_1922,N_19742,N_19758);
nor UO_1923 (O_1923,N_19892,N_19932);
and UO_1924 (O_1924,N_19667,N_19898);
or UO_1925 (O_1925,N_19885,N_19719);
or UO_1926 (O_1926,N_19763,N_19658);
nor UO_1927 (O_1927,N_19746,N_19679);
xor UO_1928 (O_1928,N_19634,N_19614);
nor UO_1929 (O_1929,N_19715,N_19703);
and UO_1930 (O_1930,N_19771,N_19800);
nand UO_1931 (O_1931,N_19799,N_19771);
and UO_1932 (O_1932,N_19843,N_19684);
or UO_1933 (O_1933,N_19841,N_19707);
xor UO_1934 (O_1934,N_19881,N_19741);
and UO_1935 (O_1935,N_19905,N_19790);
nor UO_1936 (O_1936,N_19637,N_19724);
nor UO_1937 (O_1937,N_19750,N_19732);
nor UO_1938 (O_1938,N_19874,N_19912);
nand UO_1939 (O_1939,N_19690,N_19907);
nand UO_1940 (O_1940,N_19792,N_19916);
nand UO_1941 (O_1941,N_19681,N_19827);
or UO_1942 (O_1942,N_19971,N_19758);
nor UO_1943 (O_1943,N_19754,N_19718);
xor UO_1944 (O_1944,N_19844,N_19854);
xnor UO_1945 (O_1945,N_19971,N_19825);
nor UO_1946 (O_1946,N_19891,N_19698);
or UO_1947 (O_1947,N_19987,N_19797);
and UO_1948 (O_1948,N_19886,N_19863);
and UO_1949 (O_1949,N_19660,N_19780);
or UO_1950 (O_1950,N_19967,N_19865);
nor UO_1951 (O_1951,N_19844,N_19997);
and UO_1952 (O_1952,N_19675,N_19665);
nor UO_1953 (O_1953,N_19967,N_19701);
nor UO_1954 (O_1954,N_19829,N_19606);
or UO_1955 (O_1955,N_19996,N_19845);
nand UO_1956 (O_1956,N_19766,N_19835);
nand UO_1957 (O_1957,N_19793,N_19621);
and UO_1958 (O_1958,N_19798,N_19715);
nand UO_1959 (O_1959,N_19933,N_19741);
or UO_1960 (O_1960,N_19883,N_19827);
and UO_1961 (O_1961,N_19693,N_19766);
or UO_1962 (O_1962,N_19856,N_19979);
or UO_1963 (O_1963,N_19708,N_19625);
nand UO_1964 (O_1964,N_19822,N_19938);
or UO_1965 (O_1965,N_19731,N_19791);
and UO_1966 (O_1966,N_19862,N_19733);
and UO_1967 (O_1967,N_19863,N_19676);
or UO_1968 (O_1968,N_19865,N_19977);
nor UO_1969 (O_1969,N_19796,N_19861);
nor UO_1970 (O_1970,N_19818,N_19770);
or UO_1971 (O_1971,N_19858,N_19787);
or UO_1972 (O_1972,N_19918,N_19949);
nor UO_1973 (O_1973,N_19698,N_19708);
xor UO_1974 (O_1974,N_19877,N_19987);
and UO_1975 (O_1975,N_19946,N_19663);
nand UO_1976 (O_1976,N_19706,N_19965);
nor UO_1977 (O_1977,N_19906,N_19892);
or UO_1978 (O_1978,N_19921,N_19948);
nand UO_1979 (O_1979,N_19963,N_19705);
nor UO_1980 (O_1980,N_19757,N_19900);
nor UO_1981 (O_1981,N_19695,N_19822);
xor UO_1982 (O_1982,N_19804,N_19615);
nand UO_1983 (O_1983,N_19829,N_19628);
nor UO_1984 (O_1984,N_19913,N_19940);
nand UO_1985 (O_1985,N_19984,N_19727);
and UO_1986 (O_1986,N_19854,N_19913);
and UO_1987 (O_1987,N_19681,N_19608);
nand UO_1988 (O_1988,N_19718,N_19774);
nor UO_1989 (O_1989,N_19740,N_19672);
or UO_1990 (O_1990,N_19811,N_19996);
nand UO_1991 (O_1991,N_19858,N_19835);
nand UO_1992 (O_1992,N_19638,N_19869);
nor UO_1993 (O_1993,N_19662,N_19810);
and UO_1994 (O_1994,N_19833,N_19897);
nor UO_1995 (O_1995,N_19924,N_19796);
nand UO_1996 (O_1996,N_19601,N_19925);
nor UO_1997 (O_1997,N_19898,N_19630);
xor UO_1998 (O_1998,N_19704,N_19825);
nor UO_1999 (O_1999,N_19975,N_19858);
xor UO_2000 (O_2000,N_19677,N_19927);
nand UO_2001 (O_2001,N_19669,N_19790);
or UO_2002 (O_2002,N_19709,N_19658);
xor UO_2003 (O_2003,N_19894,N_19600);
nand UO_2004 (O_2004,N_19672,N_19976);
nand UO_2005 (O_2005,N_19603,N_19688);
nand UO_2006 (O_2006,N_19885,N_19691);
xnor UO_2007 (O_2007,N_19671,N_19602);
or UO_2008 (O_2008,N_19874,N_19692);
nand UO_2009 (O_2009,N_19670,N_19974);
and UO_2010 (O_2010,N_19973,N_19697);
or UO_2011 (O_2011,N_19713,N_19876);
and UO_2012 (O_2012,N_19870,N_19678);
xor UO_2013 (O_2013,N_19929,N_19883);
and UO_2014 (O_2014,N_19797,N_19793);
nor UO_2015 (O_2015,N_19875,N_19648);
and UO_2016 (O_2016,N_19804,N_19760);
xor UO_2017 (O_2017,N_19681,N_19956);
xnor UO_2018 (O_2018,N_19685,N_19698);
and UO_2019 (O_2019,N_19994,N_19867);
nor UO_2020 (O_2020,N_19835,N_19763);
xnor UO_2021 (O_2021,N_19952,N_19762);
and UO_2022 (O_2022,N_19940,N_19877);
and UO_2023 (O_2023,N_19894,N_19761);
nand UO_2024 (O_2024,N_19694,N_19817);
nand UO_2025 (O_2025,N_19760,N_19607);
nor UO_2026 (O_2026,N_19634,N_19975);
nor UO_2027 (O_2027,N_19696,N_19929);
nor UO_2028 (O_2028,N_19758,N_19791);
xor UO_2029 (O_2029,N_19908,N_19657);
nor UO_2030 (O_2030,N_19802,N_19975);
or UO_2031 (O_2031,N_19763,N_19616);
or UO_2032 (O_2032,N_19621,N_19774);
xor UO_2033 (O_2033,N_19851,N_19625);
and UO_2034 (O_2034,N_19726,N_19870);
or UO_2035 (O_2035,N_19776,N_19766);
and UO_2036 (O_2036,N_19735,N_19908);
and UO_2037 (O_2037,N_19648,N_19971);
or UO_2038 (O_2038,N_19843,N_19733);
nor UO_2039 (O_2039,N_19659,N_19967);
xor UO_2040 (O_2040,N_19663,N_19658);
nand UO_2041 (O_2041,N_19932,N_19948);
nand UO_2042 (O_2042,N_19692,N_19791);
or UO_2043 (O_2043,N_19946,N_19995);
or UO_2044 (O_2044,N_19682,N_19735);
or UO_2045 (O_2045,N_19992,N_19833);
or UO_2046 (O_2046,N_19630,N_19690);
and UO_2047 (O_2047,N_19705,N_19623);
xor UO_2048 (O_2048,N_19631,N_19929);
nand UO_2049 (O_2049,N_19624,N_19674);
nand UO_2050 (O_2050,N_19756,N_19976);
and UO_2051 (O_2051,N_19800,N_19627);
nor UO_2052 (O_2052,N_19721,N_19664);
or UO_2053 (O_2053,N_19936,N_19788);
nand UO_2054 (O_2054,N_19909,N_19831);
nor UO_2055 (O_2055,N_19976,N_19688);
and UO_2056 (O_2056,N_19937,N_19715);
or UO_2057 (O_2057,N_19622,N_19762);
or UO_2058 (O_2058,N_19819,N_19984);
xnor UO_2059 (O_2059,N_19931,N_19915);
xor UO_2060 (O_2060,N_19909,N_19693);
or UO_2061 (O_2061,N_19668,N_19858);
nand UO_2062 (O_2062,N_19997,N_19803);
nand UO_2063 (O_2063,N_19661,N_19856);
nor UO_2064 (O_2064,N_19750,N_19821);
or UO_2065 (O_2065,N_19603,N_19966);
or UO_2066 (O_2066,N_19807,N_19967);
nand UO_2067 (O_2067,N_19619,N_19716);
nand UO_2068 (O_2068,N_19925,N_19750);
nor UO_2069 (O_2069,N_19950,N_19636);
nor UO_2070 (O_2070,N_19874,N_19978);
and UO_2071 (O_2071,N_19895,N_19933);
or UO_2072 (O_2072,N_19705,N_19610);
or UO_2073 (O_2073,N_19828,N_19816);
and UO_2074 (O_2074,N_19737,N_19718);
or UO_2075 (O_2075,N_19676,N_19792);
nand UO_2076 (O_2076,N_19842,N_19657);
xor UO_2077 (O_2077,N_19935,N_19718);
xnor UO_2078 (O_2078,N_19614,N_19635);
or UO_2079 (O_2079,N_19688,N_19849);
nor UO_2080 (O_2080,N_19806,N_19666);
and UO_2081 (O_2081,N_19691,N_19992);
xnor UO_2082 (O_2082,N_19871,N_19756);
xor UO_2083 (O_2083,N_19908,N_19649);
or UO_2084 (O_2084,N_19641,N_19715);
xnor UO_2085 (O_2085,N_19805,N_19737);
nor UO_2086 (O_2086,N_19630,N_19783);
and UO_2087 (O_2087,N_19740,N_19858);
xnor UO_2088 (O_2088,N_19977,N_19834);
nor UO_2089 (O_2089,N_19623,N_19977);
or UO_2090 (O_2090,N_19868,N_19790);
nor UO_2091 (O_2091,N_19728,N_19835);
or UO_2092 (O_2092,N_19763,N_19896);
nor UO_2093 (O_2093,N_19601,N_19716);
nor UO_2094 (O_2094,N_19921,N_19698);
and UO_2095 (O_2095,N_19978,N_19703);
nand UO_2096 (O_2096,N_19899,N_19902);
nand UO_2097 (O_2097,N_19684,N_19880);
nor UO_2098 (O_2098,N_19745,N_19977);
nor UO_2099 (O_2099,N_19717,N_19634);
xnor UO_2100 (O_2100,N_19700,N_19674);
xor UO_2101 (O_2101,N_19637,N_19928);
nand UO_2102 (O_2102,N_19899,N_19880);
xor UO_2103 (O_2103,N_19736,N_19665);
nand UO_2104 (O_2104,N_19728,N_19613);
xor UO_2105 (O_2105,N_19772,N_19884);
nor UO_2106 (O_2106,N_19996,N_19757);
nor UO_2107 (O_2107,N_19898,N_19728);
xor UO_2108 (O_2108,N_19746,N_19938);
nand UO_2109 (O_2109,N_19680,N_19650);
or UO_2110 (O_2110,N_19829,N_19825);
and UO_2111 (O_2111,N_19818,N_19874);
and UO_2112 (O_2112,N_19647,N_19753);
and UO_2113 (O_2113,N_19621,N_19994);
nand UO_2114 (O_2114,N_19638,N_19786);
nand UO_2115 (O_2115,N_19609,N_19797);
or UO_2116 (O_2116,N_19803,N_19719);
or UO_2117 (O_2117,N_19751,N_19823);
and UO_2118 (O_2118,N_19701,N_19807);
xor UO_2119 (O_2119,N_19839,N_19857);
or UO_2120 (O_2120,N_19693,N_19689);
nand UO_2121 (O_2121,N_19831,N_19792);
xnor UO_2122 (O_2122,N_19795,N_19925);
and UO_2123 (O_2123,N_19636,N_19828);
nand UO_2124 (O_2124,N_19844,N_19710);
or UO_2125 (O_2125,N_19849,N_19853);
and UO_2126 (O_2126,N_19852,N_19915);
or UO_2127 (O_2127,N_19896,N_19825);
and UO_2128 (O_2128,N_19929,N_19911);
and UO_2129 (O_2129,N_19811,N_19812);
nand UO_2130 (O_2130,N_19710,N_19799);
xor UO_2131 (O_2131,N_19975,N_19783);
nor UO_2132 (O_2132,N_19908,N_19935);
nor UO_2133 (O_2133,N_19707,N_19944);
or UO_2134 (O_2134,N_19924,N_19766);
xnor UO_2135 (O_2135,N_19871,N_19704);
and UO_2136 (O_2136,N_19913,N_19984);
xor UO_2137 (O_2137,N_19728,N_19740);
nand UO_2138 (O_2138,N_19718,N_19796);
and UO_2139 (O_2139,N_19848,N_19660);
or UO_2140 (O_2140,N_19796,N_19765);
nor UO_2141 (O_2141,N_19716,N_19994);
xnor UO_2142 (O_2142,N_19732,N_19788);
nand UO_2143 (O_2143,N_19997,N_19889);
xor UO_2144 (O_2144,N_19631,N_19827);
nand UO_2145 (O_2145,N_19638,N_19702);
nor UO_2146 (O_2146,N_19670,N_19730);
or UO_2147 (O_2147,N_19862,N_19686);
nor UO_2148 (O_2148,N_19958,N_19968);
nor UO_2149 (O_2149,N_19931,N_19606);
xor UO_2150 (O_2150,N_19694,N_19943);
and UO_2151 (O_2151,N_19740,N_19762);
and UO_2152 (O_2152,N_19827,N_19909);
nand UO_2153 (O_2153,N_19661,N_19778);
nand UO_2154 (O_2154,N_19893,N_19847);
or UO_2155 (O_2155,N_19841,N_19615);
nor UO_2156 (O_2156,N_19837,N_19813);
nand UO_2157 (O_2157,N_19679,N_19633);
or UO_2158 (O_2158,N_19873,N_19639);
or UO_2159 (O_2159,N_19911,N_19943);
and UO_2160 (O_2160,N_19662,N_19906);
xor UO_2161 (O_2161,N_19858,N_19662);
and UO_2162 (O_2162,N_19979,N_19607);
xnor UO_2163 (O_2163,N_19762,N_19855);
and UO_2164 (O_2164,N_19834,N_19925);
xor UO_2165 (O_2165,N_19806,N_19909);
and UO_2166 (O_2166,N_19861,N_19782);
and UO_2167 (O_2167,N_19670,N_19641);
xnor UO_2168 (O_2168,N_19699,N_19935);
xor UO_2169 (O_2169,N_19670,N_19649);
xor UO_2170 (O_2170,N_19807,N_19799);
or UO_2171 (O_2171,N_19880,N_19836);
nor UO_2172 (O_2172,N_19667,N_19968);
or UO_2173 (O_2173,N_19666,N_19964);
and UO_2174 (O_2174,N_19684,N_19750);
nand UO_2175 (O_2175,N_19993,N_19685);
and UO_2176 (O_2176,N_19973,N_19739);
xnor UO_2177 (O_2177,N_19801,N_19943);
or UO_2178 (O_2178,N_19902,N_19610);
xnor UO_2179 (O_2179,N_19816,N_19762);
nor UO_2180 (O_2180,N_19940,N_19848);
nor UO_2181 (O_2181,N_19659,N_19858);
xor UO_2182 (O_2182,N_19744,N_19633);
xnor UO_2183 (O_2183,N_19933,N_19901);
and UO_2184 (O_2184,N_19654,N_19785);
and UO_2185 (O_2185,N_19743,N_19619);
or UO_2186 (O_2186,N_19641,N_19619);
or UO_2187 (O_2187,N_19802,N_19796);
or UO_2188 (O_2188,N_19732,N_19798);
or UO_2189 (O_2189,N_19771,N_19682);
and UO_2190 (O_2190,N_19675,N_19674);
xnor UO_2191 (O_2191,N_19746,N_19821);
or UO_2192 (O_2192,N_19759,N_19677);
nor UO_2193 (O_2193,N_19697,N_19777);
nand UO_2194 (O_2194,N_19905,N_19704);
xnor UO_2195 (O_2195,N_19704,N_19697);
xnor UO_2196 (O_2196,N_19619,N_19727);
nand UO_2197 (O_2197,N_19957,N_19721);
or UO_2198 (O_2198,N_19831,N_19671);
nor UO_2199 (O_2199,N_19723,N_19847);
xor UO_2200 (O_2200,N_19866,N_19824);
nand UO_2201 (O_2201,N_19932,N_19991);
nor UO_2202 (O_2202,N_19627,N_19837);
and UO_2203 (O_2203,N_19766,N_19671);
and UO_2204 (O_2204,N_19912,N_19926);
xnor UO_2205 (O_2205,N_19676,N_19801);
xnor UO_2206 (O_2206,N_19770,N_19683);
nand UO_2207 (O_2207,N_19946,N_19881);
nand UO_2208 (O_2208,N_19848,N_19931);
xor UO_2209 (O_2209,N_19602,N_19916);
nand UO_2210 (O_2210,N_19842,N_19916);
or UO_2211 (O_2211,N_19852,N_19871);
nor UO_2212 (O_2212,N_19998,N_19691);
xor UO_2213 (O_2213,N_19841,N_19692);
nor UO_2214 (O_2214,N_19775,N_19773);
xnor UO_2215 (O_2215,N_19617,N_19627);
and UO_2216 (O_2216,N_19884,N_19838);
or UO_2217 (O_2217,N_19609,N_19672);
nand UO_2218 (O_2218,N_19602,N_19819);
or UO_2219 (O_2219,N_19778,N_19917);
nand UO_2220 (O_2220,N_19733,N_19697);
xor UO_2221 (O_2221,N_19919,N_19968);
or UO_2222 (O_2222,N_19802,N_19811);
or UO_2223 (O_2223,N_19706,N_19741);
xor UO_2224 (O_2224,N_19619,N_19961);
nor UO_2225 (O_2225,N_19769,N_19658);
nand UO_2226 (O_2226,N_19711,N_19895);
nor UO_2227 (O_2227,N_19864,N_19770);
or UO_2228 (O_2228,N_19918,N_19832);
nor UO_2229 (O_2229,N_19669,N_19837);
nand UO_2230 (O_2230,N_19957,N_19666);
nor UO_2231 (O_2231,N_19725,N_19694);
and UO_2232 (O_2232,N_19807,N_19615);
or UO_2233 (O_2233,N_19711,N_19850);
xnor UO_2234 (O_2234,N_19834,N_19984);
nand UO_2235 (O_2235,N_19641,N_19605);
nor UO_2236 (O_2236,N_19697,N_19827);
nor UO_2237 (O_2237,N_19849,N_19607);
xor UO_2238 (O_2238,N_19936,N_19819);
nor UO_2239 (O_2239,N_19893,N_19783);
xnor UO_2240 (O_2240,N_19819,N_19795);
and UO_2241 (O_2241,N_19828,N_19670);
xnor UO_2242 (O_2242,N_19726,N_19937);
nor UO_2243 (O_2243,N_19635,N_19673);
or UO_2244 (O_2244,N_19629,N_19782);
nand UO_2245 (O_2245,N_19914,N_19870);
nand UO_2246 (O_2246,N_19947,N_19974);
xnor UO_2247 (O_2247,N_19897,N_19718);
and UO_2248 (O_2248,N_19726,N_19872);
and UO_2249 (O_2249,N_19785,N_19896);
and UO_2250 (O_2250,N_19755,N_19824);
nand UO_2251 (O_2251,N_19652,N_19882);
or UO_2252 (O_2252,N_19995,N_19629);
or UO_2253 (O_2253,N_19824,N_19956);
xnor UO_2254 (O_2254,N_19837,N_19677);
and UO_2255 (O_2255,N_19998,N_19992);
xnor UO_2256 (O_2256,N_19838,N_19865);
and UO_2257 (O_2257,N_19714,N_19608);
nor UO_2258 (O_2258,N_19615,N_19732);
nor UO_2259 (O_2259,N_19900,N_19931);
nor UO_2260 (O_2260,N_19736,N_19898);
nor UO_2261 (O_2261,N_19879,N_19685);
xor UO_2262 (O_2262,N_19771,N_19653);
nor UO_2263 (O_2263,N_19777,N_19975);
and UO_2264 (O_2264,N_19712,N_19602);
and UO_2265 (O_2265,N_19751,N_19794);
xor UO_2266 (O_2266,N_19815,N_19965);
nand UO_2267 (O_2267,N_19832,N_19815);
or UO_2268 (O_2268,N_19860,N_19720);
xnor UO_2269 (O_2269,N_19833,N_19609);
xor UO_2270 (O_2270,N_19999,N_19706);
xnor UO_2271 (O_2271,N_19823,N_19611);
xnor UO_2272 (O_2272,N_19703,N_19905);
xnor UO_2273 (O_2273,N_19623,N_19970);
or UO_2274 (O_2274,N_19794,N_19811);
and UO_2275 (O_2275,N_19675,N_19994);
xnor UO_2276 (O_2276,N_19918,N_19923);
nor UO_2277 (O_2277,N_19994,N_19982);
and UO_2278 (O_2278,N_19762,N_19656);
nand UO_2279 (O_2279,N_19921,N_19950);
or UO_2280 (O_2280,N_19711,N_19775);
nand UO_2281 (O_2281,N_19940,N_19872);
nand UO_2282 (O_2282,N_19843,N_19941);
or UO_2283 (O_2283,N_19636,N_19622);
nand UO_2284 (O_2284,N_19894,N_19949);
nand UO_2285 (O_2285,N_19695,N_19968);
nor UO_2286 (O_2286,N_19687,N_19847);
and UO_2287 (O_2287,N_19963,N_19612);
nor UO_2288 (O_2288,N_19852,N_19780);
nand UO_2289 (O_2289,N_19768,N_19813);
xor UO_2290 (O_2290,N_19653,N_19764);
and UO_2291 (O_2291,N_19743,N_19883);
and UO_2292 (O_2292,N_19950,N_19869);
nor UO_2293 (O_2293,N_19780,N_19762);
and UO_2294 (O_2294,N_19818,N_19641);
nor UO_2295 (O_2295,N_19763,N_19700);
nand UO_2296 (O_2296,N_19822,N_19835);
xnor UO_2297 (O_2297,N_19942,N_19986);
nor UO_2298 (O_2298,N_19652,N_19656);
nor UO_2299 (O_2299,N_19650,N_19675);
and UO_2300 (O_2300,N_19613,N_19755);
and UO_2301 (O_2301,N_19868,N_19724);
xnor UO_2302 (O_2302,N_19895,N_19878);
and UO_2303 (O_2303,N_19732,N_19686);
and UO_2304 (O_2304,N_19821,N_19717);
xor UO_2305 (O_2305,N_19939,N_19839);
or UO_2306 (O_2306,N_19785,N_19665);
and UO_2307 (O_2307,N_19766,N_19860);
and UO_2308 (O_2308,N_19898,N_19842);
and UO_2309 (O_2309,N_19661,N_19876);
nand UO_2310 (O_2310,N_19975,N_19981);
xor UO_2311 (O_2311,N_19822,N_19688);
and UO_2312 (O_2312,N_19701,N_19844);
or UO_2313 (O_2313,N_19848,N_19697);
nor UO_2314 (O_2314,N_19705,N_19833);
xnor UO_2315 (O_2315,N_19611,N_19890);
nor UO_2316 (O_2316,N_19993,N_19881);
nand UO_2317 (O_2317,N_19963,N_19907);
or UO_2318 (O_2318,N_19751,N_19781);
xor UO_2319 (O_2319,N_19989,N_19955);
nor UO_2320 (O_2320,N_19877,N_19986);
and UO_2321 (O_2321,N_19744,N_19778);
or UO_2322 (O_2322,N_19603,N_19914);
nor UO_2323 (O_2323,N_19685,N_19992);
xnor UO_2324 (O_2324,N_19956,N_19678);
and UO_2325 (O_2325,N_19673,N_19828);
and UO_2326 (O_2326,N_19800,N_19992);
or UO_2327 (O_2327,N_19905,N_19806);
xor UO_2328 (O_2328,N_19787,N_19661);
or UO_2329 (O_2329,N_19682,N_19717);
nand UO_2330 (O_2330,N_19807,N_19926);
xor UO_2331 (O_2331,N_19630,N_19616);
xor UO_2332 (O_2332,N_19714,N_19993);
and UO_2333 (O_2333,N_19655,N_19743);
xnor UO_2334 (O_2334,N_19917,N_19705);
nand UO_2335 (O_2335,N_19780,N_19666);
nor UO_2336 (O_2336,N_19603,N_19785);
nor UO_2337 (O_2337,N_19943,N_19716);
and UO_2338 (O_2338,N_19823,N_19888);
xor UO_2339 (O_2339,N_19774,N_19784);
nand UO_2340 (O_2340,N_19989,N_19899);
and UO_2341 (O_2341,N_19946,N_19619);
xnor UO_2342 (O_2342,N_19994,N_19938);
or UO_2343 (O_2343,N_19934,N_19608);
and UO_2344 (O_2344,N_19995,N_19737);
nor UO_2345 (O_2345,N_19602,N_19717);
nand UO_2346 (O_2346,N_19991,N_19672);
xor UO_2347 (O_2347,N_19649,N_19880);
or UO_2348 (O_2348,N_19965,N_19665);
xor UO_2349 (O_2349,N_19999,N_19976);
and UO_2350 (O_2350,N_19674,N_19803);
or UO_2351 (O_2351,N_19682,N_19704);
nand UO_2352 (O_2352,N_19727,N_19914);
and UO_2353 (O_2353,N_19604,N_19984);
or UO_2354 (O_2354,N_19794,N_19819);
nand UO_2355 (O_2355,N_19988,N_19951);
xnor UO_2356 (O_2356,N_19800,N_19735);
nor UO_2357 (O_2357,N_19699,N_19920);
nor UO_2358 (O_2358,N_19946,N_19804);
and UO_2359 (O_2359,N_19890,N_19910);
nand UO_2360 (O_2360,N_19681,N_19666);
and UO_2361 (O_2361,N_19932,N_19794);
or UO_2362 (O_2362,N_19814,N_19897);
and UO_2363 (O_2363,N_19970,N_19761);
nor UO_2364 (O_2364,N_19754,N_19658);
nand UO_2365 (O_2365,N_19842,N_19683);
xor UO_2366 (O_2366,N_19665,N_19890);
xnor UO_2367 (O_2367,N_19713,N_19826);
xor UO_2368 (O_2368,N_19982,N_19652);
nor UO_2369 (O_2369,N_19941,N_19874);
or UO_2370 (O_2370,N_19909,N_19985);
and UO_2371 (O_2371,N_19850,N_19733);
xnor UO_2372 (O_2372,N_19628,N_19621);
nor UO_2373 (O_2373,N_19841,N_19741);
xnor UO_2374 (O_2374,N_19992,N_19855);
or UO_2375 (O_2375,N_19754,N_19604);
nand UO_2376 (O_2376,N_19867,N_19734);
nor UO_2377 (O_2377,N_19721,N_19746);
nand UO_2378 (O_2378,N_19742,N_19628);
or UO_2379 (O_2379,N_19669,N_19985);
and UO_2380 (O_2380,N_19792,N_19930);
nor UO_2381 (O_2381,N_19762,N_19684);
nand UO_2382 (O_2382,N_19931,N_19842);
nand UO_2383 (O_2383,N_19612,N_19994);
nor UO_2384 (O_2384,N_19655,N_19859);
xnor UO_2385 (O_2385,N_19856,N_19692);
and UO_2386 (O_2386,N_19623,N_19902);
and UO_2387 (O_2387,N_19640,N_19999);
and UO_2388 (O_2388,N_19698,N_19824);
nor UO_2389 (O_2389,N_19797,N_19781);
or UO_2390 (O_2390,N_19946,N_19694);
nor UO_2391 (O_2391,N_19806,N_19703);
nand UO_2392 (O_2392,N_19941,N_19655);
nand UO_2393 (O_2393,N_19661,N_19733);
nand UO_2394 (O_2394,N_19777,N_19767);
nor UO_2395 (O_2395,N_19769,N_19730);
or UO_2396 (O_2396,N_19644,N_19760);
or UO_2397 (O_2397,N_19608,N_19972);
or UO_2398 (O_2398,N_19776,N_19953);
nor UO_2399 (O_2399,N_19933,N_19717);
or UO_2400 (O_2400,N_19680,N_19965);
xnor UO_2401 (O_2401,N_19766,N_19644);
nand UO_2402 (O_2402,N_19606,N_19985);
and UO_2403 (O_2403,N_19877,N_19723);
nor UO_2404 (O_2404,N_19659,N_19704);
nor UO_2405 (O_2405,N_19636,N_19750);
nand UO_2406 (O_2406,N_19970,N_19644);
nor UO_2407 (O_2407,N_19903,N_19868);
and UO_2408 (O_2408,N_19803,N_19846);
nor UO_2409 (O_2409,N_19726,N_19939);
and UO_2410 (O_2410,N_19687,N_19834);
and UO_2411 (O_2411,N_19657,N_19654);
nor UO_2412 (O_2412,N_19773,N_19705);
nor UO_2413 (O_2413,N_19988,N_19990);
nor UO_2414 (O_2414,N_19792,N_19872);
nand UO_2415 (O_2415,N_19892,N_19863);
nand UO_2416 (O_2416,N_19738,N_19656);
xor UO_2417 (O_2417,N_19892,N_19778);
and UO_2418 (O_2418,N_19646,N_19815);
nor UO_2419 (O_2419,N_19719,N_19854);
nand UO_2420 (O_2420,N_19738,N_19725);
or UO_2421 (O_2421,N_19696,N_19785);
nor UO_2422 (O_2422,N_19828,N_19939);
xnor UO_2423 (O_2423,N_19744,N_19975);
and UO_2424 (O_2424,N_19757,N_19660);
nand UO_2425 (O_2425,N_19973,N_19978);
xnor UO_2426 (O_2426,N_19732,N_19707);
nor UO_2427 (O_2427,N_19967,N_19692);
xor UO_2428 (O_2428,N_19772,N_19955);
and UO_2429 (O_2429,N_19798,N_19919);
or UO_2430 (O_2430,N_19646,N_19810);
and UO_2431 (O_2431,N_19890,N_19990);
or UO_2432 (O_2432,N_19934,N_19964);
and UO_2433 (O_2433,N_19764,N_19793);
nand UO_2434 (O_2434,N_19714,N_19911);
xor UO_2435 (O_2435,N_19631,N_19838);
and UO_2436 (O_2436,N_19752,N_19769);
and UO_2437 (O_2437,N_19815,N_19661);
xor UO_2438 (O_2438,N_19984,N_19846);
xnor UO_2439 (O_2439,N_19689,N_19661);
nand UO_2440 (O_2440,N_19819,N_19744);
nand UO_2441 (O_2441,N_19601,N_19970);
nand UO_2442 (O_2442,N_19732,N_19904);
xor UO_2443 (O_2443,N_19610,N_19856);
nand UO_2444 (O_2444,N_19740,N_19968);
and UO_2445 (O_2445,N_19808,N_19937);
xnor UO_2446 (O_2446,N_19919,N_19986);
nor UO_2447 (O_2447,N_19825,N_19968);
xor UO_2448 (O_2448,N_19985,N_19982);
xor UO_2449 (O_2449,N_19724,N_19743);
nor UO_2450 (O_2450,N_19847,N_19913);
nand UO_2451 (O_2451,N_19627,N_19784);
nand UO_2452 (O_2452,N_19934,N_19704);
xor UO_2453 (O_2453,N_19954,N_19760);
nand UO_2454 (O_2454,N_19816,N_19612);
xnor UO_2455 (O_2455,N_19858,N_19914);
nor UO_2456 (O_2456,N_19719,N_19852);
or UO_2457 (O_2457,N_19698,N_19954);
nor UO_2458 (O_2458,N_19611,N_19709);
nor UO_2459 (O_2459,N_19762,N_19736);
and UO_2460 (O_2460,N_19636,N_19787);
nor UO_2461 (O_2461,N_19998,N_19676);
and UO_2462 (O_2462,N_19641,N_19877);
nand UO_2463 (O_2463,N_19960,N_19812);
nand UO_2464 (O_2464,N_19845,N_19903);
nor UO_2465 (O_2465,N_19947,N_19636);
or UO_2466 (O_2466,N_19885,N_19932);
and UO_2467 (O_2467,N_19880,N_19941);
and UO_2468 (O_2468,N_19937,N_19865);
nor UO_2469 (O_2469,N_19818,N_19925);
xor UO_2470 (O_2470,N_19974,N_19913);
nand UO_2471 (O_2471,N_19800,N_19939);
nor UO_2472 (O_2472,N_19631,N_19909);
and UO_2473 (O_2473,N_19640,N_19867);
or UO_2474 (O_2474,N_19938,N_19693);
or UO_2475 (O_2475,N_19796,N_19915);
or UO_2476 (O_2476,N_19872,N_19620);
nand UO_2477 (O_2477,N_19714,N_19935);
nand UO_2478 (O_2478,N_19918,N_19980);
nand UO_2479 (O_2479,N_19658,N_19623);
nor UO_2480 (O_2480,N_19883,N_19783);
nand UO_2481 (O_2481,N_19922,N_19998);
xnor UO_2482 (O_2482,N_19864,N_19880);
xor UO_2483 (O_2483,N_19842,N_19926);
nor UO_2484 (O_2484,N_19883,N_19839);
or UO_2485 (O_2485,N_19948,N_19906);
or UO_2486 (O_2486,N_19712,N_19716);
and UO_2487 (O_2487,N_19990,N_19650);
or UO_2488 (O_2488,N_19837,N_19699);
or UO_2489 (O_2489,N_19943,N_19745);
nand UO_2490 (O_2490,N_19678,N_19851);
nand UO_2491 (O_2491,N_19605,N_19794);
nor UO_2492 (O_2492,N_19612,N_19690);
nand UO_2493 (O_2493,N_19897,N_19775);
or UO_2494 (O_2494,N_19983,N_19749);
nor UO_2495 (O_2495,N_19871,N_19876);
nor UO_2496 (O_2496,N_19987,N_19984);
and UO_2497 (O_2497,N_19822,N_19898);
or UO_2498 (O_2498,N_19750,N_19950);
nor UO_2499 (O_2499,N_19699,N_19948);
endmodule