module basic_3000_30000_3500_20_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_354,In_2212);
xnor U1 (N_1,In_1887,In_2438);
nand U2 (N_2,In_2375,In_1732);
nand U3 (N_3,In_1465,In_2678);
nor U4 (N_4,In_2394,In_2634);
or U5 (N_5,In_2293,In_2819);
and U6 (N_6,In_1260,In_1855);
and U7 (N_7,In_592,In_1312);
xor U8 (N_8,In_1988,In_74);
nor U9 (N_9,In_1379,In_2268);
xnor U10 (N_10,In_1675,In_703);
and U11 (N_11,In_1481,In_1576);
or U12 (N_12,In_1021,In_1181);
and U13 (N_13,In_1192,In_1534);
or U14 (N_14,In_568,In_1536);
xnor U15 (N_15,In_753,In_201);
xnor U16 (N_16,In_483,In_321);
and U17 (N_17,In_1259,In_1822);
xor U18 (N_18,In_2183,In_2361);
and U19 (N_19,In_2686,In_2692);
nand U20 (N_20,In_1839,In_1191);
nand U21 (N_21,In_784,In_370);
or U22 (N_22,In_424,In_2170);
or U23 (N_23,In_115,In_1281);
nor U24 (N_24,In_2453,In_33);
nor U25 (N_25,In_941,In_39);
and U26 (N_26,In_913,In_478);
xor U27 (N_27,In_1370,In_1299);
or U28 (N_28,In_1507,In_2858);
or U29 (N_29,In_396,In_439);
and U30 (N_30,In_1199,In_2639);
nand U31 (N_31,In_1118,In_1439);
or U32 (N_32,In_1375,In_1940);
nor U33 (N_33,In_1339,In_2315);
nor U34 (N_34,In_672,In_1078);
and U35 (N_35,In_1566,In_205);
xnor U36 (N_36,In_812,In_1937);
nand U37 (N_37,In_63,In_352);
nand U38 (N_38,In_258,In_2613);
or U39 (N_39,In_2231,In_195);
nand U40 (N_40,In_1275,In_2216);
or U41 (N_41,In_799,In_13);
and U42 (N_42,In_2680,In_1911);
nand U43 (N_43,In_1698,In_374);
nand U44 (N_44,In_297,In_1955);
and U45 (N_45,In_1458,In_890);
xor U46 (N_46,In_1431,In_877);
or U47 (N_47,In_234,In_184);
xnor U48 (N_48,In_1564,In_2380);
and U49 (N_49,In_2500,In_2984);
nor U50 (N_50,In_2239,In_1349);
or U51 (N_51,In_612,In_2079);
nor U52 (N_52,In_2395,In_754);
nor U53 (N_53,In_1969,In_246);
and U54 (N_54,In_698,In_1217);
or U55 (N_55,In_323,In_269);
or U56 (N_56,In_2952,In_1622);
and U57 (N_57,In_1309,In_2103);
nand U58 (N_58,In_1963,In_2448);
nand U59 (N_59,In_2367,In_2476);
nor U60 (N_60,In_1501,In_1502);
nand U61 (N_61,In_1215,In_143);
and U62 (N_62,In_2196,In_2875);
xor U63 (N_63,In_405,In_80);
and U64 (N_64,In_249,In_908);
xor U65 (N_65,In_2527,In_2768);
xor U66 (N_66,In_440,In_712);
or U67 (N_67,In_1594,In_2757);
nand U68 (N_68,In_1610,In_1306);
nor U69 (N_69,In_2495,In_418);
and U70 (N_70,In_1877,In_789);
nand U71 (N_71,In_1210,In_1122);
nor U72 (N_72,In_2646,In_2581);
nand U73 (N_73,In_845,In_180);
xnor U74 (N_74,In_1952,In_2415);
nand U75 (N_75,In_2083,In_846);
and U76 (N_76,In_1853,In_35);
nor U77 (N_77,In_1561,In_1512);
or U78 (N_78,In_1117,In_2568);
nor U79 (N_79,In_1523,In_2508);
xor U80 (N_80,In_410,In_1520);
nor U81 (N_81,In_1335,In_574);
nor U82 (N_82,In_2166,In_2266);
xor U83 (N_83,In_2350,In_1825);
nor U84 (N_84,In_818,In_2140);
and U85 (N_85,In_2718,In_2082);
or U86 (N_86,In_891,In_1320);
nand U87 (N_87,In_1796,In_2635);
nor U88 (N_88,In_2398,In_874);
nand U89 (N_89,In_2328,In_2431);
xor U90 (N_90,In_618,In_1279);
or U91 (N_91,In_1452,In_1263);
and U92 (N_92,In_779,In_1637);
nand U93 (N_93,In_1999,In_815);
or U94 (N_94,In_2969,In_947);
or U95 (N_95,In_1090,In_1683);
nand U96 (N_96,In_2993,In_2533);
nor U97 (N_97,In_2782,In_512);
nor U98 (N_98,In_2254,In_1100);
xnor U99 (N_99,In_2110,In_121);
nand U100 (N_100,In_2545,In_1112);
xnor U101 (N_101,In_442,In_900);
or U102 (N_102,In_606,In_2296);
nor U103 (N_103,In_2576,In_1129);
nand U104 (N_104,In_2649,In_484);
and U105 (N_105,In_2209,In_2619);
and U106 (N_106,In_2148,In_811);
nor U107 (N_107,In_1466,In_2679);
and U108 (N_108,In_2674,In_1961);
or U109 (N_109,In_746,In_1945);
nor U110 (N_110,In_1124,In_542);
or U111 (N_111,In_1904,In_1020);
nor U112 (N_112,In_2488,In_1667);
or U113 (N_113,In_1696,In_2187);
or U114 (N_114,In_1885,In_579);
xnor U115 (N_115,In_2567,In_481);
xnor U116 (N_116,In_128,In_1156);
and U117 (N_117,In_960,In_675);
and U118 (N_118,In_2849,In_373);
nand U119 (N_119,In_622,In_2735);
xnor U120 (N_120,In_43,In_2316);
or U121 (N_121,In_2552,In_2566);
nand U122 (N_122,In_2624,In_589);
nand U123 (N_123,In_2366,In_2549);
and U124 (N_124,In_262,In_925);
xnor U125 (N_125,In_1066,In_1775);
and U126 (N_126,In_2317,In_1503);
nor U127 (N_127,In_2672,In_2155);
nand U128 (N_128,In_2075,In_767);
and U129 (N_129,In_1454,In_2242);
xnor U130 (N_130,In_267,In_2949);
nor U131 (N_131,In_1302,In_1892);
nor U132 (N_132,In_404,In_2588);
nor U133 (N_133,In_1073,In_2131);
nor U134 (N_134,In_2972,In_2353);
nand U135 (N_135,In_2825,In_700);
nor U136 (N_136,In_780,In_1074);
and U137 (N_137,In_52,In_515);
and U138 (N_138,In_1803,In_2682);
xnor U139 (N_139,In_1994,In_2026);
xor U140 (N_140,In_1120,In_2404);
or U141 (N_141,In_2062,In_1453);
nand U142 (N_142,In_2199,In_1041);
nand U143 (N_143,In_29,In_2863);
nor U144 (N_144,In_2313,In_1926);
or U145 (N_145,In_556,In_487);
and U146 (N_146,In_2294,In_1906);
nand U147 (N_147,In_907,In_2911);
nor U148 (N_148,In_601,In_1437);
xor U149 (N_149,In_1258,In_607);
and U150 (N_150,In_1462,In_2287);
and U151 (N_151,In_96,In_957);
nor U152 (N_152,In_2388,In_2805);
and U153 (N_153,In_317,In_26);
nand U154 (N_154,In_1901,In_2421);
and U155 (N_155,In_2464,In_2539);
xnor U156 (N_156,In_1827,In_2893);
and U157 (N_157,In_881,In_2164);
nand U158 (N_158,In_572,In_855);
nor U159 (N_159,In_537,In_1135);
and U160 (N_160,In_1671,In_2876);
xor U161 (N_161,In_1017,In_1652);
or U162 (N_162,In_2073,In_2561);
or U163 (N_163,In_518,In_1939);
nor U164 (N_164,In_231,In_2710);
nand U165 (N_165,In_1209,In_318);
and U166 (N_166,In_1096,In_4);
xnor U167 (N_167,In_1282,In_2990);
nor U168 (N_168,In_669,In_1704);
nand U169 (N_169,In_1088,In_350);
nand U170 (N_170,In_1674,In_1089);
and U171 (N_171,In_1542,In_2031);
or U172 (N_172,In_1693,In_2900);
nor U173 (N_173,In_1980,In_1322);
or U174 (N_174,In_507,In_1527);
nor U175 (N_175,In_463,In_641);
nor U176 (N_176,In_1278,In_1574);
nand U177 (N_177,In_2493,In_2470);
nor U178 (N_178,In_1085,In_1037);
nand U179 (N_179,In_2355,In_1552);
and U180 (N_180,In_1024,In_1551);
xor U181 (N_181,In_462,In_1011);
nor U182 (N_182,In_1423,In_787);
or U183 (N_183,In_539,In_1603);
and U184 (N_184,In_1075,In_2924);
xnor U185 (N_185,In_224,In_1947);
nand U186 (N_186,In_998,In_1076);
nor U187 (N_187,In_132,In_673);
xor U188 (N_188,In_173,In_2618);
and U189 (N_189,In_492,In_2905);
xor U190 (N_190,In_2102,In_2886);
or U191 (N_191,In_682,In_118);
nand U192 (N_192,In_1055,In_886);
or U193 (N_193,In_2694,In_2705);
and U194 (N_194,In_788,In_2486);
or U195 (N_195,In_795,In_803);
and U196 (N_196,In_1558,In_1457);
xor U197 (N_197,In_2336,In_166);
nor U198 (N_198,In_2450,In_285);
or U199 (N_199,In_1966,In_1851);
xor U200 (N_200,In_752,In_2363);
nor U201 (N_201,In_2163,In_367);
nand U202 (N_202,In_516,In_561);
xnor U203 (N_203,In_841,In_705);
nand U204 (N_204,In_2124,In_2114);
and U205 (N_205,In_1202,In_1162);
nor U206 (N_206,In_2841,In_375);
nor U207 (N_207,In_451,In_959);
nand U208 (N_208,In_2097,In_2746);
xnor U209 (N_209,In_320,In_1747);
xor U210 (N_210,In_808,In_1758);
and U211 (N_211,In_1060,In_1863);
and U212 (N_212,In_168,In_2788);
and U213 (N_213,In_500,In_1658);
and U214 (N_214,In_1004,In_2414);
or U215 (N_215,In_2643,In_804);
xor U216 (N_216,In_1972,In_809);
xnor U217 (N_217,In_2116,In_1170);
nand U218 (N_218,In_384,In_1480);
nor U219 (N_219,In_2880,In_2853);
nor U220 (N_220,In_600,In_963);
xor U221 (N_221,In_2338,In_232);
and U222 (N_222,In_726,In_2335);
nand U223 (N_223,In_2071,In_1139);
xor U224 (N_224,In_1500,In_1585);
xor U225 (N_225,In_54,In_415);
nor U226 (N_226,In_1266,In_1811);
or U227 (N_227,In_1705,In_2481);
or U228 (N_228,In_657,In_1183);
nor U229 (N_229,In_69,In_1272);
nor U230 (N_230,In_2751,In_2227);
or U231 (N_231,In_78,In_2530);
or U232 (N_232,In_72,In_873);
or U233 (N_233,In_1915,In_362);
nand U234 (N_234,In_1201,In_1657);
nand U235 (N_235,In_2354,In_599);
nand U236 (N_236,In_697,In_2191);
or U237 (N_237,In_1922,In_2241);
and U238 (N_238,In_2501,In_1097);
or U239 (N_239,In_2745,In_2654);
nor U240 (N_240,In_1896,In_2748);
nand U241 (N_241,In_526,In_1932);
nor U242 (N_242,In_2659,In_151);
nor U243 (N_243,In_316,In_402);
nor U244 (N_244,In_2010,In_903);
xor U245 (N_245,In_1185,In_1736);
nor U246 (N_246,In_2771,In_762);
nand U247 (N_247,In_2340,In_626);
or U248 (N_248,In_2428,In_2273);
nor U249 (N_249,In_1713,In_2221);
nor U250 (N_250,In_668,In_1575);
and U251 (N_251,In_2332,In_2295);
xnor U252 (N_252,In_1759,In_608);
xor U253 (N_253,In_2383,In_560);
nor U254 (N_254,In_508,In_2714);
and U255 (N_255,In_117,In_2756);
nor U256 (N_256,In_1164,In_1848);
and U257 (N_257,In_1921,In_1391);
nor U258 (N_258,In_984,In_2507);
or U259 (N_259,In_1236,In_2057);
or U260 (N_260,In_1269,In_1095);
nand U261 (N_261,In_2312,In_2277);
or U262 (N_262,In_338,In_441);
nand U263 (N_263,In_2726,In_421);
nand U264 (N_264,In_2234,In_1353);
and U265 (N_265,In_2218,In_167);
nand U266 (N_266,In_2593,In_1402);
and U267 (N_267,In_1948,In_2167);
and U268 (N_268,In_2783,In_2696);
nor U269 (N_269,In_1376,In_2046);
or U270 (N_270,In_220,In_2836);
or U271 (N_271,In_1860,In_830);
and U272 (N_272,In_2025,In_334);
and U273 (N_273,In_1769,In_2769);
xnor U274 (N_274,In_1451,In_98);
nor U275 (N_275,In_1250,In_2645);
and U276 (N_276,In_319,In_2651);
or U277 (N_277,In_620,In_41);
and U278 (N_278,In_307,In_296);
nor U279 (N_279,In_2220,In_196);
xnor U280 (N_280,In_2877,In_264);
nand U281 (N_281,In_1242,In_2105);
or U282 (N_282,In_2292,In_1418);
xnor U283 (N_283,In_1742,In_2667);
and U284 (N_284,In_1783,In_2707);
or U285 (N_285,In_1509,In_58);
xor U286 (N_286,In_1583,In_2349);
nand U287 (N_287,In_2675,In_2490);
xnor U288 (N_288,In_2406,In_1408);
or U289 (N_289,In_1599,In_2542);
xnor U290 (N_290,In_486,In_2120);
xor U291 (N_291,In_386,In_2740);
and U292 (N_292,In_422,In_1161);
and U293 (N_293,In_2407,In_152);
xor U294 (N_294,In_394,In_2232);
or U295 (N_295,In_1363,In_2719);
nand U296 (N_296,In_1790,In_2637);
xnor U297 (N_297,In_1433,In_684);
xnor U298 (N_298,In_2595,In_342);
or U299 (N_299,In_2118,In_2846);
xnor U300 (N_300,In_1256,In_2784);
nand U301 (N_301,In_2405,In_2504);
and U302 (N_302,In_2011,In_635);
nor U303 (N_303,In_663,In_828);
and U304 (N_304,In_2325,In_1560);
nand U305 (N_305,In_1590,In_2016);
and U306 (N_306,In_1337,In_2061);
nand U307 (N_307,In_227,In_1265);
or U308 (N_308,In_2633,In_2460);
and U309 (N_309,In_2134,In_47);
or U310 (N_310,In_2629,In_2240);
and U311 (N_311,In_1013,In_2895);
nand U312 (N_312,In_2224,In_329);
nand U313 (N_313,In_1111,In_208);
and U314 (N_314,In_692,In_1329);
nor U315 (N_315,In_793,In_2200);
nor U316 (N_316,In_708,In_1989);
xnor U317 (N_317,In_688,In_2898);
or U318 (N_318,In_1608,In_1600);
nor U319 (N_319,In_938,In_751);
xnor U320 (N_320,In_885,In_2289);
nor U321 (N_321,In_411,In_2014);
xnor U322 (N_322,In_2699,In_1795);
and U323 (N_323,In_2891,In_2485);
or U324 (N_324,In_1018,In_810);
xnor U325 (N_325,In_948,In_2092);
nor U326 (N_326,In_1328,In_188);
xor U327 (N_327,In_1800,In_2766);
or U328 (N_328,In_1725,In_2797);
and U329 (N_329,In_980,In_981);
or U330 (N_330,In_123,In_813);
nor U331 (N_331,In_2474,In_1861);
and U332 (N_332,In_1837,In_2456);
or U333 (N_333,In_2838,In_1717);
xor U334 (N_334,In_2435,In_2729);
or U335 (N_335,In_1058,In_1008);
or U336 (N_336,In_1787,In_251);
xnor U337 (N_337,In_2653,In_2562);
and U338 (N_338,In_1031,In_1455);
nand U339 (N_339,In_1276,In_615);
nand U340 (N_340,In_1193,In_1160);
or U341 (N_341,In_679,In_2081);
xnor U342 (N_342,In_412,In_315);
or U343 (N_343,In_1186,In_1680);
and U344 (N_344,In_2440,In_2845);
xnor U345 (N_345,In_503,In_1548);
nor U346 (N_346,In_1214,In_1753);
or U347 (N_347,In_2319,In_936);
or U348 (N_348,In_1425,In_674);
and U349 (N_349,In_369,In_2144);
nor U350 (N_350,In_2462,In_1155);
and U351 (N_351,In_717,In_2973);
or U352 (N_352,In_255,In_2871);
and U353 (N_353,In_1721,In_339);
nor U354 (N_354,In_2150,In_897);
nand U355 (N_355,In_671,In_2824);
or U356 (N_356,In_2641,In_860);
nor U357 (N_357,In_1687,In_119);
and U358 (N_358,In_2798,In_67);
nand U359 (N_359,In_453,In_1812);
xnor U360 (N_360,In_313,In_979);
xor U361 (N_361,In_216,In_156);
or U362 (N_362,In_1581,In_1879);
nor U363 (N_363,In_2712,In_1629);
and U364 (N_364,In_2555,In_178);
xnor U365 (N_365,In_736,In_2760);
xnor U366 (N_366,In_1189,In_1356);
or U367 (N_367,In_2205,In_2777);
or U368 (N_368,In_2622,In_2035);
nand U369 (N_369,In_2934,In_2019);
and U370 (N_370,In_77,In_892);
and U371 (N_371,In_609,In_546);
and U372 (N_372,In_2070,In_2452);
and U373 (N_373,In_870,In_433);
or U374 (N_374,In_1805,In_1247);
and U375 (N_375,In_164,In_1981);
nand U376 (N_376,In_1472,In_2283);
xnor U377 (N_377,In_2517,In_2970);
nand U378 (N_378,In_2104,In_2430);
xor U379 (N_379,In_357,In_2827);
and U380 (N_380,In_2506,In_1146);
xnor U381 (N_381,In_934,In_2357);
or U382 (N_382,In_2575,In_1638);
and U383 (N_383,In_1173,In_2171);
and U384 (N_384,In_2711,In_732);
xor U385 (N_385,In_409,In_1832);
nand U386 (N_386,In_1959,In_848);
and U387 (N_387,In_2724,In_1211);
and U388 (N_388,In_2180,In_1044);
xnor U389 (N_389,In_2706,In_2484);
nand U390 (N_390,In_1615,In_2147);
nor U391 (N_391,In_1182,In_2179);
or U392 (N_392,In_2479,In_2376);
nor U393 (N_393,In_277,In_1145);
nor U394 (N_394,In_2612,In_1977);
nor U395 (N_395,In_1559,In_1491);
nand U396 (N_396,In_521,In_104);
nor U397 (N_397,In_221,In_1533);
or U398 (N_398,In_744,In_1461);
xnor U399 (N_399,In_1970,In_83);
xor U400 (N_400,In_929,In_862);
or U401 (N_401,In_1577,In_376);
nor U402 (N_402,In_344,In_1562);
nor U403 (N_403,In_1369,In_584);
or U404 (N_404,In_1227,In_2620);
xnor U405 (N_405,In_1749,In_1751);
xor U406 (N_406,In_2802,In_1131);
and U407 (N_407,In_2812,In_1627);
and U408 (N_408,In_2975,In_53);
or U409 (N_409,In_435,In_1025);
xor U410 (N_410,In_2408,In_2586);
or U411 (N_411,In_2856,In_529);
and U412 (N_412,In_2941,In_2677);
and U413 (N_413,In_802,In_226);
nand U414 (N_414,In_644,In_2207);
nor U415 (N_415,In_493,In_1184);
and U416 (N_416,In_2072,In_209);
and U417 (N_417,In_2791,In_2933);
or U418 (N_418,In_276,In_1808);
or U419 (N_419,In_1110,In_868);
nand U420 (N_420,In_2377,In_294);
nand U421 (N_421,In_992,In_449);
nand U422 (N_422,In_127,In_1893);
xor U423 (N_423,In_1300,In_1746);
xnor U424 (N_424,In_1043,In_2360);
xor U425 (N_425,In_968,In_1332);
and U426 (N_426,In_2915,In_2458);
nor U427 (N_427,In_2799,In_1);
xor U428 (N_428,In_2865,In_197);
and U429 (N_429,In_2931,In_1718);
nor U430 (N_430,In_634,In_1126);
or U431 (N_431,In_171,In_1621);
nor U432 (N_432,In_1083,In_884);
and U433 (N_433,In_1213,In_1469);
or U434 (N_434,In_743,In_982);
or U435 (N_435,In_770,In_1382);
nor U436 (N_436,In_1023,In_2288);
xor U437 (N_437,In_85,In_2094);
or U438 (N_438,In_1572,In_495);
nor U439 (N_439,In_102,In_527);
nor U440 (N_440,In_969,In_1814);
or U441 (N_441,In_1059,In_1065);
or U442 (N_442,In_966,In_1648);
or U443 (N_443,In_2473,In_1381);
nand U444 (N_444,In_1828,In_777);
or U445 (N_445,In_1168,In_1728);
xnor U446 (N_446,In_1578,In_932);
nand U447 (N_447,In_1149,In_7);
nand U448 (N_448,In_807,In_1582);
or U449 (N_449,In_2976,In_990);
or U450 (N_450,In_2400,In_2045);
nand U451 (N_451,In_1862,In_1815);
or U452 (N_452,In_389,In_2099);
and U453 (N_453,In_1388,In_1804);
nor U454 (N_454,In_1119,In_2433);
and U455 (N_455,In_311,In_408);
nor U456 (N_456,In_653,In_2559);
or U457 (N_457,In_1350,In_1544);
or U458 (N_458,In_2152,In_134);
xnor U459 (N_459,In_1398,In_2971);
xnor U460 (N_460,In_1748,In_1829);
nand U461 (N_461,In_1488,In_90);
nor U462 (N_462,In_1310,In_875);
or U463 (N_463,In_340,In_1077);
xnor U464 (N_464,In_585,In_365);
and U465 (N_465,In_1340,In_272);
xnor U466 (N_466,In_850,In_632);
and U467 (N_467,In_856,In_1556);
nor U468 (N_468,In_1802,In_863);
nand U469 (N_469,In_836,In_747);
nand U470 (N_470,In_2246,In_2806);
or U471 (N_471,In_460,In_68);
or U472 (N_472,In_2992,In_2808);
or U473 (N_473,In_2785,In_2442);
and U474 (N_474,In_2119,In_1956);
xnor U475 (N_475,In_2889,In_2922);
nor U476 (N_476,In_1688,In_603);
nor U477 (N_477,In_2912,In_1738);
xnor U478 (N_478,In_2940,In_1246);
nor U479 (N_479,In_2747,In_878);
xnor U480 (N_480,In_942,In_452);
and U481 (N_481,In_2663,In_1773);
xnor U482 (N_482,In_1856,In_829);
nand U483 (N_483,In_1785,In_1428);
or U484 (N_484,In_48,In_1127);
nand U485 (N_485,In_2233,In_596);
or U486 (N_486,In_2257,In_2058);
xnor U487 (N_487,In_681,In_926);
and U488 (N_488,In_1733,In_1053);
and U489 (N_489,In_2813,In_1891);
nor U490 (N_490,In_2664,In_225);
nand U491 (N_491,In_773,In_287);
and U492 (N_492,In_2708,In_2307);
and U493 (N_493,In_1756,In_1132);
and U494 (N_494,In_309,In_1419);
nand U495 (N_495,In_400,In_2850);
and U496 (N_496,In_1788,In_1040);
nand U497 (N_497,In_1639,In_2122);
or U498 (N_498,In_2602,In_598);
or U499 (N_499,In_1056,In_656);
or U500 (N_500,In_1793,In_1499);
nor U501 (N_501,In_1591,In_1516);
or U502 (N_502,In_1767,In_1002);
or U503 (N_503,In_2090,In_241);
nor U504 (N_504,In_2265,In_1253);
xnor U505 (N_505,In_2632,In_2723);
nand U506 (N_506,In_2550,In_2786);
nand U507 (N_507,In_1495,In_1798);
and U508 (N_508,In_2173,In_2510);
nor U509 (N_509,In_2851,In_2763);
or U510 (N_510,In_1943,In_587);
xor U511 (N_511,In_2702,In_1859);
or U512 (N_512,In_2796,In_1968);
or U513 (N_513,In_1358,In_536);
and U514 (N_514,In_790,In_2631);
nor U515 (N_515,In_2611,In_640);
nand U516 (N_516,In_9,In_2512);
nor U517 (N_517,In_2499,In_1715);
nor U518 (N_518,In_950,In_2267);
nor U519 (N_519,In_139,In_1845);
nand U520 (N_520,In_206,In_1526);
nand U521 (N_521,In_956,In_786);
nor U522 (N_522,In_2413,In_2480);
and U523 (N_523,In_1172,In_1087);
nand U524 (N_524,In_466,In_1664);
nand U525 (N_525,In_2899,In_1684);
nand U526 (N_526,In_511,In_2725);
nand U527 (N_527,In_2461,In_1410);
xnor U528 (N_528,In_2676,In_525);
xor U529 (N_529,In_243,In_1262);
nand U530 (N_530,In_1571,In_1916);
and U531 (N_531,In_1338,In_2610);
xor U532 (N_532,In_1128,In_2917);
nor U533 (N_533,In_764,In_1195);
or U534 (N_534,In_2096,In_575);
xnor U535 (N_535,In_1498,In_1285);
nor U536 (N_536,In_2491,In_588);
or U537 (N_537,In_2960,In_2954);
and U538 (N_538,In_56,In_1656);
or U539 (N_539,In_1801,In_1305);
nor U540 (N_540,In_1318,In_1539);
xor U541 (N_541,In_1745,In_1686);
or U542 (N_542,In_1665,In_1331);
or U543 (N_543,In_837,In_2772);
nand U544 (N_544,In_1712,In_765);
or U545 (N_545,In_1768,In_2926);
or U546 (N_546,In_145,In_2505);
nand U547 (N_547,In_558,In_2883);
or U548 (N_548,In_1616,In_2857);
nand U549 (N_549,In_490,In_581);
xnor U550 (N_550,In_2792,In_2158);
or U551 (N_551,In_2938,In_2585);
or U552 (N_552,In_42,In_253);
nor U553 (N_553,In_2089,In_1228);
nor U554 (N_554,In_1150,In_1316);
xor U555 (N_555,In_2457,In_2280);
nand U556 (N_556,In_648,In_2195);
and U557 (N_557,In_2615,In_2348);
or U558 (N_558,In_177,In_785);
nor U559 (N_559,In_444,In_731);
and U560 (N_560,In_879,In_946);
and U561 (N_561,In_975,In_1084);
nand U562 (N_562,In_1057,In_445);
and U563 (N_563,In_2211,In_1550);
xnor U564 (N_564,In_686,In_2432);
and U565 (N_565,In_1470,In_1573);
xnor U566 (N_566,In_126,In_2184);
or U567 (N_567,In_710,In_157);
xnor U568 (N_568,In_395,In_2425);
and U569 (N_569,In_1907,In_2522);
xnor U570 (N_570,In_1511,In_655);
nor U571 (N_571,In_2314,In_2811);
or U572 (N_572,In_1833,In_1143);
or U573 (N_573,In_1399,In_40);
nand U574 (N_574,In_2318,In_1654);
xor U575 (N_575,In_431,In_1528);
and U576 (N_576,In_1292,In_796);
or U577 (N_577,In_1604,In_2832);
nor U578 (N_578,In_280,In_1971);
nand U579 (N_579,In_2733,In_2217);
nor U580 (N_580,In_2423,In_2968);
or U581 (N_581,In_1995,In_2868);
nor U582 (N_582,In_2112,In_355);
or U583 (N_583,In_1525,In_1876);
nor U584 (N_584,In_2697,In_2983);
nand U585 (N_585,In_1412,In_1401);
and U586 (N_586,In_1010,In_2732);
xnor U587 (N_587,In_2959,In_1248);
nand U588 (N_588,In_1367,In_2957);
nand U589 (N_589,In_213,In_2299);
nand U590 (N_590,In_210,In_2310);
and U591 (N_591,In_1403,In_1846);
xor U592 (N_592,In_1755,In_1842);
nand U593 (N_593,In_720,In_2053);
nand U594 (N_594,In_2182,In_1429);
nand U595 (N_595,In_110,In_1261);
and U596 (N_596,In_2607,In_1770);
nor U597 (N_597,In_2359,In_685);
nand U598 (N_598,In_2995,In_1739);
and U599 (N_599,In_1086,In_1270);
nand U600 (N_600,In_2821,In_1597);
nor U601 (N_601,In_1858,In_2862);
nand U602 (N_602,In_1677,In_2955);
xor U603 (N_603,In_633,In_428);
or U604 (N_604,In_533,In_2962);
xor U605 (N_605,In_2471,In_325);
nor U606 (N_606,In_379,In_920);
nor U607 (N_607,In_2894,In_2002);
nor U608 (N_608,In_239,In_1899);
nor U609 (N_609,In_2468,In_477);
and U610 (N_610,In_1957,In_1485);
nand U611 (N_611,In_2346,In_1447);
or U612 (N_612,In_2867,In_1941);
and U613 (N_613,In_1840,In_8);
and U614 (N_614,In_1831,In_1456);
nor U615 (N_615,In_1644,In_1116);
and U616 (N_616,In_2015,In_2793);
nand U617 (N_617,In_1998,In_2642);
and U618 (N_618,In_203,In_567);
nand U619 (N_619,In_2126,In_1807);
nand U620 (N_620,In_488,In_2778);
nand U621 (N_621,In_725,In_2580);
nand U622 (N_622,In_666,In_212);
nor U623 (N_623,In_305,In_985);
nand U624 (N_624,In_70,In_22);
nor U625 (N_625,In_1479,In_937);
nor U626 (N_626,In_1958,In_2592);
nor U627 (N_627,In_602,In_2737);
nor U628 (N_628,In_2151,In_2320);
nor U629 (N_629,In_775,In_755);
nor U630 (N_630,In_2932,In_1314);
xnor U631 (N_631,In_2498,In_2410);
xor U632 (N_632,In_1813,In_2172);
xnor U633 (N_633,In_791,In_1563);
and U634 (N_634,In_2986,In_1225);
nand U635 (N_635,In_19,In_2929);
xor U636 (N_636,In_1178,In_1203);
xor U637 (N_637,In_2441,In_550);
xor U638 (N_638,In_821,In_2519);
nand U639 (N_639,In_763,In_2154);
and U640 (N_640,In_1875,In_922);
nor U641 (N_641,In_443,In_716);
nand U642 (N_642,In_1586,In_489);
and U643 (N_643,In_1826,In_911);
nor U644 (N_644,In_2193,In_353);
and U645 (N_645,In_2927,In_566);
or U646 (N_646,In_759,In_853);
or U647 (N_647,In_1490,In_2901);
xor U648 (N_648,In_1177,In_954);
nor U649 (N_649,In_38,In_1426);
or U650 (N_650,In_702,In_1938);
xnor U651 (N_651,In_2573,In_689);
or U652 (N_652,In_2091,In_729);
xnor U653 (N_653,In_1019,In_1543);
nor U654 (N_654,In_1103,In_831);
or U655 (N_655,In_2656,In_304);
nand U656 (N_656,In_683,In_2381);
xor U657 (N_657,In_2101,In_1974);
nor U658 (N_658,In_149,In_2701);
and U659 (N_659,In_2009,In_1619);
nand U660 (N_660,In_1238,In_1778);
and U661 (N_661,In_538,In_2673);
and U662 (N_662,In_2032,In_332);
xor U663 (N_663,In_2621,In_851);
nor U664 (N_664,In_2238,In_2243);
and U665 (N_665,In_2762,In_2703);
xnor U666 (N_666,In_2981,In_1819);
xor U667 (N_667,In_1626,In_491);
nor U668 (N_668,In_32,In_20);
xor U669 (N_669,In_1857,In_989);
or U670 (N_670,In_677,In_678);
nand U671 (N_671,In_2655,In_1741);
xor U672 (N_672,In_2284,In_1205);
or U673 (N_673,In_2225,In_214);
nor U674 (N_674,In_2214,In_2537);
xnor U675 (N_675,In_1460,In_2160);
xnor U676 (N_676,In_1268,In_1070);
and U677 (N_677,In_310,In_189);
or U678 (N_678,In_328,In_509);
or U679 (N_679,In_624,In_2362);
nand U680 (N_680,In_630,In_1960);
xor U681 (N_681,In_983,In_343);
nand U682 (N_682,In_1496,In_2076);
nor U683 (N_683,In_1237,In_893);
nor U684 (N_684,In_2055,In_2256);
and U685 (N_685,In_469,In_2117);
nor U686 (N_686,In_1450,In_1537);
xor U687 (N_687,In_2463,In_1514);
nand U688 (N_688,In_1930,In_1710);
or U689 (N_689,In_2742,In_1593);
or U690 (N_690,In_2178,In_2436);
nor U691 (N_691,In_498,In_1873);
and U692 (N_692,In_905,In_721);
or U693 (N_693,In_1620,In_1894);
or U694 (N_694,In_594,In_1874);
and U695 (N_695,In_1006,In_970);
or U696 (N_696,In_2311,In_1866);
and U697 (N_697,In_2928,In_1786);
and U698 (N_698,In_1761,In_2693);
and U699 (N_699,In_2475,In_2948);
or U700 (N_700,In_1400,In_2717);
or U701 (N_701,In_965,In_207);
xor U702 (N_702,In_2222,In_1427);
nand U703 (N_703,In_819,In_2291);
or U704 (N_704,In_1368,In_944);
xnor U705 (N_705,In_282,In_99);
nor U706 (N_706,In_921,In_939);
and U707 (N_707,In_2323,In_2597);
xnor U708 (N_708,In_380,In_2532);
or U709 (N_709,In_547,In_591);
nand U710 (N_710,In_1390,In_2252);
or U711 (N_711,In_918,In_680);
nor U712 (N_712,In_1524,In_186);
nor U713 (N_713,In_420,In_1662);
xor U714 (N_714,In_286,In_825);
or U715 (N_715,In_2028,In_2982);
or U716 (N_716,In_2030,In_2781);
or U717 (N_717,In_768,In_2910);
or U718 (N_718,In_2903,In_366);
and U719 (N_719,In_2132,In_2197);
xnor U720 (N_720,In_1727,In_2190);
or U721 (N_721,In_738,In_578);
xor U722 (N_722,In_1611,In_528);
and U723 (N_723,In_834,In_2988);
nand U724 (N_724,In_1125,In_563);
nor U725 (N_725,In_1791,In_2235);
xor U726 (N_726,In_1280,In_2303);
or U727 (N_727,In_198,In_1295);
nor U728 (N_728,In_1612,In_1473);
nor U729 (N_729,In_1650,In_501);
xnor U730 (N_730,In_549,In_887);
nand U731 (N_731,In_1308,In_1165);
and U732 (N_732,In_772,In_2967);
nand U733 (N_733,In_1510,In_2088);
xor U734 (N_734,In_867,In_610);
xor U735 (N_735,In_1976,In_437);
xnor U736 (N_736,In_1438,In_1641);
xnor U737 (N_737,In_1809,In_1030);
xnor U738 (N_738,In_2963,In_223);
nand U739 (N_739,In_1816,In_111);
nor U740 (N_740,In_2828,In_2077);
xor U741 (N_741,In_446,In_1504);
and U742 (N_742,In_1682,In_275);
or U743 (N_743,In_1513,In_2095);
xnor U744 (N_744,In_1468,In_2874);
or U745 (N_745,In_211,In_2794);
xor U746 (N_746,In_293,In_423);
xnor U747 (N_747,In_430,In_573);
and U748 (N_748,In_1406,In_163);
nand U749 (N_749,In_552,In_1106);
xnor U750 (N_750,In_1154,In_695);
xnor U751 (N_751,In_2005,In_2882);
nor U752 (N_752,In_540,In_222);
or U753 (N_753,In_1218,In_2966);
or U754 (N_754,In_1883,In_2467);
nand U755 (N_755,In_1554,In_1661);
nand U756 (N_756,In_506,In_345);
and U757 (N_757,In_2810,In_977);
or U758 (N_758,In_2715,In_510);
and U759 (N_759,In_742,In_783);
nor U760 (N_760,In_1046,In_1483);
nor U761 (N_761,In_923,In_1982);
nor U762 (N_762,In_1175,In_1924);
nand U763 (N_763,In_1167,In_401);
nor U764 (N_764,In_183,In_2569);
nand U765 (N_765,In_2958,In_378);
and U766 (N_766,In_2213,In_771);
nor U767 (N_767,In_2129,In_1944);
and U768 (N_768,In_504,In_1492);
nand U769 (N_769,In_16,In_1417);
xnor U770 (N_770,In_2689,In_2066);
or U771 (N_771,In_1022,In_1459);
nor U772 (N_772,In_2892,In_1865);
nor U773 (N_773,In_2761,In_1007);
xor U774 (N_774,In_1042,In_65);
or U775 (N_775,In_346,In_368);
nand U776 (N_776,In_351,In_1341);
nor U777 (N_777,In_1163,In_1864);
xor U778 (N_778,In_801,In_426);
nor U779 (N_779,In_2616,In_2989);
nand U780 (N_780,In_930,In_2153);
nor U781 (N_781,In_1521,In_2052);
and U782 (N_782,In_284,In_2039);
nor U783 (N_783,In_2779,In_2574);
or U784 (N_784,In_931,In_470);
nand U785 (N_785,In_854,In_883);
nor U786 (N_786,In_12,In_524);
nor U787 (N_787,In_2700,In_2625);
xnor U788 (N_788,In_2272,In_496);
or U789 (N_789,In_1771,In_146);
xor U790 (N_790,In_403,In_1487);
nor U791 (N_791,In_650,In_1588);
and U792 (N_792,In_1506,In_2730);
nand U793 (N_793,In_973,In_2127);
nand U794 (N_794,In_381,In_2918);
xor U795 (N_795,In_1734,In_2051);
xor U796 (N_796,In_1121,In_1197);
nor U797 (N_797,In_576,In_1766);
and U798 (N_798,In_1869,In_1151);
nand U799 (N_799,In_2695,In_2965);
or U800 (N_800,In_2852,In_1878);
nor U801 (N_801,In_1694,In_2137);
nand U802 (N_802,In_1047,In_290);
xor U803 (N_803,In_457,In_1180);
nand U804 (N_804,In_2086,In_2449);
nand U805 (N_805,In_1784,In_147);
or U806 (N_806,In_1200,In_2397);
xnor U807 (N_807,In_1061,In_112);
and U808 (N_808,In_55,In_2041);
nand U809 (N_809,In_2327,In_2731);
xor U810 (N_810,In_1365,In_419);
and U811 (N_811,In_1762,In_2276);
nand U812 (N_812,In_2543,In_1393);
nor U813 (N_813,In_1171,In_137);
xor U814 (N_814,In_2420,In_1655);
and U815 (N_815,In_2861,In_2080);
nand U816 (N_816,In_2996,In_1936);
nand U817 (N_817,In_281,In_179);
nand U818 (N_818,In_1529,In_1048);
or U819 (N_819,In_1206,In_1441);
nor U820 (N_820,In_2004,In_87);
nor U821 (N_821,In_341,In_124);
and U822 (N_822,In_2060,In_2048);
nand U823 (N_823,In_175,In_1613);
nand U824 (N_824,In_2412,In_2878);
and U825 (N_825,In_1001,In_499);
or U826 (N_826,In_2606,In_1434);
nor U827 (N_827,In_383,In_2583);
nor U828 (N_828,In_1950,In_604);
and U829 (N_829,In_1834,In_1910);
xor U830 (N_830,In_153,In_737);
nor U831 (N_831,In_1394,In_502);
and U832 (N_832,In_1700,In_130);
nor U833 (N_833,In_2764,In_707);
nand U834 (N_834,In_2603,In_871);
nor U835 (N_835,In_1806,In_2524);
xnor U836 (N_836,In_649,In_2194);
or U837 (N_837,In_728,In_1632);
and U838 (N_838,In_2831,In_2584);
or U839 (N_839,In_2626,In_360);
or U840 (N_840,In_994,In_1912);
nand U841 (N_841,In_1868,In_1123);
and U842 (N_842,In_1668,In_2084);
nand U843 (N_843,In_1986,In_545);
or U844 (N_844,In_1050,In_2558);
or U845 (N_845,In_300,In_2364);
and U846 (N_846,In_1494,In_1634);
nor U847 (N_847,In_544,In_1902);
nand U848 (N_848,In_1797,In_715);
xor U849 (N_849,In_1607,In_1326);
and U850 (N_850,In_1933,In_2455);
and U851 (N_851,In_2833,In_1942);
or U852 (N_852,In_1476,In_2713);
nor U853 (N_853,In_1416,In_2249);
xnor U854 (N_854,In_2204,In_2890);
or U855 (N_855,In_2219,In_1882);
xnor U856 (N_856,In_399,In_2775);
xnor U857 (N_857,In_2459,In_1697);
nor U858 (N_858,In_2690,In_1094);
xor U859 (N_859,In_1405,In_1062);
nand U860 (N_860,In_2373,In_1273);
nand U861 (N_861,In_2630,In_1222);
xnor U862 (N_862,In_1144,In_5);
xor U863 (N_863,In_158,In_2688);
xor U864 (N_864,In_1716,In_2914);
or U865 (N_865,In_2609,In_2999);
nor U866 (N_866,In_2341,In_1646);
and U867 (N_867,In_295,In_872);
or U868 (N_868,In_2042,In_11);
or U869 (N_869,In_1692,In_2345);
nand U870 (N_870,In_2835,In_2773);
xor U871 (N_871,In_2437,In_2554);
nor U872 (N_872,In_1038,In_565);
xnor U873 (N_873,In_274,In_2503);
and U874 (N_874,In_2547,In_2146);
nor U875 (N_875,In_2446,In_432);
xor U876 (N_876,In_1993,In_1446);
xor U877 (N_877,In_1954,In_1235);
or U878 (N_878,In_557,In_1230);
nand U879 (N_879,In_1781,In_1835);
nand U880 (N_880,In_2599,In_2226);
xnor U881 (N_881,In_1169,In_2752);
xnor U882 (N_882,In_1484,In_2188);
nand U883 (N_883,In_2837,In_1541);
nand U884 (N_884,In_1900,In_2774);
and U885 (N_885,In_135,In_2264);
or U886 (N_886,In_2445,In_735);
nand U887 (N_887,In_2417,In_129);
nand U888 (N_888,In_2881,In_1288);
and U889 (N_889,In_2477,In_2176);
nand U890 (N_890,In_2520,In_336);
nand U891 (N_891,In_2356,In_181);
or U892 (N_892,In_2451,In_2820);
and U893 (N_893,In_79,In_2006);
and U894 (N_894,In_1997,In_888);
xor U895 (N_895,In_1174,In_1389);
or U896 (N_896,In_303,In_2873);
nor U897 (N_897,In_519,In_2426);
xnor U898 (N_898,In_257,In_2021);
nor U899 (N_899,In_1689,In_10);
or U900 (N_900,In_2145,In_543);
nand U901 (N_901,In_1678,In_141);
or U902 (N_902,In_1729,In_676);
or U903 (N_903,In_2443,In_2496);
xor U904 (N_904,In_28,In_2738);
xnor U905 (N_905,In_1424,In_1413);
or U906 (N_906,In_2333,In_450);
nand U907 (N_907,In_2465,In_2258);
nor U908 (N_908,In_1780,In_2872);
and U909 (N_909,In_1625,In_497);
or U910 (N_910,In_1141,In_382);
or U911 (N_911,In_2047,In_2301);
xor U912 (N_912,In_1517,In_1824);
nor U913 (N_913,In_2135,In_1929);
nor U914 (N_914,In_427,In_1204);
nor U915 (N_915,In_1449,In_358);
nor U916 (N_916,In_306,In_1754);
xor U917 (N_917,In_21,In_1378);
xor U918 (N_918,In_2108,In_125);
nor U919 (N_919,In_494,In_71);
nand U920 (N_920,In_1990,In_292);
or U921 (N_921,In_2698,In_229);
nand U922 (N_922,In_337,In_2546);
xnor U923 (N_923,In_100,In_1254);
nor U924 (N_924,In_2384,In_82);
nor U925 (N_925,In_37,In_2050);
nand U926 (N_926,In_434,In_916);
or U927 (N_927,In_2330,In_645);
nand U928 (N_928,In_2511,In_1052);
or U929 (N_929,In_2250,In_76);
or U930 (N_930,In_2141,In_1415);
nor U931 (N_931,In_2847,In_454);
and U932 (N_932,In_2754,In_472);
nand U933 (N_933,In_1992,In_1290);
and U934 (N_934,In_2947,In_2565);
nand U935 (N_935,In_1699,In_1435);
nor U936 (N_936,In_1301,In_1372);
nor U937 (N_937,In_185,In_1991);
xnor U938 (N_938,In_894,In_215);
and U939 (N_939,In_2668,In_991);
and U940 (N_940,In_1701,In_1414);
and U941 (N_941,In_2201,In_586);
xnor U942 (N_942,In_2065,In_2230);
and U943 (N_943,In_2556,In_359);
xor U944 (N_944,In_1034,In_2815);
nor U945 (N_945,In_2665,In_2727);
or U946 (N_946,In_833,In_2271);
and U947 (N_947,In_1142,In_169);
xor U948 (N_948,In_97,In_60);
and U949 (N_949,In_2419,In_1898);
nand U950 (N_950,In_2669,In_1649);
xor U951 (N_951,In_174,In_2925);
xor U952 (N_952,In_1241,In_2049);
nor U953 (N_953,In_106,In_133);
nand U954 (N_954,In_1546,In_1303);
or U955 (N_955,In_406,In_2337);
or U956 (N_956,In_2036,In_2157);
nand U957 (N_957,In_302,In_2444);
xor U958 (N_958,In_2809,In_301);
xnor U959 (N_959,In_1244,In_1841);
or U960 (N_960,In_1881,In_899);
and U961 (N_961,In_2640,In_1430);
nand U962 (N_962,In_2638,In_1690);
nor U963 (N_963,In_2896,In_1448);
and U964 (N_964,In_2022,In_84);
and U965 (N_965,In_388,In_1148);
xnor U966 (N_966,In_822,In_2024);
and U967 (N_967,In_103,In_660);
xnor U968 (N_968,In_244,In_2027);
xnor U969 (N_969,In_1157,In_505);
and U970 (N_970,In_176,In_2270);
nand U971 (N_971,In_324,In_327);
nor U972 (N_972,In_2308,In_88);
and U973 (N_973,In_2902,In_1467);
nor U974 (N_974,In_2770,In_758);
nor U975 (N_975,In_1714,In_1810);
or U976 (N_976,In_2758,In_1764);
nand U977 (N_977,In_1219,In_1109);
nor U978 (N_978,In_1679,In_730);
nand U979 (N_979,In_2596,In_1036);
xnor U980 (N_980,In_827,In_1220);
nand U981 (N_981,In_172,In_2870);
nor U982 (N_982,In_840,In_1567);
or U983 (N_983,In_49,In_138);
and U984 (N_984,In_909,In_326);
xor U985 (N_985,In_1000,In_2168);
nor U986 (N_986,In_1927,In_393);
or U987 (N_987,In_160,In_1224);
or U988 (N_988,In_1935,In_1631);
nor U989 (N_989,In_2623,In_1092);
nor U990 (N_990,In_2023,In_1792);
or U991 (N_991,In_2652,In_1188);
nor U992 (N_992,In_1763,In_465);
nand U993 (N_993,In_2994,In_880);
xor U994 (N_994,In_2750,In_2306);
nor U995 (N_995,In_2842,In_2269);
xnor U996 (N_996,In_2540,In_1039);
and U997 (N_997,In_34,In_798);
and U998 (N_998,In_17,In_734);
nor U999 (N_999,In_2078,In_1730);
nor U1000 (N_1000,In_839,In_2884);
nor U1001 (N_1001,In_1296,In_1914);
nor U1002 (N_1002,In_2950,In_291);
nand U1003 (N_1003,In_2133,In_611);
or U1004 (N_1004,In_776,In_2571);
nor U1005 (N_1005,In_661,In_1436);
xor U1006 (N_1006,In_1115,In_237);
and U1007 (N_1007,In_2907,In_279);
or U1008 (N_1008,In_73,In_904);
and U1009 (N_1009,In_2657,In_1722);
nand U1010 (N_1010,In_2223,In_1505);
xor U1011 (N_1011,In_1029,In_398);
or U1012 (N_1012,In_2647,In_823);
and U1013 (N_1013,In_1380,In_1847);
nor U1014 (N_1014,In_2720,In_535);
or U1015 (N_1015,In_2411,In_1681);
xor U1016 (N_1016,In_1606,In_461);
or U1017 (N_1017,In_458,In_2829);
xor U1018 (N_1018,In_1190,In_2013);
nand U1019 (N_1019,In_2297,In_1012);
nand U1020 (N_1020,In_2391,In_2570);
nand U1021 (N_1021,In_2780,In_1596);
nor U1022 (N_1022,In_199,In_1386);
nand U1023 (N_1023,In_817,In_1849);
nor U1024 (N_1024,In_252,In_2666);
and U1025 (N_1025,In_377,In_480);
nand U1026 (N_1026,In_1361,In_1395);
and U1027 (N_1027,In_2594,In_2953);
xnor U1028 (N_1028,In_2123,In_1334);
nor U1029 (N_1029,In_2139,In_2681);
nand U1030 (N_1030,In_2921,In_1602);
or U1031 (N_1031,In_1670,In_2401);
nand U1032 (N_1032,In_372,In_1348);
and U1033 (N_1033,In_1079,In_2253);
nand U1034 (N_1034,In_142,In_1104);
nand U1035 (N_1035,In_2617,In_2553);
nand U1036 (N_1036,In_701,In_2687);
and U1037 (N_1037,In_2251,In_2716);
and U1038 (N_1038,In_1216,In_27);
nor U1039 (N_1039,In_745,In_1645);
xor U1040 (N_1040,In_1231,In_722);
and U1041 (N_1041,In_1794,In_2403);
and U1042 (N_1042,In_1232,In_1362);
nand U1043 (N_1043,In_2803,In_1377);
or U1044 (N_1044,In_541,In_927);
nor U1045 (N_1045,In_1311,In_2563);
xor U1046 (N_1046,In_2386,In_1568);
nand U1047 (N_1047,In_2093,In_2260);
nor U1048 (N_1048,In_0,In_1482);
and U1049 (N_1049,In_2290,In_749);
and U1050 (N_1050,In_425,In_2371);
and U1051 (N_1051,In_1315,In_2536);
and U1052 (N_1052,In_64,In_1324);
xor U1053 (N_1053,In_2578,In_1444);
and U1054 (N_1054,In_2113,In_2840);
nand U1055 (N_1055,In_202,In_1333);
nor U1056 (N_1056,In_2392,In_2165);
or U1057 (N_1057,In_1913,In_2008);
xnor U1058 (N_1058,In_1028,In_235);
and U1059 (N_1059,In_1355,In_271);
nand U1060 (N_1060,In_2069,In_2244);
xor U1061 (N_1061,In_1702,In_2143);
nand U1062 (N_1062,In_2904,In_2590);
xnor U1063 (N_1063,In_555,In_2210);
xor U1064 (N_1064,In_800,In_170);
or U1065 (N_1065,In_654,In_1880);
xnor U1066 (N_1066,In_2115,In_1903);
nor U1067 (N_1067,In_2382,In_814);
xor U1068 (N_1068,In_2228,In_2186);
nand U1069 (N_1069,In_1016,In_1965);
nand U1070 (N_1070,In_832,In_473);
and U1071 (N_1071,In_2424,In_30);
xor U1072 (N_1072,In_2822,In_1618);
nor U1073 (N_1073,In_2285,In_261);
and U1074 (N_1074,In_690,In_1884);
xnor U1075 (N_1075,In_651,In_2854);
nor U1076 (N_1076,In_1653,In_1737);
nand U1077 (N_1077,In_2826,In_46);
and U1078 (N_1078,In_637,In_866);
nor U1079 (N_1079,In_670,In_2721);
nand U1080 (N_1080,In_270,In_643);
or U1081 (N_1081,In_1666,In_706);
xnor U1082 (N_1082,In_910,In_1357);
xor U1083 (N_1083,In_1844,In_843);
or U1084 (N_1084,In_1064,In_1321);
xnor U1085 (N_1085,In_2572,In_1515);
xnor U1086 (N_1086,In_289,In_876);
or U1087 (N_1087,In_2125,In_1093);
nand U1088 (N_1088,In_1723,In_1443);
nor U1089 (N_1089,In_371,In_2447);
nor U1090 (N_1090,In_1635,In_2935);
nand U1091 (N_1091,In_1015,In_204);
and U1092 (N_1092,In_2,In_1069);
xor U1093 (N_1093,In_59,In_2393);
or U1094 (N_1094,In_805,In_964);
and U1095 (N_1095,In_1249,In_2521);
nor U1096 (N_1096,In_2262,In_1345);
and U1097 (N_1097,In_2259,In_2304);
xor U1098 (N_1098,In_1975,In_718);
or U1099 (N_1099,In_769,In_2192);
xor U1100 (N_1100,In_1890,In_756);
xor U1101 (N_1101,In_2389,In_2162);
and U1102 (N_1102,In_233,In_474);
xnor U1103 (N_1103,In_2535,In_299);
nor U1104 (N_1104,In_2100,In_1871);
xnor U1105 (N_1105,In_1760,In_958);
xnor U1106 (N_1106,In_2804,In_23);
or U1107 (N_1107,In_2787,In_1931);
nor U1108 (N_1108,In_1530,In_347);
or U1109 (N_1109,In_1478,In_967);
or U1110 (N_1110,In_1895,In_2368);
or U1111 (N_1111,In_760,In_459);
nand U1112 (N_1112,In_972,In_2908);
xor U1113 (N_1113,In_1277,In_1726);
and U1114 (N_1114,In_1905,In_1027);
xnor U1115 (N_1115,In_1676,In_613);
or U1116 (N_1116,In_2261,In_1464);
and U1117 (N_1117,In_122,In_2523);
or U1118 (N_1118,In_2056,In_1159);
nor U1119 (N_1119,In_2469,In_2279);
nand U1120 (N_1120,In_2670,In_2483);
nor U1121 (N_1121,In_2577,In_2321);
nor U1122 (N_1122,In_951,In_1818);
and U1123 (N_1123,In_1925,In_2043);
or U1124 (N_1124,In_696,In_1067);
xor U1125 (N_1125,In_1508,In_2528);
or U1126 (N_1126,In_658,In_2807);
nor U1127 (N_1127,In_194,In_1923);
nand U1128 (N_1128,In_2736,In_1908);
xor U1129 (N_1129,In_260,In_349);
and U1130 (N_1130,In_1854,In_647);
nor U1131 (N_1131,In_2068,In_605);
nand U1132 (N_1132,In_1817,In_531);
and U1133 (N_1133,In_2644,In_1724);
or U1134 (N_1134,In_2946,In_2879);
xor U1135 (N_1135,In_2334,In_1071);
nor U1136 (N_1136,In_2352,In_247);
xnor U1137 (N_1137,In_952,In_1772);
and U1138 (N_1138,In_2961,In_191);
nand U1139 (N_1139,In_464,In_1920);
xnor U1140 (N_1140,In_2591,In_2795);
and U1141 (N_1141,In_2937,In_1836);
nand U1142 (N_1142,In_2956,In_2044);
nor U1143 (N_1143,In_593,In_2074);
nor U1144 (N_1144,In_154,In_766);
or U1145 (N_1145,In_595,In_81);
nand U1146 (N_1146,In_2177,In_436);
nor U1147 (N_1147,In_364,In_2038);
xnor U1148 (N_1148,In_2885,In_2029);
or U1149 (N_1149,In_109,In_333);
nand U1150 (N_1150,In_1962,In_2789);
or U1151 (N_1151,In_2281,In_1005);
nor U1152 (N_1152,In_724,In_148);
and U1153 (N_1153,In_978,In_1918);
nor U1154 (N_1154,In_2662,In_816);
xor U1155 (N_1155,In_1996,In_953);
nor U1156 (N_1156,In_2286,In_1838);
and U1157 (N_1157,In_1187,In_1707);
and U1158 (N_1158,In_699,In_1226);
xnor U1159 (N_1159,In_2358,In_2627);
nand U1160 (N_1160,In_2169,In_1385);
nand U1161 (N_1161,In_636,In_2343);
and U1162 (N_1162,In_625,In_2020);
nand U1163 (N_1163,In_1293,In_1432);
and U1164 (N_1164,In_617,In_1973);
or U1165 (N_1165,In_2991,In_534);
and U1166 (N_1166,In_314,In_159);
or U1167 (N_1167,In_2342,In_1489);
nor U1168 (N_1168,In_2245,In_614);
nand U1169 (N_1169,In_2860,In_882);
xnor U1170 (N_1170,In_1267,In_986);
xnor U1171 (N_1171,In_1789,In_1352);
xor U1172 (N_1172,In_1243,In_1628);
and U1173 (N_1173,In_438,In_532);
or U1174 (N_1174,In_2755,In_1695);
and U1175 (N_1175,In_2385,In_14);
or U1176 (N_1176,In_471,In_1663);
xor U1177 (N_1177,In_467,In_2790);
nor U1178 (N_1178,In_719,In_961);
nor U1179 (N_1179,In_2541,In_1373);
nor U1180 (N_1180,In_2396,In_2909);
or U1181 (N_1181,In_1872,In_859);
nand U1182 (N_1182,In_2660,In_1445);
nor U1183 (N_1183,In_517,In_1371);
nand U1184 (N_1184,In_1063,In_86);
xnor U1185 (N_1185,In_219,In_2605);
nand U1186 (N_1186,In_2943,In_2749);
or U1187 (N_1187,In_2274,In_1917);
and U1188 (N_1188,In_1518,In_1617);
and U1189 (N_1189,In_1497,In_1538);
nand U1190 (N_1190,In_2636,In_1397);
or U1191 (N_1191,In_1033,In_1317);
or U1192 (N_1192,In_629,In_569);
and U1193 (N_1193,In_2000,In_1685);
xor U1194 (N_1194,In_2454,In_1820);
or U1195 (N_1195,In_2548,In_2823);
nor U1196 (N_1196,In_2351,In_1422);
xor U1197 (N_1197,In_2059,In_1099);
and U1198 (N_1198,In_638,In_2923);
nand U1199 (N_1199,In_2331,In_826);
nand U1200 (N_1200,In_1889,In_849);
and U1201 (N_1201,In_468,In_2685);
and U1202 (N_1202,In_331,In_1323);
and U1203 (N_1203,In_105,In_1407);
or U1204 (N_1204,In_523,In_1257);
or U1205 (N_1205,In_639,In_1614);
nor U1206 (N_1206,In_155,In_1051);
or U1207 (N_1207,In_1477,In_971);
nor U1208 (N_1208,In_2628,In_847);
xor U1209 (N_1209,In_1387,In_1313);
and U1210 (N_1210,In_1642,In_2579);
xor U1211 (N_1211,In_513,In_2344);
nor U1212 (N_1212,In_1984,In_741);
or U1213 (N_1213,In_2744,In_865);
and U1214 (N_1214,In_62,In_2614);
and U1215 (N_1215,In_2001,In_727);
or U1216 (N_1216,In_1421,In_1752);
and U1217 (N_1217,In_915,In_2302);
nor U1218 (N_1218,In_548,In_1153);
nor U1219 (N_1219,In_1196,In_2608);
nand U1220 (N_1220,In_659,In_559);
nor U1221 (N_1221,In_245,In_844);
and U1222 (N_1222,In_89,In_387);
and U1223 (N_1223,In_933,In_2418);
or U1224 (N_1224,In_475,In_949);
nor U1225 (N_1225,In_631,In_1221);
nor U1226 (N_1226,In_627,In_92);
xnor U1227 (N_1227,In_2324,In_2843);
and U1228 (N_1228,In_1251,In_864);
nor U1229 (N_1229,In_397,In_1179);
xor U1230 (N_1230,In_217,In_1152);
or U1231 (N_1231,In_2534,In_1519);
nor U1232 (N_1232,In_2839,In_842);
xnor U1233 (N_1233,In_1396,In_91);
and U1234 (N_1234,In_2369,In_238);
xnor U1235 (N_1235,In_1327,In_577);
nand U1236 (N_1236,In_1553,In_2339);
nand U1237 (N_1237,In_2704,In_1068);
nand U1238 (N_1238,In_838,In_1643);
nand U1239 (N_1239,In_2237,In_2107);
nand U1240 (N_1240,In_987,In_820);
or U1241 (N_1241,In_2434,In_1531);
or U1242 (N_1242,In_479,In_2215);
nor U1243 (N_1243,In_242,In_2589);
nand U1244 (N_1244,In_898,In_1102);
or U1245 (N_1245,In_1240,In_335);
and U1246 (N_1246,In_456,In_2012);
and U1247 (N_1247,In_1587,In_1366);
or U1248 (N_1248,In_15,In_711);
and U1249 (N_1249,In_2709,In_150);
nand U1250 (N_1250,In_955,In_520);
and U1251 (N_1251,In_781,In_1579);
and U1252 (N_1252,In_2305,In_943);
xor U1253 (N_1253,In_2897,In_2978);
and U1254 (N_1254,In_935,In_356);
or U1255 (N_1255,In_2248,In_2159);
and U1256 (N_1256,In_2834,In_278);
xor U1257 (N_1257,In_3,In_2136);
nor U1258 (N_1258,In_265,In_2255);
xnor U1259 (N_1259,In_2329,In_1669);
and U1260 (N_1260,In_642,In_2944);
and U1261 (N_1261,In_693,In_144);
or U1262 (N_1262,In_2526,In_2198);
nand U1263 (N_1263,In_1354,In_2390);
xnor U1264 (N_1264,In_2913,In_1383);
xor U1265 (N_1265,In_1985,In_564);
and U1266 (N_1266,In_914,In_1735);
and U1267 (N_1267,In_1471,In_861);
or U1268 (N_1268,In_1208,In_919);
nand U1269 (N_1269,In_2765,In_1870);
or U1270 (N_1270,In_2951,In_1949);
xnor U1271 (N_1271,In_2818,In_448);
or U1272 (N_1272,In_1080,In_824);
nor U1273 (N_1273,In_906,In_2439);
nand U1274 (N_1274,In_806,In_1909);
nor U1275 (N_1275,In_288,In_778);
xor U1276 (N_1276,In_1081,In_192);
nor U1277 (N_1277,In_2658,In_2156);
nand U1278 (N_1278,In_1660,In_24);
or U1279 (N_1279,In_2661,In_385);
xor U1280 (N_1280,In_120,In_1342);
and U1281 (N_1281,In_2387,In_230);
nand U1282 (N_1282,In_1239,In_1360);
and U1283 (N_1283,In_995,In_704);
nor U1284 (N_1284,In_1343,In_485);
and U1285 (N_1285,In_646,In_619);
xnor U1286 (N_1286,In_94,In_2977);
nor U1287 (N_1287,In_2759,In_1946);
nand U1288 (N_1288,In_554,In_50);
and U1289 (N_1289,In_2203,In_1098);
nand U1290 (N_1290,In_1072,In_1105);
and U1291 (N_1291,In_2130,In_928);
and U1292 (N_1292,In_962,In_392);
or U1293 (N_1293,In_2017,In_2482);
and U1294 (N_1294,In_1176,In_268);
xor U1295 (N_1295,In_1003,In_2370);
nor U1296 (N_1296,In_694,In_2416);
nand U1297 (N_1297,In_1346,In_1708);
nand U1298 (N_1298,In_2587,In_835);
or U1299 (N_1299,In_1009,In_1166);
nor U1300 (N_1300,In_2181,In_2409);
nor U1301 (N_1301,In_2298,In_1953);
nor U1302 (N_1302,In_2844,In_1404);
or U1303 (N_1303,In_31,In_113);
xnor U1304 (N_1304,In_1101,In_2604);
nor U1305 (N_1305,In_36,In_44);
and U1306 (N_1306,In_901,In_997);
nor U1307 (N_1307,In_218,In_2916);
and U1308 (N_1308,In_2087,In_2650);
and U1309 (N_1309,In_2229,In_162);
and U1310 (N_1310,In_2309,In_2551);
nor U1311 (N_1311,In_782,In_240);
nor U1312 (N_1312,In_1967,In_1867);
nand U1313 (N_1313,In_1140,In_794);
nor U1314 (N_1314,In_1136,In_1821);
or U1315 (N_1315,In_61,In_1134);
or U1316 (N_1316,In_273,In_757);
and U1317 (N_1317,In_748,In_2054);
nor U1318 (N_1318,In_530,In_1886);
nand U1319 (N_1319,In_1799,In_1351);
xnor U1320 (N_1320,In_902,In_988);
or U1321 (N_1321,In_107,In_455);
xnor U1322 (N_1322,In_1731,In_652);
or U1323 (N_1323,In_1107,In_1194);
xnor U1324 (N_1324,In_2098,In_2399);
and U1325 (N_1325,In_996,In_298);
xor U1326 (N_1326,In_2208,In_416);
or U1327 (N_1327,In_1595,In_1659);
nor U1328 (N_1328,In_193,In_2855);
and U1329 (N_1329,In_2516,In_447);
xor U1330 (N_1330,In_739,In_1298);
nor U1331 (N_1331,In_2801,In_664);
xor U1332 (N_1332,In_75,In_1284);
nor U1333 (N_1333,In_18,In_1252);
and U1334 (N_1334,In_2174,In_283);
xor U1335 (N_1335,In_522,In_895);
nand U1336 (N_1336,In_1549,In_1601);
and U1337 (N_1337,In_2598,In_1651);
or U1338 (N_1338,In_1522,In_330);
nor U1339 (N_1339,In_2472,In_1442);
xor U1340 (N_1340,In_2557,In_57);
nor U1341 (N_1341,In_2033,In_266);
nor U1342 (N_1342,In_2888,In_312);
or U1343 (N_1343,In_25,In_1691);
and U1344 (N_1344,In_1711,In_2322);
nor U1345 (N_1345,In_2275,In_2149);
xnor U1346 (N_1346,In_924,In_390);
nor U1347 (N_1347,In_940,In_1557);
nor U1348 (N_1348,In_1673,In_1547);
nor U1349 (N_1349,In_1420,In_1297);
nand U1350 (N_1350,In_2502,In_1709);
or U1351 (N_1351,In_1130,In_2974);
nor U1352 (N_1352,In_852,In_116);
nand U1353 (N_1353,In_1919,In_1580);
nor U1354 (N_1354,In_1706,In_429);
nand U1355 (N_1355,In_1198,In_1271);
nor U1356 (N_1356,In_1463,In_190);
or U1357 (N_1357,In_761,In_2743);
xor U1358 (N_1358,In_2509,In_1364);
or U1359 (N_1359,In_1719,In_945);
or U1360 (N_1360,In_140,In_1532);
nor U1361 (N_1361,In_2063,In_476);
and U1362 (N_1362,In_1592,In_482);
or U1363 (N_1363,In_2997,In_1133);
and U1364 (N_1364,In_1987,In_1274);
nor U1365 (N_1365,In_2939,In_2998);
xnor U1366 (N_1366,In_687,In_1623);
xor U1367 (N_1367,In_2919,In_256);
nand U1368 (N_1368,In_45,In_1750);
or U1369 (N_1369,In_792,In_248);
nor U1370 (N_1370,In_2372,In_1743);
or U1371 (N_1371,In_2374,In_2600);
xor U1372 (N_1372,In_2648,In_1640);
and U1373 (N_1373,In_740,In_2263);
xnor U1374 (N_1374,In_2037,In_254);
and U1375 (N_1375,In_2427,In_774);
nand U1376 (N_1376,In_551,In_2300);
nand U1377 (N_1377,In_2722,In_66);
nand U1378 (N_1378,In_912,In_1082);
nor U1379 (N_1379,In_2601,In_623);
xor U1380 (N_1380,In_2942,In_2866);
nand U1381 (N_1381,In_361,In_2734);
or U1382 (N_1382,In_1951,In_570);
or U1383 (N_1383,In_2379,In_1934);
and U1384 (N_1384,In_236,In_2887);
nand U1385 (N_1385,In_391,In_2365);
nor U1386 (N_1386,In_1609,In_628);
nand U1387 (N_1387,In_1049,In_228);
nand U1388 (N_1388,In_2518,In_1264);
nor U1389 (N_1389,In_200,In_1565);
xnor U1390 (N_1390,In_1014,In_2691);
or U1391 (N_1391,In_1569,In_667);
or U1392 (N_1392,In_1114,In_2175);
or U1393 (N_1393,In_2945,In_114);
and U1394 (N_1394,In_1744,In_1545);
or U1395 (N_1395,In_2538,In_2936);
nor U1396 (N_1396,In_2582,In_2429);
and U1397 (N_1397,In_1605,In_1026);
and U1398 (N_1398,In_93,In_2106);
nand U1399 (N_1399,In_1113,In_2767);
or U1400 (N_1400,In_2859,In_108);
and U1401 (N_1401,In_2282,In_1287);
or U1402 (N_1402,In_1589,In_2034);
nand U1403 (N_1403,In_1852,In_976);
and U1404 (N_1404,In_1158,In_709);
nand U1405 (N_1405,In_1540,In_1535);
xnor U1406 (N_1406,In_414,In_1289);
and U1407 (N_1407,In_1978,In_917);
xnor U1408 (N_1408,In_2514,In_583);
xnor U1409 (N_1409,In_2064,In_2544);
nand U1410 (N_1410,In_2111,In_2185);
and U1411 (N_1411,In_2525,In_797);
xor U1412 (N_1412,In_1374,In_1319);
or U1413 (N_1413,In_6,In_2776);
xnor U1414 (N_1414,In_2489,In_1138);
xnor U1415 (N_1415,In_1555,In_553);
nor U1416 (N_1416,In_95,In_2869);
or U1417 (N_1417,In_1336,In_2739);
nand U1418 (N_1418,In_2347,In_1347);
and U1419 (N_1419,In_1979,In_2085);
nand U1420 (N_1420,In_1330,In_1765);
xnor U1421 (N_1421,In_1212,In_1630);
and U1422 (N_1422,In_259,In_1774);
xnor U1423 (N_1423,In_1779,In_2018);
xnor U1424 (N_1424,In_363,In_1234);
or U1425 (N_1425,In_1035,In_187);
nor U1426 (N_1426,In_2040,In_1703);
or U1427 (N_1427,In_1344,In_417);
and U1428 (N_1428,In_2728,In_1888);
xor U1429 (N_1429,In_2067,In_582);
nand U1430 (N_1430,In_2930,In_571);
or U1431 (N_1431,In_1624,In_1245);
xor U1432 (N_1432,In_2138,In_665);
or U1433 (N_1433,In_2478,In_2466);
nand U1434 (N_1434,In_869,In_974);
or U1435 (N_1435,In_2492,In_2987);
nor U1436 (N_1436,In_2487,In_2830);
nand U1437 (N_1437,In_1229,In_2920);
nand U1438 (N_1438,In_2402,In_1325);
or U1439 (N_1439,In_2161,In_348);
xor U1440 (N_1440,In_1823,In_1304);
and U1441 (N_1441,In_2980,In_562);
nand U1442 (N_1442,In_1286,In_1411);
or U1443 (N_1443,In_621,In_2985);
xor U1444 (N_1444,In_2003,In_1223);
and U1445 (N_1445,In_2378,In_165);
nor U1446 (N_1446,In_1782,In_101);
or U1447 (N_1447,In_2531,In_1392);
or U1448 (N_1448,In_1255,In_1633);
and U1449 (N_1449,In_1283,In_1647);
and U1450 (N_1450,In_51,In_2753);
xnor U1451 (N_1451,In_1928,In_733);
xor U1452 (N_1452,In_1777,In_2247);
and U1453 (N_1453,In_2848,In_993);
or U1454 (N_1454,In_580,In_136);
nand U1455 (N_1455,In_2202,In_1207);
xnor U1456 (N_1456,In_2741,In_723);
nand U1457 (N_1457,In_999,In_2671);
nor U1458 (N_1458,In_713,In_1830);
nand U1459 (N_1459,In_250,In_1843);
and U1460 (N_1460,In_2128,In_1032);
and U1461 (N_1461,In_131,In_616);
xor U1462 (N_1462,In_2906,In_714);
nand U1463 (N_1463,In_590,In_2278);
nor U1464 (N_1464,In_2326,In_1233);
or U1465 (N_1465,In_1384,In_2964);
xor U1466 (N_1466,In_1045,In_1493);
nand U1467 (N_1467,In_1776,In_2007);
and U1468 (N_1468,In_1291,In_2515);
and U1469 (N_1469,In_1964,In_161);
and U1470 (N_1470,In_1091,In_1672);
nand U1471 (N_1471,In_2800,In_1054);
xnor U1472 (N_1472,In_2142,In_1584);
xnor U1473 (N_1473,In_2189,In_2814);
nor U1474 (N_1474,In_1359,In_2513);
nand U1475 (N_1475,In_2684,In_1570);
or U1476 (N_1476,In_597,In_1983);
or U1477 (N_1477,In_2817,In_1475);
nor U1478 (N_1478,In_1850,In_1720);
nor U1479 (N_1479,In_691,In_2422);
or U1480 (N_1480,In_308,In_2206);
and U1481 (N_1481,In_182,In_2816);
nand U1482 (N_1482,In_2529,In_407);
xor U1483 (N_1483,In_1474,In_2109);
nand U1484 (N_1484,In_2560,In_1147);
xor U1485 (N_1485,In_1294,In_750);
nand U1486 (N_1486,In_322,In_1409);
or U1487 (N_1487,In_857,In_2121);
nand U1488 (N_1488,In_1598,In_889);
nand U1489 (N_1489,In_1440,In_1740);
and U1490 (N_1490,In_2864,In_896);
and U1491 (N_1491,In_2236,In_2683);
and U1492 (N_1492,In_2497,In_1757);
nor U1493 (N_1493,In_263,In_2979);
xor U1494 (N_1494,In_662,In_1108);
xor U1495 (N_1495,In_413,In_2564);
xnor U1496 (N_1496,In_2494,In_514);
nand U1497 (N_1497,In_858,In_1636);
nor U1498 (N_1498,In_1486,In_1897);
and U1499 (N_1499,In_1307,In_1137);
or U1500 (N_1500,N_274,N_1218);
nor U1501 (N_1501,N_1473,N_388);
or U1502 (N_1502,N_883,N_224);
xnor U1503 (N_1503,N_61,N_252);
or U1504 (N_1504,N_1337,N_10);
and U1505 (N_1505,N_1274,N_1076);
and U1506 (N_1506,N_912,N_936);
nand U1507 (N_1507,N_1153,N_266);
nand U1508 (N_1508,N_147,N_921);
nor U1509 (N_1509,N_194,N_401);
nor U1510 (N_1510,N_1312,N_1290);
or U1511 (N_1511,N_228,N_17);
xnor U1512 (N_1512,N_521,N_1224);
nand U1513 (N_1513,N_569,N_57);
nand U1514 (N_1514,N_1383,N_781);
and U1515 (N_1515,N_1061,N_817);
and U1516 (N_1516,N_518,N_530);
xor U1517 (N_1517,N_144,N_1059);
or U1518 (N_1518,N_986,N_1227);
or U1519 (N_1519,N_201,N_141);
and U1520 (N_1520,N_1198,N_565);
nand U1521 (N_1521,N_773,N_353);
nor U1522 (N_1522,N_453,N_1089);
nand U1523 (N_1523,N_1318,N_68);
or U1524 (N_1524,N_1474,N_1382);
or U1525 (N_1525,N_435,N_1499);
or U1526 (N_1526,N_696,N_6);
nor U1527 (N_1527,N_1207,N_1292);
or U1528 (N_1528,N_957,N_1284);
xnor U1529 (N_1529,N_498,N_944);
nor U1530 (N_1530,N_778,N_750);
xnor U1531 (N_1531,N_1273,N_272);
or U1532 (N_1532,N_64,N_1239);
nor U1533 (N_1533,N_841,N_164);
xnor U1534 (N_1534,N_1323,N_1495);
xor U1535 (N_1535,N_1168,N_737);
and U1536 (N_1536,N_1389,N_1062);
nand U1537 (N_1537,N_803,N_1392);
and U1538 (N_1538,N_859,N_605);
or U1539 (N_1539,N_223,N_1080);
nor U1540 (N_1540,N_710,N_1232);
xor U1541 (N_1541,N_262,N_475);
and U1542 (N_1542,N_765,N_374);
or U1543 (N_1543,N_1331,N_1391);
nor U1544 (N_1544,N_1357,N_465);
and U1545 (N_1545,N_395,N_29);
nand U1546 (N_1546,N_776,N_175);
and U1547 (N_1547,N_1065,N_60);
or U1548 (N_1548,N_914,N_84);
and U1549 (N_1549,N_1333,N_1395);
xor U1550 (N_1550,N_768,N_990);
xnor U1551 (N_1551,N_1370,N_1070);
nor U1552 (N_1552,N_83,N_1088);
nand U1553 (N_1553,N_20,N_685);
xor U1554 (N_1554,N_153,N_1260);
and U1555 (N_1555,N_1275,N_51);
nor U1556 (N_1556,N_1004,N_1172);
nor U1557 (N_1557,N_563,N_1121);
or U1558 (N_1558,N_1226,N_1481);
or U1559 (N_1559,N_327,N_71);
and U1560 (N_1560,N_92,N_805);
nor U1561 (N_1561,N_377,N_42);
and U1562 (N_1562,N_1064,N_995);
or U1563 (N_1563,N_671,N_203);
nand U1564 (N_1564,N_1210,N_1092);
nor U1565 (N_1565,N_472,N_634);
nor U1566 (N_1566,N_451,N_344);
xor U1567 (N_1567,N_1072,N_221);
xnor U1568 (N_1568,N_1068,N_1487);
or U1569 (N_1569,N_31,N_938);
nor U1570 (N_1570,N_1354,N_705);
xnor U1571 (N_1571,N_976,N_1456);
nand U1572 (N_1572,N_67,N_370);
or U1573 (N_1573,N_1302,N_298);
nor U1574 (N_1574,N_180,N_522);
nor U1575 (N_1575,N_1316,N_503);
nor U1576 (N_1576,N_1240,N_507);
nor U1577 (N_1577,N_933,N_1016);
or U1578 (N_1578,N_647,N_242);
nand U1579 (N_1579,N_430,N_948);
nor U1580 (N_1580,N_1155,N_1025);
nand U1581 (N_1581,N_861,N_1222);
nor U1582 (N_1582,N_244,N_992);
xnor U1583 (N_1583,N_1005,N_693);
nor U1584 (N_1584,N_512,N_222);
xnor U1585 (N_1585,N_18,N_1291);
and U1586 (N_1586,N_850,N_1398);
nand U1587 (N_1587,N_1196,N_586);
and U1588 (N_1588,N_429,N_1431);
nand U1589 (N_1589,N_954,N_645);
nand U1590 (N_1590,N_162,N_1235);
and U1591 (N_1591,N_1242,N_580);
nor U1592 (N_1592,N_1037,N_744);
xnor U1593 (N_1593,N_903,N_959);
xor U1594 (N_1594,N_732,N_1493);
nand U1595 (N_1595,N_230,N_269);
and U1596 (N_1596,N_13,N_932);
xnor U1597 (N_1597,N_1165,N_366);
or U1598 (N_1598,N_1148,N_1256);
nand U1599 (N_1599,N_177,N_205);
xor U1600 (N_1600,N_546,N_913);
nor U1601 (N_1601,N_39,N_253);
nor U1602 (N_1602,N_606,N_1458);
xnor U1603 (N_1603,N_785,N_978);
nand U1604 (N_1604,N_434,N_484);
or U1605 (N_1605,N_1255,N_440);
xnor U1606 (N_1606,N_1454,N_432);
nand U1607 (N_1607,N_1018,N_1369);
or U1608 (N_1608,N_247,N_927);
and U1609 (N_1609,N_243,N_720);
nor U1610 (N_1610,N_980,N_418);
xor U1611 (N_1611,N_759,N_1156);
xor U1612 (N_1612,N_22,N_456);
or U1613 (N_1613,N_1073,N_90);
nor U1614 (N_1614,N_209,N_404);
nor U1615 (N_1615,N_641,N_760);
xnor U1616 (N_1616,N_753,N_103);
nand U1617 (N_1617,N_1390,N_246);
or U1618 (N_1618,N_931,N_206);
xor U1619 (N_1619,N_1099,N_746);
or U1620 (N_1620,N_1342,N_1447);
xnor U1621 (N_1621,N_1332,N_183);
nand U1622 (N_1622,N_469,N_1243);
xor U1623 (N_1623,N_731,N_1125);
xnor U1624 (N_1624,N_493,N_545);
or U1625 (N_1625,N_33,N_1405);
xnor U1626 (N_1626,N_322,N_89);
nand U1627 (N_1627,N_952,N_66);
or U1628 (N_1628,N_1325,N_820);
nor U1629 (N_1629,N_899,N_400);
nand U1630 (N_1630,N_702,N_268);
xnor U1631 (N_1631,N_277,N_195);
or U1632 (N_1632,N_558,N_91);
nor U1633 (N_1633,N_1010,N_158);
and U1634 (N_1634,N_1414,N_681);
or U1635 (N_1635,N_80,N_1434);
or U1636 (N_1636,N_176,N_801);
xor U1637 (N_1637,N_112,N_1330);
and U1638 (N_1638,N_544,N_1338);
xor U1639 (N_1639,N_939,N_1321);
nand U1640 (N_1640,N_853,N_624);
nor U1641 (N_1641,N_791,N_682);
nor U1642 (N_1642,N_282,N_998);
xor U1643 (N_1643,N_1409,N_72);
nor U1644 (N_1644,N_1228,N_1281);
nor U1645 (N_1645,N_1415,N_220);
nor U1646 (N_1646,N_630,N_387);
nor U1647 (N_1647,N_725,N_1287);
xnor U1648 (N_1648,N_114,N_55);
or U1649 (N_1649,N_74,N_1253);
xnor U1650 (N_1650,N_1490,N_982);
xnor U1651 (N_1651,N_1028,N_782);
or U1652 (N_1652,N_863,N_45);
or U1653 (N_1653,N_734,N_751);
or U1654 (N_1654,N_113,N_1223);
and U1655 (N_1655,N_467,N_1124);
nand U1656 (N_1656,N_1297,N_28);
nand U1657 (N_1657,N_1241,N_384);
nand U1658 (N_1658,N_1047,N_1497);
and U1659 (N_1659,N_1254,N_822);
xor U1660 (N_1660,N_208,N_1277);
and U1661 (N_1661,N_455,N_738);
and U1662 (N_1662,N_1400,N_1257);
or U1663 (N_1663,N_1324,N_550);
xor U1664 (N_1664,N_52,N_819);
and U1665 (N_1665,N_542,N_286);
or U1666 (N_1666,N_811,N_894);
nand U1667 (N_1667,N_1095,N_187);
nor U1668 (N_1668,N_470,N_721);
nand U1669 (N_1669,N_733,N_1205);
and U1670 (N_1670,N_1211,N_1445);
xnor U1671 (N_1671,N_191,N_623);
xor U1672 (N_1672,N_1074,N_1430);
nor U1673 (N_1673,N_412,N_800);
nor U1674 (N_1674,N_504,N_1426);
nand U1675 (N_1675,N_829,N_895);
nor U1676 (N_1676,N_735,N_163);
nor U1677 (N_1677,N_362,N_5);
and U1678 (N_1678,N_905,N_1105);
and U1679 (N_1679,N_761,N_136);
nor U1680 (N_1680,N_873,N_173);
and U1681 (N_1681,N_1336,N_238);
xnor U1682 (N_1682,N_302,N_1424);
and U1683 (N_1683,N_834,N_123);
nand U1684 (N_1684,N_310,N_1294);
nor U1685 (N_1685,N_178,N_1109);
nand U1686 (N_1686,N_1160,N_24);
nand U1687 (N_1687,N_446,N_452);
and U1688 (N_1688,N_359,N_334);
nor U1689 (N_1689,N_288,N_474);
nand U1690 (N_1690,N_716,N_701);
and U1691 (N_1691,N_528,N_379);
nand U1692 (N_1692,N_1317,N_41);
and U1693 (N_1693,N_248,N_576);
or U1694 (N_1694,N_239,N_76);
or U1695 (N_1695,N_240,N_1233);
nor U1696 (N_1696,N_887,N_494);
nand U1697 (N_1697,N_572,N_1491);
or U1698 (N_1698,N_145,N_1163);
and U1699 (N_1699,N_532,N_1451);
nand U1700 (N_1700,N_762,N_922);
nor U1701 (N_1701,N_1219,N_1345);
or U1702 (N_1702,N_795,N_852);
nand U1703 (N_1703,N_742,N_602);
xnor U1704 (N_1704,N_78,N_1249);
or U1705 (N_1705,N_381,N_506);
and U1706 (N_1706,N_666,N_851);
nand U1707 (N_1707,N_642,N_981);
xor U1708 (N_1708,N_1286,N_308);
xor U1709 (N_1709,N_1149,N_613);
xnor U1710 (N_1710,N_1278,N_133);
xnor U1711 (N_1711,N_622,N_984);
and U1712 (N_1712,N_254,N_447);
and U1713 (N_1713,N_1268,N_1334);
or U1714 (N_1714,N_295,N_390);
and U1715 (N_1715,N_961,N_1230);
nor U1716 (N_1716,N_367,N_1011);
and U1717 (N_1717,N_798,N_407);
or U1718 (N_1718,N_1050,N_146);
and U1719 (N_1719,N_871,N_174);
or U1720 (N_1720,N_1134,N_307);
or U1721 (N_1721,N_448,N_1195);
and U1722 (N_1722,N_140,N_758);
or U1723 (N_1723,N_797,N_293);
nor U1724 (N_1724,N_1102,N_391);
nand U1725 (N_1725,N_166,N_462);
nor U1726 (N_1726,N_98,N_49);
nor U1727 (N_1727,N_481,N_637);
or U1728 (N_1728,N_1387,N_424);
and U1729 (N_1729,N_996,N_1193);
xnor U1730 (N_1730,N_499,N_101);
nor U1731 (N_1731,N_336,N_265);
nor U1732 (N_1732,N_321,N_331);
xnor U1733 (N_1733,N_1478,N_290);
and U1734 (N_1734,N_697,N_58);
or U1735 (N_1735,N_593,N_1267);
nor U1736 (N_1736,N_468,N_309);
xnor U1737 (N_1737,N_1271,N_38);
nor U1738 (N_1738,N_1049,N_584);
and U1739 (N_1739,N_655,N_1192);
xnor U1740 (N_1740,N_923,N_1107);
and U1741 (N_1741,N_699,N_1280);
or U1742 (N_1742,N_263,N_1335);
nand U1743 (N_1743,N_1351,N_81);
nor U1744 (N_1744,N_397,N_1096);
xor U1745 (N_1745,N_790,N_943);
nand U1746 (N_1746,N_385,N_405);
xnor U1747 (N_1747,N_445,N_1410);
xnor U1748 (N_1748,N_1470,N_715);
and U1749 (N_1749,N_333,N_100);
nand U1750 (N_1750,N_116,N_457);
xor U1751 (N_1751,N_568,N_1123);
or U1752 (N_1752,N_599,N_1375);
xor U1753 (N_1753,N_488,N_712);
or U1754 (N_1754,N_1413,N_1475);
nand U1755 (N_1755,N_1270,N_1307);
nor U1756 (N_1756,N_1457,N_1311);
or U1757 (N_1757,N_1194,N_1182);
nor U1758 (N_1758,N_1175,N_1419);
or U1759 (N_1759,N_1306,N_600);
nand U1760 (N_1760,N_380,N_1485);
and U1761 (N_1761,N_1174,N_821);
nor U1762 (N_1762,N_9,N_972);
and U1763 (N_1763,N_818,N_1460);
nor U1764 (N_1764,N_1461,N_722);
and U1765 (N_1765,N_305,N_1180);
xnor U1766 (N_1766,N_150,N_571);
xor U1767 (N_1767,N_919,N_1244);
or U1768 (N_1768,N_755,N_537);
nor U1769 (N_1769,N_471,N_125);
xnor U1770 (N_1770,N_890,N_27);
nor U1771 (N_1771,N_1203,N_214);
nand U1772 (N_1772,N_1063,N_1373);
and U1773 (N_1773,N_1299,N_486);
and U1774 (N_1774,N_1450,N_1386);
and U1775 (N_1775,N_756,N_551);
nand U1776 (N_1776,N_1183,N_1197);
nand U1777 (N_1777,N_1420,N_1465);
or U1778 (N_1778,N_313,N_1399);
xor U1779 (N_1779,N_118,N_708);
nand U1780 (N_1780,N_53,N_907);
and U1781 (N_1781,N_1007,N_372);
or U1782 (N_1782,N_662,N_423);
or U1783 (N_1783,N_261,N_612);
or U1784 (N_1784,N_777,N_999);
nand U1785 (N_1785,N_170,N_607);
or U1786 (N_1786,N_433,N_591);
or U1787 (N_1787,N_65,N_349);
nor U1788 (N_1788,N_1229,N_1135);
nand U1789 (N_1789,N_496,N_842);
xnor U1790 (N_1790,N_570,N_951);
nand U1791 (N_1791,N_99,N_1116);
xnor U1792 (N_1792,N_219,N_937);
xnor U1793 (N_1793,N_611,N_562);
nand U1794 (N_1794,N_1213,N_1093);
nand U1795 (N_1795,N_659,N_1077);
nand U1796 (N_1796,N_875,N_646);
xnor U1797 (N_1797,N_1376,N_1380);
nand U1798 (N_1798,N_406,N_399);
nand U1799 (N_1799,N_698,N_1177);
nand U1800 (N_1800,N_1326,N_316);
nand U1801 (N_1801,N_1328,N_318);
nand U1802 (N_1802,N_2,N_1048);
or U1803 (N_1803,N_1439,N_1101);
nand U1804 (N_1804,N_1300,N_1122);
nor U1805 (N_1805,N_902,N_182);
nand U1806 (N_1806,N_582,N_1162);
or U1807 (N_1807,N_257,N_552);
nand U1808 (N_1808,N_121,N_635);
nand U1809 (N_1809,N_1443,N_213);
nand U1810 (N_1810,N_706,N_458);
nor U1811 (N_1811,N_414,N_1412);
and U1812 (N_1812,N_1237,N_631);
nor U1813 (N_1813,N_814,N_1388);
xnor U1814 (N_1814,N_864,N_1408);
xnor U1815 (N_1815,N_19,N_517);
xnor U1816 (N_1816,N_1138,N_704);
xor U1817 (N_1817,N_726,N_1411);
xor U1818 (N_1818,N_207,N_1120);
or U1819 (N_1819,N_199,N_216);
xor U1820 (N_1820,N_1054,N_1440);
or U1821 (N_1821,N_1362,N_840);
or U1822 (N_1822,N_843,N_700);
nand U1823 (N_1823,N_189,N_371);
nand U1824 (N_1824,N_250,N_1452);
nor U1825 (N_1825,N_849,N_1459);
or U1826 (N_1826,N_1236,N_598);
and U1827 (N_1827,N_879,N_1248);
and U1828 (N_1828,N_962,N_925);
xor U1829 (N_1829,N_1110,N_1463);
nand U1830 (N_1830,N_270,N_294);
xor U1831 (N_1831,N_1377,N_126);
nand U1832 (N_1832,N_1154,N_809);
or U1833 (N_1833,N_1191,N_1264);
or U1834 (N_1834,N_1090,N_906);
nand U1835 (N_1835,N_1350,N_916);
nor U1836 (N_1836,N_533,N_413);
nor U1837 (N_1837,N_736,N_977);
xnor U1838 (N_1838,N_691,N_1282);
or U1839 (N_1839,N_312,N_1303);
nor U1840 (N_1840,N_59,N_82);
nor U1841 (N_1841,N_36,N_709);
nor U1842 (N_1842,N_44,N_225);
nor U1843 (N_1843,N_1084,N_264);
xor U1844 (N_1844,N_363,N_421);
or U1845 (N_1845,N_870,N_1117);
nand U1846 (N_1846,N_604,N_131);
nor U1847 (N_1847,N_1114,N_994);
nor U1848 (N_1848,N_1462,N_810);
or U1849 (N_1849,N_1051,N_1140);
or U1850 (N_1850,N_956,N_1032);
nor U1851 (N_1851,N_534,N_857);
xnor U1852 (N_1852,N_945,N_1115);
xor U1853 (N_1853,N_329,N_1385);
nand U1854 (N_1854,N_652,N_1313);
xnor U1855 (N_1855,N_1471,N_459);
nor U1856 (N_1856,N_1247,N_618);
xor U1857 (N_1857,N_478,N_1441);
or U1858 (N_1858,N_1003,N_193);
or U1859 (N_1859,N_1378,N_54);
or U1860 (N_1860,N_301,N_56);
xor U1861 (N_1861,N_1170,N_644);
xor U1862 (N_1862,N_855,N_1397);
or U1863 (N_1863,N_616,N_483);
xnor U1864 (N_1864,N_276,N_947);
nand U1865 (N_1865,N_1315,N_675);
nor U1866 (N_1866,N_718,N_320);
xor U1867 (N_1867,N_93,N_1098);
or U1868 (N_1868,N_909,N_231);
or U1869 (N_1869,N_970,N_752);
or U1870 (N_1870,N_383,N_376);
nand U1871 (N_1871,N_1266,N_284);
or U1872 (N_1872,N_1329,N_1322);
nand U1873 (N_1873,N_1201,N_884);
or U1874 (N_1874,N_513,N_711);
or U1875 (N_1875,N_454,N_1019);
nand U1876 (N_1876,N_1427,N_1144);
and U1877 (N_1877,N_3,N_1480);
and U1878 (N_1878,N_1027,N_489);
and U1879 (N_1879,N_1141,N_975);
and U1880 (N_1880,N_94,N_77);
xnor U1881 (N_1881,N_32,N_826);
and U1882 (N_1882,N_345,N_573);
xor U1883 (N_1883,N_540,N_500);
xnor U1884 (N_1884,N_633,N_908);
or U1885 (N_1885,N_1171,N_1035);
nor U1886 (N_1886,N_1015,N_719);
xor U1887 (N_1887,N_1252,N_129);
nor U1888 (N_1888,N_161,N_1301);
or U1889 (N_1889,N_941,N_1094);
and U1890 (N_1890,N_583,N_523);
and U1891 (N_1891,N_210,N_514);
xnor U1892 (N_1892,N_930,N_138);
nand U1893 (N_1893,N_1130,N_767);
or U1894 (N_1894,N_63,N_694);
xor U1895 (N_1895,N_119,N_987);
and U1896 (N_1896,N_1444,N_185);
nor U1897 (N_1897,N_846,N_1021);
or U1898 (N_1898,N_564,N_1432);
and U1899 (N_1899,N_997,N_665);
and U1900 (N_1900,N_1147,N_862);
and U1901 (N_1901,N_117,N_1288);
or U1902 (N_1902,N_409,N_949);
and U1903 (N_1903,N_460,N_314);
or U1904 (N_1904,N_1104,N_1407);
xnor U1905 (N_1905,N_743,N_135);
xnor U1906 (N_1906,N_168,N_784);
xnor U1907 (N_1907,N_1179,N_215);
and U1908 (N_1908,N_292,N_26);
or U1909 (N_1909,N_0,N_46);
and U1910 (N_1910,N_788,N_640);
or U1911 (N_1911,N_520,N_1013);
and U1912 (N_1912,N_649,N_1368);
xor U1913 (N_1913,N_1359,N_1467);
xor U1914 (N_1914,N_47,N_11);
nand U1915 (N_1915,N_929,N_1214);
nand U1916 (N_1916,N_554,N_1103);
nor U1917 (N_1917,N_1043,N_969);
xnor U1918 (N_1918,N_234,N_964);
nor U1919 (N_1919,N_1418,N_110);
nor U1920 (N_1920,N_1143,N_1085);
xor U1921 (N_1921,N_154,N_1045);
xnor U1922 (N_1922,N_1261,N_73);
xor U1923 (N_1923,N_415,N_1173);
nand U1924 (N_1924,N_356,N_137);
xnor U1925 (N_1925,N_502,N_592);
nor U1926 (N_1926,N_657,N_688);
nor U1927 (N_1927,N_97,N_1285);
xnor U1928 (N_1928,N_1366,N_619);
nor U1929 (N_1929,N_1258,N_1464);
nor U1930 (N_1930,N_979,N_335);
nor U1931 (N_1931,N_425,N_212);
and U1932 (N_1932,N_654,N_771);
and U1933 (N_1933,N_297,N_886);
or U1934 (N_1934,N_326,N_62);
nand U1935 (N_1935,N_155,N_1437);
nor U1936 (N_1936,N_1029,N_687);
xor U1937 (N_1937,N_837,N_881);
nor U1938 (N_1938,N_1379,N_727);
nand U1939 (N_1939,N_1053,N_1449);
xor U1940 (N_1940,N_373,N_872);
xor U1941 (N_1941,N_196,N_747);
nand U1942 (N_1942,N_1453,N_828);
xor U1943 (N_1943,N_830,N_431);
and U1944 (N_1944,N_878,N_1157);
nand U1945 (N_1945,N_1097,N_856);
nand U1946 (N_1946,N_1221,N_1341);
xor U1947 (N_1947,N_70,N_1309);
and U1948 (N_1948,N_251,N_748);
and U1949 (N_1949,N_271,N_1052);
and U1950 (N_1950,N_749,N_1404);
xor U1951 (N_1951,N_661,N_966);
or U1952 (N_1952,N_278,N_1279);
nor U1953 (N_1953,N_764,N_197);
nor U1954 (N_1954,N_422,N_1484);
nand U1955 (N_1955,N_891,N_1381);
xnor U1956 (N_1956,N_926,N_226);
nand U1957 (N_1957,N_985,N_1202);
or U1958 (N_1958,N_1308,N_303);
and U1959 (N_1959,N_104,N_1071);
xnor U1960 (N_1960,N_621,N_296);
or U1961 (N_1961,N_786,N_1394);
nor U1962 (N_1962,N_30,N_283);
or U1963 (N_1963,N_1320,N_495);
nor U1964 (N_1964,N_23,N_588);
or U1965 (N_1965,N_1353,N_1293);
xor U1966 (N_1966,N_1340,N_325);
nand U1967 (N_1967,N_1041,N_339);
or U1968 (N_1968,N_369,N_233);
nor U1969 (N_1969,N_351,N_650);
or U1970 (N_1970,N_273,N_1129);
xnor U1971 (N_1971,N_355,N_1161);
xor U1972 (N_1972,N_449,N_1187);
xor U1973 (N_1973,N_287,N_779);
and U1974 (N_1974,N_1262,N_901);
nor U1975 (N_1975,N_143,N_1479);
and U1976 (N_1976,N_127,N_382);
nand U1977 (N_1977,N_868,N_892);
xor U1978 (N_1978,N_306,N_854);
xor U1979 (N_1979,N_280,N_561);
nand U1980 (N_1980,N_1108,N_4);
and U1981 (N_1981,N_553,N_1446);
and U1982 (N_1982,N_392,N_793);
or U1983 (N_1983,N_581,N_1000);
xor U1984 (N_1984,N_490,N_967);
xor U1985 (N_1985,N_15,N_299);
xor U1986 (N_1986,N_416,N_664);
or U1987 (N_1987,N_442,N_439);
nor U1988 (N_1988,N_482,N_1246);
nor U1989 (N_1989,N_1492,N_874);
and U1990 (N_1990,N_1006,N_1184);
and U1991 (N_1991,N_690,N_1423);
and U1992 (N_1992,N_1136,N_1269);
xnor U1993 (N_1993,N_1199,N_347);
nor U1994 (N_1994,N_858,N_466);
nor U1995 (N_1995,N_615,N_663);
nand U1996 (N_1996,N_1188,N_1489);
or U1997 (N_1997,N_1039,N_450);
or U1998 (N_1998,N_527,N_343);
nand U1999 (N_1999,N_1436,N_953);
nand U2000 (N_2000,N_539,N_845);
nor U2001 (N_2001,N_1164,N_668);
nor U2002 (N_2002,N_1057,N_1477);
xor U2003 (N_2003,N_638,N_940);
or U2004 (N_2004,N_876,N_867);
or U2005 (N_2005,N_281,N_237);
nand U2006 (N_2006,N_667,N_1361);
nand U2007 (N_2007,N_95,N_1403);
and U2008 (N_2008,N_594,N_7);
nand U2009 (N_2009,N_1416,N_1044);
or U2010 (N_2010,N_1396,N_368);
nor U2011 (N_2011,N_684,N_658);
nand U2012 (N_2012,N_656,N_245);
and U2013 (N_2013,N_780,N_556);
nor U2014 (N_2014,N_1272,N_1126);
or U2015 (N_2015,N_1139,N_896);
xor U2016 (N_2016,N_43,N_1349);
nor U2017 (N_2017,N_1014,N_596);
nand U2018 (N_2018,N_1060,N_394);
or U2019 (N_2019,N_974,N_1158);
and U2020 (N_2020,N_160,N_918);
nor U2021 (N_2021,N_838,N_1421);
and U2022 (N_2022,N_1002,N_674);
and U2023 (N_2023,N_1393,N_364);
nor U2024 (N_2024,N_559,N_186);
nand U2025 (N_2025,N_968,N_832);
or U2026 (N_2026,N_410,N_608);
or U2027 (N_2027,N_1146,N_683);
nor U2028 (N_2028,N_134,N_21);
or U2029 (N_2029,N_880,N_48);
nand U2030 (N_2030,N_1360,N_703);
and U2031 (N_2031,N_1009,N_1026);
nor U2032 (N_2032,N_1151,N_403);
and U2033 (N_2033,N_833,N_441);
and U2034 (N_2034,N_1069,N_1091);
nand U2035 (N_2035,N_1127,N_428);
xnor U2036 (N_2036,N_772,N_361);
nand U2037 (N_2037,N_802,N_35);
and U2038 (N_2038,N_156,N_549);
or U2039 (N_2039,N_1231,N_1251);
xor U2040 (N_2040,N_1428,N_511);
xor U2041 (N_2041,N_632,N_792);
nand U2042 (N_2042,N_950,N_190);
xnor U2043 (N_2043,N_695,N_882);
nor U2044 (N_2044,N_740,N_426);
nand U2045 (N_2045,N_1367,N_536);
or U2046 (N_2046,N_1131,N_476);
and U2047 (N_2047,N_516,N_1468);
nor U2048 (N_2048,N_443,N_1058);
xnor U2049 (N_2049,N_825,N_888);
or U2050 (N_2050,N_1448,N_236);
or U2051 (N_2051,N_477,N_673);
nand U2052 (N_2052,N_739,N_86);
nor U2053 (N_2053,N_165,N_807);
and U2054 (N_2054,N_519,N_1100);
or U2055 (N_2055,N_437,N_386);
nand U2056 (N_2056,N_590,N_106);
and U2057 (N_2057,N_169,N_567);
xnor U2058 (N_2058,N_12,N_839);
xor U2059 (N_2059,N_877,N_525);
nand U2060 (N_2060,N_915,N_893);
xor U2061 (N_2061,N_1020,N_1142);
xor U2062 (N_2062,N_1185,N_105);
xnor U2063 (N_2063,N_256,N_87);
or U2064 (N_2064,N_651,N_111);
xnor U2065 (N_2065,N_291,N_375);
nor U2066 (N_2066,N_1344,N_865);
nand U2067 (N_2067,N_1150,N_538);
xnor U2068 (N_2068,N_1305,N_955);
and U2069 (N_2069,N_920,N_1225);
or U2070 (N_2070,N_198,N_14);
and U2071 (N_2071,N_204,N_1310);
or U2072 (N_2072,N_796,N_323);
nand U2073 (N_2073,N_217,N_1494);
nor U2074 (N_2074,N_1078,N_1206);
xor U2075 (N_2075,N_461,N_357);
nand U2076 (N_2076,N_491,N_689);
and U2077 (N_2077,N_319,N_754);
xor U2078 (N_2078,N_1466,N_900);
nand U2079 (N_2079,N_1067,N_766);
nor U2080 (N_2080,N_1087,N_714);
nand U2081 (N_2081,N_402,N_885);
and U2082 (N_2082,N_1295,N_1215);
nand U2083 (N_2083,N_626,N_1371);
or U2084 (N_2084,N_96,N_1476);
and U2085 (N_2085,N_1438,N_844);
nor U2086 (N_2086,N_1455,N_1022);
or U2087 (N_2087,N_775,N_770);
nand U2088 (N_2088,N_255,N_1355);
nor U2089 (N_2089,N_188,N_192);
and U2090 (N_2090,N_279,N_848);
and U2091 (N_2091,N_783,N_643);
and U2092 (N_2092,N_151,N_1435);
or U2093 (N_2093,N_202,N_1469);
xor U2094 (N_2094,N_328,N_88);
nand U2095 (N_2095,N_505,N_1046);
and U2096 (N_2096,N_960,N_420);
nand U2097 (N_2097,N_317,N_1166);
or U2098 (N_2098,N_1358,N_389);
nor U2099 (N_2099,N_1245,N_229);
and U2100 (N_2100,N_835,N_1339);
nand U2101 (N_2101,N_1082,N_358);
xnor U2102 (N_2102,N_620,N_988);
nor U2103 (N_2103,N_152,N_348);
xor U2104 (N_2104,N_1001,N_1075);
nor U2105 (N_2105,N_898,N_610);
and U2106 (N_2106,N_108,N_289);
and U2107 (N_2107,N_1298,N_804);
nand U2108 (N_2108,N_232,N_1128);
nor U2109 (N_2109,N_75,N_149);
xor U2110 (N_2110,N_1356,N_813);
or U2111 (N_2111,N_1112,N_679);
nor U2112 (N_2112,N_601,N_157);
and U2113 (N_2113,N_989,N_578);
nor U2114 (N_2114,N_1289,N_774);
and U2115 (N_2115,N_1276,N_1250);
nand U2116 (N_2116,N_787,N_910);
nand U2117 (N_2117,N_1036,N_436);
or U2118 (N_2118,N_464,N_1442);
xnor U2119 (N_2119,N_120,N_692);
nand U2120 (N_2120,N_479,N_971);
or U2121 (N_2121,N_267,N_524);
nor U2122 (N_2122,N_597,N_16);
and U2123 (N_2123,N_677,N_812);
or U2124 (N_2124,N_1152,N_942);
or U2125 (N_2125,N_1023,N_1133);
nor U2126 (N_2126,N_917,N_560);
or U2127 (N_2127,N_1429,N_769);
or U2128 (N_2128,N_142,N_991);
nand U2129 (N_2129,N_1034,N_1238);
xor U2130 (N_2130,N_124,N_1384);
nand U2131 (N_2131,N_1352,N_159);
nand U2132 (N_2132,N_816,N_1024);
xor U2133 (N_2133,N_258,N_676);
or U2134 (N_2134,N_25,N_211);
nor U2135 (N_2135,N_847,N_184);
nor U2136 (N_2136,N_1204,N_107);
nor U2137 (N_2137,N_249,N_543);
xnor U2138 (N_2138,N_259,N_365);
or U2139 (N_2139,N_1217,N_1176);
and U2140 (N_2140,N_1346,N_595);
nor U2141 (N_2141,N_1422,N_1220);
xor U2142 (N_2142,N_37,N_548);
nor U2143 (N_2143,N_1017,N_492);
or U2144 (N_2144,N_1200,N_1012);
xnor U2145 (N_2145,N_928,N_672);
xor U2146 (N_2146,N_728,N_463);
and U2147 (N_2147,N_148,N_1118);
nand U2148 (N_2148,N_1283,N_398);
and U2149 (N_2149,N_869,N_408);
xnor U2150 (N_2150,N_653,N_1159);
nor U2151 (N_2151,N_627,N_338);
or U2152 (N_2152,N_958,N_1216);
xor U2153 (N_2153,N_1402,N_575);
nand U2154 (N_2154,N_1486,N_1083);
or U2155 (N_2155,N_1343,N_628);
xor U2156 (N_2156,N_85,N_648);
xnor U2157 (N_2157,N_337,N_179);
and U2158 (N_2158,N_181,N_547);
and U2159 (N_2159,N_1433,N_480);
or U2160 (N_2160,N_324,N_745);
and U2161 (N_2161,N_1365,N_332);
nand U2162 (N_2162,N_167,N_227);
nand U2163 (N_2163,N_1406,N_799);
nor U2164 (N_2164,N_1263,N_427);
xor U2165 (N_2165,N_1038,N_1472);
and U2166 (N_2166,N_485,N_1042);
nand U2167 (N_2167,N_577,N_330);
and U2168 (N_2168,N_241,N_1234);
nand U2169 (N_2169,N_1304,N_973);
or U2170 (N_2170,N_411,N_535);
xnor U2171 (N_2171,N_311,N_1372);
nand U2172 (N_2172,N_122,N_1364);
and U2173 (N_2173,N_686,N_889);
and U2174 (N_2174,N_350,N_1167);
and U2175 (N_2175,N_1259,N_1488);
xnor U2176 (N_2176,N_1327,N_1137);
nand U2177 (N_2177,N_1079,N_393);
or U2178 (N_2178,N_680,N_200);
or U2179 (N_2179,N_574,N_132);
and U2180 (N_2180,N_935,N_1319);
nand U2181 (N_2181,N_1483,N_1209);
nor U2182 (N_2182,N_510,N_717);
nand U2183 (N_2183,N_815,N_603);
nand U2184 (N_2184,N_8,N_794);
or U2185 (N_2185,N_617,N_354);
nand U2186 (N_2186,N_636,N_109);
and U2187 (N_2187,N_757,N_260);
xnor U2188 (N_2188,N_585,N_763);
nor U2189 (N_2189,N_529,N_713);
nor U2190 (N_2190,N_139,N_670);
and U2191 (N_2191,N_730,N_508);
or U2192 (N_2192,N_1031,N_526);
nand U2193 (N_2193,N_69,N_924);
and U2194 (N_2194,N_1119,N_1401);
nor U2195 (N_2195,N_419,N_808);
xor U2196 (N_2196,N_487,N_589);
nand U2197 (N_2197,N_1496,N_515);
or U2198 (N_2198,N_235,N_1132);
xnor U2199 (N_2199,N_360,N_300);
xor U2200 (N_2200,N_218,N_315);
nor U2201 (N_2201,N_724,N_342);
or U2202 (N_2202,N_1030,N_172);
and U2203 (N_2203,N_824,N_1498);
xor U2204 (N_2204,N_275,N_625);
and U2205 (N_2205,N_823,N_806);
xor U2206 (N_2206,N_396,N_1189);
or U2207 (N_2207,N_444,N_993);
xnor U2208 (N_2208,N_1066,N_1314);
nand U2209 (N_2209,N_1208,N_566);
nand U2210 (N_2210,N_1348,N_965);
nand U2211 (N_2211,N_1055,N_827);
or U2212 (N_2212,N_934,N_678);
or U2213 (N_2213,N_340,N_378);
or U2214 (N_2214,N_1056,N_1111);
and U2215 (N_2215,N_963,N_741);
and U2216 (N_2216,N_1265,N_946);
nor U2217 (N_2217,N_831,N_557);
nor U2218 (N_2218,N_587,N_130);
xnor U2219 (N_2219,N_1113,N_79);
xor U2220 (N_2220,N_1482,N_438);
xor U2221 (N_2221,N_115,N_473);
and U2222 (N_2222,N_1,N_497);
and U2223 (N_2223,N_866,N_285);
and U2224 (N_2224,N_501,N_1145);
nand U2225 (N_2225,N_789,N_128);
nor U2226 (N_2226,N_304,N_660);
xnor U2227 (N_2227,N_897,N_1106);
nand U2228 (N_2228,N_1181,N_609);
or U2229 (N_2229,N_1212,N_531);
xnor U2230 (N_2230,N_669,N_1425);
or U2231 (N_2231,N_1374,N_1190);
and U2232 (N_2232,N_1296,N_1081);
nand U2233 (N_2233,N_1363,N_836);
xor U2234 (N_2234,N_860,N_1040);
or U2235 (N_2235,N_509,N_1169);
and U2236 (N_2236,N_40,N_639);
or U2237 (N_2237,N_352,N_1008);
and U2238 (N_2238,N_1347,N_555);
nor U2239 (N_2239,N_1033,N_707);
and U2240 (N_2240,N_34,N_1417);
or U2241 (N_2241,N_911,N_723);
nor U2242 (N_2242,N_904,N_1178);
nand U2243 (N_2243,N_102,N_1086);
xnor U2244 (N_2244,N_50,N_729);
or U2245 (N_2245,N_541,N_983);
and U2246 (N_2246,N_341,N_629);
and U2247 (N_2247,N_417,N_614);
and U2248 (N_2248,N_579,N_346);
and U2249 (N_2249,N_171,N_1186);
xor U2250 (N_2250,N_894,N_483);
nand U2251 (N_2251,N_911,N_1358);
nand U2252 (N_2252,N_744,N_858);
xor U2253 (N_2253,N_1348,N_1451);
nand U2254 (N_2254,N_1329,N_1295);
or U2255 (N_2255,N_1100,N_648);
nor U2256 (N_2256,N_225,N_1197);
xnor U2257 (N_2257,N_1069,N_957);
nor U2258 (N_2258,N_1255,N_1338);
nand U2259 (N_2259,N_222,N_274);
nor U2260 (N_2260,N_263,N_561);
nand U2261 (N_2261,N_398,N_625);
and U2262 (N_2262,N_1498,N_1114);
or U2263 (N_2263,N_956,N_873);
xor U2264 (N_2264,N_308,N_1189);
nor U2265 (N_2265,N_486,N_1121);
nor U2266 (N_2266,N_1284,N_699);
or U2267 (N_2267,N_605,N_520);
nor U2268 (N_2268,N_1394,N_1108);
xnor U2269 (N_2269,N_578,N_1354);
or U2270 (N_2270,N_1343,N_225);
and U2271 (N_2271,N_366,N_1437);
nor U2272 (N_2272,N_220,N_992);
and U2273 (N_2273,N_1029,N_696);
and U2274 (N_2274,N_864,N_1223);
nand U2275 (N_2275,N_1170,N_561);
nand U2276 (N_2276,N_784,N_307);
and U2277 (N_2277,N_609,N_140);
nand U2278 (N_2278,N_953,N_103);
and U2279 (N_2279,N_440,N_808);
or U2280 (N_2280,N_867,N_458);
nor U2281 (N_2281,N_920,N_1049);
nand U2282 (N_2282,N_785,N_1407);
xor U2283 (N_2283,N_574,N_355);
nor U2284 (N_2284,N_1256,N_134);
or U2285 (N_2285,N_1341,N_837);
nand U2286 (N_2286,N_479,N_1429);
nand U2287 (N_2287,N_1196,N_1172);
xnor U2288 (N_2288,N_363,N_762);
or U2289 (N_2289,N_1407,N_350);
or U2290 (N_2290,N_889,N_1053);
nand U2291 (N_2291,N_1248,N_1082);
nand U2292 (N_2292,N_180,N_598);
nor U2293 (N_2293,N_497,N_1462);
and U2294 (N_2294,N_1264,N_761);
nand U2295 (N_2295,N_779,N_807);
and U2296 (N_2296,N_170,N_1013);
and U2297 (N_2297,N_548,N_1226);
or U2298 (N_2298,N_1040,N_1141);
xnor U2299 (N_2299,N_805,N_1044);
nand U2300 (N_2300,N_1004,N_667);
xor U2301 (N_2301,N_508,N_822);
and U2302 (N_2302,N_709,N_1460);
nor U2303 (N_2303,N_562,N_1412);
nor U2304 (N_2304,N_1387,N_134);
or U2305 (N_2305,N_1284,N_240);
nor U2306 (N_2306,N_639,N_300);
or U2307 (N_2307,N_804,N_962);
and U2308 (N_2308,N_672,N_598);
nor U2309 (N_2309,N_1491,N_1361);
and U2310 (N_2310,N_561,N_974);
and U2311 (N_2311,N_844,N_181);
xnor U2312 (N_2312,N_1113,N_961);
nor U2313 (N_2313,N_390,N_1485);
or U2314 (N_2314,N_429,N_708);
nor U2315 (N_2315,N_1013,N_1027);
or U2316 (N_2316,N_675,N_563);
nand U2317 (N_2317,N_201,N_2);
or U2318 (N_2318,N_762,N_734);
xnor U2319 (N_2319,N_673,N_406);
and U2320 (N_2320,N_1222,N_1472);
xnor U2321 (N_2321,N_566,N_573);
nor U2322 (N_2322,N_335,N_1109);
and U2323 (N_2323,N_1052,N_525);
and U2324 (N_2324,N_1264,N_301);
nor U2325 (N_2325,N_1420,N_194);
or U2326 (N_2326,N_1421,N_255);
nor U2327 (N_2327,N_553,N_338);
xor U2328 (N_2328,N_1403,N_451);
nand U2329 (N_2329,N_1476,N_142);
nand U2330 (N_2330,N_1423,N_202);
nor U2331 (N_2331,N_694,N_660);
or U2332 (N_2332,N_1300,N_984);
nand U2333 (N_2333,N_877,N_640);
xnor U2334 (N_2334,N_369,N_914);
xor U2335 (N_2335,N_1405,N_49);
xnor U2336 (N_2336,N_1425,N_41);
nand U2337 (N_2337,N_548,N_709);
nand U2338 (N_2338,N_1085,N_59);
or U2339 (N_2339,N_804,N_83);
and U2340 (N_2340,N_628,N_951);
nand U2341 (N_2341,N_320,N_1412);
nand U2342 (N_2342,N_443,N_1185);
nor U2343 (N_2343,N_1032,N_935);
or U2344 (N_2344,N_344,N_186);
nor U2345 (N_2345,N_49,N_190);
nand U2346 (N_2346,N_815,N_507);
or U2347 (N_2347,N_1307,N_774);
nand U2348 (N_2348,N_1079,N_1099);
xor U2349 (N_2349,N_820,N_1015);
nor U2350 (N_2350,N_1436,N_1146);
xnor U2351 (N_2351,N_1172,N_435);
and U2352 (N_2352,N_799,N_1375);
or U2353 (N_2353,N_1439,N_1332);
nand U2354 (N_2354,N_103,N_68);
nand U2355 (N_2355,N_145,N_1102);
nand U2356 (N_2356,N_533,N_787);
nand U2357 (N_2357,N_1232,N_974);
and U2358 (N_2358,N_550,N_169);
or U2359 (N_2359,N_425,N_516);
or U2360 (N_2360,N_907,N_380);
and U2361 (N_2361,N_286,N_467);
xor U2362 (N_2362,N_150,N_358);
nor U2363 (N_2363,N_172,N_408);
xor U2364 (N_2364,N_1019,N_956);
or U2365 (N_2365,N_217,N_37);
xnor U2366 (N_2366,N_919,N_339);
nand U2367 (N_2367,N_512,N_633);
or U2368 (N_2368,N_1345,N_650);
xnor U2369 (N_2369,N_388,N_1459);
and U2370 (N_2370,N_1229,N_44);
and U2371 (N_2371,N_39,N_1276);
xor U2372 (N_2372,N_229,N_187);
and U2373 (N_2373,N_387,N_895);
xnor U2374 (N_2374,N_1051,N_323);
xnor U2375 (N_2375,N_78,N_303);
and U2376 (N_2376,N_411,N_313);
or U2377 (N_2377,N_552,N_612);
xor U2378 (N_2378,N_536,N_744);
nor U2379 (N_2379,N_1192,N_1332);
and U2380 (N_2380,N_925,N_848);
or U2381 (N_2381,N_265,N_684);
xor U2382 (N_2382,N_1479,N_973);
xnor U2383 (N_2383,N_350,N_1073);
nand U2384 (N_2384,N_336,N_177);
nand U2385 (N_2385,N_1288,N_1447);
nand U2386 (N_2386,N_557,N_112);
nand U2387 (N_2387,N_1339,N_1025);
and U2388 (N_2388,N_825,N_47);
and U2389 (N_2389,N_1390,N_208);
nor U2390 (N_2390,N_422,N_1429);
or U2391 (N_2391,N_740,N_251);
nor U2392 (N_2392,N_1341,N_1429);
xnor U2393 (N_2393,N_88,N_771);
xor U2394 (N_2394,N_675,N_297);
xor U2395 (N_2395,N_802,N_882);
xor U2396 (N_2396,N_1458,N_235);
nand U2397 (N_2397,N_279,N_1381);
and U2398 (N_2398,N_1294,N_1485);
nor U2399 (N_2399,N_1497,N_765);
xor U2400 (N_2400,N_1234,N_546);
or U2401 (N_2401,N_651,N_1163);
and U2402 (N_2402,N_659,N_119);
nor U2403 (N_2403,N_1434,N_454);
and U2404 (N_2404,N_1494,N_1199);
nand U2405 (N_2405,N_895,N_1375);
nor U2406 (N_2406,N_1117,N_297);
or U2407 (N_2407,N_1220,N_1257);
nor U2408 (N_2408,N_617,N_875);
xor U2409 (N_2409,N_1130,N_82);
and U2410 (N_2410,N_362,N_140);
and U2411 (N_2411,N_844,N_644);
or U2412 (N_2412,N_899,N_22);
nand U2413 (N_2413,N_544,N_182);
nor U2414 (N_2414,N_870,N_1307);
and U2415 (N_2415,N_863,N_386);
and U2416 (N_2416,N_1198,N_1456);
nand U2417 (N_2417,N_1348,N_1447);
and U2418 (N_2418,N_995,N_3);
and U2419 (N_2419,N_97,N_902);
or U2420 (N_2420,N_1488,N_573);
xnor U2421 (N_2421,N_1482,N_1394);
xor U2422 (N_2422,N_635,N_620);
or U2423 (N_2423,N_960,N_627);
nor U2424 (N_2424,N_1323,N_1203);
xor U2425 (N_2425,N_630,N_745);
nor U2426 (N_2426,N_437,N_252);
xor U2427 (N_2427,N_528,N_274);
or U2428 (N_2428,N_909,N_635);
xor U2429 (N_2429,N_122,N_376);
and U2430 (N_2430,N_421,N_916);
or U2431 (N_2431,N_1430,N_1460);
or U2432 (N_2432,N_466,N_591);
nand U2433 (N_2433,N_30,N_1418);
or U2434 (N_2434,N_225,N_562);
or U2435 (N_2435,N_1071,N_837);
or U2436 (N_2436,N_414,N_246);
and U2437 (N_2437,N_1022,N_1337);
nor U2438 (N_2438,N_1494,N_492);
nand U2439 (N_2439,N_119,N_678);
xor U2440 (N_2440,N_1204,N_24);
or U2441 (N_2441,N_181,N_1022);
and U2442 (N_2442,N_850,N_662);
and U2443 (N_2443,N_1329,N_667);
and U2444 (N_2444,N_907,N_293);
nand U2445 (N_2445,N_857,N_444);
or U2446 (N_2446,N_522,N_549);
or U2447 (N_2447,N_619,N_214);
and U2448 (N_2448,N_422,N_533);
nand U2449 (N_2449,N_366,N_755);
nor U2450 (N_2450,N_416,N_707);
nor U2451 (N_2451,N_875,N_934);
nor U2452 (N_2452,N_763,N_845);
or U2453 (N_2453,N_310,N_400);
xnor U2454 (N_2454,N_113,N_398);
or U2455 (N_2455,N_397,N_463);
or U2456 (N_2456,N_413,N_1378);
nor U2457 (N_2457,N_796,N_1162);
or U2458 (N_2458,N_1347,N_1100);
xnor U2459 (N_2459,N_234,N_695);
nand U2460 (N_2460,N_1415,N_903);
xnor U2461 (N_2461,N_1380,N_387);
nand U2462 (N_2462,N_1008,N_1047);
nand U2463 (N_2463,N_1311,N_620);
or U2464 (N_2464,N_30,N_618);
and U2465 (N_2465,N_340,N_215);
xor U2466 (N_2466,N_1169,N_120);
and U2467 (N_2467,N_394,N_362);
or U2468 (N_2468,N_1024,N_587);
and U2469 (N_2469,N_165,N_831);
nor U2470 (N_2470,N_1487,N_791);
xor U2471 (N_2471,N_274,N_784);
nand U2472 (N_2472,N_1184,N_387);
xnor U2473 (N_2473,N_839,N_700);
nor U2474 (N_2474,N_1113,N_759);
or U2475 (N_2475,N_703,N_542);
or U2476 (N_2476,N_604,N_43);
or U2477 (N_2477,N_1096,N_607);
nor U2478 (N_2478,N_762,N_607);
or U2479 (N_2479,N_172,N_1353);
nand U2480 (N_2480,N_377,N_227);
xor U2481 (N_2481,N_231,N_176);
or U2482 (N_2482,N_1138,N_1426);
and U2483 (N_2483,N_731,N_765);
and U2484 (N_2484,N_1008,N_1301);
and U2485 (N_2485,N_1428,N_583);
nand U2486 (N_2486,N_965,N_530);
nor U2487 (N_2487,N_1065,N_1162);
xnor U2488 (N_2488,N_151,N_159);
or U2489 (N_2489,N_708,N_764);
nand U2490 (N_2490,N_306,N_595);
xnor U2491 (N_2491,N_1493,N_650);
and U2492 (N_2492,N_555,N_203);
or U2493 (N_2493,N_1460,N_916);
and U2494 (N_2494,N_1132,N_5);
and U2495 (N_2495,N_949,N_444);
nor U2496 (N_2496,N_517,N_808);
and U2497 (N_2497,N_61,N_943);
xnor U2498 (N_2498,N_168,N_1247);
nor U2499 (N_2499,N_481,N_42);
nor U2500 (N_2500,N_721,N_101);
nand U2501 (N_2501,N_100,N_852);
xor U2502 (N_2502,N_1232,N_448);
or U2503 (N_2503,N_776,N_1484);
and U2504 (N_2504,N_1025,N_1204);
or U2505 (N_2505,N_755,N_126);
xor U2506 (N_2506,N_511,N_398);
or U2507 (N_2507,N_1407,N_1164);
and U2508 (N_2508,N_1313,N_1427);
or U2509 (N_2509,N_73,N_850);
and U2510 (N_2510,N_46,N_1351);
nor U2511 (N_2511,N_454,N_1193);
and U2512 (N_2512,N_524,N_1275);
nor U2513 (N_2513,N_101,N_590);
and U2514 (N_2514,N_636,N_403);
xor U2515 (N_2515,N_1438,N_990);
xnor U2516 (N_2516,N_1350,N_166);
nor U2517 (N_2517,N_1089,N_243);
or U2518 (N_2518,N_1091,N_1333);
nand U2519 (N_2519,N_1223,N_8);
nor U2520 (N_2520,N_1423,N_1280);
nand U2521 (N_2521,N_68,N_158);
nand U2522 (N_2522,N_1198,N_286);
xnor U2523 (N_2523,N_1395,N_721);
nand U2524 (N_2524,N_376,N_1440);
xnor U2525 (N_2525,N_515,N_752);
and U2526 (N_2526,N_389,N_1337);
or U2527 (N_2527,N_195,N_1065);
and U2528 (N_2528,N_869,N_358);
or U2529 (N_2529,N_1435,N_1408);
xor U2530 (N_2530,N_1194,N_1199);
nand U2531 (N_2531,N_507,N_605);
nor U2532 (N_2532,N_979,N_306);
or U2533 (N_2533,N_1223,N_10);
nand U2534 (N_2534,N_1325,N_68);
nand U2535 (N_2535,N_9,N_1164);
or U2536 (N_2536,N_808,N_102);
or U2537 (N_2537,N_1024,N_1293);
nand U2538 (N_2538,N_1270,N_965);
xor U2539 (N_2539,N_588,N_689);
and U2540 (N_2540,N_972,N_426);
xor U2541 (N_2541,N_934,N_110);
or U2542 (N_2542,N_534,N_903);
and U2543 (N_2543,N_959,N_547);
nor U2544 (N_2544,N_1232,N_1468);
or U2545 (N_2545,N_1164,N_250);
xor U2546 (N_2546,N_330,N_1020);
xor U2547 (N_2547,N_174,N_414);
or U2548 (N_2548,N_240,N_468);
xnor U2549 (N_2549,N_1468,N_886);
xnor U2550 (N_2550,N_1047,N_969);
and U2551 (N_2551,N_225,N_1286);
and U2552 (N_2552,N_933,N_847);
and U2553 (N_2553,N_144,N_778);
nand U2554 (N_2554,N_1310,N_116);
xor U2555 (N_2555,N_1376,N_546);
xor U2556 (N_2556,N_523,N_356);
nand U2557 (N_2557,N_1079,N_794);
nand U2558 (N_2558,N_851,N_495);
xnor U2559 (N_2559,N_1331,N_846);
nand U2560 (N_2560,N_1164,N_1420);
or U2561 (N_2561,N_1247,N_664);
and U2562 (N_2562,N_757,N_970);
nand U2563 (N_2563,N_885,N_1018);
xnor U2564 (N_2564,N_132,N_790);
or U2565 (N_2565,N_1049,N_869);
and U2566 (N_2566,N_207,N_1001);
nand U2567 (N_2567,N_253,N_1015);
or U2568 (N_2568,N_1466,N_609);
and U2569 (N_2569,N_1464,N_1314);
and U2570 (N_2570,N_1485,N_590);
or U2571 (N_2571,N_1450,N_726);
xnor U2572 (N_2572,N_1315,N_41);
or U2573 (N_2573,N_434,N_1383);
xnor U2574 (N_2574,N_826,N_1273);
nor U2575 (N_2575,N_571,N_868);
xnor U2576 (N_2576,N_837,N_1078);
and U2577 (N_2577,N_565,N_980);
nor U2578 (N_2578,N_598,N_250);
xnor U2579 (N_2579,N_596,N_1166);
or U2580 (N_2580,N_666,N_871);
or U2581 (N_2581,N_689,N_439);
and U2582 (N_2582,N_251,N_989);
nand U2583 (N_2583,N_780,N_1031);
nor U2584 (N_2584,N_793,N_1158);
nor U2585 (N_2585,N_286,N_1129);
nor U2586 (N_2586,N_736,N_609);
nand U2587 (N_2587,N_894,N_0);
or U2588 (N_2588,N_653,N_819);
xnor U2589 (N_2589,N_157,N_617);
xnor U2590 (N_2590,N_905,N_101);
and U2591 (N_2591,N_838,N_1254);
nand U2592 (N_2592,N_624,N_935);
nand U2593 (N_2593,N_492,N_781);
xnor U2594 (N_2594,N_1083,N_1491);
xor U2595 (N_2595,N_11,N_1068);
and U2596 (N_2596,N_1339,N_1302);
and U2597 (N_2597,N_630,N_610);
nor U2598 (N_2598,N_224,N_773);
xnor U2599 (N_2599,N_805,N_1072);
nand U2600 (N_2600,N_1451,N_90);
xnor U2601 (N_2601,N_865,N_227);
or U2602 (N_2602,N_593,N_754);
and U2603 (N_2603,N_1451,N_370);
or U2604 (N_2604,N_1327,N_227);
or U2605 (N_2605,N_774,N_1355);
nor U2606 (N_2606,N_1403,N_197);
xnor U2607 (N_2607,N_584,N_233);
and U2608 (N_2608,N_258,N_1046);
xnor U2609 (N_2609,N_389,N_1345);
xor U2610 (N_2610,N_509,N_1255);
and U2611 (N_2611,N_365,N_1406);
and U2612 (N_2612,N_1345,N_746);
or U2613 (N_2613,N_632,N_280);
nor U2614 (N_2614,N_1235,N_421);
xnor U2615 (N_2615,N_898,N_68);
nor U2616 (N_2616,N_1137,N_605);
nor U2617 (N_2617,N_98,N_1194);
xor U2618 (N_2618,N_840,N_735);
xnor U2619 (N_2619,N_1313,N_221);
and U2620 (N_2620,N_1160,N_663);
and U2621 (N_2621,N_341,N_1484);
nand U2622 (N_2622,N_115,N_875);
xor U2623 (N_2623,N_1211,N_62);
or U2624 (N_2624,N_717,N_1079);
nand U2625 (N_2625,N_413,N_1195);
xor U2626 (N_2626,N_333,N_820);
or U2627 (N_2627,N_337,N_159);
and U2628 (N_2628,N_1444,N_772);
nand U2629 (N_2629,N_434,N_733);
nor U2630 (N_2630,N_247,N_393);
nand U2631 (N_2631,N_117,N_1333);
xor U2632 (N_2632,N_271,N_125);
and U2633 (N_2633,N_371,N_814);
and U2634 (N_2634,N_401,N_942);
nor U2635 (N_2635,N_1183,N_544);
and U2636 (N_2636,N_376,N_283);
nand U2637 (N_2637,N_968,N_248);
nand U2638 (N_2638,N_1053,N_1003);
nand U2639 (N_2639,N_664,N_156);
nor U2640 (N_2640,N_1231,N_220);
nor U2641 (N_2641,N_276,N_1208);
nand U2642 (N_2642,N_1355,N_1179);
nor U2643 (N_2643,N_705,N_473);
nor U2644 (N_2644,N_386,N_1254);
xnor U2645 (N_2645,N_1264,N_1305);
xnor U2646 (N_2646,N_321,N_722);
xor U2647 (N_2647,N_260,N_219);
nand U2648 (N_2648,N_743,N_784);
or U2649 (N_2649,N_525,N_399);
xor U2650 (N_2650,N_1081,N_843);
nand U2651 (N_2651,N_372,N_772);
and U2652 (N_2652,N_158,N_121);
xor U2653 (N_2653,N_267,N_924);
or U2654 (N_2654,N_249,N_532);
nor U2655 (N_2655,N_863,N_1223);
nand U2656 (N_2656,N_718,N_910);
and U2657 (N_2657,N_820,N_45);
and U2658 (N_2658,N_330,N_611);
xnor U2659 (N_2659,N_896,N_613);
nor U2660 (N_2660,N_1231,N_110);
nand U2661 (N_2661,N_1,N_1481);
nand U2662 (N_2662,N_472,N_912);
nand U2663 (N_2663,N_958,N_791);
xnor U2664 (N_2664,N_393,N_1384);
xor U2665 (N_2665,N_102,N_1265);
xor U2666 (N_2666,N_734,N_68);
and U2667 (N_2667,N_776,N_252);
nor U2668 (N_2668,N_1402,N_608);
and U2669 (N_2669,N_1440,N_354);
and U2670 (N_2670,N_1340,N_640);
and U2671 (N_2671,N_261,N_173);
or U2672 (N_2672,N_490,N_1294);
xor U2673 (N_2673,N_1176,N_82);
xor U2674 (N_2674,N_162,N_499);
or U2675 (N_2675,N_433,N_39);
nand U2676 (N_2676,N_511,N_178);
nor U2677 (N_2677,N_478,N_1301);
xor U2678 (N_2678,N_680,N_917);
nor U2679 (N_2679,N_453,N_924);
xor U2680 (N_2680,N_1106,N_339);
xnor U2681 (N_2681,N_1037,N_1099);
nor U2682 (N_2682,N_276,N_1224);
or U2683 (N_2683,N_982,N_1341);
xor U2684 (N_2684,N_1407,N_338);
nand U2685 (N_2685,N_626,N_488);
nor U2686 (N_2686,N_1102,N_400);
and U2687 (N_2687,N_1495,N_1094);
xnor U2688 (N_2688,N_125,N_1031);
nand U2689 (N_2689,N_664,N_1053);
nand U2690 (N_2690,N_91,N_478);
xnor U2691 (N_2691,N_1167,N_159);
or U2692 (N_2692,N_102,N_1080);
xnor U2693 (N_2693,N_879,N_574);
nor U2694 (N_2694,N_1411,N_199);
or U2695 (N_2695,N_91,N_564);
and U2696 (N_2696,N_179,N_372);
xnor U2697 (N_2697,N_1129,N_1382);
nand U2698 (N_2698,N_970,N_434);
and U2699 (N_2699,N_1249,N_794);
or U2700 (N_2700,N_1219,N_547);
or U2701 (N_2701,N_1413,N_1483);
nand U2702 (N_2702,N_957,N_765);
nand U2703 (N_2703,N_164,N_133);
nor U2704 (N_2704,N_311,N_1430);
nand U2705 (N_2705,N_857,N_191);
xnor U2706 (N_2706,N_269,N_1240);
or U2707 (N_2707,N_1018,N_165);
and U2708 (N_2708,N_414,N_57);
nand U2709 (N_2709,N_653,N_1430);
nor U2710 (N_2710,N_1316,N_682);
nor U2711 (N_2711,N_306,N_1208);
and U2712 (N_2712,N_517,N_947);
or U2713 (N_2713,N_514,N_954);
xnor U2714 (N_2714,N_822,N_518);
xor U2715 (N_2715,N_1368,N_631);
nor U2716 (N_2716,N_63,N_629);
nand U2717 (N_2717,N_1189,N_1242);
and U2718 (N_2718,N_166,N_801);
nor U2719 (N_2719,N_19,N_1357);
nand U2720 (N_2720,N_1102,N_1302);
or U2721 (N_2721,N_698,N_747);
and U2722 (N_2722,N_409,N_204);
nor U2723 (N_2723,N_1340,N_382);
or U2724 (N_2724,N_277,N_582);
nor U2725 (N_2725,N_229,N_660);
or U2726 (N_2726,N_487,N_1111);
xnor U2727 (N_2727,N_980,N_1355);
xnor U2728 (N_2728,N_1096,N_1026);
or U2729 (N_2729,N_1015,N_529);
nor U2730 (N_2730,N_99,N_1010);
nor U2731 (N_2731,N_1106,N_715);
xnor U2732 (N_2732,N_57,N_712);
nor U2733 (N_2733,N_839,N_158);
nor U2734 (N_2734,N_592,N_358);
xor U2735 (N_2735,N_513,N_314);
xor U2736 (N_2736,N_150,N_1174);
and U2737 (N_2737,N_1084,N_1118);
nand U2738 (N_2738,N_983,N_1107);
xor U2739 (N_2739,N_1122,N_294);
nand U2740 (N_2740,N_809,N_987);
and U2741 (N_2741,N_1267,N_240);
and U2742 (N_2742,N_1367,N_364);
or U2743 (N_2743,N_1286,N_457);
nor U2744 (N_2744,N_62,N_286);
xnor U2745 (N_2745,N_1211,N_1371);
and U2746 (N_2746,N_92,N_251);
nand U2747 (N_2747,N_40,N_604);
xnor U2748 (N_2748,N_1200,N_489);
nor U2749 (N_2749,N_980,N_901);
xor U2750 (N_2750,N_569,N_372);
nand U2751 (N_2751,N_1491,N_275);
and U2752 (N_2752,N_1454,N_1480);
nor U2753 (N_2753,N_1089,N_89);
and U2754 (N_2754,N_603,N_1141);
nand U2755 (N_2755,N_1301,N_798);
and U2756 (N_2756,N_754,N_715);
nor U2757 (N_2757,N_1077,N_1294);
and U2758 (N_2758,N_1110,N_873);
nand U2759 (N_2759,N_883,N_1366);
and U2760 (N_2760,N_120,N_269);
nand U2761 (N_2761,N_1473,N_1144);
or U2762 (N_2762,N_1081,N_864);
xor U2763 (N_2763,N_872,N_1209);
or U2764 (N_2764,N_1128,N_715);
and U2765 (N_2765,N_4,N_1402);
xnor U2766 (N_2766,N_1296,N_933);
nor U2767 (N_2767,N_773,N_910);
nand U2768 (N_2768,N_71,N_300);
nand U2769 (N_2769,N_660,N_1315);
nor U2770 (N_2770,N_326,N_1288);
and U2771 (N_2771,N_433,N_1098);
and U2772 (N_2772,N_237,N_475);
and U2773 (N_2773,N_758,N_134);
or U2774 (N_2774,N_745,N_965);
or U2775 (N_2775,N_617,N_885);
or U2776 (N_2776,N_312,N_820);
xor U2777 (N_2777,N_760,N_590);
nor U2778 (N_2778,N_926,N_817);
or U2779 (N_2779,N_1377,N_25);
and U2780 (N_2780,N_574,N_864);
xor U2781 (N_2781,N_764,N_959);
nor U2782 (N_2782,N_1080,N_1046);
xnor U2783 (N_2783,N_418,N_1405);
nor U2784 (N_2784,N_130,N_1366);
nand U2785 (N_2785,N_835,N_867);
nand U2786 (N_2786,N_711,N_293);
and U2787 (N_2787,N_1435,N_466);
and U2788 (N_2788,N_275,N_999);
nand U2789 (N_2789,N_125,N_1015);
nor U2790 (N_2790,N_892,N_77);
nand U2791 (N_2791,N_509,N_1467);
nor U2792 (N_2792,N_964,N_524);
xnor U2793 (N_2793,N_396,N_811);
or U2794 (N_2794,N_1,N_472);
or U2795 (N_2795,N_1286,N_808);
nor U2796 (N_2796,N_1012,N_584);
nor U2797 (N_2797,N_1487,N_551);
or U2798 (N_2798,N_1064,N_277);
nor U2799 (N_2799,N_835,N_1111);
xor U2800 (N_2800,N_180,N_26);
nand U2801 (N_2801,N_961,N_1104);
and U2802 (N_2802,N_648,N_309);
nand U2803 (N_2803,N_618,N_1402);
nor U2804 (N_2804,N_117,N_884);
or U2805 (N_2805,N_776,N_1497);
and U2806 (N_2806,N_695,N_1137);
or U2807 (N_2807,N_337,N_1179);
xnor U2808 (N_2808,N_654,N_914);
nor U2809 (N_2809,N_67,N_96);
nand U2810 (N_2810,N_301,N_594);
nor U2811 (N_2811,N_1483,N_640);
nand U2812 (N_2812,N_906,N_1333);
xnor U2813 (N_2813,N_254,N_55);
and U2814 (N_2814,N_1388,N_1479);
or U2815 (N_2815,N_425,N_685);
xor U2816 (N_2816,N_1088,N_1263);
or U2817 (N_2817,N_1430,N_1095);
or U2818 (N_2818,N_177,N_884);
nor U2819 (N_2819,N_534,N_588);
nand U2820 (N_2820,N_141,N_1482);
nand U2821 (N_2821,N_619,N_633);
or U2822 (N_2822,N_1066,N_1008);
and U2823 (N_2823,N_137,N_1327);
or U2824 (N_2824,N_353,N_653);
nand U2825 (N_2825,N_944,N_1495);
nor U2826 (N_2826,N_1066,N_53);
nor U2827 (N_2827,N_1145,N_456);
nand U2828 (N_2828,N_1177,N_1134);
or U2829 (N_2829,N_1212,N_749);
or U2830 (N_2830,N_1456,N_375);
xor U2831 (N_2831,N_61,N_605);
nand U2832 (N_2832,N_8,N_1173);
or U2833 (N_2833,N_492,N_1251);
xnor U2834 (N_2834,N_1117,N_804);
nand U2835 (N_2835,N_772,N_1333);
and U2836 (N_2836,N_988,N_1271);
nand U2837 (N_2837,N_1192,N_39);
or U2838 (N_2838,N_474,N_1172);
nand U2839 (N_2839,N_185,N_957);
xnor U2840 (N_2840,N_318,N_1316);
xor U2841 (N_2841,N_1066,N_1296);
or U2842 (N_2842,N_240,N_1025);
nand U2843 (N_2843,N_1289,N_204);
and U2844 (N_2844,N_797,N_855);
or U2845 (N_2845,N_1247,N_724);
xnor U2846 (N_2846,N_1278,N_779);
and U2847 (N_2847,N_1102,N_537);
nand U2848 (N_2848,N_883,N_946);
or U2849 (N_2849,N_1086,N_621);
and U2850 (N_2850,N_791,N_429);
nand U2851 (N_2851,N_1215,N_684);
nand U2852 (N_2852,N_463,N_581);
nor U2853 (N_2853,N_359,N_245);
and U2854 (N_2854,N_769,N_1279);
and U2855 (N_2855,N_947,N_219);
xor U2856 (N_2856,N_598,N_1204);
and U2857 (N_2857,N_1442,N_986);
xor U2858 (N_2858,N_1495,N_777);
nand U2859 (N_2859,N_889,N_194);
nor U2860 (N_2860,N_693,N_485);
nand U2861 (N_2861,N_835,N_821);
xor U2862 (N_2862,N_210,N_1365);
or U2863 (N_2863,N_1378,N_817);
nand U2864 (N_2864,N_250,N_371);
and U2865 (N_2865,N_1269,N_247);
or U2866 (N_2866,N_596,N_36);
nand U2867 (N_2867,N_865,N_1373);
nand U2868 (N_2868,N_1224,N_424);
and U2869 (N_2869,N_348,N_989);
and U2870 (N_2870,N_668,N_1446);
nor U2871 (N_2871,N_320,N_551);
nor U2872 (N_2872,N_783,N_559);
or U2873 (N_2873,N_1358,N_350);
nor U2874 (N_2874,N_1016,N_41);
xor U2875 (N_2875,N_37,N_466);
and U2876 (N_2876,N_748,N_876);
nor U2877 (N_2877,N_1325,N_399);
nand U2878 (N_2878,N_516,N_1459);
and U2879 (N_2879,N_554,N_885);
nor U2880 (N_2880,N_812,N_196);
nand U2881 (N_2881,N_431,N_1221);
xor U2882 (N_2882,N_325,N_90);
or U2883 (N_2883,N_677,N_1387);
xor U2884 (N_2884,N_1132,N_1003);
nand U2885 (N_2885,N_1343,N_1127);
or U2886 (N_2886,N_887,N_154);
and U2887 (N_2887,N_558,N_896);
and U2888 (N_2888,N_1053,N_1152);
xnor U2889 (N_2889,N_955,N_1225);
or U2890 (N_2890,N_674,N_940);
and U2891 (N_2891,N_821,N_976);
nand U2892 (N_2892,N_1166,N_1105);
nor U2893 (N_2893,N_496,N_398);
and U2894 (N_2894,N_518,N_793);
xor U2895 (N_2895,N_414,N_1480);
or U2896 (N_2896,N_725,N_392);
xor U2897 (N_2897,N_808,N_127);
or U2898 (N_2898,N_794,N_35);
and U2899 (N_2899,N_577,N_1102);
nor U2900 (N_2900,N_820,N_514);
nand U2901 (N_2901,N_1210,N_498);
and U2902 (N_2902,N_1418,N_1454);
nor U2903 (N_2903,N_1317,N_468);
and U2904 (N_2904,N_1399,N_1257);
xnor U2905 (N_2905,N_1105,N_1013);
and U2906 (N_2906,N_509,N_1496);
or U2907 (N_2907,N_1185,N_1468);
nand U2908 (N_2908,N_1077,N_803);
or U2909 (N_2909,N_396,N_628);
or U2910 (N_2910,N_1100,N_284);
and U2911 (N_2911,N_1218,N_650);
nor U2912 (N_2912,N_145,N_1177);
nand U2913 (N_2913,N_671,N_1220);
nor U2914 (N_2914,N_1451,N_1384);
or U2915 (N_2915,N_979,N_1100);
xnor U2916 (N_2916,N_1401,N_633);
nand U2917 (N_2917,N_1426,N_1428);
or U2918 (N_2918,N_73,N_391);
and U2919 (N_2919,N_296,N_297);
and U2920 (N_2920,N_692,N_391);
and U2921 (N_2921,N_1393,N_207);
or U2922 (N_2922,N_1277,N_928);
or U2923 (N_2923,N_612,N_1144);
nand U2924 (N_2924,N_1181,N_427);
or U2925 (N_2925,N_659,N_667);
xnor U2926 (N_2926,N_264,N_959);
nand U2927 (N_2927,N_914,N_545);
xor U2928 (N_2928,N_813,N_116);
nand U2929 (N_2929,N_557,N_1104);
xnor U2930 (N_2930,N_1075,N_579);
nor U2931 (N_2931,N_749,N_658);
nand U2932 (N_2932,N_42,N_520);
xnor U2933 (N_2933,N_130,N_501);
xnor U2934 (N_2934,N_385,N_93);
or U2935 (N_2935,N_503,N_1199);
nand U2936 (N_2936,N_187,N_696);
or U2937 (N_2937,N_292,N_1208);
xnor U2938 (N_2938,N_1134,N_981);
xnor U2939 (N_2939,N_1249,N_877);
xnor U2940 (N_2940,N_1346,N_1314);
xnor U2941 (N_2941,N_1067,N_322);
nand U2942 (N_2942,N_769,N_1052);
and U2943 (N_2943,N_149,N_256);
nor U2944 (N_2944,N_521,N_411);
and U2945 (N_2945,N_1309,N_1303);
nor U2946 (N_2946,N_1422,N_766);
or U2947 (N_2947,N_1338,N_952);
or U2948 (N_2948,N_1361,N_757);
and U2949 (N_2949,N_835,N_1291);
xor U2950 (N_2950,N_300,N_488);
xor U2951 (N_2951,N_1177,N_1446);
nand U2952 (N_2952,N_344,N_880);
or U2953 (N_2953,N_891,N_983);
xor U2954 (N_2954,N_1309,N_1200);
and U2955 (N_2955,N_310,N_549);
xor U2956 (N_2956,N_1072,N_1155);
xor U2957 (N_2957,N_1453,N_418);
xor U2958 (N_2958,N_214,N_1050);
nand U2959 (N_2959,N_962,N_625);
nand U2960 (N_2960,N_1276,N_810);
xnor U2961 (N_2961,N_594,N_931);
nor U2962 (N_2962,N_1481,N_24);
and U2963 (N_2963,N_1244,N_679);
nand U2964 (N_2964,N_246,N_1474);
nand U2965 (N_2965,N_1112,N_533);
nor U2966 (N_2966,N_1461,N_1033);
nand U2967 (N_2967,N_677,N_13);
or U2968 (N_2968,N_759,N_18);
nor U2969 (N_2969,N_440,N_701);
nor U2970 (N_2970,N_1406,N_166);
or U2971 (N_2971,N_836,N_552);
or U2972 (N_2972,N_1321,N_909);
xnor U2973 (N_2973,N_854,N_1472);
xnor U2974 (N_2974,N_1169,N_924);
or U2975 (N_2975,N_872,N_103);
nand U2976 (N_2976,N_80,N_1308);
nand U2977 (N_2977,N_527,N_1031);
nand U2978 (N_2978,N_738,N_411);
or U2979 (N_2979,N_564,N_645);
xor U2980 (N_2980,N_77,N_1417);
xnor U2981 (N_2981,N_1030,N_996);
nand U2982 (N_2982,N_465,N_834);
and U2983 (N_2983,N_451,N_754);
and U2984 (N_2984,N_860,N_924);
nor U2985 (N_2985,N_176,N_694);
nand U2986 (N_2986,N_1421,N_1290);
nand U2987 (N_2987,N_784,N_227);
nand U2988 (N_2988,N_1083,N_1009);
nand U2989 (N_2989,N_61,N_1100);
nand U2990 (N_2990,N_848,N_1134);
and U2991 (N_2991,N_32,N_490);
nor U2992 (N_2992,N_195,N_980);
nand U2993 (N_2993,N_592,N_363);
or U2994 (N_2994,N_191,N_271);
nand U2995 (N_2995,N_1329,N_1426);
and U2996 (N_2996,N_153,N_1028);
xor U2997 (N_2997,N_698,N_1441);
and U2998 (N_2998,N_1230,N_393);
and U2999 (N_2999,N_1398,N_365);
xor U3000 (N_3000,N_2950,N_2621);
and U3001 (N_3001,N_2116,N_2643);
and U3002 (N_3002,N_2473,N_2465);
nand U3003 (N_3003,N_2359,N_1589);
nor U3004 (N_3004,N_2449,N_2106);
nor U3005 (N_3005,N_2401,N_2934);
nand U3006 (N_3006,N_2572,N_2534);
nand U3007 (N_3007,N_2707,N_2113);
nand U3008 (N_3008,N_2609,N_1931);
xor U3009 (N_3009,N_2331,N_2618);
xor U3010 (N_3010,N_2515,N_2959);
or U3011 (N_3011,N_1746,N_2144);
xor U3012 (N_3012,N_1677,N_2670);
nand U3013 (N_3013,N_2311,N_1747);
and U3014 (N_3014,N_1606,N_2952);
nor U3015 (N_3015,N_1961,N_2900);
and U3016 (N_3016,N_2591,N_1713);
and U3017 (N_3017,N_2736,N_1521);
and U3018 (N_3018,N_2958,N_1941);
or U3019 (N_3019,N_2564,N_2842);
nor U3020 (N_3020,N_2257,N_2972);
nand U3021 (N_3021,N_2989,N_1624);
xor U3022 (N_3022,N_2565,N_2471);
or U3023 (N_3023,N_1541,N_1987);
or U3024 (N_3024,N_1623,N_2273);
and U3025 (N_3025,N_2576,N_1972);
nand U3026 (N_3026,N_2650,N_2190);
xor U3027 (N_3027,N_2675,N_2852);
nand U3028 (N_3028,N_2503,N_2236);
nand U3029 (N_3029,N_2129,N_2248);
xnor U3030 (N_3030,N_2688,N_2745);
or U3031 (N_3031,N_2508,N_1580);
nand U3032 (N_3032,N_1852,N_2151);
or U3033 (N_3033,N_2255,N_2336);
and U3034 (N_3034,N_2603,N_2747);
or U3035 (N_3035,N_2637,N_2481);
xnor U3036 (N_3036,N_2362,N_2494);
and U3037 (N_3037,N_2325,N_2220);
and U3038 (N_3038,N_1764,N_2810);
xnor U3039 (N_3039,N_1913,N_2376);
xnor U3040 (N_3040,N_1691,N_2077);
and U3041 (N_3041,N_1500,N_1681);
and U3042 (N_3042,N_2601,N_2916);
nand U3043 (N_3043,N_2291,N_2766);
xor U3044 (N_3044,N_2509,N_2974);
nor U3045 (N_3045,N_2356,N_1649);
xor U3046 (N_3046,N_1607,N_1594);
nand U3047 (N_3047,N_2904,N_2804);
nand U3048 (N_3048,N_2991,N_2647);
xor U3049 (N_3049,N_1598,N_2429);
xnor U3050 (N_3050,N_2155,N_2046);
and U3051 (N_3051,N_2094,N_2301);
nand U3052 (N_3052,N_2853,N_2308);
nor U3053 (N_3053,N_1563,N_1978);
nor U3054 (N_3054,N_1809,N_2809);
xor U3055 (N_3055,N_1638,N_1516);
or U3056 (N_3056,N_2548,N_1923);
or U3057 (N_3057,N_2462,N_1816);
nor U3058 (N_3058,N_1576,N_2044);
and U3059 (N_3059,N_1860,N_2890);
xor U3060 (N_3060,N_2138,N_1878);
nand U3061 (N_3061,N_2289,N_1612);
and U3062 (N_3062,N_2612,N_2268);
xnor U3063 (N_3063,N_2798,N_2998);
or U3064 (N_3064,N_2121,N_1502);
nand U3065 (N_3065,N_2474,N_1748);
and U3066 (N_3066,N_1507,N_1896);
xor U3067 (N_3067,N_2568,N_1814);
nor U3068 (N_3068,N_1868,N_1585);
or U3069 (N_3069,N_1633,N_2370);
nor U3070 (N_3070,N_1513,N_2536);
nor U3071 (N_3071,N_2454,N_2379);
and U3072 (N_3072,N_1562,N_2657);
nand U3073 (N_3073,N_2250,N_2286);
or U3074 (N_3074,N_2186,N_1862);
nor U3075 (N_3075,N_2953,N_2872);
and U3076 (N_3076,N_2263,N_2933);
nand U3077 (N_3077,N_1726,N_1900);
nor U3078 (N_3078,N_2394,N_1671);
or U3079 (N_3079,N_1985,N_1737);
and U3080 (N_3080,N_2724,N_2101);
xor U3081 (N_3081,N_2850,N_2856);
xnor U3082 (N_3082,N_2718,N_1722);
or U3083 (N_3083,N_2467,N_1880);
nor U3084 (N_3084,N_1789,N_1718);
and U3085 (N_3085,N_2001,N_2528);
xor U3086 (N_3086,N_2269,N_1924);
nand U3087 (N_3087,N_2491,N_2205);
or U3088 (N_3088,N_2954,N_2924);
and U3089 (N_3089,N_2104,N_2701);
nand U3090 (N_3090,N_1955,N_1772);
xnor U3091 (N_3091,N_2107,N_1905);
nand U3092 (N_3092,N_2170,N_2187);
and U3093 (N_3093,N_2150,N_2658);
xor U3094 (N_3094,N_1518,N_2898);
nand U3095 (N_3095,N_1965,N_2738);
or U3096 (N_3096,N_2585,N_2600);
and U3097 (N_3097,N_1927,N_2351);
xor U3098 (N_3098,N_1794,N_2469);
and U3099 (N_3099,N_1926,N_2669);
or U3100 (N_3100,N_2493,N_2010);
nor U3101 (N_3101,N_2648,N_2789);
and U3102 (N_3102,N_2360,N_1573);
nor U3103 (N_3103,N_1546,N_2247);
nor U3104 (N_3104,N_1835,N_2328);
nor U3105 (N_3105,N_1865,N_2968);
xnor U3106 (N_3106,N_2475,N_2049);
xnor U3107 (N_3107,N_1815,N_2426);
or U3108 (N_3108,N_2277,N_2184);
nor U3109 (N_3109,N_2751,N_2708);
and U3110 (N_3110,N_2870,N_2791);
nor U3111 (N_3111,N_1797,N_1855);
or U3112 (N_3112,N_2605,N_1954);
xor U3113 (N_3113,N_2677,N_2397);
or U3114 (N_3114,N_2721,N_1637);
nor U3115 (N_3115,N_2759,N_2188);
or U3116 (N_3116,N_1720,N_2817);
or U3117 (N_3117,N_1861,N_2499);
xnor U3118 (N_3118,N_1631,N_2782);
xnor U3119 (N_3119,N_1668,N_2667);
nand U3120 (N_3120,N_2369,N_1807);
nand U3121 (N_3121,N_2181,N_1841);
and U3122 (N_3122,N_2278,N_2877);
nand U3123 (N_3123,N_2013,N_1729);
and U3124 (N_3124,N_1949,N_2057);
nor U3125 (N_3125,N_1790,N_2655);
xnor U3126 (N_3126,N_1662,N_2735);
nand U3127 (N_3127,N_2338,N_2073);
or U3128 (N_3128,N_2774,N_2693);
and U3129 (N_3129,N_2540,N_2251);
nand U3130 (N_3130,N_1682,N_1544);
nor U3131 (N_3131,N_1520,N_1572);
nor U3132 (N_3132,N_1577,N_2773);
nand U3133 (N_3133,N_2378,N_2003);
nand U3134 (N_3134,N_2048,N_2552);
nand U3135 (N_3135,N_2395,N_2293);
nand U3136 (N_3136,N_2757,N_2321);
nor U3137 (N_3137,N_2862,N_1917);
xnor U3138 (N_3138,N_2501,N_1626);
nor U3139 (N_3139,N_1916,N_2832);
nand U3140 (N_3140,N_2239,N_2297);
xnor U3141 (N_3141,N_1990,N_2149);
or U3142 (N_3142,N_2694,N_2442);
nor U3143 (N_3143,N_2981,N_1773);
nor U3144 (N_3144,N_2925,N_2796);
nand U3145 (N_3145,N_2119,N_1986);
and U3146 (N_3146,N_1714,N_2267);
xor U3147 (N_3147,N_2203,N_2818);
or U3148 (N_3148,N_2005,N_1539);
nand U3149 (N_3149,N_2302,N_1724);
xor U3150 (N_3150,N_2678,N_1717);
and U3151 (N_3151,N_2713,N_1886);
nor U3152 (N_3152,N_2866,N_2089);
nor U3153 (N_3153,N_2522,N_1937);
and U3154 (N_3154,N_1727,N_2517);
xor U3155 (N_3155,N_1834,N_2533);
nor U3156 (N_3156,N_2771,N_1599);
xnor U3157 (N_3157,N_1586,N_2733);
nand U3158 (N_3158,N_2165,N_1750);
nand U3159 (N_3159,N_2148,N_2802);
xor U3160 (N_3160,N_2445,N_2435);
or U3161 (N_3161,N_2691,N_1540);
and U3162 (N_3162,N_1603,N_2606);
or U3163 (N_3163,N_2995,N_2768);
and U3164 (N_3164,N_2135,N_2711);
and U3165 (N_3165,N_1524,N_2319);
nor U3166 (N_3166,N_2446,N_1575);
or U3167 (N_3167,N_2801,N_2583);
nand U3168 (N_3168,N_1556,N_2452);
xor U3169 (N_3169,N_2537,N_2034);
nor U3170 (N_3170,N_1515,N_2091);
and U3171 (N_3171,N_2207,N_2525);
and U3172 (N_3172,N_2368,N_1695);
or U3173 (N_3173,N_2894,N_1582);
and U3174 (N_3174,N_2000,N_2306);
and U3175 (N_3175,N_2640,N_1509);
nor U3176 (N_3176,N_2416,N_1652);
or U3177 (N_3177,N_2975,N_1596);
and U3178 (N_3178,N_2566,N_1780);
nand U3179 (N_3179,N_2437,N_2324);
or U3180 (N_3180,N_2161,N_1616);
xnor U3181 (N_3181,N_1735,N_2489);
xor U3182 (N_3182,N_1665,N_2593);
nor U3183 (N_3183,N_1592,N_2617);
nand U3184 (N_3184,N_2392,N_2811);
nand U3185 (N_3185,N_2709,N_2276);
and U3186 (N_3186,N_2202,N_2404);
nor U3187 (N_3187,N_2403,N_1538);
nand U3188 (N_3188,N_2743,N_2256);
nor U3189 (N_3189,N_2696,N_2871);
nand U3190 (N_3190,N_1526,N_1553);
and U3191 (N_3191,N_2117,N_1968);
xnor U3192 (N_3192,N_1784,N_2366);
nor U3193 (N_3193,N_1774,N_1688);
and U3194 (N_3194,N_2948,N_2915);
or U3195 (N_3195,N_2619,N_1891);
xnor U3196 (N_3196,N_1762,N_2180);
nand U3197 (N_3197,N_2795,N_2706);
nor U3198 (N_3198,N_2727,N_2663);
and U3199 (N_3199,N_2596,N_1734);
and U3200 (N_3200,N_2420,N_2361);
nand U3201 (N_3201,N_2042,N_2069);
and U3202 (N_3202,N_2892,N_2698);
nand U3203 (N_3203,N_1706,N_2065);
nor U3204 (N_3204,N_1745,N_2532);
xnor U3205 (N_3205,N_2843,N_1622);
nand U3206 (N_3206,N_1890,N_2062);
or U3207 (N_3207,N_2191,N_2938);
xnor U3208 (N_3208,N_2036,N_1543);
nor U3209 (N_3209,N_2122,N_1527);
or U3210 (N_3210,N_2754,N_1699);
xor U3211 (N_3211,N_2635,N_1579);
nand U3212 (N_3212,N_2819,N_2625);
and U3213 (N_3213,N_1545,N_2334);
or U3214 (N_3214,N_2056,N_2805);
and U3215 (N_3215,N_2204,N_2345);
xor U3216 (N_3216,N_2615,N_2799);
and U3217 (N_3217,N_2623,N_1752);
nor U3218 (N_3218,N_2837,N_1531);
and U3219 (N_3219,N_2895,N_1588);
and U3220 (N_3220,N_2216,N_2611);
xor U3221 (N_3221,N_2164,N_1832);
or U3222 (N_3222,N_2851,N_1731);
nor U3223 (N_3223,N_2323,N_1992);
and U3224 (N_3224,N_2407,N_2340);
nand U3225 (N_3225,N_1888,N_2884);
nand U3226 (N_3226,N_2863,N_1966);
nor U3227 (N_3227,N_2982,N_2423);
and U3228 (N_3228,N_1995,N_1758);
nor U3229 (N_3229,N_2422,N_2006);
and U3230 (N_3230,N_2788,N_2405);
nor U3231 (N_3231,N_2039,N_1963);
xnor U3232 (N_3232,N_1889,N_2740);
xor U3233 (N_3233,N_2868,N_2775);
nor U3234 (N_3234,N_1863,N_2127);
nor U3235 (N_3235,N_2758,N_2303);
xnor U3236 (N_3236,N_1853,N_2704);
nand U3237 (N_3237,N_2641,N_2339);
xor U3238 (N_3238,N_1838,N_2573);
and U3239 (N_3239,N_2053,N_2730);
or U3240 (N_3240,N_1604,N_2910);
or U3241 (N_3241,N_2942,N_2919);
xnor U3242 (N_3242,N_2874,N_1519);
nand U3243 (N_3243,N_1974,N_2578);
and U3244 (N_3244,N_1970,N_2189);
and U3245 (N_3245,N_1804,N_1740);
nor U3246 (N_3246,N_2235,N_2285);
nor U3247 (N_3247,N_2020,N_1934);
or U3248 (N_3248,N_2153,N_2451);
nor U3249 (N_3249,N_2438,N_2544);
nor U3250 (N_3250,N_2957,N_2307);
nor U3251 (N_3251,N_1640,N_2440);
or U3252 (N_3252,N_2780,N_2484);
nor U3253 (N_3253,N_2705,N_2133);
or U3254 (N_3254,N_1552,N_2068);
nand U3255 (N_3255,N_1628,N_2026);
and U3256 (N_3256,N_2019,N_1567);
nand U3257 (N_3257,N_2265,N_2719);
and U3258 (N_3258,N_1991,N_2728);
nand U3259 (N_3259,N_2200,N_2364);
xor U3260 (N_3260,N_2608,N_2266);
nand U3261 (N_3261,N_1802,N_2315);
nand U3262 (N_3262,N_2676,N_2487);
nor U3263 (N_3263,N_2906,N_2098);
nand U3264 (N_3264,N_2185,N_2665);
and U3265 (N_3265,N_2059,N_1833);
or U3266 (N_3266,N_2529,N_1897);
and U3267 (N_3267,N_1769,N_2985);
nand U3268 (N_3268,N_2028,N_2283);
or U3269 (N_3269,N_2346,N_2947);
and U3270 (N_3270,N_1581,N_2316);
and U3271 (N_3271,N_2502,N_2622);
xnor U3272 (N_3272,N_1503,N_2914);
or U3273 (N_3273,N_2604,N_2997);
xor U3274 (N_3274,N_2889,N_2146);
and U3275 (N_3275,N_2275,N_2996);
nor U3276 (N_3276,N_2697,N_2342);
or U3277 (N_3277,N_1803,N_2374);
and U3278 (N_3278,N_2715,N_2541);
or U3279 (N_3279,N_2966,N_1754);
xnor U3280 (N_3280,N_2903,N_1997);
xor U3281 (N_3281,N_1756,N_1812);
nor U3282 (N_3282,N_2781,N_2241);
and U3283 (N_3283,N_2222,N_2549);
nor U3284 (N_3284,N_1982,N_2179);
nand U3285 (N_3285,N_1698,N_2031);
or U3286 (N_3286,N_1882,N_2826);
xnor U3287 (N_3287,N_2692,N_1565);
nand U3288 (N_3288,N_2993,N_2546);
nand U3289 (N_3289,N_2777,N_2066);
nor U3290 (N_3290,N_1873,N_2457);
and U3291 (N_3291,N_1919,N_2977);
xor U3292 (N_3292,N_1825,N_2946);
nor U3293 (N_3293,N_2685,N_2383);
nor U3294 (N_3294,N_2274,N_2047);
nor U3295 (N_3295,N_2986,N_1999);
nor U3296 (N_3296,N_1885,N_1843);
or U3297 (N_3297,N_1817,N_2097);
xnor U3298 (N_3298,N_1620,N_2980);
xnor U3299 (N_3299,N_2803,N_1942);
and U3300 (N_3300,N_2720,N_2498);
and U3301 (N_3301,N_2662,N_1736);
and U3302 (N_3302,N_2433,N_2393);
nand U3303 (N_3303,N_2582,N_2074);
xor U3304 (N_3304,N_2105,N_2926);
and U3305 (N_3305,N_1710,N_2602);
xnor U3306 (N_3306,N_1829,N_1898);
nand U3307 (N_3307,N_2761,N_1902);
nor U3308 (N_3308,N_1669,N_1791);
xor U3309 (N_3309,N_2869,N_2830);
or U3310 (N_3310,N_2584,N_1511);
and U3311 (N_3311,N_2159,N_2835);
xnor U3312 (N_3312,N_2058,N_2806);
nand U3313 (N_3313,N_2375,N_2822);
or U3314 (N_3314,N_2299,N_1879);
xnor U3315 (N_3315,N_2626,N_2624);
xor U3316 (N_3316,N_1738,N_2358);
or U3317 (N_3317,N_1667,N_2922);
nand U3318 (N_3318,N_2664,N_2246);
and U3319 (N_3319,N_2237,N_2381);
and U3320 (N_3320,N_1697,N_2110);
nor U3321 (N_3321,N_2973,N_2939);
and U3322 (N_3322,N_1808,N_2660);
or U3323 (N_3323,N_2571,N_2464);
nand U3324 (N_3324,N_2913,N_1508);
and U3325 (N_3325,N_1525,N_2211);
xnor U3326 (N_3326,N_1561,N_2343);
and U3327 (N_3327,N_2710,N_2955);
nand U3328 (N_3328,N_2551,N_1528);
and U3329 (N_3329,N_1950,N_2163);
nor U3330 (N_3330,N_2310,N_1685);
xor U3331 (N_3331,N_1778,N_2787);
nand U3332 (N_3332,N_1884,N_2666);
and U3333 (N_3333,N_1785,N_2518);
or U3334 (N_3334,N_1630,N_2861);
and U3335 (N_3335,N_2849,N_1881);
nand U3336 (N_3336,N_1895,N_2786);
nand U3337 (N_3337,N_2313,N_2304);
nand U3338 (N_3338,N_2553,N_2243);
or U3339 (N_3339,N_2231,N_2168);
xnor U3340 (N_3340,N_2590,N_1981);
and U3341 (N_3341,N_2225,N_2923);
and U3342 (N_3342,N_1887,N_2045);
nor U3343 (N_3343,N_2970,N_2579);
or U3344 (N_3344,N_1989,N_2734);
nor U3345 (N_3345,N_2723,N_2936);
nor U3346 (N_3346,N_1973,N_2260);
nor U3347 (N_3347,N_1583,N_1948);
or U3348 (N_3348,N_2380,N_2907);
or U3349 (N_3349,N_1848,N_1674);
and U3350 (N_3350,N_2638,N_1930);
and U3351 (N_3351,N_2088,N_1940);
nand U3352 (N_3352,N_1979,N_2563);
xor U3353 (N_3353,N_2103,N_2415);
or U3354 (N_3354,N_2654,N_2964);
or U3355 (N_3355,N_1615,N_1798);
xnor U3356 (N_3356,N_1601,N_1811);
nand U3357 (N_3357,N_1828,N_1909);
nor U3358 (N_3358,N_2879,N_2322);
nand U3359 (N_3359,N_1801,N_2009);
nand U3360 (N_3360,N_2102,N_2022);
or U3361 (N_3361,N_2245,N_2167);
and U3362 (N_3362,N_2086,N_2460);
nor U3363 (N_3363,N_2332,N_2002);
nor U3364 (N_3364,N_2253,N_1793);
nor U3365 (N_3365,N_2015,N_2821);
xor U3366 (N_3366,N_1907,N_1823);
and U3367 (N_3367,N_2687,N_2885);
xor U3368 (N_3368,N_2425,N_2613);
or U3369 (N_3369,N_2470,N_2496);
nand U3370 (N_3370,N_2223,N_1864);
nor U3371 (N_3371,N_1639,N_2411);
or U3372 (N_3372,N_1704,N_2838);
nand U3373 (N_3373,N_2545,N_2109);
nand U3374 (N_3374,N_2512,N_1683);
xor U3375 (N_3375,N_1730,N_2586);
and U3376 (N_3376,N_1657,N_2240);
and U3377 (N_3377,N_2037,N_2961);
and U3378 (N_3378,N_2232,N_2447);
or U3379 (N_3379,N_1578,N_2854);
and U3380 (N_3380,N_2506,N_1749);
and U3381 (N_3381,N_2620,N_1787);
and U3382 (N_3382,N_2134,N_2427);
xor U3383 (N_3383,N_2413,N_2535);
nor U3384 (N_3384,N_2547,N_1558);
or U3385 (N_3385,N_2314,N_1943);
nor U3386 (N_3386,N_2215,N_2156);
nor U3387 (N_3387,N_2318,N_2194);
and U3388 (N_3388,N_2949,N_2329);
nand U3389 (N_3389,N_1768,N_1642);
nand U3390 (N_3390,N_1723,N_2388);
nand U3391 (N_3391,N_1799,N_2770);
xnor U3392 (N_3392,N_2330,N_2282);
xnor U3393 (N_3393,N_2399,N_2444);
and U3394 (N_3394,N_2371,N_1693);
nor U3395 (N_3395,N_2032,N_1658);
xnor U3396 (N_3396,N_2505,N_1928);
nand U3397 (N_3397,N_2390,N_2178);
or U3398 (N_3398,N_2254,N_2960);
nand U3399 (N_3399,N_2355,N_1857);
nand U3400 (N_3400,N_2560,N_2929);
nor U3401 (N_3401,N_1532,N_2616);
or U3402 (N_3402,N_1960,N_2114);
xnor U3403 (N_3403,N_2043,N_2279);
or U3404 (N_3404,N_2287,N_2510);
xor U3405 (N_3405,N_2607,N_2384);
nor U3406 (N_3406,N_1851,N_1962);
nand U3407 (N_3407,N_1744,N_2927);
or U3408 (N_3408,N_2305,N_2672);
and U3409 (N_3409,N_2023,N_2417);
nand U3410 (N_3410,N_2944,N_2599);
or U3411 (N_3411,N_2829,N_2999);
nand U3412 (N_3412,N_2259,N_1956);
xor U3413 (N_3413,N_2815,N_2911);
or U3414 (N_3414,N_2466,N_2645);
xnor U3415 (N_3415,N_2406,N_2051);
or U3416 (N_3416,N_2472,N_1732);
and U3417 (N_3417,N_2352,N_1547);
xnor U3418 (N_3418,N_1977,N_2887);
nand U3419 (N_3419,N_1805,N_2206);
xnor U3420 (N_3420,N_2865,N_2271);
nor U3421 (N_3421,N_1783,N_2453);
or U3422 (N_3422,N_1666,N_2531);
and U3423 (N_3423,N_2468,N_2492);
nor U3424 (N_3424,N_1600,N_2965);
nand U3425 (N_3425,N_2176,N_2886);
or U3426 (N_3426,N_1670,N_2382);
xor U3427 (N_3427,N_1921,N_2079);
nor U3428 (N_3428,N_1796,N_2681);
nor U3429 (N_3429,N_2555,N_2507);
nand U3430 (N_3430,N_2524,N_1654);
nor U3431 (N_3431,N_1844,N_2700);
or U3432 (N_3432,N_1757,N_1771);
nor U3433 (N_3433,N_1692,N_2476);
xor U3434 (N_3434,N_1846,N_2831);
xor U3435 (N_3435,N_2410,N_2846);
nor U3436 (N_3436,N_2347,N_2523);
nor U3437 (N_3437,N_1788,N_1703);
or U3438 (N_3438,N_1661,N_1996);
and U3439 (N_3439,N_1554,N_2882);
or U3440 (N_3440,N_1929,N_2908);
and U3441 (N_3441,N_2012,N_1705);
or U3442 (N_3442,N_2050,N_2920);
and U3443 (N_3443,N_2598,N_1593);
xor U3444 (N_3444,N_2350,N_2030);
nand U3445 (N_3445,N_2901,N_2295);
nor U3446 (N_3446,N_1609,N_1935);
xor U3447 (N_3447,N_2177,N_2744);
xnor U3448 (N_3448,N_2095,N_2479);
xor U3449 (N_3449,N_2649,N_2962);
and U3450 (N_3450,N_2902,N_2100);
and U3451 (N_3451,N_1914,N_2632);
nor U3452 (N_3452,N_2940,N_2270);
nand U3453 (N_3453,N_2731,N_2653);
nor U3454 (N_3454,N_2132,N_1920);
and U3455 (N_3455,N_1792,N_1510);
xor U3456 (N_3456,N_1542,N_2642);
nor U3457 (N_3457,N_2941,N_2543);
xor U3458 (N_3458,N_2171,N_2823);
or U3459 (N_3459,N_1651,N_2888);
or U3460 (N_3460,N_1533,N_1877);
xnor U3461 (N_3461,N_2634,N_2880);
nand U3462 (N_3462,N_1663,N_2061);
nor U3463 (N_3463,N_2684,N_2763);
and U3464 (N_3464,N_2441,N_2712);
nand U3465 (N_3465,N_2746,N_2398);
nand U3466 (N_3466,N_2897,N_1911);
nand U3467 (N_3467,N_2800,N_2588);
or U3468 (N_3468,N_1938,N_2480);
nand U3469 (N_3469,N_2716,N_1822);
and U3470 (N_3470,N_1983,N_2514);
and U3471 (N_3471,N_2385,N_2574);
nand U3472 (N_3472,N_1711,N_1910);
and U3473 (N_3473,N_2714,N_2978);
and U3474 (N_3474,N_2418,N_2083);
nand U3475 (N_3475,N_2244,N_2732);
nand U3476 (N_3476,N_1555,N_2595);
xnor U3477 (N_3477,N_1566,N_1632);
or U3478 (N_3478,N_1743,N_2807);
and U3479 (N_3479,N_1522,N_2208);
or U3480 (N_3480,N_2141,N_2118);
nand U3481 (N_3481,N_1587,N_2765);
or U3482 (N_3482,N_2828,N_2414);
or U3483 (N_3483,N_2041,N_2630);
and U3484 (N_3484,N_2227,N_2249);
nand U3485 (N_3485,N_1786,N_1686);
xor U3486 (N_3486,N_1849,N_1850);
nand U3487 (N_3487,N_2883,N_1839);
nand U3488 (N_3488,N_1739,N_2027);
or U3489 (N_3489,N_2813,N_1613);
or U3490 (N_3490,N_1870,N_2071);
nor U3491 (N_3491,N_2157,N_2261);
or U3492 (N_3492,N_1611,N_2482);
xor U3493 (N_3493,N_1715,N_1958);
and U3494 (N_3494,N_2162,N_1994);
nor U3495 (N_3495,N_1529,N_2682);
or U3496 (N_3496,N_1602,N_2386);
and U3497 (N_3497,N_1504,N_2790);
or U3498 (N_3498,N_2126,N_1976);
xor U3499 (N_3499,N_1617,N_2567);
nand U3500 (N_3500,N_2349,N_1776);
nand U3501 (N_3501,N_1619,N_1655);
nor U3502 (N_3502,N_2090,N_1584);
nor U3503 (N_3503,N_2644,N_1858);
and U3504 (N_3504,N_2450,N_2087);
xor U3505 (N_3505,N_2326,N_1763);
nand U3506 (N_3506,N_2335,N_2158);
xor U3507 (N_3507,N_2201,N_2860);
or U3508 (N_3508,N_2363,N_1874);
nand U3509 (N_3509,N_2272,N_2750);
xnor U3510 (N_3510,N_2794,N_1899);
and U3511 (N_3511,N_1947,N_2589);
nand U3512 (N_3512,N_2172,N_2412);
or U3513 (N_3513,N_2483,N_2587);
and U3514 (N_3514,N_1953,N_1751);
nand U3515 (N_3515,N_2776,N_2984);
nor U3516 (N_3516,N_1641,N_1925);
or U3517 (N_3517,N_1741,N_2864);
xor U3518 (N_3518,N_1883,N_2317);
nor U3519 (N_3519,N_2298,N_2542);
and U3520 (N_3520,N_2783,N_2597);
nor U3521 (N_3521,N_1872,N_2402);
nand U3522 (N_3522,N_2428,N_1702);
nand U3523 (N_3523,N_2448,N_2210);
nor U3524 (N_3524,N_2909,N_2976);
xnor U3525 (N_3525,N_1760,N_2085);
and U3526 (N_3526,N_2076,N_2570);
nand U3527 (N_3527,N_2485,N_1675);
or U3528 (N_3528,N_2373,N_2921);
or U3529 (N_3529,N_2550,N_1694);
xor U3530 (N_3530,N_2559,N_2979);
xor U3531 (N_3531,N_2131,N_2284);
and U3532 (N_3532,N_1719,N_2577);
nand U3533 (N_3533,N_2169,N_2839);
and U3534 (N_3534,N_1813,N_1964);
or U3535 (N_3535,N_1980,N_1506);
nor U3536 (N_3536,N_2651,N_1836);
nor U3537 (N_3537,N_2668,N_2742);
xor U3538 (N_3538,N_1840,N_1765);
and U3539 (N_3539,N_2017,N_2337);
xor U3540 (N_3540,N_2081,N_1716);
and U3541 (N_3541,N_2785,N_1687);
xnor U3542 (N_3542,N_2912,N_2784);
nor U3543 (N_3543,N_2377,N_2530);
xnor U3544 (N_3544,N_2125,N_2702);
xor U3545 (N_3545,N_2038,N_2569);
xor U3546 (N_3546,N_2951,N_2580);
nand U3547 (N_3547,N_2857,N_2538);
nand U3548 (N_3548,N_2055,N_2029);
or U3549 (N_3549,N_1537,N_2147);
or U3550 (N_3550,N_1645,N_2899);
or U3551 (N_3551,N_2214,N_2639);
xnor U3552 (N_3552,N_1643,N_2652);
nand U3553 (N_3553,N_2836,N_2212);
xnor U3554 (N_3554,N_2881,N_1908);
xnor U3555 (N_3555,N_2928,N_1549);
and U3556 (N_3556,N_2808,N_2333);
nor U3557 (N_3557,N_1514,N_2683);
xor U3558 (N_3558,N_2520,N_2756);
xnor U3559 (N_3559,N_1530,N_2504);
and U3560 (N_3560,N_2070,N_2409);
nand U3561 (N_3561,N_2199,N_2661);
nand U3562 (N_3562,N_2527,N_2646);
nand U3563 (N_3563,N_2820,N_2463);
xor U3564 (N_3564,N_2341,N_2067);
nand U3565 (N_3565,N_2320,N_2229);
or U3566 (N_3566,N_1608,N_1782);
nor U3567 (N_3567,N_1648,N_1795);
xnor U3568 (N_3568,N_1810,N_2431);
and U3569 (N_3569,N_1627,N_2592);
or U3570 (N_3570,N_1733,N_2195);
nand U3571 (N_3571,N_2391,N_2183);
or U3572 (N_3572,N_2945,N_2008);
or U3573 (N_3573,N_2124,N_2680);
nor U3574 (N_3574,N_1550,N_2834);
or U3575 (N_3575,N_2636,N_1922);
nand U3576 (N_3576,N_1959,N_2893);
nor U3577 (N_3577,N_2230,N_1906);
and U3578 (N_3578,N_2160,N_1557);
xor U3579 (N_3579,N_2436,N_2686);
and U3580 (N_3580,N_1957,N_1517);
nor U3581 (N_3581,N_1892,N_1842);
nand U3582 (N_3582,N_2182,N_2238);
xor U3583 (N_3583,N_2497,N_1932);
and U3584 (N_3584,N_2389,N_1775);
xnor U3585 (N_3585,N_2344,N_1988);
nor U3586 (N_3586,N_2855,N_1700);
xor U3587 (N_3587,N_2490,N_2858);
nor U3588 (N_3588,N_2387,N_2659);
and U3589 (N_3589,N_2174,N_1618);
and U3590 (N_3590,N_1614,N_2792);
xnor U3591 (N_3591,N_1912,N_1696);
or U3592 (N_3592,N_1684,N_2699);
xnor U3593 (N_3593,N_2562,N_2456);
and U3594 (N_3594,N_1779,N_2778);
or U3595 (N_3595,N_2128,N_2561);
nand U3596 (N_3596,N_2033,N_2752);
and U3597 (N_3597,N_2166,N_1903);
xnor U3598 (N_3598,N_2519,N_2173);
and U3599 (N_3599,N_2461,N_1673);
and U3600 (N_3600,N_2848,N_2956);
or U3601 (N_3601,N_1827,N_1837);
nor U3602 (N_3602,N_2115,N_2099);
and U3603 (N_3603,N_1712,N_1859);
nand U3604 (N_3604,N_2967,N_2137);
nor U3605 (N_3605,N_2918,N_2140);
and U3606 (N_3606,N_1721,N_2969);
xor U3607 (N_3607,N_1770,N_2722);
xnor U3608 (N_3608,N_1672,N_2108);
nor U3609 (N_3609,N_2193,N_2063);
nand U3610 (N_3610,N_2935,N_2825);
and U3611 (N_3611,N_2007,N_2875);
nand U3612 (N_3612,N_1535,N_1559);
nand U3613 (N_3613,N_2142,N_2689);
and U3614 (N_3614,N_2354,N_2932);
or U3615 (N_3615,N_2495,N_1876);
nor U3616 (N_3616,N_2430,N_1894);
nand U3617 (N_3617,N_2833,N_1523);
and U3618 (N_3618,N_1946,N_2937);
nand U3619 (N_3619,N_2096,N_1819);
xor U3620 (N_3620,N_1551,N_2365);
or U3621 (N_3621,N_2025,N_1708);
or U3622 (N_3622,N_2459,N_1610);
or U3623 (N_3623,N_2327,N_2840);
nor U3624 (N_3624,N_1975,N_2143);
or U3625 (N_3625,N_2764,N_2695);
or U3626 (N_3626,N_1569,N_2814);
nor U3627 (N_3627,N_1647,N_2931);
nand U3628 (N_3628,N_2419,N_2120);
or U3629 (N_3629,N_2988,N_1984);
and U3630 (N_3630,N_1646,N_1701);
or U3631 (N_3631,N_2488,N_2152);
and U3632 (N_3632,N_2064,N_1564);
xor U3633 (N_3633,N_1725,N_1933);
and U3634 (N_3634,N_1660,N_2627);
nand U3635 (N_3635,N_2112,N_1847);
nor U3636 (N_3636,N_2987,N_1680);
nor U3637 (N_3637,N_2486,N_2896);
or U3638 (N_3638,N_2296,N_1952);
or U3639 (N_3639,N_2557,N_2575);
nand U3640 (N_3640,N_2312,N_2016);
nor U3641 (N_3641,N_2443,N_1629);
xor U3642 (N_3642,N_1777,N_2558);
nor U3643 (N_3643,N_1875,N_1548);
nand U3644 (N_3644,N_2252,N_2633);
or U3645 (N_3645,N_1690,N_1824);
xnor U3646 (N_3646,N_1590,N_2762);
nor U3647 (N_3647,N_2478,N_1867);
nor U3648 (N_3648,N_1664,N_2084);
nand U3649 (N_3649,N_1742,N_2281);
nand U3650 (N_3650,N_2258,N_2755);
or U3651 (N_3651,N_2779,N_1574);
or U3652 (N_3652,N_2511,N_1621);
xor U3653 (N_3653,N_2867,N_1918);
nand U3654 (N_3654,N_2614,N_2300);
and U3655 (N_3655,N_2554,N_2876);
nand U3656 (N_3656,N_2656,N_1969);
and U3657 (N_3657,N_2130,N_2075);
nor U3658 (N_3658,N_2793,N_1806);
or U3659 (N_3659,N_2294,N_2054);
nor U3660 (N_3660,N_2859,N_2963);
and U3661 (N_3661,N_2930,N_2594);
xnor U3662 (N_3662,N_2455,N_1800);
nor U3663 (N_3663,N_2209,N_2983);
and U3664 (N_3664,N_1605,N_2197);
or U3665 (N_3665,N_2400,N_1707);
or U3666 (N_3666,N_1998,N_2348);
nand U3667 (N_3667,N_2353,N_2878);
nand U3668 (N_3668,N_1845,N_2824);
nand U3669 (N_3669,N_2891,N_1597);
nand U3670 (N_3670,N_2421,N_1893);
nand U3671 (N_3671,N_2154,N_2737);
or U3672 (N_3672,N_2424,N_2816);
xor U3673 (N_3673,N_1653,N_1709);
nor U3674 (N_3674,N_1679,N_1854);
or U3675 (N_3675,N_2290,N_2753);
xor U3676 (N_3676,N_2516,N_2477);
xor U3677 (N_3677,N_1831,N_2513);
nand U3678 (N_3678,N_2703,N_2556);
and U3679 (N_3679,N_2192,N_2396);
xnor U3680 (N_3680,N_2060,N_2233);
nor U3681 (N_3681,N_1871,N_2224);
xnor U3682 (N_3682,N_1967,N_1650);
or U3683 (N_3683,N_2679,N_2213);
or U3684 (N_3684,N_2218,N_2690);
nor U3685 (N_3685,N_2217,N_2741);
nand U3686 (N_3686,N_1689,N_2040);
or U3687 (N_3687,N_1570,N_2631);
xor U3688 (N_3688,N_2943,N_2628);
nor U3689 (N_3689,N_1856,N_1625);
nand U3690 (N_3690,N_2671,N_2035);
xnor U3691 (N_3691,N_1635,N_2767);
xnor U3692 (N_3692,N_2080,N_1678);
nand U3693 (N_3693,N_1915,N_2994);
or U3694 (N_3694,N_2769,N_2196);
or U3695 (N_3695,N_2139,N_1901);
xnor U3696 (N_3696,N_1781,N_2844);
nor U3697 (N_3697,N_2797,N_1826);
nor U3698 (N_3698,N_2011,N_1568);
or U3699 (N_3699,N_2971,N_2078);
and U3700 (N_3700,N_1869,N_1656);
or U3701 (N_3701,N_2234,N_1866);
nand U3702 (N_3702,N_2748,N_1753);
xnor U3703 (N_3703,N_2228,N_2111);
nand U3704 (N_3704,N_2905,N_1944);
xnor U3705 (N_3705,N_2581,N_2827);
and U3706 (N_3706,N_2847,N_1536);
nand U3707 (N_3707,N_2521,N_1759);
or U3708 (N_3708,N_1904,N_1659);
nand U3709 (N_3709,N_2749,N_1993);
nor U3710 (N_3710,N_2082,N_1728);
nor U3711 (N_3711,N_1644,N_2990);
xor U3712 (N_3712,N_2367,N_2726);
nand U3713 (N_3713,N_1636,N_1821);
and U3714 (N_3714,N_2674,N_2004);
nand U3715 (N_3715,N_1595,N_2434);
and U3716 (N_3716,N_1505,N_2175);
xnor U3717 (N_3717,N_1951,N_1971);
or U3718 (N_3718,N_1936,N_2372);
or U3719 (N_3719,N_2014,N_2226);
and U3720 (N_3720,N_2123,N_2432);
and U3721 (N_3721,N_2841,N_2812);
xnor U3722 (N_3722,N_2145,N_2198);
nand U3723 (N_3723,N_2242,N_2629);
and U3724 (N_3724,N_2024,N_2052);
and U3725 (N_3725,N_2288,N_2739);
nand U3726 (N_3726,N_1945,N_2280);
nor U3727 (N_3727,N_2539,N_1939);
or U3728 (N_3728,N_2309,N_2092);
nand U3729 (N_3729,N_1591,N_1830);
nor U3730 (N_3730,N_2021,N_1534);
nand U3731 (N_3731,N_1766,N_2292);
nand U3732 (N_3732,N_1501,N_2018);
nand U3733 (N_3733,N_1676,N_2072);
xor U3734 (N_3734,N_1755,N_2725);
and U3735 (N_3735,N_1634,N_2093);
or U3736 (N_3736,N_2262,N_2992);
xor U3737 (N_3737,N_2264,N_2917);
and U3738 (N_3738,N_1767,N_2610);
xor U3739 (N_3739,N_1820,N_1818);
nor U3740 (N_3740,N_2845,N_2717);
and U3741 (N_3741,N_1560,N_2439);
xnor U3742 (N_3742,N_2673,N_2772);
nor U3743 (N_3743,N_2760,N_2873);
nand U3744 (N_3744,N_2500,N_1512);
nand U3745 (N_3745,N_2729,N_2526);
nand U3746 (N_3746,N_1571,N_2408);
or U3747 (N_3747,N_2458,N_1761);
nor U3748 (N_3748,N_2219,N_2221);
nor U3749 (N_3749,N_2136,N_2357);
xnor U3750 (N_3750,N_1844,N_1640);
xnor U3751 (N_3751,N_2485,N_2407);
xor U3752 (N_3752,N_2095,N_2428);
xor U3753 (N_3753,N_2122,N_1897);
nor U3754 (N_3754,N_1581,N_2706);
or U3755 (N_3755,N_2757,N_1774);
or U3756 (N_3756,N_2688,N_2345);
and U3757 (N_3757,N_2333,N_2879);
and U3758 (N_3758,N_2340,N_2625);
or U3759 (N_3759,N_2836,N_2811);
xnor U3760 (N_3760,N_1772,N_1906);
nand U3761 (N_3761,N_2443,N_2839);
and U3762 (N_3762,N_1914,N_2241);
nor U3763 (N_3763,N_2202,N_2041);
nand U3764 (N_3764,N_2455,N_1890);
xnor U3765 (N_3765,N_1898,N_2826);
or U3766 (N_3766,N_1579,N_1565);
xor U3767 (N_3767,N_2042,N_2710);
or U3768 (N_3768,N_2226,N_2654);
nand U3769 (N_3769,N_2541,N_1934);
xor U3770 (N_3770,N_2566,N_1958);
nor U3771 (N_3771,N_2646,N_2815);
and U3772 (N_3772,N_2492,N_2971);
nor U3773 (N_3773,N_2160,N_1799);
xor U3774 (N_3774,N_2453,N_2492);
nor U3775 (N_3775,N_2674,N_2375);
nor U3776 (N_3776,N_2654,N_1981);
nand U3777 (N_3777,N_1970,N_2675);
xnor U3778 (N_3778,N_2800,N_2085);
xnor U3779 (N_3779,N_2234,N_2513);
and U3780 (N_3780,N_2374,N_2533);
nor U3781 (N_3781,N_2592,N_1611);
and U3782 (N_3782,N_2466,N_2060);
and U3783 (N_3783,N_2563,N_2493);
or U3784 (N_3784,N_1562,N_1505);
or U3785 (N_3785,N_2818,N_2078);
and U3786 (N_3786,N_1547,N_2469);
nand U3787 (N_3787,N_1840,N_2394);
and U3788 (N_3788,N_2124,N_1816);
and U3789 (N_3789,N_2163,N_1807);
nor U3790 (N_3790,N_1871,N_1835);
xor U3791 (N_3791,N_2798,N_2431);
and U3792 (N_3792,N_2272,N_1921);
xor U3793 (N_3793,N_2220,N_2291);
or U3794 (N_3794,N_2474,N_1623);
and U3795 (N_3795,N_1797,N_2048);
nand U3796 (N_3796,N_2970,N_2741);
nor U3797 (N_3797,N_2084,N_2113);
nand U3798 (N_3798,N_2512,N_1530);
nor U3799 (N_3799,N_2796,N_2062);
xnor U3800 (N_3800,N_2892,N_1889);
nor U3801 (N_3801,N_1835,N_2582);
xor U3802 (N_3802,N_2343,N_2965);
nand U3803 (N_3803,N_2486,N_2348);
or U3804 (N_3804,N_2456,N_2264);
xor U3805 (N_3805,N_2224,N_2209);
and U3806 (N_3806,N_1788,N_1915);
or U3807 (N_3807,N_1539,N_1752);
xnor U3808 (N_3808,N_2469,N_2692);
or U3809 (N_3809,N_1570,N_2603);
or U3810 (N_3810,N_2156,N_2410);
or U3811 (N_3811,N_1729,N_1562);
or U3812 (N_3812,N_1871,N_1509);
nor U3813 (N_3813,N_2127,N_1918);
nor U3814 (N_3814,N_1802,N_2822);
nand U3815 (N_3815,N_1910,N_2585);
xnor U3816 (N_3816,N_2262,N_1737);
or U3817 (N_3817,N_2446,N_2572);
xor U3818 (N_3818,N_2531,N_1617);
and U3819 (N_3819,N_2893,N_1733);
or U3820 (N_3820,N_2217,N_2278);
or U3821 (N_3821,N_2112,N_2581);
and U3822 (N_3822,N_2830,N_2276);
nand U3823 (N_3823,N_2738,N_2435);
or U3824 (N_3824,N_2045,N_2787);
or U3825 (N_3825,N_2298,N_1643);
nor U3826 (N_3826,N_2676,N_1642);
nor U3827 (N_3827,N_2916,N_1712);
and U3828 (N_3828,N_2652,N_1663);
or U3829 (N_3829,N_2822,N_1987);
nand U3830 (N_3830,N_2513,N_1745);
and U3831 (N_3831,N_1776,N_1553);
xnor U3832 (N_3832,N_1761,N_2945);
or U3833 (N_3833,N_1913,N_1714);
nand U3834 (N_3834,N_2833,N_2143);
xor U3835 (N_3835,N_2690,N_1991);
xor U3836 (N_3836,N_1799,N_2719);
and U3837 (N_3837,N_2907,N_2043);
xor U3838 (N_3838,N_2333,N_1680);
nand U3839 (N_3839,N_2636,N_2589);
xnor U3840 (N_3840,N_2153,N_2916);
nor U3841 (N_3841,N_2724,N_2927);
nand U3842 (N_3842,N_1552,N_2750);
nand U3843 (N_3843,N_2444,N_1672);
or U3844 (N_3844,N_2916,N_2945);
or U3845 (N_3845,N_2160,N_1693);
nor U3846 (N_3846,N_1666,N_2060);
nand U3847 (N_3847,N_2484,N_1504);
nor U3848 (N_3848,N_1657,N_2899);
nor U3849 (N_3849,N_1866,N_2689);
xnor U3850 (N_3850,N_1639,N_2719);
xor U3851 (N_3851,N_1696,N_2571);
nand U3852 (N_3852,N_1870,N_2129);
nand U3853 (N_3853,N_2919,N_2842);
nor U3854 (N_3854,N_1738,N_2497);
and U3855 (N_3855,N_2623,N_1751);
xnor U3856 (N_3856,N_2587,N_1798);
and U3857 (N_3857,N_1852,N_1658);
xor U3858 (N_3858,N_2049,N_2456);
nor U3859 (N_3859,N_2272,N_2139);
nor U3860 (N_3860,N_2337,N_2231);
xor U3861 (N_3861,N_1828,N_2055);
xnor U3862 (N_3862,N_2654,N_2051);
and U3863 (N_3863,N_2762,N_2920);
xnor U3864 (N_3864,N_2975,N_2752);
nor U3865 (N_3865,N_2028,N_2942);
or U3866 (N_3866,N_1668,N_1509);
nand U3867 (N_3867,N_1506,N_2932);
nor U3868 (N_3868,N_2948,N_2356);
or U3869 (N_3869,N_2108,N_2779);
xor U3870 (N_3870,N_2940,N_1570);
nand U3871 (N_3871,N_2559,N_1631);
and U3872 (N_3872,N_2610,N_1950);
or U3873 (N_3873,N_1860,N_2529);
and U3874 (N_3874,N_2650,N_1559);
nor U3875 (N_3875,N_2587,N_1665);
and U3876 (N_3876,N_1587,N_2980);
and U3877 (N_3877,N_1620,N_2572);
xnor U3878 (N_3878,N_2865,N_2575);
or U3879 (N_3879,N_2673,N_1895);
nor U3880 (N_3880,N_1969,N_1668);
nor U3881 (N_3881,N_2011,N_2719);
nand U3882 (N_3882,N_2579,N_2071);
or U3883 (N_3883,N_2911,N_2460);
xor U3884 (N_3884,N_2014,N_2887);
nand U3885 (N_3885,N_2458,N_1806);
and U3886 (N_3886,N_2137,N_2266);
xnor U3887 (N_3887,N_2961,N_2424);
and U3888 (N_3888,N_2756,N_1888);
and U3889 (N_3889,N_2509,N_2120);
nor U3890 (N_3890,N_1641,N_2343);
or U3891 (N_3891,N_2763,N_2296);
nand U3892 (N_3892,N_1897,N_2909);
nor U3893 (N_3893,N_1885,N_2771);
xnor U3894 (N_3894,N_2333,N_1601);
nor U3895 (N_3895,N_1621,N_1665);
nor U3896 (N_3896,N_1667,N_2287);
or U3897 (N_3897,N_1604,N_1774);
nor U3898 (N_3898,N_2785,N_2839);
or U3899 (N_3899,N_1685,N_2030);
or U3900 (N_3900,N_2423,N_2254);
or U3901 (N_3901,N_1650,N_2737);
or U3902 (N_3902,N_2250,N_1603);
nand U3903 (N_3903,N_2651,N_2342);
nand U3904 (N_3904,N_1876,N_1506);
nand U3905 (N_3905,N_2897,N_2426);
and U3906 (N_3906,N_2508,N_2315);
or U3907 (N_3907,N_2425,N_2638);
nand U3908 (N_3908,N_2715,N_2004);
nand U3909 (N_3909,N_1547,N_2972);
nor U3910 (N_3910,N_1675,N_1857);
nand U3911 (N_3911,N_2858,N_1741);
xnor U3912 (N_3912,N_1937,N_2578);
xnor U3913 (N_3913,N_2802,N_2559);
nor U3914 (N_3914,N_1918,N_2648);
xnor U3915 (N_3915,N_2575,N_2648);
and U3916 (N_3916,N_2839,N_2441);
xnor U3917 (N_3917,N_2605,N_1988);
and U3918 (N_3918,N_1961,N_1649);
nand U3919 (N_3919,N_1551,N_2878);
xor U3920 (N_3920,N_2037,N_1574);
nand U3921 (N_3921,N_2267,N_1639);
or U3922 (N_3922,N_1924,N_2831);
xnor U3923 (N_3923,N_2801,N_1719);
or U3924 (N_3924,N_2032,N_1545);
and U3925 (N_3925,N_2747,N_1660);
or U3926 (N_3926,N_2046,N_1637);
or U3927 (N_3927,N_2892,N_2910);
xor U3928 (N_3928,N_2696,N_2120);
and U3929 (N_3929,N_2400,N_2896);
xor U3930 (N_3930,N_2264,N_2191);
xnor U3931 (N_3931,N_2877,N_2816);
xnor U3932 (N_3932,N_2840,N_2567);
and U3933 (N_3933,N_2560,N_1844);
and U3934 (N_3934,N_2188,N_1702);
nand U3935 (N_3935,N_2951,N_1662);
and U3936 (N_3936,N_1614,N_1527);
xor U3937 (N_3937,N_2428,N_1987);
and U3938 (N_3938,N_1527,N_2233);
nor U3939 (N_3939,N_1688,N_2634);
or U3940 (N_3940,N_2599,N_1853);
xnor U3941 (N_3941,N_2683,N_1824);
nand U3942 (N_3942,N_2569,N_1799);
xor U3943 (N_3943,N_1595,N_2543);
nand U3944 (N_3944,N_2925,N_2710);
nand U3945 (N_3945,N_2289,N_2665);
nand U3946 (N_3946,N_1622,N_2201);
nand U3947 (N_3947,N_1831,N_2160);
or U3948 (N_3948,N_2005,N_2159);
or U3949 (N_3949,N_2698,N_2789);
nor U3950 (N_3950,N_2033,N_1614);
nand U3951 (N_3951,N_2032,N_2835);
nor U3952 (N_3952,N_2254,N_2690);
or U3953 (N_3953,N_1864,N_2685);
and U3954 (N_3954,N_1904,N_1789);
and U3955 (N_3955,N_1500,N_2376);
nand U3956 (N_3956,N_2746,N_2246);
and U3957 (N_3957,N_2432,N_1600);
nor U3958 (N_3958,N_2518,N_2191);
and U3959 (N_3959,N_2246,N_2025);
nor U3960 (N_3960,N_2305,N_2769);
nand U3961 (N_3961,N_2292,N_2674);
nand U3962 (N_3962,N_1649,N_2864);
nor U3963 (N_3963,N_2254,N_2511);
xnor U3964 (N_3964,N_1954,N_1760);
xor U3965 (N_3965,N_2974,N_2349);
nor U3966 (N_3966,N_1645,N_1872);
xor U3967 (N_3967,N_1740,N_2304);
xor U3968 (N_3968,N_1537,N_2560);
or U3969 (N_3969,N_2326,N_2588);
nor U3970 (N_3970,N_1820,N_2822);
nor U3971 (N_3971,N_2216,N_1933);
and U3972 (N_3972,N_2300,N_1581);
nor U3973 (N_3973,N_2059,N_2649);
nor U3974 (N_3974,N_2004,N_2910);
and U3975 (N_3975,N_2744,N_2713);
nand U3976 (N_3976,N_2197,N_1655);
nand U3977 (N_3977,N_2648,N_2291);
nor U3978 (N_3978,N_2519,N_2020);
xnor U3979 (N_3979,N_2579,N_1716);
and U3980 (N_3980,N_1876,N_2836);
or U3981 (N_3981,N_2636,N_2702);
xnor U3982 (N_3982,N_2227,N_2417);
nor U3983 (N_3983,N_1508,N_2162);
xor U3984 (N_3984,N_2360,N_2362);
and U3985 (N_3985,N_2468,N_2783);
and U3986 (N_3986,N_2560,N_2543);
nor U3987 (N_3987,N_2857,N_1704);
or U3988 (N_3988,N_1854,N_1644);
nor U3989 (N_3989,N_2679,N_2403);
nor U3990 (N_3990,N_2888,N_2741);
nor U3991 (N_3991,N_2505,N_1829);
nand U3992 (N_3992,N_2892,N_2602);
nand U3993 (N_3993,N_2431,N_2680);
nand U3994 (N_3994,N_1567,N_2272);
and U3995 (N_3995,N_1507,N_2639);
nand U3996 (N_3996,N_1711,N_1691);
and U3997 (N_3997,N_1589,N_1794);
xor U3998 (N_3998,N_1829,N_2500);
and U3999 (N_3999,N_2062,N_1863);
nand U4000 (N_4000,N_2968,N_2629);
nor U4001 (N_4001,N_2559,N_1994);
and U4002 (N_4002,N_2491,N_2773);
xor U4003 (N_4003,N_2830,N_2807);
nand U4004 (N_4004,N_2196,N_1526);
nand U4005 (N_4005,N_1607,N_2953);
nor U4006 (N_4006,N_2387,N_2185);
or U4007 (N_4007,N_1914,N_2117);
nor U4008 (N_4008,N_2188,N_2933);
or U4009 (N_4009,N_2809,N_1975);
and U4010 (N_4010,N_1539,N_1796);
nand U4011 (N_4011,N_1863,N_1910);
and U4012 (N_4012,N_2805,N_2133);
nand U4013 (N_4013,N_2468,N_2859);
and U4014 (N_4014,N_1816,N_1620);
xor U4015 (N_4015,N_1675,N_2204);
nand U4016 (N_4016,N_1671,N_2587);
and U4017 (N_4017,N_2638,N_1573);
or U4018 (N_4018,N_2810,N_2393);
nor U4019 (N_4019,N_2675,N_2522);
nand U4020 (N_4020,N_2564,N_2391);
and U4021 (N_4021,N_2031,N_2421);
and U4022 (N_4022,N_2961,N_2708);
nor U4023 (N_4023,N_2668,N_1867);
nor U4024 (N_4024,N_2173,N_2405);
or U4025 (N_4025,N_1976,N_2218);
nand U4026 (N_4026,N_2930,N_1921);
and U4027 (N_4027,N_1934,N_2416);
nand U4028 (N_4028,N_2043,N_1672);
nor U4029 (N_4029,N_2312,N_1580);
and U4030 (N_4030,N_2607,N_2310);
nand U4031 (N_4031,N_2232,N_2343);
nor U4032 (N_4032,N_2171,N_1895);
and U4033 (N_4033,N_2901,N_1558);
xor U4034 (N_4034,N_2088,N_1624);
nor U4035 (N_4035,N_1631,N_2168);
nor U4036 (N_4036,N_2140,N_2761);
xor U4037 (N_4037,N_2829,N_2805);
xnor U4038 (N_4038,N_2900,N_2541);
nor U4039 (N_4039,N_2827,N_2719);
and U4040 (N_4040,N_2038,N_2156);
nand U4041 (N_4041,N_1871,N_2255);
xnor U4042 (N_4042,N_2411,N_1682);
nor U4043 (N_4043,N_2352,N_2788);
nand U4044 (N_4044,N_1773,N_1822);
and U4045 (N_4045,N_2230,N_1569);
nor U4046 (N_4046,N_1792,N_1533);
or U4047 (N_4047,N_1526,N_1708);
xnor U4048 (N_4048,N_2595,N_2437);
nand U4049 (N_4049,N_1898,N_2510);
nor U4050 (N_4050,N_1621,N_2664);
or U4051 (N_4051,N_2435,N_1641);
xor U4052 (N_4052,N_2435,N_2767);
xnor U4053 (N_4053,N_2261,N_1828);
nor U4054 (N_4054,N_2664,N_1508);
nor U4055 (N_4055,N_1861,N_1955);
nor U4056 (N_4056,N_2654,N_2777);
nor U4057 (N_4057,N_2502,N_2770);
nand U4058 (N_4058,N_2672,N_1538);
nor U4059 (N_4059,N_2621,N_2372);
nand U4060 (N_4060,N_2323,N_1962);
nand U4061 (N_4061,N_2250,N_1629);
xnor U4062 (N_4062,N_1613,N_1678);
nor U4063 (N_4063,N_2386,N_1611);
nand U4064 (N_4064,N_1741,N_2165);
or U4065 (N_4065,N_2265,N_1812);
nor U4066 (N_4066,N_1990,N_2340);
and U4067 (N_4067,N_2912,N_1619);
or U4068 (N_4068,N_2826,N_2658);
and U4069 (N_4069,N_1592,N_1524);
nor U4070 (N_4070,N_2455,N_1701);
nor U4071 (N_4071,N_2524,N_1708);
xor U4072 (N_4072,N_2476,N_2045);
and U4073 (N_4073,N_2598,N_1703);
nand U4074 (N_4074,N_2321,N_2007);
nor U4075 (N_4075,N_1811,N_1804);
xnor U4076 (N_4076,N_2384,N_2149);
nor U4077 (N_4077,N_1569,N_1771);
or U4078 (N_4078,N_2210,N_2967);
xnor U4079 (N_4079,N_2673,N_2363);
nand U4080 (N_4080,N_2811,N_1676);
and U4081 (N_4081,N_2056,N_2620);
and U4082 (N_4082,N_2731,N_2522);
or U4083 (N_4083,N_2600,N_1627);
and U4084 (N_4084,N_2180,N_2357);
nand U4085 (N_4085,N_2427,N_1660);
xnor U4086 (N_4086,N_2786,N_2328);
xnor U4087 (N_4087,N_2970,N_2904);
xnor U4088 (N_4088,N_2527,N_2136);
or U4089 (N_4089,N_2147,N_1798);
nand U4090 (N_4090,N_2067,N_2256);
nand U4091 (N_4091,N_1644,N_2419);
nand U4092 (N_4092,N_2995,N_2037);
nand U4093 (N_4093,N_2078,N_1563);
and U4094 (N_4094,N_2880,N_2015);
xor U4095 (N_4095,N_2549,N_2675);
nand U4096 (N_4096,N_2289,N_1825);
nor U4097 (N_4097,N_2804,N_2313);
and U4098 (N_4098,N_2000,N_2153);
and U4099 (N_4099,N_2127,N_2421);
or U4100 (N_4100,N_2774,N_1543);
nand U4101 (N_4101,N_2788,N_2162);
xor U4102 (N_4102,N_2999,N_1800);
nor U4103 (N_4103,N_1537,N_2186);
or U4104 (N_4104,N_1695,N_2807);
nand U4105 (N_4105,N_2496,N_2512);
and U4106 (N_4106,N_2029,N_1910);
and U4107 (N_4107,N_1969,N_1783);
nand U4108 (N_4108,N_2160,N_1643);
xnor U4109 (N_4109,N_2145,N_2291);
nor U4110 (N_4110,N_2807,N_1680);
xnor U4111 (N_4111,N_1624,N_2921);
nand U4112 (N_4112,N_2645,N_2319);
xnor U4113 (N_4113,N_2210,N_1978);
or U4114 (N_4114,N_1573,N_1618);
xnor U4115 (N_4115,N_1909,N_1534);
or U4116 (N_4116,N_2847,N_2352);
nand U4117 (N_4117,N_1933,N_1795);
or U4118 (N_4118,N_1799,N_1788);
and U4119 (N_4119,N_1934,N_1699);
xor U4120 (N_4120,N_2707,N_1967);
nand U4121 (N_4121,N_2218,N_2239);
and U4122 (N_4122,N_2630,N_2854);
and U4123 (N_4123,N_1775,N_1861);
xnor U4124 (N_4124,N_2176,N_2593);
or U4125 (N_4125,N_1703,N_2625);
nand U4126 (N_4126,N_2871,N_2571);
and U4127 (N_4127,N_2007,N_2089);
xor U4128 (N_4128,N_2338,N_2289);
xor U4129 (N_4129,N_1751,N_2801);
nand U4130 (N_4130,N_2179,N_2890);
and U4131 (N_4131,N_2401,N_2306);
or U4132 (N_4132,N_2927,N_1502);
or U4133 (N_4133,N_1994,N_2807);
or U4134 (N_4134,N_1848,N_2611);
and U4135 (N_4135,N_2126,N_1683);
nand U4136 (N_4136,N_1868,N_2693);
xnor U4137 (N_4137,N_1880,N_2944);
xnor U4138 (N_4138,N_1932,N_1599);
and U4139 (N_4139,N_2982,N_1509);
and U4140 (N_4140,N_2458,N_2363);
nor U4141 (N_4141,N_2255,N_2610);
or U4142 (N_4142,N_2502,N_1530);
and U4143 (N_4143,N_2040,N_2054);
xor U4144 (N_4144,N_1813,N_1733);
or U4145 (N_4145,N_1763,N_2547);
nor U4146 (N_4146,N_1635,N_2942);
and U4147 (N_4147,N_2361,N_2102);
and U4148 (N_4148,N_2931,N_2488);
xor U4149 (N_4149,N_2845,N_2175);
xor U4150 (N_4150,N_2380,N_2801);
xor U4151 (N_4151,N_2274,N_2858);
xor U4152 (N_4152,N_2058,N_1793);
xnor U4153 (N_4153,N_2249,N_1662);
or U4154 (N_4154,N_2319,N_2627);
and U4155 (N_4155,N_1851,N_2226);
nand U4156 (N_4156,N_1772,N_1624);
and U4157 (N_4157,N_2711,N_1978);
xor U4158 (N_4158,N_2751,N_1726);
or U4159 (N_4159,N_2669,N_2912);
or U4160 (N_4160,N_1612,N_1896);
or U4161 (N_4161,N_2905,N_2306);
nand U4162 (N_4162,N_2984,N_2061);
or U4163 (N_4163,N_2107,N_1821);
and U4164 (N_4164,N_2328,N_1785);
nor U4165 (N_4165,N_1858,N_2076);
or U4166 (N_4166,N_2276,N_1988);
nand U4167 (N_4167,N_2181,N_1748);
xnor U4168 (N_4168,N_2205,N_2984);
and U4169 (N_4169,N_1759,N_1730);
or U4170 (N_4170,N_2766,N_1660);
and U4171 (N_4171,N_2037,N_2455);
or U4172 (N_4172,N_2865,N_2655);
nor U4173 (N_4173,N_2223,N_2721);
xor U4174 (N_4174,N_2489,N_2965);
or U4175 (N_4175,N_2833,N_1525);
nand U4176 (N_4176,N_2473,N_2915);
nand U4177 (N_4177,N_1837,N_1867);
or U4178 (N_4178,N_2632,N_2536);
or U4179 (N_4179,N_2502,N_2352);
and U4180 (N_4180,N_2626,N_2579);
or U4181 (N_4181,N_1691,N_2125);
nor U4182 (N_4182,N_2170,N_2946);
and U4183 (N_4183,N_1541,N_1628);
and U4184 (N_4184,N_2396,N_2185);
nor U4185 (N_4185,N_2716,N_2835);
xor U4186 (N_4186,N_2141,N_1565);
or U4187 (N_4187,N_2681,N_1669);
nand U4188 (N_4188,N_1820,N_1929);
nand U4189 (N_4189,N_2593,N_2616);
nor U4190 (N_4190,N_2797,N_2369);
nor U4191 (N_4191,N_1557,N_2448);
nand U4192 (N_4192,N_2313,N_2395);
nor U4193 (N_4193,N_2504,N_2144);
and U4194 (N_4194,N_2065,N_2962);
nor U4195 (N_4195,N_2768,N_2399);
and U4196 (N_4196,N_1897,N_2041);
or U4197 (N_4197,N_2154,N_2089);
xor U4198 (N_4198,N_2986,N_1839);
xnor U4199 (N_4199,N_2043,N_1547);
or U4200 (N_4200,N_2403,N_2261);
xnor U4201 (N_4201,N_2423,N_2790);
nand U4202 (N_4202,N_1550,N_2712);
or U4203 (N_4203,N_1597,N_2000);
and U4204 (N_4204,N_2471,N_1893);
or U4205 (N_4205,N_2560,N_1826);
or U4206 (N_4206,N_2087,N_2984);
nor U4207 (N_4207,N_2161,N_2396);
nor U4208 (N_4208,N_1986,N_2249);
nor U4209 (N_4209,N_2980,N_2591);
xnor U4210 (N_4210,N_1537,N_1807);
or U4211 (N_4211,N_2418,N_2240);
xor U4212 (N_4212,N_2007,N_1895);
xor U4213 (N_4213,N_2049,N_1778);
xor U4214 (N_4214,N_1704,N_2309);
nand U4215 (N_4215,N_1822,N_2395);
xor U4216 (N_4216,N_2382,N_1925);
nor U4217 (N_4217,N_2839,N_1696);
nand U4218 (N_4218,N_2300,N_2613);
xor U4219 (N_4219,N_2109,N_2019);
or U4220 (N_4220,N_2162,N_2603);
xor U4221 (N_4221,N_1639,N_2095);
nand U4222 (N_4222,N_2836,N_1860);
xor U4223 (N_4223,N_1825,N_2498);
nand U4224 (N_4224,N_2027,N_2381);
nor U4225 (N_4225,N_1633,N_2183);
nor U4226 (N_4226,N_2237,N_1757);
and U4227 (N_4227,N_2684,N_2526);
or U4228 (N_4228,N_1957,N_2692);
or U4229 (N_4229,N_2244,N_2304);
xnor U4230 (N_4230,N_2566,N_2003);
xor U4231 (N_4231,N_2275,N_1637);
and U4232 (N_4232,N_2112,N_1975);
xnor U4233 (N_4233,N_1968,N_2435);
xnor U4234 (N_4234,N_1536,N_2554);
and U4235 (N_4235,N_1678,N_2816);
nor U4236 (N_4236,N_2622,N_2262);
nor U4237 (N_4237,N_2758,N_2557);
xor U4238 (N_4238,N_1880,N_2548);
xor U4239 (N_4239,N_2842,N_2962);
nand U4240 (N_4240,N_2259,N_2562);
nand U4241 (N_4241,N_1529,N_2614);
xor U4242 (N_4242,N_2961,N_2569);
xnor U4243 (N_4243,N_2982,N_2251);
xor U4244 (N_4244,N_2721,N_2155);
or U4245 (N_4245,N_2902,N_2585);
xnor U4246 (N_4246,N_2664,N_2970);
and U4247 (N_4247,N_1911,N_1641);
nand U4248 (N_4248,N_1718,N_1922);
xnor U4249 (N_4249,N_2425,N_2959);
nor U4250 (N_4250,N_1794,N_2727);
xor U4251 (N_4251,N_2338,N_1934);
nor U4252 (N_4252,N_1521,N_1596);
nor U4253 (N_4253,N_1925,N_2005);
nor U4254 (N_4254,N_1607,N_1878);
and U4255 (N_4255,N_2118,N_1986);
nand U4256 (N_4256,N_2786,N_2818);
nand U4257 (N_4257,N_2295,N_2323);
nand U4258 (N_4258,N_1640,N_1874);
and U4259 (N_4259,N_2285,N_1706);
nand U4260 (N_4260,N_1576,N_1965);
and U4261 (N_4261,N_1823,N_1918);
nor U4262 (N_4262,N_2422,N_2393);
and U4263 (N_4263,N_2242,N_2776);
nor U4264 (N_4264,N_2872,N_1628);
nor U4265 (N_4265,N_1998,N_2130);
nor U4266 (N_4266,N_2942,N_2369);
xnor U4267 (N_4267,N_1870,N_1652);
nand U4268 (N_4268,N_1857,N_1906);
and U4269 (N_4269,N_2184,N_2802);
nor U4270 (N_4270,N_1997,N_1885);
and U4271 (N_4271,N_2485,N_1948);
nor U4272 (N_4272,N_2800,N_2921);
xor U4273 (N_4273,N_1626,N_2948);
or U4274 (N_4274,N_2423,N_1958);
nor U4275 (N_4275,N_1814,N_2846);
xor U4276 (N_4276,N_2940,N_1933);
nor U4277 (N_4277,N_2894,N_2670);
xor U4278 (N_4278,N_2948,N_2569);
xnor U4279 (N_4279,N_1742,N_1957);
and U4280 (N_4280,N_1676,N_2133);
or U4281 (N_4281,N_1717,N_2953);
nand U4282 (N_4282,N_1886,N_2095);
nand U4283 (N_4283,N_2678,N_2567);
or U4284 (N_4284,N_1890,N_2484);
nand U4285 (N_4285,N_2938,N_1944);
xor U4286 (N_4286,N_2099,N_2596);
or U4287 (N_4287,N_2387,N_2100);
nor U4288 (N_4288,N_1615,N_2646);
or U4289 (N_4289,N_2776,N_1744);
nor U4290 (N_4290,N_2417,N_1867);
or U4291 (N_4291,N_1895,N_1726);
xor U4292 (N_4292,N_2908,N_2393);
nand U4293 (N_4293,N_1656,N_2039);
nand U4294 (N_4294,N_2470,N_2247);
xnor U4295 (N_4295,N_2454,N_2406);
or U4296 (N_4296,N_2583,N_2595);
nand U4297 (N_4297,N_2626,N_1938);
or U4298 (N_4298,N_1796,N_2821);
or U4299 (N_4299,N_1546,N_2510);
or U4300 (N_4300,N_1643,N_1872);
nand U4301 (N_4301,N_1764,N_2045);
nand U4302 (N_4302,N_1797,N_2139);
nor U4303 (N_4303,N_1712,N_2806);
nand U4304 (N_4304,N_1982,N_2333);
nand U4305 (N_4305,N_2160,N_1991);
nand U4306 (N_4306,N_2395,N_2022);
nor U4307 (N_4307,N_2583,N_2015);
xnor U4308 (N_4308,N_2566,N_2285);
and U4309 (N_4309,N_2766,N_2676);
nand U4310 (N_4310,N_1646,N_1865);
xnor U4311 (N_4311,N_2050,N_1636);
nand U4312 (N_4312,N_1934,N_1612);
nor U4313 (N_4313,N_2260,N_1730);
and U4314 (N_4314,N_2666,N_2381);
nor U4315 (N_4315,N_1737,N_1960);
nand U4316 (N_4316,N_1879,N_2025);
xor U4317 (N_4317,N_2173,N_2421);
nor U4318 (N_4318,N_2113,N_1545);
or U4319 (N_4319,N_2061,N_2411);
or U4320 (N_4320,N_2406,N_2716);
or U4321 (N_4321,N_1588,N_1502);
and U4322 (N_4322,N_2274,N_1565);
nor U4323 (N_4323,N_1889,N_2650);
nand U4324 (N_4324,N_2461,N_2157);
xor U4325 (N_4325,N_1626,N_2363);
and U4326 (N_4326,N_2598,N_2953);
xor U4327 (N_4327,N_2009,N_2145);
xnor U4328 (N_4328,N_1912,N_2271);
or U4329 (N_4329,N_2819,N_1601);
nor U4330 (N_4330,N_2515,N_1651);
or U4331 (N_4331,N_2578,N_1941);
or U4332 (N_4332,N_2994,N_1932);
nand U4333 (N_4333,N_1727,N_2455);
or U4334 (N_4334,N_2806,N_2420);
nor U4335 (N_4335,N_2965,N_1688);
nand U4336 (N_4336,N_1619,N_2709);
and U4337 (N_4337,N_2554,N_1952);
or U4338 (N_4338,N_2416,N_2542);
or U4339 (N_4339,N_1512,N_1700);
and U4340 (N_4340,N_2446,N_2603);
and U4341 (N_4341,N_2281,N_2653);
and U4342 (N_4342,N_2602,N_1562);
xor U4343 (N_4343,N_2936,N_2471);
and U4344 (N_4344,N_2440,N_2670);
nor U4345 (N_4345,N_2240,N_1918);
and U4346 (N_4346,N_2847,N_1669);
and U4347 (N_4347,N_2406,N_2996);
nor U4348 (N_4348,N_2890,N_2138);
and U4349 (N_4349,N_2600,N_1945);
xnor U4350 (N_4350,N_2670,N_2404);
xor U4351 (N_4351,N_1942,N_1813);
and U4352 (N_4352,N_2500,N_2051);
or U4353 (N_4353,N_1977,N_2286);
or U4354 (N_4354,N_2596,N_2412);
xnor U4355 (N_4355,N_2858,N_2208);
nand U4356 (N_4356,N_2314,N_2442);
nor U4357 (N_4357,N_2776,N_2166);
nand U4358 (N_4358,N_2431,N_2183);
xor U4359 (N_4359,N_1607,N_2344);
and U4360 (N_4360,N_1897,N_2603);
and U4361 (N_4361,N_2138,N_1571);
or U4362 (N_4362,N_2061,N_2852);
nand U4363 (N_4363,N_1967,N_1933);
nor U4364 (N_4364,N_2888,N_1743);
nand U4365 (N_4365,N_2343,N_1786);
xor U4366 (N_4366,N_2917,N_2707);
or U4367 (N_4367,N_2589,N_1615);
or U4368 (N_4368,N_2869,N_1691);
xnor U4369 (N_4369,N_1745,N_1873);
or U4370 (N_4370,N_1745,N_2334);
and U4371 (N_4371,N_1844,N_2657);
or U4372 (N_4372,N_2650,N_2801);
and U4373 (N_4373,N_1787,N_2526);
and U4374 (N_4374,N_2335,N_2117);
xor U4375 (N_4375,N_2249,N_2060);
or U4376 (N_4376,N_1827,N_1869);
nor U4377 (N_4377,N_2863,N_1714);
or U4378 (N_4378,N_2891,N_2011);
nand U4379 (N_4379,N_2145,N_1562);
and U4380 (N_4380,N_2261,N_1798);
and U4381 (N_4381,N_2792,N_2536);
nand U4382 (N_4382,N_2696,N_2834);
or U4383 (N_4383,N_2978,N_1581);
and U4384 (N_4384,N_2720,N_1937);
and U4385 (N_4385,N_2014,N_2782);
and U4386 (N_4386,N_2097,N_1510);
nand U4387 (N_4387,N_2205,N_2412);
or U4388 (N_4388,N_2324,N_2411);
or U4389 (N_4389,N_2197,N_2138);
nor U4390 (N_4390,N_2691,N_1613);
and U4391 (N_4391,N_1937,N_2516);
and U4392 (N_4392,N_1753,N_2275);
nand U4393 (N_4393,N_2261,N_1884);
nand U4394 (N_4394,N_2126,N_1841);
or U4395 (N_4395,N_2243,N_2116);
nand U4396 (N_4396,N_2442,N_1652);
and U4397 (N_4397,N_1604,N_2229);
nor U4398 (N_4398,N_2806,N_2329);
xor U4399 (N_4399,N_1843,N_2411);
or U4400 (N_4400,N_1709,N_2225);
xnor U4401 (N_4401,N_2089,N_2655);
nor U4402 (N_4402,N_2861,N_1666);
xnor U4403 (N_4403,N_1532,N_2543);
or U4404 (N_4404,N_2996,N_2433);
nor U4405 (N_4405,N_1566,N_2422);
and U4406 (N_4406,N_2916,N_2180);
nand U4407 (N_4407,N_1850,N_2820);
nor U4408 (N_4408,N_1590,N_2757);
and U4409 (N_4409,N_2761,N_2362);
xnor U4410 (N_4410,N_2520,N_2817);
xnor U4411 (N_4411,N_2115,N_2634);
and U4412 (N_4412,N_2550,N_1926);
and U4413 (N_4413,N_1587,N_2247);
nor U4414 (N_4414,N_2857,N_2608);
nor U4415 (N_4415,N_2859,N_2825);
xnor U4416 (N_4416,N_1962,N_1640);
and U4417 (N_4417,N_1832,N_1585);
or U4418 (N_4418,N_2996,N_2904);
nand U4419 (N_4419,N_2014,N_2626);
and U4420 (N_4420,N_2976,N_1789);
xnor U4421 (N_4421,N_1949,N_1725);
and U4422 (N_4422,N_1929,N_2589);
and U4423 (N_4423,N_1659,N_2187);
and U4424 (N_4424,N_2124,N_1653);
nor U4425 (N_4425,N_2839,N_2377);
nand U4426 (N_4426,N_2925,N_2353);
xnor U4427 (N_4427,N_1550,N_1768);
nor U4428 (N_4428,N_1586,N_2603);
nand U4429 (N_4429,N_2642,N_2065);
or U4430 (N_4430,N_2214,N_2411);
xor U4431 (N_4431,N_2379,N_1709);
and U4432 (N_4432,N_2903,N_2049);
nor U4433 (N_4433,N_1559,N_2005);
xnor U4434 (N_4434,N_1878,N_2737);
or U4435 (N_4435,N_1511,N_1508);
nand U4436 (N_4436,N_2598,N_2443);
and U4437 (N_4437,N_1929,N_2834);
or U4438 (N_4438,N_2504,N_2807);
xnor U4439 (N_4439,N_1645,N_2936);
nor U4440 (N_4440,N_1991,N_2070);
and U4441 (N_4441,N_2881,N_1508);
or U4442 (N_4442,N_2796,N_1917);
nor U4443 (N_4443,N_2315,N_2584);
and U4444 (N_4444,N_2546,N_1936);
xnor U4445 (N_4445,N_2574,N_1507);
xor U4446 (N_4446,N_1970,N_2382);
nor U4447 (N_4447,N_2389,N_2858);
xor U4448 (N_4448,N_2492,N_1726);
nor U4449 (N_4449,N_2522,N_2743);
and U4450 (N_4450,N_2645,N_2616);
or U4451 (N_4451,N_2785,N_1612);
and U4452 (N_4452,N_2461,N_1687);
and U4453 (N_4453,N_2014,N_1829);
nand U4454 (N_4454,N_2358,N_2781);
nand U4455 (N_4455,N_2577,N_2526);
nand U4456 (N_4456,N_1635,N_1669);
xnor U4457 (N_4457,N_2557,N_2203);
and U4458 (N_4458,N_2205,N_2193);
or U4459 (N_4459,N_1520,N_1557);
xor U4460 (N_4460,N_2782,N_2468);
or U4461 (N_4461,N_2059,N_2832);
nor U4462 (N_4462,N_1531,N_2978);
xor U4463 (N_4463,N_2226,N_2656);
and U4464 (N_4464,N_2970,N_2351);
xor U4465 (N_4465,N_2605,N_2981);
nand U4466 (N_4466,N_2609,N_2458);
or U4467 (N_4467,N_1610,N_2883);
and U4468 (N_4468,N_2067,N_2392);
nand U4469 (N_4469,N_2780,N_1561);
nor U4470 (N_4470,N_1729,N_2285);
xnor U4471 (N_4471,N_2560,N_1584);
or U4472 (N_4472,N_2763,N_2669);
xnor U4473 (N_4473,N_1940,N_2293);
and U4474 (N_4474,N_1992,N_2218);
xnor U4475 (N_4475,N_2777,N_1599);
and U4476 (N_4476,N_1503,N_2164);
xnor U4477 (N_4477,N_2677,N_1874);
xor U4478 (N_4478,N_1582,N_2150);
and U4479 (N_4479,N_1591,N_2014);
or U4480 (N_4480,N_1511,N_2613);
xnor U4481 (N_4481,N_2365,N_1765);
and U4482 (N_4482,N_1654,N_2224);
nand U4483 (N_4483,N_2717,N_2223);
nor U4484 (N_4484,N_2510,N_1537);
nand U4485 (N_4485,N_2334,N_1807);
nand U4486 (N_4486,N_2432,N_2431);
xor U4487 (N_4487,N_2398,N_1797);
xnor U4488 (N_4488,N_2311,N_2104);
or U4489 (N_4489,N_2013,N_1611);
nand U4490 (N_4490,N_1867,N_2197);
nand U4491 (N_4491,N_1562,N_1784);
and U4492 (N_4492,N_2657,N_2580);
or U4493 (N_4493,N_2034,N_2630);
xnor U4494 (N_4494,N_2255,N_2017);
or U4495 (N_4495,N_2247,N_2577);
and U4496 (N_4496,N_2059,N_2672);
nor U4497 (N_4497,N_2997,N_2260);
and U4498 (N_4498,N_1855,N_2414);
nor U4499 (N_4499,N_1641,N_1518);
or U4500 (N_4500,N_4187,N_4147);
nand U4501 (N_4501,N_3769,N_3135);
xor U4502 (N_4502,N_3829,N_3931);
nor U4503 (N_4503,N_4458,N_4144);
or U4504 (N_4504,N_3059,N_3184);
xnor U4505 (N_4505,N_3662,N_3714);
or U4506 (N_4506,N_3876,N_3070);
xor U4507 (N_4507,N_3802,N_3837);
and U4508 (N_4508,N_3191,N_3905);
or U4509 (N_4509,N_3220,N_4275);
and U4510 (N_4510,N_3508,N_3491);
xnor U4511 (N_4511,N_4169,N_3160);
xnor U4512 (N_4512,N_3418,N_4017);
xnor U4513 (N_4513,N_3056,N_4194);
and U4514 (N_4514,N_3459,N_3154);
xor U4515 (N_4515,N_3292,N_3368);
nand U4516 (N_4516,N_4047,N_4013);
or U4517 (N_4517,N_3913,N_3590);
or U4518 (N_4518,N_4197,N_3315);
nand U4519 (N_4519,N_3926,N_4201);
or U4520 (N_4520,N_3511,N_3826);
or U4521 (N_4521,N_3100,N_4494);
nand U4522 (N_4522,N_3020,N_4385);
nor U4523 (N_4523,N_3378,N_3237);
nor U4524 (N_4524,N_3813,N_3375);
nor U4525 (N_4525,N_3647,N_3705);
or U4526 (N_4526,N_4460,N_3830);
xor U4527 (N_4527,N_3514,N_4315);
or U4528 (N_4528,N_3642,N_3503);
or U4529 (N_4529,N_4272,N_4174);
nor U4530 (N_4530,N_4291,N_3602);
xnor U4531 (N_4531,N_3666,N_3189);
nor U4532 (N_4532,N_3290,N_4283);
nand U4533 (N_4533,N_4210,N_4447);
nor U4534 (N_4534,N_3472,N_3080);
nand U4535 (N_4535,N_3961,N_3079);
nor U4536 (N_4536,N_3981,N_4044);
nand U4537 (N_4537,N_3965,N_4414);
nor U4538 (N_4538,N_4025,N_3153);
nand U4539 (N_4539,N_4455,N_3739);
nor U4540 (N_4540,N_3137,N_4337);
and U4541 (N_4541,N_3027,N_3575);
nor U4542 (N_4542,N_3879,N_4005);
nor U4543 (N_4543,N_3466,N_4206);
and U4544 (N_4544,N_3619,N_3943);
nand U4545 (N_4545,N_3078,N_3163);
nor U4546 (N_4546,N_4152,N_3749);
nor U4547 (N_4547,N_3777,N_4485);
and U4548 (N_4548,N_3525,N_3316);
and U4549 (N_4549,N_3329,N_3134);
or U4550 (N_4550,N_3695,N_3013);
nand U4551 (N_4551,N_3517,N_3430);
nand U4552 (N_4552,N_3039,N_4293);
xnor U4553 (N_4553,N_3624,N_4319);
nand U4554 (N_4554,N_3089,N_3608);
nor U4555 (N_4555,N_3268,N_4223);
nor U4556 (N_4556,N_4222,N_4259);
xnor U4557 (N_4557,N_3337,N_3344);
or U4558 (N_4558,N_4381,N_3932);
or U4559 (N_4559,N_4074,N_3435);
and U4560 (N_4560,N_3983,N_3615);
and U4561 (N_4561,N_4063,N_4393);
nor U4562 (N_4562,N_3485,N_3627);
or U4563 (N_4563,N_4247,N_4466);
or U4564 (N_4564,N_3878,N_3622);
xnor U4565 (N_4565,N_3032,N_3018);
nor U4566 (N_4566,N_4190,N_4449);
or U4567 (N_4567,N_4023,N_4036);
or U4568 (N_4568,N_4295,N_3437);
and U4569 (N_4569,N_4229,N_3850);
nand U4570 (N_4570,N_3420,N_3677);
xnor U4571 (N_4571,N_4356,N_4402);
xnor U4572 (N_4572,N_3449,N_4105);
xnor U4573 (N_4573,N_4121,N_3040);
and U4574 (N_4574,N_4358,N_3409);
or U4575 (N_4575,N_4129,N_4141);
xnor U4576 (N_4576,N_3865,N_3716);
and U4577 (N_4577,N_3301,N_4200);
and U4578 (N_4578,N_3381,N_3783);
nor U4579 (N_4579,N_3360,N_3129);
and U4580 (N_4580,N_4126,N_4065);
xor U4581 (N_4581,N_4474,N_3818);
xnor U4582 (N_4582,N_4246,N_4051);
or U4583 (N_4583,N_3453,N_3112);
and U4584 (N_4584,N_4499,N_4470);
nand U4585 (N_4585,N_3574,N_3328);
nand U4586 (N_4586,N_3639,N_4438);
or U4587 (N_4587,N_4106,N_4339);
nor U4588 (N_4588,N_4101,N_4361);
nand U4589 (N_4589,N_3419,N_3086);
xnor U4590 (N_4590,N_3977,N_4367);
or U4591 (N_4591,N_3276,N_4318);
nor U4592 (N_4592,N_3683,N_3718);
xor U4593 (N_4593,N_3109,N_3335);
xor U4594 (N_4594,N_4300,N_3151);
and U4595 (N_4595,N_3580,N_3407);
nand U4596 (N_4596,N_4467,N_4083);
and U4597 (N_4597,N_4331,N_3216);
or U4598 (N_4598,N_3704,N_4120);
nor U4599 (N_4599,N_4424,N_4251);
and U4600 (N_4600,N_4456,N_4062);
and U4601 (N_4601,N_3493,N_3339);
xnor U4602 (N_4602,N_3118,N_3791);
or U4603 (N_4603,N_3728,N_3104);
xor U4604 (N_4604,N_3969,N_3022);
xor U4605 (N_4605,N_3751,N_3263);
xor U4606 (N_4606,N_3473,N_3971);
nand U4607 (N_4607,N_3637,N_3864);
and U4608 (N_4608,N_3568,N_3570);
nor U4609 (N_4609,N_4213,N_3841);
and U4610 (N_4610,N_3035,N_4400);
xor U4611 (N_4611,N_3305,N_3603);
and U4612 (N_4612,N_3550,N_4365);
nor U4613 (N_4613,N_4374,N_3656);
nand U4614 (N_4614,N_3808,N_3847);
and U4615 (N_4615,N_4451,N_3005);
nor U4616 (N_4616,N_3862,N_3959);
nand U4617 (N_4617,N_3571,N_3776);
or U4618 (N_4618,N_3589,N_4132);
or U4619 (N_4619,N_3760,N_3933);
nor U4620 (N_4620,N_4158,N_3354);
and U4621 (N_4621,N_3586,N_4294);
xor U4622 (N_4622,N_3646,N_3533);
and U4623 (N_4623,N_4420,N_3239);
nor U4624 (N_4624,N_4317,N_3441);
nand U4625 (N_4625,N_3836,N_4348);
or U4626 (N_4626,N_3029,N_3201);
xor U4627 (N_4627,N_3458,N_3256);
nand U4628 (N_4628,N_3162,N_3262);
xor U4629 (N_4629,N_4137,N_3569);
xor U4630 (N_4630,N_3417,N_3928);
or U4631 (N_4631,N_3094,N_3423);
xor U4632 (N_4632,N_4311,N_3469);
nand U4633 (N_4633,N_3840,N_3553);
nand U4634 (N_4634,N_3025,N_3966);
nand U4635 (N_4635,N_3125,N_3158);
and U4636 (N_4636,N_3413,N_3529);
nor U4637 (N_4637,N_3804,N_4382);
xnor U4638 (N_4638,N_3882,N_3003);
and U4639 (N_4639,N_3171,N_3272);
nor U4640 (N_4640,N_4279,N_3373);
and U4641 (N_4641,N_3773,N_3894);
or U4642 (N_4642,N_3009,N_3254);
or U4643 (N_4643,N_3204,N_4270);
or U4644 (N_4644,N_4482,N_4153);
nor U4645 (N_4645,N_3377,N_3400);
xor U4646 (N_4646,N_3766,N_3772);
and U4647 (N_4647,N_3004,N_3269);
and U4648 (N_4648,N_3504,N_3041);
nand U4649 (N_4649,N_3471,N_3918);
nand U4650 (N_4650,N_3787,N_3524);
or U4651 (N_4651,N_3756,N_4168);
nor U4652 (N_4652,N_3560,N_4404);
xnor U4653 (N_4653,N_3761,N_3144);
nand U4654 (N_4654,N_3576,N_3505);
xnor U4655 (N_4655,N_3730,N_4159);
or U4656 (N_4656,N_4145,N_3531);
xnor U4657 (N_4657,N_3790,N_4401);
or U4658 (N_4658,N_4292,N_3793);
xnor U4659 (N_4659,N_3600,N_4188);
or U4660 (N_4660,N_3017,N_3884);
or U4661 (N_4661,N_3340,N_3544);
nor U4662 (N_4662,N_3391,N_3701);
and U4663 (N_4663,N_3643,N_3497);
or U4664 (N_4664,N_4192,N_3426);
nand U4665 (N_4665,N_3439,N_4032);
nand U4666 (N_4666,N_3217,N_3800);
and U4667 (N_4667,N_3421,N_3215);
nand U4668 (N_4668,N_3745,N_3659);
nor U4669 (N_4669,N_4108,N_3008);
xor U4670 (N_4670,N_3287,N_3374);
xor U4671 (N_4671,N_3579,N_3443);
or U4672 (N_4672,N_3820,N_3250);
nor U4673 (N_4673,N_3597,N_3775);
xor U4674 (N_4674,N_3117,N_4091);
or U4675 (N_4675,N_4175,N_3181);
nor U4676 (N_4676,N_3518,N_4418);
and U4677 (N_4677,N_3363,N_3175);
nand U4678 (N_4678,N_3512,N_3542);
nor U4679 (N_4679,N_3521,N_4056);
and U4680 (N_4680,N_3090,N_3653);
and U4681 (N_4681,N_3149,N_3609);
or U4682 (N_4682,N_3648,N_3480);
or U4683 (N_4683,N_3330,N_4086);
and U4684 (N_4684,N_4119,N_3997);
nor U4685 (N_4685,N_3834,N_3225);
and U4686 (N_4686,N_4329,N_3910);
nand U4687 (N_4687,N_4139,N_4022);
xnor U4688 (N_4688,N_3433,N_3916);
or U4689 (N_4689,N_4314,N_3489);
and U4690 (N_4690,N_3996,N_4258);
or U4691 (N_4691,N_4262,N_3306);
xnor U4692 (N_4692,N_4233,N_4184);
nor U4693 (N_4693,N_3901,N_3177);
nand U4694 (N_4694,N_3387,N_3725);
xnor U4695 (N_4695,N_3440,N_3142);
or U4696 (N_4696,N_3388,N_3610);
nand U4697 (N_4697,N_4441,N_3385);
and U4698 (N_4698,N_3605,N_4039);
and U4699 (N_4699,N_3270,N_3582);
nand U4700 (N_4700,N_3404,N_4248);
and U4701 (N_4701,N_3281,N_4340);
xnor U4702 (N_4702,N_3405,N_3392);
nor U4703 (N_4703,N_3986,N_3084);
nor U4704 (N_4704,N_4373,N_4107);
and U4705 (N_4705,N_4443,N_3880);
xnor U4706 (N_4706,N_4488,N_4027);
and U4707 (N_4707,N_4006,N_3243);
nand U4708 (N_4708,N_3468,N_4379);
nand U4709 (N_4709,N_4109,N_3152);
nand U4710 (N_4710,N_3652,N_4312);
and U4711 (N_4711,N_4138,N_4195);
nand U4712 (N_4712,N_3801,N_3849);
xnor U4713 (N_4713,N_3541,N_3535);
nor U4714 (N_4714,N_4070,N_3563);
xor U4715 (N_4715,N_3114,N_3103);
xnor U4716 (N_4716,N_3866,N_3345);
xnor U4717 (N_4717,N_3313,N_4231);
xor U4718 (N_4718,N_3001,N_4491);
and U4719 (N_4719,N_4479,N_3155);
nand U4720 (N_4720,N_4468,N_3973);
and U4721 (N_4721,N_4478,N_4334);
nand U4722 (N_4722,N_4172,N_3617);
nand U4723 (N_4723,N_3877,N_3014);
nor U4724 (N_4724,N_4199,N_3226);
nand U4725 (N_4725,N_3554,N_3043);
nand U4726 (N_4726,N_4209,N_3785);
nor U4727 (N_4727,N_4462,N_3422);
or U4728 (N_4728,N_4046,N_4309);
and U4729 (N_4729,N_3559,N_3989);
nor U4730 (N_4730,N_3455,N_4305);
nand U4731 (N_4731,N_3537,N_4421);
nor U4732 (N_4732,N_4015,N_4186);
nor U4733 (N_4733,N_3638,N_3167);
or U4734 (N_4734,N_3719,N_4193);
xnor U4735 (N_4735,N_4324,N_3081);
xnor U4736 (N_4736,N_3976,N_3689);
or U4737 (N_4737,N_3376,N_4031);
nor U4738 (N_4738,N_3558,N_3620);
nand U4739 (N_4739,N_4030,N_3771);
and U4740 (N_4740,N_4226,N_3596);
and U4741 (N_4741,N_3173,N_3307);
xnor U4742 (N_4742,N_4266,N_4178);
nor U4743 (N_4743,N_4253,N_3900);
nand U4744 (N_4744,N_3366,N_4362);
xnor U4745 (N_4745,N_3676,N_3583);
and U4746 (N_4746,N_3046,N_3194);
nor U4747 (N_4747,N_4277,N_4207);
and U4748 (N_4748,N_3658,N_4122);
nor U4749 (N_4749,N_3630,N_3798);
nor U4750 (N_4750,N_3805,N_3737);
xnor U4751 (N_4751,N_3165,N_4183);
or U4752 (N_4752,N_4264,N_4446);
and U4753 (N_4753,N_3578,N_3494);
nor U4754 (N_4754,N_3794,N_3372);
xor U4755 (N_4755,N_3264,N_3451);
nor U4756 (N_4756,N_3229,N_4323);
and U4757 (N_4757,N_3096,N_3464);
and U4758 (N_4758,N_4067,N_4016);
or U4759 (N_4759,N_4281,N_3510);
nor U4760 (N_4760,N_3147,N_4461);
or U4761 (N_4761,N_4419,N_3105);
nand U4762 (N_4762,N_3982,N_4476);
nor U4763 (N_4763,N_4090,N_3755);
or U4764 (N_4764,N_3506,N_4492);
nor U4765 (N_4765,N_3033,N_3692);
nand U4766 (N_4766,N_4263,N_3671);
xnor U4767 (N_4767,N_4077,N_3351);
nand U4768 (N_4768,N_4313,N_3534);
and U4769 (N_4769,N_4125,N_3288);
nand U4770 (N_4770,N_4388,N_3348);
nor U4771 (N_4771,N_4408,N_4146);
or U4772 (N_4772,N_3611,N_4260);
nor U4773 (N_4773,N_4273,N_3628);
nand U4774 (N_4774,N_4290,N_3319);
xnor U4775 (N_4775,N_3899,N_3599);
xor U4776 (N_4776,N_3724,N_4073);
xnor U4777 (N_4777,N_4196,N_3050);
or U4778 (N_4778,N_4002,N_3930);
or U4779 (N_4779,N_3779,N_3467);
nor U4780 (N_4780,N_3364,N_3462);
or U4781 (N_4781,N_3807,N_3995);
or U4782 (N_4782,N_3282,N_3067);
or U4783 (N_4783,N_4116,N_3827);
and U4784 (N_4784,N_4149,N_4230);
and U4785 (N_4785,N_4413,N_3091);
nand U4786 (N_4786,N_3641,N_4332);
xnor U4787 (N_4787,N_4346,N_3161);
and U4788 (N_4788,N_3178,N_3185);
nand U4789 (N_4789,N_3012,N_3530);
xnor U4790 (N_4790,N_4475,N_3686);
xor U4791 (N_4791,N_4384,N_3871);
xnor U4792 (N_4792,N_4177,N_3828);
nand U4793 (N_4793,N_3509,N_3253);
xnor U4794 (N_4794,N_3293,N_3224);
nor U4795 (N_4795,N_3106,N_4487);
and U4796 (N_4796,N_3612,N_3206);
xor U4797 (N_4797,N_3874,N_3054);
nor U4798 (N_4798,N_4286,N_3294);
xnor U4799 (N_4799,N_3230,N_4432);
xnor U4800 (N_4800,N_3286,N_3028);
xnor U4801 (N_4801,N_3934,N_3546);
nor U4802 (N_4802,N_4472,N_4026);
and U4803 (N_4803,N_3561,N_4118);
xnor U4804 (N_4804,N_4204,N_3116);
nor U4805 (N_4805,N_3097,N_4010);
or U4806 (N_4806,N_3133,N_4437);
nor U4807 (N_4807,N_4363,N_4211);
or U4808 (N_4808,N_3334,N_4014);
nand U4809 (N_4809,N_3291,N_4161);
or U4810 (N_4810,N_3631,N_3245);
and U4811 (N_4811,N_4397,N_3551);
nand U4812 (N_4812,N_3633,N_3833);
nand U4813 (N_4813,N_3613,N_3577);
nor U4814 (N_4814,N_4060,N_4072);
or U4815 (N_4815,N_3954,N_3727);
and U4816 (N_4816,N_4350,N_3655);
or U4817 (N_4817,N_3280,N_3859);
or U4818 (N_4818,N_3703,N_3528);
nand U4819 (N_4819,N_3675,N_4299);
or U4820 (N_4820,N_4497,N_3781);
xor U4821 (N_4821,N_3350,N_3051);
nand U4822 (N_4822,N_3629,N_3031);
nand U4823 (N_4823,N_3427,N_3169);
nor U4824 (N_4824,N_3341,N_3402);
nand U4825 (N_4825,N_3732,N_3298);
or U4826 (N_4826,N_3073,N_3450);
xnor U4827 (N_4827,N_4490,N_3077);
nand U4828 (N_4828,N_3383,N_3904);
and U4829 (N_4829,N_4498,N_3297);
xor U4830 (N_4830,N_3697,N_3644);
xnor U4831 (N_4831,N_3870,N_3187);
nand U4832 (N_4832,N_3285,N_3212);
and U4833 (N_4833,N_3914,N_3353);
and U4834 (N_4834,N_3164,N_4282);
nand U4835 (N_4835,N_3278,N_3664);
and U4836 (N_4836,N_3712,N_3527);
or U4837 (N_4837,N_3102,N_4269);
nor U4838 (N_4838,N_3238,N_4463);
xor U4839 (N_4839,N_3770,N_3809);
or U4840 (N_4840,N_4321,N_4117);
xnor U4841 (N_4841,N_4355,N_4267);
xor U4842 (N_4842,N_4179,N_3030);
nor U4843 (N_4843,N_4357,N_3411);
nand U4844 (N_4844,N_3929,N_3935);
or U4845 (N_4845,N_3964,N_3907);
nor U4846 (N_4846,N_3764,N_3895);
nand U4847 (N_4847,N_3447,N_3988);
xnor U4848 (N_4848,N_3975,N_3499);
nor U4849 (N_4849,N_3592,N_4130);
or U4850 (N_4850,N_3064,N_3386);
and U4851 (N_4851,N_3516,N_4364);
and U4852 (N_4852,N_4288,N_4430);
or U4853 (N_4853,N_3598,N_4338);
xnor U4854 (N_4854,N_3816,N_3242);
xnor U4855 (N_4855,N_4349,N_3957);
or U4856 (N_4856,N_3670,N_3011);
and U4857 (N_4857,N_3072,N_3711);
or U4858 (N_4858,N_3851,N_3362);
nor U4859 (N_4859,N_3709,N_3896);
xnor U4860 (N_4860,N_3331,N_3186);
and U4861 (N_4861,N_4042,N_3352);
xnor U4862 (N_4862,N_3902,N_3673);
and U4863 (N_4863,N_4345,N_4394);
nor U4864 (N_4864,N_3890,N_4208);
or U4865 (N_4865,N_4075,N_3759);
xor U4866 (N_4866,N_4133,N_3717);
xnor U4867 (N_4867,N_3843,N_4489);
xor U4868 (N_4868,N_4111,N_3107);
or U4869 (N_4869,N_3110,N_3438);
nand U4870 (N_4870,N_3741,N_3545);
nand U4871 (N_4871,N_3338,N_3744);
nor U4872 (N_4872,N_3398,N_4354);
and U4873 (N_4873,N_3687,N_4427);
nor U4874 (N_4874,N_3721,N_3786);
and U4875 (N_4875,N_3562,N_4228);
or U4876 (N_4876,N_3758,N_4148);
and U4877 (N_4877,N_4041,N_3838);
xor U4878 (N_4878,N_3752,N_4045);
nor U4879 (N_4879,N_3240,N_3395);
and U4880 (N_4880,N_4104,N_4055);
xnor U4881 (N_4881,N_3058,N_4088);
or U4882 (N_4882,N_4422,N_3188);
xor U4883 (N_4883,N_3099,N_4054);
xnor U4884 (N_4884,N_4238,N_3415);
nor U4885 (N_4885,N_3735,N_3556);
or U4886 (N_4886,N_3461,N_4276);
xor U4887 (N_4887,N_3408,N_4096);
nand U4888 (N_4888,N_3690,N_3685);
nor U4889 (N_4889,N_3953,N_4154);
nor U4890 (N_4890,N_3765,N_3679);
nor U4891 (N_4891,N_3979,N_3795);
xnor U4892 (N_4892,N_3275,N_3621);
nand U4893 (N_4893,N_4112,N_4093);
nor U4894 (N_4894,N_3860,N_4103);
and U4895 (N_4895,N_4278,N_3784);
nand U4896 (N_4896,N_4216,N_3606);
xor U4897 (N_4897,N_4189,N_3994);
nor U4898 (N_4898,N_3604,N_3359);
nor U4899 (N_4899,N_3696,N_3640);
nand U4900 (N_4900,N_3199,N_3909);
nor U4901 (N_4901,N_3567,N_3811);
or U4902 (N_4902,N_4134,N_3049);
or U4903 (N_4903,N_4452,N_3429);
nand U4904 (N_4904,N_4143,N_3519);
and U4905 (N_4905,N_3898,N_3179);
or U4906 (N_4906,N_4391,N_3999);
nand U4907 (N_4907,N_4205,N_4100);
nor U4908 (N_4908,N_4150,N_4224);
nand U4909 (N_4909,N_4411,N_4257);
nor U4910 (N_4910,N_4048,N_3015);
nand U4911 (N_4911,N_3845,N_3132);
nand U4912 (N_4912,N_3342,N_4389);
and U4913 (N_4913,N_3266,N_3587);
xnor U4914 (N_4914,N_3057,N_3310);
nor U4915 (N_4915,N_3214,N_4429);
nor U4916 (N_4916,N_3312,N_3052);
xnor U4917 (N_4917,N_3939,N_4434);
and U4918 (N_4918,N_3356,N_4341);
nor U4919 (N_4919,N_3261,N_3343);
nand U4920 (N_4920,N_3234,N_4092);
nor U4921 (N_4921,N_4428,N_3182);
and U4922 (N_4922,N_3146,N_3034);
nand U4923 (N_4923,N_3594,N_4135);
nor U4924 (N_4924,N_4366,N_4214);
xnor U4925 (N_4925,N_4306,N_4254);
nand U4926 (N_4926,N_3024,N_3483);
and U4927 (N_4927,N_3336,N_4274);
nand U4928 (N_4928,N_4271,N_3799);
or U4929 (N_4929,N_3536,N_4221);
nor U4930 (N_4930,N_4079,N_4037);
and U4931 (N_4931,N_3889,N_3668);
nand U4932 (N_4932,N_4457,N_3349);
xor U4933 (N_4933,N_3706,N_3515);
and U4934 (N_4934,N_3564,N_3076);
and U4935 (N_4935,N_3747,N_3672);
xnor U4936 (N_4936,N_3526,N_3674);
or U4937 (N_4937,N_3825,N_3523);
or U4938 (N_4938,N_4018,N_4173);
nor U4939 (N_4939,N_3231,N_3595);
nor U4940 (N_4940,N_4308,N_3998);
or U4941 (N_4941,N_4403,N_3274);
xor U4942 (N_4942,N_4052,N_4433);
nor U4943 (N_4943,N_4212,N_4298);
xor U4944 (N_4944,N_3127,N_3476);
xor U4945 (N_4945,N_4004,N_3822);
and U4946 (N_4946,N_4021,N_3258);
xor U4947 (N_4947,N_3543,N_3919);
nand U4948 (N_4948,N_3835,N_4359);
or U4949 (N_4949,N_4435,N_3698);
or U4950 (N_4950,N_4099,N_3235);
or U4951 (N_4951,N_3498,N_3548);
or U4952 (N_4952,N_4191,N_3774);
or U4953 (N_4953,N_3252,N_3198);
nor U4954 (N_4954,N_3487,N_3037);
nor U4955 (N_4955,N_3740,N_4436);
nor U4956 (N_4956,N_3940,N_4024);
nand U4957 (N_4957,N_3681,N_3170);
and U4958 (N_4958,N_3055,N_3053);
nand U4959 (N_4959,N_3942,N_3736);
or U4960 (N_4960,N_3157,N_4336);
or U4961 (N_4961,N_3130,N_3174);
xnor U4962 (N_4962,N_3723,N_3365);
xor U4963 (N_4963,N_4335,N_3700);
nand U4964 (N_4964,N_3318,N_3205);
and U4965 (N_4965,N_3358,N_4343);
nand U4966 (N_4966,N_4087,N_3075);
nor U4967 (N_4967,N_3379,N_3814);
and U4968 (N_4968,N_3768,N_4471);
nand U4969 (N_4969,N_4453,N_3098);
and U4970 (N_4970,N_3903,N_4370);
xor U4971 (N_4971,N_3380,N_3680);
or U4972 (N_4972,N_3626,N_3951);
or U4973 (N_4973,N_3917,N_3460);
and U4974 (N_4974,N_4439,N_4007);
xor U4975 (N_4975,N_3477,N_3332);
nand U4976 (N_4976,N_4097,N_4328);
and U4977 (N_4977,N_3960,N_3684);
xnor U4978 (N_4978,N_4480,N_3944);
or U4979 (N_4979,N_3990,N_3763);
nor U4980 (N_4980,N_3200,N_3000);
and U4981 (N_4981,N_4395,N_3636);
nor U4982 (N_4982,N_4284,N_4245);
xnor U4983 (N_4983,N_3131,N_3071);
or U4984 (N_4984,N_3788,N_4296);
nand U4985 (N_4985,N_3486,N_3311);
nand U4986 (N_4986,N_3042,N_3863);
xnor U4987 (N_4987,N_4301,N_3502);
nand U4988 (N_4988,N_3555,N_4001);
nor U4989 (N_4989,N_4376,N_3767);
nand U4990 (N_4990,N_4131,N_4076);
nand U4991 (N_4991,N_3869,N_3326);
nor U4992 (N_4992,N_3573,N_4155);
and U4993 (N_4993,N_4124,N_4110);
nor U4994 (N_4994,N_4176,N_3208);
nor U4995 (N_4995,N_3962,N_4123);
nand U4996 (N_4996,N_3465,N_3852);
nor U4997 (N_4997,N_4242,N_3867);
or U4998 (N_4998,N_3403,N_3588);
xor U4999 (N_4999,N_3474,N_3950);
xor U5000 (N_5000,N_4378,N_3762);
nor U5001 (N_5001,N_4068,N_3495);
xor U5002 (N_5002,N_3065,N_4128);
or U5003 (N_5003,N_3044,N_3384);
and U5004 (N_5004,N_4082,N_3424);
nand U5005 (N_5005,N_4320,N_3304);
or U5006 (N_5006,N_3168,N_3183);
nand U5007 (N_5007,N_3432,N_4163);
or U5008 (N_5008,N_4495,N_3488);
nor U5009 (N_5009,N_3300,N_3361);
xor U5010 (N_5010,N_4493,N_4033);
nand U5011 (N_5011,N_3207,N_4285);
nand U5012 (N_5012,N_3394,N_4353);
and U5013 (N_5013,N_3842,N_4410);
xor U5014 (N_5014,N_4236,N_3984);
nand U5015 (N_5015,N_3955,N_3481);
and U5016 (N_5016,N_3092,N_3936);
nor U5017 (N_5017,N_3846,N_4162);
nor U5018 (N_5018,N_3284,N_3821);
xor U5019 (N_5019,N_3093,N_3246);
or U5020 (N_5020,N_3197,N_3945);
nor U5021 (N_5021,N_3665,N_3710);
or U5022 (N_5022,N_3729,N_3475);
nor U5023 (N_5023,N_3434,N_3713);
or U5024 (N_5024,N_4352,N_3708);
or U5025 (N_5025,N_4442,N_3321);
nor U5026 (N_5026,N_4454,N_3797);
or U5027 (N_5027,N_4166,N_3678);
or U5028 (N_5028,N_3355,N_3754);
xnor U5029 (N_5029,N_4360,N_4448);
xor U5030 (N_5030,N_3925,N_3101);
and U5031 (N_5031,N_3273,N_3143);
xnor U5032 (N_5032,N_3522,N_4220);
xnor U5033 (N_5033,N_4431,N_3399);
and U5034 (N_5034,N_4069,N_4080);
xor U5035 (N_5035,N_4181,N_3062);
nor U5036 (N_5036,N_4268,N_4053);
or U5037 (N_5037,N_3192,N_4061);
and U5038 (N_5038,N_4225,N_4265);
nand U5039 (N_5039,N_3651,N_4035);
nand U5040 (N_5040,N_3911,N_3591);
or U5041 (N_5041,N_4375,N_3844);
nand U5042 (N_5042,N_3145,N_3333);
or U5043 (N_5043,N_3317,N_4038);
xor U5044 (N_5044,N_4218,N_4084);
and U5045 (N_5045,N_3066,N_3369);
xnor U5046 (N_5046,N_3581,N_4396);
xor U5047 (N_5047,N_3557,N_3299);
and U5048 (N_5048,N_3069,N_3088);
nor U5049 (N_5049,N_3908,N_3457);
xor U5050 (N_5050,N_3211,N_4171);
xor U5051 (N_5051,N_4217,N_3949);
nor U5052 (N_5052,N_3985,N_3150);
xnor U5053 (N_5053,N_3868,N_3623);
or U5054 (N_5054,N_3748,N_4227);
and U5055 (N_5055,N_3812,N_3397);
or U5056 (N_5056,N_3823,N_3232);
xor U5057 (N_5057,N_3585,N_4459);
nor U5058 (N_5058,N_3371,N_3649);
and U5059 (N_5059,N_4372,N_3858);
xor U5060 (N_5060,N_4304,N_3906);
nor U5061 (N_5061,N_3289,N_3726);
and U5062 (N_5062,N_4003,N_3501);
nand U5063 (N_5063,N_3707,N_4043);
or U5064 (N_5064,N_3532,N_4302);
nand U5065 (N_5065,N_4250,N_4012);
xnor U5066 (N_5066,N_4333,N_4392);
nor U5067 (N_5067,N_3881,N_3314);
nor U5068 (N_5068,N_3203,N_3016);
nor U5069 (N_5069,N_4057,N_3141);
nand U5070 (N_5070,N_4369,N_3113);
nor U5071 (N_5071,N_3470,N_3691);
xor U5072 (N_5072,N_3492,N_3176);
xnor U5073 (N_5073,N_4078,N_3210);
nor U5074 (N_5074,N_3061,N_3972);
and U5075 (N_5075,N_4008,N_4440);
or U5076 (N_5076,N_3593,N_3416);
and U5077 (N_5077,N_4390,N_4185);
xnor U5078 (N_5078,N_4426,N_3121);
and U5079 (N_5079,N_4464,N_3320);
nand U5080 (N_5080,N_4028,N_4399);
xor U5081 (N_5081,N_3247,N_3886);
xor U5082 (N_5082,N_3295,N_3669);
nand U5083 (N_5083,N_3309,N_3414);
nand U5084 (N_5084,N_3271,N_3410);
nand U5085 (N_5085,N_4398,N_3442);
or U5086 (N_5086,N_3978,N_4215);
nor U5087 (N_5087,N_3249,N_4310);
xor U5088 (N_5088,N_4050,N_4102);
xnor U5089 (N_5089,N_4444,N_3888);
and U5090 (N_5090,N_4156,N_3233);
nand U5091 (N_5091,N_4483,N_3887);
and U5092 (N_5092,N_3699,N_3824);
or U5093 (N_5093,N_3139,N_4020);
nand U5094 (N_5094,N_4351,N_3540);
and U5095 (N_5095,N_3927,N_3277);
nand U5096 (N_5096,N_3660,N_3479);
nor U5097 (N_5097,N_3923,N_3490);
nor U5098 (N_5098,N_3584,N_3412);
xnor U5099 (N_5099,N_3607,N_3952);
xnor U5100 (N_5100,N_3166,N_3063);
and U5101 (N_5101,N_4011,N_3180);
or U5102 (N_5102,N_3915,N_3159);
and U5103 (N_5103,N_4252,N_3757);
xor U5104 (N_5104,N_4386,N_4330);
and U5105 (N_5105,N_3875,N_3682);
nand U5106 (N_5106,N_3782,N_3463);
nand U5107 (N_5107,N_4344,N_3993);
nand U5108 (N_5108,N_3446,N_3456);
and U5109 (N_5109,N_4114,N_4019);
nand U5110 (N_5110,N_4244,N_4180);
nor U5111 (N_5111,N_4280,N_3921);
nand U5112 (N_5112,N_3632,N_4098);
or U5113 (N_5113,N_4140,N_3625);
nor U5114 (N_5114,N_4239,N_3742);
xnor U5115 (N_5115,N_3370,N_4089);
and U5116 (N_5116,N_3236,N_3436);
or U5117 (N_5117,N_4034,N_3958);
nand U5118 (N_5118,N_3694,N_3857);
xnor U5119 (N_5119,N_4182,N_3733);
xnor U5120 (N_5120,N_4465,N_3854);
nor U5121 (N_5121,N_3810,N_4113);
nand U5122 (N_5122,N_4327,N_4289);
or U5123 (N_5123,N_3663,N_3992);
and U5124 (N_5124,N_4234,N_3279);
nand U5125 (N_5125,N_3156,N_4325);
xnor U5126 (N_5126,N_3885,N_4416);
xnor U5127 (N_5127,N_3406,N_3657);
nand U5128 (N_5128,N_4095,N_3454);
nor U5129 (N_5129,N_4415,N_3303);
nand U5130 (N_5130,N_3778,N_3484);
and U5131 (N_5131,N_3074,N_3209);
and U5132 (N_5132,N_3257,N_3792);
xor U5133 (N_5133,N_4380,N_4142);
xor U5134 (N_5134,N_3974,N_3248);
or U5135 (N_5135,N_4425,N_3861);
or U5136 (N_5136,N_3572,N_3500);
nor U5137 (N_5137,N_3115,N_3891);
nand U5138 (N_5138,N_3963,N_3832);
nor U5139 (N_5139,N_3196,N_3140);
nor U5140 (N_5140,N_4115,N_4029);
nand U5141 (N_5141,N_4307,N_3327);
nand U5142 (N_5142,N_3083,N_3912);
and U5143 (N_5143,N_3138,N_3087);
nor U5144 (N_5144,N_4243,N_4496);
or U5145 (N_5145,N_3948,N_3883);
nand U5146 (N_5146,N_3006,N_3218);
nor U5147 (N_5147,N_3722,N_4219);
nand U5148 (N_5148,N_3947,N_4417);
xor U5149 (N_5149,N_3507,N_3734);
nand U5150 (N_5150,N_3172,N_3195);
or U5151 (N_5151,N_3123,N_3667);
and U5152 (N_5152,N_3382,N_4445);
nand U5153 (N_5153,N_3126,N_3060);
nor U5154 (N_5154,N_3991,N_3539);
and U5155 (N_5155,N_4059,N_3549);
nand U5156 (N_5156,N_4423,N_4237);
or U5157 (N_5157,N_3720,N_3324);
xnor U5158 (N_5158,N_3023,N_3026);
xnor U5159 (N_5159,N_3922,N_3654);
and U5160 (N_5160,N_3325,N_3428);
nor U5161 (N_5161,N_4377,N_4127);
nand U5162 (N_5162,N_4450,N_3946);
nand U5163 (N_5163,N_3111,N_4347);
nand U5164 (N_5164,N_3746,N_3839);
xor U5165 (N_5165,N_3853,N_4407);
nor U5166 (N_5166,N_4322,N_3095);
and U5167 (N_5167,N_3715,N_3190);
and U5168 (N_5168,N_4167,N_3108);
and U5169 (N_5169,N_4160,N_3322);
or U5170 (N_5170,N_3265,N_3047);
nor U5171 (N_5171,N_4164,N_3789);
or U5172 (N_5172,N_3222,N_4287);
or U5173 (N_5173,N_3221,N_3122);
nor U5174 (N_5174,N_4249,N_3855);
and U5175 (N_5175,N_3956,N_3753);
or U5176 (N_5176,N_3202,N_3920);
xnor U5177 (N_5177,N_4469,N_3513);
nand U5178 (N_5178,N_3478,N_4170);
or U5179 (N_5179,N_4241,N_3260);
xor U5180 (N_5180,N_3119,N_4198);
nand U5181 (N_5181,N_3038,N_3445);
nor U5182 (N_5182,N_3193,N_3021);
or U5183 (N_5183,N_4203,N_3425);
xor U5184 (N_5184,N_3967,N_3120);
and U5185 (N_5185,N_3393,N_3255);
xor U5186 (N_5186,N_4165,N_4202);
or U5187 (N_5187,N_3856,N_3892);
nor U5188 (N_5188,N_4326,N_3796);
or U5189 (N_5189,N_3244,N_3743);
nand U5190 (N_5190,N_3941,N_4486);
xor U5191 (N_5191,N_3002,N_3048);
nor U5192 (N_5192,N_3346,N_4406);
xor U5193 (N_5193,N_4235,N_3634);
xor U5194 (N_5194,N_3085,N_4405);
xnor U5195 (N_5195,N_4009,N_3924);
nor U5196 (N_5196,N_3448,N_4081);
nand U5197 (N_5197,N_4071,N_3780);
nor U5198 (N_5198,N_3661,N_3396);
nor U5199 (N_5199,N_3520,N_4481);
or U5200 (N_5200,N_4297,N_4232);
or U5201 (N_5201,N_3010,N_3897);
nor U5202 (N_5202,N_3045,N_3817);
nor U5203 (N_5203,N_3614,N_3228);
nor U5204 (N_5204,N_4484,N_4066);
or U5205 (N_5205,N_3750,N_4409);
and U5206 (N_5206,N_3082,N_3645);
nor U5207 (N_5207,N_3552,N_3259);
nor U5208 (N_5208,N_4368,N_3401);
nand U5209 (N_5209,N_4240,N_3938);
and U5210 (N_5210,N_3357,N_3227);
nand U5211 (N_5211,N_3819,N_3806);
xnor U5212 (N_5212,N_4151,N_3124);
nor U5213 (N_5213,N_3223,N_3538);
or U5214 (N_5214,N_4157,N_3347);
and U5215 (N_5215,N_4303,N_3872);
xnor U5216 (N_5216,N_3616,N_4383);
nor U5217 (N_5217,N_3635,N_3431);
nor U5218 (N_5218,N_3019,N_3007);
nand U5219 (N_5219,N_3390,N_4255);
nand U5220 (N_5220,N_3389,N_3148);
xor U5221 (N_5221,N_3601,N_3937);
and U5222 (N_5222,N_3308,N_3482);
xor U5223 (N_5223,N_4342,N_3323);
nor U5224 (N_5224,N_4316,N_3803);
xnor U5225 (N_5225,N_3566,N_3738);
or U5226 (N_5226,N_3893,N_4387);
and U5227 (N_5227,N_3987,N_3068);
or U5228 (N_5228,N_3128,N_3367);
and U5229 (N_5229,N_3693,N_3970);
and U5230 (N_5230,N_3565,N_3136);
xnor U5231 (N_5231,N_4371,N_3036);
nor U5232 (N_5232,N_3213,N_4040);
and U5233 (N_5233,N_3815,N_3283);
nor U5234 (N_5234,N_3731,N_4136);
nor U5235 (N_5235,N_3968,N_4261);
or U5236 (N_5236,N_3267,N_3702);
and U5237 (N_5237,N_4256,N_3547);
and U5238 (N_5238,N_3302,N_3251);
and U5239 (N_5239,N_3650,N_3219);
nand U5240 (N_5240,N_3980,N_4049);
or U5241 (N_5241,N_4094,N_3848);
nor U5242 (N_5242,N_4000,N_3831);
or U5243 (N_5243,N_3496,N_4064);
nor U5244 (N_5244,N_3296,N_4085);
or U5245 (N_5245,N_4477,N_4058);
nand U5246 (N_5246,N_4473,N_4412);
and U5247 (N_5247,N_3688,N_3241);
nand U5248 (N_5248,N_3618,N_3444);
nand U5249 (N_5249,N_3873,N_3452);
and U5250 (N_5250,N_3723,N_3604);
and U5251 (N_5251,N_3753,N_3344);
and U5252 (N_5252,N_3211,N_4241);
xor U5253 (N_5253,N_3940,N_3188);
or U5254 (N_5254,N_3030,N_3444);
nand U5255 (N_5255,N_4147,N_3399);
xnor U5256 (N_5256,N_4293,N_3900);
nor U5257 (N_5257,N_4025,N_4069);
or U5258 (N_5258,N_4375,N_3552);
and U5259 (N_5259,N_3203,N_3979);
and U5260 (N_5260,N_3794,N_3750);
xor U5261 (N_5261,N_3116,N_4460);
or U5262 (N_5262,N_3554,N_3606);
or U5263 (N_5263,N_4448,N_3957);
xor U5264 (N_5264,N_4293,N_4367);
and U5265 (N_5265,N_4207,N_3762);
nand U5266 (N_5266,N_4426,N_3815);
xnor U5267 (N_5267,N_3474,N_3713);
nand U5268 (N_5268,N_3363,N_3040);
and U5269 (N_5269,N_4436,N_3325);
nand U5270 (N_5270,N_3783,N_3608);
nand U5271 (N_5271,N_3307,N_4308);
or U5272 (N_5272,N_3347,N_3204);
and U5273 (N_5273,N_3497,N_3353);
nand U5274 (N_5274,N_3686,N_3155);
nor U5275 (N_5275,N_3344,N_3219);
nor U5276 (N_5276,N_3610,N_4158);
nand U5277 (N_5277,N_4448,N_3188);
or U5278 (N_5278,N_4185,N_4169);
and U5279 (N_5279,N_3017,N_3987);
nor U5280 (N_5280,N_3084,N_3116);
nor U5281 (N_5281,N_3268,N_3929);
and U5282 (N_5282,N_3637,N_3003);
nand U5283 (N_5283,N_4469,N_3378);
xnor U5284 (N_5284,N_3848,N_3564);
xnor U5285 (N_5285,N_4244,N_3869);
nand U5286 (N_5286,N_3890,N_3233);
nor U5287 (N_5287,N_4126,N_4486);
and U5288 (N_5288,N_3130,N_4285);
xnor U5289 (N_5289,N_3584,N_4021);
nand U5290 (N_5290,N_4193,N_3952);
nand U5291 (N_5291,N_3691,N_3827);
nand U5292 (N_5292,N_3276,N_3870);
or U5293 (N_5293,N_3856,N_4142);
nor U5294 (N_5294,N_3760,N_3817);
nand U5295 (N_5295,N_4204,N_3630);
nand U5296 (N_5296,N_4399,N_3974);
nand U5297 (N_5297,N_3356,N_3510);
nand U5298 (N_5298,N_3987,N_4335);
nand U5299 (N_5299,N_4457,N_3646);
and U5300 (N_5300,N_4258,N_4411);
or U5301 (N_5301,N_3714,N_3915);
nor U5302 (N_5302,N_3028,N_3182);
xor U5303 (N_5303,N_3956,N_3732);
xor U5304 (N_5304,N_3871,N_4348);
or U5305 (N_5305,N_3524,N_4361);
or U5306 (N_5306,N_3383,N_3723);
nor U5307 (N_5307,N_3742,N_4442);
nor U5308 (N_5308,N_4111,N_3407);
nor U5309 (N_5309,N_3787,N_3151);
and U5310 (N_5310,N_3743,N_4300);
or U5311 (N_5311,N_4314,N_3412);
nand U5312 (N_5312,N_4047,N_3446);
nor U5313 (N_5313,N_3834,N_3929);
nand U5314 (N_5314,N_3501,N_3246);
nand U5315 (N_5315,N_3161,N_4460);
nor U5316 (N_5316,N_3687,N_3174);
or U5317 (N_5317,N_4036,N_3240);
xor U5318 (N_5318,N_3239,N_3359);
or U5319 (N_5319,N_4459,N_3334);
xnor U5320 (N_5320,N_4183,N_4107);
xnor U5321 (N_5321,N_4330,N_3600);
or U5322 (N_5322,N_4417,N_4222);
or U5323 (N_5323,N_3249,N_3081);
xor U5324 (N_5324,N_4322,N_3203);
or U5325 (N_5325,N_4179,N_3657);
nand U5326 (N_5326,N_3430,N_3622);
xor U5327 (N_5327,N_4197,N_3676);
and U5328 (N_5328,N_3817,N_4311);
or U5329 (N_5329,N_3233,N_4406);
or U5330 (N_5330,N_3098,N_3685);
and U5331 (N_5331,N_4348,N_3495);
and U5332 (N_5332,N_4433,N_4497);
xor U5333 (N_5333,N_3458,N_4372);
nor U5334 (N_5334,N_4078,N_3492);
xnor U5335 (N_5335,N_3297,N_4006);
or U5336 (N_5336,N_4450,N_3499);
xnor U5337 (N_5337,N_3469,N_3786);
and U5338 (N_5338,N_3274,N_3121);
and U5339 (N_5339,N_3650,N_3405);
and U5340 (N_5340,N_4199,N_3732);
or U5341 (N_5341,N_3275,N_3703);
or U5342 (N_5342,N_3785,N_4427);
nor U5343 (N_5343,N_3708,N_3187);
nor U5344 (N_5344,N_3692,N_3027);
xnor U5345 (N_5345,N_3991,N_3190);
or U5346 (N_5346,N_3129,N_4133);
xor U5347 (N_5347,N_4243,N_3762);
or U5348 (N_5348,N_3225,N_3232);
or U5349 (N_5349,N_3108,N_3269);
and U5350 (N_5350,N_4147,N_4173);
or U5351 (N_5351,N_4485,N_4044);
or U5352 (N_5352,N_4214,N_4268);
nor U5353 (N_5353,N_3940,N_4240);
or U5354 (N_5354,N_4215,N_3848);
xnor U5355 (N_5355,N_3063,N_3673);
or U5356 (N_5356,N_4105,N_3192);
nor U5357 (N_5357,N_3405,N_3063);
xnor U5358 (N_5358,N_4119,N_3202);
or U5359 (N_5359,N_4491,N_3979);
or U5360 (N_5360,N_3700,N_3287);
xnor U5361 (N_5361,N_3689,N_4209);
nor U5362 (N_5362,N_4162,N_4381);
nand U5363 (N_5363,N_3880,N_4487);
and U5364 (N_5364,N_4279,N_3634);
nand U5365 (N_5365,N_3060,N_4467);
or U5366 (N_5366,N_3647,N_4014);
nor U5367 (N_5367,N_4381,N_3704);
or U5368 (N_5368,N_3932,N_3557);
xor U5369 (N_5369,N_3713,N_3541);
and U5370 (N_5370,N_4299,N_3872);
or U5371 (N_5371,N_3949,N_3226);
nor U5372 (N_5372,N_4106,N_4111);
nand U5373 (N_5373,N_3512,N_3344);
nor U5374 (N_5374,N_3252,N_3736);
nand U5375 (N_5375,N_3746,N_3146);
nand U5376 (N_5376,N_3044,N_4385);
nor U5377 (N_5377,N_3485,N_4183);
nand U5378 (N_5378,N_3525,N_4207);
or U5379 (N_5379,N_4154,N_3716);
or U5380 (N_5380,N_4424,N_3042);
and U5381 (N_5381,N_4312,N_3934);
and U5382 (N_5382,N_4446,N_3962);
nand U5383 (N_5383,N_4447,N_4453);
nand U5384 (N_5384,N_4067,N_3919);
nor U5385 (N_5385,N_4184,N_4227);
nand U5386 (N_5386,N_4400,N_3799);
nand U5387 (N_5387,N_4349,N_4393);
and U5388 (N_5388,N_3052,N_3501);
or U5389 (N_5389,N_3872,N_4387);
and U5390 (N_5390,N_3153,N_3790);
or U5391 (N_5391,N_4362,N_3449);
or U5392 (N_5392,N_3490,N_3015);
nor U5393 (N_5393,N_3650,N_4164);
xnor U5394 (N_5394,N_3318,N_3556);
or U5395 (N_5395,N_4374,N_4298);
xnor U5396 (N_5396,N_3035,N_4254);
nor U5397 (N_5397,N_4045,N_4182);
or U5398 (N_5398,N_4458,N_3542);
nand U5399 (N_5399,N_3107,N_4073);
xor U5400 (N_5400,N_3471,N_4378);
nor U5401 (N_5401,N_3087,N_3639);
and U5402 (N_5402,N_3147,N_3299);
nor U5403 (N_5403,N_3590,N_3963);
xor U5404 (N_5404,N_3782,N_3444);
nor U5405 (N_5405,N_4276,N_3757);
xor U5406 (N_5406,N_4407,N_4441);
nand U5407 (N_5407,N_3627,N_4214);
or U5408 (N_5408,N_3345,N_3024);
nor U5409 (N_5409,N_4390,N_3138);
nand U5410 (N_5410,N_4363,N_3623);
nor U5411 (N_5411,N_4049,N_3233);
xnor U5412 (N_5412,N_3005,N_3385);
nor U5413 (N_5413,N_4048,N_3901);
xor U5414 (N_5414,N_3767,N_3785);
xor U5415 (N_5415,N_3992,N_3890);
or U5416 (N_5416,N_4201,N_4012);
nand U5417 (N_5417,N_3674,N_4241);
or U5418 (N_5418,N_4210,N_3733);
xor U5419 (N_5419,N_3391,N_3482);
nor U5420 (N_5420,N_3255,N_3490);
nand U5421 (N_5421,N_3041,N_3319);
or U5422 (N_5422,N_3791,N_4201);
nand U5423 (N_5423,N_3645,N_3814);
xnor U5424 (N_5424,N_3821,N_3460);
nor U5425 (N_5425,N_3794,N_3207);
xnor U5426 (N_5426,N_4119,N_4102);
nand U5427 (N_5427,N_3607,N_4129);
nor U5428 (N_5428,N_3373,N_3418);
and U5429 (N_5429,N_3481,N_3466);
nor U5430 (N_5430,N_3228,N_4332);
nor U5431 (N_5431,N_3866,N_3563);
nand U5432 (N_5432,N_4385,N_3803);
or U5433 (N_5433,N_3618,N_4493);
or U5434 (N_5434,N_4366,N_3954);
nand U5435 (N_5435,N_4296,N_3423);
nand U5436 (N_5436,N_3325,N_4024);
nor U5437 (N_5437,N_3968,N_3143);
nor U5438 (N_5438,N_4107,N_3548);
or U5439 (N_5439,N_3981,N_4448);
nor U5440 (N_5440,N_3955,N_3218);
nand U5441 (N_5441,N_3376,N_3826);
nand U5442 (N_5442,N_3976,N_3974);
and U5443 (N_5443,N_3854,N_4235);
nand U5444 (N_5444,N_3677,N_3504);
xor U5445 (N_5445,N_4238,N_4259);
or U5446 (N_5446,N_3508,N_3092);
nand U5447 (N_5447,N_3429,N_3728);
nor U5448 (N_5448,N_4170,N_3798);
nor U5449 (N_5449,N_3540,N_3755);
nor U5450 (N_5450,N_3374,N_4371);
nand U5451 (N_5451,N_3485,N_3490);
xor U5452 (N_5452,N_3450,N_3623);
and U5453 (N_5453,N_3173,N_3910);
or U5454 (N_5454,N_3170,N_3380);
nor U5455 (N_5455,N_4422,N_3647);
xor U5456 (N_5456,N_3164,N_3738);
and U5457 (N_5457,N_4425,N_3147);
and U5458 (N_5458,N_4430,N_3134);
nand U5459 (N_5459,N_3909,N_3454);
xor U5460 (N_5460,N_4016,N_3116);
and U5461 (N_5461,N_3388,N_3246);
nand U5462 (N_5462,N_3972,N_3175);
nor U5463 (N_5463,N_4261,N_3750);
nor U5464 (N_5464,N_3019,N_3323);
and U5465 (N_5465,N_3990,N_4407);
and U5466 (N_5466,N_3646,N_3929);
or U5467 (N_5467,N_4259,N_3307);
and U5468 (N_5468,N_3139,N_3089);
or U5469 (N_5469,N_4333,N_3517);
xor U5470 (N_5470,N_3000,N_4356);
or U5471 (N_5471,N_4338,N_4318);
nand U5472 (N_5472,N_3456,N_3136);
xor U5473 (N_5473,N_3892,N_3185);
xnor U5474 (N_5474,N_3702,N_3824);
or U5475 (N_5475,N_3233,N_3258);
nor U5476 (N_5476,N_3072,N_3928);
xor U5477 (N_5477,N_3818,N_4228);
nand U5478 (N_5478,N_3649,N_4319);
or U5479 (N_5479,N_3565,N_3663);
or U5480 (N_5480,N_3236,N_4030);
and U5481 (N_5481,N_3775,N_3398);
or U5482 (N_5482,N_3817,N_3026);
and U5483 (N_5483,N_3277,N_3993);
nand U5484 (N_5484,N_4311,N_3537);
and U5485 (N_5485,N_3871,N_3145);
xor U5486 (N_5486,N_3964,N_3930);
xor U5487 (N_5487,N_4222,N_4270);
xnor U5488 (N_5488,N_4245,N_3833);
or U5489 (N_5489,N_3225,N_4138);
xor U5490 (N_5490,N_3490,N_3209);
nand U5491 (N_5491,N_4305,N_3074);
nand U5492 (N_5492,N_3122,N_3822);
nor U5493 (N_5493,N_3904,N_3495);
nor U5494 (N_5494,N_3557,N_3726);
nand U5495 (N_5495,N_4489,N_3356);
nand U5496 (N_5496,N_3613,N_4194);
and U5497 (N_5497,N_3031,N_3782);
or U5498 (N_5498,N_3791,N_3181);
nor U5499 (N_5499,N_4282,N_4303);
or U5500 (N_5500,N_4341,N_3471);
xnor U5501 (N_5501,N_4420,N_3769);
or U5502 (N_5502,N_3442,N_3519);
nor U5503 (N_5503,N_4441,N_3888);
xnor U5504 (N_5504,N_4089,N_3518);
xor U5505 (N_5505,N_4460,N_3241);
xor U5506 (N_5506,N_4079,N_3198);
nand U5507 (N_5507,N_4127,N_3748);
and U5508 (N_5508,N_4290,N_3931);
or U5509 (N_5509,N_3425,N_4030);
and U5510 (N_5510,N_4414,N_3332);
or U5511 (N_5511,N_3673,N_4043);
or U5512 (N_5512,N_3660,N_3355);
nor U5513 (N_5513,N_4201,N_3870);
nand U5514 (N_5514,N_3691,N_3843);
nor U5515 (N_5515,N_3052,N_3182);
xnor U5516 (N_5516,N_3445,N_4181);
nand U5517 (N_5517,N_3373,N_4170);
nor U5518 (N_5518,N_3405,N_3353);
or U5519 (N_5519,N_3235,N_3292);
and U5520 (N_5520,N_3063,N_4214);
and U5521 (N_5521,N_4036,N_3357);
or U5522 (N_5522,N_3380,N_3932);
nor U5523 (N_5523,N_3873,N_3717);
nor U5524 (N_5524,N_3807,N_3320);
nor U5525 (N_5525,N_3503,N_4194);
or U5526 (N_5526,N_4307,N_3541);
or U5527 (N_5527,N_3791,N_3990);
and U5528 (N_5528,N_4224,N_4099);
nand U5529 (N_5529,N_3735,N_3339);
xnor U5530 (N_5530,N_4100,N_4189);
and U5531 (N_5531,N_3610,N_3598);
nor U5532 (N_5532,N_4249,N_3681);
nor U5533 (N_5533,N_4498,N_3539);
xor U5534 (N_5534,N_3312,N_4244);
nand U5535 (N_5535,N_4068,N_3078);
nor U5536 (N_5536,N_3692,N_3999);
and U5537 (N_5537,N_4052,N_3067);
and U5538 (N_5538,N_4462,N_3577);
xnor U5539 (N_5539,N_4271,N_4461);
and U5540 (N_5540,N_3765,N_3541);
or U5541 (N_5541,N_4002,N_3339);
nand U5542 (N_5542,N_3466,N_4202);
nand U5543 (N_5543,N_3171,N_3659);
nand U5544 (N_5544,N_4027,N_4419);
xor U5545 (N_5545,N_3898,N_4411);
and U5546 (N_5546,N_3039,N_4110);
or U5547 (N_5547,N_3399,N_3029);
or U5548 (N_5548,N_3372,N_3496);
nand U5549 (N_5549,N_3982,N_3794);
or U5550 (N_5550,N_3747,N_3910);
xnor U5551 (N_5551,N_3659,N_3849);
nand U5552 (N_5552,N_4107,N_4432);
and U5553 (N_5553,N_4268,N_3398);
nand U5554 (N_5554,N_3782,N_3881);
nor U5555 (N_5555,N_3609,N_4157);
xor U5556 (N_5556,N_3065,N_4252);
or U5557 (N_5557,N_3539,N_4291);
nand U5558 (N_5558,N_4386,N_4165);
nand U5559 (N_5559,N_3192,N_4232);
xnor U5560 (N_5560,N_3091,N_3049);
or U5561 (N_5561,N_3150,N_4445);
nor U5562 (N_5562,N_3757,N_3556);
xor U5563 (N_5563,N_3621,N_4314);
or U5564 (N_5564,N_3188,N_3950);
and U5565 (N_5565,N_3101,N_3107);
or U5566 (N_5566,N_3513,N_4239);
or U5567 (N_5567,N_3275,N_3628);
and U5568 (N_5568,N_3178,N_3271);
nand U5569 (N_5569,N_3443,N_4042);
or U5570 (N_5570,N_3985,N_3277);
nand U5571 (N_5571,N_4361,N_3036);
nor U5572 (N_5572,N_3797,N_3113);
nor U5573 (N_5573,N_3420,N_3303);
and U5574 (N_5574,N_3836,N_3959);
and U5575 (N_5575,N_4374,N_3694);
xor U5576 (N_5576,N_3464,N_3838);
or U5577 (N_5577,N_4124,N_4030);
nor U5578 (N_5578,N_3144,N_3141);
or U5579 (N_5579,N_3175,N_3258);
nor U5580 (N_5580,N_3852,N_3772);
nand U5581 (N_5581,N_3391,N_3765);
nor U5582 (N_5582,N_4366,N_3919);
or U5583 (N_5583,N_3305,N_4143);
nand U5584 (N_5584,N_3528,N_3490);
nor U5585 (N_5585,N_3346,N_3973);
xor U5586 (N_5586,N_3071,N_3475);
nor U5587 (N_5587,N_4397,N_4294);
nand U5588 (N_5588,N_3771,N_3840);
and U5589 (N_5589,N_3127,N_3021);
xnor U5590 (N_5590,N_3092,N_3559);
nand U5591 (N_5591,N_3369,N_3736);
xor U5592 (N_5592,N_3336,N_3272);
nor U5593 (N_5593,N_3747,N_4173);
nor U5594 (N_5594,N_3491,N_3290);
xnor U5595 (N_5595,N_3695,N_3077);
or U5596 (N_5596,N_3303,N_4396);
xor U5597 (N_5597,N_4404,N_4339);
nand U5598 (N_5598,N_4158,N_3178);
nor U5599 (N_5599,N_4455,N_3659);
nor U5600 (N_5600,N_4250,N_3703);
or U5601 (N_5601,N_4285,N_3860);
or U5602 (N_5602,N_4120,N_3484);
nand U5603 (N_5603,N_4268,N_3547);
and U5604 (N_5604,N_4063,N_4332);
and U5605 (N_5605,N_3094,N_4318);
or U5606 (N_5606,N_3668,N_3080);
nor U5607 (N_5607,N_3655,N_3618);
or U5608 (N_5608,N_3318,N_3270);
nor U5609 (N_5609,N_3386,N_4220);
nor U5610 (N_5610,N_3246,N_3223);
nor U5611 (N_5611,N_3615,N_3997);
or U5612 (N_5612,N_3803,N_3765);
or U5613 (N_5613,N_3629,N_3308);
nand U5614 (N_5614,N_3656,N_3929);
or U5615 (N_5615,N_3176,N_3013);
nor U5616 (N_5616,N_3700,N_3896);
or U5617 (N_5617,N_4019,N_4110);
xnor U5618 (N_5618,N_3226,N_3190);
nand U5619 (N_5619,N_4439,N_3801);
nand U5620 (N_5620,N_3448,N_3336);
nand U5621 (N_5621,N_4139,N_3942);
or U5622 (N_5622,N_4190,N_4031);
nand U5623 (N_5623,N_4184,N_3928);
or U5624 (N_5624,N_4272,N_3702);
and U5625 (N_5625,N_3991,N_4138);
xor U5626 (N_5626,N_3713,N_3911);
and U5627 (N_5627,N_4361,N_3073);
xnor U5628 (N_5628,N_4132,N_3383);
nor U5629 (N_5629,N_3729,N_3864);
or U5630 (N_5630,N_3822,N_3571);
or U5631 (N_5631,N_4356,N_3137);
and U5632 (N_5632,N_3244,N_3892);
and U5633 (N_5633,N_3895,N_3346);
and U5634 (N_5634,N_4036,N_3490);
and U5635 (N_5635,N_4125,N_3265);
nand U5636 (N_5636,N_4387,N_3457);
nand U5637 (N_5637,N_3504,N_3006);
or U5638 (N_5638,N_3515,N_3664);
nand U5639 (N_5639,N_3192,N_3734);
nand U5640 (N_5640,N_4342,N_3800);
xnor U5641 (N_5641,N_4270,N_4020);
and U5642 (N_5642,N_3756,N_4383);
or U5643 (N_5643,N_4398,N_3597);
or U5644 (N_5644,N_4460,N_3262);
xnor U5645 (N_5645,N_4370,N_3069);
and U5646 (N_5646,N_3555,N_4097);
nand U5647 (N_5647,N_3641,N_4105);
nor U5648 (N_5648,N_3445,N_3673);
xor U5649 (N_5649,N_3909,N_3575);
or U5650 (N_5650,N_4398,N_3721);
or U5651 (N_5651,N_3878,N_3526);
nor U5652 (N_5652,N_4108,N_4057);
xor U5653 (N_5653,N_3338,N_4155);
nand U5654 (N_5654,N_3883,N_3311);
nor U5655 (N_5655,N_4428,N_3042);
nor U5656 (N_5656,N_4367,N_4086);
or U5657 (N_5657,N_4345,N_3072);
and U5658 (N_5658,N_3562,N_3962);
xor U5659 (N_5659,N_3402,N_3445);
nor U5660 (N_5660,N_4071,N_4285);
xor U5661 (N_5661,N_3976,N_3817);
or U5662 (N_5662,N_3174,N_3499);
or U5663 (N_5663,N_4150,N_3441);
and U5664 (N_5664,N_3724,N_3266);
nand U5665 (N_5665,N_3091,N_4392);
nor U5666 (N_5666,N_3823,N_3014);
and U5667 (N_5667,N_3556,N_3500);
or U5668 (N_5668,N_4392,N_3697);
xnor U5669 (N_5669,N_4348,N_3633);
nor U5670 (N_5670,N_3571,N_3485);
and U5671 (N_5671,N_4426,N_3268);
nand U5672 (N_5672,N_3366,N_3819);
xnor U5673 (N_5673,N_4010,N_3699);
nand U5674 (N_5674,N_4372,N_4030);
xor U5675 (N_5675,N_3492,N_3620);
nor U5676 (N_5676,N_4073,N_3071);
and U5677 (N_5677,N_3395,N_4398);
or U5678 (N_5678,N_4000,N_3207);
xor U5679 (N_5679,N_3254,N_3337);
xor U5680 (N_5680,N_4332,N_3423);
nor U5681 (N_5681,N_4118,N_4324);
and U5682 (N_5682,N_3131,N_3073);
and U5683 (N_5683,N_3756,N_3677);
xnor U5684 (N_5684,N_3826,N_3008);
xnor U5685 (N_5685,N_3606,N_4276);
xor U5686 (N_5686,N_3574,N_3085);
nor U5687 (N_5687,N_4267,N_3833);
xnor U5688 (N_5688,N_3083,N_3206);
and U5689 (N_5689,N_3375,N_4384);
nand U5690 (N_5690,N_4261,N_4027);
or U5691 (N_5691,N_3774,N_3083);
or U5692 (N_5692,N_4322,N_3669);
or U5693 (N_5693,N_3653,N_3314);
xor U5694 (N_5694,N_3767,N_3081);
and U5695 (N_5695,N_3768,N_4203);
xnor U5696 (N_5696,N_3730,N_4324);
nor U5697 (N_5697,N_3338,N_3747);
and U5698 (N_5698,N_3588,N_3400);
or U5699 (N_5699,N_3009,N_4133);
nand U5700 (N_5700,N_3781,N_3337);
xor U5701 (N_5701,N_3853,N_3669);
nand U5702 (N_5702,N_4034,N_3844);
xnor U5703 (N_5703,N_3374,N_3093);
nor U5704 (N_5704,N_4475,N_4227);
or U5705 (N_5705,N_3219,N_3619);
nand U5706 (N_5706,N_3805,N_3537);
xor U5707 (N_5707,N_4287,N_3469);
nand U5708 (N_5708,N_3291,N_3983);
and U5709 (N_5709,N_3924,N_4152);
and U5710 (N_5710,N_3545,N_3679);
and U5711 (N_5711,N_3578,N_4362);
nand U5712 (N_5712,N_3360,N_3297);
or U5713 (N_5713,N_3068,N_4030);
or U5714 (N_5714,N_3819,N_3210);
xor U5715 (N_5715,N_3177,N_3276);
or U5716 (N_5716,N_3637,N_3487);
and U5717 (N_5717,N_3407,N_4223);
nand U5718 (N_5718,N_3664,N_3799);
nand U5719 (N_5719,N_3393,N_3674);
and U5720 (N_5720,N_3773,N_3485);
nor U5721 (N_5721,N_3329,N_3577);
xor U5722 (N_5722,N_4132,N_3491);
or U5723 (N_5723,N_3549,N_3021);
nor U5724 (N_5724,N_3120,N_3977);
nor U5725 (N_5725,N_4460,N_3924);
or U5726 (N_5726,N_3244,N_3958);
and U5727 (N_5727,N_4041,N_4150);
or U5728 (N_5728,N_4329,N_3132);
xor U5729 (N_5729,N_3404,N_3096);
nand U5730 (N_5730,N_3555,N_3876);
xor U5731 (N_5731,N_3194,N_3976);
nand U5732 (N_5732,N_4429,N_3450);
nand U5733 (N_5733,N_3511,N_3551);
nor U5734 (N_5734,N_3599,N_4361);
xor U5735 (N_5735,N_3605,N_4368);
and U5736 (N_5736,N_4299,N_4105);
xnor U5737 (N_5737,N_3982,N_3650);
or U5738 (N_5738,N_4430,N_3635);
xnor U5739 (N_5739,N_3537,N_3107);
nor U5740 (N_5740,N_4093,N_3761);
nand U5741 (N_5741,N_3586,N_3322);
nand U5742 (N_5742,N_4102,N_4255);
nand U5743 (N_5743,N_4200,N_3593);
nor U5744 (N_5744,N_3847,N_3975);
or U5745 (N_5745,N_3960,N_3307);
or U5746 (N_5746,N_3141,N_4363);
xor U5747 (N_5747,N_3425,N_3151);
nor U5748 (N_5748,N_3554,N_3561);
and U5749 (N_5749,N_4422,N_4121);
xnor U5750 (N_5750,N_4037,N_3043);
nand U5751 (N_5751,N_4494,N_3027);
and U5752 (N_5752,N_3809,N_3841);
nand U5753 (N_5753,N_3060,N_3871);
and U5754 (N_5754,N_4237,N_4478);
or U5755 (N_5755,N_3433,N_4316);
nor U5756 (N_5756,N_4491,N_4099);
nand U5757 (N_5757,N_3615,N_3494);
or U5758 (N_5758,N_3054,N_3486);
nand U5759 (N_5759,N_4324,N_4174);
and U5760 (N_5760,N_3199,N_4102);
or U5761 (N_5761,N_3428,N_3129);
or U5762 (N_5762,N_3313,N_3638);
nand U5763 (N_5763,N_3138,N_4193);
nor U5764 (N_5764,N_4239,N_4447);
and U5765 (N_5765,N_3229,N_3925);
and U5766 (N_5766,N_3808,N_4160);
and U5767 (N_5767,N_4458,N_3533);
nor U5768 (N_5768,N_4416,N_3204);
nand U5769 (N_5769,N_4071,N_3156);
or U5770 (N_5770,N_3603,N_3833);
nand U5771 (N_5771,N_3167,N_3222);
nand U5772 (N_5772,N_3691,N_3547);
and U5773 (N_5773,N_4109,N_4181);
and U5774 (N_5774,N_4250,N_3566);
or U5775 (N_5775,N_4004,N_3658);
nor U5776 (N_5776,N_3383,N_4425);
nor U5777 (N_5777,N_3589,N_3039);
nand U5778 (N_5778,N_3102,N_3176);
or U5779 (N_5779,N_4202,N_4460);
xor U5780 (N_5780,N_3001,N_4310);
xnor U5781 (N_5781,N_3417,N_3639);
and U5782 (N_5782,N_3726,N_4223);
nor U5783 (N_5783,N_4487,N_3155);
xnor U5784 (N_5784,N_4009,N_4207);
and U5785 (N_5785,N_4435,N_3285);
and U5786 (N_5786,N_3854,N_3491);
nor U5787 (N_5787,N_4273,N_3984);
or U5788 (N_5788,N_4379,N_3844);
nand U5789 (N_5789,N_3817,N_3424);
nand U5790 (N_5790,N_3908,N_3476);
nand U5791 (N_5791,N_4247,N_4025);
and U5792 (N_5792,N_3220,N_3045);
or U5793 (N_5793,N_3218,N_3733);
or U5794 (N_5794,N_3184,N_3527);
xnor U5795 (N_5795,N_3248,N_4216);
nand U5796 (N_5796,N_3106,N_4263);
nand U5797 (N_5797,N_3417,N_3662);
nand U5798 (N_5798,N_3939,N_3065);
and U5799 (N_5799,N_3426,N_4327);
nand U5800 (N_5800,N_4104,N_3583);
or U5801 (N_5801,N_3565,N_3641);
nand U5802 (N_5802,N_4311,N_4414);
nor U5803 (N_5803,N_3701,N_4382);
xor U5804 (N_5804,N_3232,N_3236);
or U5805 (N_5805,N_3508,N_4390);
and U5806 (N_5806,N_3924,N_3391);
xnor U5807 (N_5807,N_4123,N_3324);
and U5808 (N_5808,N_3143,N_4427);
nor U5809 (N_5809,N_4380,N_3046);
xnor U5810 (N_5810,N_3119,N_3452);
or U5811 (N_5811,N_4365,N_3183);
and U5812 (N_5812,N_4068,N_4385);
nand U5813 (N_5813,N_3936,N_3673);
xor U5814 (N_5814,N_3302,N_3885);
xor U5815 (N_5815,N_3655,N_4275);
nor U5816 (N_5816,N_3472,N_3323);
nand U5817 (N_5817,N_3846,N_3964);
nand U5818 (N_5818,N_3945,N_3952);
xnor U5819 (N_5819,N_3037,N_3712);
nand U5820 (N_5820,N_4468,N_3779);
and U5821 (N_5821,N_4230,N_3062);
xnor U5822 (N_5822,N_3873,N_3364);
and U5823 (N_5823,N_3534,N_3372);
xnor U5824 (N_5824,N_3635,N_3335);
or U5825 (N_5825,N_4300,N_4123);
xor U5826 (N_5826,N_3246,N_4335);
xor U5827 (N_5827,N_4164,N_3803);
or U5828 (N_5828,N_4450,N_3639);
nor U5829 (N_5829,N_4474,N_3400);
xnor U5830 (N_5830,N_3033,N_3079);
or U5831 (N_5831,N_3569,N_3335);
or U5832 (N_5832,N_4233,N_3279);
xnor U5833 (N_5833,N_3648,N_4014);
xor U5834 (N_5834,N_3826,N_3248);
nor U5835 (N_5835,N_3598,N_3423);
nor U5836 (N_5836,N_3319,N_3529);
or U5837 (N_5837,N_3617,N_3688);
nor U5838 (N_5838,N_3795,N_3917);
or U5839 (N_5839,N_4414,N_4454);
nor U5840 (N_5840,N_3323,N_3932);
and U5841 (N_5841,N_3587,N_4408);
xor U5842 (N_5842,N_4480,N_3859);
and U5843 (N_5843,N_3710,N_3436);
xnor U5844 (N_5844,N_3425,N_3011);
and U5845 (N_5845,N_4183,N_3984);
or U5846 (N_5846,N_4167,N_3702);
nor U5847 (N_5847,N_3737,N_4290);
or U5848 (N_5848,N_3392,N_3987);
or U5849 (N_5849,N_3885,N_3237);
nor U5850 (N_5850,N_3023,N_4373);
xnor U5851 (N_5851,N_4050,N_3629);
xor U5852 (N_5852,N_4159,N_4147);
or U5853 (N_5853,N_3310,N_3595);
or U5854 (N_5854,N_4042,N_3637);
nor U5855 (N_5855,N_3723,N_4353);
nor U5856 (N_5856,N_3426,N_3607);
and U5857 (N_5857,N_3622,N_3478);
nor U5858 (N_5858,N_3633,N_3465);
and U5859 (N_5859,N_3905,N_3825);
xor U5860 (N_5860,N_3121,N_4169);
and U5861 (N_5861,N_3152,N_3057);
and U5862 (N_5862,N_3687,N_4460);
nor U5863 (N_5863,N_3948,N_3403);
xnor U5864 (N_5864,N_3898,N_4376);
nand U5865 (N_5865,N_3719,N_3240);
and U5866 (N_5866,N_3262,N_3677);
or U5867 (N_5867,N_4195,N_4087);
and U5868 (N_5868,N_3824,N_3437);
and U5869 (N_5869,N_4090,N_4423);
nand U5870 (N_5870,N_4016,N_3585);
xnor U5871 (N_5871,N_3444,N_4490);
nor U5872 (N_5872,N_4313,N_3128);
nand U5873 (N_5873,N_3506,N_3034);
and U5874 (N_5874,N_3072,N_3508);
xnor U5875 (N_5875,N_4347,N_3173);
nand U5876 (N_5876,N_3059,N_4436);
nor U5877 (N_5877,N_4091,N_3271);
and U5878 (N_5878,N_3885,N_3048);
nand U5879 (N_5879,N_3671,N_3936);
nand U5880 (N_5880,N_3551,N_4130);
xnor U5881 (N_5881,N_4434,N_4494);
or U5882 (N_5882,N_3166,N_4347);
and U5883 (N_5883,N_3538,N_4267);
nor U5884 (N_5884,N_4182,N_3063);
and U5885 (N_5885,N_3073,N_3469);
and U5886 (N_5886,N_3535,N_4402);
and U5887 (N_5887,N_4448,N_3063);
and U5888 (N_5888,N_3241,N_3070);
xor U5889 (N_5889,N_4302,N_3460);
xnor U5890 (N_5890,N_3856,N_3165);
nor U5891 (N_5891,N_3064,N_4429);
nand U5892 (N_5892,N_3723,N_3205);
nand U5893 (N_5893,N_3981,N_3388);
nand U5894 (N_5894,N_3643,N_3208);
nand U5895 (N_5895,N_4415,N_3808);
and U5896 (N_5896,N_4046,N_3239);
and U5897 (N_5897,N_4160,N_3308);
xnor U5898 (N_5898,N_4075,N_4090);
or U5899 (N_5899,N_3462,N_3032);
and U5900 (N_5900,N_3114,N_3110);
nor U5901 (N_5901,N_3929,N_3841);
or U5902 (N_5902,N_3893,N_3201);
xor U5903 (N_5903,N_3095,N_3132);
or U5904 (N_5904,N_3669,N_3664);
nand U5905 (N_5905,N_4241,N_3018);
nor U5906 (N_5906,N_3602,N_3327);
xnor U5907 (N_5907,N_3797,N_3903);
nand U5908 (N_5908,N_3528,N_3538);
and U5909 (N_5909,N_4023,N_3568);
xor U5910 (N_5910,N_3180,N_3737);
nand U5911 (N_5911,N_3999,N_3332);
nor U5912 (N_5912,N_4455,N_4330);
nand U5913 (N_5913,N_4110,N_3734);
and U5914 (N_5914,N_3375,N_3179);
nand U5915 (N_5915,N_3000,N_3559);
nand U5916 (N_5916,N_4171,N_3555);
xnor U5917 (N_5917,N_3164,N_3212);
and U5918 (N_5918,N_4094,N_3061);
xnor U5919 (N_5919,N_3890,N_3159);
xor U5920 (N_5920,N_3128,N_4432);
nand U5921 (N_5921,N_3611,N_3744);
nor U5922 (N_5922,N_4043,N_4306);
nor U5923 (N_5923,N_3751,N_3696);
xor U5924 (N_5924,N_4494,N_3268);
or U5925 (N_5925,N_3307,N_3661);
and U5926 (N_5926,N_3212,N_4290);
or U5927 (N_5927,N_3838,N_3044);
and U5928 (N_5928,N_3786,N_3602);
nand U5929 (N_5929,N_3442,N_3451);
nand U5930 (N_5930,N_4371,N_3941);
and U5931 (N_5931,N_4439,N_3188);
nor U5932 (N_5932,N_4403,N_4492);
and U5933 (N_5933,N_3810,N_4053);
nand U5934 (N_5934,N_4307,N_3741);
xnor U5935 (N_5935,N_4475,N_4153);
and U5936 (N_5936,N_3152,N_4075);
xor U5937 (N_5937,N_3284,N_3070);
xnor U5938 (N_5938,N_4148,N_3404);
or U5939 (N_5939,N_3836,N_4321);
and U5940 (N_5940,N_4291,N_3802);
and U5941 (N_5941,N_3174,N_3960);
or U5942 (N_5942,N_3955,N_3732);
nand U5943 (N_5943,N_4346,N_4427);
or U5944 (N_5944,N_4348,N_3488);
or U5945 (N_5945,N_3501,N_3983);
nor U5946 (N_5946,N_4054,N_3467);
and U5947 (N_5947,N_3937,N_4479);
and U5948 (N_5948,N_3952,N_3252);
xnor U5949 (N_5949,N_3548,N_3415);
and U5950 (N_5950,N_4156,N_3734);
nand U5951 (N_5951,N_3764,N_4041);
xor U5952 (N_5952,N_4072,N_3190);
and U5953 (N_5953,N_4042,N_3596);
or U5954 (N_5954,N_3098,N_4353);
nand U5955 (N_5955,N_3896,N_4255);
xor U5956 (N_5956,N_3460,N_3159);
nand U5957 (N_5957,N_4287,N_4480);
and U5958 (N_5958,N_3784,N_3224);
nor U5959 (N_5959,N_4310,N_3752);
xnor U5960 (N_5960,N_3723,N_3523);
and U5961 (N_5961,N_3623,N_3014);
nor U5962 (N_5962,N_3686,N_3723);
and U5963 (N_5963,N_3449,N_3819);
nand U5964 (N_5964,N_3953,N_3423);
nor U5965 (N_5965,N_4447,N_4410);
and U5966 (N_5966,N_3845,N_3010);
and U5967 (N_5967,N_3811,N_3215);
nor U5968 (N_5968,N_3978,N_3469);
xnor U5969 (N_5969,N_4331,N_3773);
and U5970 (N_5970,N_3262,N_4198);
or U5971 (N_5971,N_3209,N_3364);
nor U5972 (N_5972,N_3848,N_3238);
or U5973 (N_5973,N_4281,N_3020);
nand U5974 (N_5974,N_4058,N_4437);
nor U5975 (N_5975,N_3702,N_3528);
nand U5976 (N_5976,N_3843,N_3489);
nor U5977 (N_5977,N_3829,N_3831);
and U5978 (N_5978,N_3994,N_3642);
or U5979 (N_5979,N_3393,N_3614);
nor U5980 (N_5980,N_3670,N_4286);
nand U5981 (N_5981,N_3929,N_3189);
nor U5982 (N_5982,N_3294,N_3818);
xnor U5983 (N_5983,N_3027,N_4339);
xor U5984 (N_5984,N_3088,N_3525);
xor U5985 (N_5985,N_3596,N_3173);
nor U5986 (N_5986,N_4243,N_3173);
or U5987 (N_5987,N_3008,N_3617);
and U5988 (N_5988,N_3174,N_4157);
nand U5989 (N_5989,N_4139,N_3548);
xnor U5990 (N_5990,N_4432,N_4266);
or U5991 (N_5991,N_4251,N_4390);
or U5992 (N_5992,N_3746,N_3652);
nand U5993 (N_5993,N_3210,N_3224);
xnor U5994 (N_5994,N_3461,N_3060);
nor U5995 (N_5995,N_3424,N_3742);
nand U5996 (N_5996,N_3826,N_3580);
nor U5997 (N_5997,N_3725,N_3670);
nand U5998 (N_5998,N_4037,N_4359);
nand U5999 (N_5999,N_3672,N_3113);
xnor U6000 (N_6000,N_4972,N_5387);
or U6001 (N_6001,N_4961,N_5269);
and U6002 (N_6002,N_5954,N_5612);
or U6003 (N_6003,N_5799,N_5152);
and U6004 (N_6004,N_4545,N_5800);
xnor U6005 (N_6005,N_5015,N_5082);
xor U6006 (N_6006,N_4600,N_5434);
nand U6007 (N_6007,N_5094,N_5348);
or U6008 (N_6008,N_5945,N_5325);
xor U6009 (N_6009,N_4875,N_4797);
and U6010 (N_6010,N_5130,N_5250);
and U6011 (N_6011,N_5390,N_5077);
xnor U6012 (N_6012,N_5406,N_4978);
nor U6013 (N_6013,N_4669,N_5843);
or U6014 (N_6014,N_5416,N_5714);
and U6015 (N_6015,N_5597,N_5711);
and U6016 (N_6016,N_5389,N_4940);
nor U6017 (N_6017,N_5541,N_5080);
nand U6018 (N_6018,N_5057,N_5039);
or U6019 (N_6019,N_5972,N_5992);
xnor U6020 (N_6020,N_4680,N_4926);
or U6021 (N_6021,N_5645,N_5575);
nand U6022 (N_6022,N_5884,N_5153);
or U6023 (N_6023,N_5326,N_4790);
xor U6024 (N_6024,N_4862,N_5088);
and U6025 (N_6025,N_5161,N_5116);
nor U6026 (N_6026,N_5079,N_5043);
or U6027 (N_6027,N_5812,N_4566);
xor U6028 (N_6028,N_5727,N_5143);
nor U6029 (N_6029,N_5038,N_4911);
xnor U6030 (N_6030,N_5911,N_5070);
or U6031 (N_6031,N_4995,N_5500);
nand U6032 (N_6032,N_5748,N_5343);
nor U6033 (N_6033,N_5223,N_5523);
nand U6034 (N_6034,N_5525,N_5664);
and U6035 (N_6035,N_4732,N_5486);
nand U6036 (N_6036,N_4725,N_5732);
nor U6037 (N_6037,N_4733,N_5696);
nand U6038 (N_6038,N_5805,N_5508);
nor U6039 (N_6039,N_4603,N_4795);
nand U6040 (N_6040,N_4611,N_5624);
and U6041 (N_6041,N_5505,N_5410);
xor U6042 (N_6042,N_5674,N_4738);
xnor U6043 (N_6043,N_5731,N_5767);
nand U6044 (N_6044,N_4787,N_5988);
nand U6045 (N_6045,N_5692,N_5099);
or U6046 (N_6046,N_5121,N_4977);
or U6047 (N_6047,N_4974,N_5234);
xnor U6048 (N_6048,N_4840,N_5435);
or U6049 (N_6049,N_5687,N_5602);
and U6050 (N_6050,N_4864,N_5912);
xor U6051 (N_6051,N_5189,N_5056);
and U6052 (N_6052,N_5149,N_5471);
nor U6053 (N_6053,N_5574,N_5160);
or U6054 (N_6054,N_4737,N_5942);
and U6055 (N_6055,N_4768,N_5529);
nand U6056 (N_6056,N_5478,N_5933);
nand U6057 (N_6057,N_5623,N_4934);
nor U6058 (N_6058,N_5924,N_5689);
and U6059 (N_6059,N_5848,N_5607);
nor U6060 (N_6060,N_5216,N_5637);
or U6061 (N_6061,N_4676,N_4783);
nand U6062 (N_6062,N_5572,N_5991);
or U6063 (N_6063,N_5789,N_4728);
nand U6064 (N_6064,N_5111,N_5853);
nor U6065 (N_6065,N_5051,N_5439);
and U6066 (N_6066,N_5141,N_4947);
and U6067 (N_6067,N_5401,N_5846);
or U6068 (N_6068,N_5113,N_5700);
nand U6069 (N_6069,N_5419,N_4785);
and U6070 (N_6070,N_5156,N_4571);
xnor U6071 (N_6071,N_5304,N_4624);
nand U6072 (N_6072,N_5879,N_5022);
nand U6073 (N_6073,N_4670,N_5453);
nand U6074 (N_6074,N_5786,N_4547);
nor U6075 (N_6075,N_4501,N_5313);
or U6076 (N_6076,N_5816,N_4761);
xnor U6077 (N_6077,N_5829,N_5772);
or U6078 (N_6078,N_4520,N_5227);
or U6079 (N_6079,N_4516,N_5517);
nor U6080 (N_6080,N_4660,N_5703);
nand U6081 (N_6081,N_4636,N_4546);
xor U6082 (N_6082,N_5134,N_5368);
or U6083 (N_6083,N_5440,N_5429);
nor U6084 (N_6084,N_5995,N_5621);
and U6085 (N_6085,N_5259,N_5707);
nor U6086 (N_6086,N_4922,N_5260);
xor U6087 (N_6087,N_4549,N_5813);
xnor U6088 (N_6088,N_4641,N_5793);
xor U6089 (N_6089,N_5874,N_4562);
xor U6090 (N_6090,N_5796,N_5809);
or U6091 (N_6091,N_5142,N_5751);
xnor U6092 (N_6092,N_5824,N_5132);
xnor U6093 (N_6093,N_4541,N_5679);
nor U6094 (N_6094,N_5923,N_5502);
xnor U6095 (N_6095,N_4882,N_5490);
nor U6096 (N_6096,N_4585,N_5203);
and U6097 (N_6097,N_5430,N_5136);
nor U6098 (N_6098,N_5006,N_5339);
or U6099 (N_6099,N_5656,N_5641);
nand U6100 (N_6100,N_5828,N_5610);
and U6101 (N_6101,N_5107,N_5364);
or U6102 (N_6102,N_5449,N_5588);
nor U6103 (N_6103,N_4906,N_5078);
and U6104 (N_6104,N_5405,N_5702);
and U6105 (N_6105,N_5569,N_5729);
nor U6106 (N_6106,N_5555,N_5404);
nor U6107 (N_6107,N_4834,N_5652);
or U6108 (N_6108,N_4716,N_5521);
nor U6109 (N_6109,N_5474,N_5739);
nor U6110 (N_6110,N_5243,N_5801);
nand U6111 (N_6111,N_4534,N_4808);
nor U6112 (N_6112,N_4807,N_4957);
xnor U6113 (N_6113,N_4837,N_5802);
nand U6114 (N_6114,N_4710,N_4945);
nor U6115 (N_6115,N_4689,N_4750);
xor U6116 (N_6116,N_5720,N_5929);
nand U6117 (N_6117,N_4765,N_5367);
and U6118 (N_6118,N_5891,N_5682);
xnor U6119 (N_6119,N_4586,N_5522);
nor U6120 (N_6120,N_5681,N_5821);
or U6121 (N_6121,N_4967,N_5164);
nor U6122 (N_6122,N_5927,N_5790);
nor U6123 (N_6123,N_5938,N_5425);
nand U6124 (N_6124,N_5279,N_4522);
nand U6125 (N_6125,N_5514,N_4561);
nand U6126 (N_6126,N_5902,N_4905);
nor U6127 (N_6127,N_5354,N_5908);
nor U6128 (N_6128,N_5571,N_4671);
and U6129 (N_6129,N_4576,N_5007);
nand U6130 (N_6130,N_4986,N_5218);
and U6131 (N_6131,N_5620,N_5186);
xnor U6132 (N_6132,N_5581,N_5297);
and U6133 (N_6133,N_5150,N_5915);
or U6134 (N_6134,N_4705,N_5666);
nor U6135 (N_6135,N_5715,N_5788);
or U6136 (N_6136,N_5646,N_5940);
and U6137 (N_6137,N_5998,N_4741);
nand U6138 (N_6138,N_4568,N_5724);
xor U6139 (N_6139,N_5746,N_5540);
or U6140 (N_6140,N_5123,N_5168);
nand U6141 (N_6141,N_5213,N_5358);
and U6142 (N_6142,N_5899,N_5454);
nand U6143 (N_6143,N_5889,N_5823);
or U6144 (N_6144,N_4865,N_5159);
xor U6145 (N_6145,N_4814,N_5238);
nand U6146 (N_6146,N_5320,N_5677);
nor U6147 (N_6147,N_4613,N_5324);
nand U6148 (N_6148,N_4718,N_4779);
and U6149 (N_6149,N_4928,N_5614);
or U6150 (N_6150,N_5378,N_5437);
or U6151 (N_6151,N_5349,N_5591);
or U6152 (N_6152,N_4572,N_4570);
and U6153 (N_6153,N_5599,N_5660);
xnor U6154 (N_6154,N_5869,N_4848);
and U6155 (N_6155,N_4871,N_5895);
nor U6156 (N_6156,N_5920,N_4850);
or U6157 (N_6157,N_5593,N_5496);
nor U6158 (N_6158,N_5157,N_4577);
xor U6159 (N_6159,N_5594,N_5752);
nand U6160 (N_6160,N_5922,N_5173);
nand U6161 (N_6161,N_4592,N_4747);
or U6162 (N_6162,N_5021,N_4910);
or U6163 (N_6163,N_4616,N_4633);
nor U6164 (N_6164,N_5636,N_5340);
xor U6165 (N_6165,N_4798,N_4897);
nor U6166 (N_6166,N_4548,N_5273);
xor U6167 (N_6167,N_4748,N_5308);
and U6168 (N_6168,N_5873,N_5040);
or U6169 (N_6169,N_5488,N_5432);
or U6170 (N_6170,N_5334,N_5838);
xor U6171 (N_6171,N_5859,N_5402);
xor U6172 (N_6172,N_4884,N_4764);
xor U6173 (N_6173,N_5462,N_5976);
xnor U6174 (N_6174,N_4951,N_5797);
xor U6175 (N_6175,N_5546,N_4885);
nor U6176 (N_6176,N_4615,N_5756);
nor U6177 (N_6177,N_5093,N_4744);
xor U6178 (N_6178,N_5341,N_5830);
xnor U6179 (N_6179,N_4789,N_5543);
and U6180 (N_6180,N_5253,N_5204);
nand U6181 (N_6181,N_5780,N_5625);
nor U6182 (N_6182,N_5698,N_5630);
or U6183 (N_6183,N_5026,N_5971);
nor U6184 (N_6184,N_5303,N_5667);
and U6185 (N_6185,N_5196,N_5925);
nor U6186 (N_6186,N_5563,N_5394);
nand U6187 (N_6187,N_4659,N_4608);
nand U6188 (N_6188,N_5857,N_4819);
and U6189 (N_6189,N_4507,N_5145);
xor U6190 (N_6190,N_4550,N_5561);
xor U6191 (N_6191,N_5570,N_5850);
and U6192 (N_6192,N_5046,N_4551);
or U6193 (N_6193,N_5955,N_5818);
nor U6194 (N_6194,N_4734,N_5956);
or U6195 (N_6195,N_4628,N_4722);
or U6196 (N_6196,N_5803,N_4573);
or U6197 (N_6197,N_5315,N_5842);
xnor U6198 (N_6198,N_5559,N_4695);
and U6199 (N_6199,N_5952,N_5301);
xor U6200 (N_6200,N_4890,N_4821);
nor U6201 (N_6201,N_4902,N_5014);
xor U6202 (N_6202,N_4588,N_5373);
nand U6203 (N_6203,N_5312,N_4575);
xor U6204 (N_6204,N_5158,N_4504);
nor U6205 (N_6205,N_4932,N_4899);
nor U6206 (N_6206,N_5458,N_4966);
xnor U6207 (N_6207,N_5648,N_4620);
or U6208 (N_6208,N_5444,N_4715);
xnor U6209 (N_6209,N_5059,N_5697);
and U6210 (N_6210,N_5680,N_5959);
nand U6211 (N_6211,N_4740,N_5208);
xor U6212 (N_6212,N_5639,N_5877);
nor U6213 (N_6213,N_4930,N_5065);
or U6214 (N_6214,N_4532,N_4529);
or U6215 (N_6215,N_5485,N_4981);
nor U6216 (N_6216,N_5701,N_5629);
nor U6217 (N_6217,N_4753,N_4602);
xor U6218 (N_6218,N_4607,N_5735);
or U6219 (N_6219,N_5578,N_5197);
nand U6220 (N_6220,N_5119,N_4505);
xnor U6221 (N_6221,N_4860,N_5381);
nand U6222 (N_6222,N_5293,N_4599);
nand U6223 (N_6223,N_5221,N_4954);
nor U6224 (N_6224,N_5089,N_5982);
xor U6225 (N_6225,N_5214,N_4601);
nand U6226 (N_6226,N_4543,N_5684);
nand U6227 (N_6227,N_5131,N_5307);
xor U6228 (N_6228,N_5820,N_4915);
and U6229 (N_6229,N_4510,N_4762);
nor U6230 (N_6230,N_4556,N_5230);
nand U6231 (N_6231,N_4836,N_4810);
or U6232 (N_6232,N_5224,N_5110);
or U6233 (N_6233,N_5254,N_5470);
xor U6234 (N_6234,N_4665,N_4528);
nand U6235 (N_6235,N_5503,N_5615);
and U6236 (N_6236,N_5835,N_4874);
or U6237 (N_6237,N_5192,N_4852);
xnor U6238 (N_6238,N_4796,N_5222);
and U6239 (N_6239,N_4640,N_5861);
nand U6240 (N_6240,N_4959,N_4820);
and U6241 (N_6241,N_5583,N_4736);
xor U6242 (N_6242,N_5519,N_5935);
xnor U6243 (N_6243,N_5447,N_4584);
and U6244 (N_6244,N_5542,N_5274);
and U6245 (N_6245,N_4908,N_5286);
nor U6246 (N_6246,N_5108,N_4567);
and U6247 (N_6247,N_5815,N_5537);
and U6248 (N_6248,N_5734,N_4609);
nand U6249 (N_6249,N_4869,N_5034);
xor U6250 (N_6250,N_4826,N_4847);
and U6251 (N_6251,N_5296,N_5690);
and U6252 (N_6252,N_5551,N_5020);
nor U6253 (N_6253,N_5202,N_4720);
and U6254 (N_6254,N_5970,N_4500);
or U6255 (N_6255,N_5412,N_5577);
and U6256 (N_6256,N_5662,N_5005);
or U6257 (N_6257,N_5609,N_4679);
or U6258 (N_6258,N_5978,N_5601);
xor U6259 (N_6259,N_4707,N_4770);
or U6260 (N_6260,N_5509,N_5352);
xor U6261 (N_6261,N_5283,N_4540);
nor U6262 (N_6262,N_5008,N_5875);
xnor U6263 (N_6263,N_5833,N_5939);
nor U6264 (N_6264,N_5492,N_5380);
nor U6265 (N_6265,N_5067,N_5579);
and U6266 (N_6266,N_5672,N_5473);
and U6267 (N_6267,N_4698,N_4511);
or U6268 (N_6268,N_4666,N_5010);
xor U6269 (N_6269,N_4788,N_5530);
xor U6270 (N_6270,N_5356,N_4539);
and U6271 (N_6271,N_5212,N_5977);
and U6272 (N_6272,N_4996,N_4927);
and U6273 (N_6273,N_5331,N_5854);
nor U6274 (N_6274,N_4622,N_4948);
nor U6275 (N_6275,N_5305,N_5170);
nor U6276 (N_6276,N_5017,N_5178);
nand U6277 (N_6277,N_4929,N_5794);
or U6278 (N_6278,N_5573,N_5271);
xnor U6279 (N_6279,N_5582,N_4883);
nor U6280 (N_6280,N_5350,N_4590);
nor U6281 (N_6281,N_5346,N_4675);
or U6282 (N_6282,N_5135,N_5058);
nand U6283 (N_6283,N_5709,N_4827);
and U6284 (N_6284,N_4839,N_5480);
nor U6285 (N_6285,N_5181,N_5921);
xnor U6286 (N_6286,N_5712,N_4763);
xnor U6287 (N_6287,N_5872,N_5946);
xor U6288 (N_6288,N_4515,N_5795);
nand U6289 (N_6289,N_5916,N_5126);
nor U6290 (N_6290,N_4527,N_5475);
or U6291 (N_6291,N_4652,N_4802);
or U6292 (N_6292,N_4681,N_5806);
nand U6293 (N_6293,N_5535,N_4727);
or U6294 (N_6294,N_5631,N_4721);
or U6295 (N_6295,N_5392,N_4782);
nor U6296 (N_6296,N_5867,N_5659);
or U6297 (N_6297,N_5060,N_4843);
xnor U6298 (N_6298,N_5035,N_5695);
or U6299 (N_6299,N_4717,N_5759);
nor U6300 (N_6300,N_5688,N_5556);
and U6301 (N_6301,N_4773,N_5750);
and U6302 (N_6302,N_4587,N_4563);
nand U6303 (N_6303,N_5281,N_4994);
and U6304 (N_6304,N_4555,N_4754);
or U6305 (N_6305,N_4702,N_4969);
and U6306 (N_6306,N_4745,N_5966);
or U6307 (N_6307,N_5691,N_5771);
or U6308 (N_6308,N_4946,N_5120);
and U6309 (N_6309,N_5675,N_5310);
or U6310 (N_6310,N_5871,N_5194);
nor U6311 (N_6311,N_4888,N_5769);
and U6312 (N_6312,N_5122,N_5774);
and U6313 (N_6313,N_5256,N_4606);
nor U6314 (N_6314,N_5968,N_5219);
nor U6315 (N_6315,N_4661,N_5317);
nand U6316 (N_6316,N_5066,N_5747);
or U6317 (N_6317,N_5584,N_5836);
nand U6318 (N_6318,N_4687,N_5958);
nor U6319 (N_6319,N_4692,N_4596);
or U6320 (N_6320,N_5777,N_5494);
and U6321 (N_6321,N_4896,N_5600);
or U6322 (N_6322,N_5288,N_5635);
nand U6323 (N_6323,N_4593,N_5163);
xnor U6324 (N_6324,N_5520,N_5866);
nor U6325 (N_6325,N_4830,N_5029);
nor U6326 (N_6326,N_5883,N_4617);
and U6327 (N_6327,N_5424,N_5644);
and U6328 (N_6328,N_5754,N_5290);
nand U6329 (N_6329,N_5264,N_5975);
xor U6330 (N_6330,N_4825,N_5811);
nor U6331 (N_6331,N_4950,N_5332);
and U6332 (N_6332,N_5558,N_5863);
and U6333 (N_6333,N_4731,N_5385);
xnor U6334 (N_6334,N_4553,N_5154);
and U6335 (N_6335,N_4956,N_5353);
xor U6336 (N_6336,N_5784,N_5657);
and U6337 (N_6337,N_5397,N_5104);
nor U6338 (N_6338,N_4746,N_4723);
nor U6339 (N_6339,N_5504,N_4699);
and U6340 (N_6340,N_4815,N_5518);
or U6341 (N_6341,N_5513,N_5418);
and U6342 (N_6342,N_4993,N_5426);
nor U6343 (N_6343,N_5890,N_4856);
nor U6344 (N_6344,N_5239,N_5294);
and U6345 (N_6345,N_4935,N_5199);
or U6346 (N_6346,N_5845,N_4751);
xor U6347 (N_6347,N_5011,N_5248);
nor U6348 (N_6348,N_5284,N_5073);
nand U6349 (N_6349,N_5495,N_5903);
xnor U6350 (N_6350,N_5819,N_4667);
or U6351 (N_6351,N_5409,N_4623);
or U6352 (N_6352,N_5919,N_5235);
nand U6353 (N_6353,N_5300,N_5210);
or U6354 (N_6354,N_5960,N_4719);
or U6355 (N_6355,N_5344,N_4806);
nand U6356 (N_6356,N_4923,N_4892);
nor U6357 (N_6357,N_5399,N_5427);
xnor U6358 (N_6358,N_5002,N_5498);
nand U6359 (N_6359,N_4938,N_5943);
or U6360 (N_6360,N_5587,N_5654);
xnor U6361 (N_6361,N_4627,N_4980);
nor U6362 (N_6362,N_5783,N_5745);
xor U6363 (N_6363,N_5706,N_4708);
or U6364 (N_6364,N_4523,N_5233);
nor U6365 (N_6365,N_4900,N_5832);
or U6366 (N_6366,N_5598,N_4517);
nand U6367 (N_6367,N_5074,N_5362);
and U6368 (N_6368,N_5616,N_5888);
xor U6369 (N_6369,N_4794,N_5768);
and U6370 (N_6370,N_5831,N_4726);
or U6371 (N_6371,N_5576,N_5876);
or U6372 (N_6372,N_5245,N_5878);
nor U6373 (N_6373,N_5277,N_5862);
nor U6374 (N_6374,N_5351,N_4822);
and U6375 (N_6375,N_5463,N_5738);
nand U6376 (N_6376,N_5102,N_4878);
and U6377 (N_6377,N_5552,N_5808);
nand U6378 (N_6378,N_5180,N_5910);
and U6379 (N_6379,N_5740,N_4706);
nor U6380 (N_6380,N_4589,N_5511);
xnor U6381 (N_6381,N_5147,N_5936);
or U6382 (N_6382,N_5270,N_4629);
xnor U6383 (N_6383,N_4987,N_5329);
and U6384 (N_6384,N_5395,N_4503);
and U6385 (N_6385,N_5628,N_5860);
xor U6386 (N_6386,N_5568,N_5133);
and U6387 (N_6387,N_4735,N_4868);
nor U6388 (N_6388,N_5357,N_5001);
and U6389 (N_6389,N_4772,N_4914);
and U6390 (N_6390,N_5338,N_4824);
nand U6391 (N_6391,N_5531,N_5117);
and U6392 (N_6392,N_4776,N_4998);
and U6393 (N_6393,N_4912,N_5603);
nor U6394 (N_6394,N_5355,N_4913);
nand U6395 (N_6395,N_5403,N_5316);
and U6396 (N_6396,N_5491,N_4635);
and U6397 (N_6397,N_5191,N_4828);
and U6398 (N_6398,N_5981,N_5778);
nor U6399 (N_6399,N_5246,N_5366);
nand U6400 (N_6400,N_4943,N_4542);
xor U6401 (N_6401,N_5171,N_5129);
and U6402 (N_6402,N_5023,N_5414);
or U6403 (N_6403,N_5757,N_4618);
nand U6404 (N_6404,N_5251,N_4792);
nand U6405 (N_6405,N_5586,N_5330);
nand U6406 (N_6406,N_5012,N_5721);
nand U6407 (N_6407,N_5420,N_5244);
or U6408 (N_6408,N_5282,N_5032);
and U6409 (N_6409,N_5114,N_4637);
and U6410 (N_6410,N_4841,N_5328);
or U6411 (N_6411,N_5337,N_4835);
and U6412 (N_6412,N_5175,N_5725);
and U6413 (N_6413,N_4809,N_5941);
and U6414 (N_6414,N_4642,N_5263);
nand U6415 (N_6415,N_5595,N_5984);
nor U6416 (N_6416,N_4964,N_5318);
or U6417 (N_6417,N_5726,N_5839);
nand U6418 (N_6418,N_4559,N_5763);
nand U6419 (N_6419,N_5247,N_5327);
or U6420 (N_6420,N_5106,N_5188);
nand U6421 (N_6421,N_5323,N_5476);
and U6422 (N_6422,N_5590,N_5388);
xnor U6423 (N_6423,N_5261,N_5847);
xor U6424 (N_6424,N_5928,N_5536);
xnor U6425 (N_6425,N_5676,N_4614);
nand U6426 (N_6426,N_4953,N_5526);
nor U6427 (N_6427,N_5018,N_5278);
and U6428 (N_6428,N_4936,N_5417);
or U6429 (N_6429,N_5773,N_4887);
nor U6430 (N_6430,N_5661,N_4903);
and U6431 (N_6431,N_4743,N_5139);
and U6432 (N_6432,N_4508,N_5383);
nand U6433 (N_6433,N_5109,N_4801);
or U6434 (N_6434,N_5200,N_5456);
and U6435 (N_6435,N_5807,N_5045);
or U6436 (N_6436,N_4989,N_4849);
nor U6437 (N_6437,N_4638,N_4684);
and U6438 (N_6438,N_4859,N_5105);
nor U6439 (N_6439,N_4519,N_4895);
nor U6440 (N_6440,N_5280,N_5155);
and U6441 (N_6441,N_5604,N_5041);
or U6442 (N_6442,N_4767,N_5983);
and U6443 (N_6443,N_5232,N_5483);
and U6444 (N_6444,N_5792,N_5554);
xor U6445 (N_6445,N_5605,N_5560);
and U6446 (N_6446,N_4968,N_4983);
nand U6447 (N_6447,N_5413,N_5003);
or U6448 (N_6448,N_4604,N_4962);
and U6449 (N_6449,N_4851,N_5167);
nor U6450 (N_6450,N_5071,N_4774);
nor U6451 (N_6451,N_5377,N_5241);
xnor U6452 (N_6452,N_4757,N_5016);
or U6453 (N_6453,N_5716,N_5371);
nor U6454 (N_6454,N_5255,N_5363);
xnor U6455 (N_6455,N_5993,N_5997);
or U6456 (N_6456,N_4678,N_4893);
nor U6457 (N_6457,N_5081,N_4696);
or U6458 (N_6458,N_5042,N_5882);
or U6459 (N_6459,N_4949,N_5632);
xnor U6460 (N_6460,N_4846,N_5087);
nor U6461 (N_6461,N_5292,N_5913);
and U6462 (N_6462,N_5127,N_5969);
xnor U6463 (N_6463,N_5484,N_5013);
xnor U6464 (N_6464,N_5653,N_5892);
nand U6465 (N_6465,N_4955,N_5027);
or U6466 (N_6466,N_5804,N_5091);
or U6467 (N_6467,N_4526,N_4630);
nand U6468 (N_6468,N_5342,N_5708);
or U6469 (N_6469,N_4578,N_4521);
xor U6470 (N_6470,N_5258,N_5717);
and U6471 (N_6471,N_4530,N_4891);
and U6472 (N_6472,N_4771,N_5441);
nand U6473 (N_6473,N_5539,N_5407);
nand U6474 (N_6474,N_4742,N_5472);
xnor U6475 (N_6475,N_5528,N_5477);
or U6476 (N_6476,N_5393,N_5887);
nor U6477 (N_6477,N_5906,N_5973);
nor U6478 (N_6478,N_4778,N_4538);
and U6479 (N_6479,N_5704,N_4691);
nand U6480 (N_6480,N_5516,N_5633);
and U6481 (N_6481,N_4973,N_4714);
or U6482 (N_6482,N_4512,N_4688);
and U6483 (N_6483,N_4863,N_5766);
or U6484 (N_6484,N_5640,N_5461);
nor U6485 (N_6485,N_4756,N_4686);
nand U6486 (N_6486,N_5979,N_5791);
and U6487 (N_6487,N_5668,N_5146);
and U6488 (N_6488,N_4963,N_5761);
nor U6489 (N_6489,N_5673,N_5365);
or U6490 (N_6490,N_4876,N_4803);
xor U6491 (N_6491,N_4749,N_4625);
and U6492 (N_6492,N_5781,N_4781);
xnor U6493 (N_6493,N_5382,N_4775);
and U6494 (N_6494,N_4760,N_4514);
nand U6495 (N_6495,N_5693,N_4648);
and U6496 (N_6496,N_4867,N_4701);
nand U6497 (N_6497,N_5897,N_5787);
nor U6498 (N_6498,N_5827,N_5686);
xor U6499 (N_6499,N_5465,N_5162);
nand U6500 (N_6500,N_4813,N_4937);
nor U6501 (N_6501,N_5231,N_5459);
or U6502 (N_6502,N_5987,N_5050);
xnor U6503 (N_6503,N_5479,N_4597);
and U6504 (N_6504,N_5347,N_5295);
nand U6505 (N_6505,N_4988,N_4557);
nand U6506 (N_6506,N_5374,N_5229);
and U6507 (N_6507,N_5125,N_4833);
nand U6508 (N_6508,N_5782,N_5333);
or U6509 (N_6509,N_5481,N_5442);
or U6510 (N_6510,N_5949,N_5626);
nor U6511 (N_6511,N_4786,N_5268);
or U6512 (N_6512,N_5421,N_5785);
and U6513 (N_6513,N_5183,N_5319);
nor U6514 (N_6514,N_4643,N_5336);
and U6515 (N_6515,N_5469,N_4952);
or U6516 (N_6516,N_5999,N_4769);
nand U6517 (N_6517,N_5986,N_4672);
nor U6518 (N_6518,N_5665,N_5638);
nand U6519 (N_6519,N_4777,N_5000);
nand U6520 (N_6520,N_5033,N_5849);
and U6521 (N_6521,N_5497,N_5926);
xnor U6522 (N_6522,N_4941,N_4700);
xnor U6523 (N_6523,N_5627,N_5967);
and U6524 (N_6524,N_5776,N_5669);
and U6525 (N_6525,N_4560,N_5762);
xnor U6526 (N_6526,N_4838,N_5515);
and U6527 (N_6527,N_5658,N_5930);
nor U6528 (N_6528,N_4866,N_5585);
xor U6529 (N_6529,N_5069,N_5914);
nand U6530 (N_6530,N_5423,N_4634);
nor U6531 (N_6531,N_5580,N_4921);
nand U6532 (N_6532,N_5095,N_4704);
and U6533 (N_6533,N_4800,N_4920);
xnor U6534 (N_6534,N_4975,N_5112);
nand U6535 (N_6535,N_5457,N_5379);
and U6536 (N_6536,N_5651,N_5527);
nor U6537 (N_6537,N_5634,N_4533);
nor U6538 (N_6538,N_5894,N_5179);
nor U6539 (N_6539,N_5683,N_5622);
xor U6540 (N_6540,N_5896,N_4965);
or U6541 (N_6541,N_5730,N_5291);
nand U6542 (N_6542,N_5309,N_4958);
and U6543 (N_6543,N_5722,N_5858);
and U6544 (N_6544,N_4697,N_4694);
xor U6545 (N_6545,N_5138,N_5881);
or U6546 (N_6546,N_4999,N_5272);
nor U6547 (N_6547,N_5723,N_5880);
nand U6548 (N_6548,N_5190,N_4854);
nor U6549 (N_6549,N_4647,N_4939);
and U6550 (N_6550,N_5817,N_5206);
and U6551 (N_6551,N_5990,N_5396);
xor U6552 (N_6552,N_5055,N_4907);
and U6553 (N_6553,N_4644,N_5855);
nand U6554 (N_6554,N_5037,N_4816);
xnor U6555 (N_6555,N_4984,N_5741);
nand U6556 (N_6556,N_5433,N_4904);
xor U6557 (N_6557,N_5207,N_4537);
nor U6558 (N_6558,N_5822,N_5671);
or U6559 (N_6559,N_4982,N_5030);
or U6560 (N_6560,N_4544,N_4942);
or U6561 (N_6561,N_5565,N_5510);
and U6562 (N_6562,N_5335,N_5524);
nand U6563 (N_6563,N_5937,N_5618);
nand U6564 (N_6564,N_4870,N_4909);
xnor U6565 (N_6565,N_4842,N_5538);
nor U6566 (N_6566,N_4976,N_5596);
or U6567 (N_6567,N_5499,N_5948);
or U6568 (N_6568,N_4690,N_5460);
nand U6569 (N_6569,N_5411,N_5195);
xor U6570 (N_6570,N_4569,N_5443);
nand U6571 (N_6571,N_5989,N_5193);
xnor U6572 (N_6572,N_4759,N_5128);
nand U6573 (N_6573,N_4755,N_4793);
or U6574 (N_6574,N_4513,N_4804);
nor U6575 (N_6575,N_5840,N_5851);
nor U6576 (N_6576,N_5466,N_5372);
xor U6577 (N_6577,N_4598,N_5464);
xor U6578 (N_6578,N_4673,N_4619);
xnor U6579 (N_6579,N_5375,N_5436);
xnor U6580 (N_6580,N_4881,N_5299);
and U6581 (N_6581,N_5151,N_4780);
nor U6582 (N_6582,N_5215,N_5611);
or U6583 (N_6583,N_4612,N_5608);
and U6584 (N_6584,N_5718,N_4626);
or U6585 (N_6585,N_4752,N_5172);
nand U6586 (N_6586,N_5140,N_5118);
nor U6587 (N_6587,N_5953,N_5918);
nor U6588 (N_6588,N_4653,N_5100);
or U6589 (N_6589,N_5137,N_4674);
and U6590 (N_6590,N_4990,N_5900);
nor U6591 (N_6591,N_5314,N_5115);
and U6592 (N_6592,N_5376,N_5166);
xnor U6593 (N_6593,N_5083,N_5209);
or U6594 (N_6594,N_4805,N_4579);
and U6595 (N_6595,N_5096,N_4931);
or U6596 (N_6596,N_5391,N_4712);
and U6597 (N_6597,N_5174,N_4709);
xor U6598 (N_6598,N_5090,N_4729);
nor U6599 (N_6599,N_5198,N_4924);
or U6600 (N_6600,N_4985,N_5592);
nand U6601 (N_6601,N_5415,N_4992);
nor U6602 (N_6602,N_5856,N_5257);
or U6603 (N_6603,N_5061,N_5678);
xnor U6604 (N_6604,N_5834,N_4916);
xnor U6605 (N_6605,N_5092,N_5252);
xnor U6606 (N_6606,N_5262,N_5994);
xor U6607 (N_6607,N_5068,N_4552);
and U6608 (N_6608,N_4855,N_4650);
and U6609 (N_6609,N_5905,N_5187);
and U6610 (N_6610,N_4531,N_4506);
xnor U6611 (N_6611,N_5980,N_4662);
nor U6612 (N_6612,N_5553,N_5886);
or U6613 (N_6613,N_5359,N_5642);
and U6614 (N_6614,N_5098,N_4558);
or U6615 (N_6615,N_5053,N_5736);
or U6616 (N_6616,N_5226,N_4580);
nor U6617 (N_6617,N_4979,N_4693);
nand U6618 (N_6618,N_5947,N_4565);
nand U6619 (N_6619,N_5031,N_4933);
or U6620 (N_6620,N_4925,N_4845);
xor U6621 (N_6621,N_5868,N_4917);
nor U6622 (N_6622,N_5028,N_4645);
or U6623 (N_6623,N_5566,N_5944);
nor U6624 (N_6624,N_5306,N_5670);
nand U6625 (N_6625,N_5176,N_5548);
nand U6626 (N_6626,N_5534,N_5951);
nor U6627 (N_6627,N_4997,N_4658);
xnor U6628 (N_6628,N_5764,N_5950);
nand U6629 (N_6629,N_4872,N_4857);
nand U6630 (N_6630,N_5322,N_4581);
xnor U6631 (N_6631,N_5148,N_5557);
or U6632 (N_6632,N_4621,N_5467);
nand U6633 (N_6633,N_5076,N_5760);
nand U6634 (N_6634,N_5220,N_5885);
xor U6635 (N_6635,N_5758,N_5742);
nand U6636 (N_6636,N_5103,N_5451);
and U6637 (N_6637,N_5361,N_5240);
or U6638 (N_6638,N_5841,N_4991);
and U6639 (N_6639,N_4823,N_4711);
nand U6640 (N_6640,N_5996,N_5506);
and U6641 (N_6641,N_5438,N_5964);
nor U6642 (N_6642,N_5985,N_4524);
xnor U6643 (N_6643,N_5455,N_4594);
or U6644 (N_6644,N_4656,N_5907);
and U6645 (N_6645,N_5810,N_5532);
nand U6646 (N_6646,N_5185,N_5649);
and U6647 (N_6647,N_5025,N_4960);
and U6648 (N_6648,N_5064,N_5468);
xor U6649 (N_6649,N_5302,N_5755);
nand U6650 (N_6650,N_4817,N_5446);
nor U6651 (N_6651,N_5719,N_5699);
xnor U6652 (N_6652,N_5072,N_5870);
xnor U6653 (N_6653,N_5825,N_5512);
nor U6654 (N_6654,N_4971,N_5369);
or U6655 (N_6655,N_4525,N_5237);
xnor U6656 (N_6656,N_5606,N_4901);
nand U6657 (N_6657,N_4632,N_4610);
xor U6658 (N_6658,N_4595,N_4509);
nand U6659 (N_6659,N_5184,N_4677);
or U6660 (N_6660,N_5965,N_4713);
nor U6661 (N_6661,N_5957,N_5097);
nor U6662 (N_6662,N_4758,N_5728);
nor U6663 (N_6663,N_4886,N_5431);
nor U6664 (N_6664,N_5408,N_4898);
nor U6665 (N_6665,N_5205,N_5398);
nand U6666 (N_6666,N_5024,N_5961);
nand U6667 (N_6667,N_4879,N_5564);
xor U6668 (N_6668,N_5663,N_5901);
nor U6669 (N_6669,N_5422,N_5452);
nor U6670 (N_6670,N_5567,N_5345);
and U6671 (N_6671,N_5019,N_4739);
xnor U6672 (N_6672,N_5201,N_4682);
and U6673 (N_6673,N_5737,N_4646);
nor U6674 (N_6674,N_4829,N_4502);
and U6675 (N_6675,N_5275,N_5744);
or U6676 (N_6676,N_5428,N_5974);
nor U6677 (N_6677,N_5384,N_4877);
nor U6678 (N_6678,N_5589,N_5779);
nor U6679 (N_6679,N_4657,N_5749);
or U6680 (N_6680,N_5507,N_5493);
or U6681 (N_6681,N_5228,N_5705);
nand U6682 (N_6682,N_5052,N_5036);
xnor U6683 (N_6683,N_4554,N_5733);
nor U6684 (N_6684,N_5963,N_5004);
or U6685 (N_6685,N_4651,N_5086);
nand U6686 (N_6686,N_5962,N_4818);
nand U6687 (N_6687,N_5289,N_5655);
nor U6688 (N_6688,N_5619,N_5169);
xnor U6689 (N_6689,N_5450,N_5049);
xor U6690 (N_6690,N_5448,N_4518);
xnor U6691 (N_6691,N_5562,N_5298);
or U6692 (N_6692,N_5550,N_4730);
nor U6693 (N_6693,N_5360,N_4649);
nand U6694 (N_6694,N_5075,N_5267);
or U6695 (N_6695,N_4858,N_4685);
or U6696 (N_6696,N_5054,N_5643);
or U6697 (N_6697,N_5826,N_4889);
xnor U6698 (N_6698,N_5694,N_4812);
or U6699 (N_6699,N_4536,N_5124);
nand U6700 (N_6700,N_5236,N_4605);
nand U6701 (N_6701,N_5650,N_5932);
nor U6702 (N_6702,N_4853,N_5893);
or U6703 (N_6703,N_5613,N_4564);
xor U6704 (N_6704,N_5852,N_5743);
or U6705 (N_6705,N_5048,N_5217);
xor U6706 (N_6706,N_5047,N_5798);
and U6707 (N_6707,N_5063,N_5545);
or U6708 (N_6708,N_4683,N_4894);
xor U6709 (N_6709,N_5864,N_4703);
xnor U6710 (N_6710,N_5144,N_4944);
xor U6711 (N_6711,N_4591,N_5482);
or U6712 (N_6712,N_5753,N_5549);
or U6713 (N_6713,N_5242,N_5685);
xor U6714 (N_6714,N_5713,N_5225);
or U6715 (N_6715,N_5547,N_4582);
xor U6716 (N_6716,N_5617,N_5165);
and U6717 (N_6717,N_4861,N_5934);
or U6718 (N_6718,N_5775,N_5710);
nor U6719 (N_6719,N_5276,N_5770);
or U6720 (N_6720,N_5287,N_5400);
and U6721 (N_6721,N_5898,N_5177);
xnor U6722 (N_6722,N_5489,N_4724);
and U6723 (N_6723,N_5266,N_5285);
xnor U6724 (N_6724,N_4639,N_4873);
xor U6725 (N_6725,N_5765,N_5085);
xor U6726 (N_6726,N_5445,N_4880);
xnor U6727 (N_6727,N_5386,N_5814);
and U6728 (N_6728,N_5909,N_5009);
xnor U6729 (N_6729,N_5931,N_4631);
nand U6730 (N_6730,N_5917,N_4831);
or U6731 (N_6731,N_5904,N_4655);
or U6732 (N_6732,N_4832,N_5211);
or U6733 (N_6733,N_5865,N_5084);
or U6734 (N_6734,N_5544,N_4574);
or U6735 (N_6735,N_4766,N_5837);
or U6736 (N_6736,N_5533,N_5487);
xnor U6737 (N_6737,N_4791,N_4535);
xnor U6738 (N_6738,N_5311,N_4583);
xnor U6739 (N_6739,N_5647,N_5501);
xor U6740 (N_6740,N_5182,N_4918);
and U6741 (N_6741,N_5844,N_4654);
and U6742 (N_6742,N_4784,N_4668);
xnor U6743 (N_6743,N_5044,N_5370);
nand U6744 (N_6744,N_5101,N_4811);
nand U6745 (N_6745,N_4844,N_4919);
or U6746 (N_6746,N_4799,N_5321);
xnor U6747 (N_6747,N_5062,N_5249);
xnor U6748 (N_6748,N_5265,N_4664);
nand U6749 (N_6749,N_4663,N_4970);
xor U6750 (N_6750,N_5750,N_5865);
nand U6751 (N_6751,N_5866,N_5072);
and U6752 (N_6752,N_5449,N_5921);
xor U6753 (N_6753,N_5914,N_5709);
nor U6754 (N_6754,N_4963,N_5655);
or U6755 (N_6755,N_4525,N_5741);
or U6756 (N_6756,N_5027,N_5291);
and U6757 (N_6757,N_5776,N_4780);
xor U6758 (N_6758,N_5263,N_5693);
nor U6759 (N_6759,N_5203,N_4646);
xnor U6760 (N_6760,N_5720,N_4667);
or U6761 (N_6761,N_5718,N_5942);
xor U6762 (N_6762,N_5393,N_5256);
nor U6763 (N_6763,N_5942,N_4996);
xnor U6764 (N_6764,N_5493,N_5623);
nor U6765 (N_6765,N_5387,N_5148);
or U6766 (N_6766,N_5371,N_5457);
and U6767 (N_6767,N_5657,N_4943);
or U6768 (N_6768,N_4804,N_5135);
or U6769 (N_6769,N_5966,N_4775);
or U6770 (N_6770,N_4790,N_5192);
xor U6771 (N_6771,N_5468,N_4862);
nor U6772 (N_6772,N_5270,N_4961);
or U6773 (N_6773,N_4891,N_5235);
nand U6774 (N_6774,N_5136,N_5023);
nor U6775 (N_6775,N_5196,N_4904);
xor U6776 (N_6776,N_5118,N_4681);
nor U6777 (N_6777,N_4553,N_5621);
and U6778 (N_6778,N_4785,N_5455);
nor U6779 (N_6779,N_4602,N_4797);
and U6780 (N_6780,N_4561,N_5200);
xnor U6781 (N_6781,N_4957,N_5577);
or U6782 (N_6782,N_5187,N_5698);
and U6783 (N_6783,N_4926,N_5039);
and U6784 (N_6784,N_5543,N_5358);
nand U6785 (N_6785,N_5936,N_5017);
or U6786 (N_6786,N_5440,N_5359);
and U6787 (N_6787,N_4615,N_4762);
xnor U6788 (N_6788,N_4999,N_5159);
and U6789 (N_6789,N_5917,N_5859);
nand U6790 (N_6790,N_5270,N_4742);
and U6791 (N_6791,N_5737,N_5009);
xnor U6792 (N_6792,N_5993,N_4782);
and U6793 (N_6793,N_5473,N_5676);
xor U6794 (N_6794,N_5741,N_5860);
and U6795 (N_6795,N_4816,N_5758);
xnor U6796 (N_6796,N_5163,N_5568);
or U6797 (N_6797,N_5194,N_5651);
nor U6798 (N_6798,N_5850,N_5765);
xor U6799 (N_6799,N_5506,N_5429);
nor U6800 (N_6800,N_5336,N_4785);
xor U6801 (N_6801,N_4925,N_5045);
or U6802 (N_6802,N_5149,N_5385);
xnor U6803 (N_6803,N_5344,N_5679);
nand U6804 (N_6804,N_5783,N_4750);
and U6805 (N_6805,N_5786,N_4501);
nor U6806 (N_6806,N_5353,N_5612);
nor U6807 (N_6807,N_5534,N_5532);
and U6808 (N_6808,N_4947,N_5263);
xnor U6809 (N_6809,N_5910,N_5897);
nand U6810 (N_6810,N_5219,N_5441);
nand U6811 (N_6811,N_5737,N_5531);
nand U6812 (N_6812,N_5176,N_5950);
or U6813 (N_6813,N_5769,N_4816);
nor U6814 (N_6814,N_5313,N_5300);
xor U6815 (N_6815,N_5191,N_5775);
and U6816 (N_6816,N_5318,N_5270);
xor U6817 (N_6817,N_5737,N_5912);
nand U6818 (N_6818,N_5543,N_5584);
or U6819 (N_6819,N_4707,N_5578);
xnor U6820 (N_6820,N_5441,N_4954);
nand U6821 (N_6821,N_4967,N_5668);
xor U6822 (N_6822,N_4857,N_5182);
and U6823 (N_6823,N_4932,N_5551);
or U6824 (N_6824,N_4585,N_5104);
nand U6825 (N_6825,N_5548,N_4760);
and U6826 (N_6826,N_5406,N_5643);
and U6827 (N_6827,N_4616,N_5078);
nand U6828 (N_6828,N_5947,N_5470);
or U6829 (N_6829,N_5723,N_5190);
nor U6830 (N_6830,N_5703,N_4840);
nand U6831 (N_6831,N_5157,N_5151);
xnor U6832 (N_6832,N_5597,N_5559);
xnor U6833 (N_6833,N_5879,N_4812);
and U6834 (N_6834,N_5646,N_5997);
nor U6835 (N_6835,N_5854,N_4683);
xnor U6836 (N_6836,N_4888,N_4612);
xor U6837 (N_6837,N_5054,N_5346);
nand U6838 (N_6838,N_4661,N_5970);
nor U6839 (N_6839,N_5137,N_5224);
or U6840 (N_6840,N_5434,N_5452);
xor U6841 (N_6841,N_5165,N_5408);
nor U6842 (N_6842,N_5910,N_5588);
and U6843 (N_6843,N_5157,N_4977);
or U6844 (N_6844,N_4525,N_5416);
or U6845 (N_6845,N_5966,N_4876);
nand U6846 (N_6846,N_4740,N_4637);
nand U6847 (N_6847,N_5838,N_5611);
or U6848 (N_6848,N_5487,N_4965);
and U6849 (N_6849,N_5440,N_5852);
or U6850 (N_6850,N_5666,N_5026);
nor U6851 (N_6851,N_4697,N_4747);
nor U6852 (N_6852,N_4924,N_5146);
nor U6853 (N_6853,N_4866,N_5132);
nand U6854 (N_6854,N_4839,N_4976);
xor U6855 (N_6855,N_5792,N_4619);
and U6856 (N_6856,N_5391,N_4828);
and U6857 (N_6857,N_5706,N_4508);
and U6858 (N_6858,N_5580,N_4915);
xor U6859 (N_6859,N_4555,N_5433);
xor U6860 (N_6860,N_5246,N_5351);
or U6861 (N_6861,N_5143,N_4778);
nor U6862 (N_6862,N_4623,N_5269);
nand U6863 (N_6863,N_5809,N_4812);
xor U6864 (N_6864,N_5777,N_5841);
nand U6865 (N_6865,N_5389,N_5065);
and U6866 (N_6866,N_4876,N_5971);
or U6867 (N_6867,N_5190,N_5804);
and U6868 (N_6868,N_4869,N_5721);
nand U6869 (N_6869,N_5940,N_4778);
or U6870 (N_6870,N_4614,N_4829);
nor U6871 (N_6871,N_5940,N_5425);
or U6872 (N_6872,N_5678,N_5932);
nand U6873 (N_6873,N_4803,N_4514);
nand U6874 (N_6874,N_5109,N_5350);
or U6875 (N_6875,N_5622,N_5756);
or U6876 (N_6876,N_5533,N_5557);
nand U6877 (N_6877,N_5239,N_5783);
nor U6878 (N_6878,N_5784,N_5147);
nand U6879 (N_6879,N_5840,N_5392);
nor U6880 (N_6880,N_4786,N_5313);
and U6881 (N_6881,N_5261,N_4644);
nor U6882 (N_6882,N_5486,N_4529);
nand U6883 (N_6883,N_5431,N_5304);
nand U6884 (N_6884,N_5883,N_5573);
xnor U6885 (N_6885,N_4542,N_5903);
nor U6886 (N_6886,N_5576,N_4881);
nand U6887 (N_6887,N_4912,N_4977);
and U6888 (N_6888,N_4694,N_5759);
nor U6889 (N_6889,N_5921,N_5068);
nand U6890 (N_6890,N_5469,N_5010);
nor U6891 (N_6891,N_4949,N_4720);
nand U6892 (N_6892,N_5310,N_4873);
nand U6893 (N_6893,N_5603,N_4618);
or U6894 (N_6894,N_4617,N_5664);
nor U6895 (N_6895,N_5531,N_5952);
nand U6896 (N_6896,N_5572,N_5090);
nor U6897 (N_6897,N_5034,N_5976);
nor U6898 (N_6898,N_5790,N_5702);
nor U6899 (N_6899,N_4614,N_4742);
or U6900 (N_6900,N_5291,N_4856);
nor U6901 (N_6901,N_5991,N_5528);
xor U6902 (N_6902,N_5316,N_5878);
and U6903 (N_6903,N_4711,N_4728);
nor U6904 (N_6904,N_5138,N_4561);
xnor U6905 (N_6905,N_5369,N_4956);
and U6906 (N_6906,N_4613,N_5770);
or U6907 (N_6907,N_5448,N_5526);
and U6908 (N_6908,N_5501,N_4804);
and U6909 (N_6909,N_4665,N_5324);
nand U6910 (N_6910,N_4936,N_4815);
and U6911 (N_6911,N_5726,N_5420);
nand U6912 (N_6912,N_5406,N_4653);
or U6913 (N_6913,N_4673,N_4729);
xnor U6914 (N_6914,N_4591,N_4751);
nor U6915 (N_6915,N_4731,N_5233);
nand U6916 (N_6916,N_5860,N_5848);
nand U6917 (N_6917,N_5984,N_5473);
nand U6918 (N_6918,N_5163,N_4864);
and U6919 (N_6919,N_4955,N_5584);
and U6920 (N_6920,N_5943,N_4556);
or U6921 (N_6921,N_5609,N_4698);
and U6922 (N_6922,N_5716,N_5868);
nand U6923 (N_6923,N_5351,N_5199);
or U6924 (N_6924,N_4613,N_4690);
xor U6925 (N_6925,N_4762,N_4736);
or U6926 (N_6926,N_5308,N_4784);
xnor U6927 (N_6927,N_5332,N_5639);
nand U6928 (N_6928,N_5865,N_5471);
xor U6929 (N_6929,N_4983,N_5827);
and U6930 (N_6930,N_5742,N_4979);
and U6931 (N_6931,N_5663,N_4862);
nand U6932 (N_6932,N_5380,N_5268);
or U6933 (N_6933,N_5442,N_4742);
nand U6934 (N_6934,N_4795,N_5409);
nor U6935 (N_6935,N_4944,N_5186);
or U6936 (N_6936,N_4514,N_4645);
nand U6937 (N_6937,N_5279,N_5639);
and U6938 (N_6938,N_4718,N_4736);
nand U6939 (N_6939,N_5460,N_5331);
and U6940 (N_6940,N_5549,N_4655);
xor U6941 (N_6941,N_5400,N_4919);
nor U6942 (N_6942,N_5099,N_4643);
and U6943 (N_6943,N_5319,N_5178);
nand U6944 (N_6944,N_5476,N_4831);
and U6945 (N_6945,N_5814,N_4690);
or U6946 (N_6946,N_5180,N_4514);
or U6947 (N_6947,N_5629,N_5128);
nand U6948 (N_6948,N_5905,N_4834);
nor U6949 (N_6949,N_4796,N_4732);
or U6950 (N_6950,N_5527,N_5260);
nor U6951 (N_6951,N_5227,N_4946);
or U6952 (N_6952,N_4560,N_4871);
nor U6953 (N_6953,N_4648,N_5824);
and U6954 (N_6954,N_4733,N_5115);
and U6955 (N_6955,N_4675,N_5224);
nand U6956 (N_6956,N_5959,N_5886);
nor U6957 (N_6957,N_4659,N_5847);
and U6958 (N_6958,N_5804,N_5783);
nand U6959 (N_6959,N_4886,N_4953);
xnor U6960 (N_6960,N_5658,N_4534);
nand U6961 (N_6961,N_5628,N_5193);
and U6962 (N_6962,N_5633,N_5542);
and U6963 (N_6963,N_5015,N_5626);
nor U6964 (N_6964,N_5891,N_5440);
xor U6965 (N_6965,N_4598,N_4673);
nand U6966 (N_6966,N_5697,N_4791);
nor U6967 (N_6967,N_4891,N_5748);
nand U6968 (N_6968,N_5375,N_5303);
nor U6969 (N_6969,N_4621,N_5435);
or U6970 (N_6970,N_5990,N_5841);
nand U6971 (N_6971,N_4761,N_5147);
and U6972 (N_6972,N_4799,N_5395);
nand U6973 (N_6973,N_5972,N_5499);
or U6974 (N_6974,N_5860,N_5880);
nor U6975 (N_6975,N_5762,N_5676);
or U6976 (N_6976,N_5688,N_5330);
or U6977 (N_6977,N_5442,N_5322);
xor U6978 (N_6978,N_5181,N_5614);
or U6979 (N_6979,N_5920,N_4839);
nand U6980 (N_6980,N_4972,N_5111);
or U6981 (N_6981,N_5544,N_4869);
nand U6982 (N_6982,N_5355,N_5039);
nor U6983 (N_6983,N_5198,N_4596);
or U6984 (N_6984,N_4509,N_4660);
or U6985 (N_6985,N_4759,N_5704);
and U6986 (N_6986,N_5499,N_5175);
and U6987 (N_6987,N_5167,N_5189);
and U6988 (N_6988,N_5071,N_5413);
and U6989 (N_6989,N_5133,N_4747);
nand U6990 (N_6990,N_5631,N_5668);
xnor U6991 (N_6991,N_4760,N_5398);
xor U6992 (N_6992,N_5566,N_5349);
or U6993 (N_6993,N_5079,N_5439);
nand U6994 (N_6994,N_5139,N_5274);
or U6995 (N_6995,N_5493,N_5591);
or U6996 (N_6996,N_5512,N_5811);
nand U6997 (N_6997,N_5937,N_4776);
xnor U6998 (N_6998,N_4787,N_4676);
and U6999 (N_6999,N_5803,N_5184);
nand U7000 (N_7000,N_5035,N_4952);
xnor U7001 (N_7001,N_5563,N_5508);
nor U7002 (N_7002,N_5443,N_4806);
xnor U7003 (N_7003,N_4913,N_5736);
nor U7004 (N_7004,N_5559,N_5682);
and U7005 (N_7005,N_4818,N_5907);
xor U7006 (N_7006,N_5625,N_5353);
xnor U7007 (N_7007,N_5129,N_5940);
nand U7008 (N_7008,N_5962,N_4546);
xnor U7009 (N_7009,N_5397,N_4555);
xnor U7010 (N_7010,N_5538,N_4787);
and U7011 (N_7011,N_4975,N_5367);
xor U7012 (N_7012,N_5398,N_5450);
xor U7013 (N_7013,N_4848,N_5476);
nor U7014 (N_7014,N_5137,N_5939);
or U7015 (N_7015,N_4509,N_5387);
or U7016 (N_7016,N_5815,N_4720);
xnor U7017 (N_7017,N_5841,N_5512);
or U7018 (N_7018,N_5577,N_4528);
nor U7019 (N_7019,N_5479,N_4658);
nor U7020 (N_7020,N_5709,N_4937);
nand U7021 (N_7021,N_5083,N_4501);
nor U7022 (N_7022,N_5413,N_5875);
nand U7023 (N_7023,N_4622,N_5164);
or U7024 (N_7024,N_4782,N_4679);
or U7025 (N_7025,N_4648,N_4849);
xor U7026 (N_7026,N_5443,N_4695);
xnor U7027 (N_7027,N_5903,N_4861);
xor U7028 (N_7028,N_5316,N_5666);
or U7029 (N_7029,N_5379,N_4800);
nor U7030 (N_7030,N_5375,N_5196);
nor U7031 (N_7031,N_5002,N_5824);
or U7032 (N_7032,N_4512,N_5200);
and U7033 (N_7033,N_4560,N_5544);
or U7034 (N_7034,N_5153,N_5610);
nand U7035 (N_7035,N_4962,N_5393);
and U7036 (N_7036,N_5415,N_4657);
and U7037 (N_7037,N_4608,N_4776);
nor U7038 (N_7038,N_4843,N_4756);
and U7039 (N_7039,N_5136,N_4731);
and U7040 (N_7040,N_5460,N_5694);
nor U7041 (N_7041,N_5330,N_4816);
nand U7042 (N_7042,N_5802,N_5231);
nor U7043 (N_7043,N_4879,N_4521);
xor U7044 (N_7044,N_5811,N_5242);
or U7045 (N_7045,N_4532,N_5333);
nand U7046 (N_7046,N_4900,N_5467);
and U7047 (N_7047,N_5813,N_5263);
or U7048 (N_7048,N_5833,N_5691);
and U7049 (N_7049,N_5526,N_5342);
or U7050 (N_7050,N_5874,N_5197);
or U7051 (N_7051,N_5907,N_4626);
nor U7052 (N_7052,N_5170,N_5177);
nor U7053 (N_7053,N_5235,N_5648);
or U7054 (N_7054,N_5741,N_5344);
and U7055 (N_7055,N_5133,N_4607);
xor U7056 (N_7056,N_5916,N_4799);
and U7057 (N_7057,N_5364,N_4921);
or U7058 (N_7058,N_4745,N_5118);
or U7059 (N_7059,N_5757,N_4911);
and U7060 (N_7060,N_5108,N_4983);
xnor U7061 (N_7061,N_4788,N_5864);
or U7062 (N_7062,N_5966,N_5597);
or U7063 (N_7063,N_5219,N_5012);
nor U7064 (N_7064,N_4618,N_4790);
nor U7065 (N_7065,N_5163,N_5609);
nor U7066 (N_7066,N_5206,N_5472);
nand U7067 (N_7067,N_5465,N_5932);
and U7068 (N_7068,N_5736,N_5117);
nand U7069 (N_7069,N_5319,N_4989);
or U7070 (N_7070,N_5099,N_4819);
and U7071 (N_7071,N_5628,N_5415);
nand U7072 (N_7072,N_5442,N_4863);
xnor U7073 (N_7073,N_4790,N_5640);
or U7074 (N_7074,N_5009,N_5661);
and U7075 (N_7075,N_4678,N_4709);
xnor U7076 (N_7076,N_5715,N_5003);
or U7077 (N_7077,N_5269,N_5758);
or U7078 (N_7078,N_4687,N_4995);
nor U7079 (N_7079,N_4976,N_5456);
nor U7080 (N_7080,N_4840,N_5609);
and U7081 (N_7081,N_4855,N_5763);
nand U7082 (N_7082,N_5693,N_5827);
xnor U7083 (N_7083,N_4567,N_5003);
xor U7084 (N_7084,N_4518,N_5029);
and U7085 (N_7085,N_5132,N_5243);
nor U7086 (N_7086,N_5883,N_5460);
or U7087 (N_7087,N_5336,N_4518);
and U7088 (N_7088,N_4834,N_5483);
nand U7089 (N_7089,N_4759,N_4644);
nor U7090 (N_7090,N_5241,N_4914);
nor U7091 (N_7091,N_5799,N_4593);
or U7092 (N_7092,N_5836,N_5763);
nor U7093 (N_7093,N_5261,N_5209);
and U7094 (N_7094,N_5038,N_5859);
nand U7095 (N_7095,N_5406,N_5610);
nor U7096 (N_7096,N_4651,N_5348);
nand U7097 (N_7097,N_5383,N_5032);
nor U7098 (N_7098,N_5359,N_5196);
xor U7099 (N_7099,N_5059,N_4772);
and U7100 (N_7100,N_5734,N_5674);
or U7101 (N_7101,N_5447,N_5742);
xor U7102 (N_7102,N_5592,N_4563);
xnor U7103 (N_7103,N_5690,N_5971);
or U7104 (N_7104,N_5250,N_4937);
nor U7105 (N_7105,N_5184,N_5590);
and U7106 (N_7106,N_5518,N_5997);
or U7107 (N_7107,N_5664,N_4917);
xor U7108 (N_7108,N_5359,N_5456);
and U7109 (N_7109,N_5927,N_5245);
nor U7110 (N_7110,N_4704,N_5925);
and U7111 (N_7111,N_4703,N_5496);
and U7112 (N_7112,N_5374,N_5784);
nand U7113 (N_7113,N_4941,N_5772);
nor U7114 (N_7114,N_5463,N_5704);
or U7115 (N_7115,N_5438,N_5266);
nor U7116 (N_7116,N_5515,N_5172);
nand U7117 (N_7117,N_5835,N_4781);
xor U7118 (N_7118,N_5620,N_5602);
or U7119 (N_7119,N_4993,N_5316);
nor U7120 (N_7120,N_5493,N_5482);
or U7121 (N_7121,N_4797,N_4969);
and U7122 (N_7122,N_5897,N_5762);
xor U7123 (N_7123,N_5994,N_5110);
and U7124 (N_7124,N_5131,N_5795);
xnor U7125 (N_7125,N_5345,N_4622);
xor U7126 (N_7126,N_4641,N_5680);
nor U7127 (N_7127,N_4580,N_5217);
nand U7128 (N_7128,N_4652,N_4823);
nand U7129 (N_7129,N_5565,N_4998);
xnor U7130 (N_7130,N_4850,N_4946);
nand U7131 (N_7131,N_5133,N_4803);
nor U7132 (N_7132,N_5112,N_5022);
and U7133 (N_7133,N_4863,N_5804);
or U7134 (N_7134,N_5399,N_5977);
or U7135 (N_7135,N_5513,N_5224);
and U7136 (N_7136,N_5695,N_5641);
xnor U7137 (N_7137,N_4879,N_5019);
nand U7138 (N_7138,N_5498,N_5924);
nand U7139 (N_7139,N_5375,N_5615);
and U7140 (N_7140,N_4652,N_5190);
and U7141 (N_7141,N_5520,N_5150);
xor U7142 (N_7142,N_5378,N_5688);
or U7143 (N_7143,N_5809,N_5650);
nor U7144 (N_7144,N_5886,N_4862);
and U7145 (N_7145,N_5224,N_5967);
nand U7146 (N_7146,N_4679,N_4685);
xor U7147 (N_7147,N_5443,N_4693);
xnor U7148 (N_7148,N_5186,N_5992);
and U7149 (N_7149,N_5868,N_5528);
and U7150 (N_7150,N_5931,N_5803);
xor U7151 (N_7151,N_5338,N_5598);
nor U7152 (N_7152,N_5452,N_5127);
nor U7153 (N_7153,N_4559,N_5937);
or U7154 (N_7154,N_4610,N_5905);
or U7155 (N_7155,N_4780,N_5763);
nor U7156 (N_7156,N_5513,N_5759);
nand U7157 (N_7157,N_5071,N_5344);
and U7158 (N_7158,N_5999,N_5151);
or U7159 (N_7159,N_5771,N_5487);
nand U7160 (N_7160,N_5974,N_5824);
nor U7161 (N_7161,N_5700,N_4621);
and U7162 (N_7162,N_5003,N_5941);
xnor U7163 (N_7163,N_5006,N_5410);
nand U7164 (N_7164,N_5483,N_4773);
and U7165 (N_7165,N_5526,N_4919);
nor U7166 (N_7166,N_5932,N_5994);
xnor U7167 (N_7167,N_5745,N_5345);
or U7168 (N_7168,N_5921,N_5766);
and U7169 (N_7169,N_4725,N_5886);
and U7170 (N_7170,N_5098,N_5401);
nand U7171 (N_7171,N_5713,N_4689);
nor U7172 (N_7172,N_4890,N_5255);
nand U7173 (N_7173,N_5523,N_5144);
nor U7174 (N_7174,N_4662,N_5353);
and U7175 (N_7175,N_5577,N_4605);
nand U7176 (N_7176,N_5290,N_4564);
nand U7177 (N_7177,N_5413,N_4823);
and U7178 (N_7178,N_5468,N_4570);
nor U7179 (N_7179,N_5044,N_5705);
or U7180 (N_7180,N_5562,N_5703);
xnor U7181 (N_7181,N_5017,N_5543);
nor U7182 (N_7182,N_5075,N_5205);
nor U7183 (N_7183,N_4854,N_5748);
xnor U7184 (N_7184,N_4611,N_5240);
nor U7185 (N_7185,N_4555,N_4730);
nor U7186 (N_7186,N_4593,N_4613);
nand U7187 (N_7187,N_5385,N_5205);
nand U7188 (N_7188,N_5733,N_5396);
or U7189 (N_7189,N_5915,N_5904);
and U7190 (N_7190,N_4671,N_4788);
xnor U7191 (N_7191,N_5158,N_5074);
or U7192 (N_7192,N_5825,N_5487);
and U7193 (N_7193,N_5838,N_4849);
or U7194 (N_7194,N_4637,N_5731);
or U7195 (N_7195,N_5252,N_5865);
or U7196 (N_7196,N_4590,N_5685);
or U7197 (N_7197,N_5337,N_4816);
and U7198 (N_7198,N_5220,N_5871);
and U7199 (N_7199,N_4886,N_4655);
nand U7200 (N_7200,N_5607,N_5686);
or U7201 (N_7201,N_4529,N_4873);
xor U7202 (N_7202,N_5044,N_5459);
nand U7203 (N_7203,N_4978,N_5249);
nand U7204 (N_7204,N_5996,N_4556);
or U7205 (N_7205,N_5324,N_4770);
or U7206 (N_7206,N_5258,N_5194);
nand U7207 (N_7207,N_5506,N_5384);
or U7208 (N_7208,N_4590,N_4775);
nor U7209 (N_7209,N_5363,N_5132);
nand U7210 (N_7210,N_5404,N_5164);
nand U7211 (N_7211,N_5405,N_4738);
nand U7212 (N_7212,N_5756,N_5775);
nand U7213 (N_7213,N_4735,N_5930);
xnor U7214 (N_7214,N_4984,N_5069);
nor U7215 (N_7215,N_4808,N_4577);
or U7216 (N_7216,N_5260,N_5161);
or U7217 (N_7217,N_4827,N_5689);
nor U7218 (N_7218,N_4616,N_4510);
or U7219 (N_7219,N_5893,N_4630);
and U7220 (N_7220,N_5096,N_5718);
nand U7221 (N_7221,N_5006,N_5993);
nand U7222 (N_7222,N_5695,N_4963);
or U7223 (N_7223,N_4663,N_5925);
nand U7224 (N_7224,N_5968,N_5810);
nor U7225 (N_7225,N_5686,N_5410);
nand U7226 (N_7226,N_5204,N_5644);
xor U7227 (N_7227,N_4511,N_4837);
or U7228 (N_7228,N_4513,N_5284);
xor U7229 (N_7229,N_5452,N_5808);
nand U7230 (N_7230,N_4838,N_4580);
xnor U7231 (N_7231,N_5425,N_5531);
xnor U7232 (N_7232,N_4895,N_5307);
or U7233 (N_7233,N_5522,N_5940);
nor U7234 (N_7234,N_4907,N_4530);
nor U7235 (N_7235,N_4544,N_5352);
nor U7236 (N_7236,N_5885,N_4959);
nor U7237 (N_7237,N_5472,N_4772);
or U7238 (N_7238,N_5842,N_5869);
nor U7239 (N_7239,N_4829,N_4504);
nor U7240 (N_7240,N_5773,N_5506);
and U7241 (N_7241,N_5556,N_5198);
nand U7242 (N_7242,N_5145,N_4657);
xnor U7243 (N_7243,N_5952,N_4747);
or U7244 (N_7244,N_5270,N_5603);
nor U7245 (N_7245,N_5263,N_5741);
or U7246 (N_7246,N_4706,N_5619);
nor U7247 (N_7247,N_5479,N_4901);
nand U7248 (N_7248,N_4997,N_4897);
xnor U7249 (N_7249,N_5715,N_5558);
nor U7250 (N_7250,N_4783,N_5380);
and U7251 (N_7251,N_5300,N_5623);
or U7252 (N_7252,N_4656,N_4991);
or U7253 (N_7253,N_5331,N_4770);
xor U7254 (N_7254,N_5555,N_5447);
or U7255 (N_7255,N_4611,N_5334);
xor U7256 (N_7256,N_5373,N_4506);
or U7257 (N_7257,N_5116,N_4527);
or U7258 (N_7258,N_5788,N_5792);
nand U7259 (N_7259,N_5733,N_4541);
nand U7260 (N_7260,N_5208,N_4888);
or U7261 (N_7261,N_5149,N_5687);
nand U7262 (N_7262,N_4884,N_4808);
xor U7263 (N_7263,N_5375,N_4993);
nand U7264 (N_7264,N_5729,N_5066);
nand U7265 (N_7265,N_5767,N_4734);
nor U7266 (N_7266,N_5303,N_5455);
nand U7267 (N_7267,N_4730,N_5178);
and U7268 (N_7268,N_4688,N_4849);
nor U7269 (N_7269,N_5440,N_5547);
and U7270 (N_7270,N_5233,N_5746);
nand U7271 (N_7271,N_5095,N_5961);
nor U7272 (N_7272,N_5737,N_5676);
nand U7273 (N_7273,N_5532,N_5328);
and U7274 (N_7274,N_5140,N_5170);
or U7275 (N_7275,N_5147,N_5254);
nand U7276 (N_7276,N_4532,N_5651);
and U7277 (N_7277,N_4800,N_4862);
xnor U7278 (N_7278,N_5770,N_5400);
xor U7279 (N_7279,N_4992,N_5640);
nor U7280 (N_7280,N_5981,N_4821);
xnor U7281 (N_7281,N_5502,N_4784);
nand U7282 (N_7282,N_4938,N_5439);
nor U7283 (N_7283,N_5658,N_5062);
nor U7284 (N_7284,N_5188,N_4782);
and U7285 (N_7285,N_5611,N_4905);
and U7286 (N_7286,N_4686,N_5436);
or U7287 (N_7287,N_5088,N_4901);
and U7288 (N_7288,N_5836,N_4909);
nand U7289 (N_7289,N_5610,N_4539);
and U7290 (N_7290,N_5416,N_4676);
xor U7291 (N_7291,N_5484,N_5951);
xnor U7292 (N_7292,N_5221,N_5228);
xor U7293 (N_7293,N_5457,N_4815);
xor U7294 (N_7294,N_4841,N_5841);
nor U7295 (N_7295,N_5336,N_5581);
and U7296 (N_7296,N_5895,N_5026);
nor U7297 (N_7297,N_4944,N_5650);
nand U7298 (N_7298,N_5786,N_4514);
and U7299 (N_7299,N_5242,N_5379);
and U7300 (N_7300,N_5548,N_4717);
xor U7301 (N_7301,N_5351,N_5787);
and U7302 (N_7302,N_5508,N_5021);
or U7303 (N_7303,N_5298,N_4576);
nor U7304 (N_7304,N_5126,N_5193);
xnor U7305 (N_7305,N_5462,N_5857);
nor U7306 (N_7306,N_5418,N_5233);
nand U7307 (N_7307,N_5687,N_5660);
nor U7308 (N_7308,N_4829,N_5728);
xor U7309 (N_7309,N_4933,N_5432);
and U7310 (N_7310,N_4583,N_4602);
and U7311 (N_7311,N_5912,N_4984);
and U7312 (N_7312,N_4699,N_5420);
nand U7313 (N_7313,N_5675,N_5516);
nor U7314 (N_7314,N_5599,N_5844);
or U7315 (N_7315,N_5146,N_5641);
and U7316 (N_7316,N_5590,N_5460);
nor U7317 (N_7317,N_5242,N_4639);
xor U7318 (N_7318,N_5019,N_5706);
nor U7319 (N_7319,N_5851,N_5910);
and U7320 (N_7320,N_5395,N_5523);
nor U7321 (N_7321,N_5655,N_5277);
or U7322 (N_7322,N_4688,N_5688);
and U7323 (N_7323,N_5744,N_4981);
and U7324 (N_7324,N_5005,N_4880);
and U7325 (N_7325,N_5726,N_4927);
xor U7326 (N_7326,N_5246,N_5841);
nor U7327 (N_7327,N_4722,N_5814);
nand U7328 (N_7328,N_5802,N_4776);
or U7329 (N_7329,N_5092,N_4819);
xor U7330 (N_7330,N_5585,N_5032);
and U7331 (N_7331,N_4595,N_5906);
nor U7332 (N_7332,N_5349,N_5308);
or U7333 (N_7333,N_5193,N_4691);
or U7334 (N_7334,N_5378,N_4990);
or U7335 (N_7335,N_5182,N_5617);
or U7336 (N_7336,N_5797,N_4777);
and U7337 (N_7337,N_4827,N_4766);
or U7338 (N_7338,N_4554,N_5706);
nand U7339 (N_7339,N_5420,N_4540);
xnor U7340 (N_7340,N_4786,N_5626);
or U7341 (N_7341,N_5358,N_5729);
or U7342 (N_7342,N_5166,N_5640);
and U7343 (N_7343,N_4665,N_5692);
nand U7344 (N_7344,N_5223,N_5506);
nand U7345 (N_7345,N_5912,N_5861);
or U7346 (N_7346,N_5189,N_5517);
xnor U7347 (N_7347,N_5596,N_4553);
nor U7348 (N_7348,N_5286,N_4901);
nand U7349 (N_7349,N_4598,N_5630);
or U7350 (N_7350,N_5050,N_4675);
or U7351 (N_7351,N_5363,N_5415);
nand U7352 (N_7352,N_5633,N_5206);
nor U7353 (N_7353,N_5870,N_5039);
and U7354 (N_7354,N_5158,N_5493);
nand U7355 (N_7355,N_5103,N_5512);
nand U7356 (N_7356,N_4561,N_5787);
and U7357 (N_7357,N_4726,N_5177);
and U7358 (N_7358,N_5864,N_4602);
xnor U7359 (N_7359,N_5418,N_5731);
nand U7360 (N_7360,N_5515,N_5689);
nor U7361 (N_7361,N_5856,N_5827);
xnor U7362 (N_7362,N_5027,N_4996);
nor U7363 (N_7363,N_5229,N_5915);
and U7364 (N_7364,N_5349,N_4642);
nand U7365 (N_7365,N_5987,N_5074);
nor U7366 (N_7366,N_4678,N_4770);
and U7367 (N_7367,N_4946,N_4690);
or U7368 (N_7368,N_5997,N_4875);
and U7369 (N_7369,N_5492,N_5429);
xnor U7370 (N_7370,N_4607,N_5214);
or U7371 (N_7371,N_5418,N_4503);
and U7372 (N_7372,N_4647,N_4875);
xnor U7373 (N_7373,N_5324,N_4628);
or U7374 (N_7374,N_4946,N_4859);
and U7375 (N_7375,N_5362,N_4609);
xor U7376 (N_7376,N_4667,N_5287);
xor U7377 (N_7377,N_5351,N_4767);
and U7378 (N_7378,N_5062,N_5958);
or U7379 (N_7379,N_5209,N_5496);
xor U7380 (N_7380,N_4988,N_5940);
xor U7381 (N_7381,N_4986,N_5676);
xnor U7382 (N_7382,N_4843,N_4967);
or U7383 (N_7383,N_4807,N_5759);
or U7384 (N_7384,N_5991,N_4723);
nor U7385 (N_7385,N_4531,N_4529);
and U7386 (N_7386,N_4578,N_5299);
nand U7387 (N_7387,N_5265,N_5289);
nand U7388 (N_7388,N_5714,N_4694);
nand U7389 (N_7389,N_5808,N_4611);
xor U7390 (N_7390,N_4996,N_5490);
xnor U7391 (N_7391,N_5327,N_5852);
nand U7392 (N_7392,N_5044,N_4989);
nor U7393 (N_7393,N_4885,N_4689);
nand U7394 (N_7394,N_5451,N_4604);
nor U7395 (N_7395,N_5956,N_5109);
nand U7396 (N_7396,N_4567,N_5991);
xnor U7397 (N_7397,N_5010,N_4625);
nor U7398 (N_7398,N_5723,N_5511);
and U7399 (N_7399,N_4812,N_4699);
or U7400 (N_7400,N_4768,N_5503);
or U7401 (N_7401,N_5972,N_4894);
and U7402 (N_7402,N_4737,N_4983);
nand U7403 (N_7403,N_4970,N_5344);
and U7404 (N_7404,N_5316,N_4811);
or U7405 (N_7405,N_4774,N_5723);
or U7406 (N_7406,N_5626,N_5845);
nor U7407 (N_7407,N_5470,N_5898);
nor U7408 (N_7408,N_5351,N_5068);
xnor U7409 (N_7409,N_5094,N_4920);
and U7410 (N_7410,N_5753,N_4711);
or U7411 (N_7411,N_5694,N_4846);
and U7412 (N_7412,N_5278,N_4721);
or U7413 (N_7413,N_5318,N_5996);
or U7414 (N_7414,N_5336,N_5738);
nor U7415 (N_7415,N_5178,N_5591);
xnor U7416 (N_7416,N_5584,N_5957);
or U7417 (N_7417,N_5514,N_4651);
nand U7418 (N_7418,N_5970,N_4863);
or U7419 (N_7419,N_5390,N_4946);
and U7420 (N_7420,N_5626,N_4928);
xor U7421 (N_7421,N_5496,N_4986);
xor U7422 (N_7422,N_4774,N_4745);
and U7423 (N_7423,N_5005,N_5069);
and U7424 (N_7424,N_5963,N_5647);
nor U7425 (N_7425,N_5237,N_4562);
nor U7426 (N_7426,N_5683,N_5580);
nand U7427 (N_7427,N_5961,N_4656);
and U7428 (N_7428,N_5552,N_5285);
or U7429 (N_7429,N_5747,N_5479);
nand U7430 (N_7430,N_5443,N_5647);
xnor U7431 (N_7431,N_5240,N_5811);
or U7432 (N_7432,N_5467,N_4756);
nand U7433 (N_7433,N_4778,N_5806);
or U7434 (N_7434,N_4703,N_4636);
nand U7435 (N_7435,N_5420,N_5923);
and U7436 (N_7436,N_5099,N_4812);
or U7437 (N_7437,N_4632,N_5629);
nand U7438 (N_7438,N_5141,N_5643);
or U7439 (N_7439,N_5092,N_5501);
xnor U7440 (N_7440,N_4734,N_5679);
nor U7441 (N_7441,N_5005,N_5102);
and U7442 (N_7442,N_5474,N_4625);
or U7443 (N_7443,N_5634,N_5020);
and U7444 (N_7444,N_4519,N_4864);
and U7445 (N_7445,N_4584,N_5738);
nor U7446 (N_7446,N_4588,N_5972);
or U7447 (N_7447,N_4791,N_5449);
nor U7448 (N_7448,N_5466,N_5390);
nor U7449 (N_7449,N_5546,N_4746);
nor U7450 (N_7450,N_4553,N_5940);
and U7451 (N_7451,N_5513,N_5719);
nand U7452 (N_7452,N_5152,N_5030);
xnor U7453 (N_7453,N_5587,N_5847);
and U7454 (N_7454,N_4589,N_4864);
and U7455 (N_7455,N_4822,N_5414);
or U7456 (N_7456,N_4939,N_5123);
nor U7457 (N_7457,N_5887,N_4628);
and U7458 (N_7458,N_5866,N_5233);
and U7459 (N_7459,N_5237,N_4684);
nand U7460 (N_7460,N_5914,N_5792);
nand U7461 (N_7461,N_5996,N_4790);
and U7462 (N_7462,N_5766,N_4890);
nor U7463 (N_7463,N_5335,N_5047);
nand U7464 (N_7464,N_4862,N_5678);
nor U7465 (N_7465,N_4601,N_5661);
or U7466 (N_7466,N_5730,N_5834);
and U7467 (N_7467,N_4892,N_4900);
nand U7468 (N_7468,N_5658,N_5477);
or U7469 (N_7469,N_4544,N_4759);
or U7470 (N_7470,N_5616,N_5295);
or U7471 (N_7471,N_5596,N_4856);
nor U7472 (N_7472,N_5265,N_5974);
and U7473 (N_7473,N_5712,N_4861);
nand U7474 (N_7474,N_4875,N_5691);
nand U7475 (N_7475,N_4909,N_5076);
or U7476 (N_7476,N_4689,N_5556);
xnor U7477 (N_7477,N_5461,N_5336);
xor U7478 (N_7478,N_4614,N_5105);
nand U7479 (N_7479,N_5178,N_5372);
or U7480 (N_7480,N_5610,N_4717);
or U7481 (N_7481,N_5753,N_5491);
nand U7482 (N_7482,N_5679,N_5626);
or U7483 (N_7483,N_5784,N_4579);
and U7484 (N_7484,N_5946,N_5724);
nand U7485 (N_7485,N_5651,N_5883);
xnor U7486 (N_7486,N_5362,N_5835);
xnor U7487 (N_7487,N_5723,N_5033);
and U7488 (N_7488,N_5795,N_5578);
nand U7489 (N_7489,N_5372,N_4848);
and U7490 (N_7490,N_4709,N_5357);
nand U7491 (N_7491,N_5346,N_5473);
and U7492 (N_7492,N_5795,N_5227);
or U7493 (N_7493,N_5346,N_5445);
or U7494 (N_7494,N_5619,N_5130);
nor U7495 (N_7495,N_5717,N_4588);
or U7496 (N_7496,N_5221,N_5797);
nand U7497 (N_7497,N_5401,N_5027);
or U7498 (N_7498,N_5394,N_5351);
and U7499 (N_7499,N_4518,N_4769);
nand U7500 (N_7500,N_7241,N_7284);
nand U7501 (N_7501,N_6943,N_6780);
or U7502 (N_7502,N_6912,N_6701);
nand U7503 (N_7503,N_6332,N_6625);
nand U7504 (N_7504,N_6156,N_7297);
or U7505 (N_7505,N_6928,N_6748);
and U7506 (N_7506,N_7039,N_6797);
and U7507 (N_7507,N_6353,N_6955);
or U7508 (N_7508,N_7364,N_6863);
xnor U7509 (N_7509,N_6679,N_6935);
and U7510 (N_7510,N_7132,N_6152);
nor U7511 (N_7511,N_6777,N_7478);
xnor U7512 (N_7512,N_6620,N_7153);
xor U7513 (N_7513,N_6639,N_6967);
nand U7514 (N_7514,N_7386,N_6263);
or U7515 (N_7515,N_6315,N_6136);
or U7516 (N_7516,N_7355,N_7472);
nand U7517 (N_7517,N_6287,N_6997);
nand U7518 (N_7518,N_6779,N_6000);
nand U7519 (N_7519,N_6272,N_6038);
nor U7520 (N_7520,N_7489,N_6586);
nand U7521 (N_7521,N_6426,N_7147);
nand U7522 (N_7522,N_6442,N_7324);
and U7523 (N_7523,N_6305,N_6560);
nand U7524 (N_7524,N_6999,N_6634);
nor U7525 (N_7525,N_7261,N_6514);
nor U7526 (N_7526,N_6933,N_7257);
nand U7527 (N_7527,N_6566,N_6145);
nor U7528 (N_7528,N_6862,N_6150);
nor U7529 (N_7529,N_7378,N_6358);
nand U7530 (N_7530,N_6444,N_6614);
nor U7531 (N_7531,N_7339,N_7363);
xor U7532 (N_7532,N_7067,N_7329);
xor U7533 (N_7533,N_6565,N_6584);
nor U7534 (N_7534,N_6839,N_6941);
or U7535 (N_7535,N_7234,N_6445);
or U7536 (N_7536,N_6237,N_6649);
nor U7537 (N_7537,N_6216,N_7471);
or U7538 (N_7538,N_7317,N_6550);
nand U7539 (N_7539,N_7128,N_6448);
and U7540 (N_7540,N_7189,N_6655);
xnor U7541 (N_7541,N_6926,N_7176);
or U7542 (N_7542,N_7409,N_7418);
or U7543 (N_7543,N_6384,N_6412);
and U7544 (N_7544,N_7008,N_7402);
or U7545 (N_7545,N_6242,N_7233);
nor U7546 (N_7546,N_7042,N_6726);
and U7547 (N_7547,N_6413,N_7025);
and U7548 (N_7548,N_6329,N_6871);
nor U7549 (N_7549,N_7163,N_6306);
and U7550 (N_7550,N_7212,N_7017);
xor U7551 (N_7551,N_6922,N_6212);
and U7552 (N_7552,N_6698,N_6292);
xor U7553 (N_7553,N_6595,N_6446);
nor U7554 (N_7554,N_6690,N_6026);
or U7555 (N_7555,N_7323,N_6399);
nand U7556 (N_7556,N_7426,N_6380);
and U7557 (N_7557,N_6015,N_7051);
nand U7558 (N_7558,N_6506,N_7457);
nor U7559 (N_7559,N_6012,N_6882);
nand U7560 (N_7560,N_7264,N_6916);
nor U7561 (N_7561,N_6682,N_7332);
nor U7562 (N_7562,N_6161,N_6141);
nand U7563 (N_7563,N_6187,N_6864);
xnor U7564 (N_7564,N_6274,N_7031);
and U7565 (N_7565,N_6155,N_6996);
nand U7566 (N_7566,N_6111,N_6061);
or U7567 (N_7567,N_7041,N_6159);
nand U7568 (N_7568,N_6712,N_6393);
nand U7569 (N_7569,N_6563,N_6889);
xor U7570 (N_7570,N_7092,N_6308);
and U7571 (N_7571,N_6110,N_7301);
or U7572 (N_7572,N_7494,N_6206);
and U7573 (N_7573,N_7349,N_7283);
xnor U7574 (N_7574,N_6587,N_7129);
or U7575 (N_7575,N_6376,N_6208);
and U7576 (N_7576,N_7159,N_6958);
xnor U7577 (N_7577,N_7398,N_6536);
or U7578 (N_7578,N_7384,N_7468);
xor U7579 (N_7579,N_7187,N_6017);
or U7580 (N_7580,N_6526,N_6806);
xor U7581 (N_7581,N_7043,N_6720);
nor U7582 (N_7582,N_6593,N_7182);
nand U7583 (N_7583,N_6611,N_7318);
xnor U7584 (N_7584,N_6607,N_6294);
nor U7585 (N_7585,N_7348,N_6387);
or U7586 (N_7586,N_6089,N_7461);
nor U7587 (N_7587,N_7367,N_7145);
and U7588 (N_7588,N_6185,N_6697);
nand U7589 (N_7589,N_6285,N_6995);
nor U7590 (N_7590,N_6092,N_6617);
or U7591 (N_7591,N_6270,N_6240);
or U7592 (N_7592,N_6836,N_6674);
nor U7593 (N_7593,N_7435,N_7298);
or U7594 (N_7594,N_6461,N_7053);
xor U7595 (N_7595,N_7079,N_6386);
nand U7596 (N_7596,N_7020,N_6661);
nor U7597 (N_7597,N_6659,N_7083);
xor U7598 (N_7598,N_7216,N_7424);
or U7599 (N_7599,N_6441,N_7350);
nor U7600 (N_7600,N_7497,N_6428);
xnor U7601 (N_7601,N_6143,N_6355);
xnor U7602 (N_7602,N_6389,N_7123);
or U7603 (N_7603,N_6415,N_6910);
nor U7604 (N_7604,N_6670,N_7203);
or U7605 (N_7605,N_6956,N_6749);
nand U7606 (N_7606,N_7458,N_7266);
xor U7607 (N_7607,N_6673,N_7094);
or U7608 (N_7608,N_6160,N_7440);
xor U7609 (N_7609,N_6282,N_6857);
xor U7610 (N_7610,N_6051,N_7412);
nand U7611 (N_7611,N_6535,N_6660);
or U7612 (N_7612,N_7286,N_7220);
xnor U7613 (N_7613,N_7427,N_7277);
nor U7614 (N_7614,N_7396,N_6072);
xor U7615 (N_7615,N_7267,N_7240);
nor U7616 (N_7616,N_6201,N_6233);
and U7617 (N_7617,N_6788,N_6018);
and U7618 (N_7618,N_6752,N_7148);
nand U7619 (N_7619,N_6744,N_6893);
nand U7620 (N_7620,N_6624,N_6909);
xor U7621 (N_7621,N_6876,N_7316);
xor U7622 (N_7622,N_6490,N_7035);
xnor U7623 (N_7623,N_7195,N_7302);
nand U7624 (N_7624,N_6829,N_6747);
nor U7625 (N_7625,N_6710,N_6957);
and U7626 (N_7626,N_7046,N_6505);
nand U7627 (N_7627,N_7484,N_7099);
xnor U7628 (N_7628,N_7401,N_7109);
nand U7629 (N_7629,N_6293,N_7420);
or U7630 (N_7630,N_7290,N_7078);
or U7631 (N_7631,N_7076,N_7496);
or U7632 (N_7632,N_6359,N_6008);
xor U7633 (N_7633,N_7219,N_6778);
nor U7634 (N_7634,N_7405,N_7107);
nand U7635 (N_7635,N_6078,N_6677);
xor U7636 (N_7636,N_6422,N_7211);
nor U7637 (N_7637,N_6960,N_6613);
and U7638 (N_7638,N_7002,N_7293);
nor U7639 (N_7639,N_7231,N_7103);
xnor U7640 (N_7640,N_6202,N_6232);
and U7641 (N_7641,N_7131,N_7421);
and U7642 (N_7642,N_6036,N_6663);
nor U7643 (N_7643,N_7030,N_6031);
nor U7644 (N_7644,N_7285,N_6372);
xnor U7645 (N_7645,N_7493,N_7397);
xor U7646 (N_7646,N_7395,N_6525);
nor U7647 (N_7647,N_6897,N_7217);
nand U7648 (N_7648,N_6672,N_6148);
and U7649 (N_7649,N_6479,N_6350);
nand U7650 (N_7650,N_6190,N_7436);
xor U7651 (N_7651,N_7001,N_7180);
or U7652 (N_7652,N_6741,N_6388);
xnor U7653 (N_7653,N_6467,N_6680);
and U7654 (N_7654,N_6302,N_7340);
xnor U7655 (N_7655,N_7487,N_6460);
nor U7656 (N_7656,N_6006,N_6654);
nand U7657 (N_7657,N_7313,N_6276);
and U7658 (N_7658,N_6303,N_7089);
or U7659 (N_7659,N_6055,N_7121);
nand U7660 (N_7660,N_7139,N_7080);
xnor U7661 (N_7661,N_7473,N_6553);
and U7662 (N_7662,N_6855,N_7292);
nor U7663 (N_7663,N_7201,N_6980);
xor U7664 (N_7664,N_6895,N_6927);
and U7665 (N_7665,N_7130,N_6675);
or U7666 (N_7666,N_6009,N_6991);
nand U7667 (N_7667,N_6043,N_6239);
xor U7668 (N_7668,N_7353,N_6068);
and U7669 (N_7669,N_7289,N_7245);
and U7670 (N_7670,N_6644,N_7357);
and U7671 (N_7671,N_6377,N_6599);
and U7672 (N_7672,N_6200,N_6794);
nor U7673 (N_7673,N_6178,N_6786);
nand U7674 (N_7674,N_7380,N_6289);
and U7675 (N_7675,N_7024,N_6948);
nor U7676 (N_7676,N_6121,N_6173);
nor U7677 (N_7677,N_6569,N_6301);
nor U7678 (N_7678,N_7171,N_6964);
xor U7679 (N_7679,N_6439,N_6851);
xor U7680 (N_7680,N_7312,N_7173);
and U7681 (N_7681,N_6312,N_6904);
or U7682 (N_7682,N_6795,N_6375);
nor U7683 (N_7683,N_6403,N_7047);
and U7684 (N_7684,N_6600,N_6420);
and U7685 (N_7685,N_6787,N_6635);
nor U7686 (N_7686,N_6382,N_6947);
xnor U7687 (N_7687,N_6222,N_6004);
xnor U7688 (N_7688,N_6572,N_6360);
nor U7689 (N_7689,N_6348,N_6229);
nand U7690 (N_7690,N_6410,N_6543);
nand U7691 (N_7691,N_6279,N_7488);
xor U7692 (N_7692,N_6182,N_6821);
or U7693 (N_7693,N_6087,N_7152);
nand U7694 (N_7694,N_6828,N_6848);
xor U7695 (N_7695,N_6260,N_6491);
or U7696 (N_7696,N_6234,N_7438);
xor U7697 (N_7697,N_6082,N_6404);
and U7698 (N_7698,N_6085,N_6522);
nand U7699 (N_7699,N_6691,N_7413);
or U7700 (N_7700,N_6773,N_7434);
nor U7701 (N_7701,N_7096,N_6913);
xnor U7702 (N_7702,N_7070,N_6715);
or U7703 (N_7703,N_7336,N_6214);
or U7704 (N_7704,N_6062,N_6583);
and U7705 (N_7705,N_6564,N_6860);
and U7706 (N_7706,N_6932,N_7375);
and U7707 (N_7707,N_7122,N_6940);
xnor U7708 (N_7708,N_7135,N_6768);
nor U7709 (N_7709,N_7098,N_7013);
xnor U7710 (N_7710,N_6502,N_6449);
xor U7711 (N_7711,N_6630,N_7144);
nand U7712 (N_7712,N_6891,N_6406);
xor U7713 (N_7713,N_6197,N_6985);
nor U7714 (N_7714,N_6112,N_7104);
and U7715 (N_7715,N_6284,N_6856);
nand U7716 (N_7716,N_6340,N_6322);
nand U7717 (N_7717,N_7015,N_7105);
and U7718 (N_7718,N_6028,N_6556);
and U7719 (N_7719,N_6845,N_7360);
xnor U7720 (N_7720,N_7066,N_7126);
nand U7721 (N_7721,N_7432,N_6215);
or U7722 (N_7722,N_6343,N_6483);
nand U7723 (N_7723,N_6604,N_7115);
xor U7724 (N_7724,N_6310,N_7251);
and U7725 (N_7725,N_6259,N_6924);
xnor U7726 (N_7726,N_6459,N_6045);
or U7727 (N_7727,N_6476,N_6013);
and U7728 (N_7728,N_6896,N_6979);
xnor U7729 (N_7729,N_7419,N_6717);
xor U7730 (N_7730,N_6751,N_7331);
nor U7731 (N_7731,N_7444,N_7101);
or U7732 (N_7732,N_6500,N_6186);
and U7733 (N_7733,N_6135,N_6665);
or U7734 (N_7734,N_6846,N_7300);
nor U7735 (N_7735,N_6369,N_6335);
or U7736 (N_7736,N_7382,N_6057);
and U7737 (N_7737,N_6189,N_7351);
nand U7738 (N_7738,N_7346,N_6849);
xor U7739 (N_7739,N_6261,N_6328);
or U7740 (N_7740,N_6247,N_6198);
xor U7741 (N_7741,N_7417,N_7106);
and U7742 (N_7742,N_6374,N_6314);
nand U7743 (N_7743,N_6154,N_6046);
or U7744 (N_7744,N_7045,N_7344);
and U7745 (N_7745,N_6825,N_7476);
and U7746 (N_7746,N_7372,N_6023);
nor U7747 (N_7747,N_6519,N_7392);
and U7748 (N_7748,N_7307,N_6496);
nand U7749 (N_7749,N_7202,N_6299);
nand U7750 (N_7750,N_6745,N_7177);
and U7751 (N_7751,N_6530,N_6983);
xnor U7752 (N_7752,N_6886,N_6364);
and U7753 (N_7753,N_7385,N_7276);
or U7754 (N_7754,N_6549,N_6923);
and U7755 (N_7755,N_7206,N_6807);
nor U7756 (N_7756,N_6067,N_7456);
nor U7757 (N_7757,N_6188,N_6694);
xor U7758 (N_7758,N_6939,N_7379);
or U7759 (N_7759,N_7425,N_7328);
xor U7760 (N_7760,N_6098,N_6703);
and U7761 (N_7761,N_7222,N_7190);
xnor U7762 (N_7762,N_6936,N_7221);
or U7763 (N_7763,N_6842,N_6758);
nand U7764 (N_7764,N_7063,N_7321);
or U7765 (N_7765,N_6914,N_6395);
nor U7766 (N_7766,N_7061,N_7170);
nand U7767 (N_7767,N_7287,N_7446);
xor U7768 (N_7768,N_7157,N_7465);
xor U7769 (N_7769,N_7183,N_6629);
or U7770 (N_7770,N_6205,N_7125);
or U7771 (N_7771,N_6988,N_7228);
nor U7772 (N_7772,N_6908,N_7081);
and U7773 (N_7773,N_7366,N_6746);
nor U7774 (N_7774,N_6327,N_6433);
and U7775 (N_7775,N_6835,N_6099);
nor U7776 (N_7776,N_6662,N_6107);
nand U7777 (N_7777,N_6493,N_6605);
and U7778 (N_7778,N_6277,N_6396);
nor U7779 (N_7779,N_6424,N_6648);
and U7780 (N_7780,N_6626,N_6298);
xor U7781 (N_7781,N_6094,N_6149);
nor U7782 (N_7782,N_6770,N_6702);
xnor U7783 (N_7783,N_6273,N_6615);
nor U7784 (N_7784,N_6664,N_6341);
and U7785 (N_7785,N_6275,N_7230);
nand U7786 (N_7786,N_7269,N_6256);
xnor U7787 (N_7787,N_7365,N_6852);
xnor U7788 (N_7788,N_6347,N_6511);
nor U7789 (N_7789,N_7012,N_6971);
xnor U7790 (N_7790,N_6077,N_7225);
and U7791 (N_7791,N_6450,N_7477);
and U7792 (N_7792,N_6090,N_6632);
nor U7793 (N_7793,N_6158,N_7389);
xor U7794 (N_7794,N_6733,N_6764);
nor U7795 (N_7795,N_6076,N_7140);
or U7796 (N_7796,N_7482,N_7091);
nand U7797 (N_7797,N_6718,N_7414);
xor U7798 (N_7798,N_7449,N_6316);
nand U7799 (N_7799,N_6575,N_6058);
nand U7800 (N_7800,N_6729,N_6126);
nand U7801 (N_7801,N_6248,N_6527);
nand U7802 (N_7802,N_7021,N_7244);
nand U7803 (N_7803,N_6739,N_6267);
xor U7804 (N_7804,N_6769,N_6693);
xor U7805 (N_7805,N_6812,N_7475);
or U7806 (N_7806,N_6978,N_6561);
xnor U7807 (N_7807,N_6066,N_7454);
xnor U7808 (N_7808,N_6040,N_6668);
and U7809 (N_7809,N_6095,N_6290);
and U7810 (N_7810,N_6492,N_7032);
nand U7811 (N_7811,N_6088,N_7097);
xor U7812 (N_7812,N_7004,N_7028);
and U7813 (N_7813,N_6165,N_6005);
or U7814 (N_7814,N_7085,N_6934);
nor U7815 (N_7815,N_6554,N_7167);
and U7816 (N_7816,N_6790,N_6859);
or U7817 (N_7817,N_6551,N_6438);
nand U7818 (N_7818,N_6603,N_6056);
xor U7819 (N_7819,N_6570,N_6942);
nor U7820 (N_7820,N_6532,N_6974);
nor U7821 (N_7821,N_6972,N_6059);
nor U7822 (N_7822,N_6765,N_7445);
and U7823 (N_7823,N_6650,N_7304);
or U7824 (N_7824,N_6249,N_7007);
nand U7825 (N_7825,N_7467,N_7439);
and U7826 (N_7826,N_6809,N_6894);
and U7827 (N_7827,N_6722,N_7305);
or U7828 (N_7828,N_7410,N_7407);
xnor U7829 (N_7829,N_7188,N_6900);
nand U7830 (N_7830,N_6499,N_7010);
and U7831 (N_7831,N_6982,N_7299);
nor U7832 (N_7832,N_6645,N_6544);
nor U7833 (N_7833,N_6919,N_6833);
nor U7834 (N_7834,N_7451,N_6497);
nand U7835 (N_7835,N_6831,N_7003);
xor U7836 (N_7836,N_6488,N_6647);
and U7837 (N_7837,N_6481,N_6138);
and U7838 (N_7838,N_6203,N_6890);
and U7839 (N_7839,N_6324,N_6478);
and U7840 (N_7840,N_7242,N_6961);
or U7841 (N_7841,N_7431,N_6808);
nand U7842 (N_7842,N_6101,N_6993);
xnor U7843 (N_7843,N_6885,N_6541);
and U7844 (N_7844,N_7019,N_6137);
and U7845 (N_7845,N_7275,N_7270);
xor U7846 (N_7846,N_6952,N_6280);
and U7847 (N_7847,N_6884,N_6122);
and U7848 (N_7848,N_6534,N_6039);
xor U7849 (N_7849,N_6021,N_6401);
nor U7850 (N_7850,N_6796,N_6210);
nand U7851 (N_7851,N_7210,N_6798);
and U7852 (N_7852,N_7200,N_7345);
nor U7853 (N_7853,N_6054,N_6177);
or U7854 (N_7854,N_6437,N_6432);
and U7855 (N_7855,N_7227,N_6255);
and U7856 (N_7856,N_6981,N_6108);
nor U7857 (N_7857,N_6041,N_6288);
nand U7858 (N_7858,N_7388,N_7483);
xnor U7859 (N_7859,N_6162,N_6368);
and U7860 (N_7860,N_6470,N_7162);
nand U7861 (N_7861,N_7358,N_6547);
or U7862 (N_7862,N_6898,N_6167);
xor U7863 (N_7863,N_6042,N_7026);
nor U7864 (N_7864,N_6431,N_6238);
xor U7865 (N_7865,N_7082,N_6120);
nor U7866 (N_7866,N_6567,N_6592);
nand U7867 (N_7867,N_7306,N_6989);
nand U7868 (N_7868,N_6881,N_6349);
or U7869 (N_7869,N_6568,N_6392);
or U7870 (N_7870,N_6002,N_6477);
xor U7871 (N_7871,N_6475,N_7214);
or U7872 (N_7872,N_6727,N_7430);
xor U7873 (N_7873,N_6192,N_6228);
or U7874 (N_7874,N_7387,N_6218);
or U7875 (N_7875,N_7172,N_7423);
nor U7876 (N_7876,N_6854,N_7156);
xor U7877 (N_7877,N_7119,N_6827);
or U7878 (N_7878,N_7110,N_6669);
nor U7879 (N_7879,N_6196,N_7209);
nor U7880 (N_7880,N_6576,N_7006);
and U7881 (N_7881,N_6016,N_6509);
nand U7882 (N_7882,N_7199,N_7460);
xor U7883 (N_7883,N_7394,N_6489);
nand U7884 (N_7884,N_7429,N_6540);
xnor U7885 (N_7885,N_6434,N_6986);
nand U7886 (N_7886,N_7086,N_7247);
nand U7887 (N_7887,N_7178,N_7433);
nand U7888 (N_7888,N_6458,N_6562);
nor U7889 (N_7889,N_6383,N_7250);
xnor U7890 (N_7890,N_6453,N_6221);
xor U7891 (N_7891,N_6671,N_6373);
and U7892 (N_7892,N_6994,N_6048);
and U7893 (N_7893,N_6105,N_7498);
or U7894 (N_7894,N_6619,N_6436);
nor U7895 (N_7895,N_6883,N_6264);
nor U7896 (N_7896,N_6657,N_6140);
and U7897 (N_7897,N_7033,N_6804);
and U7898 (N_7898,N_6774,N_6319);
nand U7899 (N_7899,N_6555,N_6802);
or U7900 (N_7900,N_7411,N_7055);
or U7901 (N_7901,N_7160,N_7111);
nand U7902 (N_7902,N_6738,N_6115);
nand U7903 (N_7903,N_7093,N_6507);
xnor U7904 (N_7904,N_7356,N_6822);
xnor U7905 (N_7905,N_6269,N_6086);
and U7906 (N_7906,N_7391,N_6874);
or U7907 (N_7907,N_6868,N_6516);
nor U7908 (N_7908,N_6937,N_6810);
xnor U7909 (N_7909,N_6905,N_6705);
and U7910 (N_7910,N_6361,N_7037);
nor U7911 (N_7911,N_7334,N_7179);
nand U7912 (N_7912,N_6296,N_6861);
or U7913 (N_7913,N_6456,N_6119);
or U7914 (N_7914,N_7065,N_7490);
and U7915 (N_7915,N_6468,N_7260);
nand U7916 (N_7916,N_7208,N_7022);
nor U7917 (N_7917,N_6799,N_6642);
and U7918 (N_7918,N_7124,N_6024);
or U7919 (N_7919,N_7265,N_6918);
nor U7920 (N_7920,N_7184,N_6538);
xor U7921 (N_7921,N_6211,N_6146);
and U7922 (N_7922,N_7237,N_6951);
and U7923 (N_7923,N_6742,N_7044);
and U7924 (N_7924,N_6371,N_6784);
nand U7925 (N_7925,N_6331,N_6899);
or U7926 (N_7926,N_6966,N_7064);
xor U7927 (N_7927,N_7133,N_6266);
and U7928 (N_7928,N_6225,N_7165);
and U7929 (N_7929,N_6447,N_7034);
nand U7930 (N_7930,N_7263,N_6580);
xor U7931 (N_7931,N_6931,N_7343);
nand U7932 (N_7932,N_6130,N_7278);
nand U7933 (N_7933,N_6651,N_6391);
nand U7934 (N_7934,N_6394,N_6019);
or U7935 (N_7935,N_6060,N_7117);
nor U7936 (N_7936,N_6243,N_6637);
or U7937 (N_7937,N_7474,N_7112);
xnor U7938 (N_7938,N_6713,N_6176);
nand U7939 (N_7939,N_6053,N_6142);
nand U7940 (N_7940,N_7174,N_7224);
and U7941 (N_7941,N_6528,N_6052);
and U7942 (N_7942,N_6628,N_6723);
nand U7943 (N_7943,N_6397,N_6171);
xnor U7944 (N_7944,N_7327,N_6954);
nand U7945 (N_7945,N_6344,N_6872);
xor U7946 (N_7946,N_6124,N_7437);
nor U7947 (N_7947,N_6291,N_7262);
nor U7948 (N_7948,N_6602,N_6826);
xnor U7949 (N_7949,N_6724,N_7072);
xor U7950 (N_7950,N_7151,N_6612);
and U7951 (N_7951,N_6144,N_7271);
or U7952 (N_7952,N_6464,N_6084);
or U7953 (N_7953,N_6945,N_7062);
nand U7954 (N_7954,N_7400,N_7056);
xor U7955 (N_7955,N_6756,N_6984);
xnor U7956 (N_7956,N_7492,N_7050);
xor U7957 (N_7957,N_6585,N_6027);
nand U7958 (N_7958,N_6257,N_6622);
nand U7959 (N_7959,N_7114,N_6887);
nand U7960 (N_7960,N_6323,N_6850);
nor U7961 (N_7961,N_6153,N_6352);
xor U7962 (N_7962,N_6325,N_6838);
and U7963 (N_7963,N_6174,N_7068);
nor U7964 (N_7964,N_7408,N_6987);
nand U7965 (N_7965,N_6181,N_6782);
and U7966 (N_7966,N_7038,N_7254);
and U7967 (N_7967,N_7404,N_7027);
nor U7968 (N_7968,N_6416,N_6684);
nor U7969 (N_7969,N_6638,N_6793);
nand U7970 (N_7970,N_7374,N_6337);
and U7971 (N_7971,N_6901,N_6097);
nand U7972 (N_7972,N_6049,N_6381);
or U7973 (N_7973,N_6102,N_6252);
nor U7974 (N_7974,N_6735,N_6351);
and U7975 (N_7975,N_6022,N_6763);
or U7976 (N_7976,N_6354,N_6253);
nand U7977 (N_7977,N_7088,N_6877);
or U7978 (N_7978,N_6646,N_6977);
xnor U7979 (N_7979,N_6096,N_6903);
or U7980 (N_7980,N_6035,N_6163);
or U7981 (N_7981,N_6818,N_6241);
nor U7982 (N_7982,N_6195,N_7294);
or U7983 (N_7983,N_6959,N_6640);
nand U7984 (N_7984,N_6334,N_6429);
nand U7985 (N_7985,N_6064,N_6254);
nand U7986 (N_7986,N_7463,N_7466);
nor U7987 (N_7987,N_6003,N_6740);
xnor U7988 (N_7988,N_6820,N_6685);
or U7989 (N_7989,N_7095,N_7282);
xor U7990 (N_7990,N_6695,N_7369);
or U7991 (N_7991,N_6631,N_6508);
or U7992 (N_7992,N_6091,N_6678);
or U7993 (N_7993,N_7090,N_6071);
and U7994 (N_7994,N_7383,N_6573);
or U7995 (N_7995,N_6771,N_6616);
and U7996 (N_7996,N_6609,N_6743);
nor U7997 (N_7997,N_7149,N_6366);
or U7998 (N_7998,N_7373,N_6157);
nand U7999 (N_7999,N_7014,N_6326);
nand U8000 (N_8000,N_6220,N_6025);
xor U8001 (N_8001,N_6462,N_6962);
nand U8002 (N_8002,N_6805,N_6251);
nor U8003 (N_8003,N_7071,N_7175);
and U8004 (N_8004,N_6286,N_7141);
nand U8005 (N_8005,N_6571,N_6976);
or U8006 (N_8006,N_6558,N_6731);
nand U8007 (N_8007,N_7281,N_7040);
or U8008 (N_8008,N_6081,N_6125);
nand U8009 (N_8009,N_6531,N_7102);
and U8010 (N_8010,N_6762,N_6168);
or U8011 (N_8011,N_6400,N_6134);
nand U8012 (N_8012,N_7322,N_6521);
nor U8013 (N_8013,N_6074,N_6482);
or U8014 (N_8014,N_6409,N_7223);
or U8015 (N_8015,N_6070,N_6953);
nor U8016 (N_8016,N_6339,N_7415);
nand U8017 (N_8017,N_6606,N_6915);
and U8018 (N_8018,N_6235,N_7049);
xor U8019 (N_8019,N_7295,N_6892);
nand U8020 (N_8020,N_6425,N_6610);
or U8021 (N_8021,N_6658,N_6517);
xor U8022 (N_8022,N_6398,N_6969);
or U8023 (N_8023,N_6594,N_7361);
nand U8024 (N_8024,N_6073,N_6333);
nand U8025 (N_8025,N_6676,N_6485);
or U8026 (N_8026,N_6484,N_6529);
nand U8027 (N_8027,N_6133,N_6283);
nor U8028 (N_8028,N_7016,N_7333);
nor U8029 (N_8029,N_6407,N_6116);
nand U8030 (N_8030,N_6421,N_6451);
and U8031 (N_8031,N_7146,N_6775);
nand U8032 (N_8032,N_6865,N_6643);
nand U8033 (N_8033,N_6250,N_6653);
nand U8034 (N_8034,N_6817,N_6330);
and U8035 (N_8035,N_7168,N_7194);
nand U8036 (N_8036,N_6824,N_7288);
nor U8037 (N_8037,N_6750,N_6963);
and U8038 (N_8038,N_7243,N_7084);
and U8039 (N_8039,N_6213,N_6103);
nand U8040 (N_8040,N_7314,N_6047);
and U8041 (N_8041,N_7253,N_7207);
xor U8042 (N_8042,N_7155,N_7142);
nand U8043 (N_8043,N_7226,N_7310);
and U8044 (N_8044,N_7268,N_6714);
xor U8045 (N_8045,N_6781,N_6472);
or U8046 (N_8046,N_6811,N_6510);
or U8047 (N_8047,N_7136,N_6069);
nor U8048 (N_8048,N_6970,N_6975);
nand U8049 (N_8049,N_7249,N_6548);
or U8050 (N_8050,N_7341,N_7005);
nand U8051 (N_8051,N_7118,N_6577);
or U8052 (N_8052,N_7443,N_7320);
nor U8053 (N_8053,N_6075,N_6297);
and U8054 (N_8054,N_6408,N_7197);
or U8055 (N_8055,N_6853,N_7428);
or U8056 (N_8056,N_7393,N_6687);
and U8057 (N_8057,N_6414,N_7073);
nand U8058 (N_8058,N_7074,N_7169);
and U8059 (N_8059,N_6029,N_6180);
and U8060 (N_8060,N_6362,N_6357);
and U8061 (N_8061,N_6440,N_6118);
and U8062 (N_8062,N_6737,N_7138);
or U8063 (N_8063,N_7422,N_6621);
xnor U8064 (N_8064,N_6929,N_6487);
nand U8065 (N_8065,N_6601,N_7485);
and U8066 (N_8066,N_6378,N_6716);
or U8067 (N_8067,N_7347,N_6656);
and U8068 (N_8068,N_6032,N_6385);
nor U8069 (N_8069,N_7403,N_7335);
or U8070 (N_8070,N_6998,N_6533);
nor U8071 (N_8071,N_6618,N_7143);
or U8072 (N_8072,N_6707,N_6405);
xor U8073 (N_8073,N_6443,N_6245);
nor U8074 (N_8074,N_7459,N_7057);
or U8075 (N_8075,N_6258,N_6231);
and U8076 (N_8076,N_6992,N_6813);
nor U8077 (N_8077,N_6494,N_7303);
and U8078 (N_8078,N_7127,N_6114);
and U8079 (N_8079,N_6199,N_7354);
nor U8080 (N_8080,N_6512,N_7376);
nand U8081 (N_8081,N_7377,N_6574);
nor U8082 (N_8082,N_7469,N_7235);
and U8083 (N_8083,N_6840,N_6520);
or U8084 (N_8084,N_7442,N_6623);
and U8085 (N_8085,N_6719,N_6641);
nor U8086 (N_8086,N_6345,N_7259);
and U8087 (N_8087,N_6834,N_6706);
nor U8088 (N_8088,N_6106,N_7150);
and U8089 (N_8089,N_6147,N_6318);
and U8090 (N_8090,N_7499,N_6503);
xor U8091 (N_8091,N_6132,N_7447);
and U8092 (N_8092,N_6129,N_7196);
or U8093 (N_8093,N_6244,N_7246);
nor U8094 (N_8094,N_7311,N_7054);
nor U8095 (N_8095,N_6906,N_6065);
xor U8096 (N_8096,N_6968,N_6873);
or U8097 (N_8097,N_6093,N_7308);
and U8098 (N_8098,N_6471,N_6816);
nor U8099 (N_8099,N_7452,N_6858);
nor U8100 (N_8100,N_7325,N_7256);
or U8101 (N_8101,N_6837,N_6841);
xor U8102 (N_8102,N_6486,N_6427);
or U8103 (N_8103,N_6342,N_6011);
xnor U8104 (N_8104,N_6815,N_6474);
xnor U8105 (N_8105,N_6792,N_6226);
or U8106 (N_8106,N_6755,N_6832);
nand U8107 (N_8107,N_6965,N_6721);
nor U8108 (N_8108,N_6597,N_6455);
nand U8109 (N_8109,N_6539,N_6552);
nand U8110 (N_8110,N_7338,N_7018);
nor U8111 (N_8111,N_6686,N_6204);
xnor U8112 (N_8112,N_6652,N_7448);
nor U8113 (N_8113,N_7279,N_7462);
nor U8114 (N_8114,N_7069,N_7370);
and U8115 (N_8115,N_7291,N_6732);
nor U8116 (N_8116,N_6917,N_6219);
or U8117 (N_8117,N_7029,N_7108);
nand U8118 (N_8118,N_6498,N_6435);
nor U8119 (N_8119,N_6271,N_7048);
nand U8120 (N_8120,N_6800,N_7406);
or U8121 (N_8121,N_6504,N_7450);
and U8122 (N_8122,N_7239,N_6417);
or U8123 (N_8123,N_6911,N_6708);
or U8124 (N_8124,N_6757,N_7273);
and U8125 (N_8125,N_7023,N_6920);
xnor U8126 (N_8126,N_6546,N_6224);
xnor U8127 (N_8127,N_7193,N_7232);
and U8128 (N_8128,N_7164,N_7296);
xor U8129 (N_8129,N_7238,N_7315);
nand U8130 (N_8130,N_6184,N_7058);
or U8131 (N_8131,N_6457,N_6246);
nand U8132 (N_8132,N_6633,N_7464);
and U8133 (N_8133,N_7186,N_6175);
xor U8134 (N_8134,N_6379,N_6080);
xor U8135 (N_8135,N_7455,N_6791);
or U8136 (N_8136,N_7154,N_7453);
nor U8137 (N_8137,N_6495,N_7100);
nand U8138 (N_8138,N_6007,N_6050);
and U8139 (N_8139,N_6700,N_6880);
nand U8140 (N_8140,N_6309,N_6079);
xnor U8141 (N_8141,N_7052,N_6627);
nand U8142 (N_8142,N_6030,N_6411);
and U8143 (N_8143,N_6390,N_6930);
nand U8144 (N_8144,N_6501,N_6524);
or U8145 (N_8145,N_6636,N_6194);
xor U8146 (N_8146,N_6867,N_6589);
xnor U8147 (N_8147,N_7486,N_6365);
or U8148 (N_8148,N_7192,N_7441);
nand U8149 (N_8149,N_7274,N_7229);
nor U8150 (N_8150,N_6725,N_7280);
or U8151 (N_8151,N_6803,N_6320);
nand U8152 (N_8152,N_6127,N_6513);
xor U8153 (N_8153,N_6033,N_6191);
or U8154 (N_8154,N_7036,N_7236);
nand U8155 (N_8155,N_6217,N_6973);
xor U8156 (N_8156,N_7060,N_7000);
and U8157 (N_8157,N_7185,N_7213);
nand U8158 (N_8158,N_6172,N_6356);
and U8159 (N_8159,N_7258,N_7359);
or U8160 (N_8160,N_6588,N_6537);
nand U8161 (N_8161,N_6783,N_6465);
or U8162 (N_8162,N_6166,N_7352);
and U8163 (N_8163,N_6902,N_6262);
nor U8164 (N_8164,N_7481,N_6317);
or U8165 (N_8165,N_6591,N_6515);
nor U8166 (N_8166,N_6169,N_6430);
or U8167 (N_8167,N_7120,N_7137);
or U8168 (N_8168,N_6295,N_6949);
nand U8169 (N_8169,N_6579,N_6418);
nand U8170 (N_8170,N_6300,N_6946);
nor U8171 (N_8171,N_6230,N_6469);
nand U8172 (N_8172,N_6598,N_6688);
nand U8173 (N_8173,N_6338,N_7134);
or U8174 (N_8174,N_6776,N_6480);
nand U8175 (N_8175,N_7330,N_6034);
or U8176 (N_8176,N_7113,N_6128);
nand U8177 (N_8177,N_6582,N_6814);
xor U8178 (N_8178,N_6151,N_6104);
nor U8179 (N_8179,N_6419,N_6875);
or U8180 (N_8180,N_6704,N_6866);
nor U8181 (N_8181,N_6754,N_7166);
or U8182 (N_8182,N_6037,N_7191);
nor U8183 (N_8183,N_6759,N_6921);
and U8184 (N_8184,N_6423,N_6123);
or U8185 (N_8185,N_6596,N_7011);
and U8186 (N_8186,N_6117,N_6692);
xnor U8187 (N_8187,N_6304,N_7215);
and U8188 (N_8188,N_7252,N_7390);
or U8189 (N_8189,N_6131,N_6063);
nand U8190 (N_8190,N_6728,N_6044);
nand U8191 (N_8191,N_6281,N_7470);
or U8192 (N_8192,N_6209,N_6321);
or U8193 (N_8193,N_6268,N_6020);
or U8194 (N_8194,N_6083,N_6311);
xor U8195 (N_8195,N_6709,N_7059);
or U8196 (N_8196,N_6518,N_7326);
or U8197 (N_8197,N_6193,N_6523);
and U8198 (N_8198,N_6753,N_7248);
or U8199 (N_8199,N_7371,N_6336);
and U8200 (N_8200,N_6681,N_7479);
or U8201 (N_8201,N_6109,N_6870);
xor U8202 (N_8202,N_6760,N_6466);
nand U8203 (N_8203,N_6363,N_6236);
xnor U8204 (N_8204,N_6183,N_6869);
nor U8205 (N_8205,N_7009,N_6878);
xnor U8206 (N_8206,N_6761,N_7368);
xor U8207 (N_8207,N_6581,N_6265);
nor U8208 (N_8208,N_6683,N_6767);
and U8209 (N_8209,N_7218,N_6844);
nor U8210 (N_8210,N_7255,N_7204);
or U8211 (N_8211,N_6463,N_6843);
and U8212 (N_8212,N_6734,N_6667);
or U8213 (N_8213,N_7272,N_6847);
or U8214 (N_8214,N_6950,N_6801);
or U8215 (N_8215,N_6278,N_6938);
xor U8216 (N_8216,N_6010,N_7399);
xnor U8217 (N_8217,N_6207,N_7075);
or U8218 (N_8218,N_7087,N_6907);
xor U8219 (N_8219,N_6307,N_6164);
xnor U8220 (N_8220,N_6823,N_6578);
nor U8221 (N_8221,N_7362,N_7416);
xnor U8222 (N_8222,N_6001,N_6370);
xor U8223 (N_8223,N_7491,N_7205);
or U8224 (N_8224,N_7309,N_6789);
xnor U8225 (N_8225,N_6608,N_6179);
and U8226 (N_8226,N_7480,N_6730);
nor U8227 (N_8227,N_6402,N_7158);
and U8228 (N_8228,N_7116,N_6772);
xor U8229 (N_8229,N_6113,N_6545);
and U8230 (N_8230,N_6139,N_6100);
nor U8231 (N_8231,N_6711,N_6766);
nand U8232 (N_8232,N_6879,N_7198);
nor U8233 (N_8233,N_6696,N_6830);
xor U8234 (N_8234,N_6223,N_6944);
and U8235 (N_8235,N_7077,N_6699);
or U8236 (N_8236,N_6666,N_7319);
nand U8237 (N_8237,N_6313,N_6542);
or U8238 (N_8238,N_7337,N_6785);
or U8239 (N_8239,N_6819,N_6888);
nor U8240 (N_8240,N_6454,N_7381);
nor U8241 (N_8241,N_7161,N_6367);
and U8242 (N_8242,N_7342,N_6227);
nor U8243 (N_8243,N_6925,N_6990);
or U8244 (N_8244,N_6170,N_6590);
nand U8245 (N_8245,N_6689,N_6346);
and U8246 (N_8246,N_7495,N_6559);
nor U8247 (N_8247,N_6473,N_6452);
and U8248 (N_8248,N_7181,N_6736);
xor U8249 (N_8249,N_6014,N_6557);
nand U8250 (N_8250,N_6341,N_6311);
nor U8251 (N_8251,N_6187,N_6156);
nand U8252 (N_8252,N_6792,N_7235);
nand U8253 (N_8253,N_6396,N_6926);
or U8254 (N_8254,N_6432,N_6365);
nand U8255 (N_8255,N_6362,N_6026);
nand U8256 (N_8256,N_6131,N_6434);
nor U8257 (N_8257,N_6838,N_7386);
nand U8258 (N_8258,N_6950,N_7128);
xor U8259 (N_8259,N_6681,N_6782);
xor U8260 (N_8260,N_7296,N_6992);
xnor U8261 (N_8261,N_7280,N_6096);
or U8262 (N_8262,N_6919,N_6004);
xor U8263 (N_8263,N_7108,N_7447);
nand U8264 (N_8264,N_6877,N_7470);
nand U8265 (N_8265,N_6297,N_6723);
nand U8266 (N_8266,N_6941,N_7072);
xnor U8267 (N_8267,N_6775,N_7371);
xnor U8268 (N_8268,N_7489,N_6205);
nor U8269 (N_8269,N_7084,N_6767);
nor U8270 (N_8270,N_7183,N_6946);
nor U8271 (N_8271,N_6921,N_6559);
nand U8272 (N_8272,N_6523,N_6980);
nand U8273 (N_8273,N_7314,N_6989);
nor U8274 (N_8274,N_6010,N_7093);
or U8275 (N_8275,N_6923,N_6369);
nor U8276 (N_8276,N_7361,N_7413);
and U8277 (N_8277,N_7318,N_6916);
nor U8278 (N_8278,N_7328,N_6282);
xor U8279 (N_8279,N_6639,N_6554);
nand U8280 (N_8280,N_6194,N_7262);
or U8281 (N_8281,N_7069,N_6420);
nor U8282 (N_8282,N_6437,N_6543);
xnor U8283 (N_8283,N_7072,N_6256);
nor U8284 (N_8284,N_7125,N_6085);
nand U8285 (N_8285,N_7268,N_6850);
xor U8286 (N_8286,N_6029,N_6387);
nand U8287 (N_8287,N_6170,N_7489);
xor U8288 (N_8288,N_7322,N_6796);
and U8289 (N_8289,N_6410,N_6425);
nor U8290 (N_8290,N_6921,N_7473);
nor U8291 (N_8291,N_6501,N_6487);
xnor U8292 (N_8292,N_6132,N_6732);
and U8293 (N_8293,N_6268,N_7460);
xor U8294 (N_8294,N_6956,N_6132);
nor U8295 (N_8295,N_6203,N_6036);
and U8296 (N_8296,N_6928,N_6025);
or U8297 (N_8297,N_6412,N_6047);
nand U8298 (N_8298,N_7404,N_6137);
or U8299 (N_8299,N_6562,N_6281);
nand U8300 (N_8300,N_6805,N_6097);
nand U8301 (N_8301,N_6002,N_6493);
xor U8302 (N_8302,N_6119,N_6555);
xnor U8303 (N_8303,N_6990,N_6500);
and U8304 (N_8304,N_6342,N_7079);
and U8305 (N_8305,N_6055,N_7362);
nand U8306 (N_8306,N_6779,N_7065);
nor U8307 (N_8307,N_6011,N_6620);
xnor U8308 (N_8308,N_6181,N_7418);
and U8309 (N_8309,N_6660,N_6172);
and U8310 (N_8310,N_6457,N_6760);
or U8311 (N_8311,N_6442,N_6506);
nor U8312 (N_8312,N_6301,N_7325);
nand U8313 (N_8313,N_6997,N_6922);
nor U8314 (N_8314,N_6509,N_7292);
nand U8315 (N_8315,N_6098,N_7164);
xor U8316 (N_8316,N_7406,N_7196);
and U8317 (N_8317,N_6370,N_6484);
and U8318 (N_8318,N_7415,N_6532);
and U8319 (N_8319,N_6885,N_6728);
nand U8320 (N_8320,N_7258,N_6142);
nor U8321 (N_8321,N_7495,N_6472);
nor U8322 (N_8322,N_6285,N_7368);
nor U8323 (N_8323,N_7083,N_7477);
and U8324 (N_8324,N_6900,N_6877);
and U8325 (N_8325,N_6499,N_7090);
nand U8326 (N_8326,N_6579,N_7457);
nand U8327 (N_8327,N_6189,N_6747);
and U8328 (N_8328,N_7086,N_7178);
xnor U8329 (N_8329,N_6850,N_7067);
xnor U8330 (N_8330,N_7151,N_7481);
nor U8331 (N_8331,N_6177,N_7181);
or U8332 (N_8332,N_6705,N_7020);
or U8333 (N_8333,N_6114,N_6673);
nor U8334 (N_8334,N_7323,N_7486);
nand U8335 (N_8335,N_6641,N_6570);
or U8336 (N_8336,N_6122,N_6451);
nand U8337 (N_8337,N_6414,N_6808);
nand U8338 (N_8338,N_6246,N_6437);
and U8339 (N_8339,N_7264,N_6198);
xor U8340 (N_8340,N_7404,N_7043);
or U8341 (N_8341,N_7223,N_6351);
nand U8342 (N_8342,N_6224,N_6333);
nand U8343 (N_8343,N_6826,N_6622);
or U8344 (N_8344,N_7184,N_6696);
and U8345 (N_8345,N_7070,N_7470);
nor U8346 (N_8346,N_6800,N_7492);
xnor U8347 (N_8347,N_7150,N_6355);
or U8348 (N_8348,N_7429,N_6883);
nor U8349 (N_8349,N_6040,N_6574);
or U8350 (N_8350,N_6513,N_6909);
xor U8351 (N_8351,N_6168,N_6825);
xnor U8352 (N_8352,N_6494,N_7416);
nor U8353 (N_8353,N_7314,N_6568);
nor U8354 (N_8354,N_6902,N_7302);
nor U8355 (N_8355,N_7127,N_7334);
nand U8356 (N_8356,N_7168,N_7285);
xnor U8357 (N_8357,N_6608,N_7244);
xor U8358 (N_8358,N_6922,N_6171);
nand U8359 (N_8359,N_7117,N_6107);
nand U8360 (N_8360,N_6928,N_7099);
or U8361 (N_8361,N_7130,N_6359);
or U8362 (N_8362,N_6629,N_6711);
nand U8363 (N_8363,N_6131,N_6466);
and U8364 (N_8364,N_6753,N_6796);
and U8365 (N_8365,N_6806,N_7346);
nor U8366 (N_8366,N_7105,N_6746);
and U8367 (N_8367,N_6512,N_6263);
and U8368 (N_8368,N_6805,N_7044);
nor U8369 (N_8369,N_7237,N_6423);
xor U8370 (N_8370,N_6270,N_6384);
nand U8371 (N_8371,N_6966,N_6628);
xnor U8372 (N_8372,N_7319,N_6268);
nor U8373 (N_8373,N_6041,N_7432);
nand U8374 (N_8374,N_6409,N_7373);
or U8375 (N_8375,N_7173,N_6057);
or U8376 (N_8376,N_7238,N_6977);
xnor U8377 (N_8377,N_7313,N_6973);
xor U8378 (N_8378,N_7000,N_6805);
nand U8379 (N_8379,N_7457,N_6729);
and U8380 (N_8380,N_7331,N_6840);
and U8381 (N_8381,N_6283,N_6400);
nor U8382 (N_8382,N_7187,N_6290);
and U8383 (N_8383,N_6881,N_6700);
nand U8384 (N_8384,N_7257,N_7447);
nand U8385 (N_8385,N_7158,N_6622);
or U8386 (N_8386,N_6912,N_6422);
nand U8387 (N_8387,N_7453,N_6489);
xor U8388 (N_8388,N_6611,N_6234);
or U8389 (N_8389,N_6851,N_7273);
nand U8390 (N_8390,N_7008,N_6285);
and U8391 (N_8391,N_6313,N_6890);
nor U8392 (N_8392,N_7038,N_7319);
nand U8393 (N_8393,N_7272,N_7284);
nor U8394 (N_8394,N_6654,N_6729);
xor U8395 (N_8395,N_6078,N_6121);
nor U8396 (N_8396,N_6892,N_6391);
or U8397 (N_8397,N_7260,N_6333);
and U8398 (N_8398,N_6388,N_6408);
or U8399 (N_8399,N_6607,N_6817);
nor U8400 (N_8400,N_6925,N_6216);
nor U8401 (N_8401,N_6502,N_6187);
and U8402 (N_8402,N_6795,N_6675);
xnor U8403 (N_8403,N_7355,N_6361);
nor U8404 (N_8404,N_6255,N_7332);
nor U8405 (N_8405,N_6918,N_6925);
nor U8406 (N_8406,N_6590,N_6369);
nor U8407 (N_8407,N_6324,N_6343);
xor U8408 (N_8408,N_6989,N_6043);
or U8409 (N_8409,N_6932,N_6627);
and U8410 (N_8410,N_6977,N_7160);
or U8411 (N_8411,N_6203,N_6384);
xor U8412 (N_8412,N_6997,N_6513);
nand U8413 (N_8413,N_6266,N_7351);
nand U8414 (N_8414,N_6885,N_6952);
and U8415 (N_8415,N_7481,N_7081);
nor U8416 (N_8416,N_7278,N_6498);
and U8417 (N_8417,N_7494,N_7242);
and U8418 (N_8418,N_6641,N_6286);
xnor U8419 (N_8419,N_7184,N_6353);
and U8420 (N_8420,N_7316,N_6330);
and U8421 (N_8421,N_6452,N_7393);
or U8422 (N_8422,N_6392,N_6100);
nand U8423 (N_8423,N_7350,N_6880);
nor U8424 (N_8424,N_6805,N_6265);
nand U8425 (N_8425,N_6890,N_7330);
xnor U8426 (N_8426,N_7343,N_6630);
or U8427 (N_8427,N_6220,N_6785);
or U8428 (N_8428,N_7159,N_6166);
and U8429 (N_8429,N_6012,N_7373);
and U8430 (N_8430,N_7165,N_6527);
or U8431 (N_8431,N_6646,N_6366);
xor U8432 (N_8432,N_6318,N_6822);
or U8433 (N_8433,N_7027,N_7479);
nor U8434 (N_8434,N_6238,N_7051);
and U8435 (N_8435,N_7211,N_6101);
or U8436 (N_8436,N_6758,N_7469);
and U8437 (N_8437,N_6326,N_6944);
nand U8438 (N_8438,N_6049,N_7420);
and U8439 (N_8439,N_7366,N_7000);
nand U8440 (N_8440,N_7326,N_7481);
nor U8441 (N_8441,N_7152,N_6891);
xor U8442 (N_8442,N_6682,N_6894);
nor U8443 (N_8443,N_6756,N_6433);
or U8444 (N_8444,N_7091,N_6539);
xnor U8445 (N_8445,N_6858,N_6494);
and U8446 (N_8446,N_7087,N_7422);
and U8447 (N_8447,N_6934,N_6938);
nor U8448 (N_8448,N_7310,N_6357);
or U8449 (N_8449,N_6207,N_6867);
xor U8450 (N_8450,N_6732,N_6183);
nor U8451 (N_8451,N_7101,N_7378);
nor U8452 (N_8452,N_6880,N_7305);
and U8453 (N_8453,N_6697,N_6961);
and U8454 (N_8454,N_6012,N_6231);
xor U8455 (N_8455,N_6307,N_6448);
nand U8456 (N_8456,N_6195,N_6316);
nor U8457 (N_8457,N_6493,N_6974);
nand U8458 (N_8458,N_7258,N_6522);
xor U8459 (N_8459,N_6316,N_7002);
nand U8460 (N_8460,N_6139,N_6067);
nand U8461 (N_8461,N_7221,N_6519);
nor U8462 (N_8462,N_7161,N_7348);
nand U8463 (N_8463,N_7462,N_6727);
xor U8464 (N_8464,N_6295,N_6873);
or U8465 (N_8465,N_6806,N_7463);
xnor U8466 (N_8466,N_6711,N_6653);
or U8467 (N_8467,N_6231,N_6125);
nor U8468 (N_8468,N_6302,N_6600);
xor U8469 (N_8469,N_7060,N_7374);
nor U8470 (N_8470,N_6790,N_6290);
xor U8471 (N_8471,N_6675,N_6925);
nor U8472 (N_8472,N_6156,N_6637);
and U8473 (N_8473,N_7440,N_7306);
and U8474 (N_8474,N_7022,N_6680);
and U8475 (N_8475,N_7000,N_6717);
nand U8476 (N_8476,N_6086,N_6515);
nand U8477 (N_8477,N_6456,N_6053);
or U8478 (N_8478,N_6358,N_7363);
nor U8479 (N_8479,N_6395,N_6935);
nand U8480 (N_8480,N_7176,N_6097);
nor U8481 (N_8481,N_7060,N_7494);
and U8482 (N_8482,N_6190,N_6632);
and U8483 (N_8483,N_6997,N_6247);
or U8484 (N_8484,N_6648,N_6470);
xnor U8485 (N_8485,N_6995,N_6112);
xor U8486 (N_8486,N_6807,N_7007);
nand U8487 (N_8487,N_6315,N_6382);
and U8488 (N_8488,N_6061,N_7245);
or U8489 (N_8489,N_6683,N_7051);
xor U8490 (N_8490,N_6287,N_6151);
xor U8491 (N_8491,N_7149,N_6488);
xor U8492 (N_8492,N_6149,N_6801);
and U8493 (N_8493,N_6388,N_7324);
nand U8494 (N_8494,N_7408,N_6340);
xnor U8495 (N_8495,N_6601,N_6600);
and U8496 (N_8496,N_7310,N_6503);
nor U8497 (N_8497,N_6709,N_6540);
and U8498 (N_8498,N_7091,N_6460);
or U8499 (N_8499,N_6968,N_6145);
nor U8500 (N_8500,N_6869,N_7262);
and U8501 (N_8501,N_6750,N_6760);
nand U8502 (N_8502,N_7254,N_6752);
or U8503 (N_8503,N_7441,N_6030);
xnor U8504 (N_8504,N_6297,N_7039);
xor U8505 (N_8505,N_6850,N_7045);
xnor U8506 (N_8506,N_7463,N_6371);
xor U8507 (N_8507,N_7306,N_6563);
nor U8508 (N_8508,N_7042,N_7375);
nor U8509 (N_8509,N_7033,N_7470);
nor U8510 (N_8510,N_7333,N_6184);
xnor U8511 (N_8511,N_6951,N_6728);
xnor U8512 (N_8512,N_7157,N_6409);
xor U8513 (N_8513,N_6562,N_7354);
and U8514 (N_8514,N_6178,N_6637);
or U8515 (N_8515,N_6689,N_6661);
or U8516 (N_8516,N_7253,N_6628);
xnor U8517 (N_8517,N_6803,N_6869);
nand U8518 (N_8518,N_7023,N_7270);
xor U8519 (N_8519,N_7042,N_6279);
or U8520 (N_8520,N_6498,N_6407);
or U8521 (N_8521,N_6373,N_6833);
nor U8522 (N_8522,N_6232,N_7118);
nand U8523 (N_8523,N_6273,N_6598);
nor U8524 (N_8524,N_6103,N_6183);
nor U8525 (N_8525,N_7466,N_6775);
xnor U8526 (N_8526,N_7174,N_7377);
or U8527 (N_8527,N_6338,N_6029);
or U8528 (N_8528,N_6431,N_7005);
and U8529 (N_8529,N_6890,N_7369);
and U8530 (N_8530,N_6901,N_7156);
and U8531 (N_8531,N_6562,N_7355);
nor U8532 (N_8532,N_7092,N_7488);
and U8533 (N_8533,N_6334,N_7107);
or U8534 (N_8534,N_6695,N_6225);
or U8535 (N_8535,N_6404,N_6857);
nor U8536 (N_8536,N_6152,N_7257);
xnor U8537 (N_8537,N_6973,N_6797);
or U8538 (N_8538,N_7239,N_6075);
nor U8539 (N_8539,N_6652,N_7435);
xor U8540 (N_8540,N_6386,N_6563);
xnor U8541 (N_8541,N_7092,N_7166);
nor U8542 (N_8542,N_7213,N_7455);
or U8543 (N_8543,N_6910,N_7444);
xor U8544 (N_8544,N_6234,N_6427);
xor U8545 (N_8545,N_6103,N_6044);
nor U8546 (N_8546,N_6150,N_6659);
xor U8547 (N_8547,N_6534,N_6267);
nor U8548 (N_8548,N_7196,N_6272);
nor U8549 (N_8549,N_7150,N_6700);
nor U8550 (N_8550,N_7067,N_6840);
nor U8551 (N_8551,N_7477,N_6256);
and U8552 (N_8552,N_7027,N_7477);
nor U8553 (N_8553,N_7332,N_7438);
nand U8554 (N_8554,N_7484,N_7170);
nor U8555 (N_8555,N_7310,N_7217);
nor U8556 (N_8556,N_7006,N_7054);
or U8557 (N_8557,N_6272,N_6974);
nor U8558 (N_8558,N_6545,N_6766);
nand U8559 (N_8559,N_6884,N_7290);
xor U8560 (N_8560,N_6311,N_7462);
and U8561 (N_8561,N_6620,N_6549);
nand U8562 (N_8562,N_6421,N_6038);
nor U8563 (N_8563,N_6975,N_7074);
nand U8564 (N_8564,N_6722,N_6114);
nand U8565 (N_8565,N_6650,N_6388);
and U8566 (N_8566,N_7017,N_6125);
nor U8567 (N_8567,N_7263,N_6457);
nor U8568 (N_8568,N_7018,N_6844);
and U8569 (N_8569,N_7147,N_6196);
nor U8570 (N_8570,N_6054,N_6999);
or U8571 (N_8571,N_7127,N_7095);
xor U8572 (N_8572,N_7069,N_7371);
nor U8573 (N_8573,N_6262,N_7043);
nand U8574 (N_8574,N_7057,N_6003);
and U8575 (N_8575,N_6449,N_6131);
nand U8576 (N_8576,N_6797,N_6993);
xnor U8577 (N_8577,N_6307,N_6455);
nand U8578 (N_8578,N_6665,N_6844);
nand U8579 (N_8579,N_7207,N_6456);
nand U8580 (N_8580,N_7284,N_6066);
xnor U8581 (N_8581,N_6582,N_6002);
xnor U8582 (N_8582,N_6779,N_6468);
and U8583 (N_8583,N_6580,N_6475);
or U8584 (N_8584,N_6378,N_6149);
nor U8585 (N_8585,N_6722,N_7396);
nand U8586 (N_8586,N_6925,N_6002);
nand U8587 (N_8587,N_6786,N_7150);
or U8588 (N_8588,N_6548,N_7122);
and U8589 (N_8589,N_6020,N_6421);
nor U8590 (N_8590,N_7001,N_7165);
nand U8591 (N_8591,N_6620,N_6974);
xor U8592 (N_8592,N_7307,N_6416);
or U8593 (N_8593,N_6548,N_7366);
or U8594 (N_8594,N_6757,N_6714);
nand U8595 (N_8595,N_6806,N_7191);
and U8596 (N_8596,N_6333,N_6973);
nand U8597 (N_8597,N_7189,N_6273);
xnor U8598 (N_8598,N_6466,N_6277);
nor U8599 (N_8599,N_6035,N_6305);
xor U8600 (N_8600,N_6392,N_6966);
xor U8601 (N_8601,N_6954,N_6633);
and U8602 (N_8602,N_6031,N_7095);
nor U8603 (N_8603,N_7454,N_6115);
nand U8604 (N_8604,N_7455,N_6828);
nor U8605 (N_8605,N_7463,N_6044);
nand U8606 (N_8606,N_6492,N_6400);
xor U8607 (N_8607,N_6490,N_7251);
and U8608 (N_8608,N_7237,N_7297);
nand U8609 (N_8609,N_7126,N_7321);
nand U8610 (N_8610,N_6550,N_6119);
and U8611 (N_8611,N_6449,N_6304);
nand U8612 (N_8612,N_7108,N_7378);
xnor U8613 (N_8613,N_6960,N_7498);
nor U8614 (N_8614,N_6661,N_6738);
or U8615 (N_8615,N_6652,N_6691);
nor U8616 (N_8616,N_7036,N_7446);
nor U8617 (N_8617,N_6077,N_7230);
and U8618 (N_8618,N_7062,N_6241);
nand U8619 (N_8619,N_6266,N_6171);
or U8620 (N_8620,N_6105,N_6769);
or U8621 (N_8621,N_6291,N_6397);
and U8622 (N_8622,N_6883,N_6758);
nor U8623 (N_8623,N_7468,N_6997);
and U8624 (N_8624,N_7279,N_7421);
xnor U8625 (N_8625,N_7169,N_6293);
or U8626 (N_8626,N_6264,N_7474);
xnor U8627 (N_8627,N_7085,N_6337);
xor U8628 (N_8628,N_6501,N_6769);
nor U8629 (N_8629,N_6159,N_6545);
or U8630 (N_8630,N_6570,N_7350);
nand U8631 (N_8631,N_6654,N_6157);
nor U8632 (N_8632,N_7088,N_6930);
or U8633 (N_8633,N_6159,N_6028);
nor U8634 (N_8634,N_6871,N_6123);
nand U8635 (N_8635,N_6301,N_6991);
or U8636 (N_8636,N_6774,N_6143);
xor U8637 (N_8637,N_6361,N_6417);
nand U8638 (N_8638,N_7239,N_6795);
nor U8639 (N_8639,N_6586,N_7485);
and U8640 (N_8640,N_6969,N_6171);
or U8641 (N_8641,N_6068,N_7156);
and U8642 (N_8642,N_6863,N_7080);
xnor U8643 (N_8643,N_6921,N_7231);
or U8644 (N_8644,N_6943,N_7053);
nand U8645 (N_8645,N_7392,N_7368);
or U8646 (N_8646,N_7463,N_6225);
xnor U8647 (N_8647,N_6963,N_7451);
nor U8648 (N_8648,N_6833,N_6402);
nor U8649 (N_8649,N_6411,N_7268);
nand U8650 (N_8650,N_6394,N_7234);
or U8651 (N_8651,N_6426,N_6608);
xor U8652 (N_8652,N_6810,N_6497);
and U8653 (N_8653,N_7019,N_6476);
nand U8654 (N_8654,N_6343,N_7268);
nand U8655 (N_8655,N_6719,N_6428);
xnor U8656 (N_8656,N_7097,N_6771);
xor U8657 (N_8657,N_6362,N_6882);
and U8658 (N_8658,N_6730,N_6259);
nor U8659 (N_8659,N_7155,N_6604);
xor U8660 (N_8660,N_7331,N_6977);
nor U8661 (N_8661,N_6095,N_6180);
nor U8662 (N_8662,N_7328,N_6053);
or U8663 (N_8663,N_6694,N_6750);
nand U8664 (N_8664,N_6358,N_6393);
xor U8665 (N_8665,N_6730,N_6681);
and U8666 (N_8666,N_6668,N_6229);
nor U8667 (N_8667,N_6094,N_7320);
and U8668 (N_8668,N_6661,N_6036);
nor U8669 (N_8669,N_6713,N_7433);
xor U8670 (N_8670,N_7334,N_6943);
or U8671 (N_8671,N_6223,N_6434);
nor U8672 (N_8672,N_7341,N_6961);
nand U8673 (N_8673,N_6408,N_6365);
and U8674 (N_8674,N_6779,N_6741);
xnor U8675 (N_8675,N_6183,N_6740);
or U8676 (N_8676,N_7285,N_6890);
and U8677 (N_8677,N_6649,N_6538);
nor U8678 (N_8678,N_7311,N_7036);
and U8679 (N_8679,N_6116,N_6908);
or U8680 (N_8680,N_6391,N_6713);
nor U8681 (N_8681,N_6949,N_6404);
nor U8682 (N_8682,N_6554,N_6856);
nand U8683 (N_8683,N_6548,N_6286);
or U8684 (N_8684,N_6144,N_6677);
nand U8685 (N_8685,N_6919,N_6925);
nor U8686 (N_8686,N_6383,N_7224);
and U8687 (N_8687,N_6882,N_6112);
or U8688 (N_8688,N_6708,N_6075);
or U8689 (N_8689,N_6510,N_7427);
nand U8690 (N_8690,N_6528,N_7441);
or U8691 (N_8691,N_6556,N_6000);
xor U8692 (N_8692,N_6711,N_6029);
xnor U8693 (N_8693,N_7121,N_7096);
nand U8694 (N_8694,N_6631,N_6766);
xor U8695 (N_8695,N_6782,N_6779);
and U8696 (N_8696,N_6370,N_7036);
nor U8697 (N_8697,N_6210,N_7418);
nand U8698 (N_8698,N_6099,N_7059);
or U8699 (N_8699,N_6426,N_6349);
or U8700 (N_8700,N_7493,N_7261);
or U8701 (N_8701,N_6069,N_7338);
and U8702 (N_8702,N_6732,N_7411);
or U8703 (N_8703,N_7223,N_6577);
or U8704 (N_8704,N_6454,N_6287);
and U8705 (N_8705,N_6879,N_7451);
xor U8706 (N_8706,N_6280,N_6606);
nor U8707 (N_8707,N_7073,N_6718);
nor U8708 (N_8708,N_6528,N_6532);
and U8709 (N_8709,N_7216,N_6233);
nor U8710 (N_8710,N_7148,N_6652);
nand U8711 (N_8711,N_6689,N_6718);
xor U8712 (N_8712,N_6531,N_6106);
or U8713 (N_8713,N_6815,N_6455);
nor U8714 (N_8714,N_7062,N_7125);
xor U8715 (N_8715,N_6051,N_6107);
nor U8716 (N_8716,N_6167,N_7310);
and U8717 (N_8717,N_7203,N_6479);
or U8718 (N_8718,N_7434,N_6274);
nor U8719 (N_8719,N_6403,N_7473);
and U8720 (N_8720,N_7331,N_7107);
nand U8721 (N_8721,N_6619,N_7168);
nor U8722 (N_8722,N_6644,N_6329);
nor U8723 (N_8723,N_6877,N_6283);
or U8724 (N_8724,N_7397,N_7264);
and U8725 (N_8725,N_6244,N_6910);
nand U8726 (N_8726,N_6163,N_6726);
xnor U8727 (N_8727,N_6428,N_7397);
and U8728 (N_8728,N_7101,N_7450);
and U8729 (N_8729,N_7326,N_6828);
and U8730 (N_8730,N_7051,N_6154);
nor U8731 (N_8731,N_7455,N_6141);
nand U8732 (N_8732,N_6337,N_6001);
xnor U8733 (N_8733,N_6045,N_7300);
and U8734 (N_8734,N_6630,N_6831);
or U8735 (N_8735,N_7472,N_7102);
nor U8736 (N_8736,N_6561,N_6886);
nor U8737 (N_8737,N_6813,N_6390);
nor U8738 (N_8738,N_6453,N_6325);
nand U8739 (N_8739,N_7156,N_7322);
nor U8740 (N_8740,N_6572,N_6941);
xnor U8741 (N_8741,N_6055,N_6374);
nor U8742 (N_8742,N_6519,N_6270);
nand U8743 (N_8743,N_6298,N_6594);
nor U8744 (N_8744,N_6524,N_6014);
and U8745 (N_8745,N_7402,N_7425);
or U8746 (N_8746,N_6872,N_6080);
or U8747 (N_8747,N_6498,N_7486);
nor U8748 (N_8748,N_6575,N_7494);
or U8749 (N_8749,N_6229,N_7142);
xor U8750 (N_8750,N_6278,N_6946);
xor U8751 (N_8751,N_6951,N_6420);
and U8752 (N_8752,N_6973,N_7352);
xnor U8753 (N_8753,N_7297,N_7381);
and U8754 (N_8754,N_6854,N_7389);
and U8755 (N_8755,N_6499,N_6097);
nand U8756 (N_8756,N_6519,N_7459);
nand U8757 (N_8757,N_7346,N_7322);
nand U8758 (N_8758,N_7469,N_6369);
xnor U8759 (N_8759,N_7183,N_6756);
or U8760 (N_8760,N_6689,N_6743);
xor U8761 (N_8761,N_6313,N_7024);
nor U8762 (N_8762,N_6969,N_6691);
nor U8763 (N_8763,N_6009,N_6135);
nor U8764 (N_8764,N_6509,N_6278);
nor U8765 (N_8765,N_6075,N_6728);
or U8766 (N_8766,N_6288,N_7479);
and U8767 (N_8767,N_6585,N_6438);
xor U8768 (N_8768,N_7041,N_6900);
nand U8769 (N_8769,N_6020,N_7177);
or U8770 (N_8770,N_7438,N_7324);
or U8771 (N_8771,N_6451,N_6083);
xnor U8772 (N_8772,N_6276,N_6110);
xnor U8773 (N_8773,N_7332,N_7041);
nand U8774 (N_8774,N_6173,N_7214);
xnor U8775 (N_8775,N_6004,N_7477);
nand U8776 (N_8776,N_6813,N_7356);
xor U8777 (N_8777,N_6839,N_6585);
and U8778 (N_8778,N_6384,N_6772);
or U8779 (N_8779,N_7102,N_7438);
or U8780 (N_8780,N_6666,N_6651);
or U8781 (N_8781,N_6180,N_7446);
nor U8782 (N_8782,N_6501,N_6141);
nand U8783 (N_8783,N_6913,N_7076);
nand U8784 (N_8784,N_6456,N_7107);
and U8785 (N_8785,N_6228,N_7010);
nor U8786 (N_8786,N_6016,N_6726);
and U8787 (N_8787,N_6341,N_7062);
nand U8788 (N_8788,N_6422,N_6072);
nand U8789 (N_8789,N_7072,N_6452);
xnor U8790 (N_8790,N_7482,N_6648);
nor U8791 (N_8791,N_7080,N_7017);
nor U8792 (N_8792,N_6173,N_7280);
and U8793 (N_8793,N_6604,N_7284);
xnor U8794 (N_8794,N_6626,N_7262);
or U8795 (N_8795,N_6794,N_7421);
nand U8796 (N_8796,N_7343,N_7405);
nand U8797 (N_8797,N_6881,N_7122);
nor U8798 (N_8798,N_6011,N_7407);
nand U8799 (N_8799,N_6631,N_6908);
or U8800 (N_8800,N_6955,N_6171);
and U8801 (N_8801,N_6818,N_6990);
or U8802 (N_8802,N_6578,N_7235);
or U8803 (N_8803,N_7356,N_7335);
nor U8804 (N_8804,N_6108,N_7307);
xnor U8805 (N_8805,N_6491,N_6430);
xor U8806 (N_8806,N_6822,N_6590);
nand U8807 (N_8807,N_7273,N_6417);
nand U8808 (N_8808,N_6314,N_7356);
or U8809 (N_8809,N_6897,N_6225);
and U8810 (N_8810,N_6523,N_7358);
or U8811 (N_8811,N_6765,N_6970);
nor U8812 (N_8812,N_7005,N_6876);
xnor U8813 (N_8813,N_7237,N_6452);
nor U8814 (N_8814,N_7144,N_7435);
or U8815 (N_8815,N_6021,N_6174);
nor U8816 (N_8816,N_6764,N_6356);
nor U8817 (N_8817,N_6391,N_7283);
or U8818 (N_8818,N_6580,N_6584);
and U8819 (N_8819,N_6611,N_7235);
nor U8820 (N_8820,N_6748,N_6774);
nand U8821 (N_8821,N_6487,N_7362);
or U8822 (N_8822,N_6900,N_6662);
or U8823 (N_8823,N_6165,N_6456);
or U8824 (N_8824,N_6483,N_7234);
or U8825 (N_8825,N_7207,N_6818);
nor U8826 (N_8826,N_6763,N_6829);
or U8827 (N_8827,N_6612,N_6607);
or U8828 (N_8828,N_6985,N_6136);
nor U8829 (N_8829,N_7130,N_6493);
xor U8830 (N_8830,N_6334,N_6297);
nor U8831 (N_8831,N_6484,N_6402);
nand U8832 (N_8832,N_6035,N_6745);
nand U8833 (N_8833,N_6993,N_6392);
or U8834 (N_8834,N_6106,N_7246);
nand U8835 (N_8835,N_6134,N_7206);
nor U8836 (N_8836,N_7170,N_7224);
and U8837 (N_8837,N_6718,N_6284);
or U8838 (N_8838,N_6715,N_6039);
nand U8839 (N_8839,N_6991,N_6567);
or U8840 (N_8840,N_7425,N_7084);
xor U8841 (N_8841,N_6640,N_7111);
or U8842 (N_8842,N_6293,N_7150);
nand U8843 (N_8843,N_6138,N_7452);
xnor U8844 (N_8844,N_6582,N_6996);
nand U8845 (N_8845,N_6192,N_6873);
xor U8846 (N_8846,N_6006,N_6351);
nand U8847 (N_8847,N_6303,N_6513);
xnor U8848 (N_8848,N_6165,N_7433);
or U8849 (N_8849,N_6328,N_6252);
nor U8850 (N_8850,N_7237,N_7081);
nor U8851 (N_8851,N_6487,N_6247);
or U8852 (N_8852,N_6804,N_6006);
nand U8853 (N_8853,N_6639,N_6170);
nand U8854 (N_8854,N_6774,N_6907);
xnor U8855 (N_8855,N_6459,N_7300);
xnor U8856 (N_8856,N_6923,N_7358);
xnor U8857 (N_8857,N_6640,N_6318);
nor U8858 (N_8858,N_6370,N_7170);
nor U8859 (N_8859,N_6927,N_6648);
or U8860 (N_8860,N_6072,N_7013);
xnor U8861 (N_8861,N_7186,N_6625);
nand U8862 (N_8862,N_6627,N_7279);
or U8863 (N_8863,N_7320,N_7048);
xnor U8864 (N_8864,N_7308,N_7011);
nand U8865 (N_8865,N_6673,N_7217);
or U8866 (N_8866,N_6514,N_6428);
nor U8867 (N_8867,N_6540,N_6863);
nand U8868 (N_8868,N_6400,N_7382);
and U8869 (N_8869,N_6508,N_6588);
nor U8870 (N_8870,N_6015,N_6371);
or U8871 (N_8871,N_6836,N_7261);
nor U8872 (N_8872,N_6843,N_6210);
xnor U8873 (N_8873,N_6560,N_6735);
nand U8874 (N_8874,N_6341,N_6919);
and U8875 (N_8875,N_7016,N_7496);
and U8876 (N_8876,N_7275,N_6668);
nor U8877 (N_8877,N_7134,N_6109);
or U8878 (N_8878,N_7466,N_7358);
nor U8879 (N_8879,N_6278,N_6241);
xor U8880 (N_8880,N_6577,N_6189);
and U8881 (N_8881,N_6176,N_6214);
nor U8882 (N_8882,N_6225,N_7423);
or U8883 (N_8883,N_6081,N_6075);
and U8884 (N_8884,N_7458,N_6636);
and U8885 (N_8885,N_7287,N_6778);
and U8886 (N_8886,N_6321,N_6525);
xor U8887 (N_8887,N_6394,N_7339);
nand U8888 (N_8888,N_6852,N_6502);
or U8889 (N_8889,N_6625,N_6681);
nand U8890 (N_8890,N_7238,N_6215);
or U8891 (N_8891,N_6526,N_6143);
nand U8892 (N_8892,N_6415,N_6179);
and U8893 (N_8893,N_7166,N_7317);
nor U8894 (N_8894,N_7387,N_6484);
or U8895 (N_8895,N_7078,N_6383);
nand U8896 (N_8896,N_6333,N_6532);
nand U8897 (N_8897,N_6063,N_6488);
and U8898 (N_8898,N_6209,N_6217);
nor U8899 (N_8899,N_6184,N_7447);
nor U8900 (N_8900,N_6998,N_6168);
or U8901 (N_8901,N_7101,N_6098);
xnor U8902 (N_8902,N_6248,N_7298);
nand U8903 (N_8903,N_7371,N_6834);
or U8904 (N_8904,N_6471,N_6140);
or U8905 (N_8905,N_6142,N_6763);
xor U8906 (N_8906,N_6385,N_7470);
nor U8907 (N_8907,N_6748,N_6185);
nor U8908 (N_8908,N_7428,N_6048);
or U8909 (N_8909,N_6567,N_6142);
or U8910 (N_8910,N_6053,N_6206);
and U8911 (N_8911,N_6150,N_6393);
xnor U8912 (N_8912,N_7407,N_6124);
and U8913 (N_8913,N_6782,N_7488);
xnor U8914 (N_8914,N_6488,N_7001);
or U8915 (N_8915,N_6636,N_6664);
and U8916 (N_8916,N_6604,N_7013);
nand U8917 (N_8917,N_6262,N_6322);
and U8918 (N_8918,N_7218,N_6562);
and U8919 (N_8919,N_6885,N_6240);
xnor U8920 (N_8920,N_7193,N_6503);
or U8921 (N_8921,N_7117,N_7010);
nand U8922 (N_8922,N_7174,N_6618);
nor U8923 (N_8923,N_6543,N_7020);
nor U8924 (N_8924,N_6437,N_6848);
or U8925 (N_8925,N_7255,N_6559);
nor U8926 (N_8926,N_7407,N_7276);
or U8927 (N_8927,N_6759,N_6414);
nand U8928 (N_8928,N_7051,N_6374);
xnor U8929 (N_8929,N_6459,N_6348);
and U8930 (N_8930,N_7146,N_7150);
xnor U8931 (N_8931,N_6506,N_6394);
nor U8932 (N_8932,N_6637,N_6840);
xor U8933 (N_8933,N_6216,N_7462);
nand U8934 (N_8934,N_6254,N_7044);
nand U8935 (N_8935,N_6292,N_7256);
nand U8936 (N_8936,N_7086,N_7217);
and U8937 (N_8937,N_7394,N_6546);
or U8938 (N_8938,N_6504,N_6805);
and U8939 (N_8939,N_6156,N_7427);
or U8940 (N_8940,N_6131,N_6923);
and U8941 (N_8941,N_6383,N_6387);
xor U8942 (N_8942,N_6781,N_6514);
xnor U8943 (N_8943,N_6419,N_7486);
and U8944 (N_8944,N_6252,N_6020);
and U8945 (N_8945,N_7099,N_6463);
nor U8946 (N_8946,N_7113,N_6849);
xor U8947 (N_8947,N_7083,N_6587);
nor U8948 (N_8948,N_6999,N_6561);
nor U8949 (N_8949,N_7288,N_7338);
xnor U8950 (N_8950,N_6908,N_6879);
or U8951 (N_8951,N_7184,N_7240);
nand U8952 (N_8952,N_6784,N_6210);
nand U8953 (N_8953,N_7059,N_6371);
or U8954 (N_8954,N_7021,N_6149);
or U8955 (N_8955,N_6302,N_6517);
xnor U8956 (N_8956,N_6871,N_6951);
and U8957 (N_8957,N_6820,N_6023);
nand U8958 (N_8958,N_6545,N_6419);
and U8959 (N_8959,N_6771,N_6009);
nand U8960 (N_8960,N_6124,N_6921);
nor U8961 (N_8961,N_7175,N_6818);
or U8962 (N_8962,N_6901,N_6631);
and U8963 (N_8963,N_6804,N_6246);
or U8964 (N_8964,N_6559,N_6103);
nor U8965 (N_8965,N_6310,N_6212);
xor U8966 (N_8966,N_7120,N_6464);
and U8967 (N_8967,N_6968,N_7103);
and U8968 (N_8968,N_6480,N_6231);
or U8969 (N_8969,N_6933,N_7292);
or U8970 (N_8970,N_7323,N_7333);
xnor U8971 (N_8971,N_6870,N_7349);
nand U8972 (N_8972,N_6679,N_7324);
nand U8973 (N_8973,N_6585,N_6620);
nor U8974 (N_8974,N_7054,N_6499);
and U8975 (N_8975,N_6903,N_7476);
nand U8976 (N_8976,N_6734,N_6304);
nand U8977 (N_8977,N_7021,N_7174);
and U8978 (N_8978,N_7127,N_7008);
xnor U8979 (N_8979,N_6113,N_6697);
nor U8980 (N_8980,N_6676,N_7287);
nor U8981 (N_8981,N_6924,N_6493);
xnor U8982 (N_8982,N_6293,N_7245);
xnor U8983 (N_8983,N_7195,N_6910);
nand U8984 (N_8984,N_6552,N_6339);
or U8985 (N_8985,N_7066,N_6343);
and U8986 (N_8986,N_7157,N_6751);
or U8987 (N_8987,N_6929,N_7113);
or U8988 (N_8988,N_7427,N_7038);
nand U8989 (N_8989,N_6432,N_6172);
or U8990 (N_8990,N_6288,N_6955);
or U8991 (N_8991,N_6995,N_6272);
or U8992 (N_8992,N_7008,N_6448);
nand U8993 (N_8993,N_7308,N_6148);
or U8994 (N_8994,N_6280,N_6363);
xor U8995 (N_8995,N_6677,N_7436);
or U8996 (N_8996,N_6398,N_6892);
nand U8997 (N_8997,N_6073,N_6239);
nor U8998 (N_8998,N_6377,N_6370);
or U8999 (N_8999,N_6350,N_6437);
xor U9000 (N_9000,N_8181,N_8753);
nand U9001 (N_9001,N_8131,N_8288);
nor U9002 (N_9002,N_8120,N_8231);
and U9003 (N_9003,N_7780,N_7836);
or U9004 (N_9004,N_8700,N_8324);
nand U9005 (N_9005,N_7825,N_8440);
nor U9006 (N_9006,N_8575,N_8207);
nor U9007 (N_9007,N_7858,N_8280);
nand U9008 (N_9008,N_7509,N_8642);
and U9009 (N_9009,N_8005,N_7711);
and U9010 (N_9010,N_8279,N_7679);
nand U9011 (N_9011,N_8540,N_7748);
xnor U9012 (N_9012,N_7642,N_7755);
xnor U9013 (N_9013,N_8070,N_7526);
nor U9014 (N_9014,N_8235,N_8460);
or U9015 (N_9015,N_7828,N_8903);
nor U9016 (N_9016,N_7518,N_8143);
nand U9017 (N_9017,N_8317,N_7523);
and U9018 (N_9018,N_7619,N_8793);
and U9019 (N_9019,N_8448,N_8441);
nand U9020 (N_9020,N_7702,N_8434);
or U9021 (N_9021,N_8619,N_8667);
and U9022 (N_9022,N_8788,N_8176);
or U9023 (N_9023,N_8305,N_8817);
or U9024 (N_9024,N_7889,N_8396);
or U9025 (N_9025,N_7637,N_7718);
or U9026 (N_9026,N_8194,N_7528);
or U9027 (N_9027,N_8772,N_8372);
xor U9028 (N_9028,N_8155,N_7513);
or U9029 (N_9029,N_7798,N_8987);
or U9030 (N_9030,N_8385,N_7613);
or U9031 (N_9031,N_8364,N_8278);
or U9032 (N_9032,N_8552,N_7882);
nand U9033 (N_9033,N_8493,N_8273);
xnor U9034 (N_9034,N_8365,N_8632);
or U9035 (N_9035,N_8560,N_8999);
or U9036 (N_9036,N_7631,N_8393);
xnor U9037 (N_9037,N_7773,N_8205);
nor U9038 (N_9038,N_7878,N_7556);
or U9039 (N_9039,N_8296,N_7598);
nand U9040 (N_9040,N_7620,N_7768);
xor U9041 (N_9041,N_8362,N_8764);
nor U9042 (N_9042,N_8369,N_8402);
xnor U9043 (N_9043,N_7895,N_8891);
nor U9044 (N_9044,N_7508,N_8554);
and U9045 (N_9045,N_7861,N_7535);
or U9046 (N_9046,N_8811,N_8929);
and U9047 (N_9047,N_8838,N_7662);
and U9048 (N_9048,N_7687,N_8931);
nand U9049 (N_9049,N_7700,N_8154);
nand U9050 (N_9050,N_7550,N_8146);
xnor U9051 (N_9051,N_8060,N_8666);
nand U9052 (N_9052,N_8675,N_8980);
nor U9053 (N_9053,N_7677,N_8341);
and U9054 (N_9054,N_8246,N_8487);
nor U9055 (N_9055,N_8130,N_8658);
nor U9056 (N_9056,N_7573,N_7717);
nor U9057 (N_9057,N_8072,N_8860);
nor U9058 (N_9058,N_8428,N_8303);
and U9059 (N_9059,N_8602,N_8300);
nor U9060 (N_9060,N_8914,N_7776);
nand U9061 (N_9061,N_8265,N_8681);
and U9062 (N_9062,N_7941,N_7582);
nor U9063 (N_9063,N_8179,N_7788);
and U9064 (N_9064,N_7971,N_7913);
and U9065 (N_9065,N_8243,N_7760);
nor U9066 (N_9066,N_7908,N_8028);
nor U9067 (N_9067,N_7705,N_8913);
xor U9068 (N_9068,N_8988,N_7854);
nand U9069 (N_9069,N_7939,N_8629);
xor U9070 (N_9070,N_8590,N_8375);
xnor U9071 (N_9071,N_8550,N_8180);
xor U9072 (N_9072,N_8345,N_7988);
nor U9073 (N_9073,N_7554,N_7749);
and U9074 (N_9074,N_8065,N_8209);
xnor U9075 (N_9075,N_7820,N_8970);
nor U9076 (N_9076,N_8486,N_8519);
nand U9077 (N_9077,N_8697,N_7622);
nor U9078 (N_9078,N_8757,N_7577);
nand U9079 (N_9079,N_7511,N_7886);
and U9080 (N_9080,N_7616,N_8570);
xor U9081 (N_9081,N_8046,N_8864);
xor U9082 (N_9082,N_8614,N_8686);
nor U9083 (N_9083,N_8342,N_7815);
nor U9084 (N_9084,N_7970,N_7512);
and U9085 (N_9085,N_8054,N_8746);
xor U9086 (N_9086,N_8249,N_7781);
and U9087 (N_9087,N_7686,N_8151);
nor U9088 (N_9088,N_7729,N_8177);
and U9089 (N_9089,N_7843,N_8832);
xor U9090 (N_9090,N_8924,N_8321);
or U9091 (N_9091,N_7990,N_8383);
and U9092 (N_9092,N_7545,N_8869);
and U9093 (N_9093,N_8261,N_8933);
nand U9094 (N_9094,N_8170,N_8233);
nand U9095 (N_9095,N_7605,N_7860);
nand U9096 (N_9096,N_8615,N_7503);
nor U9097 (N_9097,N_8014,N_8297);
and U9098 (N_9098,N_8709,N_8268);
nor U9099 (N_9099,N_7847,N_8865);
nor U9100 (N_9100,N_8171,N_8814);
and U9101 (N_9101,N_8941,N_8057);
xnor U9102 (N_9102,N_7593,N_8319);
and U9103 (N_9103,N_8359,N_8902);
xor U9104 (N_9104,N_8080,N_8756);
nand U9105 (N_9105,N_8272,N_8915);
or U9106 (N_9106,N_8670,N_7903);
nand U9107 (N_9107,N_8524,N_8527);
nand U9108 (N_9108,N_8720,N_8328);
or U9109 (N_9109,N_8985,N_8162);
or U9110 (N_9110,N_8457,N_7816);
nand U9111 (N_9111,N_7848,N_8517);
nand U9112 (N_9112,N_7692,N_8103);
nor U9113 (N_9113,N_8821,N_7698);
nor U9114 (N_9114,N_8430,N_7563);
nand U9115 (N_9115,N_8047,N_8627);
nand U9116 (N_9116,N_8888,N_7767);
and U9117 (N_9117,N_8022,N_7710);
or U9118 (N_9118,N_7694,N_8710);
nor U9119 (N_9119,N_8077,N_7562);
nor U9120 (N_9120,N_7958,N_8559);
nand U9121 (N_9121,N_8734,N_7993);
and U9122 (N_9122,N_8545,N_8168);
nand U9123 (N_9123,N_7728,N_7719);
nor U9124 (N_9124,N_8325,N_8528);
nor U9125 (N_9125,N_7510,N_8594);
xnor U9126 (N_9126,N_8290,N_7972);
and U9127 (N_9127,N_7830,N_8724);
or U9128 (N_9128,N_7532,N_7937);
and U9129 (N_9129,N_8637,N_7638);
or U9130 (N_9130,N_8073,N_8326);
and U9131 (N_9131,N_7887,N_8107);
or U9132 (N_9132,N_7880,N_8355);
nand U9133 (N_9133,N_8128,N_7560);
xor U9134 (N_9134,N_7738,N_8641);
xor U9135 (N_9135,N_8652,N_7856);
nand U9136 (N_9136,N_8908,N_8435);
and U9137 (N_9137,N_8684,N_8165);
or U9138 (N_9138,N_8271,N_8818);
and U9139 (N_9139,N_8089,N_8356);
nand U9140 (N_9140,N_8971,N_7792);
xor U9141 (N_9141,N_8648,N_8188);
nor U9142 (N_9142,N_7986,N_8683);
or U9143 (N_9143,N_8225,N_8782);
xor U9144 (N_9144,N_8537,N_8230);
or U9145 (N_9145,N_7930,N_7585);
nor U9146 (N_9146,N_8136,N_7678);
xor U9147 (N_9147,N_8877,N_8939);
and U9148 (N_9148,N_8132,N_8127);
and U9149 (N_9149,N_8783,N_7961);
and U9150 (N_9150,N_7984,N_7983);
xor U9151 (N_9151,N_8829,N_7746);
nor U9152 (N_9152,N_8714,N_8467);
xor U9153 (N_9153,N_8662,N_8639);
or U9154 (N_9154,N_7869,N_7575);
xnor U9155 (N_9155,N_7940,N_7609);
and U9156 (N_9156,N_7991,N_7826);
nor U9157 (N_9157,N_8079,N_8631);
xor U9158 (N_9158,N_8742,N_8997);
xnor U9159 (N_9159,N_8484,N_7733);
and U9160 (N_9160,N_7802,N_8518);
xor U9161 (N_9161,N_7723,N_8921);
and U9162 (N_9162,N_7516,N_8227);
nand U9163 (N_9163,N_8085,N_8718);
or U9164 (N_9164,N_8992,N_7901);
xnor U9165 (N_9165,N_7845,N_8331);
or U9166 (N_9166,N_7968,N_8160);
xnor U9167 (N_9167,N_8187,N_7963);
nor U9168 (N_9168,N_7542,N_8566);
and U9169 (N_9169,N_8938,N_8766);
and U9170 (N_9170,N_8990,N_8314);
nand U9171 (N_9171,N_7646,N_8117);
nor U9172 (N_9172,N_8466,N_8361);
xnor U9173 (N_9173,N_8056,N_8890);
nor U9174 (N_9174,N_8497,N_7994);
or U9175 (N_9175,N_8926,N_8897);
and U9176 (N_9176,N_8695,N_7641);
and U9177 (N_9177,N_7601,N_8512);
xor U9178 (N_9178,N_8565,N_8794);
nor U9179 (N_9179,N_8775,N_8911);
nor U9180 (N_9180,N_8099,N_7555);
xor U9181 (N_9181,N_7607,N_7501);
nand U9182 (N_9182,N_7800,N_7962);
or U9183 (N_9183,N_8958,N_8717);
xor U9184 (N_9184,N_7676,N_7821);
xnor U9185 (N_9185,N_8896,N_7839);
nand U9186 (N_9186,N_7929,N_8228);
xor U9187 (N_9187,N_8478,N_8124);
and U9188 (N_9188,N_7691,N_8316);
nor U9189 (N_9189,N_8687,N_8221);
or U9190 (N_9190,N_8671,N_8825);
or U9191 (N_9191,N_7649,N_7666);
or U9192 (N_9192,N_7947,N_8673);
nor U9193 (N_9193,N_8354,N_7787);
or U9194 (N_9194,N_8427,N_8691);
xor U9195 (N_9195,N_8880,N_8195);
nor U9196 (N_9196,N_7959,N_8861);
nand U9197 (N_9197,N_8000,N_8021);
nor U9198 (N_9198,N_8978,N_7852);
and U9199 (N_9199,N_8447,N_8520);
nand U9200 (N_9200,N_7714,N_7894);
nand U9201 (N_9201,N_8015,N_7942);
or U9202 (N_9202,N_8101,N_8763);
and U9203 (N_9203,N_8002,N_8031);
nor U9204 (N_9204,N_7791,N_8298);
xnor U9205 (N_9205,N_8960,N_8411);
or U9206 (N_9206,N_7978,N_8850);
nand U9207 (N_9207,N_7757,N_8586);
and U9208 (N_9208,N_8703,N_8844);
or U9209 (N_9209,N_7734,N_7965);
nor U9210 (N_9210,N_7823,N_8954);
nand U9211 (N_9211,N_7764,N_8770);
or U9212 (N_9212,N_8736,N_7627);
and U9213 (N_9213,N_8549,N_8433);
nor U9214 (N_9214,N_7864,N_7916);
xor U9215 (N_9215,N_8508,N_7932);
xor U9216 (N_9216,N_7914,N_7874);
and U9217 (N_9217,N_8175,N_8767);
nor U9218 (N_9218,N_8715,N_8287);
or U9219 (N_9219,N_8664,N_7739);
nor U9220 (N_9220,N_8848,N_8418);
xor U9221 (N_9221,N_7538,N_8100);
and U9222 (N_9222,N_8483,N_8267);
and U9223 (N_9223,N_8708,N_8682);
xnor U9224 (N_9224,N_8489,N_8725);
nor U9225 (N_9225,N_8826,N_8191);
xor U9226 (N_9226,N_8769,N_7564);
nor U9227 (N_9227,N_8285,N_7580);
nand U9228 (N_9228,N_7837,N_7979);
and U9229 (N_9229,N_7907,N_8500);
and U9230 (N_9230,N_8051,N_7911);
or U9231 (N_9231,N_8340,N_7997);
nand U9232 (N_9232,N_8410,N_8463);
and U9233 (N_9233,N_8835,N_8672);
or U9234 (N_9234,N_7547,N_8745);
and U9235 (N_9235,N_8438,N_8762);
or U9236 (N_9236,N_7969,N_8599);
nand U9237 (N_9237,N_8542,N_7838);
and U9238 (N_9238,N_8984,N_8948);
or U9239 (N_9239,N_8465,N_7587);
nor U9240 (N_9240,N_8625,N_8730);
xnor U9241 (N_9241,N_8955,N_7778);
or U9242 (N_9242,N_8828,N_7761);
and U9243 (N_9243,N_7571,N_8184);
nor U9244 (N_9244,N_8951,N_7992);
or U9245 (N_9245,N_7814,N_8561);
and U9246 (N_9246,N_8909,N_8012);
nand U9247 (N_9247,N_8059,N_8417);
nand U9248 (N_9248,N_8308,N_7630);
and U9249 (N_9249,N_7981,N_7931);
or U9250 (N_9250,N_8394,N_7899);
xor U9251 (N_9251,N_7588,N_8514);
or U9252 (N_9252,N_8957,N_8449);
nor U9253 (N_9253,N_8583,N_7656);
and U9254 (N_9254,N_7906,N_8322);
and U9255 (N_9255,N_8640,N_7996);
nand U9256 (N_9256,N_8252,N_8711);
or U9257 (N_9257,N_7989,N_8842);
and U9258 (N_9258,N_7669,N_8286);
xor U9259 (N_9259,N_8592,N_8937);
and U9260 (N_9260,N_7811,N_8238);
xor U9261 (N_9261,N_8546,N_8399);
nand U9262 (N_9262,N_8371,N_8781);
or U9263 (N_9263,N_8747,N_8858);
nand U9264 (N_9264,N_8809,N_8760);
xor U9265 (N_9265,N_8972,N_8480);
nand U9266 (N_9266,N_8502,N_8699);
xnor U9267 (N_9267,N_8579,N_7824);
xnor U9268 (N_9268,N_8704,N_7834);
nor U9269 (N_9269,N_8178,N_8650);
and U9270 (N_9270,N_7667,N_7623);
or U9271 (N_9271,N_8582,N_8907);
and U9272 (N_9272,N_7801,N_8795);
xor U9273 (N_9273,N_8962,N_8967);
or U9274 (N_9274,N_8382,N_8813);
and U9275 (N_9275,N_8019,N_7909);
nor U9276 (N_9276,N_8796,N_7592);
nor U9277 (N_9277,N_8605,N_8996);
and U9278 (N_9278,N_7877,N_8388);
or U9279 (N_9279,N_7844,N_7544);
nand U9280 (N_9280,N_7857,N_8916);
nor U9281 (N_9281,N_8645,N_8623);
or U9282 (N_9282,N_8152,N_8302);
nand U9283 (N_9283,N_8386,N_7715);
or U9284 (N_9284,N_7595,N_8917);
xor U9285 (N_9285,N_8525,N_7831);
xnor U9286 (N_9286,N_7655,N_8603);
nand U9287 (N_9287,N_7604,N_7933);
xnor U9288 (N_9288,N_7810,N_8621);
nor U9289 (N_9289,N_7974,N_8776);
nor U9290 (N_9290,N_8584,N_8475);
nand U9291 (N_9291,N_8349,N_7600);
or U9292 (N_9292,N_8462,N_8733);
nor U9293 (N_9293,N_8250,N_7704);
nand U9294 (N_9294,N_8965,N_8581);
xnor U9295 (N_9295,N_8415,N_8898);
or U9296 (N_9296,N_8805,N_8856);
xnor U9297 (N_9297,N_8368,N_8148);
and U9298 (N_9298,N_8360,N_7817);
and U9299 (N_9299,N_8443,N_8633);
and U9300 (N_9300,N_7569,N_8126);
nor U9301 (N_9301,N_8790,N_8644);
and U9302 (N_9302,N_8048,N_8562);
xnor U9303 (N_9303,N_8713,N_8490);
and U9304 (N_9304,N_8889,N_8893);
nand U9305 (N_9305,N_8919,N_7648);
and U9306 (N_9306,N_7910,N_8289);
nand U9307 (N_9307,N_8949,N_8339);
xor U9308 (N_9308,N_8665,N_7967);
nand U9309 (N_9309,N_7507,N_7625);
xnor U9310 (N_9310,N_8458,N_8208);
nand U9311 (N_9311,N_7846,N_8223);
xnor U9312 (N_9312,N_8153,N_8446);
and U9313 (N_9313,N_7559,N_8934);
nand U9314 (N_9314,N_8093,N_8616);
or U9315 (N_9315,N_8726,N_8058);
nand U9316 (N_9316,N_8845,N_8189);
nor U9317 (N_9317,N_8211,N_8589);
xor U9318 (N_9318,N_8121,N_8011);
or U9319 (N_9319,N_7918,N_7615);
nor U9320 (N_9320,N_7731,N_8569);
or U9321 (N_9321,N_8765,N_7762);
nor U9322 (N_9322,N_8214,N_8881);
or U9323 (N_9323,N_8886,N_7797);
or U9324 (N_9324,N_8017,N_8135);
xor U9325 (N_9325,N_8506,N_8329);
and U9326 (N_9326,N_7543,N_8353);
nor U9327 (N_9327,N_8815,N_8173);
nand U9328 (N_9328,N_7926,N_8118);
and U9329 (N_9329,N_8426,N_8792);
or U9330 (N_9330,N_7807,N_8139);
or U9331 (N_9331,N_8572,N_8312);
and U9332 (N_9332,N_8204,N_8306);
and U9333 (N_9333,N_8780,N_8210);
and U9334 (N_9334,N_7652,N_8875);
and U9335 (N_9335,N_8729,N_8333);
or U9336 (N_9336,N_7570,N_7644);
or U9337 (N_9337,N_7636,N_7794);
or U9338 (N_9338,N_7750,N_8738);
or U9339 (N_9339,N_8547,N_8677);
nand U9340 (N_9340,N_7870,N_8892);
xor U9341 (N_9341,N_8879,N_8778);
nand U9342 (N_9342,N_8630,N_8323);
nor U9343 (N_9343,N_8884,N_8744);
or U9344 (N_9344,N_7567,N_8609);
and U9345 (N_9345,N_8033,N_7934);
xnor U9346 (N_9346,N_8281,N_7670);
nand U9347 (N_9347,N_8218,N_8347);
and U9348 (N_9348,N_8663,N_7827);
xnor U9349 (N_9349,N_7803,N_7639);
nand U9350 (N_9350,N_7617,N_8276);
xnor U9351 (N_9351,N_8607,N_7685);
xor U9352 (N_9352,N_8313,N_7568);
nor U9353 (N_9353,N_8647,N_7660);
nand U9354 (N_9354,N_8292,N_8731);
or U9355 (N_9355,N_8025,N_8947);
and U9356 (N_9356,N_8950,N_7999);
xor U9357 (N_9357,N_8284,N_8260);
nor U9358 (N_9358,N_7551,N_8833);
nand U9359 (N_9359,N_8122,N_7779);
or U9360 (N_9360,N_8414,N_8571);
nand U9361 (N_9361,N_8679,N_8807);
nand U9362 (N_9362,N_8397,N_8548);
nand U9363 (N_9363,N_7809,N_7603);
xor U9364 (N_9364,N_8998,N_8922);
and U9365 (N_9365,N_8098,N_8544);
nand U9366 (N_9366,N_7651,N_8836);
nor U9367 (N_9367,N_8959,N_8330);
and U9368 (N_9368,N_8624,N_8001);
and U9369 (N_9369,N_8853,N_7840);
and U9370 (N_9370,N_7712,N_7995);
nor U9371 (N_9371,N_7624,N_7611);
and U9372 (N_9372,N_8854,N_8995);
nor U9373 (N_9373,N_8626,N_8654);
and U9374 (N_9374,N_7765,N_8872);
nor U9375 (N_9375,N_8351,N_8042);
nor U9376 (N_9376,N_8496,N_8004);
and U9377 (N_9377,N_8503,N_8597);
xnor U9378 (N_9378,N_7514,N_8088);
nor U9379 (N_9379,N_8161,N_8452);
and U9380 (N_9380,N_8982,N_8338);
nor U9381 (N_9381,N_8432,N_8167);
nor U9382 (N_9382,N_8588,N_8282);
nand U9383 (N_9383,N_8476,N_7835);
nor U9384 (N_9384,N_8247,N_7851);
and U9385 (N_9385,N_8138,N_7876);
or U9386 (N_9386,N_8236,N_7699);
or U9387 (N_9387,N_8901,N_7693);
xor U9388 (N_9388,N_8515,N_8930);
and U9389 (N_9389,N_8874,N_7973);
nand U9390 (N_9390,N_8852,N_8239);
xnor U9391 (N_9391,N_8083,N_8646);
or U9392 (N_9392,N_8839,N_8144);
xnor U9393 (N_9393,N_8185,N_7618);
nor U9394 (N_9394,N_8749,N_7842);
or U9395 (N_9395,N_7703,N_7813);
and U9396 (N_9396,N_8010,N_7745);
xor U9397 (N_9397,N_8606,N_7946);
xor U9398 (N_9398,N_8346,N_8202);
xnor U9399 (N_9399,N_8294,N_7945);
nor U9400 (N_9400,N_7938,N_7557);
nor U9401 (N_9401,N_8039,N_8358);
nor U9402 (N_9402,N_8304,N_7898);
xnor U9403 (N_9403,N_8116,N_8115);
and U9404 (N_9404,N_8789,N_8034);
nor U9405 (N_9405,N_7589,N_8134);
and U9406 (N_9406,N_8444,N_8963);
nor U9407 (N_9407,N_8574,N_8094);
xor U9408 (N_9408,N_7521,N_7606);
or U9409 (N_9409,N_8598,N_8327);
or U9410 (N_9410,N_8104,N_8469);
nand U9411 (N_9411,N_7708,N_7796);
and U9412 (N_9412,N_7772,N_7695);
xnor U9413 (N_9413,N_8348,N_8293);
nand U9414 (N_9414,N_8425,N_7921);
nand U9415 (N_9415,N_8029,N_8026);
or U9416 (N_9416,N_8690,N_8840);
or U9417 (N_9417,N_8197,N_7721);
or U9418 (N_9418,N_7951,N_8680);
or U9419 (N_9419,N_8332,N_8507);
and U9420 (N_9420,N_8808,N_8841);
and U9421 (N_9421,N_8092,N_8421);
nand U9422 (N_9422,N_8201,N_8451);
and U9423 (N_9423,N_8391,N_8166);
and U9424 (N_9424,N_8722,N_7892);
xor U9425 (N_9425,N_8241,N_8994);
or U9426 (N_9426,N_7789,N_7696);
or U9427 (N_9427,N_8366,N_7786);
or U9428 (N_9428,N_7752,N_7626);
and U9429 (N_9429,N_7841,N_7661);
or U9430 (N_9430,N_8991,N_7658);
or U9431 (N_9431,N_8215,N_7659);
xor U9432 (N_9432,N_8923,N_8532);
xnor U9433 (N_9433,N_7867,N_7628);
xnor U9434 (N_9434,N_7654,N_8229);
xnor U9435 (N_9435,N_7578,N_7754);
nand U9436 (N_9436,N_7832,N_7640);
or U9437 (N_9437,N_7713,N_8830);
nor U9438 (N_9438,N_7581,N_7977);
or U9439 (N_9439,N_8091,N_8419);
and U9440 (N_9440,N_8090,N_8801);
nor U9441 (N_9441,N_8946,N_8694);
nand U9442 (N_9442,N_7795,N_7665);
or U9443 (N_9443,N_8283,N_8259);
nand U9444 (N_9444,N_7922,N_8863);
nor U9445 (N_9445,N_7500,N_8245);
xor U9446 (N_9446,N_8370,N_8196);
nor U9447 (N_9447,N_8737,N_8445);
xor U9448 (N_9448,N_8310,N_7594);
xor U9449 (N_9449,N_8558,N_8169);
or U9450 (N_9450,N_8473,N_8373);
and U9451 (N_9451,N_7522,N_7849);
nand U9452 (N_9452,N_8216,N_7549);
nand U9453 (N_9453,N_8301,N_8253);
or U9454 (N_9454,N_7793,N_8470);
xor U9455 (N_9455,N_8492,N_7948);
nor U9456 (N_9456,N_8887,N_8596);
or U9457 (N_9457,N_8023,N_8538);
nand U9458 (N_9458,N_8786,N_7871);
nor U9459 (N_9459,N_8636,N_7975);
and U9460 (N_9460,N_8812,N_7740);
or U9461 (N_9461,N_8266,N_7808);
and U9462 (N_9462,N_8436,N_8405);
xnor U9463 (N_9463,N_7534,N_7769);
xnor U9464 (N_9464,N_8878,N_8871);
xor U9465 (N_9465,N_8981,N_8685);
nand U9466 (N_9466,N_8494,N_8315);
nand U9467 (N_9467,N_8078,N_7763);
nor U9468 (N_9468,N_8400,N_7736);
and U9469 (N_9469,N_8075,N_8895);
xor U9470 (N_9470,N_8217,N_8336);
or U9471 (N_9471,N_7701,N_8803);
nor U9472 (N_9472,N_8804,N_7527);
xor U9473 (N_9473,N_8940,N_8876);
and U9474 (N_9474,N_7681,N_8129);
nor U9475 (N_9475,N_8377,N_7725);
xnor U9476 (N_9476,N_8459,N_8904);
and U9477 (N_9477,N_8894,N_8741);
nor U9478 (N_9478,N_8064,N_8608);
and U9479 (N_9479,N_7683,N_8439);
nand U9480 (N_9480,N_8140,N_8563);
and U9481 (N_9481,N_8069,N_8270);
nand U9482 (N_9482,N_8193,N_8944);
xor U9483 (N_9483,N_8018,N_8989);
and U9484 (N_9484,N_8416,N_8412);
or U9485 (N_9485,N_8269,N_7684);
or U9486 (N_9486,N_8750,N_8676);
nand U9487 (N_9487,N_8032,N_8643);
and U9488 (N_9488,N_8799,N_7565);
xnor U9489 (N_9489,N_8859,N_7533);
xor U9490 (N_9490,N_7612,N_8612);
nand U9491 (N_9491,N_7915,N_7805);
xnor U9492 (N_9492,N_7596,N_8758);
and U9493 (N_9493,N_8424,N_7561);
nand U9494 (N_9494,N_8274,N_8822);
and U9495 (N_9495,N_8485,N_7632);
nand U9496 (N_9496,N_7540,N_8192);
nor U9497 (N_9497,N_7706,N_8969);
nor U9498 (N_9498,N_8513,N_8378);
nand U9499 (N_9499,N_8883,N_7980);
xnor U9500 (N_9500,N_7586,N_7576);
or U9501 (N_9501,N_8454,N_8387);
or U9502 (N_9502,N_8049,N_8510);
or U9503 (N_9503,N_8928,N_7537);
nor U9504 (N_9504,N_7897,N_8739);
nand U9505 (N_9505,N_7759,N_7863);
or U9506 (N_9506,N_7674,N_7982);
or U9507 (N_9507,N_8688,N_8707);
nand U9508 (N_9508,N_7954,N_8406);
or U9509 (N_9509,N_8488,N_8237);
nand U9510 (N_9510,N_8521,N_8106);
nand U9511 (N_9511,N_8834,N_7566);
and U9512 (N_9512,N_8016,N_8953);
nor U9513 (N_9513,N_8986,N_7673);
nor U9514 (N_9514,N_7614,N_7671);
and U9515 (N_9515,N_8668,N_8702);
or U9516 (N_9516,N_8556,N_8003);
xnor U9517 (N_9517,N_8787,N_8752);
xnor U9518 (N_9518,N_8255,N_7735);
nand U9519 (N_9519,N_8061,N_8657);
xor U9520 (N_9520,N_7790,N_8097);
nand U9521 (N_9521,N_7548,N_8785);
xnor U9522 (N_9522,N_8102,N_8450);
nand U9523 (N_9523,N_8468,N_8943);
nand U9524 (N_9524,N_8275,N_8318);
nor U9525 (N_9525,N_8063,N_8481);
and U9526 (N_9526,N_8009,N_7850);
xnor U9527 (N_9527,N_7896,N_8974);
nor U9528 (N_9528,N_8885,N_8649);
nor U9529 (N_9529,N_8299,N_8531);
nand U9530 (N_9530,N_8111,N_7955);
or U9531 (N_9531,N_8824,N_7720);
nand U9532 (N_9532,N_8855,N_8220);
xor U9533 (N_9533,N_8087,N_8867);
nor U9534 (N_9534,N_8479,N_8611);
or U9535 (N_9535,N_8041,N_7964);
and U9536 (N_9536,N_8376,N_7672);
xor U9537 (N_9537,N_8125,N_8105);
nor U9538 (N_9538,N_7885,N_7853);
xnor U9539 (N_9539,N_8748,N_8027);
xnor U9540 (N_9540,N_8291,N_8634);
and U9541 (N_9541,N_7782,N_8533);
nor U9542 (N_9542,N_8258,N_7953);
nand U9543 (N_9543,N_7529,N_8976);
nand U9544 (N_9544,N_8942,N_8784);
nor U9545 (N_9545,N_8219,N_8113);
or U9546 (N_9546,N_8975,N_7893);
xor U9547 (N_9547,N_7747,N_7985);
or U9548 (N_9548,N_7956,N_8820);
nand U9549 (N_9549,N_8081,N_7653);
nand U9550 (N_9550,N_7690,N_8123);
xnor U9551 (N_9551,N_8857,N_8761);
xor U9552 (N_9552,N_8309,N_7675);
nor U9553 (N_9553,N_7732,N_7902);
nand U9554 (N_9554,N_8638,N_8526);
and U9555 (N_9555,N_8456,N_8522);
nand U9556 (N_9556,N_8968,N_8564);
or U9557 (N_9557,N_8374,N_8257);
nor U9558 (N_9558,N_7775,N_8925);
nor U9559 (N_9559,N_8392,N_8882);
or U9560 (N_9560,N_8973,N_7919);
nor U9561 (N_9561,N_8956,N_8777);
xnor U9562 (N_9562,N_8343,N_7707);
nor U9563 (N_9563,N_7806,N_7875);
nand U9564 (N_9564,N_8910,N_8705);
nor U9565 (N_9565,N_8601,N_8203);
or U9566 (N_9566,N_8389,N_8723);
nor U9567 (N_9567,N_7645,N_8692);
xnor U9568 (N_9568,N_8568,N_7584);
nand U9569 (N_9569,N_8600,N_7771);
or U9570 (N_9570,N_8870,N_8295);
and U9571 (N_9571,N_8827,N_7998);
nand U9572 (N_9572,N_8823,N_8395);
and U9573 (N_9573,N_8076,N_8728);
xnor U9574 (N_9574,N_7697,N_8409);
or U9575 (N_9575,N_8610,N_7777);
and U9576 (N_9576,N_8906,N_8530);
or U9577 (N_9577,N_8234,N_8429);
or U9578 (N_9578,N_7572,N_8773);
or U9579 (N_9579,N_7904,N_8591);
or U9580 (N_9580,N_7944,N_8320);
xnor U9581 (N_9581,N_8240,N_7591);
xnor U9582 (N_9582,N_8068,N_7927);
nor U9583 (N_9583,N_7784,N_8363);
nor U9584 (N_9584,N_8096,N_8706);
xor U9585 (N_9585,N_7873,N_8721);
and U9586 (N_9586,N_7751,N_7531);
nand U9587 (N_9587,N_8655,N_8256);
or U9588 (N_9588,N_7891,N_8810);
xor U9589 (N_9589,N_7558,N_8403);
and U9590 (N_9590,N_8156,N_7727);
xor U9591 (N_9591,N_8653,N_8727);
nor U9592 (N_9592,N_8498,N_8350);
nor U9593 (N_9593,N_8577,N_8613);
or U9594 (N_9594,N_8798,N_8578);
nand U9595 (N_9595,N_8659,N_8661);
nand U9596 (N_9596,N_8142,N_8862);
or U9597 (N_9597,N_8847,N_8437);
nand U9598 (N_9598,N_8157,N_7633);
nor U9599 (N_9599,N_7928,N_8137);
or U9600 (N_9600,N_7758,N_8141);
nor U9601 (N_9601,N_8573,N_8453);
and U9602 (N_9602,N_8551,N_7883);
nor U9603 (N_9603,N_8420,N_8030);
and U9604 (N_9604,N_7602,N_8114);
nor U9605 (N_9605,N_7680,N_8062);
xnor U9606 (N_9606,N_8472,N_7829);
or U9607 (N_9607,N_7726,N_7539);
nand U9608 (N_9608,N_8381,N_7524);
xnor U9609 (N_9609,N_8164,N_8307);
or U9610 (N_9610,N_7804,N_8040);
xor U9611 (N_9611,N_8806,N_8719);
nand U9612 (N_9612,N_8401,N_8555);
or U9613 (N_9613,N_8660,N_8529);
nor U9614 (N_9614,N_8334,N_8379);
and U9615 (N_9615,N_8020,N_8013);
nand U9616 (N_9616,N_8344,N_7716);
nor U9617 (N_9617,N_7546,N_8491);
and U9618 (N_9618,N_8251,N_7689);
xor U9619 (N_9619,N_8771,N_8900);
nor U9620 (N_9620,N_8495,N_7536);
or U9621 (N_9621,N_8384,N_8816);
xor U9622 (N_9622,N_8471,N_7872);
nand U9623 (N_9623,N_8408,N_8993);
xnor U9624 (N_9624,N_8242,N_7879);
xnor U9625 (N_9625,N_7783,N_8053);
nor U9626 (N_9626,N_7590,N_7920);
or U9627 (N_9627,N_7774,N_8398);
or U9628 (N_9628,N_8743,N_7924);
nor U9629 (N_9629,N_8952,N_7881);
nand U9630 (N_9630,N_8635,N_8055);
xor U9631 (N_9631,N_8455,N_8678);
nand U9632 (N_9632,N_8698,N_8074);
nand U9633 (N_9633,N_7599,N_7647);
and U9634 (N_9634,N_8843,N_8751);
and U9635 (N_9635,N_7663,N_8535);
and U9636 (N_9636,N_8380,N_8595);
and U9637 (N_9637,N_8254,N_7819);
or U9638 (N_9638,N_8232,N_7976);
xor U9639 (N_9639,N_8873,N_8534);
xnor U9640 (N_9640,N_8656,N_7905);
nor U9641 (N_9641,N_8244,N_8755);
nand U9642 (N_9642,N_8404,N_8423);
and U9643 (N_9643,N_8413,N_7987);
nor U9644 (N_9644,N_8108,N_7949);
and U9645 (N_9645,N_7643,N_7515);
or U9646 (N_9646,N_8866,N_7635);
nor U9647 (N_9647,N_7682,N_7621);
xnor U9648 (N_9648,N_8620,N_7753);
and U9649 (N_9649,N_7917,N_8927);
and U9650 (N_9650,N_8932,N_8067);
nand U9651 (N_9651,N_8199,N_8905);
or U9652 (N_9652,N_8851,N_8604);
nand U9653 (N_9653,N_8086,N_8802);
xor U9654 (N_9654,N_8918,N_8936);
and U9655 (N_9655,N_7668,N_8147);
or U9656 (N_9656,N_8200,N_8553);
or U9657 (N_9657,N_8759,N_8696);
xor U9658 (N_9658,N_7756,N_7770);
nor U9659 (N_9659,N_8567,N_7743);
nand U9660 (N_9660,N_8335,N_8899);
or U9661 (N_9661,N_8779,N_8264);
or U9662 (N_9662,N_7634,N_7504);
nor U9663 (N_9663,N_8158,N_8367);
and U9664 (N_9664,N_7688,N_7530);
and U9665 (N_9665,N_8499,N_8226);
xnor U9666 (N_9666,N_8474,N_8071);
nand U9667 (N_9667,N_8800,N_8222);
or U9668 (N_9668,N_8689,N_7541);
nor U9669 (N_9669,N_7610,N_7966);
nand U9670 (N_9670,N_7502,N_8935);
nor U9671 (N_9671,N_8593,N_8669);
xnor U9672 (N_9672,N_8516,N_8212);
and U9673 (N_9673,N_8224,N_8585);
nand U9674 (N_9674,N_7950,N_7923);
and U9675 (N_9675,N_7957,N_7737);
xor U9676 (N_9676,N_8159,N_8543);
nor U9677 (N_9677,N_8868,N_8112);
xor U9678 (N_9678,N_8119,N_7552);
xnor U9679 (N_9679,N_8109,N_8819);
nand U9680 (N_9680,N_7866,N_8050);
nor U9681 (N_9681,N_7884,N_8431);
nor U9682 (N_9682,N_8052,N_8066);
xnor U9683 (N_9683,N_7664,N_8557);
nand U9684 (N_9684,N_8037,N_8044);
nand U9685 (N_9685,N_8277,N_8774);
xor U9686 (N_9686,N_8110,N_8150);
nor U9687 (N_9687,N_8024,N_8198);
nor U9688 (N_9688,N_7519,N_8183);
and U9689 (N_9689,N_7855,N_7865);
or U9690 (N_9690,N_8912,N_8045);
xnor U9691 (N_9691,N_8190,N_8754);
nand U9692 (N_9692,N_7517,N_7900);
nand U9693 (N_9693,N_7868,N_8357);
and U9694 (N_9694,N_8213,N_8311);
and U9695 (N_9695,N_8541,N_7657);
or U9696 (N_9696,N_8082,N_7766);
and U9697 (N_9697,N_7812,N_8482);
or U9698 (N_9698,N_7741,N_7822);
and U9699 (N_9699,N_7583,N_8983);
nor U9700 (N_9700,N_8422,N_7629);
or U9701 (N_9701,N_8133,N_7935);
nor U9702 (N_9702,N_8172,N_8920);
or U9703 (N_9703,N_8174,N_8038);
and U9704 (N_9704,N_8442,N_8964);
and U9705 (N_9705,N_8035,N_8961);
or U9706 (N_9706,N_8337,N_8618);
or U9707 (N_9707,N_7597,N_8539);
xnor U9708 (N_9708,N_7833,N_8979);
nand U9709 (N_9709,N_8740,N_8505);
or U9710 (N_9710,N_7744,N_8735);
or U9711 (N_9711,N_8407,N_7742);
and U9712 (N_9712,N_7859,N_8701);
or U9713 (N_9713,N_8511,N_8263);
and U9714 (N_9714,N_8006,N_8617);
or U9715 (N_9715,N_7730,N_8163);
nand U9716 (N_9716,N_8651,N_8477);
xor U9717 (N_9717,N_7506,N_8509);
or U9718 (N_9718,N_7818,N_8712);
nor U9719 (N_9719,N_8791,N_7862);
nand U9720 (N_9720,N_8622,N_7650);
nor U9721 (N_9721,N_8145,N_8390);
and U9722 (N_9722,N_7520,N_8580);
and U9723 (N_9723,N_7722,N_8523);
xnor U9724 (N_9724,N_8504,N_7912);
xnor U9725 (N_9725,N_8461,N_8536);
nand U9726 (N_9726,N_8464,N_8628);
and U9727 (N_9727,N_7505,N_8095);
xnor U9728 (N_9728,N_8008,N_7960);
xnor U9729 (N_9729,N_8206,N_8262);
and U9730 (N_9730,N_8945,N_7525);
or U9731 (N_9731,N_8977,N_8966);
xnor U9732 (N_9732,N_7724,N_7709);
and U9733 (N_9733,N_8693,N_8084);
xnor U9734 (N_9734,N_8186,N_8036);
or U9735 (N_9735,N_7579,N_8248);
nand U9736 (N_9736,N_7936,N_7890);
nand U9737 (N_9737,N_8043,N_7943);
nand U9738 (N_9738,N_8587,N_8576);
xnor U9739 (N_9739,N_8501,N_8716);
and U9740 (N_9740,N_7952,N_8831);
xor U9741 (N_9741,N_8674,N_7553);
nor U9742 (N_9742,N_7925,N_8007);
xor U9743 (N_9743,N_8846,N_7574);
nand U9744 (N_9744,N_8797,N_8732);
nand U9745 (N_9745,N_8837,N_8768);
or U9746 (N_9746,N_7888,N_8149);
nor U9747 (N_9747,N_8352,N_8849);
xor U9748 (N_9748,N_7799,N_8182);
and U9749 (N_9749,N_7608,N_7785);
and U9750 (N_9750,N_8640,N_8209);
nand U9751 (N_9751,N_8924,N_7655);
nand U9752 (N_9752,N_8083,N_7838);
nor U9753 (N_9753,N_8670,N_8062);
or U9754 (N_9754,N_7969,N_8385);
and U9755 (N_9755,N_7630,N_7638);
xnor U9756 (N_9756,N_7701,N_8304);
and U9757 (N_9757,N_7726,N_8840);
nand U9758 (N_9758,N_7892,N_8815);
xnor U9759 (N_9759,N_8664,N_7670);
nor U9760 (N_9760,N_7502,N_7824);
xor U9761 (N_9761,N_8793,N_8988);
or U9762 (N_9762,N_8666,N_8965);
or U9763 (N_9763,N_8181,N_8580);
and U9764 (N_9764,N_8283,N_7542);
nor U9765 (N_9765,N_8688,N_7558);
xnor U9766 (N_9766,N_7624,N_8259);
and U9767 (N_9767,N_8020,N_7520);
or U9768 (N_9768,N_8010,N_7647);
or U9769 (N_9769,N_8464,N_8803);
xor U9770 (N_9770,N_8033,N_7512);
nand U9771 (N_9771,N_8990,N_7975);
or U9772 (N_9772,N_7625,N_8536);
or U9773 (N_9773,N_8811,N_8869);
nand U9774 (N_9774,N_7800,N_7718);
nor U9775 (N_9775,N_7653,N_8782);
or U9776 (N_9776,N_7560,N_7793);
nand U9777 (N_9777,N_8092,N_8625);
nand U9778 (N_9778,N_8544,N_8692);
nor U9779 (N_9779,N_8498,N_7507);
and U9780 (N_9780,N_8434,N_7527);
and U9781 (N_9781,N_8628,N_7741);
and U9782 (N_9782,N_8114,N_8773);
xnor U9783 (N_9783,N_8277,N_8969);
nand U9784 (N_9784,N_8470,N_8033);
and U9785 (N_9785,N_8312,N_7658);
nand U9786 (N_9786,N_7921,N_7896);
or U9787 (N_9787,N_8787,N_8014);
or U9788 (N_9788,N_8081,N_8748);
and U9789 (N_9789,N_8324,N_8876);
nand U9790 (N_9790,N_7781,N_8969);
xnor U9791 (N_9791,N_8172,N_8378);
and U9792 (N_9792,N_7766,N_7634);
and U9793 (N_9793,N_7878,N_7848);
and U9794 (N_9794,N_8652,N_7662);
nand U9795 (N_9795,N_8105,N_7862);
and U9796 (N_9796,N_8860,N_8916);
xnor U9797 (N_9797,N_8036,N_7839);
nand U9798 (N_9798,N_8298,N_8463);
nor U9799 (N_9799,N_8271,N_8325);
or U9800 (N_9800,N_8051,N_8527);
and U9801 (N_9801,N_8974,N_8600);
and U9802 (N_9802,N_7860,N_8541);
nand U9803 (N_9803,N_8691,N_8113);
nor U9804 (N_9804,N_8960,N_8551);
xnor U9805 (N_9805,N_7704,N_8036);
or U9806 (N_9806,N_7854,N_8544);
or U9807 (N_9807,N_8673,N_8543);
nand U9808 (N_9808,N_8867,N_8960);
xor U9809 (N_9809,N_8259,N_7902);
and U9810 (N_9810,N_8327,N_7915);
nand U9811 (N_9811,N_8269,N_7870);
nor U9812 (N_9812,N_8197,N_8365);
nor U9813 (N_9813,N_8741,N_8270);
and U9814 (N_9814,N_8590,N_8803);
xor U9815 (N_9815,N_7603,N_7619);
nand U9816 (N_9816,N_8485,N_8526);
xnor U9817 (N_9817,N_8501,N_8865);
nand U9818 (N_9818,N_8036,N_8090);
and U9819 (N_9819,N_8501,N_8934);
and U9820 (N_9820,N_8692,N_7798);
or U9821 (N_9821,N_8146,N_8075);
or U9822 (N_9822,N_8739,N_7953);
or U9823 (N_9823,N_8535,N_8252);
or U9824 (N_9824,N_8402,N_7606);
xor U9825 (N_9825,N_8047,N_8301);
nand U9826 (N_9826,N_8870,N_7934);
nand U9827 (N_9827,N_8625,N_7531);
nor U9828 (N_9828,N_8214,N_7928);
and U9829 (N_9829,N_8262,N_8039);
nor U9830 (N_9830,N_8385,N_7819);
nand U9831 (N_9831,N_8285,N_8091);
and U9832 (N_9832,N_8253,N_8975);
nor U9833 (N_9833,N_8461,N_7633);
nand U9834 (N_9834,N_8178,N_7663);
nor U9835 (N_9835,N_8892,N_7755);
nor U9836 (N_9836,N_8754,N_8270);
and U9837 (N_9837,N_7939,N_7682);
nand U9838 (N_9838,N_8969,N_8485);
and U9839 (N_9839,N_8604,N_7528);
nor U9840 (N_9840,N_7642,N_8122);
and U9841 (N_9841,N_8141,N_8948);
nor U9842 (N_9842,N_8902,N_8347);
or U9843 (N_9843,N_7903,N_8417);
xnor U9844 (N_9844,N_7580,N_8381);
nor U9845 (N_9845,N_8092,N_8357);
and U9846 (N_9846,N_7600,N_8147);
or U9847 (N_9847,N_8103,N_7852);
or U9848 (N_9848,N_7975,N_8442);
nand U9849 (N_9849,N_7894,N_7659);
xnor U9850 (N_9850,N_7876,N_8114);
and U9851 (N_9851,N_7836,N_7667);
or U9852 (N_9852,N_8721,N_8404);
and U9853 (N_9853,N_8898,N_7791);
xor U9854 (N_9854,N_8065,N_8617);
or U9855 (N_9855,N_8709,N_8830);
or U9856 (N_9856,N_7998,N_8484);
nor U9857 (N_9857,N_8305,N_7954);
xor U9858 (N_9858,N_7924,N_8396);
and U9859 (N_9859,N_8522,N_7845);
nor U9860 (N_9860,N_8586,N_7933);
nor U9861 (N_9861,N_8423,N_8018);
nor U9862 (N_9862,N_8398,N_8568);
nand U9863 (N_9863,N_7516,N_8290);
and U9864 (N_9864,N_7568,N_8201);
nand U9865 (N_9865,N_8171,N_7552);
and U9866 (N_9866,N_8002,N_8915);
nor U9867 (N_9867,N_8465,N_8907);
xor U9868 (N_9868,N_8858,N_8609);
nand U9869 (N_9869,N_7762,N_8139);
nand U9870 (N_9870,N_8247,N_8741);
nand U9871 (N_9871,N_8805,N_8989);
or U9872 (N_9872,N_8469,N_8086);
or U9873 (N_9873,N_8094,N_8280);
or U9874 (N_9874,N_8721,N_7786);
nor U9875 (N_9875,N_7912,N_8568);
nor U9876 (N_9876,N_8967,N_7657);
or U9877 (N_9877,N_7589,N_7895);
nand U9878 (N_9878,N_7879,N_8936);
xor U9879 (N_9879,N_8199,N_8228);
nand U9880 (N_9880,N_8596,N_8275);
and U9881 (N_9881,N_7524,N_8558);
xnor U9882 (N_9882,N_8291,N_8374);
nor U9883 (N_9883,N_8494,N_8046);
nand U9884 (N_9884,N_8931,N_8682);
xor U9885 (N_9885,N_7679,N_8955);
or U9886 (N_9886,N_8562,N_8055);
nor U9887 (N_9887,N_8927,N_8633);
nor U9888 (N_9888,N_8255,N_8857);
nand U9889 (N_9889,N_7602,N_7786);
xor U9890 (N_9890,N_7516,N_8172);
nor U9891 (N_9891,N_8028,N_7597);
nand U9892 (N_9892,N_7578,N_8327);
and U9893 (N_9893,N_8144,N_7888);
and U9894 (N_9894,N_8130,N_8958);
and U9895 (N_9895,N_7571,N_8924);
or U9896 (N_9896,N_8212,N_7846);
nand U9897 (N_9897,N_7682,N_7575);
and U9898 (N_9898,N_7589,N_7867);
nor U9899 (N_9899,N_7930,N_8783);
and U9900 (N_9900,N_8886,N_8150);
and U9901 (N_9901,N_7847,N_8704);
nor U9902 (N_9902,N_8326,N_8350);
nand U9903 (N_9903,N_7871,N_8290);
nor U9904 (N_9904,N_8124,N_8907);
and U9905 (N_9905,N_8438,N_7510);
or U9906 (N_9906,N_8827,N_8106);
xnor U9907 (N_9907,N_8592,N_8608);
nor U9908 (N_9908,N_8319,N_8053);
and U9909 (N_9909,N_8667,N_7794);
or U9910 (N_9910,N_8503,N_8742);
and U9911 (N_9911,N_8100,N_8824);
nand U9912 (N_9912,N_8675,N_8697);
nand U9913 (N_9913,N_8091,N_7892);
xor U9914 (N_9914,N_7579,N_8310);
and U9915 (N_9915,N_8978,N_8422);
or U9916 (N_9916,N_7714,N_8514);
xnor U9917 (N_9917,N_8277,N_8323);
and U9918 (N_9918,N_7552,N_8194);
nand U9919 (N_9919,N_8324,N_8368);
or U9920 (N_9920,N_8457,N_8473);
or U9921 (N_9921,N_8340,N_7955);
and U9922 (N_9922,N_7651,N_8325);
nor U9923 (N_9923,N_8568,N_8030);
nand U9924 (N_9924,N_8761,N_8548);
and U9925 (N_9925,N_8159,N_7657);
and U9926 (N_9926,N_8803,N_8157);
xnor U9927 (N_9927,N_8079,N_8392);
nor U9928 (N_9928,N_8192,N_8828);
and U9929 (N_9929,N_7751,N_7778);
or U9930 (N_9930,N_8823,N_7842);
xor U9931 (N_9931,N_8328,N_8574);
nor U9932 (N_9932,N_7949,N_8605);
or U9933 (N_9933,N_8362,N_7591);
xor U9934 (N_9934,N_7967,N_8167);
nand U9935 (N_9935,N_8032,N_8091);
xnor U9936 (N_9936,N_8124,N_8691);
nor U9937 (N_9937,N_8060,N_7710);
nor U9938 (N_9938,N_8670,N_8033);
nand U9939 (N_9939,N_7665,N_8607);
nand U9940 (N_9940,N_7633,N_8814);
and U9941 (N_9941,N_7852,N_8089);
nor U9942 (N_9942,N_8740,N_8295);
xor U9943 (N_9943,N_8596,N_7734);
and U9944 (N_9944,N_8167,N_8328);
and U9945 (N_9945,N_7617,N_8975);
or U9946 (N_9946,N_7930,N_8886);
nor U9947 (N_9947,N_8741,N_8415);
nand U9948 (N_9948,N_7533,N_7644);
xnor U9949 (N_9949,N_8455,N_7564);
nor U9950 (N_9950,N_8358,N_8875);
or U9951 (N_9951,N_8619,N_7892);
xnor U9952 (N_9952,N_7759,N_8832);
nand U9953 (N_9953,N_7652,N_8885);
nor U9954 (N_9954,N_7944,N_7831);
nand U9955 (N_9955,N_7653,N_8741);
xnor U9956 (N_9956,N_7920,N_7999);
nor U9957 (N_9957,N_8423,N_7898);
nor U9958 (N_9958,N_7895,N_8126);
nor U9959 (N_9959,N_8948,N_8829);
xor U9960 (N_9960,N_8174,N_7611);
nor U9961 (N_9961,N_7616,N_8520);
or U9962 (N_9962,N_7943,N_8024);
or U9963 (N_9963,N_8942,N_8192);
xnor U9964 (N_9964,N_8738,N_8414);
or U9965 (N_9965,N_8456,N_8723);
nor U9966 (N_9966,N_8156,N_8204);
nor U9967 (N_9967,N_8539,N_8200);
nor U9968 (N_9968,N_8489,N_8274);
or U9969 (N_9969,N_7985,N_8555);
nor U9970 (N_9970,N_8633,N_8478);
or U9971 (N_9971,N_7573,N_8302);
xor U9972 (N_9972,N_8662,N_7640);
or U9973 (N_9973,N_8331,N_7835);
or U9974 (N_9974,N_8473,N_7725);
nand U9975 (N_9975,N_8199,N_8841);
and U9976 (N_9976,N_8644,N_8480);
xnor U9977 (N_9977,N_7967,N_8197);
or U9978 (N_9978,N_8894,N_8214);
nor U9979 (N_9979,N_8269,N_8482);
nor U9980 (N_9980,N_8379,N_7840);
nor U9981 (N_9981,N_8834,N_8443);
nand U9982 (N_9982,N_8840,N_7550);
xnor U9983 (N_9983,N_7807,N_8371);
xnor U9984 (N_9984,N_7931,N_7886);
xor U9985 (N_9985,N_7847,N_8371);
nor U9986 (N_9986,N_8998,N_7785);
xor U9987 (N_9987,N_8885,N_8729);
nor U9988 (N_9988,N_7639,N_8115);
xnor U9989 (N_9989,N_7929,N_8230);
nand U9990 (N_9990,N_8155,N_7900);
or U9991 (N_9991,N_8903,N_7631);
nand U9992 (N_9992,N_8120,N_8175);
nor U9993 (N_9993,N_8903,N_7938);
xnor U9994 (N_9994,N_8285,N_7756);
and U9995 (N_9995,N_8375,N_7823);
xnor U9996 (N_9996,N_7990,N_7913);
xor U9997 (N_9997,N_8043,N_8024);
nor U9998 (N_9998,N_8795,N_8661);
or U9999 (N_9999,N_8698,N_8368);
nand U10000 (N_10000,N_8201,N_7768);
nor U10001 (N_10001,N_7902,N_7803);
and U10002 (N_10002,N_7605,N_8321);
or U10003 (N_10003,N_7761,N_8078);
or U10004 (N_10004,N_7723,N_8307);
and U10005 (N_10005,N_7917,N_8605);
xnor U10006 (N_10006,N_8949,N_8699);
nor U10007 (N_10007,N_8036,N_8284);
nor U10008 (N_10008,N_8745,N_8189);
xor U10009 (N_10009,N_7530,N_8367);
or U10010 (N_10010,N_8179,N_8543);
nor U10011 (N_10011,N_7631,N_7668);
and U10012 (N_10012,N_8249,N_8401);
xnor U10013 (N_10013,N_8903,N_8853);
nand U10014 (N_10014,N_7898,N_8922);
nor U10015 (N_10015,N_8501,N_7689);
and U10016 (N_10016,N_8123,N_8769);
nor U10017 (N_10017,N_8310,N_8189);
nor U10018 (N_10018,N_7584,N_8569);
and U10019 (N_10019,N_8630,N_7577);
or U10020 (N_10020,N_7657,N_7781);
nor U10021 (N_10021,N_7614,N_8093);
or U10022 (N_10022,N_8708,N_7580);
nor U10023 (N_10023,N_7811,N_8332);
nand U10024 (N_10024,N_8927,N_8404);
xor U10025 (N_10025,N_7605,N_8612);
nor U10026 (N_10026,N_8776,N_7663);
nor U10027 (N_10027,N_7905,N_8865);
or U10028 (N_10028,N_8131,N_8218);
and U10029 (N_10029,N_8355,N_7608);
xnor U10030 (N_10030,N_7506,N_8381);
nand U10031 (N_10031,N_7749,N_8344);
xor U10032 (N_10032,N_7836,N_8900);
or U10033 (N_10033,N_8154,N_7929);
nor U10034 (N_10034,N_8509,N_8407);
or U10035 (N_10035,N_8087,N_7915);
nor U10036 (N_10036,N_8363,N_7681);
or U10037 (N_10037,N_8116,N_8156);
or U10038 (N_10038,N_8011,N_8007);
and U10039 (N_10039,N_7686,N_7966);
xnor U10040 (N_10040,N_7558,N_8157);
and U10041 (N_10041,N_8095,N_8455);
nand U10042 (N_10042,N_7633,N_7541);
nand U10043 (N_10043,N_8928,N_8600);
xnor U10044 (N_10044,N_7838,N_8072);
nor U10045 (N_10045,N_8613,N_8091);
or U10046 (N_10046,N_7646,N_8035);
nand U10047 (N_10047,N_7539,N_8440);
nor U10048 (N_10048,N_7548,N_8358);
xor U10049 (N_10049,N_8512,N_8267);
or U10050 (N_10050,N_8815,N_7698);
and U10051 (N_10051,N_7630,N_7682);
xnor U10052 (N_10052,N_7903,N_8837);
or U10053 (N_10053,N_7946,N_7935);
nand U10054 (N_10054,N_8372,N_8058);
nor U10055 (N_10055,N_7507,N_8115);
or U10056 (N_10056,N_8647,N_8357);
xnor U10057 (N_10057,N_7678,N_7818);
xor U10058 (N_10058,N_8400,N_8321);
nor U10059 (N_10059,N_8204,N_8858);
xor U10060 (N_10060,N_7696,N_7931);
and U10061 (N_10061,N_8070,N_7705);
xnor U10062 (N_10062,N_7818,N_8648);
or U10063 (N_10063,N_8629,N_8172);
or U10064 (N_10064,N_8360,N_8601);
or U10065 (N_10065,N_8522,N_8881);
and U10066 (N_10066,N_8208,N_8277);
or U10067 (N_10067,N_7581,N_8180);
and U10068 (N_10068,N_7767,N_7956);
nor U10069 (N_10069,N_8050,N_7821);
and U10070 (N_10070,N_7964,N_8238);
nand U10071 (N_10071,N_8913,N_8168);
or U10072 (N_10072,N_7930,N_7995);
nand U10073 (N_10073,N_8339,N_8830);
nor U10074 (N_10074,N_7655,N_8666);
nand U10075 (N_10075,N_7937,N_7993);
or U10076 (N_10076,N_7976,N_8980);
nor U10077 (N_10077,N_7965,N_8060);
or U10078 (N_10078,N_7593,N_7869);
or U10079 (N_10079,N_8642,N_8777);
xor U10080 (N_10080,N_8321,N_8167);
or U10081 (N_10081,N_7590,N_8051);
or U10082 (N_10082,N_8267,N_7925);
and U10083 (N_10083,N_8685,N_8723);
nand U10084 (N_10084,N_8081,N_7816);
xor U10085 (N_10085,N_8250,N_8879);
or U10086 (N_10086,N_8207,N_7717);
or U10087 (N_10087,N_7763,N_8985);
or U10088 (N_10088,N_7596,N_7645);
xor U10089 (N_10089,N_8012,N_8858);
and U10090 (N_10090,N_8221,N_8696);
nand U10091 (N_10091,N_8686,N_7701);
and U10092 (N_10092,N_8320,N_8838);
or U10093 (N_10093,N_7592,N_8920);
nand U10094 (N_10094,N_8006,N_8738);
nand U10095 (N_10095,N_7755,N_7839);
xor U10096 (N_10096,N_8686,N_8335);
xnor U10097 (N_10097,N_7773,N_7812);
or U10098 (N_10098,N_7513,N_8052);
nand U10099 (N_10099,N_8901,N_8589);
and U10100 (N_10100,N_8034,N_7733);
nor U10101 (N_10101,N_8712,N_8362);
nor U10102 (N_10102,N_7974,N_8769);
and U10103 (N_10103,N_8373,N_8568);
xor U10104 (N_10104,N_8775,N_7578);
xnor U10105 (N_10105,N_8845,N_8960);
nor U10106 (N_10106,N_7502,N_8458);
and U10107 (N_10107,N_8628,N_8890);
nor U10108 (N_10108,N_8657,N_8502);
or U10109 (N_10109,N_7589,N_8336);
and U10110 (N_10110,N_7531,N_8506);
and U10111 (N_10111,N_8520,N_8462);
nand U10112 (N_10112,N_8660,N_8499);
nand U10113 (N_10113,N_8051,N_7900);
nor U10114 (N_10114,N_7741,N_8953);
nand U10115 (N_10115,N_7536,N_8189);
xor U10116 (N_10116,N_7523,N_8924);
nand U10117 (N_10117,N_7509,N_7658);
xor U10118 (N_10118,N_8220,N_8973);
or U10119 (N_10119,N_8037,N_8839);
xnor U10120 (N_10120,N_8747,N_8344);
nand U10121 (N_10121,N_8825,N_8775);
and U10122 (N_10122,N_8134,N_7744);
and U10123 (N_10123,N_7849,N_8167);
nor U10124 (N_10124,N_7539,N_7671);
nor U10125 (N_10125,N_7962,N_8050);
nor U10126 (N_10126,N_8885,N_8156);
and U10127 (N_10127,N_7764,N_7579);
nor U10128 (N_10128,N_7639,N_7962);
xnor U10129 (N_10129,N_8114,N_7689);
nand U10130 (N_10130,N_7619,N_8865);
and U10131 (N_10131,N_8674,N_8184);
or U10132 (N_10132,N_8468,N_8110);
nand U10133 (N_10133,N_7816,N_8176);
xnor U10134 (N_10134,N_8564,N_8072);
or U10135 (N_10135,N_8932,N_8844);
and U10136 (N_10136,N_8338,N_8340);
xor U10137 (N_10137,N_8118,N_8330);
xor U10138 (N_10138,N_8499,N_7727);
or U10139 (N_10139,N_7941,N_8207);
and U10140 (N_10140,N_8272,N_8411);
xor U10141 (N_10141,N_8965,N_7894);
nand U10142 (N_10142,N_8139,N_8799);
nand U10143 (N_10143,N_8184,N_8466);
nand U10144 (N_10144,N_8027,N_8753);
xor U10145 (N_10145,N_7792,N_7903);
or U10146 (N_10146,N_8648,N_7770);
xnor U10147 (N_10147,N_7657,N_8457);
nor U10148 (N_10148,N_8017,N_8964);
xor U10149 (N_10149,N_7788,N_8314);
xor U10150 (N_10150,N_7798,N_8243);
nand U10151 (N_10151,N_7650,N_8776);
or U10152 (N_10152,N_7506,N_8856);
nand U10153 (N_10153,N_8524,N_7562);
and U10154 (N_10154,N_7721,N_8981);
nor U10155 (N_10155,N_8589,N_7780);
nand U10156 (N_10156,N_8668,N_8474);
nor U10157 (N_10157,N_8236,N_7692);
and U10158 (N_10158,N_8493,N_8179);
or U10159 (N_10159,N_8064,N_8455);
and U10160 (N_10160,N_7564,N_8321);
nor U10161 (N_10161,N_7869,N_8222);
and U10162 (N_10162,N_7557,N_7504);
and U10163 (N_10163,N_8652,N_7599);
nor U10164 (N_10164,N_7689,N_7754);
nor U10165 (N_10165,N_7927,N_8655);
and U10166 (N_10166,N_7624,N_8621);
and U10167 (N_10167,N_8457,N_7797);
and U10168 (N_10168,N_7869,N_8361);
or U10169 (N_10169,N_8513,N_8273);
and U10170 (N_10170,N_8531,N_8586);
and U10171 (N_10171,N_7550,N_8467);
nor U10172 (N_10172,N_8954,N_8980);
or U10173 (N_10173,N_8249,N_8503);
and U10174 (N_10174,N_8936,N_7627);
nand U10175 (N_10175,N_8910,N_8275);
nor U10176 (N_10176,N_8279,N_8386);
or U10177 (N_10177,N_7827,N_8847);
xor U10178 (N_10178,N_7789,N_8702);
nand U10179 (N_10179,N_7953,N_8654);
or U10180 (N_10180,N_7747,N_7790);
nor U10181 (N_10181,N_8501,N_7824);
nand U10182 (N_10182,N_8080,N_8301);
nor U10183 (N_10183,N_7593,N_7895);
or U10184 (N_10184,N_8673,N_8986);
xor U10185 (N_10185,N_8050,N_8188);
nor U10186 (N_10186,N_8326,N_8898);
and U10187 (N_10187,N_7501,N_7660);
nand U10188 (N_10188,N_8916,N_7902);
and U10189 (N_10189,N_8603,N_8274);
xnor U10190 (N_10190,N_8998,N_8913);
xor U10191 (N_10191,N_8255,N_7775);
nand U10192 (N_10192,N_8528,N_8224);
xnor U10193 (N_10193,N_8198,N_7804);
or U10194 (N_10194,N_8042,N_7689);
or U10195 (N_10195,N_7687,N_7668);
or U10196 (N_10196,N_8795,N_8173);
and U10197 (N_10197,N_8268,N_8023);
nand U10198 (N_10198,N_8327,N_8226);
and U10199 (N_10199,N_7700,N_8551);
nand U10200 (N_10200,N_7606,N_8098);
or U10201 (N_10201,N_8880,N_8101);
and U10202 (N_10202,N_7737,N_8342);
nor U10203 (N_10203,N_8550,N_8641);
xor U10204 (N_10204,N_8199,N_7634);
and U10205 (N_10205,N_7970,N_7847);
or U10206 (N_10206,N_8953,N_7687);
and U10207 (N_10207,N_8820,N_8355);
nor U10208 (N_10208,N_7897,N_7808);
and U10209 (N_10209,N_8718,N_8505);
nand U10210 (N_10210,N_8996,N_7838);
and U10211 (N_10211,N_8696,N_7723);
nand U10212 (N_10212,N_8523,N_8377);
xnor U10213 (N_10213,N_8776,N_8131);
nor U10214 (N_10214,N_8734,N_8483);
xnor U10215 (N_10215,N_8114,N_8087);
xnor U10216 (N_10216,N_8534,N_8402);
and U10217 (N_10217,N_8647,N_8314);
and U10218 (N_10218,N_8155,N_8194);
nor U10219 (N_10219,N_8979,N_8094);
and U10220 (N_10220,N_8295,N_8519);
or U10221 (N_10221,N_7704,N_8909);
and U10222 (N_10222,N_8041,N_7818);
nor U10223 (N_10223,N_8084,N_7828);
or U10224 (N_10224,N_8654,N_8197);
or U10225 (N_10225,N_7696,N_8521);
or U10226 (N_10226,N_8674,N_8698);
xnor U10227 (N_10227,N_7563,N_7540);
or U10228 (N_10228,N_7954,N_7759);
and U10229 (N_10229,N_8636,N_8219);
nand U10230 (N_10230,N_8807,N_7646);
nor U10231 (N_10231,N_8724,N_7679);
nor U10232 (N_10232,N_8412,N_7721);
or U10233 (N_10233,N_8097,N_7620);
xor U10234 (N_10234,N_8903,N_8108);
xnor U10235 (N_10235,N_8875,N_7907);
nand U10236 (N_10236,N_8420,N_8696);
nand U10237 (N_10237,N_8808,N_7860);
xnor U10238 (N_10238,N_8402,N_7703);
or U10239 (N_10239,N_8920,N_8635);
nand U10240 (N_10240,N_7884,N_8854);
xnor U10241 (N_10241,N_8633,N_7892);
xor U10242 (N_10242,N_8642,N_8140);
nor U10243 (N_10243,N_8755,N_8255);
xnor U10244 (N_10244,N_8013,N_7588);
nand U10245 (N_10245,N_8668,N_8954);
nor U10246 (N_10246,N_8827,N_7969);
nand U10247 (N_10247,N_8996,N_8377);
and U10248 (N_10248,N_8600,N_8963);
and U10249 (N_10249,N_8344,N_7678);
nor U10250 (N_10250,N_8302,N_7936);
or U10251 (N_10251,N_8816,N_8669);
nand U10252 (N_10252,N_7656,N_7950);
and U10253 (N_10253,N_8097,N_8381);
xor U10254 (N_10254,N_8578,N_8358);
xnor U10255 (N_10255,N_8018,N_8780);
and U10256 (N_10256,N_8012,N_7603);
nor U10257 (N_10257,N_8772,N_7787);
nand U10258 (N_10258,N_8124,N_8266);
xnor U10259 (N_10259,N_8273,N_7516);
xnor U10260 (N_10260,N_8883,N_7639);
or U10261 (N_10261,N_8675,N_8009);
xnor U10262 (N_10262,N_7758,N_8995);
and U10263 (N_10263,N_8598,N_8193);
and U10264 (N_10264,N_8348,N_7559);
xor U10265 (N_10265,N_8985,N_8635);
xor U10266 (N_10266,N_7677,N_8245);
nand U10267 (N_10267,N_7972,N_8534);
and U10268 (N_10268,N_7574,N_8996);
nand U10269 (N_10269,N_8010,N_8359);
and U10270 (N_10270,N_8099,N_8645);
nor U10271 (N_10271,N_8063,N_7667);
or U10272 (N_10272,N_8538,N_7796);
nor U10273 (N_10273,N_8808,N_8921);
or U10274 (N_10274,N_8851,N_7984);
nor U10275 (N_10275,N_8865,N_8822);
and U10276 (N_10276,N_8239,N_7970);
nand U10277 (N_10277,N_8846,N_7863);
or U10278 (N_10278,N_8901,N_8970);
nand U10279 (N_10279,N_7644,N_7616);
nor U10280 (N_10280,N_8191,N_8808);
xor U10281 (N_10281,N_8099,N_7699);
or U10282 (N_10282,N_8440,N_7845);
and U10283 (N_10283,N_8199,N_8969);
xnor U10284 (N_10284,N_8434,N_7728);
nand U10285 (N_10285,N_8092,N_8259);
nor U10286 (N_10286,N_8538,N_8452);
nand U10287 (N_10287,N_8494,N_7891);
and U10288 (N_10288,N_8791,N_8302);
nand U10289 (N_10289,N_7729,N_7628);
or U10290 (N_10290,N_8967,N_8248);
and U10291 (N_10291,N_8051,N_8013);
xor U10292 (N_10292,N_8980,N_8885);
and U10293 (N_10293,N_7895,N_8112);
or U10294 (N_10294,N_8169,N_8050);
and U10295 (N_10295,N_7849,N_8964);
and U10296 (N_10296,N_8038,N_8217);
or U10297 (N_10297,N_8613,N_7704);
and U10298 (N_10298,N_8612,N_8557);
xnor U10299 (N_10299,N_8879,N_8716);
nand U10300 (N_10300,N_8804,N_7866);
or U10301 (N_10301,N_8071,N_8386);
nand U10302 (N_10302,N_8848,N_8842);
nor U10303 (N_10303,N_7620,N_8749);
xnor U10304 (N_10304,N_8016,N_8756);
nor U10305 (N_10305,N_7665,N_8356);
and U10306 (N_10306,N_7665,N_8253);
nand U10307 (N_10307,N_8338,N_8455);
nor U10308 (N_10308,N_8540,N_8062);
nor U10309 (N_10309,N_7523,N_7531);
nor U10310 (N_10310,N_7786,N_7944);
xnor U10311 (N_10311,N_8820,N_8837);
nand U10312 (N_10312,N_8732,N_8692);
nand U10313 (N_10313,N_8730,N_7851);
nor U10314 (N_10314,N_7824,N_7954);
xor U10315 (N_10315,N_8167,N_8098);
nor U10316 (N_10316,N_8146,N_8989);
nand U10317 (N_10317,N_8305,N_8719);
nor U10318 (N_10318,N_8851,N_8427);
or U10319 (N_10319,N_8180,N_8373);
nor U10320 (N_10320,N_8415,N_7856);
xnor U10321 (N_10321,N_8737,N_8374);
or U10322 (N_10322,N_8155,N_8091);
nand U10323 (N_10323,N_8968,N_8214);
or U10324 (N_10324,N_7615,N_8660);
and U10325 (N_10325,N_8908,N_7545);
nand U10326 (N_10326,N_8010,N_8000);
and U10327 (N_10327,N_8876,N_7932);
nand U10328 (N_10328,N_8068,N_8768);
nor U10329 (N_10329,N_7955,N_8170);
nor U10330 (N_10330,N_8553,N_8490);
and U10331 (N_10331,N_7910,N_8667);
or U10332 (N_10332,N_8267,N_7868);
nor U10333 (N_10333,N_8782,N_7689);
nand U10334 (N_10334,N_7733,N_8798);
and U10335 (N_10335,N_7778,N_8468);
or U10336 (N_10336,N_8134,N_8709);
nand U10337 (N_10337,N_8201,N_7605);
and U10338 (N_10338,N_8890,N_8195);
and U10339 (N_10339,N_7751,N_8355);
xnor U10340 (N_10340,N_7858,N_8835);
nand U10341 (N_10341,N_8401,N_7671);
or U10342 (N_10342,N_8896,N_8043);
or U10343 (N_10343,N_7741,N_7616);
nand U10344 (N_10344,N_8396,N_8722);
nand U10345 (N_10345,N_8804,N_7785);
xnor U10346 (N_10346,N_8014,N_8020);
nand U10347 (N_10347,N_8764,N_8160);
nor U10348 (N_10348,N_8408,N_8266);
nand U10349 (N_10349,N_8691,N_7819);
nand U10350 (N_10350,N_7708,N_8613);
nor U10351 (N_10351,N_7865,N_8997);
nor U10352 (N_10352,N_8429,N_8962);
or U10353 (N_10353,N_8676,N_8654);
nand U10354 (N_10354,N_8407,N_8833);
nand U10355 (N_10355,N_8189,N_7847);
or U10356 (N_10356,N_8934,N_7567);
and U10357 (N_10357,N_8988,N_8269);
xnor U10358 (N_10358,N_8036,N_8941);
xor U10359 (N_10359,N_7689,N_8737);
xnor U10360 (N_10360,N_7605,N_8003);
and U10361 (N_10361,N_8368,N_8149);
or U10362 (N_10362,N_7750,N_8330);
nor U10363 (N_10363,N_8000,N_8649);
nand U10364 (N_10364,N_7911,N_8349);
xnor U10365 (N_10365,N_8552,N_7919);
and U10366 (N_10366,N_8998,N_8765);
and U10367 (N_10367,N_8499,N_8752);
nand U10368 (N_10368,N_8916,N_8465);
or U10369 (N_10369,N_8352,N_8017);
nor U10370 (N_10370,N_8761,N_8047);
nand U10371 (N_10371,N_8772,N_7868);
nand U10372 (N_10372,N_7753,N_8481);
nand U10373 (N_10373,N_7634,N_8108);
nor U10374 (N_10374,N_7625,N_8125);
xor U10375 (N_10375,N_8881,N_7659);
nor U10376 (N_10376,N_8949,N_8538);
or U10377 (N_10377,N_8835,N_7998);
xnor U10378 (N_10378,N_8137,N_7706);
and U10379 (N_10379,N_8761,N_7571);
nand U10380 (N_10380,N_8497,N_8087);
nor U10381 (N_10381,N_8168,N_8671);
nand U10382 (N_10382,N_8643,N_8114);
or U10383 (N_10383,N_8013,N_8228);
xor U10384 (N_10384,N_7778,N_7660);
nand U10385 (N_10385,N_8517,N_8687);
nor U10386 (N_10386,N_8383,N_8853);
nor U10387 (N_10387,N_8895,N_8059);
xnor U10388 (N_10388,N_8453,N_8885);
and U10389 (N_10389,N_8788,N_8246);
or U10390 (N_10390,N_7615,N_7579);
and U10391 (N_10391,N_8701,N_7786);
nand U10392 (N_10392,N_8039,N_8176);
xor U10393 (N_10393,N_7725,N_8307);
nor U10394 (N_10394,N_7842,N_7714);
xnor U10395 (N_10395,N_8999,N_8523);
or U10396 (N_10396,N_8039,N_8446);
xor U10397 (N_10397,N_7965,N_8626);
and U10398 (N_10398,N_8116,N_8266);
xor U10399 (N_10399,N_7838,N_8575);
and U10400 (N_10400,N_7665,N_8111);
nand U10401 (N_10401,N_8452,N_7813);
xor U10402 (N_10402,N_7690,N_8110);
and U10403 (N_10403,N_8426,N_7586);
and U10404 (N_10404,N_8221,N_8816);
and U10405 (N_10405,N_7995,N_8767);
nor U10406 (N_10406,N_8903,N_7887);
or U10407 (N_10407,N_7908,N_7975);
nand U10408 (N_10408,N_8466,N_8630);
nand U10409 (N_10409,N_8385,N_8312);
or U10410 (N_10410,N_8781,N_8511);
xnor U10411 (N_10411,N_8882,N_8283);
nand U10412 (N_10412,N_8142,N_8143);
and U10413 (N_10413,N_7523,N_8826);
and U10414 (N_10414,N_8829,N_8722);
xnor U10415 (N_10415,N_8337,N_7632);
nand U10416 (N_10416,N_8148,N_8086);
xnor U10417 (N_10417,N_8069,N_7585);
nand U10418 (N_10418,N_8371,N_8415);
nand U10419 (N_10419,N_8927,N_8946);
xor U10420 (N_10420,N_7731,N_8405);
nor U10421 (N_10421,N_8668,N_7623);
nor U10422 (N_10422,N_8241,N_8542);
nand U10423 (N_10423,N_7698,N_7941);
and U10424 (N_10424,N_8705,N_8670);
nor U10425 (N_10425,N_7749,N_7572);
and U10426 (N_10426,N_8212,N_8886);
and U10427 (N_10427,N_8383,N_8471);
or U10428 (N_10428,N_7773,N_8407);
or U10429 (N_10429,N_7727,N_8857);
nand U10430 (N_10430,N_8445,N_7580);
and U10431 (N_10431,N_7816,N_8542);
xor U10432 (N_10432,N_8428,N_7652);
or U10433 (N_10433,N_8808,N_8382);
or U10434 (N_10434,N_8918,N_8980);
xor U10435 (N_10435,N_8003,N_8440);
xor U10436 (N_10436,N_8814,N_7965);
nor U10437 (N_10437,N_7719,N_8103);
xnor U10438 (N_10438,N_8252,N_8522);
nand U10439 (N_10439,N_7844,N_8044);
nor U10440 (N_10440,N_8593,N_7646);
or U10441 (N_10441,N_7934,N_8809);
or U10442 (N_10442,N_7575,N_7632);
nor U10443 (N_10443,N_7966,N_8587);
xor U10444 (N_10444,N_8012,N_8296);
xor U10445 (N_10445,N_8095,N_8217);
nor U10446 (N_10446,N_8456,N_7952);
or U10447 (N_10447,N_8888,N_8965);
nand U10448 (N_10448,N_8197,N_8403);
or U10449 (N_10449,N_7703,N_7994);
xor U10450 (N_10450,N_8214,N_8453);
nor U10451 (N_10451,N_8353,N_8606);
and U10452 (N_10452,N_8957,N_8904);
nand U10453 (N_10453,N_7844,N_8277);
or U10454 (N_10454,N_8254,N_8715);
nor U10455 (N_10455,N_8890,N_7952);
and U10456 (N_10456,N_8209,N_8429);
nor U10457 (N_10457,N_8953,N_8155);
nand U10458 (N_10458,N_8040,N_8575);
xor U10459 (N_10459,N_8675,N_7797);
xor U10460 (N_10460,N_8001,N_7815);
and U10461 (N_10461,N_7793,N_8773);
nor U10462 (N_10462,N_7904,N_8173);
or U10463 (N_10463,N_8580,N_8003);
nand U10464 (N_10464,N_8438,N_8629);
or U10465 (N_10465,N_8084,N_8952);
and U10466 (N_10466,N_8261,N_8830);
nor U10467 (N_10467,N_8949,N_8573);
nand U10468 (N_10468,N_7765,N_8607);
xnor U10469 (N_10469,N_8683,N_8763);
and U10470 (N_10470,N_7762,N_8783);
or U10471 (N_10471,N_8462,N_8182);
and U10472 (N_10472,N_8044,N_8663);
and U10473 (N_10473,N_8782,N_7957);
or U10474 (N_10474,N_8002,N_8144);
or U10475 (N_10475,N_8079,N_7655);
and U10476 (N_10476,N_8893,N_8904);
nand U10477 (N_10477,N_8710,N_8285);
nor U10478 (N_10478,N_8236,N_8114);
and U10479 (N_10479,N_8247,N_7894);
nor U10480 (N_10480,N_8375,N_7982);
nand U10481 (N_10481,N_8404,N_8741);
or U10482 (N_10482,N_8203,N_8157);
xor U10483 (N_10483,N_8416,N_8780);
nor U10484 (N_10484,N_8811,N_8501);
and U10485 (N_10485,N_8607,N_7628);
nand U10486 (N_10486,N_7906,N_8475);
and U10487 (N_10487,N_7637,N_8349);
or U10488 (N_10488,N_8616,N_8675);
xor U10489 (N_10489,N_7562,N_8997);
nor U10490 (N_10490,N_8497,N_8892);
and U10491 (N_10491,N_7713,N_7518);
xor U10492 (N_10492,N_8559,N_7567);
nand U10493 (N_10493,N_8523,N_7753);
or U10494 (N_10494,N_8307,N_8536);
xnor U10495 (N_10495,N_7828,N_7819);
and U10496 (N_10496,N_7557,N_8346);
xnor U10497 (N_10497,N_8771,N_8054);
or U10498 (N_10498,N_8878,N_7767);
nand U10499 (N_10499,N_7786,N_7987);
nand U10500 (N_10500,N_10068,N_9798);
and U10501 (N_10501,N_9873,N_9556);
nor U10502 (N_10502,N_10376,N_9153);
nand U10503 (N_10503,N_10316,N_9668);
xor U10504 (N_10504,N_10370,N_9657);
and U10505 (N_10505,N_9550,N_9065);
nor U10506 (N_10506,N_9846,N_9324);
nor U10507 (N_10507,N_9654,N_10191);
and U10508 (N_10508,N_9316,N_10061);
nand U10509 (N_10509,N_9639,N_9537);
and U10510 (N_10510,N_9515,N_10317);
xnor U10511 (N_10511,N_9723,N_9385);
xnor U10512 (N_10512,N_9584,N_10287);
nor U10513 (N_10513,N_10037,N_9301);
and U10514 (N_10514,N_9880,N_10236);
or U10515 (N_10515,N_9501,N_9405);
or U10516 (N_10516,N_9703,N_9136);
nand U10517 (N_10517,N_9431,N_9403);
nand U10518 (N_10518,N_10426,N_9650);
and U10519 (N_10519,N_9706,N_9117);
nor U10520 (N_10520,N_9937,N_10147);
nor U10521 (N_10521,N_9666,N_9623);
and U10522 (N_10522,N_9057,N_9251);
xor U10523 (N_10523,N_9868,N_10223);
nor U10524 (N_10524,N_9946,N_10255);
nand U10525 (N_10525,N_9180,N_9157);
xnor U10526 (N_10526,N_10108,N_9128);
and U10527 (N_10527,N_9216,N_9156);
xnor U10528 (N_10528,N_9903,N_9532);
nand U10529 (N_10529,N_10380,N_9595);
and U10530 (N_10530,N_9634,N_9827);
nand U10531 (N_10531,N_9508,N_10084);
nor U10532 (N_10532,N_10286,N_9488);
nand U10533 (N_10533,N_10275,N_10135);
nor U10534 (N_10534,N_9226,N_9265);
and U10535 (N_10535,N_9466,N_10077);
xnor U10536 (N_10536,N_10285,N_9204);
or U10537 (N_10537,N_10356,N_9683);
and U10538 (N_10538,N_10076,N_9383);
nor U10539 (N_10539,N_9496,N_9600);
xor U10540 (N_10540,N_9871,N_9037);
or U10541 (N_10541,N_9625,N_9296);
nand U10542 (N_10542,N_9667,N_9140);
xor U10543 (N_10543,N_9949,N_9074);
xor U10544 (N_10544,N_9984,N_10014);
or U10545 (N_10545,N_9413,N_9356);
nor U10546 (N_10546,N_10273,N_10162);
and U10547 (N_10547,N_9304,N_9217);
or U10548 (N_10548,N_10470,N_9255);
and U10549 (N_10549,N_10253,N_10214);
nand U10550 (N_10550,N_9404,N_10419);
and U10551 (N_10551,N_10199,N_10182);
xor U10552 (N_10552,N_9738,N_10143);
xor U10553 (N_10553,N_10060,N_10302);
nor U10554 (N_10554,N_9622,N_9328);
and U10555 (N_10555,N_10119,N_10159);
and U10556 (N_10556,N_9451,N_10123);
and U10557 (N_10557,N_9010,N_9805);
or U10558 (N_10558,N_9977,N_9961);
nor U10559 (N_10559,N_10128,N_9271);
and U10560 (N_10560,N_9219,N_10374);
and U10561 (N_10561,N_9808,N_9305);
and U10562 (N_10562,N_10237,N_9778);
nor U10563 (N_10563,N_9620,N_9450);
and U10564 (N_10564,N_10212,N_9347);
and U10565 (N_10565,N_9360,N_10217);
or U10566 (N_10566,N_10100,N_9154);
and U10567 (N_10567,N_9765,N_10321);
or U10568 (N_10568,N_9237,N_10194);
nor U10569 (N_10569,N_9746,N_9744);
and U10570 (N_10570,N_10091,N_10291);
nor U10571 (N_10571,N_10283,N_9343);
nand U10572 (N_10572,N_10368,N_10114);
xnor U10573 (N_10573,N_9139,N_9097);
or U10574 (N_10574,N_9740,N_10111);
or U10575 (N_10575,N_9875,N_10067);
xnor U10576 (N_10576,N_9281,N_9710);
and U10577 (N_10577,N_9190,N_9215);
nor U10578 (N_10578,N_9321,N_10101);
or U10579 (N_10579,N_10028,N_9959);
nand U10580 (N_10580,N_9919,N_9366);
xor U10581 (N_10581,N_10475,N_10030);
and U10582 (N_10582,N_9252,N_9241);
or U10583 (N_10583,N_10274,N_9303);
and U10584 (N_10584,N_10152,N_9454);
nand U10585 (N_10585,N_9588,N_9837);
nand U10586 (N_10586,N_10297,N_9194);
xnor U10587 (N_10587,N_9349,N_10467);
nand U10588 (N_10588,N_9016,N_9292);
and U10589 (N_10589,N_9045,N_9986);
xnor U10590 (N_10590,N_9771,N_9815);
nor U10591 (N_10591,N_9464,N_9784);
or U10592 (N_10592,N_10427,N_9373);
or U10593 (N_10593,N_10282,N_10125);
xor U10594 (N_10594,N_9202,N_9574);
xnor U10595 (N_10595,N_10337,N_9598);
and U10596 (N_10596,N_9049,N_10340);
or U10597 (N_10597,N_9544,N_9963);
xnor U10598 (N_10598,N_9182,N_9663);
nand U10599 (N_10599,N_9952,N_9053);
nand U10600 (N_10600,N_10322,N_9175);
xnor U10601 (N_10601,N_9865,N_9842);
nand U10602 (N_10602,N_10139,N_9857);
xnor U10603 (N_10603,N_10130,N_10088);
nand U10604 (N_10604,N_9593,N_9422);
nor U10605 (N_10605,N_10145,N_10314);
nor U10606 (N_10606,N_9106,N_10423);
or U10607 (N_10607,N_9633,N_10203);
nor U10608 (N_10608,N_10023,N_9525);
xnor U10609 (N_10609,N_10010,N_9551);
or U10610 (N_10610,N_9341,N_10411);
xor U10611 (N_10611,N_9661,N_9186);
and U10612 (N_10612,N_9181,N_9036);
xnor U10613 (N_10613,N_9424,N_10184);
and U10614 (N_10614,N_9239,N_9981);
and U10615 (N_10615,N_9264,N_9462);
nand U10616 (N_10616,N_9856,N_9026);
or U10617 (N_10617,N_9232,N_9086);
and U10618 (N_10618,N_9656,N_9870);
or U10619 (N_10619,N_10174,N_9660);
nand U10620 (N_10620,N_9312,N_10464);
and U10621 (N_10621,N_9354,N_9928);
and U10622 (N_10622,N_9495,N_10220);
and U10623 (N_10623,N_9258,N_9726);
and U10624 (N_10624,N_10041,N_10228);
xnor U10625 (N_10625,N_9119,N_9849);
or U10626 (N_10626,N_10185,N_9018);
and U10627 (N_10627,N_10490,N_9695);
and U10628 (N_10628,N_9262,N_9612);
nand U10629 (N_10629,N_9665,N_10264);
xnor U10630 (N_10630,N_10434,N_9229);
and U10631 (N_10631,N_10346,N_10124);
or U10632 (N_10632,N_9836,N_10158);
xnor U10633 (N_10633,N_9320,N_9131);
xnor U10634 (N_10634,N_9279,N_9528);
nor U10635 (N_10635,N_10105,N_9460);
and U10636 (N_10636,N_10201,N_9013);
or U10637 (N_10637,N_9887,N_9969);
nor U10638 (N_10638,N_9783,N_10004);
or U10639 (N_10639,N_9915,N_10318);
nand U10640 (N_10640,N_9171,N_10462);
nand U10641 (N_10641,N_10449,N_9114);
and U10642 (N_10642,N_9280,N_9192);
xor U10643 (N_10643,N_9021,N_10446);
nor U10644 (N_10644,N_9944,N_10357);
xor U10645 (N_10645,N_10213,N_9769);
or U10646 (N_10646,N_9902,N_9147);
or U10647 (N_10647,N_9160,N_9134);
xor U10648 (N_10648,N_9306,N_10062);
and U10649 (N_10649,N_9375,N_10326);
nor U10650 (N_10650,N_10360,N_10024);
and U10651 (N_10651,N_9244,N_9372);
xor U10652 (N_10652,N_9091,N_10366);
xor U10653 (N_10653,N_10053,N_9084);
or U10654 (N_10654,N_9813,N_9407);
nand U10655 (N_10655,N_9945,N_10293);
or U10656 (N_10656,N_9749,N_9956);
nor U10657 (N_10657,N_10226,N_10261);
nor U10658 (N_10658,N_10052,N_9035);
nand U10659 (N_10659,N_10136,N_9874);
and U10660 (N_10660,N_9882,N_9076);
nand U10661 (N_10661,N_9910,N_9253);
xnor U10662 (N_10662,N_9811,N_9402);
nor U10663 (N_10663,N_9398,N_9075);
or U10664 (N_10664,N_10042,N_10328);
and U10665 (N_10665,N_9061,N_9393);
nor U10666 (N_10666,N_9092,N_10015);
nand U10667 (N_10667,N_9031,N_9884);
and U10668 (N_10668,N_9812,N_9287);
nor U10669 (N_10669,N_9472,N_9187);
or U10670 (N_10670,N_9497,N_9731);
and U10671 (N_10671,N_9334,N_9697);
or U10672 (N_10672,N_9499,N_9770);
or U10673 (N_10673,N_9705,N_9209);
and U10674 (N_10674,N_9379,N_9476);
nand U10675 (N_10675,N_9965,N_10421);
and U10676 (N_10676,N_10477,N_9776);
and U10677 (N_10677,N_9392,N_9012);
xnor U10678 (N_10678,N_9170,N_9901);
nor U10679 (N_10679,N_10187,N_10150);
nor U10680 (N_10680,N_9767,N_10412);
or U10681 (N_10681,N_10339,N_10485);
xor U10682 (N_10682,N_9917,N_9469);
nand U10683 (N_10683,N_9823,N_9121);
and U10684 (N_10684,N_10252,N_9979);
nand U10685 (N_10685,N_10190,N_9432);
and U10686 (N_10686,N_10402,N_10106);
and U10687 (N_10687,N_10035,N_10375);
xnor U10688 (N_10688,N_9526,N_9921);
nor U10689 (N_10689,N_10054,N_10081);
or U10690 (N_10690,N_9573,N_9135);
xor U10691 (N_10691,N_9889,N_9032);
and U10692 (N_10692,N_9835,N_10065);
and U10693 (N_10693,N_10040,N_9067);
nand U10694 (N_10694,N_9250,N_10395);
nor U10695 (N_10695,N_9803,N_10183);
and U10696 (N_10696,N_9617,N_10401);
nor U10697 (N_10697,N_10113,N_10151);
nor U10698 (N_10698,N_9548,N_10071);
or U10699 (N_10699,N_9090,N_9955);
nor U10700 (N_10700,N_9742,N_10117);
xor U10701 (N_10701,N_10079,N_10029);
xnor U10702 (N_10702,N_10096,N_10300);
or U10703 (N_10703,N_9947,N_10486);
or U10704 (N_10704,N_9231,N_10243);
nor U10705 (N_10705,N_9631,N_10144);
nand U10706 (N_10706,N_10355,N_10176);
and U10707 (N_10707,N_10116,N_10109);
or U10708 (N_10708,N_9756,N_10180);
nand U10709 (N_10709,N_9640,N_9096);
nand U10710 (N_10710,N_10371,N_10221);
or U10711 (N_10711,N_9143,N_9381);
nand U10712 (N_10712,N_9781,N_9580);
nand U10713 (N_10713,N_10444,N_9315);
xnor U10714 (N_10714,N_9234,N_10379);
nand U10715 (N_10715,N_10189,N_9310);
xnor U10716 (N_10716,N_9970,N_10383);
xor U10717 (N_10717,N_9042,N_9210);
nand U10718 (N_10718,N_10348,N_9411);
or U10719 (N_10719,N_9483,N_9758);
nor U10720 (N_10720,N_9072,N_9369);
nor U10721 (N_10721,N_9093,N_10160);
and U10722 (N_10722,N_9809,N_9897);
and U10723 (N_10723,N_10384,N_10127);
xor U10724 (N_10724,N_9927,N_9712);
nor U10725 (N_10725,N_10095,N_9885);
nor U10726 (N_10726,N_9879,N_9430);
and U10727 (N_10727,N_9943,N_9958);
xor U10728 (N_10728,N_10456,N_9440);
and U10729 (N_10729,N_9862,N_10409);
nand U10730 (N_10730,N_10057,N_10197);
xor U10731 (N_10731,N_9282,N_9579);
nor U10732 (N_10732,N_10126,N_9230);
or U10733 (N_10733,N_9174,N_9912);
xnor U10734 (N_10734,N_10051,N_9124);
and U10735 (N_10735,N_9954,N_10206);
and U10736 (N_10736,N_10262,N_10138);
and U10737 (N_10737,N_9218,N_9883);
and U10738 (N_10738,N_10205,N_10025);
nand U10739 (N_10739,N_9060,N_9427);
or U10740 (N_10740,N_9213,N_10089);
nand U10741 (N_10741,N_10155,N_9750);
xor U10742 (N_10742,N_10045,N_9044);
nand U10743 (N_10743,N_9277,N_10393);
nor U10744 (N_10744,N_10167,N_9960);
nand U10745 (N_10745,N_10069,N_9980);
xor U10746 (N_10746,N_9384,N_9452);
xor U10747 (N_10747,N_9289,N_9892);
nand U10748 (N_10748,N_9833,N_9167);
nand U10749 (N_10749,N_9487,N_9975);
nand U10750 (N_10750,N_9391,N_10372);
xor U10751 (N_10751,N_9618,N_9342);
xor U10752 (N_10752,N_9177,N_9468);
and U10753 (N_10753,N_9322,N_9481);
xor U10754 (N_10754,N_9913,N_9535);
nor U10755 (N_10755,N_9141,N_9085);
nor U10756 (N_10756,N_9717,N_10031);
or U10757 (N_10757,N_9957,N_9329);
nor U10758 (N_10758,N_10198,N_9396);
xor U10759 (N_10759,N_9212,N_9939);
nor U10760 (N_10760,N_9056,N_10195);
nand U10761 (N_10761,N_10229,N_9794);
xnor U10762 (N_10762,N_9534,N_9138);
nor U10763 (N_10763,N_9736,N_10087);
xor U10764 (N_10764,N_9626,N_9721);
nand U10765 (N_10765,N_9102,N_9199);
nand U10766 (N_10766,N_9520,N_9118);
nand U10767 (N_10767,N_10440,N_9364);
xor U10768 (N_10768,N_9557,N_9936);
nand U10769 (N_10769,N_9014,N_9570);
nand U10770 (N_10770,N_9380,N_9779);
nor U10771 (N_10771,N_10272,N_9048);
nor U10772 (N_10772,N_10487,N_9168);
nand U10773 (N_10773,N_9333,N_10492);
nor U10774 (N_10774,N_9704,N_10331);
nor U10775 (N_10775,N_9877,N_9637);
or U10776 (N_10776,N_9005,N_9493);
and U10777 (N_10777,N_9261,N_9554);
xor U10778 (N_10778,N_9467,N_10344);
nand U10779 (N_10779,N_9890,N_10333);
or U10780 (N_10780,N_9169,N_9071);
or U10781 (N_10781,N_9011,N_9519);
or U10782 (N_10782,N_9340,N_9604);
or U10783 (N_10783,N_9966,N_9299);
xnor U10784 (N_10784,N_10334,N_10323);
xnor U10785 (N_10785,N_9094,N_9995);
nor U10786 (N_10786,N_9638,N_10244);
and U10787 (N_10787,N_9068,N_10034);
nor U10788 (N_10788,N_10361,N_10407);
or U10789 (N_10789,N_9516,N_9636);
and U10790 (N_10790,N_10265,N_9500);
nand U10791 (N_10791,N_9715,N_9517);
xnor U10792 (N_10792,N_10394,N_10161);
nor U10793 (N_10793,N_9144,N_10473);
nor U10794 (N_10794,N_9616,N_9964);
and U10795 (N_10795,N_9188,N_9103);
and U10796 (N_10796,N_9807,N_9577);
or U10797 (N_10797,N_9429,N_10258);
nor U10798 (N_10798,N_9308,N_9669);
or U10799 (N_10799,N_10168,N_9564);
xnor U10800 (N_10800,N_9020,N_9410);
nor U10801 (N_10801,N_10238,N_9678);
or U10802 (N_10802,N_10442,N_9270);
nand U10803 (N_10803,N_10141,N_9034);
nand U10804 (N_10804,N_9567,N_10211);
and U10805 (N_10805,N_10064,N_10164);
nor U10806 (N_10806,N_9694,N_9614);
xnor U10807 (N_10807,N_9368,N_9569);
xnor U10808 (N_10808,N_9069,N_9689);
xnor U10809 (N_10809,N_9681,N_10173);
and U10810 (N_10810,N_10294,N_9498);
or U10811 (N_10811,N_9932,N_9482);
nor U10812 (N_10812,N_10315,N_10112);
nand U10813 (N_10813,N_10204,N_9473);
or U10814 (N_10814,N_9233,N_9129);
and U10815 (N_10815,N_9365,N_9571);
xnor U10816 (N_10816,N_9540,N_9938);
and U10817 (N_10817,N_10157,N_10165);
xnor U10818 (N_10818,N_10169,N_9109);
xnor U10819 (N_10819,N_9001,N_9825);
nand U10820 (N_10820,N_9235,N_10471);
nor U10821 (N_10821,N_10432,N_9853);
or U10822 (N_10822,N_9733,N_9796);
or U10823 (N_10823,N_10260,N_9415);
xor U10824 (N_10824,N_9337,N_10072);
nand U10825 (N_10825,N_9855,N_9759);
or U10826 (N_10826,N_9552,N_9772);
and U10827 (N_10827,N_9539,N_10278);
nor U10828 (N_10828,N_9492,N_10098);
nand U10829 (N_10829,N_10306,N_10484);
nor U10830 (N_10830,N_9562,N_10248);
nand U10831 (N_10831,N_9200,N_10429);
xor U10832 (N_10832,N_9635,N_10082);
xor U10833 (N_10833,N_10312,N_10202);
xor U10834 (N_10834,N_9486,N_9110);
or U10835 (N_10835,N_9459,N_10468);
xor U10836 (N_10836,N_9941,N_9457);
or U10837 (N_10837,N_9576,N_9257);
or U10838 (N_10838,N_10320,N_9309);
or U10839 (N_10839,N_10092,N_10269);
nor U10840 (N_10840,N_9568,N_9824);
nand U10841 (N_10841,N_9732,N_9127);
and U10842 (N_10842,N_9437,N_9418);
nand U10843 (N_10843,N_9693,N_9133);
nor U10844 (N_10844,N_9659,N_9791);
nor U10845 (N_10845,N_9330,N_10452);
or U10846 (N_10846,N_9080,N_9256);
nand U10847 (N_10847,N_9353,N_9420);
nor U10848 (N_10848,N_10296,N_9630);
nand U10849 (N_10849,N_9345,N_9926);
and U10850 (N_10850,N_9185,N_10377);
nor U10851 (N_10851,N_9030,N_9839);
and U10852 (N_10852,N_10016,N_10418);
nor U10853 (N_10853,N_9435,N_9007);
or U10854 (N_10854,N_9191,N_9445);
xnor U10855 (N_10855,N_10120,N_9920);
nor U10856 (N_10856,N_10043,N_10002);
nand U10857 (N_10857,N_9652,N_9298);
xnor U10858 (N_10858,N_9649,N_9672);
nor U10859 (N_10859,N_10324,N_9613);
xor U10860 (N_10860,N_9931,N_9505);
nand U10861 (N_10861,N_10122,N_9083);
xor U10862 (N_10862,N_9530,N_9647);
and U10863 (N_10863,N_10078,N_9948);
and U10864 (N_10864,N_9696,N_10048);
nand U10865 (N_10865,N_9872,N_9115);
or U10866 (N_10866,N_9722,N_9173);
nand U10867 (N_10867,N_9867,N_9426);
xor U10868 (N_10868,N_9850,N_10259);
or U10869 (N_10869,N_9602,N_9909);
nor U10870 (N_10870,N_9019,N_9490);
xor U10871 (N_10871,N_10365,N_9719);
xnor U10872 (N_10872,N_10066,N_9120);
nand U10873 (N_10873,N_9852,N_9455);
nand U10874 (N_10874,N_9822,N_9692);
nor U10875 (N_10875,N_9940,N_9549);
nor U10876 (N_10876,N_10140,N_9240);
nand U10877 (N_10877,N_9739,N_9997);
xnor U10878 (N_10878,N_10461,N_9972);
and U10879 (N_10879,N_9848,N_9967);
or U10880 (N_10880,N_10424,N_9448);
nor U10881 (N_10881,N_10307,N_9082);
nor U10882 (N_10882,N_10225,N_9918);
xnor U10883 (N_10883,N_10235,N_9336);
and U10884 (N_10884,N_9601,N_9155);
nor U10885 (N_10885,N_9433,N_10389);
nor U10886 (N_10886,N_9023,N_9728);
xor U10887 (N_10887,N_10329,N_10270);
nor U10888 (N_10888,N_9687,N_10441);
xor U10889 (N_10889,N_9542,N_9914);
nor U10890 (N_10890,N_9698,N_9254);
and U10891 (N_10891,N_10428,N_9859);
or U10892 (N_10892,N_9793,N_9243);
nand U10893 (N_10893,N_10257,N_10335);
nor U10894 (N_10894,N_10055,N_10404);
or U10895 (N_10895,N_10142,N_9294);
nor U10896 (N_10896,N_10149,N_10347);
and U10897 (N_10897,N_9161,N_9362);
nand U10898 (N_10898,N_9610,N_10290);
or U10899 (N_10899,N_10247,N_10364);
nor U10900 (N_10900,N_9286,N_10304);
nor U10901 (N_10901,N_10063,N_10494);
nand U10902 (N_10902,N_10436,N_9751);
nand U10903 (N_10903,N_9307,N_9589);
xor U10904 (N_10904,N_10398,N_10415);
nand U10905 (N_10905,N_10222,N_9348);
or U10906 (N_10906,N_10354,N_10121);
or U10907 (N_10907,N_9220,N_10070);
and U10908 (N_10908,N_10110,N_9607);
or U10909 (N_10909,N_9363,N_10209);
xor U10910 (N_10910,N_9806,N_10420);
or U10911 (N_10911,N_9866,N_10489);
nand U10912 (N_10912,N_9295,N_9198);
or U10913 (N_10913,N_9123,N_9810);
or U10914 (N_10914,N_9406,N_9148);
nor U10915 (N_10915,N_9831,N_10455);
nor U10916 (N_10916,N_9050,N_10496);
xnor U10917 (N_10917,N_9400,N_10133);
and U10918 (N_10918,N_10026,N_10457);
nand U10919 (N_10919,N_9325,N_9709);
nand U10920 (N_10920,N_9895,N_10478);
and U10921 (N_10921,N_9560,N_9502);
and U10922 (N_10922,N_9269,N_10430);
nand U10923 (N_10923,N_9592,N_9300);
nand U10924 (N_10924,N_9088,N_9971);
and U10925 (N_10925,N_9205,N_9522);
and U10926 (N_10926,N_9339,N_9527);
xor U10927 (N_10927,N_9260,N_10414);
nor U10928 (N_10928,N_9477,N_9463);
nand U10929 (N_10929,N_10388,N_10367);
nor U10930 (N_10930,N_9283,N_9078);
nand U10931 (N_10931,N_9099,N_9988);
xor U10932 (N_10932,N_10097,N_9101);
nand U10933 (N_10933,N_9272,N_9566);
xor U10934 (N_10934,N_9290,N_9925);
nor U10935 (N_10935,N_9775,N_10207);
nor U10936 (N_10936,N_10232,N_9438);
and U10937 (N_10937,N_10482,N_9046);
nor U10938 (N_10938,N_9670,N_9236);
and U10939 (N_10939,N_10341,N_9189);
xnor U10940 (N_10940,N_9025,N_9878);
nor U10941 (N_10941,N_9478,N_9624);
nor U10942 (N_10942,N_10309,N_9399);
xnor U10943 (N_10943,N_9052,N_9331);
and U10944 (N_10944,N_10179,N_9844);
and U10945 (N_10945,N_10186,N_9905);
nor U10946 (N_10946,N_9471,N_10327);
and U10947 (N_10947,N_9314,N_10483);
or U10948 (N_10948,N_10305,N_9323);
xor U10949 (N_10949,N_10338,N_9165);
xor U10950 (N_10950,N_9183,N_9070);
nand U10951 (N_10951,N_10463,N_9382);
xnor U10952 (N_10952,N_9291,N_9730);
or U10953 (N_10953,N_9374,N_10387);
nand U10954 (N_10954,N_9802,N_9105);
and U10955 (N_10955,N_9465,N_10210);
xor U10956 (N_10956,N_9644,N_9397);
or U10957 (N_10957,N_9058,N_9685);
and U10958 (N_10958,N_10094,N_9263);
nand U10959 (N_10959,N_10153,N_9196);
or U10960 (N_10960,N_9475,N_10378);
and U10961 (N_10961,N_9801,N_9524);
and U10962 (N_10962,N_9355,N_10242);
nand U10963 (N_10963,N_9686,N_10188);
nor U10964 (N_10964,N_9900,N_10299);
or U10965 (N_10965,N_9081,N_10200);
xnor U10966 (N_10966,N_9511,N_10170);
nor U10967 (N_10967,N_9000,N_9387);
nor U10968 (N_10968,N_9389,N_9934);
xor U10969 (N_10969,N_9484,N_10454);
nand U10970 (N_10970,N_9273,N_10218);
or U10971 (N_10971,N_10403,N_9159);
nor U10972 (N_10972,N_10268,N_9763);
nor U10973 (N_10973,N_9512,N_10074);
nor U10974 (N_10974,N_9461,N_9267);
and U10975 (N_10975,N_10480,N_9605);
xor U10976 (N_10976,N_10018,N_9821);
nor U10977 (N_10977,N_9725,N_9377);
nand U10978 (N_10978,N_9747,N_9278);
and U10979 (N_10979,N_9766,N_9676);
and U10980 (N_10980,N_9409,N_9641);
nor U10981 (N_10981,N_9223,N_9158);
and U10982 (N_10982,N_9628,N_9752);
and U10983 (N_10983,N_9022,N_9024);
nor U10984 (N_10984,N_9591,N_9788);
and U10985 (N_10985,N_9782,N_10271);
and U10986 (N_10986,N_9619,N_10005);
or U10987 (N_10987,N_9054,N_9350);
or U10988 (N_10988,N_9107,N_9439);
or U10989 (N_10989,N_9819,N_9606);
nor U10990 (N_10990,N_9436,N_9891);
or U10991 (N_10991,N_9442,N_10192);
and U10992 (N_10992,N_10391,N_9108);
nor U10993 (N_10993,N_9679,N_9015);
xor U10994 (N_10994,N_10311,N_9428);
or U10995 (N_10995,N_9906,N_9100);
nor U10996 (N_10996,N_9843,N_9063);
and U10997 (N_10997,N_9713,N_9646);
or U10998 (N_10998,N_9820,N_9829);
nand U10999 (N_10999,N_9126,N_10358);
and U11000 (N_11000,N_10090,N_9122);
nor U11001 (N_11001,N_10433,N_9449);
or U11002 (N_11002,N_10003,N_10488);
nand U11003 (N_11003,N_9043,N_9597);
and U11004 (N_11004,N_9583,N_9506);
nand U11005 (N_11005,N_9653,N_9688);
nor U11006 (N_11006,N_10313,N_10154);
or U11007 (N_11007,N_9737,N_9533);
nor U11008 (N_11008,N_10437,N_9987);
nor U11009 (N_11009,N_10396,N_9179);
and U11010 (N_11010,N_10413,N_10336);
or U11011 (N_11011,N_9266,N_9164);
or U11012 (N_11012,N_9590,N_9951);
or U11013 (N_11013,N_9543,N_9311);
nand U11014 (N_11014,N_9335,N_10239);
nor U11015 (N_11015,N_10406,N_9359);
and U11016 (N_11016,N_9792,N_10448);
xnor U11017 (N_11017,N_9861,N_9609);
nor U11018 (N_11018,N_10493,N_9994);
nor U11019 (N_11019,N_9645,N_9923);
nand U11020 (N_11020,N_9033,N_10319);
xor U11021 (N_11021,N_10075,N_10039);
and U11022 (N_11022,N_10330,N_10129);
and U11023 (N_11023,N_10298,N_9546);
xor U11024 (N_11024,N_9149,N_9673);
nor U11025 (N_11025,N_10224,N_9968);
nand U11026 (N_11026,N_9474,N_10103);
xnor U11027 (N_11027,N_10006,N_10156);
nand U11028 (N_11028,N_9864,N_10416);
or U11029 (N_11029,N_9774,N_10310);
xor U11030 (N_11030,N_10178,N_9565);
nand U11031 (N_11031,N_10137,N_9834);
and U11032 (N_11032,N_10342,N_9586);
and U11033 (N_11033,N_9990,N_9150);
nand U11034 (N_11034,N_9648,N_9748);
nor U11035 (N_11035,N_10499,N_9064);
or U11036 (N_11036,N_9699,N_9051);
and U11037 (N_11037,N_9434,N_9351);
xnor U11038 (N_11038,N_9494,N_9547);
nand U11039 (N_11039,N_9581,N_9112);
and U11040 (N_11040,N_9203,N_10284);
nor U11041 (N_11041,N_9211,N_9006);
or U11042 (N_11042,N_9992,N_9225);
or U11043 (N_11043,N_10451,N_10058);
or U11044 (N_11044,N_10086,N_9089);
and U11045 (N_11045,N_9425,N_10102);
xnor U11046 (N_11046,N_9621,N_9248);
nand U11047 (N_11047,N_9735,N_9394);
nor U11048 (N_11048,N_10425,N_9675);
nor U11049 (N_11049,N_9041,N_10465);
or U11050 (N_11050,N_9453,N_10175);
nand U11051 (N_11051,N_10280,N_9346);
nor U11052 (N_11052,N_9146,N_9275);
and U11053 (N_11053,N_9587,N_9017);
xnor U11054 (N_11054,N_9814,N_9184);
nand U11055 (N_11055,N_9274,N_10399);
and U11056 (N_11056,N_9376,N_9858);
xor U11057 (N_11057,N_10115,N_9197);
nor U11058 (N_11058,N_10256,N_10009);
or U11059 (N_11059,N_9896,N_9854);
or U11060 (N_11060,N_10104,N_9677);
or U11061 (N_11061,N_10472,N_9242);
and U11062 (N_11062,N_9922,N_10001);
nor U11063 (N_11063,N_9662,N_9991);
and U11064 (N_11064,N_9222,N_10474);
nand U11065 (N_11065,N_9458,N_9982);
xor U11066 (N_11066,N_9104,N_9840);
or U11067 (N_11067,N_9816,N_9830);
or U11068 (N_11068,N_9757,N_9038);
nor U11069 (N_11069,N_10231,N_10215);
and U11070 (N_11070,N_10343,N_9326);
xor U11071 (N_11071,N_9847,N_10359);
or U11072 (N_11072,N_9441,N_9536);
or U11073 (N_11073,N_9790,N_9111);
nor U11074 (N_11074,N_9838,N_9930);
xnor U11075 (N_11075,N_9302,N_9327);
and U11076 (N_11076,N_9443,N_10012);
xor U11077 (N_11077,N_9996,N_9352);
nor U11078 (N_11078,N_10007,N_10352);
nand U11079 (N_11079,N_9414,N_9828);
nand U11080 (N_11080,N_10438,N_10292);
or U11081 (N_11081,N_9582,N_10193);
xor U11082 (N_11082,N_9538,N_9974);
xnor U11083 (N_11083,N_9313,N_9888);
nor U11084 (N_11084,N_9743,N_9004);
nand U11085 (N_11085,N_9386,N_10353);
and U11086 (N_11086,N_9983,N_9594);
nand U11087 (N_11087,N_10046,N_10373);
xnor U11088 (N_11088,N_10107,N_9087);
nor U11089 (N_11089,N_9332,N_9077);
or U11090 (N_11090,N_9800,N_10118);
nor U11091 (N_11091,N_10431,N_9561);
xor U11092 (N_11092,N_9768,N_9412);
and U11093 (N_11093,N_9716,N_10369);
xnor U11094 (N_11094,N_10350,N_9247);
and U11095 (N_11095,N_9059,N_9416);
or U11096 (N_11096,N_10234,N_9116);
nand U11097 (N_11097,N_10022,N_9444);
xnor U11098 (N_11098,N_9447,N_9764);
or U11099 (N_11099,N_10230,N_10219);
xnor U11100 (N_11100,N_9417,N_9761);
and U11101 (N_11101,N_9978,N_9221);
and U11102 (N_11102,N_9818,N_9259);
and U11103 (N_11103,N_10332,N_10080);
nand U11104 (N_11104,N_9344,N_9367);
nor U11105 (N_11105,N_9338,N_9615);
or U11106 (N_11106,N_9249,N_9762);
nand U11107 (N_11107,N_9572,N_9976);
nor U11108 (N_11108,N_9207,N_9456);
nand U11109 (N_11109,N_9370,N_9817);
xor U11110 (N_11110,N_9632,N_9028);
and U11111 (N_11111,N_9777,N_10196);
nor U11112 (N_11112,N_10134,N_9664);
and U11113 (N_11113,N_10417,N_9655);
or U11114 (N_11114,N_9073,N_9388);
nor U11115 (N_11115,N_9113,N_9419);
and U11116 (N_11116,N_10093,N_9390);
nor U11117 (N_11117,N_9787,N_10013);
or U11118 (N_11118,N_9132,N_10277);
xnor U11119 (N_11119,N_10439,N_10363);
nor U11120 (N_11120,N_9507,N_9040);
xnor U11121 (N_11121,N_9700,N_10146);
and U11122 (N_11122,N_9993,N_9690);
or U11123 (N_11123,N_10245,N_10249);
nand U11124 (N_11124,N_10445,N_9529);
nand U11125 (N_11125,N_9989,N_9489);
nor U11126 (N_11126,N_9479,N_9718);
xnor U11127 (N_11127,N_9371,N_10251);
nand U11128 (N_11128,N_9734,N_9729);
and U11129 (N_11129,N_10021,N_9708);
xnor U11130 (N_11130,N_9780,N_9575);
nor U11131 (N_11131,N_10288,N_9985);
and U11132 (N_11132,N_10033,N_9795);
nand U11133 (N_11133,N_9470,N_9916);
xor U11134 (N_11134,N_9904,N_10227);
or U11135 (N_11135,N_9898,N_10410);
nor U11136 (N_11136,N_9029,N_10386);
xor U11137 (N_11137,N_9785,N_9682);
or U11138 (N_11138,N_10241,N_10056);
nor U11139 (N_11139,N_10020,N_9886);
xor U11140 (N_11140,N_10466,N_10351);
or U11141 (N_11141,N_9238,N_10163);
or U11142 (N_11142,N_9066,N_9055);
or U11143 (N_11143,N_9585,N_9559);
or U11144 (N_11144,N_9518,N_9714);
or U11145 (N_11145,N_9707,N_10397);
nand U11146 (N_11146,N_10345,N_9753);
and U11147 (N_11147,N_9727,N_9876);
nor U11148 (N_11148,N_9227,N_9629);
nor U11149 (N_11149,N_9268,N_9541);
and U11150 (N_11150,N_10038,N_10405);
nor U11151 (N_11151,N_9671,N_10132);
xor U11152 (N_11152,N_9881,N_9642);
nand U11153 (N_11153,N_10263,N_10019);
nand U11154 (N_11154,N_10008,N_9095);
xnor U11155 (N_11155,N_10308,N_9702);
nor U11156 (N_11156,N_9851,N_9224);
nor U11157 (N_11157,N_10295,N_9962);
and U11158 (N_11158,N_9523,N_10099);
xnor U11159 (N_11159,N_9401,N_10250);
or U11160 (N_11160,N_9950,N_9172);
or U11161 (N_11161,N_9924,N_9786);
and U11162 (N_11162,N_10131,N_9293);
nand U11163 (N_11163,N_10276,N_10497);
and U11164 (N_11164,N_9627,N_9893);
nor U11165 (N_11165,N_9485,N_9908);
nor U11166 (N_11166,N_9658,N_10050);
and U11167 (N_11167,N_9423,N_10000);
nor U11168 (N_11168,N_10177,N_9701);
xnor U11169 (N_11169,N_9228,N_10083);
and U11170 (N_11170,N_9285,N_10458);
and U11171 (N_11171,N_10400,N_9142);
or U11172 (N_11172,N_10381,N_9684);
nor U11173 (N_11173,N_9599,N_9008);
xnor U11174 (N_11174,N_9491,N_10047);
and U11175 (N_11175,N_10281,N_9039);
nand U11176 (N_11176,N_10011,N_9002);
nor U11177 (N_11177,N_10362,N_9510);
or U11178 (N_11178,N_10246,N_9563);
nor U11179 (N_11179,N_9276,N_9894);
xnor U11180 (N_11180,N_9062,N_10148);
or U11181 (N_11181,N_9166,N_9973);
xor U11182 (N_11182,N_9395,N_10233);
and U11183 (N_11183,N_10303,N_10479);
nor U11184 (N_11184,N_9755,N_10032);
nand U11185 (N_11185,N_10459,N_10481);
xor U11186 (N_11186,N_10469,N_9999);
or U11187 (N_11187,N_9832,N_10349);
xnor U11188 (N_11188,N_9578,N_9521);
or U11189 (N_11189,N_9804,N_10325);
nand U11190 (N_11190,N_9361,N_9152);
or U11191 (N_11191,N_9317,N_9079);
xor U11192 (N_11192,N_9509,N_10443);
nor U11193 (N_11193,N_10085,N_9773);
or U11194 (N_11194,N_10476,N_9288);
nand U11195 (N_11195,N_10453,N_10460);
nor U11196 (N_11196,N_10017,N_9193);
xnor U11197 (N_11197,N_10172,N_9942);
xor U11198 (N_11198,N_10216,N_9214);
xor U11199 (N_11199,N_9125,N_9378);
and U11200 (N_11200,N_10240,N_9680);
or U11201 (N_11201,N_9319,N_9480);
nor U11202 (N_11202,N_10266,N_9643);
or U11203 (N_11203,N_9799,N_9137);
xnor U11204 (N_11204,N_9408,N_9284);
or U11205 (N_11205,N_9929,N_9503);
nand U11206 (N_11206,N_9130,N_9953);
xnor U11207 (N_11207,N_9608,N_10392);
nand U11208 (N_11208,N_9720,N_9651);
and U11209 (N_11209,N_9206,N_9009);
xnor U11210 (N_11210,N_9674,N_10073);
xor U11211 (N_11211,N_9933,N_9826);
nand U11212 (N_11212,N_9098,N_9297);
nor U11213 (N_11213,N_10027,N_9178);
or U11214 (N_11214,N_10181,N_9145);
xnor U11215 (N_11215,N_9754,N_10408);
xor U11216 (N_11216,N_10208,N_9797);
nor U11217 (N_11217,N_10447,N_9558);
xor U11218 (N_11218,N_9907,N_9553);
xor U11219 (N_11219,N_10044,N_10390);
or U11220 (N_11220,N_9208,N_10301);
xor U11221 (N_11221,N_9195,N_9899);
nor U11222 (N_11222,N_9504,N_9531);
xor U11223 (N_11223,N_9935,N_10171);
nand U11224 (N_11224,N_9514,N_9745);
nand U11225 (N_11225,N_9162,N_9446);
or U11226 (N_11226,N_10049,N_9151);
nor U11227 (N_11227,N_10450,N_9869);
nand U11228 (N_11228,N_10254,N_9911);
xnor U11229 (N_11229,N_10435,N_9027);
and U11230 (N_11230,N_9358,N_9789);
xnor U11231 (N_11231,N_9860,N_10166);
xor U11232 (N_11232,N_9596,N_9760);
nor U11233 (N_11233,N_9555,N_9513);
or U11234 (N_11234,N_9711,N_9421);
xnor U11235 (N_11235,N_9724,N_9545);
xnor U11236 (N_11236,N_9603,N_9863);
or U11237 (N_11237,N_9318,N_10059);
and U11238 (N_11238,N_10422,N_10385);
nand U11239 (N_11239,N_9246,N_10289);
xnor U11240 (N_11240,N_9691,N_10382);
or U11241 (N_11241,N_9047,N_10495);
xor U11242 (N_11242,N_10279,N_9357);
xor U11243 (N_11243,N_9201,N_9611);
and U11244 (N_11244,N_9176,N_9741);
and U11245 (N_11245,N_9998,N_9163);
xnor U11246 (N_11246,N_10036,N_10491);
and U11247 (N_11247,N_9245,N_9845);
nand U11248 (N_11248,N_9841,N_9003);
or U11249 (N_11249,N_10267,N_10498);
or U11250 (N_11250,N_9086,N_10342);
nand U11251 (N_11251,N_9231,N_9959);
or U11252 (N_11252,N_10131,N_9839);
or U11253 (N_11253,N_9723,N_9507);
and U11254 (N_11254,N_9879,N_9196);
nand U11255 (N_11255,N_10313,N_10051);
and U11256 (N_11256,N_9117,N_9523);
or U11257 (N_11257,N_9559,N_9831);
xor U11258 (N_11258,N_10432,N_9201);
and U11259 (N_11259,N_10231,N_9060);
nand U11260 (N_11260,N_10098,N_9831);
xor U11261 (N_11261,N_9082,N_10257);
nor U11262 (N_11262,N_9116,N_10188);
and U11263 (N_11263,N_9812,N_10161);
nor U11264 (N_11264,N_10064,N_9009);
or U11265 (N_11265,N_9137,N_10207);
nor U11266 (N_11266,N_10338,N_10046);
nor U11267 (N_11267,N_9265,N_9379);
or U11268 (N_11268,N_9750,N_9041);
xnor U11269 (N_11269,N_9102,N_10327);
nand U11270 (N_11270,N_9607,N_9382);
and U11271 (N_11271,N_9465,N_9596);
nand U11272 (N_11272,N_9675,N_9826);
xnor U11273 (N_11273,N_9483,N_10220);
nand U11274 (N_11274,N_9106,N_9180);
or U11275 (N_11275,N_10135,N_9004);
and U11276 (N_11276,N_9901,N_9371);
nand U11277 (N_11277,N_9948,N_10495);
or U11278 (N_11278,N_10104,N_9880);
xor U11279 (N_11279,N_9444,N_10381);
xnor U11280 (N_11280,N_10455,N_9827);
xor U11281 (N_11281,N_10324,N_9422);
and U11282 (N_11282,N_9989,N_10410);
nor U11283 (N_11283,N_9677,N_9902);
or U11284 (N_11284,N_10143,N_9595);
and U11285 (N_11285,N_9247,N_9419);
nand U11286 (N_11286,N_10121,N_9072);
nand U11287 (N_11287,N_9978,N_10136);
nand U11288 (N_11288,N_10100,N_9978);
nand U11289 (N_11289,N_9538,N_9246);
or U11290 (N_11290,N_9067,N_10374);
nor U11291 (N_11291,N_9044,N_9720);
and U11292 (N_11292,N_9151,N_9913);
or U11293 (N_11293,N_10241,N_10466);
or U11294 (N_11294,N_9653,N_10321);
xnor U11295 (N_11295,N_9970,N_10414);
xnor U11296 (N_11296,N_9167,N_10497);
xnor U11297 (N_11297,N_9657,N_10479);
and U11298 (N_11298,N_9390,N_9282);
xor U11299 (N_11299,N_10017,N_9935);
or U11300 (N_11300,N_9505,N_9166);
nor U11301 (N_11301,N_9244,N_9835);
or U11302 (N_11302,N_9190,N_9925);
or U11303 (N_11303,N_10028,N_9975);
nor U11304 (N_11304,N_9032,N_10281);
and U11305 (N_11305,N_9043,N_10487);
nand U11306 (N_11306,N_9095,N_9357);
nor U11307 (N_11307,N_10204,N_9643);
nor U11308 (N_11308,N_10024,N_9742);
or U11309 (N_11309,N_9197,N_9656);
and U11310 (N_11310,N_9584,N_9228);
nor U11311 (N_11311,N_10260,N_10286);
or U11312 (N_11312,N_9514,N_10072);
and U11313 (N_11313,N_9696,N_10227);
and U11314 (N_11314,N_9158,N_9035);
xnor U11315 (N_11315,N_10326,N_9437);
and U11316 (N_11316,N_10067,N_9641);
nand U11317 (N_11317,N_9547,N_10437);
and U11318 (N_11318,N_9344,N_9136);
xnor U11319 (N_11319,N_10326,N_9265);
nor U11320 (N_11320,N_10232,N_9915);
nor U11321 (N_11321,N_9978,N_10163);
and U11322 (N_11322,N_9300,N_9019);
xor U11323 (N_11323,N_9255,N_10289);
nand U11324 (N_11324,N_9378,N_10352);
nor U11325 (N_11325,N_10296,N_9921);
xor U11326 (N_11326,N_9310,N_9462);
or U11327 (N_11327,N_10223,N_10425);
nand U11328 (N_11328,N_9202,N_9834);
xnor U11329 (N_11329,N_10376,N_10387);
and U11330 (N_11330,N_10156,N_9192);
or U11331 (N_11331,N_9833,N_10297);
nor U11332 (N_11332,N_10321,N_9329);
and U11333 (N_11333,N_9673,N_10136);
nand U11334 (N_11334,N_9446,N_10262);
or U11335 (N_11335,N_10448,N_10321);
nor U11336 (N_11336,N_9633,N_9974);
xor U11337 (N_11337,N_9553,N_9570);
xor U11338 (N_11338,N_10153,N_10340);
or U11339 (N_11339,N_9290,N_9939);
or U11340 (N_11340,N_9356,N_9362);
and U11341 (N_11341,N_9526,N_9956);
or U11342 (N_11342,N_9087,N_9847);
or U11343 (N_11343,N_9140,N_10429);
xnor U11344 (N_11344,N_10256,N_10151);
xor U11345 (N_11345,N_10287,N_9786);
or U11346 (N_11346,N_9338,N_9129);
and U11347 (N_11347,N_10022,N_9388);
nand U11348 (N_11348,N_9675,N_10432);
xnor U11349 (N_11349,N_10206,N_10291);
or U11350 (N_11350,N_10060,N_9954);
xor U11351 (N_11351,N_9964,N_9908);
and U11352 (N_11352,N_10242,N_9363);
xor U11353 (N_11353,N_9506,N_9845);
and U11354 (N_11354,N_10152,N_9589);
nor U11355 (N_11355,N_9268,N_9028);
or U11356 (N_11356,N_9871,N_9087);
and U11357 (N_11357,N_9298,N_10279);
xnor U11358 (N_11358,N_9139,N_9786);
xnor U11359 (N_11359,N_10140,N_9917);
and U11360 (N_11360,N_9693,N_9189);
or U11361 (N_11361,N_9664,N_9567);
nor U11362 (N_11362,N_10258,N_9955);
nand U11363 (N_11363,N_9027,N_9707);
xor U11364 (N_11364,N_10096,N_10285);
nand U11365 (N_11365,N_10045,N_10124);
nor U11366 (N_11366,N_9237,N_9764);
xnor U11367 (N_11367,N_9501,N_9503);
nor U11368 (N_11368,N_9940,N_10349);
nand U11369 (N_11369,N_9036,N_9919);
xor U11370 (N_11370,N_9004,N_9097);
nor U11371 (N_11371,N_9986,N_10386);
or U11372 (N_11372,N_10480,N_9380);
or U11373 (N_11373,N_9706,N_9197);
xnor U11374 (N_11374,N_9356,N_9297);
nor U11375 (N_11375,N_10497,N_9867);
xnor U11376 (N_11376,N_9322,N_9204);
and U11377 (N_11377,N_10427,N_10271);
or U11378 (N_11378,N_9812,N_9056);
xor U11379 (N_11379,N_10261,N_10195);
or U11380 (N_11380,N_9743,N_10152);
or U11381 (N_11381,N_9753,N_9257);
or U11382 (N_11382,N_9385,N_10103);
and U11383 (N_11383,N_9034,N_9416);
or U11384 (N_11384,N_9087,N_9717);
and U11385 (N_11385,N_10208,N_9203);
xor U11386 (N_11386,N_10137,N_9763);
or U11387 (N_11387,N_10399,N_9835);
and U11388 (N_11388,N_10158,N_9988);
nor U11389 (N_11389,N_10135,N_9860);
or U11390 (N_11390,N_10409,N_9578);
nand U11391 (N_11391,N_10036,N_10074);
or U11392 (N_11392,N_9911,N_9957);
and U11393 (N_11393,N_10109,N_9490);
or U11394 (N_11394,N_9877,N_9197);
nand U11395 (N_11395,N_9862,N_9872);
and U11396 (N_11396,N_9696,N_9385);
xor U11397 (N_11397,N_9902,N_9660);
and U11398 (N_11398,N_9481,N_10228);
xor U11399 (N_11399,N_10018,N_9261);
xnor U11400 (N_11400,N_9126,N_9637);
nand U11401 (N_11401,N_9743,N_9816);
nor U11402 (N_11402,N_9576,N_9206);
or U11403 (N_11403,N_9351,N_9212);
xor U11404 (N_11404,N_9575,N_9117);
and U11405 (N_11405,N_9178,N_9094);
or U11406 (N_11406,N_9402,N_9604);
xnor U11407 (N_11407,N_9656,N_10104);
and U11408 (N_11408,N_9321,N_10003);
xnor U11409 (N_11409,N_9280,N_9885);
xnor U11410 (N_11410,N_9358,N_9475);
nor U11411 (N_11411,N_9551,N_9108);
or U11412 (N_11412,N_9096,N_9212);
nand U11413 (N_11413,N_9757,N_10465);
nor U11414 (N_11414,N_10269,N_9906);
nor U11415 (N_11415,N_9051,N_10272);
or U11416 (N_11416,N_9964,N_10354);
and U11417 (N_11417,N_9488,N_10205);
xor U11418 (N_11418,N_10043,N_9376);
nand U11419 (N_11419,N_9114,N_9514);
and U11420 (N_11420,N_10258,N_10415);
nand U11421 (N_11421,N_9663,N_9375);
xor U11422 (N_11422,N_9187,N_9686);
nor U11423 (N_11423,N_9293,N_9686);
nor U11424 (N_11424,N_9796,N_9701);
xor U11425 (N_11425,N_9592,N_9350);
xor U11426 (N_11426,N_10332,N_9716);
xor U11427 (N_11427,N_10123,N_9242);
or U11428 (N_11428,N_9703,N_9807);
nand U11429 (N_11429,N_10095,N_10169);
nor U11430 (N_11430,N_9622,N_9774);
nand U11431 (N_11431,N_9251,N_9391);
nor U11432 (N_11432,N_10487,N_9713);
xor U11433 (N_11433,N_9454,N_10389);
or U11434 (N_11434,N_9208,N_9596);
nand U11435 (N_11435,N_9860,N_9620);
nand U11436 (N_11436,N_10422,N_10095);
nand U11437 (N_11437,N_9405,N_10334);
or U11438 (N_11438,N_9979,N_10393);
and U11439 (N_11439,N_10363,N_10017);
nor U11440 (N_11440,N_9198,N_9767);
nand U11441 (N_11441,N_9075,N_10118);
nor U11442 (N_11442,N_9048,N_9523);
nand U11443 (N_11443,N_9717,N_9261);
nand U11444 (N_11444,N_9593,N_9224);
nand U11445 (N_11445,N_9691,N_10106);
and U11446 (N_11446,N_10078,N_9544);
nand U11447 (N_11447,N_9632,N_9568);
nand U11448 (N_11448,N_10145,N_9283);
and U11449 (N_11449,N_9038,N_10363);
nor U11450 (N_11450,N_9307,N_10446);
nand U11451 (N_11451,N_9666,N_10185);
xor U11452 (N_11452,N_9347,N_9330);
xor U11453 (N_11453,N_9400,N_10012);
and U11454 (N_11454,N_9356,N_9723);
nand U11455 (N_11455,N_10413,N_9318);
nor U11456 (N_11456,N_9944,N_9552);
nor U11457 (N_11457,N_10305,N_10054);
or U11458 (N_11458,N_9058,N_10452);
or U11459 (N_11459,N_9289,N_9885);
nor U11460 (N_11460,N_10260,N_9045);
nand U11461 (N_11461,N_9757,N_9054);
and U11462 (N_11462,N_9235,N_9244);
or U11463 (N_11463,N_9547,N_9605);
nor U11464 (N_11464,N_9417,N_9791);
nor U11465 (N_11465,N_9942,N_10299);
xor U11466 (N_11466,N_10370,N_9348);
xnor U11467 (N_11467,N_9085,N_9763);
and U11468 (N_11468,N_9111,N_9269);
xnor U11469 (N_11469,N_9213,N_9346);
and U11470 (N_11470,N_10451,N_9725);
nand U11471 (N_11471,N_9216,N_10323);
xor U11472 (N_11472,N_9019,N_10172);
and U11473 (N_11473,N_9243,N_9833);
or U11474 (N_11474,N_10352,N_10171);
xnor U11475 (N_11475,N_9928,N_9217);
and U11476 (N_11476,N_10397,N_9285);
xor U11477 (N_11477,N_10238,N_10061);
and U11478 (N_11478,N_9428,N_9729);
and U11479 (N_11479,N_9602,N_9224);
nor U11480 (N_11480,N_10221,N_10335);
and U11481 (N_11481,N_9555,N_9292);
or U11482 (N_11482,N_9679,N_10057);
or U11483 (N_11483,N_10415,N_10422);
or U11484 (N_11484,N_10192,N_10212);
nand U11485 (N_11485,N_10493,N_9623);
nor U11486 (N_11486,N_10020,N_10035);
nor U11487 (N_11487,N_9268,N_9101);
nor U11488 (N_11488,N_9289,N_10494);
nand U11489 (N_11489,N_10399,N_10043);
nand U11490 (N_11490,N_9374,N_9778);
or U11491 (N_11491,N_9793,N_9515);
and U11492 (N_11492,N_9069,N_10141);
and U11493 (N_11493,N_10077,N_10489);
or U11494 (N_11494,N_10263,N_10439);
xnor U11495 (N_11495,N_9239,N_9703);
nor U11496 (N_11496,N_9118,N_9177);
and U11497 (N_11497,N_10000,N_9827);
or U11498 (N_11498,N_10365,N_9055);
and U11499 (N_11499,N_10147,N_9808);
xnor U11500 (N_11500,N_9279,N_10398);
and U11501 (N_11501,N_9890,N_9807);
nor U11502 (N_11502,N_10111,N_9721);
nor U11503 (N_11503,N_9017,N_9579);
nor U11504 (N_11504,N_10314,N_9915);
xor U11505 (N_11505,N_9921,N_9644);
or U11506 (N_11506,N_9086,N_9426);
and U11507 (N_11507,N_9392,N_9258);
nand U11508 (N_11508,N_9729,N_9662);
xnor U11509 (N_11509,N_9423,N_9848);
xor U11510 (N_11510,N_9551,N_9704);
nand U11511 (N_11511,N_9587,N_9244);
nor U11512 (N_11512,N_9282,N_10247);
xnor U11513 (N_11513,N_9833,N_9513);
and U11514 (N_11514,N_10057,N_9790);
and U11515 (N_11515,N_9784,N_9079);
or U11516 (N_11516,N_9588,N_9021);
nor U11517 (N_11517,N_9226,N_9577);
xor U11518 (N_11518,N_9030,N_9259);
or U11519 (N_11519,N_9069,N_10280);
nand U11520 (N_11520,N_9929,N_10471);
nand U11521 (N_11521,N_9098,N_9394);
xnor U11522 (N_11522,N_9097,N_9986);
nor U11523 (N_11523,N_9855,N_10398);
xnor U11524 (N_11524,N_9361,N_9688);
and U11525 (N_11525,N_9736,N_9172);
or U11526 (N_11526,N_10161,N_9880);
nor U11527 (N_11527,N_10042,N_10016);
nor U11528 (N_11528,N_9693,N_9994);
and U11529 (N_11529,N_9059,N_9288);
xnor U11530 (N_11530,N_9672,N_9050);
nor U11531 (N_11531,N_10332,N_9615);
and U11532 (N_11532,N_9763,N_9191);
nor U11533 (N_11533,N_9839,N_10228);
nor U11534 (N_11534,N_9144,N_9944);
xnor U11535 (N_11535,N_10027,N_9330);
nor U11536 (N_11536,N_10096,N_9763);
nor U11537 (N_11537,N_9569,N_10428);
or U11538 (N_11538,N_10025,N_9178);
nand U11539 (N_11539,N_9260,N_9862);
nand U11540 (N_11540,N_10432,N_9697);
or U11541 (N_11541,N_9381,N_9287);
nand U11542 (N_11542,N_9476,N_9016);
or U11543 (N_11543,N_9749,N_10145);
nor U11544 (N_11544,N_9080,N_9405);
nand U11545 (N_11545,N_10037,N_9317);
nor U11546 (N_11546,N_9623,N_9652);
nor U11547 (N_11547,N_9861,N_10020);
nand U11548 (N_11548,N_10339,N_9638);
nor U11549 (N_11549,N_10350,N_9927);
and U11550 (N_11550,N_9238,N_9960);
and U11551 (N_11551,N_9211,N_9274);
nor U11552 (N_11552,N_9411,N_10144);
nor U11553 (N_11553,N_10464,N_9428);
nor U11554 (N_11554,N_9994,N_9765);
nand U11555 (N_11555,N_9699,N_9053);
nor U11556 (N_11556,N_9504,N_9056);
or U11557 (N_11557,N_9514,N_9477);
nor U11558 (N_11558,N_10406,N_10155);
nor U11559 (N_11559,N_9478,N_9874);
nand U11560 (N_11560,N_10111,N_10120);
and U11561 (N_11561,N_10206,N_10331);
or U11562 (N_11562,N_9642,N_10000);
nand U11563 (N_11563,N_9621,N_10007);
or U11564 (N_11564,N_9985,N_9423);
and U11565 (N_11565,N_9034,N_10423);
or U11566 (N_11566,N_9789,N_9423);
nor U11567 (N_11567,N_9676,N_9635);
xnor U11568 (N_11568,N_9264,N_9518);
or U11569 (N_11569,N_9476,N_9580);
and U11570 (N_11570,N_9048,N_10229);
nand U11571 (N_11571,N_10460,N_9091);
xnor U11572 (N_11572,N_9774,N_9493);
or U11573 (N_11573,N_9908,N_9608);
or U11574 (N_11574,N_9204,N_9761);
or U11575 (N_11575,N_9147,N_9069);
xnor U11576 (N_11576,N_9765,N_9301);
nor U11577 (N_11577,N_10319,N_9874);
nor U11578 (N_11578,N_9125,N_10365);
nand U11579 (N_11579,N_9810,N_9797);
nor U11580 (N_11580,N_10221,N_10490);
nor U11581 (N_11581,N_9145,N_9837);
nor U11582 (N_11582,N_10488,N_10241);
and U11583 (N_11583,N_9801,N_9571);
or U11584 (N_11584,N_10358,N_10124);
and U11585 (N_11585,N_9501,N_10188);
or U11586 (N_11586,N_9633,N_9887);
nor U11587 (N_11587,N_9948,N_9217);
nand U11588 (N_11588,N_9409,N_10310);
nor U11589 (N_11589,N_10426,N_9265);
nor U11590 (N_11590,N_9885,N_9921);
nand U11591 (N_11591,N_10090,N_10120);
or U11592 (N_11592,N_10468,N_9546);
nor U11593 (N_11593,N_9884,N_9824);
xor U11594 (N_11594,N_9450,N_9212);
nand U11595 (N_11595,N_9633,N_10011);
and U11596 (N_11596,N_10432,N_9669);
or U11597 (N_11597,N_9708,N_9211);
or U11598 (N_11598,N_9009,N_9166);
or U11599 (N_11599,N_10163,N_9602);
nand U11600 (N_11600,N_9537,N_9441);
nor U11601 (N_11601,N_10270,N_9550);
and U11602 (N_11602,N_10147,N_9391);
and U11603 (N_11603,N_9425,N_9878);
xnor U11604 (N_11604,N_9615,N_9572);
and U11605 (N_11605,N_9388,N_10214);
and U11606 (N_11606,N_9279,N_10304);
nor U11607 (N_11607,N_9611,N_9687);
nand U11608 (N_11608,N_9052,N_9998);
xor U11609 (N_11609,N_9844,N_9001);
and U11610 (N_11610,N_10192,N_9563);
and U11611 (N_11611,N_9427,N_9072);
xor U11612 (N_11612,N_9839,N_9102);
or U11613 (N_11613,N_9609,N_9879);
xnor U11614 (N_11614,N_9064,N_9231);
xor U11615 (N_11615,N_10238,N_9528);
xor U11616 (N_11616,N_9552,N_10424);
nor U11617 (N_11617,N_9915,N_10345);
and U11618 (N_11618,N_9837,N_9765);
xnor U11619 (N_11619,N_9827,N_9306);
nand U11620 (N_11620,N_9696,N_10277);
nand U11621 (N_11621,N_9664,N_10253);
nor U11622 (N_11622,N_10269,N_9883);
and U11623 (N_11623,N_9886,N_10355);
or U11624 (N_11624,N_9627,N_9054);
and U11625 (N_11625,N_10238,N_9509);
or U11626 (N_11626,N_9466,N_10138);
and U11627 (N_11627,N_9273,N_9637);
and U11628 (N_11628,N_9546,N_10247);
nand U11629 (N_11629,N_9079,N_9637);
nand U11630 (N_11630,N_10153,N_9484);
nand U11631 (N_11631,N_10150,N_9074);
nand U11632 (N_11632,N_9188,N_9763);
nand U11633 (N_11633,N_10416,N_10472);
nor U11634 (N_11634,N_9479,N_10058);
and U11635 (N_11635,N_9822,N_9811);
xor U11636 (N_11636,N_9328,N_9503);
xnor U11637 (N_11637,N_9058,N_9745);
xnor U11638 (N_11638,N_9436,N_9922);
xor U11639 (N_11639,N_9222,N_9975);
and U11640 (N_11640,N_9257,N_9259);
and U11641 (N_11641,N_9420,N_10347);
and U11642 (N_11642,N_10108,N_9013);
and U11643 (N_11643,N_9522,N_10103);
and U11644 (N_11644,N_9242,N_9341);
and U11645 (N_11645,N_9581,N_9769);
xor U11646 (N_11646,N_10290,N_9842);
or U11647 (N_11647,N_10251,N_9884);
or U11648 (N_11648,N_9472,N_9122);
or U11649 (N_11649,N_9240,N_10406);
xnor U11650 (N_11650,N_9061,N_10078);
nor U11651 (N_11651,N_9189,N_9843);
and U11652 (N_11652,N_9726,N_9192);
nand U11653 (N_11653,N_9588,N_10274);
nand U11654 (N_11654,N_9958,N_10024);
xor U11655 (N_11655,N_9537,N_9044);
nor U11656 (N_11656,N_9957,N_9471);
xor U11657 (N_11657,N_9424,N_10316);
or U11658 (N_11658,N_9968,N_10417);
nor U11659 (N_11659,N_9196,N_9201);
nand U11660 (N_11660,N_9785,N_9718);
nand U11661 (N_11661,N_9933,N_10445);
nor U11662 (N_11662,N_9981,N_10007);
nand U11663 (N_11663,N_10109,N_10305);
and U11664 (N_11664,N_9977,N_10286);
nor U11665 (N_11665,N_9266,N_9256);
and U11666 (N_11666,N_10330,N_9494);
nor U11667 (N_11667,N_9653,N_9378);
xor U11668 (N_11668,N_9090,N_9666);
or U11669 (N_11669,N_9543,N_9220);
or U11670 (N_11670,N_9308,N_10375);
and U11671 (N_11671,N_10351,N_10483);
nand U11672 (N_11672,N_9188,N_9661);
xor U11673 (N_11673,N_10072,N_9855);
nor U11674 (N_11674,N_9817,N_10255);
nor U11675 (N_11675,N_9812,N_9889);
nor U11676 (N_11676,N_9565,N_10499);
xor U11677 (N_11677,N_9941,N_10064);
or U11678 (N_11678,N_10203,N_10272);
and U11679 (N_11679,N_9958,N_10014);
and U11680 (N_11680,N_9613,N_9281);
or U11681 (N_11681,N_9345,N_10401);
xnor U11682 (N_11682,N_9326,N_9773);
and U11683 (N_11683,N_9941,N_9545);
nand U11684 (N_11684,N_9724,N_10384);
or U11685 (N_11685,N_9867,N_9040);
and U11686 (N_11686,N_9823,N_10245);
xnor U11687 (N_11687,N_9965,N_10070);
xnor U11688 (N_11688,N_10460,N_10346);
and U11689 (N_11689,N_9264,N_9770);
and U11690 (N_11690,N_10243,N_9310);
and U11691 (N_11691,N_9503,N_9793);
or U11692 (N_11692,N_10451,N_9494);
or U11693 (N_11693,N_10114,N_9489);
nor U11694 (N_11694,N_9632,N_10169);
xnor U11695 (N_11695,N_10362,N_9920);
xor U11696 (N_11696,N_9901,N_9701);
and U11697 (N_11697,N_10183,N_9463);
nor U11698 (N_11698,N_9012,N_9163);
xor U11699 (N_11699,N_9135,N_9087);
and U11700 (N_11700,N_9632,N_9550);
xor U11701 (N_11701,N_9152,N_9376);
xnor U11702 (N_11702,N_9425,N_10042);
xor U11703 (N_11703,N_10043,N_9949);
and U11704 (N_11704,N_10258,N_9970);
nand U11705 (N_11705,N_9925,N_9590);
xnor U11706 (N_11706,N_10263,N_10404);
xnor U11707 (N_11707,N_9723,N_10175);
and U11708 (N_11708,N_9538,N_9224);
xor U11709 (N_11709,N_9771,N_10256);
and U11710 (N_11710,N_9238,N_10279);
xnor U11711 (N_11711,N_9791,N_10111);
or U11712 (N_11712,N_10372,N_10299);
nand U11713 (N_11713,N_9390,N_9936);
nand U11714 (N_11714,N_9623,N_9985);
nand U11715 (N_11715,N_10459,N_9693);
xnor U11716 (N_11716,N_9042,N_9371);
nor U11717 (N_11717,N_9799,N_9159);
or U11718 (N_11718,N_10090,N_10105);
xnor U11719 (N_11719,N_9008,N_9567);
nand U11720 (N_11720,N_9807,N_10065);
nor U11721 (N_11721,N_9848,N_9297);
or U11722 (N_11722,N_9598,N_9322);
or U11723 (N_11723,N_10379,N_9839);
nor U11724 (N_11724,N_9702,N_9382);
or U11725 (N_11725,N_9470,N_10333);
nand U11726 (N_11726,N_9153,N_9524);
xor U11727 (N_11727,N_9515,N_9705);
nand U11728 (N_11728,N_9855,N_9169);
nand U11729 (N_11729,N_9882,N_9001);
or U11730 (N_11730,N_9536,N_9300);
and U11731 (N_11731,N_10090,N_10293);
xor U11732 (N_11732,N_9571,N_9314);
or U11733 (N_11733,N_10121,N_9649);
or U11734 (N_11734,N_9384,N_9406);
or U11735 (N_11735,N_9226,N_10302);
and U11736 (N_11736,N_9898,N_9219);
or U11737 (N_11737,N_9759,N_10301);
nand U11738 (N_11738,N_9644,N_9518);
nand U11739 (N_11739,N_10002,N_10473);
xor U11740 (N_11740,N_10284,N_10143);
or U11741 (N_11741,N_10154,N_9550);
and U11742 (N_11742,N_9133,N_9700);
and U11743 (N_11743,N_9428,N_9335);
nand U11744 (N_11744,N_10493,N_9868);
nor U11745 (N_11745,N_9107,N_10172);
nor U11746 (N_11746,N_9679,N_9004);
and U11747 (N_11747,N_9361,N_9030);
and U11748 (N_11748,N_9074,N_9528);
nor U11749 (N_11749,N_9325,N_10030);
nand U11750 (N_11750,N_9817,N_9013);
nor U11751 (N_11751,N_9101,N_9665);
nand U11752 (N_11752,N_9389,N_10441);
xor U11753 (N_11753,N_9523,N_9564);
xor U11754 (N_11754,N_10400,N_10345);
nor U11755 (N_11755,N_9994,N_9894);
nand U11756 (N_11756,N_10394,N_9165);
nand U11757 (N_11757,N_9554,N_10437);
nor U11758 (N_11758,N_9596,N_9683);
xor U11759 (N_11759,N_9790,N_10187);
xnor U11760 (N_11760,N_9627,N_10085);
nand U11761 (N_11761,N_10147,N_10444);
xor U11762 (N_11762,N_9643,N_9379);
or U11763 (N_11763,N_9826,N_9662);
or U11764 (N_11764,N_9359,N_9425);
and U11765 (N_11765,N_9406,N_9713);
or U11766 (N_11766,N_10203,N_9492);
nor U11767 (N_11767,N_9396,N_9548);
nor U11768 (N_11768,N_9283,N_9988);
nor U11769 (N_11769,N_10231,N_10271);
nor U11770 (N_11770,N_9521,N_9221);
xnor U11771 (N_11771,N_9080,N_9728);
nand U11772 (N_11772,N_9554,N_10094);
xor U11773 (N_11773,N_9526,N_9422);
nand U11774 (N_11774,N_10393,N_9843);
and U11775 (N_11775,N_9150,N_9831);
nor U11776 (N_11776,N_9542,N_9563);
and U11777 (N_11777,N_10304,N_9635);
nand U11778 (N_11778,N_10470,N_9360);
nor U11779 (N_11779,N_10136,N_10281);
xor U11780 (N_11780,N_9214,N_9628);
and U11781 (N_11781,N_9318,N_9863);
and U11782 (N_11782,N_9439,N_9891);
xor U11783 (N_11783,N_9461,N_9797);
xnor U11784 (N_11784,N_9229,N_9204);
nand U11785 (N_11785,N_10191,N_9634);
or U11786 (N_11786,N_9769,N_9233);
and U11787 (N_11787,N_9644,N_9401);
or U11788 (N_11788,N_9489,N_9494);
nor U11789 (N_11789,N_9169,N_10374);
or U11790 (N_11790,N_10337,N_9467);
and U11791 (N_11791,N_9844,N_10186);
and U11792 (N_11792,N_9388,N_9505);
or U11793 (N_11793,N_9395,N_10381);
nor U11794 (N_11794,N_10464,N_10374);
xor U11795 (N_11795,N_9247,N_10223);
nor U11796 (N_11796,N_9031,N_9334);
nand U11797 (N_11797,N_10350,N_9846);
xnor U11798 (N_11798,N_10308,N_9473);
nor U11799 (N_11799,N_10204,N_9358);
nand U11800 (N_11800,N_9671,N_9667);
or U11801 (N_11801,N_10431,N_9877);
or U11802 (N_11802,N_9590,N_9263);
nand U11803 (N_11803,N_9603,N_10497);
nand U11804 (N_11804,N_9268,N_9534);
or U11805 (N_11805,N_10166,N_10444);
nand U11806 (N_11806,N_9481,N_10401);
or U11807 (N_11807,N_9026,N_9448);
nand U11808 (N_11808,N_9645,N_10264);
or U11809 (N_11809,N_9474,N_10126);
or U11810 (N_11810,N_9160,N_9971);
and U11811 (N_11811,N_10373,N_9385);
and U11812 (N_11812,N_9674,N_10210);
nor U11813 (N_11813,N_10477,N_10370);
nor U11814 (N_11814,N_10122,N_10402);
nand U11815 (N_11815,N_10178,N_9677);
and U11816 (N_11816,N_9535,N_9852);
nand U11817 (N_11817,N_9152,N_9499);
or U11818 (N_11818,N_10015,N_10434);
xor U11819 (N_11819,N_10472,N_9184);
nand U11820 (N_11820,N_9176,N_9598);
or U11821 (N_11821,N_10059,N_10103);
or U11822 (N_11822,N_9466,N_9952);
and U11823 (N_11823,N_9457,N_9310);
nand U11824 (N_11824,N_9153,N_10458);
and U11825 (N_11825,N_9897,N_9274);
nor U11826 (N_11826,N_9099,N_9594);
nand U11827 (N_11827,N_10124,N_9645);
and U11828 (N_11828,N_9796,N_9030);
or U11829 (N_11829,N_9948,N_9945);
and U11830 (N_11830,N_10423,N_9771);
nand U11831 (N_11831,N_9241,N_9337);
or U11832 (N_11832,N_9736,N_9199);
or U11833 (N_11833,N_9103,N_10259);
nand U11834 (N_11834,N_9225,N_9698);
xor U11835 (N_11835,N_9760,N_9133);
nor U11836 (N_11836,N_10255,N_10465);
nor U11837 (N_11837,N_10218,N_9676);
nor U11838 (N_11838,N_10292,N_9977);
nor U11839 (N_11839,N_10211,N_9078);
or U11840 (N_11840,N_9194,N_9366);
nand U11841 (N_11841,N_9099,N_9569);
or U11842 (N_11842,N_9976,N_10140);
and U11843 (N_11843,N_10158,N_9849);
nor U11844 (N_11844,N_10421,N_9779);
nor U11845 (N_11845,N_9999,N_9987);
and U11846 (N_11846,N_10312,N_9785);
nand U11847 (N_11847,N_9051,N_9586);
or U11848 (N_11848,N_9398,N_9337);
nor U11849 (N_11849,N_9445,N_10330);
nor U11850 (N_11850,N_9753,N_9306);
nor U11851 (N_11851,N_9877,N_9527);
nor U11852 (N_11852,N_9914,N_10436);
or U11853 (N_11853,N_9751,N_9683);
nor U11854 (N_11854,N_9439,N_10392);
or U11855 (N_11855,N_9896,N_9598);
nand U11856 (N_11856,N_9145,N_9940);
or U11857 (N_11857,N_9229,N_10098);
nor U11858 (N_11858,N_9212,N_9124);
and U11859 (N_11859,N_10215,N_10327);
or U11860 (N_11860,N_9600,N_10325);
nand U11861 (N_11861,N_10021,N_10242);
or U11862 (N_11862,N_10119,N_10138);
nand U11863 (N_11863,N_9699,N_10253);
nand U11864 (N_11864,N_9101,N_9412);
xor U11865 (N_11865,N_9069,N_9755);
and U11866 (N_11866,N_9437,N_9638);
nand U11867 (N_11867,N_10091,N_10174);
nor U11868 (N_11868,N_9410,N_9166);
nand U11869 (N_11869,N_9974,N_9142);
nand U11870 (N_11870,N_9966,N_10130);
nor U11871 (N_11871,N_9633,N_9773);
nor U11872 (N_11872,N_10272,N_10017);
and U11873 (N_11873,N_10355,N_9545);
xor U11874 (N_11874,N_9288,N_10358);
or U11875 (N_11875,N_9891,N_9600);
nor U11876 (N_11876,N_9206,N_9622);
or U11877 (N_11877,N_9425,N_9708);
nor U11878 (N_11878,N_9292,N_9001);
or U11879 (N_11879,N_10169,N_9192);
and U11880 (N_11880,N_10137,N_10447);
nand U11881 (N_11881,N_10195,N_9572);
and U11882 (N_11882,N_10010,N_10360);
nor U11883 (N_11883,N_9399,N_10118);
and U11884 (N_11884,N_9805,N_9358);
nor U11885 (N_11885,N_9468,N_10252);
xnor U11886 (N_11886,N_10336,N_9472);
xnor U11887 (N_11887,N_10344,N_10168);
xnor U11888 (N_11888,N_9539,N_9919);
and U11889 (N_11889,N_10036,N_9127);
and U11890 (N_11890,N_10276,N_9097);
or U11891 (N_11891,N_9166,N_9582);
nand U11892 (N_11892,N_9064,N_10101);
xor U11893 (N_11893,N_9702,N_9732);
and U11894 (N_11894,N_9836,N_9585);
and U11895 (N_11895,N_10160,N_9231);
and U11896 (N_11896,N_9518,N_9824);
nor U11897 (N_11897,N_9243,N_9139);
xnor U11898 (N_11898,N_10020,N_9513);
and U11899 (N_11899,N_10186,N_9229);
xnor U11900 (N_11900,N_9892,N_10123);
nor U11901 (N_11901,N_10037,N_10000);
and U11902 (N_11902,N_10407,N_9627);
and U11903 (N_11903,N_9946,N_10457);
and U11904 (N_11904,N_9427,N_10277);
and U11905 (N_11905,N_10030,N_9076);
or U11906 (N_11906,N_9508,N_9369);
xnor U11907 (N_11907,N_9193,N_9298);
and U11908 (N_11908,N_10143,N_9995);
or U11909 (N_11909,N_10312,N_9596);
nor U11910 (N_11910,N_10024,N_9503);
or U11911 (N_11911,N_10466,N_9821);
nor U11912 (N_11912,N_9049,N_9733);
nor U11913 (N_11913,N_9949,N_10258);
or U11914 (N_11914,N_9398,N_9298);
or U11915 (N_11915,N_9935,N_9230);
xnor U11916 (N_11916,N_9928,N_9360);
nor U11917 (N_11917,N_10053,N_10012);
nand U11918 (N_11918,N_9256,N_9576);
xor U11919 (N_11919,N_9777,N_9536);
nor U11920 (N_11920,N_10185,N_9762);
nand U11921 (N_11921,N_9827,N_10499);
nand U11922 (N_11922,N_9644,N_9134);
nand U11923 (N_11923,N_9073,N_9850);
nand U11924 (N_11924,N_10445,N_10311);
nor U11925 (N_11925,N_10031,N_10382);
nor U11926 (N_11926,N_10199,N_9543);
and U11927 (N_11927,N_10294,N_10318);
nor U11928 (N_11928,N_9940,N_9529);
nand U11929 (N_11929,N_10295,N_9282);
or U11930 (N_11930,N_9284,N_9008);
nand U11931 (N_11931,N_10461,N_9477);
nor U11932 (N_11932,N_9384,N_9595);
xor U11933 (N_11933,N_10301,N_9868);
or U11934 (N_11934,N_9884,N_9514);
or U11935 (N_11935,N_10132,N_9420);
and U11936 (N_11936,N_9320,N_10233);
nand U11937 (N_11937,N_9375,N_10358);
nand U11938 (N_11938,N_9940,N_9290);
and U11939 (N_11939,N_9642,N_9096);
and U11940 (N_11940,N_9029,N_9683);
nor U11941 (N_11941,N_10398,N_9986);
or U11942 (N_11942,N_9235,N_9942);
or U11943 (N_11943,N_10050,N_9474);
nor U11944 (N_11944,N_9596,N_10478);
and U11945 (N_11945,N_10095,N_10245);
and U11946 (N_11946,N_10390,N_9417);
nor U11947 (N_11947,N_9463,N_9461);
xnor U11948 (N_11948,N_10406,N_9261);
xor U11949 (N_11949,N_10415,N_9656);
nor U11950 (N_11950,N_9494,N_9193);
nand U11951 (N_11951,N_9962,N_9470);
and U11952 (N_11952,N_10078,N_9722);
or U11953 (N_11953,N_9668,N_10164);
nor U11954 (N_11954,N_10401,N_10050);
and U11955 (N_11955,N_10197,N_9122);
nor U11956 (N_11956,N_9567,N_9767);
or U11957 (N_11957,N_9185,N_10124);
and U11958 (N_11958,N_9633,N_10271);
nand U11959 (N_11959,N_9823,N_9126);
nand U11960 (N_11960,N_10286,N_9109);
xor U11961 (N_11961,N_9354,N_9215);
xor U11962 (N_11962,N_9424,N_10210);
nand U11963 (N_11963,N_10308,N_9366);
xnor U11964 (N_11964,N_9247,N_9183);
nand U11965 (N_11965,N_10125,N_10061);
and U11966 (N_11966,N_9561,N_9238);
and U11967 (N_11967,N_9698,N_9780);
and U11968 (N_11968,N_9270,N_9692);
nor U11969 (N_11969,N_9543,N_9042);
nand U11970 (N_11970,N_10054,N_9375);
and U11971 (N_11971,N_9148,N_9035);
nand U11972 (N_11972,N_9136,N_9026);
xor U11973 (N_11973,N_9659,N_10060);
and U11974 (N_11974,N_9998,N_9624);
and U11975 (N_11975,N_9645,N_10237);
nor U11976 (N_11976,N_9726,N_9702);
or U11977 (N_11977,N_9738,N_9361);
nor U11978 (N_11978,N_10124,N_9030);
or U11979 (N_11979,N_9154,N_9918);
and U11980 (N_11980,N_9166,N_9338);
xnor U11981 (N_11981,N_9205,N_9288);
or U11982 (N_11982,N_9100,N_9403);
nand U11983 (N_11983,N_10080,N_9638);
nand U11984 (N_11984,N_9148,N_9337);
nand U11985 (N_11985,N_9792,N_9354);
nand U11986 (N_11986,N_9200,N_9873);
nand U11987 (N_11987,N_9210,N_10101);
and U11988 (N_11988,N_9963,N_9754);
nor U11989 (N_11989,N_9132,N_10185);
and U11990 (N_11990,N_10266,N_9170);
nand U11991 (N_11991,N_9422,N_10010);
and U11992 (N_11992,N_10408,N_9046);
or U11993 (N_11993,N_9753,N_9705);
xnor U11994 (N_11994,N_10141,N_10413);
or U11995 (N_11995,N_10132,N_9821);
xor U11996 (N_11996,N_9472,N_9597);
and U11997 (N_11997,N_9482,N_9259);
and U11998 (N_11998,N_9797,N_10306);
and U11999 (N_11999,N_9676,N_9815);
nand U12000 (N_12000,N_11207,N_11861);
nor U12001 (N_12001,N_10610,N_11382);
nand U12002 (N_12002,N_11587,N_11124);
nor U12003 (N_12003,N_11695,N_11626);
or U12004 (N_12004,N_10694,N_11858);
nor U12005 (N_12005,N_10739,N_11167);
or U12006 (N_12006,N_10619,N_11015);
nor U12007 (N_12007,N_10886,N_10862);
nor U12008 (N_12008,N_10945,N_10579);
or U12009 (N_12009,N_11939,N_10741);
nand U12010 (N_12010,N_10680,N_11044);
and U12011 (N_12011,N_10690,N_10667);
nand U12012 (N_12012,N_10730,N_11938);
nor U12013 (N_12013,N_10659,N_11490);
xnor U12014 (N_12014,N_11312,N_10750);
nor U12015 (N_12015,N_10900,N_11025);
xnor U12016 (N_12016,N_11842,N_10996);
or U12017 (N_12017,N_11914,N_10705);
nor U12018 (N_12018,N_10774,N_11008);
xor U12019 (N_12019,N_11867,N_11644);
xnor U12020 (N_12020,N_11792,N_10989);
and U12021 (N_12021,N_11331,N_10547);
and U12022 (N_12022,N_10829,N_11708);
xor U12023 (N_12023,N_10695,N_11463);
or U12024 (N_12024,N_10798,N_11972);
or U12025 (N_12025,N_11170,N_11298);
xnor U12026 (N_12026,N_11163,N_11229);
nand U12027 (N_12027,N_11430,N_10646);
nor U12028 (N_12028,N_11558,N_10832);
or U12029 (N_12029,N_11397,N_11948);
and U12030 (N_12030,N_11234,N_10558);
and U12031 (N_12031,N_10870,N_10743);
nand U12032 (N_12032,N_11789,N_11760);
nor U12033 (N_12033,N_11765,N_11955);
nor U12034 (N_12034,N_11053,N_11109);
or U12035 (N_12035,N_11050,N_11403);
or U12036 (N_12036,N_11685,N_10665);
xor U12037 (N_12037,N_11546,N_10561);
nand U12038 (N_12038,N_11652,N_10985);
xnor U12039 (N_12039,N_11970,N_11641);
nand U12040 (N_12040,N_11992,N_10863);
nor U12041 (N_12041,N_10508,N_10591);
xnor U12042 (N_12042,N_11359,N_11636);
xor U12043 (N_12043,N_10633,N_11584);
nor U12044 (N_12044,N_10556,N_11432);
or U12045 (N_12045,N_10766,N_11889);
or U12046 (N_12046,N_11217,N_10930);
nor U12047 (N_12047,N_11950,N_11277);
and U12048 (N_12048,N_10603,N_11780);
xor U12049 (N_12049,N_11774,N_11705);
xor U12050 (N_12050,N_11758,N_11521);
nor U12051 (N_12051,N_11005,N_11306);
or U12052 (N_12052,N_10772,N_10907);
or U12053 (N_12053,N_10581,N_10614);
nand U12054 (N_12054,N_11986,N_11173);
and U12055 (N_12055,N_11850,N_10967);
or U12056 (N_12056,N_11085,N_11341);
or U12057 (N_12057,N_11784,N_11667);
nor U12058 (N_12058,N_11425,N_10947);
and U12059 (N_12059,N_11419,N_10812);
or U12060 (N_12060,N_11872,N_11535);
or U12061 (N_12061,N_11480,N_11391);
or U12062 (N_12062,N_11960,N_11361);
nor U12063 (N_12063,N_11372,N_11037);
xnor U12064 (N_12064,N_11912,N_11804);
and U12065 (N_12065,N_11334,N_11832);
or U12066 (N_12066,N_11296,N_10532);
xor U12067 (N_12067,N_10575,N_11866);
nand U12068 (N_12068,N_11919,N_11937);
or U12069 (N_12069,N_11568,N_11639);
nand U12070 (N_12070,N_10510,N_11056);
nor U12071 (N_12071,N_11544,N_10613);
xor U12072 (N_12072,N_11379,N_11615);
nor U12073 (N_12073,N_11893,N_10745);
and U12074 (N_12074,N_11766,N_11770);
or U12075 (N_12075,N_11680,N_11886);
and U12076 (N_12076,N_10800,N_11930);
nand U12077 (N_12077,N_11745,N_11001);
nand U12078 (N_12078,N_10987,N_11625);
nand U12079 (N_12079,N_10854,N_10871);
and U12080 (N_12080,N_11579,N_11031);
and U12081 (N_12081,N_10894,N_10818);
nand U12082 (N_12082,N_10916,N_11859);
nand U12083 (N_12083,N_10938,N_10615);
nor U12084 (N_12084,N_10569,N_11997);
and U12085 (N_12085,N_11420,N_11462);
and U12086 (N_12086,N_10504,N_11483);
and U12087 (N_12087,N_11357,N_11895);
nand U12088 (N_12088,N_11876,N_11197);
and U12089 (N_12089,N_11437,N_10757);
or U12090 (N_12090,N_10568,N_11089);
or U12091 (N_12091,N_11291,N_10632);
and U12092 (N_12092,N_11776,N_10959);
nor U12093 (N_12093,N_11840,N_11367);
or U12094 (N_12094,N_11067,N_10681);
or U12095 (N_12095,N_11487,N_11057);
xor U12096 (N_12096,N_11346,N_10605);
xor U12097 (N_12097,N_11692,N_11389);
nor U12098 (N_12098,N_11900,N_10551);
nand U12099 (N_12099,N_11714,N_11473);
xor U12100 (N_12100,N_10697,N_11035);
and U12101 (N_12101,N_11848,N_11278);
xnor U12102 (N_12102,N_11009,N_11923);
or U12103 (N_12103,N_11141,N_10597);
nand U12104 (N_12104,N_10638,N_10618);
nor U12105 (N_12105,N_11325,N_11801);
nor U12106 (N_12106,N_10767,N_11024);
or U12107 (N_12107,N_10785,N_11411);
xor U12108 (N_12108,N_11777,N_11402);
and U12109 (N_12109,N_11224,N_11538);
and U12110 (N_12110,N_11469,N_11570);
nand U12111 (N_12111,N_10627,N_11059);
or U12112 (N_12112,N_10554,N_11012);
or U12113 (N_12113,N_10761,N_11604);
nor U12114 (N_12114,N_11511,N_10799);
xnor U12115 (N_12115,N_11308,N_10736);
nand U12116 (N_12116,N_11103,N_11808);
nand U12117 (N_12117,N_11246,N_11724);
nor U12118 (N_12118,N_11622,N_11450);
and U12119 (N_12119,N_11655,N_11128);
and U12120 (N_12120,N_11703,N_10587);
nand U12121 (N_12121,N_11201,N_11710);
xor U12122 (N_12122,N_11422,N_11356);
xnor U12123 (N_12123,N_11623,N_11534);
xor U12124 (N_12124,N_11581,N_10816);
and U12125 (N_12125,N_11415,N_11529);
xnor U12126 (N_12126,N_11360,N_10570);
xnor U12127 (N_12127,N_10981,N_10713);
or U12128 (N_12128,N_10949,N_11741);
nor U12129 (N_12129,N_11821,N_11845);
nor U12130 (N_12130,N_10759,N_11275);
xnor U12131 (N_12131,N_11018,N_11851);
and U12132 (N_12132,N_10727,N_11995);
nor U12133 (N_12133,N_11384,N_10936);
nor U12134 (N_12134,N_10715,N_10563);
nand U12135 (N_12135,N_10545,N_11152);
xnor U12136 (N_12136,N_10933,N_11079);
xor U12137 (N_12137,N_10887,N_11916);
or U12138 (N_12138,N_11526,N_10926);
nand U12139 (N_12139,N_11971,N_11349);
or U12140 (N_12140,N_10540,N_11922);
and U12141 (N_12141,N_11294,N_10884);
and U12142 (N_12142,N_11879,N_10523);
and U12143 (N_12143,N_11310,N_10837);
nand U12144 (N_12144,N_11525,N_11825);
and U12145 (N_12145,N_11449,N_10789);
and U12146 (N_12146,N_10566,N_11027);
or U12147 (N_12147,N_11178,N_11390);
nand U12148 (N_12148,N_11728,N_11934);
and U12149 (N_12149,N_11385,N_11907);
nand U12150 (N_12150,N_10534,N_11678);
nor U12151 (N_12151,N_11899,N_10795);
nand U12152 (N_12152,N_11863,N_11259);
or U12153 (N_12153,N_11701,N_11924);
nor U12154 (N_12154,N_11453,N_11285);
xor U12155 (N_12155,N_11691,N_10904);
or U12156 (N_12156,N_11965,N_10686);
nor U12157 (N_12157,N_11102,N_11738);
xor U12158 (N_12158,N_11654,N_10637);
nor U12159 (N_12159,N_10892,N_10973);
nor U12160 (N_12160,N_11989,N_10920);
and U12161 (N_12161,N_10810,N_11022);
xnor U12162 (N_12162,N_11495,N_11790);
nand U12163 (N_12163,N_10879,N_10675);
and U12164 (N_12164,N_11265,N_11322);
nand U12165 (N_12165,N_11504,N_11052);
xnor U12166 (N_12166,N_11693,N_11286);
and U12167 (N_12167,N_10762,N_11198);
nand U12168 (N_12168,N_10919,N_10609);
xor U12169 (N_12169,N_11806,N_10662);
nand U12170 (N_12170,N_11497,N_11836);
or U12171 (N_12171,N_11439,N_11176);
or U12172 (N_12172,N_11248,N_11093);
nand U12173 (N_12173,N_11061,N_10738);
xnor U12174 (N_12174,N_10527,N_11958);
nor U12175 (N_12175,N_11250,N_11712);
nor U12176 (N_12176,N_10602,N_11864);
and U12177 (N_12177,N_11110,N_10855);
xor U12178 (N_12178,N_11791,N_11984);
nand U12179 (N_12179,N_11470,N_11206);
nand U12180 (N_12180,N_11720,N_11146);
and U12181 (N_12181,N_10714,N_11540);
nor U12182 (N_12182,N_11795,N_11165);
xor U12183 (N_12183,N_11560,N_11476);
xor U12184 (N_12184,N_11660,N_11139);
or U12185 (N_12185,N_11394,N_11976);
or U12186 (N_12186,N_10806,N_10895);
nand U12187 (N_12187,N_10807,N_11066);
and U12188 (N_12188,N_11663,N_11253);
or U12189 (N_12189,N_10903,N_11761);
and U12190 (N_12190,N_11877,N_11466);
xnor U12191 (N_12191,N_11751,N_10625);
nand U12192 (N_12192,N_10507,N_11162);
xnor U12193 (N_12193,N_10629,N_11482);
or U12194 (N_12194,N_11562,N_11287);
or U12195 (N_12195,N_10771,N_11004);
and U12196 (N_12196,N_10636,N_10653);
nand U12197 (N_12197,N_11078,N_11671);
and U12198 (N_12198,N_11120,N_11313);
xnor U12199 (N_12199,N_11664,N_10849);
nand U12200 (N_12200,N_10931,N_10525);
nor U12201 (N_12201,N_11441,N_10984);
nor U12202 (N_12202,N_10639,N_10821);
xor U12203 (N_12203,N_11177,N_11068);
or U12204 (N_12204,N_10817,N_10823);
and U12205 (N_12205,N_11537,N_10850);
xnor U12206 (N_12206,N_10711,N_11682);
nand U12207 (N_12207,N_11672,N_11396);
or U12208 (N_12208,N_11953,N_11817);
or U12209 (N_12209,N_10994,N_11943);
nand U12210 (N_12210,N_11301,N_11918);
and U12211 (N_12211,N_11576,N_10718);
xor U12212 (N_12212,N_11481,N_11326);
nand U12213 (N_12213,N_11247,N_11041);
xnor U12214 (N_12214,N_11257,N_11557);
or U12215 (N_12215,N_11764,N_11181);
or U12216 (N_12216,N_10642,N_10872);
or U12217 (N_12217,N_11029,N_11589);
xor U12218 (N_12218,N_11266,N_10852);
or U12219 (N_12219,N_11122,N_11147);
xor U12220 (N_12220,N_11271,N_11186);
nand U12221 (N_12221,N_11548,N_10943);
and U12222 (N_12222,N_11182,N_11945);
xnor U12223 (N_12223,N_11952,N_11405);
nor U12224 (N_12224,N_11552,N_10896);
nand U12225 (N_12225,N_10873,N_11601);
xnor U12226 (N_12226,N_10623,N_10787);
and U12227 (N_12227,N_11588,N_11594);
nand U12228 (N_12228,N_11319,N_11330);
xnor U12229 (N_12229,N_11602,N_10924);
and U12230 (N_12230,N_11797,N_11375);
xor U12231 (N_12231,N_11135,N_11794);
nor U12232 (N_12232,N_11125,N_10600);
nor U12233 (N_12233,N_11966,N_11737);
xor U12234 (N_12234,N_11489,N_11337);
nor U12235 (N_12235,N_11169,N_10846);
xnor U12236 (N_12236,N_11456,N_11716);
xnor U12237 (N_12237,N_11670,N_11071);
nor U12238 (N_12238,N_11095,N_10997);
nor U12239 (N_12239,N_11688,N_11108);
nor U12240 (N_12240,N_10780,N_11957);
xor U12241 (N_12241,N_10788,N_11718);
xor U12242 (N_12242,N_11827,N_11216);
and U12243 (N_12243,N_11392,N_10840);
xnor U12244 (N_12244,N_10669,N_10932);
nand U12245 (N_12245,N_10797,N_11669);
nand U12246 (N_12246,N_10670,N_10564);
nand U12247 (N_12247,N_10515,N_11807);
xor U12248 (N_12248,N_11896,N_11111);
or U12249 (N_12249,N_11339,N_11857);
xnor U12250 (N_12250,N_11533,N_11947);
and U12251 (N_12251,N_11767,N_10843);
nor U12252 (N_12252,N_11309,N_10918);
nor U12253 (N_12253,N_11157,N_10604);
xnor U12254 (N_12254,N_10553,N_11969);
and U12255 (N_12255,N_10781,N_11909);
and U12256 (N_12256,N_11689,N_11846);
nand U12257 (N_12257,N_11129,N_11276);
or U12258 (N_12258,N_10988,N_11028);
nand U12259 (N_12259,N_11898,N_11903);
and U12260 (N_12260,N_11818,N_11661);
nor U12261 (N_12261,N_11320,N_11475);
or U12262 (N_12262,N_10733,N_10687);
nand U12263 (N_12263,N_11090,N_11344);
or U12264 (N_12264,N_11782,N_11822);
nand U12265 (N_12265,N_10684,N_11399);
xnor U12266 (N_12266,N_11648,N_11561);
xor U12267 (N_12267,N_10595,N_10502);
and U12268 (N_12268,N_11510,N_11179);
xor U12269 (N_12269,N_11200,N_10572);
and U12270 (N_12270,N_11016,N_11532);
xor U12271 (N_12271,N_10722,N_10844);
and U12272 (N_12272,N_11920,N_11666);
xnor U12273 (N_12273,N_11910,N_11263);
nor U12274 (N_12274,N_11940,N_11023);
nor U12275 (N_12275,N_10869,N_11335);
or U12276 (N_12276,N_11500,N_11964);
or U12277 (N_12277,N_11184,N_11904);
nand U12278 (N_12278,N_10897,N_11161);
and U12279 (N_12279,N_11355,N_10702);
xor U12280 (N_12280,N_10803,N_11395);
or U12281 (N_12281,N_11743,N_11192);
and U12282 (N_12282,N_10954,N_10822);
nor U12283 (N_12283,N_11010,N_10899);
nor U12284 (N_12284,N_11194,N_11084);
or U12285 (N_12285,N_11032,N_11815);
nand U12286 (N_12286,N_10674,N_11739);
nor U12287 (N_12287,N_11871,N_11047);
nand U12288 (N_12288,N_11119,N_10891);
nand U12289 (N_12289,N_10972,N_11921);
or U12290 (N_12290,N_11592,N_11779);
nand U12291 (N_12291,N_11932,N_11150);
xor U12292 (N_12292,N_11569,N_10621);
nand U12293 (N_12293,N_11933,N_10731);
xnor U12294 (N_12294,N_11172,N_11493);
and U12295 (N_12295,N_11811,N_11731);
nand U12296 (N_12296,N_10965,N_11034);
xor U12297 (N_12297,N_11369,N_10616);
nand U12298 (N_12298,N_10875,N_11987);
nor U12299 (N_12299,N_10848,N_11843);
xnor U12300 (N_12300,N_11781,N_10533);
and U12301 (N_12301,N_10598,N_10866);
or U12302 (N_12302,N_11892,N_11599);
nand U12303 (N_12303,N_11347,N_10661);
nand U12304 (N_12304,N_10951,N_11171);
nand U12305 (N_12305,N_11227,N_10881);
nor U12306 (N_12306,N_10794,N_10939);
and U12307 (N_12307,N_11824,N_11734);
nand U12308 (N_12308,N_11088,N_11222);
or U12309 (N_12309,N_11293,N_11830);
nand U12310 (N_12310,N_10631,N_11282);
xnor U12311 (N_12311,N_11659,N_10728);
or U12312 (N_12312,N_11515,N_11798);
xnor U12313 (N_12313,N_10503,N_10763);
nor U12314 (N_12314,N_11638,N_11199);
nand U12315 (N_12315,N_11613,N_11645);
nor U12316 (N_12316,N_10970,N_11160);
nor U12317 (N_12317,N_10912,N_10580);
or U12318 (N_12318,N_11284,N_10864);
xor U12319 (N_12319,N_10856,N_11702);
nor U12320 (N_12320,N_11144,N_11094);
xor U12321 (N_12321,N_11017,N_10567);
or U12322 (N_12322,N_11273,N_11438);
nand U12323 (N_12323,N_10543,N_11077);
nor U12324 (N_12324,N_11772,N_11193);
and U12325 (N_12325,N_11829,N_10833);
nand U12326 (N_12326,N_10660,N_11956);
xor U12327 (N_12327,N_10805,N_11563);
and U12328 (N_12328,N_11793,N_11646);
nor U12329 (N_12329,N_11267,N_11598);
nor U12330 (N_12330,N_11611,N_11926);
nor U12331 (N_12331,N_11106,N_10557);
or U12332 (N_12332,N_10548,N_11358);
xnor U12333 (N_12333,N_11819,N_11255);
or U12334 (N_12334,N_10992,N_10902);
xor U12335 (N_12335,N_11474,N_11136);
nand U12336 (N_12336,N_10993,N_10699);
nand U12337 (N_12337,N_10808,N_11556);
nor U12338 (N_12338,N_10878,N_11159);
and U12339 (N_12339,N_10905,N_10544);
nand U12340 (N_12340,N_11074,N_10768);
or U12341 (N_12341,N_10647,N_11468);
or U12342 (N_12342,N_11985,N_10552);
and U12343 (N_12343,N_11213,N_11058);
nand U12344 (N_12344,N_10673,N_11060);
or U12345 (N_12345,N_11762,N_11244);
nand U12346 (N_12346,N_11049,N_11467);
and U12347 (N_12347,N_10783,N_10980);
nor U12348 (N_12348,N_11913,N_11717);
nor U12349 (N_12349,N_11501,N_11874);
nor U12350 (N_12350,N_11578,N_10860);
and U12351 (N_12351,N_11917,N_10644);
and U12352 (N_12352,N_11107,N_10550);
and U12353 (N_12353,N_11214,N_10958);
xnor U12354 (N_12354,N_10582,N_11342);
nor U12355 (N_12355,N_10546,N_11885);
nor U12356 (N_12356,N_11547,N_11826);
nor U12357 (N_12357,N_11911,N_11404);
xnor U12358 (N_12358,N_11513,N_10979);
nand U12359 (N_12359,N_11567,N_11749);
nand U12360 (N_12360,N_11092,N_10672);
nor U12361 (N_12361,N_11366,N_11834);
xnor U12362 (N_12362,N_11585,N_11318);
or U12363 (N_12363,N_11021,N_11443);
nor U12364 (N_12364,N_11086,N_11831);
xnor U12365 (N_12365,N_11388,N_11407);
nor U12366 (N_12366,N_10682,N_10769);
xnor U12367 (N_12367,N_10804,N_11145);
nor U12368 (N_12368,N_10782,N_11423);
nand U12369 (N_12369,N_10671,N_11706);
or U12370 (N_12370,N_10778,N_11502);
and U12371 (N_12371,N_10758,N_10594);
or U12372 (N_12372,N_11778,N_11097);
xor U12373 (N_12373,N_10836,N_11590);
and U12374 (N_12374,N_11980,N_11897);
nor U12375 (N_12375,N_10536,N_10748);
nor U12376 (N_12376,N_11302,N_10953);
xnor U12377 (N_12377,N_11460,N_11414);
xnor U12378 (N_12378,N_10668,N_10754);
nand U12379 (N_12379,N_11498,N_11454);
or U12380 (N_12380,N_11240,N_10940);
xor U12381 (N_12381,N_10574,N_10773);
or U12382 (N_12382,N_10793,N_11055);
nor U12383 (N_12383,N_10971,N_11100);
nor U12384 (N_12384,N_11632,N_11307);
nand U12385 (N_12385,N_11329,N_11252);
and U12386 (N_12386,N_11249,N_11769);
or U12387 (N_12387,N_11101,N_11512);
and U12388 (N_12388,N_10652,N_10877);
xnor U12389 (N_12389,N_11202,N_11225);
or U12390 (N_12390,N_11870,N_11583);
nand U12391 (N_12391,N_10968,N_10654);
nand U12392 (N_12392,N_10624,N_11812);
nand U12393 (N_12393,N_10530,N_10952);
xnor U12394 (N_12394,N_10964,N_10732);
or U12395 (N_12395,N_11137,N_11694);
nor U12396 (N_12396,N_10683,N_11428);
nand U12397 (N_12397,N_10937,N_11542);
nand U12398 (N_12398,N_11541,N_11205);
nor U12399 (N_12399,N_10995,N_11555);
xor U12400 (N_12400,N_11756,N_11378);
or U12401 (N_12401,N_11455,N_11154);
or U12402 (N_12402,N_11131,N_10542);
xor U12403 (N_12403,N_11148,N_10801);
or U12404 (N_12404,N_11317,N_11123);
nand U12405 (N_12405,N_11297,N_10664);
xor U12406 (N_12406,N_11096,N_11727);
nor U12407 (N_12407,N_11003,N_11775);
or U12408 (N_12408,N_11478,N_11506);
nor U12409 (N_12409,N_11323,N_11573);
xor U12410 (N_12410,N_10607,N_11890);
and U12411 (N_12411,N_11783,N_11961);
and U12412 (N_12412,N_10893,N_11571);
nor U12413 (N_12413,N_11753,N_11603);
nor U12414 (N_12414,N_11233,N_11303);
nor U12415 (N_12415,N_10723,N_10990);
xor U12416 (N_12416,N_10790,N_11721);
xnor U12417 (N_12417,N_10847,N_10706);
or U12418 (N_12418,N_10961,N_10719);
or U12419 (N_12419,N_10634,N_11410);
xnor U12420 (N_12420,N_10578,N_11854);
nand U12421 (N_12421,N_11963,N_11990);
xor U12422 (N_12422,N_11536,N_11994);
xor U12423 (N_12423,N_11528,N_11674);
nand U12424 (N_12424,N_11545,N_10565);
and U12425 (N_12425,N_10679,N_10962);
or U12426 (N_12426,N_11998,N_11882);
nand U12427 (N_12427,N_10744,N_11290);
or U12428 (N_12428,N_10776,N_10608);
nand U12429 (N_12429,N_11746,N_11757);
xor U12430 (N_12430,N_11187,N_11189);
xor U12431 (N_12431,N_10906,N_11374);
nand U12432 (N_12432,N_10651,N_11733);
nand U12433 (N_12433,N_11183,N_11973);
nor U12434 (N_12434,N_11458,N_10599);
or U12435 (N_12435,N_10658,N_11577);
and U12436 (N_12436,N_10588,N_10859);
nand U12437 (N_12437,N_10858,N_11949);
xor U12438 (N_12438,N_10648,N_11098);
xor U12439 (N_12439,N_11518,N_11231);
or U12440 (N_12440,N_11531,N_11386);
and U12441 (N_12441,N_10838,N_11036);
nand U12442 (N_12442,N_11002,N_10538);
and U12443 (N_12443,N_10617,N_11988);
xor U12444 (N_12444,N_11559,N_11127);
nor U12445 (N_12445,N_10868,N_11232);
xnor U12446 (N_12446,N_11699,N_10888);
xnor U12447 (N_12447,N_10576,N_10571);
xor U12448 (N_12448,N_11763,N_10590);
nand U12449 (N_12449,N_11376,N_11915);
or U12450 (N_12450,N_11091,N_10882);
nor U12451 (N_12451,N_11087,N_10535);
xnor U12452 (N_12452,N_11353,N_11316);
nand U12453 (N_12453,N_10917,N_10825);
and U12454 (N_12454,N_11979,N_11311);
and U12455 (N_12455,N_11281,N_11243);
xor U12456 (N_12456,N_11099,N_11524);
or U12457 (N_12457,N_10622,N_11993);
nand U12458 (N_12458,N_10955,N_11925);
or U12459 (N_12459,N_10819,N_11019);
and U12460 (N_12460,N_10883,N_10640);
nor U12461 (N_12461,N_10746,N_10779);
xnor U12462 (N_12462,N_11853,N_10764);
or U12463 (N_12463,N_10531,N_10885);
nor U12464 (N_12464,N_10676,N_10941);
nand U12465 (N_12465,N_11413,N_10977);
and U12466 (N_12466,N_10645,N_11288);
and U12467 (N_12467,N_10708,N_11477);
or U12468 (N_12468,N_10611,N_11427);
nor U12469 (N_12469,N_11787,N_11735);
or U12470 (N_12470,N_11596,N_11006);
xnor U12471 (N_12471,N_11505,N_11928);
nor U12472 (N_12472,N_11212,N_10606);
or U12473 (N_12473,N_11865,N_11722);
and U12474 (N_12474,N_10693,N_10721);
nor U12475 (N_12475,N_11042,N_11190);
xor U12476 (N_12476,N_10720,N_11838);
or U12477 (N_12477,N_11408,N_10512);
nor U12478 (N_12478,N_11595,N_11813);
and U12479 (N_12479,N_10513,N_10975);
nand U12480 (N_12480,N_10963,N_11332);
and U12481 (N_12481,N_11637,N_11543);
and U12482 (N_12482,N_11434,N_11241);
and U12483 (N_12483,N_11673,N_11070);
and U12484 (N_12484,N_11605,N_10505);
nand U12485 (N_12485,N_10974,N_10890);
or U12486 (N_12486,N_10630,N_11698);
nor U12487 (N_12487,N_11891,N_11550);
xnor U12488 (N_12488,N_11251,N_10519);
and U12489 (N_12489,N_11618,N_10830);
or U12490 (N_12490,N_11429,N_11616);
nor U12491 (N_12491,N_10841,N_11747);
and U12492 (N_12492,N_10559,N_11340);
nand U12493 (N_12493,N_11732,N_11981);
nand U12494 (N_12494,N_11196,N_11686);
nor U12495 (N_12495,N_10691,N_11884);
nor U12496 (N_12496,N_11508,N_10751);
and U12497 (N_12497,N_11447,N_10641);
xor U12498 (N_12498,N_11677,N_11038);
nand U12499 (N_12499,N_11647,N_10696);
nand U12500 (N_12500,N_11941,N_11270);
nand U12501 (N_12501,N_10593,N_11054);
nor U12502 (N_12502,N_11610,N_11640);
nand U12503 (N_12503,N_10735,N_11448);
and U12504 (N_12504,N_11218,N_11314);
nor U12505 (N_12505,N_10982,N_11363);
nand U12506 (N_12506,N_11479,N_10726);
nor U12507 (N_12507,N_11580,N_11264);
and U12508 (N_12508,N_10677,N_11723);
or U12509 (N_12509,N_11959,N_11082);
or U12510 (N_12510,N_11968,N_10700);
nor U12511 (N_12511,N_11011,N_10539);
nor U12512 (N_12512,N_10827,N_11445);
nand U12513 (N_12513,N_11658,N_10983);
xor U12514 (N_12514,N_11700,N_11612);
and U12515 (N_12515,N_11676,N_10585);
nand U12516 (N_12516,N_10524,N_10560);
nor U12517 (N_12517,N_11954,N_11522);
and U12518 (N_12518,N_11065,N_10922);
nor U12519 (N_12519,N_11174,N_11156);
and U12520 (N_12520,N_11802,N_11209);
nor U12521 (N_12521,N_11878,N_11839);
nand U12522 (N_12522,N_11138,N_10712);
and U12523 (N_12523,N_11486,N_10724);
nor U12524 (N_12524,N_11299,N_11304);
xor U12525 (N_12525,N_11553,N_11155);
nand U12526 (N_12526,N_11268,N_11345);
or U12527 (N_12527,N_11383,N_11642);
xor U12528 (N_12528,N_10709,N_10826);
and U12529 (N_12529,N_11327,N_11503);
and U12530 (N_12530,N_10635,N_11237);
nor U12531 (N_12531,N_11837,N_10620);
xor U12532 (N_12532,N_11143,N_11869);
nor U12533 (N_12533,N_10824,N_10752);
nand U12534 (N_12534,N_10784,N_11412);
or U12535 (N_12535,N_11064,N_10876);
nor U12536 (N_12536,N_10689,N_11684);
and U12537 (N_12537,N_11204,N_11080);
xor U12538 (N_12538,N_11768,N_11130);
xnor U12539 (N_12539,N_11725,N_11219);
xnor U12540 (N_12540,N_11653,N_11983);
xnor U12541 (N_12541,N_11507,N_10555);
xnor U12542 (N_12542,N_11628,N_11230);
or U12543 (N_12543,N_11444,N_11440);
and U12544 (N_12544,N_11112,N_10537);
or U12545 (N_12545,N_11452,N_10734);
and U12546 (N_12546,N_10901,N_10857);
nand U12547 (N_12547,N_10928,N_11185);
nand U12548 (N_12548,N_11880,N_11081);
and U12549 (N_12549,N_11352,N_10612);
xnor U12550 (N_12550,N_10520,N_11117);
or U12551 (N_12551,N_11816,N_11788);
xor U12552 (N_12552,N_11690,N_11364);
nor U12553 (N_12553,N_11539,N_11274);
or U12554 (N_12554,N_11514,N_10957);
nor U12555 (N_12555,N_10521,N_11868);
or U12556 (N_12556,N_11075,N_11292);
and U12557 (N_12557,N_11350,N_10655);
nand U12558 (N_12558,N_11351,N_10865);
or U12559 (N_12559,N_11063,N_11828);
and U12560 (N_12560,N_10811,N_11697);
nand U12561 (N_12561,N_10678,N_10909);
or U12562 (N_12562,N_11226,N_11841);
or U12563 (N_12563,N_10742,N_10944);
and U12564 (N_12564,N_11683,N_11617);
nor U12565 (N_12565,N_11134,N_11272);
nand U12566 (N_12566,N_10913,N_11707);
or U12567 (N_12567,N_10946,N_11643);
nor U12568 (N_12568,N_11755,N_11208);
xor U12569 (N_12569,N_11606,N_11121);
and U12570 (N_12570,N_10908,N_11814);
nand U12571 (N_12571,N_11368,N_10737);
and U12572 (N_12572,N_11013,N_10889);
or U12573 (N_12573,N_11348,N_11175);
or U12574 (N_12574,N_11381,N_11696);
nor U12575 (N_12575,N_10813,N_10991);
or U12576 (N_12576,N_11373,N_11554);
xor U12577 (N_12577,N_10948,N_10506);
or U12578 (N_12578,N_11810,N_11754);
xnor U12579 (N_12579,N_10749,N_11051);
or U12580 (N_12580,N_11315,N_11262);
nand U12581 (N_12581,N_10835,N_10969);
or U12582 (N_12582,N_11711,N_10925);
or U12583 (N_12583,N_11069,N_11215);
xor U12584 (N_12584,N_11888,N_11852);
nor U12585 (N_12585,N_11681,N_11883);
xor U12586 (N_12586,N_10529,N_11902);
nand U12587 (N_12587,N_11847,N_11936);
and U12588 (N_12588,N_10915,N_10592);
and U12589 (N_12589,N_11750,N_11211);
nand U12590 (N_12590,N_11709,N_11740);
nor U12591 (N_12591,N_11354,N_11607);
nor U12592 (N_12592,N_11730,N_11043);
and U12593 (N_12593,N_11849,N_10786);
or U12594 (N_12594,N_11083,N_11860);
xor U12595 (N_12595,N_11844,N_10729);
and U12596 (N_12596,N_10562,N_11978);
and U12597 (N_12597,N_10802,N_11343);
and U12598 (N_12598,N_11665,N_10921);
nand U12599 (N_12599,N_11223,N_11856);
or U12600 (N_12600,N_10956,N_10753);
and U12601 (N_12601,N_11191,N_11283);
nor U12602 (N_12602,N_11457,N_11239);
and U12603 (N_12603,N_11338,N_11180);
nand U12604 (N_12604,N_11908,N_11321);
xnor U12605 (N_12605,N_11236,N_11336);
nand U12606 (N_12606,N_10511,N_10927);
nand U12607 (N_12607,N_11105,N_10760);
or U12608 (N_12608,N_10522,N_11574);
or U12609 (N_12609,N_11530,N_11729);
nand U12610 (N_12610,N_11046,N_11962);
nand U12611 (N_12611,N_11220,N_10791);
xnor U12612 (N_12612,N_11551,N_10584);
or U12613 (N_12613,N_11142,N_10626);
nor U12614 (N_12614,N_10500,N_11158);
xor U12615 (N_12615,N_10777,N_11629);
nor U12616 (N_12616,N_11188,N_10716);
or U12617 (N_12617,N_11786,N_11591);
nand U12618 (N_12618,N_10692,N_11951);
nand U12619 (N_12619,N_11370,N_11803);
or U12620 (N_12620,N_11115,N_10950);
and U12621 (N_12621,N_11494,N_10831);
nand U12622 (N_12622,N_11472,N_11651);
nor U12623 (N_12623,N_10628,N_11417);
or U12624 (N_12624,N_11221,N_11609);
xnor U12625 (N_12625,N_10986,N_10725);
xnor U12626 (N_12626,N_10828,N_10853);
xnor U12627 (N_12627,N_11333,N_11045);
and U12628 (N_12628,N_11238,N_11401);
nor U12629 (N_12629,N_10516,N_11881);
or U12630 (N_12630,N_11446,N_11195);
nor U12631 (N_12631,N_11305,N_11873);
or U12632 (N_12632,N_10526,N_10842);
xnor U12633 (N_12633,N_11593,N_11631);
and U12634 (N_12634,N_11149,N_11451);
nand U12635 (N_12635,N_11151,N_11855);
nor U12636 (N_12636,N_10707,N_10698);
or U12637 (N_12637,N_11901,N_11736);
nor U12638 (N_12638,N_10861,N_10704);
and U12639 (N_12639,N_11000,N_11280);
nand U12640 (N_12640,N_11991,N_10549);
or U12641 (N_12641,N_11635,N_10663);
or U12642 (N_12642,N_11471,N_11796);
or U12643 (N_12643,N_10851,N_10650);
nand U12644 (N_12644,N_11668,N_11398);
and U12645 (N_12645,N_11715,N_11906);
nand U12646 (N_12646,N_11935,N_11759);
or U12647 (N_12647,N_11033,N_10509);
xnor U12648 (N_12648,N_11624,N_11833);
nand U12649 (N_12649,N_11228,N_11619);
nand U12650 (N_12650,N_11809,N_11627);
nor U12651 (N_12651,N_10914,N_10589);
xor U12652 (N_12652,N_11377,N_11620);
or U12653 (N_12653,N_10910,N_11805);
and U12654 (N_12654,N_11324,N_11662);
or U12655 (N_12655,N_11527,N_10796);
and U12656 (N_12656,N_11929,N_10815);
nor U12657 (N_12657,N_10685,N_11650);
xnor U12658 (N_12658,N_11153,N_11656);
or U12659 (N_12659,N_11118,N_11210);
nor U12660 (N_12660,N_10656,N_11927);
or U12661 (N_12661,N_11279,N_11488);
or U12662 (N_12662,N_11630,N_11800);
xnor U12663 (N_12663,N_11752,N_11835);
or U12664 (N_12664,N_11742,N_11164);
nand U12665 (N_12665,N_10960,N_11600);
nor U12666 (N_12666,N_11975,N_11967);
nor U12667 (N_12667,N_11424,N_10688);
xnor U12668 (N_12668,N_11076,N_11492);
and U12669 (N_12669,N_10765,N_11242);
or U12670 (N_12670,N_11362,N_11744);
nor U12671 (N_12671,N_11862,N_11942);
and U12672 (N_12672,N_11726,N_11977);
nand U12673 (N_12673,N_10649,N_11235);
or U12674 (N_12674,N_11256,N_11426);
nor U12675 (N_12675,N_11999,N_11565);
xnor U12676 (N_12676,N_11328,N_11114);
nand U12677 (N_12677,N_10999,N_10966);
and U12678 (N_12678,N_10717,N_11416);
xnor U12679 (N_12679,N_11549,N_11431);
nand U12680 (N_12680,N_11436,N_11409);
nor U12681 (N_12681,N_11944,N_10703);
nor U12682 (N_12682,N_10775,N_10756);
xor U12683 (N_12683,N_10701,N_10935);
nand U12684 (N_12684,N_11499,N_11260);
or U12685 (N_12685,N_10976,N_10929);
or U12686 (N_12686,N_11614,N_11300);
and U12687 (N_12687,N_11597,N_11982);
or U12688 (N_12688,N_11258,N_10710);
nor U12689 (N_12689,N_11823,N_10596);
or U12690 (N_12690,N_11713,N_11048);
and U12691 (N_12691,N_11435,N_11771);
xnor U12692 (N_12692,N_11104,N_10586);
and U12693 (N_12693,N_10583,N_10740);
nor U12694 (N_12694,N_11026,N_11657);
nor U12695 (N_12695,N_10867,N_11687);
or U12696 (N_12696,N_11039,N_11406);
nand U12697 (N_12697,N_11289,N_10501);
xnor U12698 (N_12698,N_11464,N_11523);
and U12699 (N_12699,N_11675,N_11894);
nor U12700 (N_12700,N_11014,N_11931);
nor U12701 (N_12701,N_11203,N_11621);
xor U12702 (N_12702,N_10942,N_11633);
xnor U12703 (N_12703,N_11132,N_11484);
nand U12704 (N_12704,N_10792,N_11461);
or U12705 (N_12705,N_11365,N_10517);
xor U12706 (N_12706,N_10747,N_10814);
nor U12707 (N_12707,N_11887,N_11073);
nor U12708 (N_12708,N_11072,N_10514);
xor U12709 (N_12709,N_10934,N_10923);
xor U12710 (N_12710,N_10528,N_11400);
nor U12711 (N_12711,N_10573,N_10755);
nor U12712 (N_12712,N_11785,N_11519);
or U12713 (N_12713,N_11261,N_10911);
nor U12714 (N_12714,N_11380,N_10820);
nor U12715 (N_12715,N_11295,N_11704);
nor U12716 (N_12716,N_11799,N_11418);
xnor U12717 (N_12717,N_11421,N_11996);
xor U12718 (N_12718,N_11126,N_11564);
nand U12719 (N_12719,N_11974,N_10839);
xnor U12720 (N_12720,N_11168,N_11245);
or U12721 (N_12721,N_11133,N_11634);
xnor U12722 (N_12722,N_11433,N_11371);
xor U12723 (N_12723,N_11459,N_11905);
and U12724 (N_12724,N_11520,N_11491);
nor U12725 (N_12725,N_10601,N_10998);
xor U12726 (N_12726,N_11608,N_11387);
or U12727 (N_12727,N_11040,N_11113);
or U12728 (N_12728,N_11820,N_11465);
and U12729 (N_12729,N_10577,N_11020);
nand U12730 (N_12730,N_11679,N_10657);
nor U12731 (N_12731,N_11586,N_11166);
nand U12732 (N_12732,N_11269,N_11649);
and U12733 (N_12733,N_10770,N_10666);
nand U12734 (N_12734,N_10518,N_11030);
nor U12735 (N_12735,N_11509,N_11062);
nand U12736 (N_12736,N_11140,N_10809);
or U12737 (N_12737,N_11566,N_11254);
nand U12738 (N_12738,N_11393,N_11496);
xor U12739 (N_12739,N_10874,N_10643);
xnor U12740 (N_12740,N_10834,N_11748);
nand U12741 (N_12741,N_11485,N_11517);
xnor U12742 (N_12742,N_11875,N_11946);
and U12743 (N_12743,N_11572,N_10845);
xor U12744 (N_12744,N_10978,N_10541);
and U12745 (N_12745,N_11442,N_10880);
nand U12746 (N_12746,N_11007,N_11582);
xor U12747 (N_12747,N_11719,N_11773);
nand U12748 (N_12748,N_11516,N_11116);
nor U12749 (N_12749,N_10898,N_11575);
nand U12750 (N_12750,N_11302,N_10655);
or U12751 (N_12751,N_10844,N_11269);
and U12752 (N_12752,N_11281,N_11913);
and U12753 (N_12753,N_11524,N_11555);
xnor U12754 (N_12754,N_11117,N_10582);
nand U12755 (N_12755,N_10522,N_11390);
nand U12756 (N_12756,N_10768,N_11582);
or U12757 (N_12757,N_10996,N_11918);
nor U12758 (N_12758,N_11455,N_11477);
xor U12759 (N_12759,N_10934,N_11687);
and U12760 (N_12760,N_10674,N_11764);
and U12761 (N_12761,N_11885,N_11399);
nand U12762 (N_12762,N_11306,N_11898);
and U12763 (N_12763,N_11922,N_11387);
nand U12764 (N_12764,N_11354,N_11421);
xnor U12765 (N_12765,N_10624,N_10793);
nand U12766 (N_12766,N_10823,N_11137);
xor U12767 (N_12767,N_11491,N_11249);
or U12768 (N_12768,N_11103,N_10527);
nor U12769 (N_12769,N_11836,N_11263);
and U12770 (N_12770,N_11443,N_11872);
nand U12771 (N_12771,N_11178,N_11938);
nor U12772 (N_12772,N_10586,N_11916);
nor U12773 (N_12773,N_11522,N_11608);
nand U12774 (N_12774,N_11625,N_10938);
and U12775 (N_12775,N_11757,N_11076);
or U12776 (N_12776,N_10543,N_10729);
nor U12777 (N_12777,N_11824,N_10765);
or U12778 (N_12778,N_11962,N_11328);
and U12779 (N_12779,N_11683,N_10681);
and U12780 (N_12780,N_11350,N_11805);
nor U12781 (N_12781,N_10776,N_10964);
nor U12782 (N_12782,N_10553,N_11055);
and U12783 (N_12783,N_10644,N_11375);
nor U12784 (N_12784,N_11114,N_11357);
nor U12785 (N_12785,N_11913,N_11525);
or U12786 (N_12786,N_10694,N_10696);
and U12787 (N_12787,N_11257,N_11861);
or U12788 (N_12788,N_10911,N_11210);
nor U12789 (N_12789,N_10989,N_11083);
nor U12790 (N_12790,N_11561,N_10711);
xnor U12791 (N_12791,N_11159,N_11009);
nand U12792 (N_12792,N_10837,N_10725);
or U12793 (N_12793,N_11978,N_11376);
and U12794 (N_12794,N_11662,N_10706);
nand U12795 (N_12795,N_11779,N_10626);
nor U12796 (N_12796,N_11561,N_11443);
nor U12797 (N_12797,N_11834,N_11004);
xor U12798 (N_12798,N_11504,N_11073);
and U12799 (N_12799,N_10537,N_11170);
nor U12800 (N_12800,N_11984,N_10670);
xor U12801 (N_12801,N_11204,N_11096);
nand U12802 (N_12802,N_10997,N_11321);
nand U12803 (N_12803,N_11441,N_11485);
xor U12804 (N_12804,N_10829,N_11884);
xor U12805 (N_12805,N_11297,N_10902);
nand U12806 (N_12806,N_11646,N_11799);
or U12807 (N_12807,N_11252,N_11985);
nand U12808 (N_12808,N_11544,N_10921);
xnor U12809 (N_12809,N_11302,N_11884);
and U12810 (N_12810,N_11298,N_11312);
nand U12811 (N_12811,N_10720,N_11416);
and U12812 (N_12812,N_11719,N_11223);
xnor U12813 (N_12813,N_10553,N_11778);
nand U12814 (N_12814,N_11980,N_11877);
and U12815 (N_12815,N_10503,N_11995);
and U12816 (N_12816,N_11721,N_11339);
xnor U12817 (N_12817,N_11381,N_10712);
nand U12818 (N_12818,N_11780,N_10787);
xnor U12819 (N_12819,N_10907,N_11759);
and U12820 (N_12820,N_11322,N_10580);
and U12821 (N_12821,N_11486,N_11520);
or U12822 (N_12822,N_11701,N_10944);
nand U12823 (N_12823,N_10763,N_10813);
or U12824 (N_12824,N_11049,N_11779);
nand U12825 (N_12825,N_10979,N_10998);
or U12826 (N_12826,N_11723,N_10514);
and U12827 (N_12827,N_11151,N_10586);
xnor U12828 (N_12828,N_10729,N_11816);
or U12829 (N_12829,N_11943,N_10743);
nand U12830 (N_12830,N_11694,N_11416);
nand U12831 (N_12831,N_10868,N_11513);
or U12832 (N_12832,N_11138,N_11101);
nand U12833 (N_12833,N_11770,N_10515);
nor U12834 (N_12834,N_11064,N_10513);
nor U12835 (N_12835,N_11849,N_11471);
nand U12836 (N_12836,N_10501,N_11506);
and U12837 (N_12837,N_10734,N_11456);
and U12838 (N_12838,N_11061,N_10644);
xnor U12839 (N_12839,N_11782,N_11694);
or U12840 (N_12840,N_11830,N_10678);
nor U12841 (N_12841,N_10804,N_11687);
nor U12842 (N_12842,N_11985,N_10610);
or U12843 (N_12843,N_10773,N_11452);
nor U12844 (N_12844,N_11515,N_10540);
and U12845 (N_12845,N_11673,N_10851);
nand U12846 (N_12846,N_10699,N_11303);
xor U12847 (N_12847,N_11477,N_11537);
and U12848 (N_12848,N_11949,N_11321);
nand U12849 (N_12849,N_11264,N_10653);
xnor U12850 (N_12850,N_11880,N_11995);
nand U12851 (N_12851,N_11750,N_11820);
xnor U12852 (N_12852,N_11757,N_10519);
or U12853 (N_12853,N_11784,N_11111);
or U12854 (N_12854,N_11375,N_11022);
and U12855 (N_12855,N_11857,N_11602);
xnor U12856 (N_12856,N_11301,N_11093);
nand U12857 (N_12857,N_10573,N_10864);
nand U12858 (N_12858,N_11541,N_10951);
nand U12859 (N_12859,N_11455,N_10649);
nand U12860 (N_12860,N_11092,N_10838);
nor U12861 (N_12861,N_11121,N_11198);
and U12862 (N_12862,N_11092,N_10716);
and U12863 (N_12863,N_10660,N_11445);
xnor U12864 (N_12864,N_11330,N_11152);
nor U12865 (N_12865,N_11578,N_10702);
nand U12866 (N_12866,N_11611,N_11211);
xnor U12867 (N_12867,N_10962,N_11969);
or U12868 (N_12868,N_10780,N_11402);
nand U12869 (N_12869,N_11507,N_10515);
and U12870 (N_12870,N_11462,N_10539);
nand U12871 (N_12871,N_11891,N_11869);
xnor U12872 (N_12872,N_11814,N_10920);
nor U12873 (N_12873,N_11833,N_10540);
or U12874 (N_12874,N_11616,N_10743);
or U12875 (N_12875,N_11883,N_10554);
or U12876 (N_12876,N_11501,N_11195);
nand U12877 (N_12877,N_10769,N_11411);
xor U12878 (N_12878,N_11029,N_11275);
nor U12879 (N_12879,N_11160,N_11742);
xor U12880 (N_12880,N_10623,N_10897);
and U12881 (N_12881,N_11162,N_11673);
or U12882 (N_12882,N_11501,N_11860);
nor U12883 (N_12883,N_10565,N_10604);
or U12884 (N_12884,N_11855,N_11552);
nand U12885 (N_12885,N_10785,N_10764);
nand U12886 (N_12886,N_11685,N_11208);
nand U12887 (N_12887,N_11220,N_11800);
nor U12888 (N_12888,N_11036,N_11524);
and U12889 (N_12889,N_10600,N_11927);
nor U12890 (N_12890,N_10680,N_11104);
nor U12891 (N_12891,N_11773,N_11178);
nor U12892 (N_12892,N_10904,N_11076);
xnor U12893 (N_12893,N_10686,N_11942);
and U12894 (N_12894,N_11861,N_11699);
xor U12895 (N_12895,N_11289,N_11093);
nand U12896 (N_12896,N_11694,N_11082);
xnor U12897 (N_12897,N_11931,N_11527);
nand U12898 (N_12898,N_11871,N_11479);
and U12899 (N_12899,N_11964,N_11990);
nand U12900 (N_12900,N_10831,N_11995);
xnor U12901 (N_12901,N_11381,N_11626);
and U12902 (N_12902,N_11958,N_10714);
and U12903 (N_12903,N_10566,N_11433);
or U12904 (N_12904,N_10748,N_11509);
and U12905 (N_12905,N_11115,N_11533);
nor U12906 (N_12906,N_11040,N_11082);
xnor U12907 (N_12907,N_10763,N_11536);
nor U12908 (N_12908,N_10823,N_11197);
or U12909 (N_12909,N_11801,N_10727);
or U12910 (N_12910,N_11750,N_11059);
nor U12911 (N_12911,N_11764,N_11708);
or U12912 (N_12912,N_11767,N_11873);
nand U12913 (N_12913,N_11204,N_10784);
xnor U12914 (N_12914,N_11904,N_11171);
nand U12915 (N_12915,N_10884,N_10801);
nor U12916 (N_12916,N_10850,N_10867);
nor U12917 (N_12917,N_10555,N_10582);
nor U12918 (N_12918,N_11178,N_10677);
xor U12919 (N_12919,N_11697,N_11090);
and U12920 (N_12920,N_11961,N_11780);
or U12921 (N_12921,N_11486,N_11424);
nand U12922 (N_12922,N_10685,N_10963);
nor U12923 (N_12923,N_11049,N_11767);
nand U12924 (N_12924,N_11086,N_10705);
nand U12925 (N_12925,N_11575,N_11175);
and U12926 (N_12926,N_11210,N_11231);
xnor U12927 (N_12927,N_10937,N_10898);
nand U12928 (N_12928,N_10995,N_10960);
nor U12929 (N_12929,N_10786,N_10654);
and U12930 (N_12930,N_10502,N_10724);
and U12931 (N_12931,N_11471,N_11992);
or U12932 (N_12932,N_11894,N_10771);
nand U12933 (N_12933,N_11757,N_11595);
xnor U12934 (N_12934,N_11479,N_11272);
nor U12935 (N_12935,N_10874,N_11078);
nand U12936 (N_12936,N_11434,N_10618);
nand U12937 (N_12937,N_11392,N_10665);
and U12938 (N_12938,N_11377,N_10997);
nand U12939 (N_12939,N_11532,N_11838);
and U12940 (N_12940,N_11743,N_11092);
nor U12941 (N_12941,N_11563,N_10826);
nand U12942 (N_12942,N_11905,N_10873);
or U12943 (N_12943,N_10518,N_11198);
xnor U12944 (N_12944,N_11264,N_11529);
nor U12945 (N_12945,N_11592,N_11987);
nor U12946 (N_12946,N_11925,N_11719);
nor U12947 (N_12947,N_11562,N_11440);
or U12948 (N_12948,N_11999,N_11794);
or U12949 (N_12949,N_11590,N_11068);
or U12950 (N_12950,N_11963,N_11729);
nand U12951 (N_12951,N_11801,N_11539);
nand U12952 (N_12952,N_11576,N_11593);
or U12953 (N_12953,N_11671,N_11455);
nand U12954 (N_12954,N_11793,N_11521);
and U12955 (N_12955,N_11974,N_11318);
nand U12956 (N_12956,N_11930,N_11834);
nand U12957 (N_12957,N_10587,N_10832);
xor U12958 (N_12958,N_11715,N_11168);
nor U12959 (N_12959,N_11917,N_10795);
and U12960 (N_12960,N_11516,N_11885);
xor U12961 (N_12961,N_10999,N_10926);
and U12962 (N_12962,N_10609,N_11429);
or U12963 (N_12963,N_10793,N_10913);
nand U12964 (N_12964,N_11710,N_11278);
and U12965 (N_12965,N_10650,N_10528);
or U12966 (N_12966,N_10500,N_10618);
nor U12967 (N_12967,N_10580,N_11248);
or U12968 (N_12968,N_11196,N_10868);
xnor U12969 (N_12969,N_11191,N_11342);
nor U12970 (N_12970,N_11026,N_11020);
or U12971 (N_12971,N_11110,N_10879);
nor U12972 (N_12972,N_10843,N_11785);
xnor U12973 (N_12973,N_10504,N_11201);
xor U12974 (N_12974,N_10734,N_11619);
or U12975 (N_12975,N_10847,N_11943);
and U12976 (N_12976,N_10817,N_11549);
nand U12977 (N_12977,N_11072,N_11428);
and U12978 (N_12978,N_11238,N_11359);
and U12979 (N_12979,N_11223,N_10791);
xor U12980 (N_12980,N_10674,N_11024);
nor U12981 (N_12981,N_11961,N_11953);
and U12982 (N_12982,N_11887,N_10680);
and U12983 (N_12983,N_11141,N_11108);
and U12984 (N_12984,N_11138,N_11584);
nand U12985 (N_12985,N_11982,N_10900);
and U12986 (N_12986,N_11805,N_11881);
nand U12987 (N_12987,N_11425,N_11675);
and U12988 (N_12988,N_11795,N_11438);
and U12989 (N_12989,N_10803,N_11711);
nor U12990 (N_12990,N_10738,N_11151);
nor U12991 (N_12991,N_11024,N_11831);
nor U12992 (N_12992,N_11990,N_11425);
or U12993 (N_12993,N_11372,N_11252);
and U12994 (N_12994,N_11251,N_11057);
xor U12995 (N_12995,N_11489,N_11963);
xnor U12996 (N_12996,N_11698,N_10703);
xor U12997 (N_12997,N_11028,N_11758);
nand U12998 (N_12998,N_11798,N_10918);
and U12999 (N_12999,N_10814,N_11588);
xor U13000 (N_13000,N_11409,N_11552);
and U13001 (N_13001,N_11360,N_10572);
or U13002 (N_13002,N_11291,N_10617);
and U13003 (N_13003,N_11270,N_11700);
nor U13004 (N_13004,N_11277,N_11909);
nor U13005 (N_13005,N_11512,N_11258);
nand U13006 (N_13006,N_11864,N_10505);
xnor U13007 (N_13007,N_11435,N_11600);
or U13008 (N_13008,N_10674,N_10898);
and U13009 (N_13009,N_10507,N_11917);
nor U13010 (N_13010,N_11934,N_11130);
nand U13011 (N_13011,N_11695,N_10648);
xnor U13012 (N_13012,N_10972,N_11933);
xor U13013 (N_13013,N_10858,N_11628);
nor U13014 (N_13014,N_11300,N_11651);
nand U13015 (N_13015,N_11783,N_11079);
nor U13016 (N_13016,N_11630,N_10880);
xor U13017 (N_13017,N_11656,N_11860);
xnor U13018 (N_13018,N_11575,N_11726);
and U13019 (N_13019,N_11337,N_10560);
xnor U13020 (N_13020,N_11464,N_11558);
or U13021 (N_13021,N_11866,N_11651);
xor U13022 (N_13022,N_11648,N_11818);
or U13023 (N_13023,N_11674,N_10636);
xor U13024 (N_13024,N_11702,N_10952);
and U13025 (N_13025,N_10987,N_11661);
nand U13026 (N_13026,N_10710,N_11712);
nor U13027 (N_13027,N_11412,N_11131);
and U13028 (N_13028,N_11140,N_11172);
nor U13029 (N_13029,N_10770,N_11589);
nor U13030 (N_13030,N_11817,N_11250);
or U13031 (N_13031,N_11166,N_11045);
and U13032 (N_13032,N_10702,N_10989);
or U13033 (N_13033,N_11425,N_10990);
xnor U13034 (N_13034,N_10694,N_11703);
nor U13035 (N_13035,N_11160,N_10679);
nor U13036 (N_13036,N_11231,N_10733);
xnor U13037 (N_13037,N_11695,N_10642);
nand U13038 (N_13038,N_10635,N_11859);
nand U13039 (N_13039,N_11386,N_11996);
nand U13040 (N_13040,N_11285,N_11298);
xor U13041 (N_13041,N_11148,N_11548);
nor U13042 (N_13042,N_11059,N_11936);
nand U13043 (N_13043,N_11628,N_11161);
nor U13044 (N_13044,N_11353,N_11712);
and U13045 (N_13045,N_11828,N_11818);
xnor U13046 (N_13046,N_11301,N_10632);
nor U13047 (N_13047,N_11167,N_10805);
xor U13048 (N_13048,N_11538,N_11822);
or U13049 (N_13049,N_10993,N_11813);
and U13050 (N_13050,N_10686,N_11534);
or U13051 (N_13051,N_11940,N_10641);
or U13052 (N_13052,N_11110,N_11315);
nor U13053 (N_13053,N_11633,N_10893);
xor U13054 (N_13054,N_11737,N_11360);
xnor U13055 (N_13055,N_11581,N_11549);
or U13056 (N_13056,N_11837,N_11568);
nor U13057 (N_13057,N_11623,N_11166);
nand U13058 (N_13058,N_11973,N_10519);
nand U13059 (N_13059,N_11528,N_11050);
or U13060 (N_13060,N_11337,N_11343);
nand U13061 (N_13061,N_10872,N_11798);
xnor U13062 (N_13062,N_10511,N_11077);
nor U13063 (N_13063,N_11742,N_10528);
and U13064 (N_13064,N_11211,N_11422);
nand U13065 (N_13065,N_10704,N_11573);
xor U13066 (N_13066,N_11717,N_10720);
and U13067 (N_13067,N_10708,N_10928);
and U13068 (N_13068,N_11114,N_10627);
xnor U13069 (N_13069,N_11613,N_11577);
and U13070 (N_13070,N_11379,N_10597);
or U13071 (N_13071,N_10853,N_11752);
nand U13072 (N_13072,N_10879,N_11516);
and U13073 (N_13073,N_10854,N_11694);
nor U13074 (N_13074,N_11976,N_11255);
and U13075 (N_13075,N_11718,N_11701);
nand U13076 (N_13076,N_11282,N_11790);
nand U13077 (N_13077,N_11600,N_10891);
xor U13078 (N_13078,N_11968,N_11932);
and U13079 (N_13079,N_10832,N_10511);
nand U13080 (N_13080,N_11159,N_11471);
nor U13081 (N_13081,N_11237,N_11715);
nand U13082 (N_13082,N_11515,N_10678);
nand U13083 (N_13083,N_11728,N_11758);
nand U13084 (N_13084,N_11545,N_11986);
nand U13085 (N_13085,N_11378,N_11666);
nor U13086 (N_13086,N_11628,N_11859);
nor U13087 (N_13087,N_11135,N_11334);
or U13088 (N_13088,N_10697,N_11961);
nor U13089 (N_13089,N_11519,N_10969);
xor U13090 (N_13090,N_10656,N_10732);
or U13091 (N_13091,N_10961,N_11425);
nor U13092 (N_13092,N_10646,N_10578);
xnor U13093 (N_13093,N_11572,N_11517);
nand U13094 (N_13094,N_10914,N_10972);
and U13095 (N_13095,N_11216,N_11858);
or U13096 (N_13096,N_11367,N_11801);
and U13097 (N_13097,N_10622,N_11428);
nand U13098 (N_13098,N_11637,N_10746);
xor U13099 (N_13099,N_10699,N_11089);
xor U13100 (N_13100,N_10843,N_11094);
xnor U13101 (N_13101,N_10834,N_11095);
or U13102 (N_13102,N_11284,N_11977);
nand U13103 (N_13103,N_11902,N_10798);
or U13104 (N_13104,N_10584,N_11265);
nand U13105 (N_13105,N_11669,N_11672);
xor U13106 (N_13106,N_11725,N_11856);
xor U13107 (N_13107,N_11473,N_11943);
or U13108 (N_13108,N_10743,N_11418);
or U13109 (N_13109,N_10635,N_10702);
xor U13110 (N_13110,N_10804,N_11736);
nor U13111 (N_13111,N_11454,N_11720);
and U13112 (N_13112,N_11465,N_10550);
and U13113 (N_13113,N_11494,N_10617);
or U13114 (N_13114,N_11453,N_11390);
nand U13115 (N_13115,N_11760,N_11509);
and U13116 (N_13116,N_11692,N_11907);
and U13117 (N_13117,N_11213,N_11737);
xnor U13118 (N_13118,N_10515,N_10944);
and U13119 (N_13119,N_10694,N_11851);
xor U13120 (N_13120,N_11814,N_10959);
xnor U13121 (N_13121,N_11456,N_10826);
or U13122 (N_13122,N_11430,N_10841);
nor U13123 (N_13123,N_10855,N_11187);
and U13124 (N_13124,N_11641,N_11006);
nor U13125 (N_13125,N_10814,N_11467);
nand U13126 (N_13126,N_10608,N_10795);
or U13127 (N_13127,N_11787,N_10599);
and U13128 (N_13128,N_10668,N_11394);
nor U13129 (N_13129,N_10834,N_11368);
nand U13130 (N_13130,N_10676,N_11478);
or U13131 (N_13131,N_11453,N_10574);
and U13132 (N_13132,N_11018,N_11830);
nor U13133 (N_13133,N_11277,N_10910);
nor U13134 (N_13134,N_10706,N_11576);
nand U13135 (N_13135,N_10655,N_11380);
xor U13136 (N_13136,N_10919,N_10561);
and U13137 (N_13137,N_11338,N_11299);
nand U13138 (N_13138,N_10805,N_10556);
xor U13139 (N_13139,N_10765,N_10866);
nand U13140 (N_13140,N_10845,N_11125);
xor U13141 (N_13141,N_10886,N_11677);
nand U13142 (N_13142,N_11082,N_11607);
nor U13143 (N_13143,N_11496,N_11751);
nand U13144 (N_13144,N_10741,N_11805);
and U13145 (N_13145,N_11662,N_10895);
xor U13146 (N_13146,N_11916,N_10844);
xnor U13147 (N_13147,N_10636,N_11776);
nor U13148 (N_13148,N_11661,N_11379);
or U13149 (N_13149,N_10783,N_11434);
nand U13150 (N_13150,N_11700,N_11734);
nor U13151 (N_13151,N_10935,N_10622);
nand U13152 (N_13152,N_10613,N_11740);
xor U13153 (N_13153,N_11291,N_10661);
nand U13154 (N_13154,N_11507,N_11310);
nand U13155 (N_13155,N_10861,N_11489);
and U13156 (N_13156,N_10863,N_11604);
xor U13157 (N_13157,N_11154,N_10930);
xor U13158 (N_13158,N_11136,N_10784);
xor U13159 (N_13159,N_10599,N_11057);
nor U13160 (N_13160,N_11632,N_11970);
and U13161 (N_13161,N_10520,N_10529);
nor U13162 (N_13162,N_10904,N_11835);
or U13163 (N_13163,N_11778,N_11390);
xor U13164 (N_13164,N_11996,N_10951);
xnor U13165 (N_13165,N_11677,N_10500);
nand U13166 (N_13166,N_11566,N_11690);
or U13167 (N_13167,N_11359,N_10711);
or U13168 (N_13168,N_11640,N_11635);
xor U13169 (N_13169,N_11265,N_11717);
xor U13170 (N_13170,N_11921,N_10896);
nor U13171 (N_13171,N_11595,N_10652);
and U13172 (N_13172,N_11284,N_11309);
xnor U13173 (N_13173,N_11081,N_11157);
xor U13174 (N_13174,N_11684,N_10929);
xnor U13175 (N_13175,N_10529,N_11059);
nand U13176 (N_13176,N_11686,N_11667);
or U13177 (N_13177,N_10978,N_11793);
nand U13178 (N_13178,N_10623,N_11926);
nor U13179 (N_13179,N_11727,N_10962);
and U13180 (N_13180,N_10836,N_11968);
xnor U13181 (N_13181,N_11958,N_11919);
or U13182 (N_13182,N_11533,N_10801);
nor U13183 (N_13183,N_10895,N_10770);
nand U13184 (N_13184,N_11674,N_10693);
or U13185 (N_13185,N_10524,N_11567);
nor U13186 (N_13186,N_10902,N_11304);
and U13187 (N_13187,N_10945,N_11752);
xnor U13188 (N_13188,N_11858,N_11469);
or U13189 (N_13189,N_11189,N_11420);
xnor U13190 (N_13190,N_10538,N_11377);
xnor U13191 (N_13191,N_11782,N_11362);
and U13192 (N_13192,N_11140,N_11070);
xor U13193 (N_13193,N_11610,N_11766);
and U13194 (N_13194,N_11446,N_11255);
xnor U13195 (N_13195,N_11444,N_10994);
xnor U13196 (N_13196,N_10621,N_10729);
xor U13197 (N_13197,N_11698,N_11968);
nor U13198 (N_13198,N_11421,N_10851);
and U13199 (N_13199,N_11741,N_11860);
xnor U13200 (N_13200,N_10512,N_10647);
or U13201 (N_13201,N_10679,N_11408);
nand U13202 (N_13202,N_11098,N_11862);
nand U13203 (N_13203,N_11274,N_11562);
and U13204 (N_13204,N_10792,N_11951);
or U13205 (N_13205,N_11646,N_11116);
xnor U13206 (N_13206,N_11072,N_11304);
nor U13207 (N_13207,N_11326,N_10967);
nand U13208 (N_13208,N_10550,N_10885);
xor U13209 (N_13209,N_11833,N_11768);
nor U13210 (N_13210,N_11340,N_11985);
or U13211 (N_13211,N_10689,N_10775);
or U13212 (N_13212,N_11517,N_10974);
and U13213 (N_13213,N_11594,N_10628);
nor U13214 (N_13214,N_11027,N_11835);
nor U13215 (N_13215,N_11190,N_11990);
or U13216 (N_13216,N_10969,N_11310);
and U13217 (N_13217,N_11218,N_11736);
or U13218 (N_13218,N_11419,N_11528);
nand U13219 (N_13219,N_11325,N_11100);
and U13220 (N_13220,N_10675,N_10988);
and U13221 (N_13221,N_11062,N_11550);
xnor U13222 (N_13222,N_11203,N_11660);
or U13223 (N_13223,N_10768,N_11871);
nand U13224 (N_13224,N_11601,N_10691);
and U13225 (N_13225,N_10809,N_11385);
xor U13226 (N_13226,N_11188,N_11272);
xor U13227 (N_13227,N_11419,N_11828);
or U13228 (N_13228,N_10567,N_10699);
or U13229 (N_13229,N_11561,N_11273);
or U13230 (N_13230,N_11482,N_11225);
nand U13231 (N_13231,N_11295,N_11495);
nand U13232 (N_13232,N_11764,N_11499);
nand U13233 (N_13233,N_10926,N_11343);
nor U13234 (N_13234,N_11405,N_10614);
xor U13235 (N_13235,N_11488,N_10694);
or U13236 (N_13236,N_11938,N_11114);
or U13237 (N_13237,N_11704,N_11454);
nand U13238 (N_13238,N_10899,N_11995);
and U13239 (N_13239,N_11795,N_11835);
nor U13240 (N_13240,N_10745,N_10824);
nand U13241 (N_13241,N_11608,N_11397);
or U13242 (N_13242,N_11835,N_10748);
nor U13243 (N_13243,N_11642,N_11615);
nand U13244 (N_13244,N_11853,N_11757);
nand U13245 (N_13245,N_10611,N_11030);
and U13246 (N_13246,N_10891,N_11421);
nor U13247 (N_13247,N_11713,N_11118);
nor U13248 (N_13248,N_10789,N_11337);
nor U13249 (N_13249,N_10954,N_11681);
nand U13250 (N_13250,N_11471,N_10702);
or U13251 (N_13251,N_11570,N_10594);
xnor U13252 (N_13252,N_11649,N_11505);
nor U13253 (N_13253,N_10647,N_10681);
or U13254 (N_13254,N_11002,N_11183);
nor U13255 (N_13255,N_10643,N_11232);
nor U13256 (N_13256,N_11860,N_11369);
and U13257 (N_13257,N_11782,N_10528);
nand U13258 (N_13258,N_11082,N_10820);
xor U13259 (N_13259,N_11966,N_11524);
and U13260 (N_13260,N_11484,N_10556);
xnor U13261 (N_13261,N_10968,N_10845);
and U13262 (N_13262,N_11784,N_11480);
nand U13263 (N_13263,N_11359,N_10912);
nor U13264 (N_13264,N_10735,N_10513);
xor U13265 (N_13265,N_11971,N_11739);
and U13266 (N_13266,N_11704,N_11332);
and U13267 (N_13267,N_10716,N_11485);
nand U13268 (N_13268,N_11149,N_11318);
or U13269 (N_13269,N_11098,N_11083);
xnor U13270 (N_13270,N_11446,N_11186);
or U13271 (N_13271,N_11294,N_10705);
or U13272 (N_13272,N_11274,N_10664);
xnor U13273 (N_13273,N_10711,N_10769);
or U13274 (N_13274,N_11689,N_11969);
xor U13275 (N_13275,N_10797,N_11403);
nor U13276 (N_13276,N_11834,N_11827);
and U13277 (N_13277,N_10870,N_11796);
or U13278 (N_13278,N_11837,N_11889);
nand U13279 (N_13279,N_11882,N_10966);
or U13280 (N_13280,N_10728,N_11500);
nor U13281 (N_13281,N_11098,N_10686);
or U13282 (N_13282,N_11087,N_11459);
nor U13283 (N_13283,N_10895,N_10919);
and U13284 (N_13284,N_11705,N_10859);
and U13285 (N_13285,N_11124,N_10984);
or U13286 (N_13286,N_11395,N_11546);
xnor U13287 (N_13287,N_11459,N_11467);
and U13288 (N_13288,N_11211,N_11007);
xnor U13289 (N_13289,N_10892,N_10939);
and U13290 (N_13290,N_10538,N_10736);
and U13291 (N_13291,N_11963,N_11076);
xor U13292 (N_13292,N_11310,N_11689);
or U13293 (N_13293,N_11688,N_11417);
and U13294 (N_13294,N_11030,N_10808);
xor U13295 (N_13295,N_11398,N_11682);
xnor U13296 (N_13296,N_11089,N_10952);
nand U13297 (N_13297,N_11026,N_11932);
and U13298 (N_13298,N_11533,N_11380);
and U13299 (N_13299,N_10953,N_10536);
and U13300 (N_13300,N_11211,N_11296);
and U13301 (N_13301,N_10931,N_10531);
xor U13302 (N_13302,N_10722,N_11081);
nand U13303 (N_13303,N_11680,N_11078);
or U13304 (N_13304,N_10943,N_11185);
and U13305 (N_13305,N_11956,N_10586);
xnor U13306 (N_13306,N_10929,N_11008);
nand U13307 (N_13307,N_10541,N_11354);
nand U13308 (N_13308,N_10661,N_11648);
nand U13309 (N_13309,N_10510,N_10943);
nor U13310 (N_13310,N_10884,N_10636);
or U13311 (N_13311,N_10857,N_11517);
or U13312 (N_13312,N_11588,N_11784);
nor U13313 (N_13313,N_11321,N_11497);
or U13314 (N_13314,N_11327,N_11158);
nor U13315 (N_13315,N_11763,N_10844);
nor U13316 (N_13316,N_11784,N_11119);
nand U13317 (N_13317,N_10629,N_10977);
xnor U13318 (N_13318,N_11661,N_11304);
and U13319 (N_13319,N_11038,N_11970);
xnor U13320 (N_13320,N_11551,N_10899);
or U13321 (N_13321,N_11764,N_11671);
or U13322 (N_13322,N_10703,N_10848);
xnor U13323 (N_13323,N_10744,N_11258);
and U13324 (N_13324,N_11324,N_11738);
or U13325 (N_13325,N_10887,N_10795);
and U13326 (N_13326,N_10776,N_11943);
and U13327 (N_13327,N_11788,N_11920);
or U13328 (N_13328,N_11701,N_11282);
nand U13329 (N_13329,N_11307,N_11347);
xor U13330 (N_13330,N_10571,N_11524);
xor U13331 (N_13331,N_11536,N_11581);
and U13332 (N_13332,N_11720,N_11976);
nand U13333 (N_13333,N_11177,N_11805);
nand U13334 (N_13334,N_11976,N_11431);
and U13335 (N_13335,N_10621,N_10956);
or U13336 (N_13336,N_11953,N_11337);
and U13337 (N_13337,N_11615,N_11257);
and U13338 (N_13338,N_11364,N_10994);
nor U13339 (N_13339,N_11982,N_10830);
and U13340 (N_13340,N_11766,N_10535);
and U13341 (N_13341,N_10701,N_11683);
nand U13342 (N_13342,N_10930,N_11335);
or U13343 (N_13343,N_11389,N_11231);
nor U13344 (N_13344,N_11306,N_11273);
xor U13345 (N_13345,N_11997,N_11200);
nand U13346 (N_13346,N_11764,N_11453);
and U13347 (N_13347,N_11051,N_11020);
xor U13348 (N_13348,N_11127,N_11667);
and U13349 (N_13349,N_11351,N_11646);
or U13350 (N_13350,N_11974,N_11068);
xnor U13351 (N_13351,N_11125,N_11116);
or U13352 (N_13352,N_11648,N_11133);
and U13353 (N_13353,N_11508,N_11766);
and U13354 (N_13354,N_11078,N_11941);
or U13355 (N_13355,N_11886,N_11273);
and U13356 (N_13356,N_11005,N_11392);
nor U13357 (N_13357,N_10859,N_11718);
nor U13358 (N_13358,N_11952,N_11823);
or U13359 (N_13359,N_10882,N_11977);
nor U13360 (N_13360,N_11802,N_11696);
nor U13361 (N_13361,N_10701,N_11224);
xor U13362 (N_13362,N_11278,N_10931);
xnor U13363 (N_13363,N_10811,N_11418);
nand U13364 (N_13364,N_11051,N_11992);
nand U13365 (N_13365,N_10799,N_11047);
or U13366 (N_13366,N_11975,N_11197);
nand U13367 (N_13367,N_10557,N_11551);
xor U13368 (N_13368,N_11235,N_11870);
xnor U13369 (N_13369,N_11866,N_10529);
and U13370 (N_13370,N_11554,N_11958);
nand U13371 (N_13371,N_11889,N_10628);
xnor U13372 (N_13372,N_11275,N_11472);
nand U13373 (N_13373,N_10995,N_11113);
or U13374 (N_13374,N_10552,N_11756);
xor U13375 (N_13375,N_11571,N_10531);
xnor U13376 (N_13376,N_11816,N_11061);
or U13377 (N_13377,N_11413,N_11646);
nand U13378 (N_13378,N_10986,N_10902);
nor U13379 (N_13379,N_11926,N_11614);
nor U13380 (N_13380,N_11445,N_10797);
nand U13381 (N_13381,N_11057,N_10773);
xor U13382 (N_13382,N_11475,N_10920);
or U13383 (N_13383,N_11568,N_11448);
or U13384 (N_13384,N_10559,N_10712);
nand U13385 (N_13385,N_10535,N_11946);
and U13386 (N_13386,N_11597,N_11572);
xor U13387 (N_13387,N_11785,N_11498);
or U13388 (N_13388,N_11027,N_11661);
nand U13389 (N_13389,N_11076,N_11118);
xnor U13390 (N_13390,N_11236,N_11767);
nand U13391 (N_13391,N_11181,N_11404);
nand U13392 (N_13392,N_11040,N_11429);
and U13393 (N_13393,N_10804,N_11156);
or U13394 (N_13394,N_11043,N_11720);
xor U13395 (N_13395,N_10767,N_11792);
nand U13396 (N_13396,N_10694,N_11334);
and U13397 (N_13397,N_10544,N_11746);
nor U13398 (N_13398,N_11947,N_11352);
xnor U13399 (N_13399,N_10838,N_11965);
nor U13400 (N_13400,N_11958,N_10750);
xnor U13401 (N_13401,N_10581,N_11518);
and U13402 (N_13402,N_11163,N_11520);
nor U13403 (N_13403,N_11062,N_10731);
or U13404 (N_13404,N_11146,N_10540);
or U13405 (N_13405,N_11955,N_11195);
or U13406 (N_13406,N_11411,N_11466);
or U13407 (N_13407,N_11088,N_10610);
and U13408 (N_13408,N_11268,N_10686);
nor U13409 (N_13409,N_11291,N_10757);
xor U13410 (N_13410,N_10911,N_10826);
xnor U13411 (N_13411,N_11853,N_10722);
xnor U13412 (N_13412,N_11201,N_10714);
or U13413 (N_13413,N_11643,N_10854);
and U13414 (N_13414,N_11406,N_11405);
nor U13415 (N_13415,N_11185,N_11913);
xor U13416 (N_13416,N_11126,N_11859);
and U13417 (N_13417,N_10993,N_11822);
nand U13418 (N_13418,N_11928,N_10820);
nand U13419 (N_13419,N_11790,N_10692);
nor U13420 (N_13420,N_11311,N_10604);
or U13421 (N_13421,N_11276,N_11260);
nand U13422 (N_13422,N_10560,N_10606);
or U13423 (N_13423,N_10952,N_11026);
nand U13424 (N_13424,N_10544,N_11433);
or U13425 (N_13425,N_10886,N_11188);
nor U13426 (N_13426,N_11909,N_11897);
nor U13427 (N_13427,N_11279,N_11140);
nand U13428 (N_13428,N_10504,N_11925);
nand U13429 (N_13429,N_10747,N_11647);
nand U13430 (N_13430,N_11315,N_11038);
nand U13431 (N_13431,N_11203,N_10928);
nand U13432 (N_13432,N_11335,N_10996);
or U13433 (N_13433,N_11789,N_11729);
or U13434 (N_13434,N_11416,N_10799);
nand U13435 (N_13435,N_10697,N_11466);
nor U13436 (N_13436,N_10696,N_11964);
nor U13437 (N_13437,N_10817,N_10675);
nor U13438 (N_13438,N_11113,N_11168);
or U13439 (N_13439,N_11262,N_11316);
or U13440 (N_13440,N_11176,N_11055);
xor U13441 (N_13441,N_10946,N_10882);
nand U13442 (N_13442,N_11113,N_10562);
or U13443 (N_13443,N_10856,N_10920);
xnor U13444 (N_13444,N_11376,N_10920);
xor U13445 (N_13445,N_10776,N_10944);
xor U13446 (N_13446,N_11417,N_10809);
nand U13447 (N_13447,N_11949,N_11312);
nand U13448 (N_13448,N_10741,N_10939);
or U13449 (N_13449,N_10567,N_11594);
xor U13450 (N_13450,N_11765,N_10980);
and U13451 (N_13451,N_11438,N_10730);
nand U13452 (N_13452,N_11716,N_10679);
or U13453 (N_13453,N_11625,N_11052);
xor U13454 (N_13454,N_11379,N_10689);
xor U13455 (N_13455,N_10537,N_11336);
xnor U13456 (N_13456,N_11524,N_10858);
and U13457 (N_13457,N_11079,N_11573);
nor U13458 (N_13458,N_11482,N_10628);
xnor U13459 (N_13459,N_11454,N_10908);
xnor U13460 (N_13460,N_11785,N_11903);
nand U13461 (N_13461,N_11692,N_10921);
xor U13462 (N_13462,N_11280,N_10744);
and U13463 (N_13463,N_10732,N_10703);
xnor U13464 (N_13464,N_11242,N_11954);
nor U13465 (N_13465,N_11997,N_10823);
and U13466 (N_13466,N_11302,N_11517);
nor U13467 (N_13467,N_10847,N_11576);
or U13468 (N_13468,N_11591,N_10584);
xnor U13469 (N_13469,N_10684,N_11745);
nor U13470 (N_13470,N_10981,N_10528);
or U13471 (N_13471,N_11505,N_11859);
nor U13472 (N_13472,N_11285,N_10512);
nand U13473 (N_13473,N_10812,N_11469);
or U13474 (N_13474,N_11774,N_11630);
nor U13475 (N_13475,N_11274,N_11402);
xnor U13476 (N_13476,N_10680,N_10846);
xnor U13477 (N_13477,N_11550,N_10500);
nand U13478 (N_13478,N_10870,N_10508);
nor U13479 (N_13479,N_10662,N_10886);
nor U13480 (N_13480,N_11009,N_11186);
nor U13481 (N_13481,N_11528,N_10598);
and U13482 (N_13482,N_11835,N_11789);
and U13483 (N_13483,N_11930,N_11466);
nand U13484 (N_13484,N_11837,N_10766);
xnor U13485 (N_13485,N_11278,N_11937);
nand U13486 (N_13486,N_10962,N_11978);
and U13487 (N_13487,N_11257,N_10517);
nand U13488 (N_13488,N_11369,N_10774);
nand U13489 (N_13489,N_11954,N_11313);
xor U13490 (N_13490,N_11033,N_11174);
and U13491 (N_13491,N_10518,N_10816);
or U13492 (N_13492,N_10613,N_11187);
nand U13493 (N_13493,N_10945,N_10813);
nor U13494 (N_13494,N_11147,N_10762);
xor U13495 (N_13495,N_11631,N_11771);
nor U13496 (N_13496,N_11374,N_10953);
nand U13497 (N_13497,N_11792,N_11163);
nor U13498 (N_13498,N_10564,N_11053);
or U13499 (N_13499,N_10585,N_11788);
xnor U13500 (N_13500,N_12452,N_13345);
nor U13501 (N_13501,N_12656,N_13127);
and U13502 (N_13502,N_12991,N_12136);
xor U13503 (N_13503,N_12607,N_13167);
nand U13504 (N_13504,N_12780,N_12082);
and U13505 (N_13505,N_13060,N_13148);
and U13506 (N_13506,N_13419,N_12603);
nor U13507 (N_13507,N_12554,N_13204);
xnor U13508 (N_13508,N_12071,N_12726);
nor U13509 (N_13509,N_12759,N_13066);
nor U13510 (N_13510,N_13331,N_12447);
xor U13511 (N_13511,N_12856,N_12496);
nand U13512 (N_13512,N_12464,N_12491);
or U13513 (N_13513,N_12631,N_13416);
and U13514 (N_13514,N_12530,N_13260);
or U13515 (N_13515,N_13139,N_12133);
xor U13516 (N_13516,N_13267,N_12242);
or U13517 (N_13517,N_13284,N_12016);
and U13518 (N_13518,N_13336,N_13128);
nand U13519 (N_13519,N_13003,N_12134);
or U13520 (N_13520,N_12694,N_12436);
nor U13521 (N_13521,N_12213,N_13394);
and U13522 (N_13522,N_12534,N_12976);
nand U13523 (N_13523,N_12728,N_13326);
or U13524 (N_13524,N_12186,N_13070);
or U13525 (N_13525,N_12426,N_13374);
nand U13526 (N_13526,N_12825,N_13401);
or U13527 (N_13527,N_13112,N_13485);
nand U13528 (N_13528,N_12766,N_12178);
nor U13529 (N_13529,N_13322,N_12386);
and U13530 (N_13530,N_13147,N_13094);
nand U13531 (N_13531,N_12244,N_12281);
nand U13532 (N_13532,N_12828,N_12095);
or U13533 (N_13533,N_13275,N_13019);
or U13534 (N_13534,N_12654,N_13467);
and U13535 (N_13535,N_13212,N_12472);
xnor U13536 (N_13536,N_12476,N_12589);
and U13537 (N_13537,N_12936,N_13365);
nand U13538 (N_13538,N_12255,N_12636);
and U13539 (N_13539,N_12968,N_12091);
nor U13540 (N_13540,N_12762,N_12323);
nand U13541 (N_13541,N_13218,N_12669);
nor U13542 (N_13542,N_12943,N_12684);
nand U13543 (N_13543,N_12751,N_12522);
xor U13544 (N_13544,N_13122,N_12482);
xor U13545 (N_13545,N_13107,N_12532);
or U13546 (N_13546,N_12785,N_13214);
and U13547 (N_13547,N_12754,N_13192);
or U13548 (N_13548,N_12682,N_12526);
nor U13549 (N_13549,N_12864,N_12911);
and U13550 (N_13550,N_12270,N_13347);
or U13551 (N_13551,N_12744,N_13186);
nand U13552 (N_13552,N_13451,N_12583);
and U13553 (N_13553,N_13184,N_13030);
nor U13554 (N_13554,N_12229,N_12498);
nand U13555 (N_13555,N_13156,N_12641);
xnor U13556 (N_13556,N_12233,N_13454);
xor U13557 (N_13557,N_12110,N_13450);
or U13558 (N_13558,N_13093,N_12351);
nor U13559 (N_13559,N_12942,N_13382);
or U13560 (N_13560,N_12548,N_13348);
xnor U13561 (N_13561,N_13325,N_13288);
and U13562 (N_13562,N_12542,N_12143);
nor U13563 (N_13563,N_12411,N_12459);
nand U13564 (N_13564,N_12346,N_12468);
and U13565 (N_13565,N_13163,N_12531);
and U13566 (N_13566,N_12153,N_13061);
and U13567 (N_13567,N_12981,N_12937);
nand U13568 (N_13568,N_12378,N_13209);
and U13569 (N_13569,N_13023,N_12608);
nand U13570 (N_13570,N_12695,N_13228);
xnor U13571 (N_13571,N_12356,N_13125);
nand U13572 (N_13572,N_12433,N_12929);
or U13573 (N_13573,N_12147,N_13010);
xnor U13574 (N_13574,N_12615,N_13299);
and U13575 (N_13575,N_13463,N_13196);
and U13576 (N_13576,N_13311,N_13152);
and U13577 (N_13577,N_12502,N_12814);
xnor U13578 (N_13578,N_13303,N_13457);
or U13579 (N_13579,N_12135,N_13466);
and U13580 (N_13580,N_12348,N_12473);
nand U13581 (N_13581,N_13042,N_12341);
and U13582 (N_13582,N_12232,N_12019);
or U13583 (N_13583,N_12500,N_13333);
nand U13584 (N_13584,N_12646,N_12081);
nor U13585 (N_13585,N_12432,N_12121);
nor U13586 (N_13586,N_12183,N_13404);
xor U13587 (N_13587,N_13358,N_12793);
nor U13588 (N_13588,N_12797,N_12268);
nor U13589 (N_13589,N_12640,N_12375);
or U13590 (N_13590,N_12558,N_12563);
or U13591 (N_13591,N_13216,N_12553);
nor U13592 (N_13592,N_12803,N_12519);
nor U13593 (N_13593,N_12959,N_12127);
nor U13594 (N_13594,N_12090,N_13320);
xnor U13595 (N_13595,N_12827,N_12696);
nor U13596 (N_13596,N_12824,N_13271);
and U13597 (N_13597,N_12345,N_12400);
nor U13598 (N_13598,N_12863,N_12679);
and U13599 (N_13599,N_12945,N_12484);
nor U13600 (N_13600,N_13161,N_12499);
and U13601 (N_13601,N_12449,N_13488);
or U13602 (N_13602,N_12822,N_12344);
nand U13603 (N_13603,N_12381,N_12077);
and U13604 (N_13604,N_13343,N_12117);
nand U13605 (N_13605,N_12601,N_12466);
or U13606 (N_13606,N_12703,N_12750);
or U13607 (N_13607,N_12957,N_13048);
xor U13608 (N_13608,N_12140,N_12755);
xor U13609 (N_13609,N_12031,N_13040);
nor U13610 (N_13610,N_12283,N_12892);
and U13611 (N_13611,N_12560,N_13084);
nor U13612 (N_13612,N_12561,N_13472);
or U13613 (N_13613,N_13460,N_12758);
xor U13614 (N_13614,N_13428,N_12632);
xor U13615 (N_13615,N_13456,N_12108);
nand U13616 (N_13616,N_12357,N_12152);
xnor U13617 (N_13617,N_12439,N_12673);
or U13618 (N_13618,N_13033,N_12305);
nor U13619 (N_13619,N_12141,N_13424);
nand U13620 (N_13620,N_12844,N_12312);
nor U13621 (N_13621,N_13407,N_12708);
or U13622 (N_13622,N_13123,N_13235);
nor U13623 (N_13623,N_12602,N_12579);
nor U13624 (N_13624,N_12799,N_12124);
xor U13625 (N_13625,N_12955,N_13130);
xnor U13626 (N_13626,N_12018,N_13285);
or U13627 (N_13627,N_12711,N_12410);
nand U13628 (N_13628,N_13195,N_12321);
nor U13629 (N_13629,N_12768,N_12836);
nor U13630 (N_13630,N_12774,N_12198);
or U13631 (N_13631,N_13118,N_13441);
or U13632 (N_13632,N_12585,N_12985);
nand U13633 (N_13633,N_12670,N_13124);
and U13634 (N_13634,N_13254,N_13263);
nand U13635 (N_13635,N_12061,N_12393);
nor U13636 (N_13636,N_12609,N_12201);
xnor U13637 (N_13637,N_12886,N_13402);
nand U13638 (N_13638,N_12672,N_12131);
xnor U13639 (N_13639,N_12079,N_13140);
nand U13640 (N_13640,N_13363,N_13221);
nor U13641 (N_13641,N_12279,N_12928);
nand U13642 (N_13642,N_12064,N_13206);
and U13643 (N_13643,N_12027,N_12816);
nand U13644 (N_13644,N_13442,N_12159);
or U13645 (N_13645,N_12635,N_12848);
and U13646 (N_13646,N_12083,N_13051);
xnor U13647 (N_13647,N_12151,N_12315);
nand U13648 (N_13648,N_12835,N_13266);
nor U13649 (N_13649,N_12205,N_12474);
xor U13650 (N_13650,N_12123,N_13079);
and U13651 (N_13651,N_12457,N_12555);
nor U13652 (N_13652,N_13487,N_12479);
xnor U13653 (N_13653,N_12330,N_13001);
xor U13654 (N_13654,N_12389,N_13421);
or U13655 (N_13655,N_13312,N_12206);
or U13656 (N_13656,N_12919,N_12567);
nor U13657 (N_13657,N_12597,N_12072);
and U13658 (N_13658,N_13222,N_12811);
nand U13659 (N_13659,N_12663,N_12256);
nand U13660 (N_13660,N_12409,N_12382);
or U13661 (N_13661,N_12508,N_13117);
and U13662 (N_13662,N_12450,N_13335);
xor U13663 (N_13663,N_12442,N_12873);
or U13664 (N_13664,N_12295,N_13364);
nor U13665 (N_13665,N_12009,N_12053);
or U13666 (N_13666,N_13174,N_12782);
nand U13667 (N_13667,N_13317,N_13481);
or U13668 (N_13668,N_13020,N_13141);
and U13669 (N_13669,N_12714,N_13352);
xnor U13670 (N_13670,N_12240,N_13330);
nand U13671 (N_13671,N_12717,N_12846);
and U13672 (N_13672,N_12556,N_12493);
nand U13673 (N_13673,N_12462,N_12520);
nor U13674 (N_13674,N_12986,N_13415);
nand U13675 (N_13675,N_12172,N_13302);
nor U13676 (N_13676,N_12176,N_13080);
and U13677 (N_13677,N_13110,N_12252);
or U13678 (N_13678,N_13439,N_13376);
or U13679 (N_13679,N_12819,N_12149);
nor U13680 (N_13680,N_12495,N_12595);
and U13681 (N_13681,N_12035,N_13381);
or U13682 (N_13682,N_13314,N_13417);
xor U13683 (N_13683,N_12817,N_13341);
xnor U13684 (N_13684,N_12210,N_13101);
or U13685 (N_13685,N_12277,N_12710);
nand U13686 (N_13686,N_12999,N_13105);
and U13687 (N_13687,N_12199,N_12021);
or U13688 (N_13688,N_12598,N_13461);
nand U13689 (N_13689,N_13159,N_12851);
xnor U13690 (N_13690,N_12309,N_12207);
xnor U13691 (N_13691,N_12823,N_12327);
xor U13692 (N_13692,N_12756,N_13129);
or U13693 (N_13693,N_12842,N_12338);
nor U13694 (N_13694,N_13445,N_12625);
or U13695 (N_13695,N_12700,N_12461);
or U13696 (N_13696,N_12888,N_13274);
nand U13697 (N_13697,N_12939,N_12644);
xnor U13698 (N_13698,N_12322,N_12593);
nand U13699 (N_13699,N_12078,N_12723);
or U13700 (N_13700,N_12221,N_12329);
nor U13701 (N_13701,N_13191,N_12773);
xor U13702 (N_13702,N_12489,N_13351);
and U13703 (N_13703,N_12852,N_12118);
xnor U13704 (N_13704,N_13058,N_12818);
xnor U13705 (N_13705,N_12107,N_13241);
or U13706 (N_13706,N_12249,N_13111);
nand U13707 (N_13707,N_12293,N_12834);
nor U13708 (N_13708,N_12045,N_12342);
or U13709 (N_13709,N_12582,N_12666);
nor U13710 (N_13710,N_12794,N_12926);
xor U13711 (N_13711,N_12676,N_13075);
or U13712 (N_13712,N_13057,N_12062);
and U13713 (N_13713,N_12866,N_12550);
nand U13714 (N_13714,N_13065,N_12047);
and U13715 (N_13715,N_12171,N_12004);
and U13716 (N_13716,N_12390,N_12421);
nand U13717 (N_13717,N_13164,N_13183);
and U13718 (N_13718,N_12306,N_12246);
nand U13719 (N_13719,N_13479,N_12335);
xnor U13720 (N_13720,N_13115,N_12704);
or U13721 (N_13721,N_12182,N_12282);
xor U13722 (N_13722,N_12689,N_12286);
xnor U13723 (N_13723,N_13046,N_12931);
xor U13724 (N_13724,N_12529,N_13091);
and U13725 (N_13725,N_12158,N_12006);
or U13726 (N_13726,N_12565,N_12397);
xor U13727 (N_13727,N_12285,N_12612);
nor U13728 (N_13728,N_12138,N_13484);
and U13729 (N_13729,N_12333,N_13283);
nor U13730 (N_13730,N_13398,N_12005);
nor U13731 (N_13731,N_12099,N_12022);
nand U13732 (N_13732,N_12362,N_12647);
or U13733 (N_13733,N_12320,N_13294);
xnor U13734 (N_13734,N_13410,N_12465);
and U13735 (N_13735,N_12494,N_12060);
and U13736 (N_13736,N_12645,N_12648);
nor U13737 (N_13737,N_13496,N_12103);
nor U13738 (N_13738,N_12687,N_12094);
nor U13739 (N_13739,N_12961,N_12254);
nand U13740 (N_13740,N_13012,N_12174);
or U13741 (N_13741,N_13025,N_13493);
xnor U13742 (N_13742,N_12874,N_12604);
xnor U13743 (N_13743,N_13366,N_13249);
and U13744 (N_13744,N_12829,N_12146);
and U13745 (N_13745,N_13154,N_13386);
or U13746 (N_13746,N_13006,N_12039);
or U13747 (N_13747,N_12288,N_12317);
or U13748 (N_13748,N_12020,N_12982);
nand U13749 (N_13749,N_12900,N_13134);
and U13750 (N_13750,N_12801,N_12313);
xor U13751 (N_13751,N_12787,N_12216);
or U13752 (N_13752,N_13319,N_13405);
nand U13753 (N_13753,N_12303,N_12169);
nor U13754 (N_13754,N_12841,N_13047);
nand U13755 (N_13755,N_13432,N_12741);
nand U13756 (N_13756,N_12838,N_12408);
or U13757 (N_13757,N_12188,N_12840);
nand U13758 (N_13758,N_13232,N_13328);
nand U13759 (N_13759,N_12055,N_13096);
or U13760 (N_13760,N_13280,N_12148);
xnor U13761 (N_13761,N_12506,N_12651);
nand U13762 (N_13762,N_12964,N_13272);
nor U13763 (N_13763,N_12092,N_13197);
and U13764 (N_13764,N_12879,N_12638);
xor U13765 (N_13765,N_12332,N_12424);
nand U13766 (N_13766,N_13226,N_13473);
xnor U13767 (N_13767,N_12273,N_13138);
or U13768 (N_13768,N_13434,N_13056);
xnor U13769 (N_13769,N_13356,N_12853);
and U13770 (N_13770,N_12951,N_13172);
and U13771 (N_13771,N_12969,N_12440);
or U13772 (N_13772,N_12056,N_13081);
nand U13773 (N_13773,N_12738,N_12260);
xnor U13774 (N_13774,N_12671,N_12865);
or U13775 (N_13775,N_12847,N_13339);
nor U13776 (N_13776,N_13009,N_12620);
or U13777 (N_13777,N_12521,N_13413);
or U13778 (N_13778,N_12992,N_13305);
xnor U13779 (N_13779,N_12264,N_12403);
nor U13780 (N_13780,N_12924,N_12425);
xor U13781 (N_13781,N_12204,N_12513);
nor U13782 (N_13782,N_12517,N_12231);
xor U13783 (N_13783,N_13106,N_12328);
nor U13784 (N_13784,N_13470,N_13492);
and U13785 (N_13785,N_12105,N_12987);
and U13786 (N_13786,N_12516,N_12225);
nor U13787 (N_13787,N_12340,N_12114);
and U13788 (N_13788,N_12736,N_12034);
or U13789 (N_13789,N_12958,N_12184);
or U13790 (N_13790,N_13121,N_12952);
or U13791 (N_13791,N_12074,N_13286);
nand U13792 (N_13792,N_12990,N_12463);
xnor U13793 (N_13793,N_12680,N_13227);
and U13794 (N_13794,N_12239,N_12668);
and U13795 (N_13795,N_12798,N_12012);
nand U13796 (N_13796,N_12324,N_13368);
nor U13797 (N_13797,N_12524,N_12549);
nand U13798 (N_13798,N_13022,N_12456);
or U13799 (N_13799,N_13133,N_13225);
xnor U13800 (N_13800,N_13002,N_12304);
and U13801 (N_13801,N_13392,N_12434);
nor U13802 (N_13802,N_13211,N_12490);
nor U13803 (N_13803,N_12831,N_12525);
nand U13804 (N_13804,N_12407,N_12975);
nand U13805 (N_13805,N_12977,N_12483);
xor U13806 (N_13806,N_12956,N_12712);
or U13807 (N_13807,N_12308,N_12788);
nor U13808 (N_13808,N_13433,N_13114);
nor U13809 (N_13809,N_12963,N_12245);
or U13810 (N_13810,N_12259,N_13248);
and U13811 (N_13811,N_13449,N_12940);
xor U13812 (N_13812,N_13074,N_13373);
nand U13813 (N_13813,N_12692,N_12705);
xor U13814 (N_13814,N_12298,N_13372);
nand U13815 (N_13815,N_13188,N_12454);
nor U13816 (N_13816,N_12112,N_12241);
and U13817 (N_13817,N_12528,N_12997);
xor U13818 (N_13818,N_12545,N_12037);
and U13819 (N_13819,N_13296,N_13068);
and U13820 (N_13820,N_12301,N_13168);
nand U13821 (N_13821,N_12272,N_12427);
xnor U13822 (N_13822,N_12059,N_12721);
xnor U13823 (N_13823,N_12278,N_12869);
or U13824 (N_13824,N_12574,N_12302);
or U13825 (N_13825,N_12420,N_12935);
and U13826 (N_13826,N_13256,N_12808);
or U13827 (N_13827,N_12032,N_12753);
and U13828 (N_13828,N_12748,N_12209);
nand U13829 (N_13829,N_12139,N_12662);
or U13830 (N_13830,N_13032,N_12876);
or U13831 (N_13831,N_13090,N_12292);
xnor U13832 (N_13832,N_13116,N_13202);
or U13833 (N_13833,N_12104,N_13474);
or U13834 (N_13834,N_12129,N_12170);
and U13835 (N_13835,N_12683,N_12938);
nor U13836 (N_13836,N_12445,N_12331);
nor U13837 (N_13837,N_13119,N_12591);
nor U13838 (N_13838,N_12984,N_12097);
or U13839 (N_13839,N_13420,N_12236);
nand U13840 (N_13840,N_13471,N_12578);
and U13841 (N_13841,N_12419,N_13224);
nor U13842 (N_13842,N_13108,N_12967);
or U13843 (N_13843,N_12781,N_13189);
nor U13844 (N_13844,N_13077,N_12802);
and U13845 (N_13845,N_12966,N_13327);
and U13846 (N_13846,N_12622,N_12540);
nand U13847 (N_13847,N_13013,N_12894);
and U13848 (N_13848,N_12533,N_12353);
nand U13849 (N_13849,N_13017,N_13099);
xor U13850 (N_13850,N_12150,N_13337);
nand U13851 (N_13851,N_12905,N_12181);
nand U13852 (N_13852,N_13103,N_12718);
and U13853 (N_13853,N_12763,N_12993);
or U13854 (N_13854,N_12891,N_13045);
xor U13855 (N_13855,N_12383,N_13403);
nand U13856 (N_13856,N_13092,N_13478);
nand U13857 (N_13857,N_12971,N_13237);
nand U13858 (N_13858,N_12478,N_12460);
nand U13859 (N_13859,N_13321,N_12044);
and U13860 (N_13860,N_12996,N_12510);
or U13861 (N_13861,N_13253,N_12180);
or U13862 (N_13862,N_12610,N_12568);
nor U13863 (N_13863,N_12566,N_12994);
or U13864 (N_13864,N_12211,N_13464);
or U13865 (N_13865,N_12222,N_12435);
xnor U13866 (N_13866,N_12551,N_12889);
or U13867 (N_13867,N_12675,N_13295);
nand U13868 (N_13868,N_12230,N_12477);
nand U13869 (N_13869,N_12821,N_13397);
nor U13870 (N_13870,N_12480,N_12275);
nand U13871 (N_13871,N_13297,N_12605);
and U13872 (N_13872,N_13465,N_12024);
nand U13873 (N_13873,N_12248,N_13126);
nor U13874 (N_13874,N_12458,N_12161);
or U13875 (N_13875,N_12194,N_12901);
and U13876 (N_13876,N_12227,N_12953);
nor U13877 (N_13877,N_13483,N_12623);
or U13878 (N_13878,N_13037,N_13458);
or U13879 (N_13879,N_12202,N_12757);
nand U13880 (N_13880,N_12902,N_13005);
or U13881 (N_13881,N_12843,N_12405);
nand U13882 (N_13882,N_12734,N_12980);
and U13883 (N_13883,N_12890,N_12946);
nor U13884 (N_13884,N_13257,N_13088);
nand U13885 (N_13885,N_12065,N_12310);
or U13886 (N_13886,N_12041,N_13477);
nand U13887 (N_13887,N_13313,N_13323);
xnor U13888 (N_13888,N_12287,N_13053);
and U13889 (N_13889,N_12339,N_13166);
nand U13890 (N_13890,N_13059,N_12747);
nand U13891 (N_13891,N_12057,N_12974);
or U13892 (N_13892,N_13318,N_12307);
and U13893 (N_13893,N_12862,N_12810);
nor U13894 (N_13894,N_13316,N_12882);
or U13895 (N_13895,N_12572,N_13446);
and U13896 (N_13896,N_13043,N_13499);
xnor U13897 (N_13897,N_13004,N_12155);
xnor U13898 (N_13898,N_12897,N_12637);
or U13899 (N_13899,N_13269,N_12514);
and U13900 (N_13900,N_12617,N_13264);
xor U13901 (N_13901,N_12970,N_13489);
nor U13902 (N_13902,N_13052,N_12923);
xnor U13903 (N_13903,N_12903,N_12337);
xor U13904 (N_13904,N_12707,N_12515);
and U13905 (N_13905,N_12765,N_12173);
and U13906 (N_13906,N_12557,N_12665);
and U13907 (N_13907,N_12523,N_12850);
or U13908 (N_13908,N_13438,N_12014);
or U13909 (N_13909,N_12167,N_13007);
or U13910 (N_13910,N_13422,N_12789);
nor U13911 (N_13911,N_12664,N_12126);
and U13912 (N_13912,N_13262,N_12311);
xor U13913 (N_13913,N_12412,N_12978);
nand U13914 (N_13914,N_12616,N_12350);
or U13915 (N_13915,N_12359,N_12051);
and U13916 (N_13916,N_12261,N_12237);
or U13917 (N_13917,N_12069,N_12373);
and U13918 (N_13918,N_12577,N_13360);
xor U13919 (N_13919,N_12394,N_12701);
and U13920 (N_13920,N_12415,N_12196);
xnor U13921 (N_13921,N_12830,N_12659);
nand U13922 (N_13922,N_12366,N_12475);
nor U13923 (N_13923,N_12764,N_13246);
or U13924 (N_13924,N_13137,N_13095);
or U13925 (N_13925,N_12446,N_12581);
nor U13926 (N_13926,N_13389,N_12076);
and U13927 (N_13927,N_12398,N_13251);
xor U13928 (N_13928,N_12989,N_13086);
nand U13929 (N_13929,N_13359,N_12179);
xor U13930 (N_13930,N_13200,N_12621);
nor U13931 (N_13931,N_13240,N_12404);
nor U13932 (N_13932,N_12336,N_13062);
nor U13933 (N_13933,N_12023,N_12538);
nand U13934 (N_13934,N_12226,N_12049);
nor U13935 (N_13935,N_12733,N_12907);
and U13936 (N_13936,N_12029,N_13270);
or U13937 (N_13937,N_12401,N_13245);
and U13938 (N_13938,N_12085,N_13089);
nand U13939 (N_13939,N_12909,N_12776);
and U13940 (N_13940,N_12354,N_12297);
and U13941 (N_13941,N_13076,N_12002);
xor U13942 (N_13942,N_12507,N_13354);
xnor U13943 (N_13943,N_12017,N_12594);
xnor U13944 (N_13944,N_12068,N_13193);
and U13945 (N_13945,N_13063,N_12391);
or U13946 (N_13946,N_12742,N_12629);
and U13947 (N_13947,N_13252,N_13082);
nor U13948 (N_13948,N_12347,N_12699);
and U13949 (N_13949,N_12932,N_12486);
or U13950 (N_13950,N_12364,N_12492);
or U13951 (N_13951,N_12904,N_12887);
xnor U13952 (N_13952,N_13338,N_13170);
nor U13953 (N_13953,N_13036,N_12715);
and U13954 (N_13954,N_13306,N_12387);
nor U13955 (N_13955,N_12786,N_12043);
or U13956 (N_13956,N_12284,N_13379);
xnor U13957 (N_13957,N_13038,N_12485);
and U13958 (N_13958,N_12535,N_12238);
nor U13959 (N_13959,N_12512,N_12451);
or U13960 (N_13960,N_13437,N_12916);
and U13961 (N_13961,N_12693,N_12655);
nand U13962 (N_13962,N_12455,N_13250);
xnor U13963 (N_13963,N_13243,N_12036);
xor U13964 (N_13964,N_12368,N_12294);
nor U13965 (N_13965,N_12193,N_12208);
xor U13966 (N_13966,N_12243,N_13162);
and U13967 (N_13967,N_12849,N_12125);
nand U13968 (N_13968,N_13255,N_13229);
xor U13969 (N_13969,N_13261,N_13165);
and U13970 (N_13970,N_12716,N_12326);
xor U13971 (N_13971,N_12487,N_13380);
or U13972 (N_13972,N_12509,N_13021);
or U13973 (N_13973,N_12875,N_13355);
or U13974 (N_13974,N_12089,N_12767);
nor U13975 (N_13975,N_12720,N_12428);
and U13976 (N_13976,N_12195,N_12224);
or U13977 (N_13977,N_12070,N_13220);
nand U13978 (N_13978,N_12571,N_12883);
nand U13979 (N_13979,N_13178,N_12973);
and U13980 (N_13980,N_12437,N_12795);
xor U13981 (N_13981,N_12732,N_12026);
and U13982 (N_13982,N_12417,N_13034);
or U13983 (N_13983,N_13334,N_12448);
nor U13984 (N_13984,N_12011,N_13155);
nand U13985 (N_13985,N_12779,N_12592);
nand U13986 (N_13986,N_13342,N_13072);
or U13987 (N_13987,N_12947,N_12925);
nor U13988 (N_13988,N_12380,N_12395);
and U13989 (N_13989,N_12584,N_12422);
nor U13990 (N_13990,N_13390,N_13149);
and U13991 (N_13991,N_13406,N_13375);
and U13992 (N_13992,N_12769,N_13055);
nor U13993 (N_13993,N_12719,N_13026);
nand U13994 (N_13994,N_13370,N_13219);
nand U13995 (N_13995,N_13304,N_13011);
or U13996 (N_13996,N_13287,N_13169);
or U13997 (N_13997,N_12771,N_12086);
nor U13998 (N_13998,N_13495,N_12739);
nand U13999 (N_13999,N_12343,N_12423);
nand U14000 (N_14000,N_13367,N_13015);
xor U14001 (N_14001,N_13497,N_12015);
and U14002 (N_14002,N_12300,N_12948);
xor U14003 (N_14003,N_13244,N_12003);
and U14004 (N_14004,N_13258,N_13447);
xor U14005 (N_14005,N_12511,N_12804);
xor U14006 (N_14006,N_12972,N_13029);
nand U14007 (N_14007,N_13289,N_12730);
nand U14008 (N_14008,N_12096,N_12861);
nand U14009 (N_14009,N_12737,N_13215);
and U14010 (N_14010,N_12652,N_13292);
xnor U14011 (N_14011,N_12618,N_12219);
nor U14012 (N_14012,N_12677,N_13230);
and U14013 (N_14013,N_13131,N_13309);
nand U14014 (N_14014,N_13078,N_13282);
xor U14015 (N_14015,N_12745,N_12575);
or U14016 (N_14016,N_12546,N_13435);
and U14017 (N_14017,N_12899,N_12441);
xnor U14018 (N_14018,N_12042,N_12130);
nand U14019 (N_14019,N_12590,N_13344);
or U14020 (N_14020,N_12087,N_12746);
nor U14021 (N_14021,N_12257,N_12376);
nand U14022 (N_14022,N_12467,N_12918);
or U14023 (N_14023,N_12430,N_12469);
or U14024 (N_14024,N_12291,N_13350);
or U14025 (N_14025,N_12267,N_12740);
nand U14026 (N_14026,N_12218,N_13357);
or U14027 (N_14027,N_12010,N_13377);
nor U14028 (N_14028,N_12253,N_13102);
and U14029 (N_14029,N_12541,N_13098);
xnor U14030 (N_14030,N_12895,N_12361);
xor U14031 (N_14031,N_12318,N_13028);
or U14032 (N_14032,N_12262,N_13194);
or U14033 (N_14033,N_13073,N_13361);
nand U14034 (N_14034,N_12377,N_12743);
nor U14035 (N_14035,N_13332,N_12367);
or U14036 (N_14036,N_12352,N_12860);
nor U14037 (N_14037,N_12634,N_13423);
or U14038 (N_14038,N_12429,N_12806);
nand U14039 (N_14039,N_12690,N_12633);
and U14040 (N_14040,N_12698,N_13329);
nand U14041 (N_14041,N_13018,N_13412);
or U14042 (N_14042,N_12325,N_12599);
nand U14043 (N_14043,N_12413,N_12443);
and U14044 (N_14044,N_12100,N_12772);
and U14045 (N_14045,N_12922,N_13238);
nor U14046 (N_14046,N_12163,N_12657);
or U14047 (N_14047,N_12885,N_12867);
nor U14048 (N_14048,N_12630,N_12667);
nand U14049 (N_14049,N_12674,N_12431);
xor U14050 (N_14050,N_12562,N_13378);
and U14051 (N_14051,N_12438,N_13181);
nor U14052 (N_14052,N_12857,N_12685);
nor U14053 (N_14053,N_12000,N_12688);
nand U14054 (N_14054,N_13024,N_13418);
and U14055 (N_14055,N_12950,N_12223);
nor U14056 (N_14056,N_13400,N_12912);
nor U14057 (N_14057,N_12777,N_12576);
nand U14058 (N_14058,N_13486,N_13468);
xnor U14059 (N_14059,N_12709,N_12722);
or U14060 (N_14060,N_13031,N_12274);
and U14061 (N_14061,N_13340,N_13016);
or U14062 (N_14062,N_13279,N_12063);
nand U14063 (N_14063,N_12067,N_13490);
nor U14064 (N_14064,N_12185,N_12266);
nand U14065 (N_14065,N_12775,N_12941);
or U14066 (N_14066,N_12796,N_12543);
and U14067 (N_14067,N_12770,N_12586);
nor U14068 (N_14068,N_13462,N_12157);
or U14069 (N_14069,N_13187,N_12119);
nor U14070 (N_14070,N_13476,N_12388);
xnor U14071 (N_14071,N_13213,N_12639);
and U14072 (N_14072,N_12080,N_12660);
or U14073 (N_14073,N_12212,N_13157);
or U14074 (N_14074,N_12833,N_13039);
and U14075 (N_14075,N_12858,N_12058);
and U14076 (N_14076,N_12691,N_13071);
and U14077 (N_14077,N_12289,N_12501);
and U14078 (N_14078,N_12162,N_13298);
or U14079 (N_14079,N_12215,N_13498);
nor U14080 (N_14080,N_13310,N_13158);
and U14081 (N_14081,N_13315,N_12109);
nor U14082 (N_14082,N_12142,N_13049);
and U14083 (N_14083,N_13411,N_12156);
nand U14084 (N_14084,N_13277,N_13436);
xnor U14085 (N_14085,N_12600,N_12790);
and U14086 (N_14086,N_12132,N_13480);
or U14087 (N_14087,N_12536,N_13180);
or U14088 (N_14088,N_13145,N_12896);
and U14089 (N_14089,N_13324,N_12048);
and U14090 (N_14090,N_12872,N_12650);
nor U14091 (N_14091,N_12760,N_13143);
nand U14092 (N_14092,N_12372,N_13268);
or U14093 (N_14093,N_12234,N_13455);
xnor U14094 (N_14094,N_12191,N_13459);
xor U14095 (N_14095,N_12166,N_12653);
nor U14096 (N_14096,N_12220,N_13199);
nand U14097 (N_14097,N_13430,N_12778);
nor U14098 (N_14098,N_13142,N_12933);
xor U14099 (N_14099,N_13231,N_12649);
and U14100 (N_14100,N_12878,N_12392);
nand U14101 (N_14101,N_12877,N_12137);
xnor U14102 (N_14102,N_12122,N_13469);
and U14103 (N_14103,N_12559,N_12954);
xnor U14104 (N_14104,N_13205,N_13395);
nand U14105 (N_14105,N_12265,N_12399);
xnor U14106 (N_14106,N_13069,N_12374);
nor U14107 (N_14107,N_12111,N_12627);
xnor U14108 (N_14108,N_12235,N_12870);
nor U14109 (N_14109,N_12573,N_13239);
nor U14110 (N_14110,N_12809,N_12661);
nand U14111 (N_14111,N_13083,N_12093);
or U14112 (N_14112,N_12488,N_13427);
nand U14113 (N_14113,N_13388,N_12370);
xnor U14114 (N_14114,N_12624,N_12190);
nor U14115 (N_14115,N_13431,N_12033);
nor U14116 (N_14116,N_13097,N_13217);
and U14117 (N_14117,N_12921,N_13000);
nand U14118 (N_14118,N_13050,N_12731);
nand U14119 (N_14119,N_13176,N_13444);
nor U14120 (N_14120,N_13475,N_12930);
and U14121 (N_14121,N_13369,N_12839);
nand U14122 (N_14122,N_13175,N_12815);
or U14123 (N_14123,N_12406,N_12416);
xor U14124 (N_14124,N_12914,N_13399);
nor U14125 (N_14125,N_12098,N_12396);
nor U14126 (N_14126,N_12503,N_12314);
and U14127 (N_14127,N_13113,N_12832);
nor U14128 (N_14128,N_13136,N_12168);
and U14129 (N_14129,N_12552,N_13210);
and U14130 (N_14130,N_12363,N_12013);
or U14131 (N_14131,N_12518,N_13008);
nand U14132 (N_14132,N_12588,N_12038);
nor U14133 (N_14133,N_12197,N_12547);
or U14134 (N_14134,N_12702,N_12564);
nor U14135 (N_14135,N_12725,N_13385);
nand U14136 (N_14136,N_12189,N_12250);
nor U14137 (N_14137,N_13179,N_12881);
nor U14138 (N_14138,N_12028,N_12784);
or U14139 (N_14139,N_13426,N_13160);
xnor U14140 (N_14140,N_12884,N_12384);
nand U14141 (N_14141,N_13393,N_13391);
nor U14142 (N_14142,N_12379,N_12800);
nand U14143 (N_14143,N_12481,N_13120);
or U14144 (N_14144,N_13035,N_12713);
and U14145 (N_14145,N_12606,N_12596);
and U14146 (N_14146,N_12101,N_13054);
and U14147 (N_14147,N_12871,N_13198);
xor U14148 (N_14148,N_13109,N_13100);
nand U14149 (N_14149,N_13182,N_13353);
nand U14150 (N_14150,N_12812,N_13201);
nor U14151 (N_14151,N_12537,N_13276);
nor U14152 (N_14152,N_12263,N_12910);
xor U14153 (N_14153,N_12965,N_12106);
nand U14154 (N_14154,N_12280,N_13234);
or U14155 (N_14155,N_12115,N_13087);
xor U14156 (N_14156,N_12418,N_12187);
or U14157 (N_14157,N_12102,N_12820);
nor U14158 (N_14158,N_12073,N_12160);
or U14159 (N_14159,N_12355,N_12611);
or U14160 (N_14160,N_12128,N_12030);
nor U14161 (N_14161,N_13247,N_12007);
and U14162 (N_14162,N_12228,N_13135);
and U14163 (N_14163,N_13085,N_12807);
xnor U14164 (N_14164,N_12749,N_12251);
xnor U14165 (N_14165,N_12165,N_12983);
and U14166 (N_14166,N_13104,N_13223);
or U14167 (N_14167,N_12628,N_13185);
and U14168 (N_14168,N_12052,N_12658);
nand U14169 (N_14169,N_12920,N_12619);
xor U14170 (N_14170,N_12761,N_13408);
or U14171 (N_14171,N_13064,N_12040);
xor U14172 (N_14172,N_12296,N_12360);
and U14173 (N_14173,N_12614,N_12643);
or U14174 (N_14174,N_12706,N_12358);
nand U14175 (N_14175,N_12046,N_12164);
nor U14176 (N_14176,N_12505,N_13281);
and U14177 (N_14177,N_12893,N_12995);
and U14178 (N_14178,N_12001,N_12203);
or U14179 (N_14179,N_12470,N_12783);
nor U14180 (N_14180,N_12686,N_12913);
or U14181 (N_14181,N_12845,N_13425);
or U14182 (N_14182,N_13293,N_12414);
nor U14183 (N_14183,N_12949,N_13429);
nor U14184 (N_14184,N_12544,N_12580);
nor U14185 (N_14185,N_13414,N_12144);
or U14186 (N_14186,N_13259,N_12681);
nor U14187 (N_14187,N_12217,N_12587);
nor U14188 (N_14188,N_12570,N_12247);
nor U14189 (N_14189,N_12050,N_12154);
xnor U14190 (N_14190,N_13242,N_13173);
or U14191 (N_14191,N_12319,N_13396);
xnor U14192 (N_14192,N_13494,N_13291);
nand U14193 (N_14193,N_13409,N_13265);
or U14194 (N_14194,N_13290,N_12290);
nor U14195 (N_14195,N_12444,N_12539);
xnor U14196 (N_14196,N_12258,N_12402);
or U14197 (N_14197,N_13177,N_12120);
nand U14198 (N_14198,N_12979,N_12276);
nor U14199 (N_14199,N_12504,N_12678);
or U14200 (N_14200,N_12088,N_13371);
xor U14201 (N_14201,N_12497,N_12214);
or U14202 (N_14202,N_12697,N_12271);
and U14203 (N_14203,N_12385,N_13383);
xnor U14204 (N_14204,N_13482,N_13452);
and U14205 (N_14205,N_12906,N_12880);
xnor U14206 (N_14206,N_12349,N_13233);
nor U14207 (N_14207,N_12724,N_12962);
nor U14208 (N_14208,N_13308,N_12116);
nand U14209 (N_14209,N_12145,N_12898);
xor U14210 (N_14210,N_12066,N_13132);
or U14211 (N_14211,N_12369,N_13387);
nor U14212 (N_14212,N_13346,N_12200);
xnor U14213 (N_14213,N_13027,N_12113);
xor U14214 (N_14214,N_13044,N_12177);
nor U14215 (N_14215,N_12805,N_12752);
nand U14216 (N_14216,N_12371,N_13153);
nand U14217 (N_14217,N_12334,N_12915);
nand U14218 (N_14218,N_13491,N_12084);
and U14219 (N_14219,N_13448,N_12453);
nand U14220 (N_14220,N_13453,N_13150);
nand U14221 (N_14221,N_13144,N_12569);
xor U14222 (N_14222,N_12729,N_12859);
and U14223 (N_14223,N_12008,N_13307);
or U14224 (N_14224,N_13203,N_12365);
nor U14225 (N_14225,N_12054,N_13041);
xor U14226 (N_14226,N_12917,N_13014);
or U14227 (N_14227,N_12855,N_13273);
and U14228 (N_14228,N_12626,N_12727);
nand U14229 (N_14229,N_13146,N_12471);
and U14230 (N_14230,N_12316,N_13349);
and U14231 (N_14231,N_12642,N_12988);
or U14232 (N_14232,N_13151,N_12792);
nor U14233 (N_14233,N_12868,N_13443);
nand U14234 (N_14234,N_13440,N_12613);
and U14235 (N_14235,N_12998,N_13236);
nand U14236 (N_14236,N_12175,N_12025);
or U14237 (N_14237,N_12927,N_12735);
or U14238 (N_14238,N_13300,N_12791);
nand U14239 (N_14239,N_13384,N_12527);
xor U14240 (N_14240,N_13171,N_12075);
nand U14241 (N_14241,N_12826,N_12934);
nand U14242 (N_14242,N_12854,N_12908);
xor U14243 (N_14243,N_13301,N_12813);
nand U14244 (N_14244,N_12944,N_12269);
nor U14245 (N_14245,N_13190,N_12299);
nor U14246 (N_14246,N_12192,N_13362);
or U14247 (N_14247,N_13278,N_13207);
nand U14248 (N_14248,N_12960,N_13067);
or U14249 (N_14249,N_13208,N_12837);
nor U14250 (N_14250,N_12738,N_12761);
nand U14251 (N_14251,N_12647,N_12524);
or U14252 (N_14252,N_13147,N_12038);
nand U14253 (N_14253,N_12784,N_12047);
and U14254 (N_14254,N_13168,N_12977);
and U14255 (N_14255,N_12552,N_13092);
and U14256 (N_14256,N_12535,N_12458);
or U14257 (N_14257,N_12622,N_12444);
nor U14258 (N_14258,N_13069,N_13203);
xnor U14259 (N_14259,N_13441,N_12855);
and U14260 (N_14260,N_12542,N_13192);
and U14261 (N_14261,N_12742,N_12096);
nor U14262 (N_14262,N_12833,N_12194);
nor U14263 (N_14263,N_12116,N_12907);
or U14264 (N_14264,N_13391,N_13298);
nand U14265 (N_14265,N_12027,N_12433);
nand U14266 (N_14266,N_12560,N_12483);
nor U14267 (N_14267,N_13228,N_12915);
and U14268 (N_14268,N_13277,N_12718);
and U14269 (N_14269,N_12079,N_12402);
or U14270 (N_14270,N_13481,N_13193);
or U14271 (N_14271,N_12568,N_12470);
nand U14272 (N_14272,N_12228,N_13083);
nor U14273 (N_14273,N_12585,N_13366);
nor U14274 (N_14274,N_12526,N_13318);
xnor U14275 (N_14275,N_12529,N_12686);
nor U14276 (N_14276,N_12738,N_12601);
xnor U14277 (N_14277,N_12349,N_12669);
xnor U14278 (N_14278,N_13385,N_12434);
or U14279 (N_14279,N_12494,N_12910);
nor U14280 (N_14280,N_13407,N_13202);
nor U14281 (N_14281,N_12650,N_12952);
and U14282 (N_14282,N_12322,N_13080);
or U14283 (N_14283,N_12318,N_12576);
or U14284 (N_14284,N_12225,N_12432);
or U14285 (N_14285,N_13497,N_13014);
xnor U14286 (N_14286,N_13401,N_12519);
nand U14287 (N_14287,N_12379,N_12502);
nor U14288 (N_14288,N_12368,N_13203);
xor U14289 (N_14289,N_12501,N_12909);
and U14290 (N_14290,N_13138,N_12849);
or U14291 (N_14291,N_12949,N_12543);
nand U14292 (N_14292,N_13072,N_12929);
xor U14293 (N_14293,N_12822,N_13337);
or U14294 (N_14294,N_13194,N_13162);
nand U14295 (N_14295,N_12251,N_12420);
nand U14296 (N_14296,N_12605,N_12389);
nor U14297 (N_14297,N_12296,N_13334);
or U14298 (N_14298,N_13074,N_13227);
and U14299 (N_14299,N_12133,N_12260);
and U14300 (N_14300,N_13037,N_12653);
and U14301 (N_14301,N_12062,N_12757);
nor U14302 (N_14302,N_12736,N_12526);
nand U14303 (N_14303,N_13158,N_12737);
nand U14304 (N_14304,N_13366,N_13452);
and U14305 (N_14305,N_12951,N_12326);
and U14306 (N_14306,N_13195,N_13129);
or U14307 (N_14307,N_12696,N_12461);
and U14308 (N_14308,N_13358,N_12872);
or U14309 (N_14309,N_12022,N_12984);
nand U14310 (N_14310,N_12435,N_12966);
nand U14311 (N_14311,N_12462,N_12219);
xnor U14312 (N_14312,N_13004,N_12869);
nor U14313 (N_14313,N_12401,N_12814);
and U14314 (N_14314,N_13051,N_12687);
and U14315 (N_14315,N_13095,N_12640);
or U14316 (N_14316,N_12291,N_12881);
or U14317 (N_14317,N_13272,N_12575);
nor U14318 (N_14318,N_13396,N_12143);
or U14319 (N_14319,N_12177,N_13395);
nand U14320 (N_14320,N_12290,N_12319);
or U14321 (N_14321,N_13496,N_12681);
nor U14322 (N_14322,N_12271,N_12005);
or U14323 (N_14323,N_12409,N_13491);
nand U14324 (N_14324,N_12774,N_12087);
and U14325 (N_14325,N_13035,N_12333);
nand U14326 (N_14326,N_13138,N_12230);
nor U14327 (N_14327,N_12987,N_12841);
or U14328 (N_14328,N_12592,N_12303);
nand U14329 (N_14329,N_13230,N_12375);
and U14330 (N_14330,N_12308,N_12894);
and U14331 (N_14331,N_12108,N_12524);
xor U14332 (N_14332,N_13232,N_12183);
nand U14333 (N_14333,N_12247,N_13018);
and U14334 (N_14334,N_12159,N_12429);
nor U14335 (N_14335,N_12135,N_12450);
or U14336 (N_14336,N_12762,N_13451);
xnor U14337 (N_14337,N_12158,N_13088);
nand U14338 (N_14338,N_12672,N_12680);
nor U14339 (N_14339,N_12656,N_13480);
and U14340 (N_14340,N_12271,N_12672);
xor U14341 (N_14341,N_13259,N_13099);
and U14342 (N_14342,N_13080,N_12235);
nor U14343 (N_14343,N_13379,N_12859);
xor U14344 (N_14344,N_13384,N_12191);
or U14345 (N_14345,N_12465,N_12193);
nand U14346 (N_14346,N_12955,N_12750);
xor U14347 (N_14347,N_12727,N_13023);
and U14348 (N_14348,N_12981,N_12338);
or U14349 (N_14349,N_12879,N_13440);
xnor U14350 (N_14350,N_12679,N_12169);
and U14351 (N_14351,N_13418,N_13408);
nor U14352 (N_14352,N_13052,N_12027);
nor U14353 (N_14353,N_12138,N_13327);
xnor U14354 (N_14354,N_12494,N_13237);
nand U14355 (N_14355,N_13247,N_13485);
xor U14356 (N_14356,N_12815,N_12463);
nor U14357 (N_14357,N_13156,N_13352);
nor U14358 (N_14358,N_12875,N_13262);
nand U14359 (N_14359,N_12228,N_13323);
or U14360 (N_14360,N_12776,N_12375);
nand U14361 (N_14361,N_12188,N_12654);
xor U14362 (N_14362,N_12350,N_12971);
xor U14363 (N_14363,N_12983,N_12476);
or U14364 (N_14364,N_12048,N_12703);
xor U14365 (N_14365,N_12767,N_12235);
nor U14366 (N_14366,N_12451,N_12349);
or U14367 (N_14367,N_12198,N_13435);
and U14368 (N_14368,N_12076,N_12115);
nor U14369 (N_14369,N_13404,N_12156);
nand U14370 (N_14370,N_13014,N_12058);
nand U14371 (N_14371,N_12790,N_12089);
nand U14372 (N_14372,N_13268,N_12997);
xor U14373 (N_14373,N_12444,N_12246);
xor U14374 (N_14374,N_13236,N_12857);
nor U14375 (N_14375,N_13349,N_12400);
or U14376 (N_14376,N_12949,N_13185);
nor U14377 (N_14377,N_13223,N_12373);
nand U14378 (N_14378,N_12443,N_13377);
nor U14379 (N_14379,N_13424,N_12165);
xnor U14380 (N_14380,N_13076,N_12937);
xnor U14381 (N_14381,N_12802,N_12954);
or U14382 (N_14382,N_13158,N_13009);
and U14383 (N_14383,N_13255,N_13006);
or U14384 (N_14384,N_12630,N_13234);
nand U14385 (N_14385,N_13056,N_12807);
and U14386 (N_14386,N_13211,N_13136);
or U14387 (N_14387,N_12355,N_12758);
nor U14388 (N_14388,N_12496,N_12880);
nor U14389 (N_14389,N_12816,N_12892);
nand U14390 (N_14390,N_12604,N_12609);
or U14391 (N_14391,N_12203,N_13132);
xnor U14392 (N_14392,N_12143,N_12603);
nand U14393 (N_14393,N_13449,N_13092);
nand U14394 (N_14394,N_13366,N_12615);
xnor U14395 (N_14395,N_12094,N_12640);
xnor U14396 (N_14396,N_12006,N_12533);
nor U14397 (N_14397,N_12210,N_12539);
nor U14398 (N_14398,N_12881,N_12767);
nand U14399 (N_14399,N_12856,N_12112);
xor U14400 (N_14400,N_12926,N_12893);
or U14401 (N_14401,N_12856,N_12463);
xnor U14402 (N_14402,N_12887,N_12687);
and U14403 (N_14403,N_12815,N_12296);
nand U14404 (N_14404,N_12403,N_12219);
or U14405 (N_14405,N_12162,N_12000);
and U14406 (N_14406,N_12972,N_12174);
or U14407 (N_14407,N_12094,N_12005);
or U14408 (N_14408,N_12924,N_12101);
or U14409 (N_14409,N_13347,N_12915);
xnor U14410 (N_14410,N_12865,N_12455);
or U14411 (N_14411,N_13141,N_13251);
nand U14412 (N_14412,N_12301,N_12506);
nor U14413 (N_14413,N_12761,N_13381);
and U14414 (N_14414,N_12489,N_12172);
nand U14415 (N_14415,N_13211,N_13080);
nor U14416 (N_14416,N_12485,N_12459);
nor U14417 (N_14417,N_12460,N_12051);
nand U14418 (N_14418,N_13149,N_12693);
nor U14419 (N_14419,N_13344,N_12070);
and U14420 (N_14420,N_13445,N_12358);
xnor U14421 (N_14421,N_12181,N_12589);
nand U14422 (N_14422,N_13454,N_13127);
nand U14423 (N_14423,N_13029,N_12967);
nor U14424 (N_14424,N_12087,N_12402);
and U14425 (N_14425,N_12434,N_13216);
and U14426 (N_14426,N_12739,N_13234);
or U14427 (N_14427,N_13163,N_12521);
and U14428 (N_14428,N_13196,N_13263);
and U14429 (N_14429,N_12894,N_12023);
xnor U14430 (N_14430,N_12428,N_12418);
or U14431 (N_14431,N_12831,N_12483);
or U14432 (N_14432,N_13122,N_12568);
and U14433 (N_14433,N_12303,N_13253);
and U14434 (N_14434,N_13372,N_12771);
nor U14435 (N_14435,N_12362,N_13477);
nor U14436 (N_14436,N_12170,N_12993);
nor U14437 (N_14437,N_12822,N_13191);
nor U14438 (N_14438,N_12556,N_12471);
and U14439 (N_14439,N_13344,N_13244);
nor U14440 (N_14440,N_12395,N_13390);
or U14441 (N_14441,N_13373,N_12259);
xor U14442 (N_14442,N_13475,N_12657);
nand U14443 (N_14443,N_12932,N_12998);
nand U14444 (N_14444,N_13391,N_12736);
and U14445 (N_14445,N_12672,N_13182);
nand U14446 (N_14446,N_13052,N_12154);
and U14447 (N_14447,N_12173,N_12418);
or U14448 (N_14448,N_12711,N_12374);
and U14449 (N_14449,N_13232,N_13269);
and U14450 (N_14450,N_13493,N_12082);
or U14451 (N_14451,N_12911,N_12959);
xor U14452 (N_14452,N_12662,N_13119);
or U14453 (N_14453,N_13042,N_12020);
or U14454 (N_14454,N_12146,N_12236);
and U14455 (N_14455,N_12530,N_12533);
and U14456 (N_14456,N_12325,N_12954);
nand U14457 (N_14457,N_12126,N_12330);
nand U14458 (N_14458,N_12240,N_12789);
nand U14459 (N_14459,N_13244,N_12938);
and U14460 (N_14460,N_13166,N_12993);
and U14461 (N_14461,N_12190,N_13317);
and U14462 (N_14462,N_13478,N_12821);
and U14463 (N_14463,N_13494,N_12527);
nand U14464 (N_14464,N_12769,N_12231);
xnor U14465 (N_14465,N_12878,N_12263);
nand U14466 (N_14466,N_12556,N_12497);
and U14467 (N_14467,N_12264,N_12593);
or U14468 (N_14468,N_12737,N_12756);
nor U14469 (N_14469,N_13498,N_13031);
or U14470 (N_14470,N_12096,N_12012);
and U14471 (N_14471,N_13213,N_13359);
xor U14472 (N_14472,N_13401,N_12373);
and U14473 (N_14473,N_12114,N_13022);
and U14474 (N_14474,N_13359,N_12663);
nand U14475 (N_14475,N_13063,N_12048);
and U14476 (N_14476,N_12074,N_13469);
xnor U14477 (N_14477,N_13167,N_12470);
nand U14478 (N_14478,N_12207,N_12823);
xor U14479 (N_14479,N_12069,N_12241);
and U14480 (N_14480,N_12031,N_12010);
and U14481 (N_14481,N_12930,N_12235);
or U14482 (N_14482,N_13246,N_12450);
nor U14483 (N_14483,N_12635,N_12957);
xnor U14484 (N_14484,N_12239,N_12231);
xor U14485 (N_14485,N_12002,N_12480);
or U14486 (N_14486,N_12771,N_12797);
xnor U14487 (N_14487,N_13456,N_13422);
or U14488 (N_14488,N_12456,N_12125);
or U14489 (N_14489,N_13399,N_13448);
or U14490 (N_14490,N_13373,N_13399);
nor U14491 (N_14491,N_13058,N_12564);
nor U14492 (N_14492,N_12037,N_12532);
xor U14493 (N_14493,N_13325,N_12104);
nand U14494 (N_14494,N_12276,N_12874);
and U14495 (N_14495,N_12670,N_13467);
xor U14496 (N_14496,N_12443,N_12499);
or U14497 (N_14497,N_13091,N_12173);
or U14498 (N_14498,N_13226,N_12610);
nor U14499 (N_14499,N_12996,N_13102);
xor U14500 (N_14500,N_13176,N_12167);
or U14501 (N_14501,N_13085,N_12607);
and U14502 (N_14502,N_13438,N_12545);
xor U14503 (N_14503,N_12609,N_13055);
or U14504 (N_14504,N_12497,N_12883);
or U14505 (N_14505,N_13119,N_13071);
nand U14506 (N_14506,N_12048,N_12021);
nand U14507 (N_14507,N_13167,N_13458);
nand U14508 (N_14508,N_12495,N_12900);
and U14509 (N_14509,N_12574,N_12284);
nor U14510 (N_14510,N_12710,N_13057);
xnor U14511 (N_14511,N_12382,N_13275);
xor U14512 (N_14512,N_12924,N_12998);
nand U14513 (N_14513,N_12082,N_13211);
nand U14514 (N_14514,N_12747,N_12165);
nand U14515 (N_14515,N_13124,N_13071);
xor U14516 (N_14516,N_12081,N_12876);
xor U14517 (N_14517,N_12329,N_12080);
or U14518 (N_14518,N_12330,N_12589);
and U14519 (N_14519,N_12285,N_12236);
nor U14520 (N_14520,N_12028,N_12246);
or U14521 (N_14521,N_12744,N_12777);
nand U14522 (N_14522,N_12730,N_12569);
nand U14523 (N_14523,N_13436,N_12299);
xnor U14524 (N_14524,N_13491,N_13304);
and U14525 (N_14525,N_12830,N_12873);
nor U14526 (N_14526,N_12804,N_13109);
nand U14527 (N_14527,N_13219,N_12271);
nor U14528 (N_14528,N_12954,N_12592);
nor U14529 (N_14529,N_12135,N_13348);
and U14530 (N_14530,N_12034,N_12416);
or U14531 (N_14531,N_13012,N_12624);
and U14532 (N_14532,N_12434,N_13155);
or U14533 (N_14533,N_13433,N_13319);
or U14534 (N_14534,N_13221,N_13296);
nor U14535 (N_14535,N_13128,N_12506);
xor U14536 (N_14536,N_12833,N_12658);
nor U14537 (N_14537,N_12103,N_12510);
nand U14538 (N_14538,N_12594,N_12452);
and U14539 (N_14539,N_12783,N_12872);
or U14540 (N_14540,N_13419,N_12179);
xor U14541 (N_14541,N_13282,N_13174);
xor U14542 (N_14542,N_13309,N_12552);
and U14543 (N_14543,N_12018,N_12414);
or U14544 (N_14544,N_12495,N_12411);
nor U14545 (N_14545,N_12485,N_12940);
nand U14546 (N_14546,N_12789,N_12113);
xnor U14547 (N_14547,N_12811,N_12165);
and U14548 (N_14548,N_12880,N_12028);
nand U14549 (N_14549,N_12550,N_12154);
or U14550 (N_14550,N_12331,N_13374);
or U14551 (N_14551,N_12217,N_12663);
nand U14552 (N_14552,N_12443,N_12354);
nor U14553 (N_14553,N_12839,N_13127);
and U14554 (N_14554,N_13079,N_12184);
nand U14555 (N_14555,N_12336,N_12951);
xnor U14556 (N_14556,N_12162,N_12309);
xnor U14557 (N_14557,N_12084,N_12407);
nand U14558 (N_14558,N_12587,N_12946);
and U14559 (N_14559,N_12717,N_12963);
xnor U14560 (N_14560,N_13180,N_12241);
xor U14561 (N_14561,N_12441,N_13231);
xor U14562 (N_14562,N_13333,N_12751);
nor U14563 (N_14563,N_13238,N_12944);
nor U14564 (N_14564,N_13100,N_13488);
nand U14565 (N_14565,N_13367,N_13298);
or U14566 (N_14566,N_12918,N_12152);
nand U14567 (N_14567,N_12756,N_12640);
nand U14568 (N_14568,N_12353,N_12913);
and U14569 (N_14569,N_12511,N_13195);
nor U14570 (N_14570,N_12827,N_12997);
xnor U14571 (N_14571,N_12769,N_13259);
nand U14572 (N_14572,N_12699,N_12375);
xnor U14573 (N_14573,N_12954,N_13103);
and U14574 (N_14574,N_12386,N_12586);
or U14575 (N_14575,N_12216,N_12814);
nor U14576 (N_14576,N_12240,N_13253);
nand U14577 (N_14577,N_12353,N_12936);
xor U14578 (N_14578,N_13288,N_13022);
nand U14579 (N_14579,N_12933,N_12960);
or U14580 (N_14580,N_12232,N_12616);
or U14581 (N_14581,N_12356,N_12764);
and U14582 (N_14582,N_13261,N_12670);
nand U14583 (N_14583,N_12735,N_13152);
nand U14584 (N_14584,N_12862,N_12446);
nand U14585 (N_14585,N_12467,N_12931);
or U14586 (N_14586,N_12381,N_12949);
nand U14587 (N_14587,N_12402,N_12224);
xnor U14588 (N_14588,N_12759,N_12051);
nand U14589 (N_14589,N_12350,N_13089);
nor U14590 (N_14590,N_13415,N_12812);
and U14591 (N_14591,N_13210,N_12432);
nand U14592 (N_14592,N_12830,N_12069);
and U14593 (N_14593,N_12196,N_12366);
or U14594 (N_14594,N_13455,N_13332);
nor U14595 (N_14595,N_12058,N_13432);
nor U14596 (N_14596,N_13448,N_12281);
xnor U14597 (N_14597,N_13360,N_12392);
nand U14598 (N_14598,N_13128,N_12809);
nor U14599 (N_14599,N_12977,N_13224);
and U14600 (N_14600,N_12420,N_12009);
nand U14601 (N_14601,N_12851,N_12544);
nand U14602 (N_14602,N_12290,N_12705);
nor U14603 (N_14603,N_12276,N_12037);
and U14604 (N_14604,N_12097,N_13356);
nand U14605 (N_14605,N_12154,N_12480);
or U14606 (N_14606,N_12078,N_13279);
xnor U14607 (N_14607,N_12040,N_12806);
nor U14608 (N_14608,N_12994,N_13222);
and U14609 (N_14609,N_12090,N_13044);
xnor U14610 (N_14610,N_12906,N_12530);
nand U14611 (N_14611,N_12193,N_13345);
nand U14612 (N_14612,N_12345,N_13426);
or U14613 (N_14613,N_12794,N_12788);
or U14614 (N_14614,N_13392,N_13063);
nand U14615 (N_14615,N_12840,N_12710);
nor U14616 (N_14616,N_12776,N_13162);
nand U14617 (N_14617,N_12425,N_12006);
and U14618 (N_14618,N_12343,N_12853);
or U14619 (N_14619,N_13000,N_12945);
nor U14620 (N_14620,N_12833,N_12823);
nand U14621 (N_14621,N_12454,N_12048);
and U14622 (N_14622,N_13096,N_12117);
xnor U14623 (N_14623,N_12972,N_13275);
xor U14624 (N_14624,N_12026,N_13284);
and U14625 (N_14625,N_13022,N_12847);
and U14626 (N_14626,N_12853,N_13068);
nand U14627 (N_14627,N_13335,N_12639);
or U14628 (N_14628,N_12060,N_12454);
nand U14629 (N_14629,N_13223,N_12435);
and U14630 (N_14630,N_12126,N_13281);
nand U14631 (N_14631,N_12591,N_12129);
xnor U14632 (N_14632,N_12789,N_13106);
or U14633 (N_14633,N_12047,N_13488);
xor U14634 (N_14634,N_12423,N_13119);
xnor U14635 (N_14635,N_13411,N_13450);
nand U14636 (N_14636,N_12391,N_12255);
nand U14637 (N_14637,N_12812,N_12537);
or U14638 (N_14638,N_13244,N_12140);
nor U14639 (N_14639,N_13126,N_13321);
xor U14640 (N_14640,N_12280,N_12538);
nor U14641 (N_14641,N_12047,N_12304);
xor U14642 (N_14642,N_13401,N_12771);
xor U14643 (N_14643,N_12468,N_12816);
or U14644 (N_14644,N_12335,N_12529);
nor U14645 (N_14645,N_12541,N_12880);
nand U14646 (N_14646,N_12046,N_12215);
nor U14647 (N_14647,N_13451,N_12759);
and U14648 (N_14648,N_13108,N_12341);
xnor U14649 (N_14649,N_13157,N_12862);
xor U14650 (N_14650,N_13483,N_13384);
and U14651 (N_14651,N_13309,N_12123);
xor U14652 (N_14652,N_12693,N_12774);
xor U14653 (N_14653,N_12674,N_12789);
nand U14654 (N_14654,N_12088,N_13248);
nand U14655 (N_14655,N_12717,N_13495);
or U14656 (N_14656,N_13311,N_12301);
or U14657 (N_14657,N_12124,N_13155);
nand U14658 (N_14658,N_12666,N_12986);
and U14659 (N_14659,N_13103,N_12832);
xnor U14660 (N_14660,N_13380,N_12371);
or U14661 (N_14661,N_12973,N_12456);
and U14662 (N_14662,N_13158,N_12351);
and U14663 (N_14663,N_12453,N_12374);
nor U14664 (N_14664,N_13391,N_12316);
or U14665 (N_14665,N_13145,N_12268);
or U14666 (N_14666,N_12668,N_13014);
and U14667 (N_14667,N_12203,N_12621);
and U14668 (N_14668,N_13368,N_12878);
and U14669 (N_14669,N_12336,N_13133);
and U14670 (N_14670,N_12848,N_12607);
nor U14671 (N_14671,N_12942,N_12136);
or U14672 (N_14672,N_12636,N_12072);
or U14673 (N_14673,N_12952,N_12542);
and U14674 (N_14674,N_12526,N_13177);
nor U14675 (N_14675,N_12261,N_12502);
nand U14676 (N_14676,N_12073,N_12582);
nor U14677 (N_14677,N_13124,N_13377);
and U14678 (N_14678,N_13296,N_13188);
nor U14679 (N_14679,N_12469,N_13472);
xor U14680 (N_14680,N_12597,N_12471);
or U14681 (N_14681,N_12713,N_12953);
nand U14682 (N_14682,N_12233,N_13470);
nand U14683 (N_14683,N_12048,N_12457);
nand U14684 (N_14684,N_12875,N_12446);
and U14685 (N_14685,N_12196,N_12733);
and U14686 (N_14686,N_12473,N_12378);
or U14687 (N_14687,N_12819,N_12177);
nand U14688 (N_14688,N_13132,N_13355);
and U14689 (N_14689,N_13420,N_12271);
xor U14690 (N_14690,N_13253,N_13374);
nor U14691 (N_14691,N_12492,N_12814);
xor U14692 (N_14692,N_13470,N_12331);
nand U14693 (N_14693,N_13203,N_13358);
xnor U14694 (N_14694,N_13010,N_12707);
nand U14695 (N_14695,N_12088,N_12646);
nand U14696 (N_14696,N_13027,N_12294);
nand U14697 (N_14697,N_13087,N_12973);
or U14698 (N_14698,N_12464,N_13208);
and U14699 (N_14699,N_12219,N_12957);
xnor U14700 (N_14700,N_13267,N_12011);
nand U14701 (N_14701,N_12938,N_12826);
and U14702 (N_14702,N_12579,N_13034);
nand U14703 (N_14703,N_12179,N_12557);
or U14704 (N_14704,N_13385,N_12579);
xnor U14705 (N_14705,N_12940,N_12419);
nand U14706 (N_14706,N_13031,N_12926);
nand U14707 (N_14707,N_12370,N_12442);
nor U14708 (N_14708,N_12345,N_13190);
or U14709 (N_14709,N_12879,N_12062);
xnor U14710 (N_14710,N_12689,N_12092);
or U14711 (N_14711,N_13126,N_13075);
xor U14712 (N_14712,N_12205,N_13097);
xor U14713 (N_14713,N_13390,N_12408);
or U14714 (N_14714,N_12374,N_13209);
or U14715 (N_14715,N_12402,N_12926);
xor U14716 (N_14716,N_12964,N_13327);
or U14717 (N_14717,N_13436,N_12646);
and U14718 (N_14718,N_12065,N_12568);
nand U14719 (N_14719,N_12206,N_12289);
xnor U14720 (N_14720,N_12802,N_12956);
or U14721 (N_14721,N_12593,N_12476);
nand U14722 (N_14722,N_12050,N_12660);
or U14723 (N_14723,N_13270,N_12199);
nor U14724 (N_14724,N_12354,N_12551);
nand U14725 (N_14725,N_12649,N_13496);
nor U14726 (N_14726,N_12031,N_13059);
nor U14727 (N_14727,N_12132,N_12344);
or U14728 (N_14728,N_12754,N_13194);
nor U14729 (N_14729,N_13442,N_13263);
and U14730 (N_14730,N_12715,N_12814);
or U14731 (N_14731,N_12553,N_12385);
nor U14732 (N_14732,N_13378,N_12581);
nand U14733 (N_14733,N_13301,N_12802);
xnor U14734 (N_14734,N_12819,N_12505);
nor U14735 (N_14735,N_12865,N_13100);
nand U14736 (N_14736,N_13069,N_13389);
and U14737 (N_14737,N_13358,N_12376);
nor U14738 (N_14738,N_12543,N_13365);
and U14739 (N_14739,N_12250,N_12180);
and U14740 (N_14740,N_12691,N_12286);
xnor U14741 (N_14741,N_12391,N_12156);
or U14742 (N_14742,N_12299,N_12694);
or U14743 (N_14743,N_12812,N_12940);
or U14744 (N_14744,N_13305,N_12292);
and U14745 (N_14745,N_13459,N_12890);
xnor U14746 (N_14746,N_12899,N_12171);
or U14747 (N_14747,N_12666,N_12969);
and U14748 (N_14748,N_12806,N_12924);
and U14749 (N_14749,N_12350,N_13111);
and U14750 (N_14750,N_12007,N_12086);
nand U14751 (N_14751,N_12208,N_13182);
nor U14752 (N_14752,N_13002,N_12481);
xnor U14753 (N_14753,N_12202,N_12826);
or U14754 (N_14754,N_13004,N_12754);
nor U14755 (N_14755,N_12605,N_12091);
and U14756 (N_14756,N_12615,N_12500);
nor U14757 (N_14757,N_12312,N_13239);
and U14758 (N_14758,N_12787,N_12426);
or U14759 (N_14759,N_12457,N_12387);
nand U14760 (N_14760,N_13289,N_12944);
nand U14761 (N_14761,N_13140,N_12397);
nand U14762 (N_14762,N_13209,N_13258);
nand U14763 (N_14763,N_13026,N_12863);
nor U14764 (N_14764,N_12936,N_13178);
and U14765 (N_14765,N_12199,N_12836);
and U14766 (N_14766,N_12978,N_13082);
xor U14767 (N_14767,N_13471,N_12608);
and U14768 (N_14768,N_13413,N_12306);
nor U14769 (N_14769,N_13126,N_13041);
and U14770 (N_14770,N_12290,N_12054);
nor U14771 (N_14771,N_13033,N_12016);
nor U14772 (N_14772,N_12675,N_13107);
nand U14773 (N_14773,N_13194,N_12895);
nor U14774 (N_14774,N_12690,N_12724);
nor U14775 (N_14775,N_12768,N_13455);
or U14776 (N_14776,N_13274,N_12070);
and U14777 (N_14777,N_12016,N_12957);
xor U14778 (N_14778,N_12767,N_13400);
nand U14779 (N_14779,N_13384,N_13018);
nand U14780 (N_14780,N_12474,N_12903);
and U14781 (N_14781,N_12097,N_12771);
nand U14782 (N_14782,N_12956,N_12243);
or U14783 (N_14783,N_12996,N_13469);
nor U14784 (N_14784,N_13468,N_12779);
nand U14785 (N_14785,N_12115,N_12569);
xor U14786 (N_14786,N_12114,N_12951);
nand U14787 (N_14787,N_12551,N_12765);
xnor U14788 (N_14788,N_12761,N_13447);
nor U14789 (N_14789,N_13369,N_13135);
nand U14790 (N_14790,N_13081,N_12924);
nand U14791 (N_14791,N_12900,N_12438);
nor U14792 (N_14792,N_12117,N_12703);
nor U14793 (N_14793,N_12485,N_12294);
and U14794 (N_14794,N_12432,N_13143);
nor U14795 (N_14795,N_13469,N_12270);
and U14796 (N_14796,N_12117,N_12730);
nor U14797 (N_14797,N_12192,N_12718);
nand U14798 (N_14798,N_13007,N_13120);
xnor U14799 (N_14799,N_12940,N_12499);
or U14800 (N_14800,N_12041,N_13327);
and U14801 (N_14801,N_13478,N_12524);
nand U14802 (N_14802,N_12073,N_12444);
nor U14803 (N_14803,N_12288,N_12458);
nand U14804 (N_14804,N_12345,N_13056);
nand U14805 (N_14805,N_12006,N_13454);
nor U14806 (N_14806,N_13215,N_13116);
nand U14807 (N_14807,N_13002,N_13372);
or U14808 (N_14808,N_12969,N_12601);
nor U14809 (N_14809,N_13460,N_12968);
or U14810 (N_14810,N_13300,N_12039);
nand U14811 (N_14811,N_13424,N_12536);
nand U14812 (N_14812,N_12862,N_13310);
nand U14813 (N_14813,N_12216,N_12397);
nor U14814 (N_14814,N_12634,N_12322);
or U14815 (N_14815,N_13454,N_12078);
xnor U14816 (N_14816,N_12723,N_13162);
and U14817 (N_14817,N_13281,N_12021);
nor U14818 (N_14818,N_12571,N_13198);
and U14819 (N_14819,N_12310,N_12264);
nor U14820 (N_14820,N_12619,N_12532);
and U14821 (N_14821,N_12788,N_12611);
xor U14822 (N_14822,N_13367,N_12173);
nand U14823 (N_14823,N_12487,N_12970);
and U14824 (N_14824,N_12658,N_12060);
and U14825 (N_14825,N_13062,N_12173);
or U14826 (N_14826,N_13191,N_12296);
and U14827 (N_14827,N_12268,N_12933);
or U14828 (N_14828,N_12241,N_12469);
or U14829 (N_14829,N_12150,N_12848);
and U14830 (N_14830,N_12648,N_12159);
or U14831 (N_14831,N_12551,N_12838);
xnor U14832 (N_14832,N_13006,N_13034);
and U14833 (N_14833,N_12194,N_12935);
nand U14834 (N_14834,N_13008,N_12517);
nor U14835 (N_14835,N_12683,N_12680);
and U14836 (N_14836,N_13241,N_12652);
nor U14837 (N_14837,N_13308,N_12495);
xnor U14838 (N_14838,N_13159,N_12133);
or U14839 (N_14839,N_13461,N_12338);
nand U14840 (N_14840,N_12364,N_12651);
or U14841 (N_14841,N_12005,N_12346);
xor U14842 (N_14842,N_12844,N_12007);
xor U14843 (N_14843,N_12240,N_12178);
and U14844 (N_14844,N_12035,N_12882);
and U14845 (N_14845,N_13027,N_13283);
xnor U14846 (N_14846,N_12173,N_13089);
and U14847 (N_14847,N_12390,N_12621);
nor U14848 (N_14848,N_13166,N_12005);
or U14849 (N_14849,N_12720,N_12850);
nor U14850 (N_14850,N_12529,N_12513);
and U14851 (N_14851,N_12786,N_12620);
xnor U14852 (N_14852,N_12872,N_12430);
nor U14853 (N_14853,N_13287,N_12347);
xnor U14854 (N_14854,N_13245,N_13387);
xnor U14855 (N_14855,N_12642,N_12632);
nand U14856 (N_14856,N_13017,N_13126);
and U14857 (N_14857,N_12168,N_13323);
nor U14858 (N_14858,N_12520,N_13209);
xor U14859 (N_14859,N_12993,N_12798);
and U14860 (N_14860,N_12799,N_12023);
nor U14861 (N_14861,N_13039,N_12156);
nor U14862 (N_14862,N_12578,N_12446);
or U14863 (N_14863,N_12127,N_12310);
nand U14864 (N_14864,N_13015,N_12503);
and U14865 (N_14865,N_13052,N_12117);
and U14866 (N_14866,N_12856,N_13312);
nor U14867 (N_14867,N_12491,N_13253);
xor U14868 (N_14868,N_12184,N_13467);
and U14869 (N_14869,N_12602,N_12404);
nor U14870 (N_14870,N_12092,N_12779);
and U14871 (N_14871,N_13428,N_13296);
nand U14872 (N_14872,N_12269,N_12505);
nand U14873 (N_14873,N_13074,N_12495);
or U14874 (N_14874,N_13072,N_12920);
xnor U14875 (N_14875,N_13124,N_12484);
or U14876 (N_14876,N_12353,N_13281);
nand U14877 (N_14877,N_13033,N_13369);
xor U14878 (N_14878,N_12478,N_13363);
nor U14879 (N_14879,N_13375,N_12687);
or U14880 (N_14880,N_12618,N_12163);
or U14881 (N_14881,N_12681,N_12558);
nand U14882 (N_14882,N_12865,N_12917);
nand U14883 (N_14883,N_12040,N_12322);
nand U14884 (N_14884,N_12487,N_13455);
and U14885 (N_14885,N_12195,N_12242);
and U14886 (N_14886,N_12544,N_13046);
nand U14887 (N_14887,N_13053,N_12265);
and U14888 (N_14888,N_12075,N_12304);
and U14889 (N_14889,N_12303,N_12266);
nor U14890 (N_14890,N_13303,N_12252);
nand U14891 (N_14891,N_13491,N_12169);
nand U14892 (N_14892,N_13057,N_12591);
nand U14893 (N_14893,N_12211,N_12814);
nor U14894 (N_14894,N_13171,N_12119);
nand U14895 (N_14895,N_13461,N_12506);
nand U14896 (N_14896,N_12737,N_12223);
or U14897 (N_14897,N_12223,N_12310);
and U14898 (N_14898,N_12957,N_12174);
or U14899 (N_14899,N_12909,N_12780);
or U14900 (N_14900,N_12483,N_12767);
and U14901 (N_14901,N_12731,N_13283);
nor U14902 (N_14902,N_12543,N_12317);
nand U14903 (N_14903,N_13300,N_13217);
nor U14904 (N_14904,N_12497,N_12291);
xor U14905 (N_14905,N_12468,N_12875);
nor U14906 (N_14906,N_13241,N_12871);
nor U14907 (N_14907,N_13340,N_13108);
nand U14908 (N_14908,N_12366,N_12888);
nor U14909 (N_14909,N_12575,N_12882);
nand U14910 (N_14910,N_13055,N_12686);
nand U14911 (N_14911,N_12191,N_13463);
xnor U14912 (N_14912,N_12256,N_13309);
or U14913 (N_14913,N_12738,N_13107);
or U14914 (N_14914,N_12982,N_13115);
xor U14915 (N_14915,N_13438,N_12428);
or U14916 (N_14916,N_13387,N_13325);
nor U14917 (N_14917,N_13114,N_12542);
and U14918 (N_14918,N_12121,N_13244);
nor U14919 (N_14919,N_12288,N_12160);
nor U14920 (N_14920,N_12942,N_12672);
nand U14921 (N_14921,N_12080,N_12954);
and U14922 (N_14922,N_13227,N_12606);
or U14923 (N_14923,N_12458,N_12178);
xor U14924 (N_14924,N_13422,N_12572);
and U14925 (N_14925,N_12561,N_13347);
and U14926 (N_14926,N_12240,N_12448);
or U14927 (N_14927,N_12350,N_12655);
or U14928 (N_14928,N_12907,N_13193);
and U14929 (N_14929,N_12170,N_13398);
nor U14930 (N_14930,N_12747,N_12754);
and U14931 (N_14931,N_12440,N_13143);
and U14932 (N_14932,N_12517,N_12475);
nor U14933 (N_14933,N_12168,N_13269);
nand U14934 (N_14934,N_13156,N_13237);
nor U14935 (N_14935,N_13486,N_13465);
or U14936 (N_14936,N_12917,N_13202);
nand U14937 (N_14937,N_12226,N_12638);
xnor U14938 (N_14938,N_13169,N_12002);
nor U14939 (N_14939,N_12117,N_13087);
nor U14940 (N_14940,N_12386,N_13055);
and U14941 (N_14941,N_13414,N_12266);
and U14942 (N_14942,N_12115,N_13404);
xnor U14943 (N_14943,N_12375,N_12568);
xnor U14944 (N_14944,N_12109,N_13145);
or U14945 (N_14945,N_12836,N_13036);
xnor U14946 (N_14946,N_12454,N_13400);
nor U14947 (N_14947,N_13152,N_13027);
xor U14948 (N_14948,N_13020,N_12915);
xnor U14949 (N_14949,N_12298,N_12825);
nand U14950 (N_14950,N_12020,N_12493);
nor U14951 (N_14951,N_13414,N_12711);
xor U14952 (N_14952,N_13310,N_12560);
xnor U14953 (N_14953,N_12651,N_12332);
nor U14954 (N_14954,N_13474,N_12679);
and U14955 (N_14955,N_13394,N_12307);
xor U14956 (N_14956,N_12395,N_12097);
xor U14957 (N_14957,N_13247,N_12514);
xor U14958 (N_14958,N_13299,N_12398);
and U14959 (N_14959,N_12970,N_12149);
and U14960 (N_14960,N_12688,N_13206);
or U14961 (N_14961,N_12600,N_13011);
nor U14962 (N_14962,N_12396,N_12449);
xor U14963 (N_14963,N_12421,N_12162);
nand U14964 (N_14964,N_12674,N_12616);
nand U14965 (N_14965,N_13315,N_13305);
xor U14966 (N_14966,N_13153,N_13144);
and U14967 (N_14967,N_12504,N_12998);
xor U14968 (N_14968,N_12084,N_12065);
and U14969 (N_14969,N_12641,N_13382);
nor U14970 (N_14970,N_12504,N_12051);
and U14971 (N_14971,N_13120,N_12812);
and U14972 (N_14972,N_12794,N_12258);
or U14973 (N_14973,N_13310,N_12733);
nor U14974 (N_14974,N_12631,N_12948);
and U14975 (N_14975,N_12404,N_12519);
xnor U14976 (N_14976,N_13387,N_13473);
nor U14977 (N_14977,N_12330,N_12577);
xnor U14978 (N_14978,N_12529,N_12988);
xor U14979 (N_14979,N_13283,N_12922);
nor U14980 (N_14980,N_12795,N_12069);
xor U14981 (N_14981,N_13340,N_13370);
or U14982 (N_14982,N_12489,N_13373);
nor U14983 (N_14983,N_12817,N_12366);
nor U14984 (N_14984,N_13337,N_12741);
nand U14985 (N_14985,N_12314,N_12345);
xnor U14986 (N_14986,N_13013,N_12665);
xnor U14987 (N_14987,N_12827,N_12602);
nand U14988 (N_14988,N_12990,N_13236);
nand U14989 (N_14989,N_12848,N_13040);
and U14990 (N_14990,N_13176,N_12409);
xor U14991 (N_14991,N_13290,N_12065);
xnor U14992 (N_14992,N_12636,N_13387);
nor U14993 (N_14993,N_12927,N_12266);
nor U14994 (N_14994,N_12637,N_12574);
nand U14995 (N_14995,N_12666,N_12215);
nor U14996 (N_14996,N_13239,N_12658);
nand U14997 (N_14997,N_12769,N_13039);
nand U14998 (N_14998,N_12460,N_13019);
xnor U14999 (N_14999,N_12646,N_12958);
xor U15000 (N_15000,N_14127,N_14721);
xnor U15001 (N_15001,N_13978,N_13748);
and U15002 (N_15002,N_14468,N_14068);
and U15003 (N_15003,N_14602,N_14409);
and U15004 (N_15004,N_13618,N_14508);
xor U15005 (N_15005,N_13865,N_14199);
or U15006 (N_15006,N_14330,N_13859);
nand U15007 (N_15007,N_14911,N_14306);
and U15008 (N_15008,N_14170,N_13598);
or U15009 (N_15009,N_14537,N_14646);
nand U15010 (N_15010,N_14975,N_14805);
and U15011 (N_15011,N_14279,N_14774);
xor U15012 (N_15012,N_13746,N_14828);
or U15013 (N_15013,N_13557,N_13797);
or U15014 (N_15014,N_14801,N_14533);
nand U15015 (N_15015,N_14981,N_14147);
nor U15016 (N_15016,N_14861,N_14006);
nand U15017 (N_15017,N_13632,N_14315);
nand U15018 (N_15018,N_14386,N_14282);
nand U15019 (N_15019,N_14806,N_14344);
nor U15020 (N_15020,N_14091,N_14361);
or U15021 (N_15021,N_13884,N_14454);
or U15022 (N_15022,N_13585,N_14631);
nor U15023 (N_15023,N_13900,N_14848);
or U15024 (N_15024,N_14613,N_14335);
or U15025 (N_15025,N_13868,N_14145);
nand U15026 (N_15026,N_14957,N_13801);
and U15027 (N_15027,N_14519,N_14162);
nor U15028 (N_15028,N_13812,N_14615);
nor U15029 (N_15029,N_14525,N_14994);
xor U15030 (N_15030,N_14466,N_13969);
nor U15031 (N_15031,N_14870,N_14134);
nand U15032 (N_15032,N_14191,N_14835);
xor U15033 (N_15033,N_14484,N_13916);
nand U15034 (N_15034,N_14236,N_14844);
and U15035 (N_15035,N_13661,N_14363);
xnor U15036 (N_15036,N_13860,N_14657);
nand U15037 (N_15037,N_14651,N_14252);
and U15038 (N_15038,N_13780,N_14637);
nand U15039 (N_15039,N_14942,N_14624);
nand U15040 (N_15040,N_14024,N_14211);
nor U15041 (N_15041,N_14836,N_14784);
or U15042 (N_15042,N_14207,N_14966);
nand U15043 (N_15043,N_14338,N_14909);
nand U15044 (N_15044,N_14316,N_14218);
xnor U15045 (N_15045,N_13994,N_13825);
xor U15046 (N_15046,N_13712,N_13663);
xnor U15047 (N_15047,N_13941,N_13891);
nor U15048 (N_15048,N_13711,N_13533);
xnor U15049 (N_15049,N_14952,N_14358);
xor U15050 (N_15050,N_14810,N_14062);
or U15051 (N_15051,N_13814,N_14877);
or U15052 (N_15052,N_13788,N_14736);
or U15053 (N_15053,N_14665,N_13658);
nand U15054 (N_15054,N_14054,N_14532);
xor U15055 (N_15055,N_13959,N_14716);
xnor U15056 (N_15056,N_13875,N_13699);
or U15057 (N_15057,N_13953,N_14635);
and U15058 (N_15058,N_13521,N_14057);
xor U15059 (N_15059,N_14827,N_14572);
xnor U15060 (N_15060,N_14056,N_13680);
xnor U15061 (N_15061,N_14895,N_13623);
nor U15062 (N_15062,N_14822,N_14689);
or U15063 (N_15063,N_14460,N_14408);
and U15064 (N_15064,N_13731,N_13727);
xor U15065 (N_15065,N_14186,N_13792);
and U15066 (N_15066,N_13958,N_14198);
xor U15067 (N_15067,N_14729,N_14132);
nand U15068 (N_15068,N_14833,N_14890);
or U15069 (N_15069,N_14115,N_14259);
or U15070 (N_15070,N_13595,N_13781);
and U15071 (N_15071,N_14340,N_14770);
nor U15072 (N_15072,N_14766,N_13744);
nor U15073 (N_15073,N_13582,N_13679);
or U15074 (N_15074,N_14286,N_14712);
nor U15075 (N_15075,N_13576,N_13614);
or U15076 (N_15076,N_14217,N_13855);
nand U15077 (N_15077,N_14791,N_13822);
xor U15078 (N_15078,N_14742,N_14333);
and U15079 (N_15079,N_14552,N_14104);
xnor U15080 (N_15080,N_14595,N_14061);
or U15081 (N_15081,N_14244,N_13904);
or U15082 (N_15082,N_14432,N_14510);
nor U15083 (N_15083,N_14593,N_14254);
and U15084 (N_15084,N_14448,N_13724);
or U15085 (N_15085,N_14906,N_14824);
nor U15086 (N_15086,N_14893,N_13827);
nor U15087 (N_15087,N_13560,N_14083);
nor U15088 (N_15088,N_14167,N_14264);
or U15089 (N_15089,N_13730,N_14314);
xor U15090 (N_15090,N_13654,N_14714);
nor U15091 (N_15091,N_14856,N_14782);
and U15092 (N_15092,N_13615,N_14123);
xor U15093 (N_15093,N_14853,N_14171);
nor U15094 (N_15094,N_14417,N_14165);
and U15095 (N_15095,N_14614,N_13723);
or U15096 (N_15096,N_14379,N_14487);
or U15097 (N_15097,N_13770,N_14378);
nor U15098 (N_15098,N_14430,N_14859);
and U15099 (N_15099,N_13688,N_13807);
and U15100 (N_15100,N_14415,N_14079);
or U15101 (N_15101,N_14087,N_14028);
or U15102 (N_15102,N_14747,N_13698);
or U15103 (N_15103,N_14385,N_14016);
nand U15104 (N_15104,N_13898,N_13503);
nor U15105 (N_15105,N_13539,N_13913);
and U15106 (N_15106,N_13725,N_13518);
or U15107 (N_15107,N_14954,N_13504);
and U15108 (N_15108,N_14265,N_14871);
and U15109 (N_15109,N_14857,N_14985);
or U15110 (N_15110,N_13877,N_14494);
xnor U15111 (N_15111,N_13774,N_13776);
or U15112 (N_15112,N_14888,N_14974);
and U15113 (N_15113,N_14462,N_14339);
nand U15114 (N_15114,N_13640,N_14464);
xor U15115 (N_15115,N_14040,N_14045);
xnor U15116 (N_15116,N_14809,N_14804);
nor U15117 (N_15117,N_14281,N_13753);
and U15118 (N_15118,N_14310,N_14089);
nor U15119 (N_15119,N_14013,N_14880);
and U15120 (N_15120,N_14023,N_14032);
nand U15121 (N_15121,N_14991,N_14029);
nand U15122 (N_15122,N_13667,N_13785);
nand U15123 (N_15123,N_13506,N_14192);
nand U15124 (N_15124,N_14958,N_13851);
and U15125 (N_15125,N_14564,N_13512);
nor U15126 (N_15126,N_14908,N_14493);
and U15127 (N_15127,N_13649,N_13988);
xor U15128 (N_15128,N_13756,N_13659);
xnor U15129 (N_15129,N_14465,N_14507);
xnor U15130 (N_15130,N_13972,N_14148);
or U15131 (N_15131,N_13968,N_14458);
or U15132 (N_15132,N_14597,N_14256);
or U15133 (N_15133,N_14577,N_14461);
nor U15134 (N_15134,N_13519,N_13980);
nor U15135 (N_15135,N_13566,N_13951);
nor U15136 (N_15136,N_14422,N_13786);
or U15137 (N_15137,N_13713,N_13752);
nand U15138 (N_15138,N_14195,N_13960);
xor U15139 (N_15139,N_14977,N_13908);
nor U15140 (N_15140,N_14661,N_14154);
or U15141 (N_15141,N_14072,N_14868);
or U15142 (N_15142,N_14001,N_13709);
xor U15143 (N_15143,N_14578,N_14108);
nor U15144 (N_15144,N_14764,N_14321);
xor U15145 (N_15145,N_13772,N_13849);
or U15146 (N_15146,N_14247,N_14299);
and U15147 (N_15147,N_14730,N_13665);
nor U15148 (N_15148,N_13981,N_14753);
or U15149 (N_15149,N_13845,N_14584);
xor U15150 (N_15150,N_13842,N_14400);
nand U15151 (N_15151,N_14190,N_14085);
nand U15152 (N_15152,N_14049,N_14768);
and U15153 (N_15153,N_13601,N_13630);
nand U15154 (N_15154,N_14092,N_13769);
and U15155 (N_15155,N_14086,N_13929);
or U15156 (N_15156,N_14727,N_14803);
nand U15157 (N_15157,N_14122,N_14926);
nand U15158 (N_15158,N_14864,N_14622);
nor U15159 (N_15159,N_14421,N_14093);
nand U15160 (N_15160,N_14555,N_13500);
xor U15161 (N_15161,N_13992,N_14542);
xnor U15162 (N_15162,N_14825,N_14869);
xor U15163 (N_15163,N_13950,N_14955);
and U15164 (N_15164,N_13826,N_13626);
and U15165 (N_15165,N_14474,N_13743);
or U15166 (N_15166,N_13973,N_14326);
nand U15167 (N_15167,N_13570,N_13655);
nor U15168 (N_15168,N_14617,N_14371);
nand U15169 (N_15169,N_14808,N_14639);
and U15170 (N_15170,N_13672,N_13926);
nor U15171 (N_15171,N_14664,N_13998);
or U15172 (N_15172,N_13502,N_14566);
and U15173 (N_15173,N_14789,N_14188);
xnor U15174 (N_15174,N_13946,N_14775);
or U15175 (N_15175,N_14343,N_13841);
xnor U15176 (N_15176,N_13810,N_14963);
xor U15177 (N_15177,N_13754,N_14969);
or U15178 (N_15178,N_14875,N_14823);
nor U15179 (N_15179,N_14680,N_13811);
or U15180 (N_15180,N_13757,N_13952);
xor U15181 (N_15181,N_14523,N_14457);
nand U15182 (N_15182,N_13983,N_14722);
xnor U15183 (N_15183,N_13840,N_14696);
nand U15184 (N_15184,N_14036,N_13915);
or U15185 (N_15185,N_13603,N_14773);
or U15186 (N_15186,N_13599,N_14200);
or U15187 (N_15187,N_14155,N_13716);
xor U15188 (N_15188,N_14075,N_13629);
xor U15189 (N_15189,N_14887,N_14368);
xnor U15190 (N_15190,N_14435,N_14944);
nand U15191 (N_15191,N_14241,N_14351);
nand U15192 (N_15192,N_14724,N_13578);
and U15193 (N_15193,N_14682,N_13580);
or U15194 (N_15194,N_14705,N_14130);
or U15195 (N_15195,N_14360,N_13828);
nand U15196 (N_15196,N_14142,N_14874);
nor U15197 (N_15197,N_14129,N_14272);
and U15198 (N_15198,N_13948,N_13821);
and U15199 (N_15199,N_14546,N_13676);
and U15200 (N_15200,N_14238,N_14488);
xor U15201 (N_15201,N_14173,N_14348);
or U15202 (N_15202,N_14703,N_13925);
xnor U15203 (N_15203,N_14139,N_14568);
nor U15204 (N_15204,N_14711,N_13571);
nand U15205 (N_15205,N_14674,N_14972);
nor U15206 (N_15206,N_14596,N_13871);
nor U15207 (N_15207,N_13600,N_14081);
xnor U15208 (N_15208,N_14399,N_14224);
nand U15209 (N_15209,N_14976,N_14381);
nand U15210 (N_15210,N_13848,N_14878);
nor U15211 (N_15211,N_13954,N_13525);
nand U15212 (N_15212,N_14425,N_14169);
nand U15213 (N_15213,N_14756,N_14755);
or U15214 (N_15214,N_14166,N_14373);
and U15215 (N_15215,N_13516,N_14492);
or U15216 (N_15216,N_14838,N_14387);
nand U15217 (N_15217,N_13717,N_13761);
nand U15218 (N_15218,N_13540,N_14987);
and U15219 (N_15219,N_14504,N_13509);
xor U15220 (N_15220,N_14565,N_14485);
nor U15221 (N_15221,N_14688,N_13588);
xnor U15222 (N_15222,N_14133,N_13764);
and U15223 (N_15223,N_13760,N_14496);
xor U15224 (N_15224,N_14196,N_14411);
nor U15225 (N_15225,N_14959,N_14126);
or U15226 (N_15226,N_14815,N_13933);
xnor U15227 (N_15227,N_14796,N_14209);
xnor U15228 (N_15228,N_13616,N_14495);
xor U15229 (N_15229,N_14915,N_14284);
and U15230 (N_15230,N_14843,N_13837);
or U15231 (N_15231,N_14881,N_13847);
xor U15232 (N_15232,N_14841,N_14151);
and U15233 (N_15233,N_14106,N_14135);
or U15234 (N_15234,N_14189,N_13895);
xnor U15235 (N_15235,N_13642,N_13624);
xor U15236 (N_15236,N_14840,N_14516);
nand U15237 (N_15237,N_14051,N_13647);
nor U15238 (N_15238,N_14660,N_14372);
xor U15239 (N_15239,N_13873,N_13685);
nor U15240 (N_15240,N_14066,N_14471);
xnor U15241 (N_15241,N_14929,N_14772);
and U15242 (N_15242,N_14158,N_14228);
xor U15243 (N_15243,N_14512,N_14301);
nor U15244 (N_15244,N_14459,N_14786);
nand U15245 (N_15245,N_14502,N_14852);
and U15246 (N_15246,N_14745,N_14011);
nand U15247 (N_15247,N_14862,N_14754);
and U15248 (N_15248,N_13902,N_14102);
or U15249 (N_15249,N_14992,N_14490);
or U15250 (N_15250,N_14978,N_14594);
nor U15251 (N_15251,N_14666,N_14118);
xnor U15252 (N_15252,N_14744,N_13707);
nand U15253 (N_15253,N_13886,N_13579);
nor U15254 (N_15254,N_14033,N_13613);
nor U15255 (N_15255,N_14788,N_14395);
nand U15256 (N_15256,N_14563,N_14047);
and U15257 (N_15257,N_14912,N_13681);
nor U15258 (N_15258,N_14034,N_13638);
or U15259 (N_15259,N_14900,N_13894);
nand U15260 (N_15260,N_14500,N_14821);
nor U15261 (N_15261,N_14947,N_14860);
nand U15262 (N_15262,N_13735,N_14936);
nand U15263 (N_15263,N_14832,N_14866);
nand U15264 (N_15264,N_13664,N_14463);
nor U15265 (N_15265,N_14365,N_14026);
nor U15266 (N_15266,N_14076,N_14609);
nand U15267 (N_15267,N_14573,N_14226);
nor U15268 (N_15268,N_13870,N_13920);
and U15269 (N_15269,N_13550,N_14305);
xnor U15270 (N_15270,N_13574,N_14554);
or U15271 (N_15271,N_14020,N_14867);
nor U15272 (N_15272,N_13700,N_14579);
and U15273 (N_15273,N_14585,N_14748);
nand U15274 (N_15274,N_13892,N_14090);
or U15275 (N_15275,N_13543,N_14433);
xor U15276 (N_15276,N_14670,N_13936);
nand U15277 (N_15277,N_13921,N_14356);
or U15278 (N_15278,N_13893,N_14948);
xnor U15279 (N_15279,N_14232,N_14181);
and U15280 (N_15280,N_14873,N_13697);
or U15281 (N_15281,N_14476,N_14826);
xnor U15282 (N_15282,N_14644,N_14658);
and U15283 (N_15283,N_13721,N_14923);
nor U15284 (N_15284,N_14248,N_13701);
or U15285 (N_15285,N_13888,N_13612);
nor U15286 (N_15286,N_14675,N_14312);
nand U15287 (N_15287,N_13912,N_14920);
and U15288 (N_15288,N_14479,N_14964);
nand U15289 (N_15289,N_13985,N_14116);
xor U15290 (N_15290,N_14048,N_14851);
nand U15291 (N_15291,N_14928,N_14113);
and U15292 (N_15292,N_14612,N_14679);
nand U15293 (N_15293,N_14019,N_14777);
and U15294 (N_15294,N_13971,N_13702);
xnor U15295 (N_15295,N_14800,N_14634);
and U15296 (N_15296,N_13534,N_14831);
xor U15297 (N_15297,N_14550,N_13937);
nand U15298 (N_15298,N_14121,N_14879);
nand U15299 (N_15299,N_14478,N_13947);
xnor U15300 (N_15300,N_13621,N_13651);
nand U15301 (N_15301,N_13779,N_14710);
nor U15302 (N_15302,N_13800,N_14416);
xor U15303 (N_15303,N_14213,N_13634);
nor U15304 (N_15304,N_13819,N_13787);
nor U15305 (N_15305,N_14038,N_14491);
and U15306 (N_15306,N_14561,N_14337);
xor U15307 (N_15307,N_14998,N_14790);
nand U15308 (N_15308,N_14009,N_14961);
or U15309 (N_15309,N_14349,N_14497);
nor U15310 (N_15310,N_14277,N_13989);
and U15311 (N_15311,N_14600,N_14184);
or U15312 (N_15312,N_14010,N_14898);
or U15313 (N_15313,N_14536,N_14776);
and U15314 (N_15314,N_13637,N_14088);
xnor U15315 (N_15315,N_13962,N_14761);
nand U15316 (N_15316,N_13899,N_14683);
nor U15317 (N_15317,N_14896,N_14341);
nor U15318 (N_15318,N_14640,N_14642);
xnor U15319 (N_15319,N_14146,N_14979);
nor U15320 (N_15320,N_13949,N_13965);
nand U15321 (N_15321,N_14551,N_13817);
and U15322 (N_15322,N_14545,N_14424);
or U15323 (N_15323,N_14672,N_14787);
or U15324 (N_15324,N_14302,N_14164);
nor U15325 (N_15325,N_13690,N_13706);
nand U15326 (N_15326,N_14380,N_14903);
nor U15327 (N_15327,N_14230,N_14541);
or U15328 (N_15328,N_14074,N_14183);
or U15329 (N_15329,N_14509,N_14390);
or U15330 (N_15330,N_14935,N_14785);
and U15331 (N_15331,N_14517,N_14287);
or U15332 (N_15332,N_14261,N_14111);
and U15333 (N_15333,N_14222,N_14726);
nor U15334 (N_15334,N_14918,N_14863);
or U15335 (N_15335,N_14697,N_14534);
nand U15336 (N_15336,N_14280,N_13832);
nor U15337 (N_15337,N_14819,N_14515);
and U15338 (N_15338,N_13589,N_14160);
xnor U15339 (N_15339,N_14663,N_14289);
and U15340 (N_15340,N_14233,N_14353);
or U15341 (N_15341,N_14950,N_13556);
or U15342 (N_15342,N_13793,N_13631);
xor U15343 (N_15343,N_13695,N_13656);
nor U15344 (N_15344,N_14673,N_14447);
and U15345 (N_15345,N_14253,N_13704);
xor U15346 (N_15346,N_14669,N_13719);
nand U15347 (N_15347,N_14701,N_14441);
nand U15348 (N_15348,N_14505,N_13545);
or U15349 (N_15349,N_14520,N_14706);
nor U15350 (N_15350,N_14237,N_14262);
nor U15351 (N_15351,N_14778,N_13565);
nand U15352 (N_15352,N_14275,N_14293);
and U15353 (N_15353,N_14625,N_14535);
xnor U15354 (N_15354,N_13522,N_14548);
nor U15355 (N_15355,N_14499,N_14807);
or U15356 (N_15356,N_14168,N_14098);
nor U15357 (N_15357,N_14452,N_13869);
or U15358 (N_15358,N_14197,N_14694);
nand U15359 (N_15359,N_14374,N_14608);
nor U15360 (N_15360,N_13955,N_14014);
xor U15361 (N_15361,N_14728,N_14932);
nor U15362 (N_15362,N_14205,N_14375);
or U15363 (N_15363,N_13586,N_13677);
nor U15364 (N_15364,N_14910,N_13741);
nor U15365 (N_15365,N_14251,N_14619);
and U15366 (N_15366,N_14446,N_13732);
nor U15367 (N_15367,N_14618,N_14159);
nand U15368 (N_15368,N_13806,N_13605);
or U15369 (N_15369,N_14157,N_14941);
and U15370 (N_15370,N_14357,N_14140);
or U15371 (N_15371,N_14605,N_13867);
nor U15372 (N_15372,N_13728,N_13765);
nor U15373 (N_15373,N_13515,N_14025);
nor U15374 (N_15374,N_14731,N_13767);
or U15375 (N_15375,N_14760,N_14570);
or U15376 (N_15376,N_14971,N_14175);
or U15377 (N_15377,N_13733,N_14144);
nand U15378 (N_15378,N_14715,N_14527);
nor U15379 (N_15379,N_13944,N_14583);
nand U15380 (N_15380,N_13804,N_14560);
and U15381 (N_15381,N_14143,N_14290);
xnor U15382 (N_15382,N_13606,N_14069);
xnor U15383 (N_15383,N_13694,N_14413);
and U15384 (N_15384,N_14041,N_14636);
and U15385 (N_15385,N_14781,N_13755);
nand U15386 (N_15386,N_14820,N_14276);
nand U15387 (N_15387,N_13584,N_14346);
or U15388 (N_15388,N_13597,N_13609);
and U15389 (N_15389,N_14070,N_14131);
nand U15390 (N_15390,N_14052,N_14470);
or U15391 (N_15391,N_14547,N_14216);
or U15392 (N_15392,N_14429,N_14423);
nor U15393 (N_15393,N_14983,N_14362);
and U15394 (N_15394,N_13878,N_14627);
and U15395 (N_15395,N_14355,N_14719);
nand U15396 (N_15396,N_13999,N_14996);
or U15397 (N_15397,N_13740,N_14153);
and U15398 (N_15398,N_14391,N_13782);
xnor U15399 (N_15399,N_14394,N_13789);
and U15400 (N_15400,N_14481,N_14643);
nand U15401 (N_15401,N_14426,N_13824);
or U15402 (N_15402,N_14404,N_14693);
xnor U15403 (N_15403,N_14329,N_14472);
and U15404 (N_15404,N_13604,N_13669);
nand U15405 (N_15405,N_13854,N_14318);
or U15406 (N_15406,N_13718,N_13957);
nor U15407 (N_15407,N_13919,N_14558);
or U15408 (N_15408,N_14176,N_13808);
or U15409 (N_15409,N_14749,N_13853);
xor U15410 (N_15410,N_13538,N_14304);
or U15411 (N_15411,N_14812,N_14334);
nor U15412 (N_15412,N_14037,N_14325);
and U15413 (N_15413,N_13938,N_14292);
nor U15414 (N_15414,N_14587,N_14498);
and U15415 (N_15415,N_13762,N_14849);
nor U15416 (N_15416,N_14846,N_14633);
and U15417 (N_15417,N_14654,N_14141);
or U15418 (N_15418,N_14556,N_14229);
or U15419 (N_15419,N_13511,N_14406);
nand U15420 (N_15420,N_14973,N_13970);
and U15421 (N_15421,N_14837,N_14393);
and U15422 (N_15422,N_13524,N_13905);
xnor U15423 (N_15423,N_14943,N_14575);
or U15424 (N_15424,N_14420,N_14311);
nand U15425 (N_15425,N_14842,N_14647);
nand U15426 (N_15426,N_14179,N_14586);
nor U15427 (N_15427,N_14000,N_14638);
nor U15428 (N_15428,N_14607,N_14590);
xnor U15429 (N_15429,N_13773,N_14172);
nor U15430 (N_15430,N_13771,N_13883);
nor U15431 (N_15431,N_14419,N_14601);
nand U15432 (N_15432,N_14702,N_14817);
nor U15433 (N_15433,N_14997,N_14469);
xor U15434 (N_15434,N_14328,N_13979);
and U15435 (N_15435,N_14506,N_14737);
and U15436 (N_15436,N_14802,N_14592);
xnor U15437 (N_15437,N_14970,N_14704);
xor U15438 (N_15438,N_14758,N_13657);
nand U15439 (N_15439,N_14152,N_13880);
and U15440 (N_15440,N_14792,N_14267);
xnor U15441 (N_15441,N_14892,N_14746);
or U15442 (N_15442,N_14125,N_13567);
nand U15443 (N_15443,N_13914,N_14811);
xor U15444 (N_15444,N_14720,N_14214);
and U15445 (N_15445,N_14050,N_14053);
or U15446 (N_15446,N_13763,N_14891);
and U15447 (N_15447,N_14589,N_14927);
nor U15448 (N_15448,N_13758,N_14255);
xnor U15449 (N_15449,N_14797,N_14044);
or U15450 (N_15450,N_14114,N_14201);
or U15451 (N_15451,N_14816,N_13876);
nand U15452 (N_15452,N_14342,N_13749);
or U15453 (N_15453,N_13517,N_13996);
and U15454 (N_15454,N_14513,N_14606);
nor U15455 (N_15455,N_13611,N_14793);
xor U15456 (N_15456,N_13838,N_14250);
nor U15457 (N_15457,N_14208,N_14482);
and U15458 (N_15458,N_14440,N_14531);
and U15459 (N_15459,N_13818,N_14215);
xnor U15460 (N_15460,N_13889,N_14269);
or U15461 (N_15461,N_13858,N_14757);
or U15462 (N_15462,N_14765,N_14691);
or U15463 (N_15463,N_14002,N_14798);
and U15464 (N_15464,N_13548,N_14580);
nand U15465 (N_15465,N_14156,N_14194);
xnor U15466 (N_15466,N_13967,N_14352);
xnor U15467 (N_15467,N_13796,N_14933);
nor U15468 (N_15468,N_13549,N_13650);
and U15469 (N_15469,N_14919,N_14071);
nor U15470 (N_15470,N_13572,N_13552);
or U15471 (N_15471,N_14307,N_14437);
and U15472 (N_15472,N_14354,N_14616);
nor U15473 (N_15473,N_13885,N_13984);
or U15474 (N_15474,N_14968,N_13563);
nand U15475 (N_15475,N_13617,N_14193);
nand U15476 (N_15476,N_13696,N_13689);
xor U15477 (N_15477,N_14219,N_13766);
nand U15478 (N_15478,N_14100,N_14855);
and U15479 (N_15479,N_14403,N_14569);
nor U15480 (N_15480,N_13729,N_14137);
or U15481 (N_15481,N_13546,N_13874);
or U15482 (N_15482,N_13918,N_13863);
and U15483 (N_15483,N_14741,N_14902);
xor U15484 (N_15484,N_14931,N_14369);
xor U15485 (N_15485,N_14684,N_14514);
nor U15486 (N_15486,N_13935,N_13986);
nand U15487 (N_15487,N_14008,N_14687);
nand U15488 (N_15488,N_13662,N_14949);
or U15489 (N_15489,N_14763,N_14924);
and U15490 (N_15490,N_13652,N_13625);
or U15491 (N_15491,N_13705,N_13583);
or U15492 (N_15492,N_14177,N_13610);
nor U15493 (N_15493,N_13686,N_13783);
nand U15494 (N_15494,N_13551,N_14834);
or U15495 (N_15495,N_13607,N_13726);
nand U15496 (N_15496,N_14734,N_14414);
and U15497 (N_15497,N_13737,N_14847);
xor U15498 (N_15498,N_13594,N_14161);
and U15499 (N_15499,N_14323,N_14303);
nor U15500 (N_15500,N_13879,N_13541);
and U15501 (N_15501,N_13683,N_14243);
nand U15502 (N_15502,N_14645,N_13738);
and U15503 (N_15503,N_14382,N_13514);
xor U15504 (N_15504,N_13653,N_14376);
and U15505 (N_15505,N_14940,N_14240);
nand U15506 (N_15506,N_13671,N_13993);
xor U15507 (N_15507,N_14080,N_14231);
nand U15508 (N_15508,N_13940,N_14540);
and U15509 (N_15509,N_14885,N_14872);
xor U15510 (N_15510,N_13856,N_13844);
or U15511 (N_15511,N_14438,N_14124);
nand U15512 (N_15512,N_14246,N_14431);
nand U15513 (N_15513,N_14007,N_13901);
and U15514 (N_15514,N_14031,N_14539);
or U15515 (N_15515,N_14528,N_14922);
nor U15516 (N_15516,N_14109,N_14598);
and U15517 (N_15517,N_14245,N_14242);
and U15518 (N_15518,N_13526,N_14916);
or U15519 (N_15519,N_14956,N_13660);
nor U15520 (N_15520,N_13692,N_13839);
xnor U15521 (N_15521,N_13799,N_13564);
or U15522 (N_15522,N_14591,N_14543);
xor U15523 (N_15523,N_13553,N_14984);
or U15524 (N_15524,N_14182,N_14951);
nor U15525 (N_15525,N_14995,N_13708);
and U15526 (N_15526,N_13644,N_14204);
and U15527 (N_15527,N_13910,N_14518);
and U15528 (N_15528,N_14336,N_14574);
nand U15529 (N_15529,N_13852,N_14449);
nand U15530 (N_15530,N_14084,N_14345);
xnor U15531 (N_15531,N_14676,N_13619);
nor U15532 (N_15532,N_14967,N_13974);
nor U15533 (N_15533,N_14830,N_14603);
nand U15534 (N_15534,N_14698,N_14210);
xnor U15535 (N_15535,N_13759,N_14043);
xnor U15536 (N_15536,N_13666,N_13547);
and U15537 (N_15537,N_14538,N_14652);
xor U15538 (N_15538,N_14553,N_14629);
or U15539 (N_15539,N_14750,N_13975);
or U15540 (N_15540,N_13745,N_14599);
nand U15541 (N_15541,N_14930,N_14626);
and U15542 (N_15542,N_13768,N_14389);
xnor U15543 (N_15543,N_14298,N_14022);
xor U15544 (N_15544,N_13573,N_14882);
nor U15545 (N_15545,N_14621,N_14925);
nor U15546 (N_15546,N_13561,N_13674);
or U15547 (N_15547,N_14467,N_14767);
nand U15548 (N_15548,N_14273,N_14858);
nand U15549 (N_15549,N_13593,N_14524);
nor U15550 (N_15550,N_13608,N_14383);
and U15551 (N_15551,N_14692,N_14119);
xnor U15552 (N_15552,N_14078,N_14271);
nand U15553 (N_15553,N_14384,N_13641);
and U15554 (N_15554,N_13501,N_13932);
and U15555 (N_15555,N_14096,N_14850);
or U15556 (N_15556,N_13923,N_13739);
and U15557 (N_15557,N_14656,N_13555);
and U15558 (N_15558,N_14752,N_14138);
and U15559 (N_15559,N_13636,N_14610);
and U15560 (N_15560,N_14946,N_14443);
and U15561 (N_15561,N_14428,N_14794);
xnor U15562 (N_15562,N_14300,N_14632);
or U15563 (N_15563,N_14263,N_14012);
xnor U15564 (N_15564,N_14986,N_14163);
or U15565 (N_15565,N_14653,N_13620);
xnor U15566 (N_15566,N_14567,N_14988);
and U15567 (N_15567,N_14718,N_14450);
xnor U15568 (N_15568,N_14659,N_13881);
nand U15569 (N_15569,N_14529,N_14901);
xnor U15570 (N_15570,N_13976,N_13829);
or U15571 (N_15571,N_13648,N_14270);
nand U15572 (N_15572,N_13961,N_14055);
and U15573 (N_15573,N_14107,N_14260);
and U15574 (N_15574,N_13627,N_13850);
xor U15575 (N_15575,N_14212,N_14320);
and U15576 (N_15576,N_14101,N_13592);
xor U15577 (N_15577,N_13535,N_13815);
nand U15578 (N_15578,N_14511,N_13802);
xnor U15579 (N_15579,N_13836,N_14544);
nor U15580 (N_15580,N_14960,N_14649);
nor U15581 (N_15581,N_14628,N_14576);
nor U15582 (N_15582,N_13687,N_14021);
nand U15583 (N_15583,N_14678,N_14060);
and U15584 (N_15584,N_14953,N_13720);
or U15585 (N_15585,N_14917,N_13668);
or U15586 (N_15586,N_14377,N_14455);
nand U15587 (N_15587,N_13750,N_13531);
xor U15588 (N_15588,N_14064,N_13835);
and U15589 (N_15589,N_13639,N_14297);
nand U15590 (N_15590,N_14557,N_14324);
or U15591 (N_15591,N_13587,N_13942);
nand U15592 (N_15592,N_13513,N_14681);
nor U15593 (N_15593,N_14668,N_14067);
xor U15594 (N_15594,N_14799,N_14477);
or U15595 (N_15595,N_14667,N_14717);
or U15596 (N_15596,N_14671,N_14480);
xnor U15597 (N_15597,N_13742,N_14677);
and U15598 (N_15598,N_14396,N_14082);
nor U15599 (N_15599,N_14099,N_14221);
xor U15600 (N_15600,N_13510,N_13896);
nand U15601 (N_15601,N_13715,N_13581);
and U15602 (N_15602,N_14296,N_14723);
nor U15603 (N_15603,N_13897,N_14897);
nor U15604 (N_15604,N_13890,N_14266);
xor U15605 (N_15605,N_14876,N_13537);
and U15606 (N_15606,N_13529,N_13956);
xor U15607 (N_15607,N_14884,N_14865);
nor U15608 (N_15608,N_13917,N_14442);
nor U15609 (N_15609,N_13736,N_13903);
nor U15610 (N_15610,N_14854,N_13577);
and U15611 (N_15611,N_14889,N_14738);
and U15612 (N_15612,N_13803,N_13934);
and U15613 (N_15613,N_14740,N_13673);
and U15614 (N_15614,N_14453,N_14483);
nor U15615 (N_15615,N_14110,N_14965);
or U15616 (N_15616,N_14695,N_14206);
and U15617 (N_15617,N_14030,N_14743);
nand U15618 (N_15618,N_14128,N_13622);
or U15619 (N_15619,N_14015,N_13882);
nor U15620 (N_15620,N_13982,N_13945);
xnor U15621 (N_15621,N_13857,N_14283);
nand U15622 (N_15622,N_13862,N_13784);
nor U15623 (N_15623,N_13798,N_13939);
xor U15624 (N_15624,N_14989,N_14769);
nand U15625 (N_15625,N_13966,N_13795);
nor U15626 (N_15626,N_14288,N_13554);
nand U15627 (N_15627,N_14364,N_14223);
nor U15628 (N_15628,N_13562,N_14366);
nand U15629 (N_15629,N_14732,N_14003);
xor U15630 (N_15630,N_13911,N_14436);
xnor U15631 (N_15631,N_14559,N_13987);
nor U15632 (N_15632,N_14883,N_14700);
nor U15633 (N_15633,N_14017,N_14521);
xnor U15634 (N_15634,N_14401,N_14347);
xor U15635 (N_15635,N_13575,N_13964);
nor U15636 (N_15636,N_14814,N_13823);
nor U15637 (N_15637,N_14641,N_14402);
and U15638 (N_15638,N_14370,N_13507);
xor U15639 (N_15639,N_14412,N_13536);
and U15640 (N_15640,N_13931,N_13887);
nor U15641 (N_15641,N_14937,N_13643);
and U15642 (N_15642,N_14451,N_14225);
nand U15643 (N_15643,N_14501,N_14398);
nand U15644 (N_15644,N_14699,N_13628);
xnor U15645 (N_15645,N_14990,N_13527);
or U15646 (N_15646,N_14899,N_13559);
xor U15647 (N_15647,N_13520,N_14405);
nand U15648 (N_15648,N_14203,N_14686);
xnor U15649 (N_15649,N_13703,N_13775);
and U15650 (N_15650,N_14239,N_13722);
xor U15651 (N_15651,N_14220,N_14503);
xor U15652 (N_15652,N_13691,N_14407);
nor U15653 (N_15653,N_14285,N_14894);
xnor U15654 (N_15654,N_13596,N_13872);
nand U15655 (N_15655,N_14473,N_14707);
nand U15656 (N_15656,N_13528,N_14392);
and U15657 (N_15657,N_14839,N_13778);
nor U15658 (N_15658,N_14783,N_13990);
or U15659 (N_15659,N_14004,N_14709);
xor U15660 (N_15660,N_14294,N_14063);
and U15661 (N_15661,N_14549,N_14439);
or U15662 (N_15662,N_14934,N_14112);
or U15663 (N_15663,N_13591,N_14410);
nor U15664 (N_15664,N_14886,N_14999);
nor U15665 (N_15665,N_14308,N_14907);
nor U15666 (N_15666,N_14904,N_13813);
nand U15667 (N_15667,N_14818,N_13508);
nand U15668 (N_15668,N_14094,N_14434);
nand U15669 (N_15669,N_14258,N_14257);
or U15670 (N_15670,N_13684,N_14249);
and U15671 (N_15671,N_14278,N_14982);
nand U15672 (N_15672,N_14103,N_14655);
xnor U15673 (N_15673,N_13568,N_13834);
xor U15674 (N_15674,N_14185,N_14309);
and U15675 (N_15675,N_13602,N_13963);
nor U15676 (N_15676,N_13927,N_14571);
xnor U15677 (N_15677,N_13693,N_14588);
nand U15678 (N_15678,N_13670,N_13922);
nor U15679 (N_15679,N_13635,N_14095);
or U15680 (N_15680,N_14105,N_13590);
xor U15681 (N_15681,N_14174,N_14486);
and U15682 (N_15682,N_14073,N_14962);
nor U15683 (N_15683,N_13991,N_14562);
or U15684 (N_15684,N_14708,N_14444);
nor U15685 (N_15685,N_14327,N_14733);
nor U15686 (N_15686,N_14713,N_13831);
and U15687 (N_15687,N_14418,N_14227);
and U15688 (N_15688,N_13906,N_14178);
nand U15689 (N_15689,N_14739,N_13544);
nor U15690 (N_15690,N_14180,N_13675);
and U15691 (N_15691,N_14526,N_14018);
xor U15692 (N_15692,N_14367,N_14780);
nor U15693 (N_15693,N_13924,N_14779);
and U15694 (N_15694,N_14945,N_14905);
nand U15695 (N_15695,N_14319,N_14456);
and U15696 (N_15696,N_13532,N_13816);
xnor U15697 (N_15697,N_14268,N_14202);
xnor U15698 (N_15698,N_13805,N_14993);
and U15699 (N_15699,N_13864,N_13977);
and U15700 (N_15700,N_14650,N_14187);
and U15701 (N_15701,N_13710,N_14427);
and U15702 (N_15702,N_14938,N_14322);
or U15703 (N_15703,N_14295,N_14751);
and U15704 (N_15704,N_13794,N_14725);
nand U15705 (N_15705,N_14077,N_14149);
nand U15706 (N_15706,N_14136,N_14317);
xor U15707 (N_15707,N_14771,N_14235);
nand U15708 (N_15708,N_14046,N_13682);
xor U15709 (N_15709,N_13558,N_14921);
xor U15710 (N_15710,N_14058,N_13633);
and U15711 (N_15711,N_13747,N_13523);
and U15712 (N_15712,N_13569,N_14117);
and U15713 (N_15713,N_13995,N_13530);
nor U15714 (N_15714,N_14845,N_13833);
xnor U15715 (N_15715,N_14685,N_14234);
or U15716 (N_15716,N_14291,N_13790);
or U15717 (N_15717,N_14913,N_14604);
nand U15718 (N_15718,N_14813,N_13645);
nor U15719 (N_15719,N_13943,N_14759);
xor U15720 (N_15720,N_13997,N_14690);
or U15721 (N_15721,N_13809,N_14475);
xnor U15722 (N_15722,N_13843,N_14630);
and U15723 (N_15723,N_14039,N_14620);
nor U15724 (N_15724,N_14980,N_14611);
nand U15725 (N_15725,N_14939,N_13505);
nand U15726 (N_15726,N_13846,N_14530);
or U15727 (N_15727,N_14829,N_13734);
nor U15728 (N_15728,N_13928,N_14489);
xor U15729 (N_15729,N_14648,N_13830);
or U15730 (N_15730,N_14735,N_14097);
or U15731 (N_15731,N_14059,N_14005);
and U15732 (N_15732,N_14065,N_14035);
and U15733 (N_15733,N_14150,N_13909);
nor U15734 (N_15734,N_13820,N_14332);
or U15735 (N_15735,N_14274,N_13714);
nor U15736 (N_15736,N_14522,N_14662);
xnor U15737 (N_15737,N_13777,N_13930);
xor U15738 (N_15738,N_14350,N_13646);
xnor U15739 (N_15739,N_14359,N_14623);
nor U15740 (N_15740,N_14445,N_13791);
nor U15741 (N_15741,N_14914,N_14120);
or U15742 (N_15742,N_14582,N_13861);
nor U15743 (N_15743,N_13866,N_14762);
nand U15744 (N_15744,N_14388,N_14042);
or U15745 (N_15745,N_14581,N_13542);
nand U15746 (N_15746,N_14331,N_13751);
nand U15747 (N_15747,N_14027,N_14397);
or U15748 (N_15748,N_14313,N_13907);
or U15749 (N_15749,N_14795,N_13678);
nand U15750 (N_15750,N_14303,N_14718);
nor U15751 (N_15751,N_13990,N_13905);
nor U15752 (N_15752,N_13935,N_14525);
and U15753 (N_15753,N_14513,N_14770);
xnor U15754 (N_15754,N_13778,N_14192);
or U15755 (N_15755,N_13527,N_13532);
or U15756 (N_15756,N_14004,N_14210);
and U15757 (N_15757,N_14741,N_13579);
and U15758 (N_15758,N_14690,N_14318);
or U15759 (N_15759,N_14133,N_14042);
or U15760 (N_15760,N_14436,N_14350);
xnor U15761 (N_15761,N_14285,N_14100);
or U15762 (N_15762,N_14290,N_14986);
or U15763 (N_15763,N_14995,N_13826);
and U15764 (N_15764,N_13794,N_14452);
and U15765 (N_15765,N_14814,N_13549);
and U15766 (N_15766,N_13812,N_13640);
and U15767 (N_15767,N_13971,N_14091);
nand U15768 (N_15768,N_13975,N_14635);
xnor U15769 (N_15769,N_14920,N_14897);
nand U15770 (N_15770,N_14097,N_14754);
xor U15771 (N_15771,N_14223,N_13895);
and U15772 (N_15772,N_14620,N_14178);
or U15773 (N_15773,N_13773,N_14845);
and U15774 (N_15774,N_14279,N_13639);
nor U15775 (N_15775,N_14875,N_14969);
nor U15776 (N_15776,N_14455,N_14048);
or U15777 (N_15777,N_14171,N_14189);
nand U15778 (N_15778,N_14481,N_13563);
or U15779 (N_15779,N_14603,N_13889);
nand U15780 (N_15780,N_14601,N_14739);
xor U15781 (N_15781,N_13533,N_13628);
xor U15782 (N_15782,N_14012,N_14104);
or U15783 (N_15783,N_13690,N_13750);
nor U15784 (N_15784,N_13643,N_14100);
xor U15785 (N_15785,N_14446,N_14963);
nor U15786 (N_15786,N_13777,N_14779);
nand U15787 (N_15787,N_14771,N_14575);
nand U15788 (N_15788,N_13518,N_13854);
xor U15789 (N_15789,N_14539,N_14199);
nand U15790 (N_15790,N_13755,N_14289);
and U15791 (N_15791,N_14905,N_14627);
nand U15792 (N_15792,N_14159,N_14353);
nor U15793 (N_15793,N_14355,N_14512);
and U15794 (N_15794,N_14302,N_14621);
nor U15795 (N_15795,N_14508,N_14078);
or U15796 (N_15796,N_14970,N_14443);
nand U15797 (N_15797,N_14639,N_13709);
nand U15798 (N_15798,N_14708,N_13979);
nor U15799 (N_15799,N_14455,N_14117);
xor U15800 (N_15800,N_14233,N_14134);
nor U15801 (N_15801,N_13876,N_14849);
xnor U15802 (N_15802,N_14035,N_14269);
or U15803 (N_15803,N_14480,N_14395);
and U15804 (N_15804,N_13872,N_14846);
and U15805 (N_15805,N_13933,N_13503);
xor U15806 (N_15806,N_14575,N_14871);
nor U15807 (N_15807,N_14234,N_14239);
nand U15808 (N_15808,N_14415,N_14982);
or U15809 (N_15809,N_14641,N_13826);
xor U15810 (N_15810,N_13892,N_13840);
nand U15811 (N_15811,N_14119,N_13940);
or U15812 (N_15812,N_14275,N_13937);
and U15813 (N_15813,N_13991,N_13574);
xnor U15814 (N_15814,N_14164,N_14381);
xor U15815 (N_15815,N_14920,N_14071);
or U15816 (N_15816,N_13933,N_13685);
and U15817 (N_15817,N_14723,N_14313);
and U15818 (N_15818,N_14976,N_14101);
nand U15819 (N_15819,N_13792,N_14590);
nand U15820 (N_15820,N_13692,N_13945);
and U15821 (N_15821,N_13962,N_14175);
xor U15822 (N_15822,N_13537,N_14156);
and U15823 (N_15823,N_14887,N_13900);
nand U15824 (N_15824,N_14770,N_13657);
xor U15825 (N_15825,N_14657,N_14370);
nand U15826 (N_15826,N_14538,N_13529);
nor U15827 (N_15827,N_14411,N_13576);
or U15828 (N_15828,N_14872,N_14910);
nor U15829 (N_15829,N_14604,N_14537);
xnor U15830 (N_15830,N_13765,N_14789);
nand U15831 (N_15831,N_14306,N_14062);
or U15832 (N_15832,N_13896,N_14348);
xor U15833 (N_15833,N_14419,N_14815);
nor U15834 (N_15834,N_14100,N_13757);
or U15835 (N_15835,N_14348,N_14976);
nand U15836 (N_15836,N_14012,N_14264);
or U15837 (N_15837,N_14144,N_14243);
and U15838 (N_15838,N_14064,N_13907);
nand U15839 (N_15839,N_13938,N_13895);
nor U15840 (N_15840,N_13691,N_13837);
nor U15841 (N_15841,N_14384,N_13754);
nor U15842 (N_15842,N_13638,N_14812);
xnor U15843 (N_15843,N_14393,N_14952);
or U15844 (N_15844,N_14223,N_14972);
nor U15845 (N_15845,N_13960,N_14557);
and U15846 (N_15846,N_13868,N_14105);
xnor U15847 (N_15847,N_13801,N_13562);
nand U15848 (N_15848,N_13716,N_13925);
xor U15849 (N_15849,N_13789,N_14822);
xnor U15850 (N_15850,N_14390,N_14337);
or U15851 (N_15851,N_13809,N_14901);
or U15852 (N_15852,N_14872,N_13979);
nand U15853 (N_15853,N_14531,N_13603);
xor U15854 (N_15854,N_14737,N_14015);
nand U15855 (N_15855,N_14192,N_14136);
xnor U15856 (N_15856,N_13817,N_14846);
nor U15857 (N_15857,N_14026,N_14564);
nand U15858 (N_15858,N_14147,N_14037);
nand U15859 (N_15859,N_14143,N_14693);
or U15860 (N_15860,N_14647,N_13978);
nor U15861 (N_15861,N_13968,N_13681);
and U15862 (N_15862,N_14504,N_14546);
and U15863 (N_15863,N_13761,N_14880);
xnor U15864 (N_15864,N_14275,N_13714);
and U15865 (N_15865,N_14342,N_13772);
nand U15866 (N_15866,N_14863,N_14890);
or U15867 (N_15867,N_14205,N_13664);
or U15868 (N_15868,N_14934,N_13589);
xnor U15869 (N_15869,N_14718,N_14858);
or U15870 (N_15870,N_13636,N_14611);
or U15871 (N_15871,N_13579,N_14611);
xnor U15872 (N_15872,N_14834,N_14159);
nor U15873 (N_15873,N_14018,N_13948);
nor U15874 (N_15874,N_13891,N_13882);
nand U15875 (N_15875,N_14587,N_14010);
nand U15876 (N_15876,N_14632,N_14523);
and U15877 (N_15877,N_13930,N_14411);
nand U15878 (N_15878,N_14537,N_14017);
xnor U15879 (N_15879,N_14027,N_14959);
or U15880 (N_15880,N_14755,N_13814);
xnor U15881 (N_15881,N_13845,N_14940);
nor U15882 (N_15882,N_14272,N_14189);
or U15883 (N_15883,N_13667,N_13565);
and U15884 (N_15884,N_14364,N_14800);
xor U15885 (N_15885,N_14130,N_14527);
or U15886 (N_15886,N_13701,N_13801);
or U15887 (N_15887,N_14818,N_14616);
nand U15888 (N_15888,N_13992,N_14897);
nor U15889 (N_15889,N_14315,N_14834);
xor U15890 (N_15890,N_14231,N_14677);
or U15891 (N_15891,N_14104,N_14293);
nand U15892 (N_15892,N_13917,N_14032);
xnor U15893 (N_15893,N_13564,N_14661);
and U15894 (N_15894,N_14545,N_13640);
and U15895 (N_15895,N_14890,N_13953);
nor U15896 (N_15896,N_14483,N_14738);
and U15897 (N_15897,N_14642,N_14797);
xor U15898 (N_15898,N_13963,N_14372);
nand U15899 (N_15899,N_14532,N_13500);
xnor U15900 (N_15900,N_13988,N_14565);
or U15901 (N_15901,N_14026,N_14395);
nand U15902 (N_15902,N_13901,N_14966);
or U15903 (N_15903,N_14549,N_13920);
or U15904 (N_15904,N_14525,N_13950);
nand U15905 (N_15905,N_13766,N_14674);
nor U15906 (N_15906,N_14066,N_13953);
or U15907 (N_15907,N_13545,N_14867);
or U15908 (N_15908,N_14169,N_14929);
or U15909 (N_15909,N_14783,N_14085);
nor U15910 (N_15910,N_13870,N_14404);
nor U15911 (N_15911,N_14118,N_14443);
and U15912 (N_15912,N_14554,N_14270);
or U15913 (N_15913,N_14992,N_14425);
and U15914 (N_15914,N_13551,N_13816);
xor U15915 (N_15915,N_13608,N_14523);
nor U15916 (N_15916,N_14332,N_14293);
or U15917 (N_15917,N_13722,N_13503);
and U15918 (N_15918,N_13775,N_14767);
nor U15919 (N_15919,N_13633,N_14189);
nand U15920 (N_15920,N_14103,N_14250);
nand U15921 (N_15921,N_14919,N_14231);
or U15922 (N_15922,N_13964,N_14991);
or U15923 (N_15923,N_14158,N_13558);
or U15924 (N_15924,N_13558,N_14261);
nor U15925 (N_15925,N_14016,N_14695);
and U15926 (N_15926,N_13972,N_13541);
nor U15927 (N_15927,N_14597,N_14423);
nor U15928 (N_15928,N_14259,N_14432);
and U15929 (N_15929,N_14722,N_14296);
nor U15930 (N_15930,N_14661,N_14736);
nor U15931 (N_15931,N_14814,N_14633);
and U15932 (N_15932,N_13862,N_14734);
nand U15933 (N_15933,N_14929,N_14171);
and U15934 (N_15934,N_13639,N_14342);
nor U15935 (N_15935,N_14930,N_13916);
xnor U15936 (N_15936,N_14725,N_14023);
nand U15937 (N_15937,N_14268,N_13658);
xor U15938 (N_15938,N_14543,N_14204);
and U15939 (N_15939,N_13848,N_14959);
or U15940 (N_15940,N_14067,N_13937);
and U15941 (N_15941,N_13743,N_14453);
xnor U15942 (N_15942,N_14595,N_13869);
or U15943 (N_15943,N_14791,N_14071);
or U15944 (N_15944,N_13995,N_14845);
or U15945 (N_15945,N_13670,N_13705);
nor U15946 (N_15946,N_14017,N_14306);
and U15947 (N_15947,N_14924,N_14137);
or U15948 (N_15948,N_14902,N_13678);
nand U15949 (N_15949,N_14391,N_13529);
or U15950 (N_15950,N_14113,N_14926);
or U15951 (N_15951,N_14557,N_14136);
xor U15952 (N_15952,N_13828,N_13728);
nor U15953 (N_15953,N_14608,N_14009);
nor U15954 (N_15954,N_13650,N_13935);
nand U15955 (N_15955,N_14782,N_14507);
and U15956 (N_15956,N_14627,N_14492);
or U15957 (N_15957,N_13831,N_14404);
nor U15958 (N_15958,N_13602,N_14620);
nor U15959 (N_15959,N_14782,N_14629);
and U15960 (N_15960,N_13568,N_13935);
nand U15961 (N_15961,N_14865,N_14328);
xor U15962 (N_15962,N_13707,N_14229);
nor U15963 (N_15963,N_14764,N_13926);
nand U15964 (N_15964,N_14823,N_13572);
xor U15965 (N_15965,N_14366,N_14973);
nand U15966 (N_15966,N_14604,N_13778);
and U15967 (N_15967,N_13996,N_14131);
nand U15968 (N_15968,N_13501,N_13980);
and U15969 (N_15969,N_13728,N_14235);
xor U15970 (N_15970,N_14197,N_14500);
nor U15971 (N_15971,N_14121,N_14443);
and U15972 (N_15972,N_14457,N_13655);
xnor U15973 (N_15973,N_14848,N_14573);
and U15974 (N_15974,N_14260,N_14667);
or U15975 (N_15975,N_14393,N_13801);
and U15976 (N_15976,N_14800,N_14675);
and U15977 (N_15977,N_14751,N_13962);
nand U15978 (N_15978,N_13809,N_13610);
and U15979 (N_15979,N_14561,N_14670);
and U15980 (N_15980,N_14315,N_14020);
nand U15981 (N_15981,N_13632,N_13823);
or U15982 (N_15982,N_14991,N_14142);
nand U15983 (N_15983,N_14788,N_14858);
and U15984 (N_15984,N_13838,N_14431);
nand U15985 (N_15985,N_14863,N_14944);
or U15986 (N_15986,N_14352,N_13651);
xnor U15987 (N_15987,N_14486,N_14552);
xnor U15988 (N_15988,N_14384,N_14627);
nor U15989 (N_15989,N_14545,N_13531);
nand U15990 (N_15990,N_14118,N_13787);
or U15991 (N_15991,N_14493,N_13680);
nor U15992 (N_15992,N_14641,N_14807);
nand U15993 (N_15993,N_14115,N_14821);
xor U15994 (N_15994,N_14625,N_14267);
nand U15995 (N_15995,N_14970,N_14777);
or U15996 (N_15996,N_14264,N_13738);
or U15997 (N_15997,N_14795,N_14176);
or U15998 (N_15998,N_13951,N_14863);
or U15999 (N_15999,N_13945,N_13845);
and U16000 (N_16000,N_14014,N_13794);
or U16001 (N_16001,N_14192,N_13799);
nand U16002 (N_16002,N_14838,N_14195);
nor U16003 (N_16003,N_14480,N_14413);
nor U16004 (N_16004,N_13924,N_14132);
or U16005 (N_16005,N_13558,N_13853);
nand U16006 (N_16006,N_13742,N_14141);
nor U16007 (N_16007,N_13613,N_13802);
nand U16008 (N_16008,N_14766,N_14634);
and U16009 (N_16009,N_14085,N_14774);
or U16010 (N_16010,N_14057,N_14916);
xor U16011 (N_16011,N_14475,N_13513);
nand U16012 (N_16012,N_14653,N_14681);
xnor U16013 (N_16013,N_14877,N_13515);
or U16014 (N_16014,N_14909,N_14775);
xor U16015 (N_16015,N_14836,N_14530);
nor U16016 (N_16016,N_14110,N_14489);
nand U16017 (N_16017,N_14400,N_14113);
and U16018 (N_16018,N_14059,N_14390);
or U16019 (N_16019,N_14822,N_13612);
or U16020 (N_16020,N_13735,N_13793);
or U16021 (N_16021,N_13641,N_13940);
xnor U16022 (N_16022,N_13646,N_14519);
and U16023 (N_16023,N_14017,N_14459);
nor U16024 (N_16024,N_14299,N_13769);
or U16025 (N_16025,N_14631,N_14374);
xor U16026 (N_16026,N_14311,N_13556);
xnor U16027 (N_16027,N_14682,N_14505);
nand U16028 (N_16028,N_13834,N_14593);
nor U16029 (N_16029,N_13734,N_14389);
xor U16030 (N_16030,N_14813,N_14111);
xnor U16031 (N_16031,N_14744,N_14145);
nor U16032 (N_16032,N_14544,N_13890);
or U16033 (N_16033,N_14271,N_14653);
and U16034 (N_16034,N_13536,N_14808);
nor U16035 (N_16035,N_14929,N_14506);
or U16036 (N_16036,N_14399,N_14237);
nand U16037 (N_16037,N_14871,N_14563);
nand U16038 (N_16038,N_14333,N_13786);
nor U16039 (N_16039,N_14663,N_14568);
nand U16040 (N_16040,N_14291,N_14958);
and U16041 (N_16041,N_14966,N_13977);
or U16042 (N_16042,N_14026,N_13781);
nand U16043 (N_16043,N_13779,N_13573);
xor U16044 (N_16044,N_13891,N_13525);
or U16045 (N_16045,N_14477,N_14421);
or U16046 (N_16046,N_13536,N_14182);
nor U16047 (N_16047,N_14211,N_14463);
or U16048 (N_16048,N_13913,N_13979);
nand U16049 (N_16049,N_13761,N_14284);
nor U16050 (N_16050,N_14571,N_14422);
nand U16051 (N_16051,N_14370,N_14110);
nor U16052 (N_16052,N_14707,N_14664);
and U16053 (N_16053,N_14101,N_13686);
and U16054 (N_16054,N_14012,N_14642);
or U16055 (N_16055,N_13888,N_14699);
or U16056 (N_16056,N_14920,N_14375);
and U16057 (N_16057,N_14151,N_14256);
and U16058 (N_16058,N_14401,N_14073);
xor U16059 (N_16059,N_14522,N_14137);
nand U16060 (N_16060,N_14799,N_14350);
xor U16061 (N_16061,N_14354,N_14701);
nand U16062 (N_16062,N_13969,N_13771);
or U16063 (N_16063,N_14662,N_14684);
and U16064 (N_16064,N_14272,N_14005);
and U16065 (N_16065,N_14671,N_14330);
nand U16066 (N_16066,N_14202,N_14734);
nor U16067 (N_16067,N_14177,N_14910);
nand U16068 (N_16068,N_13837,N_13764);
nand U16069 (N_16069,N_14690,N_14511);
or U16070 (N_16070,N_14662,N_14467);
or U16071 (N_16071,N_14318,N_14963);
nand U16072 (N_16072,N_13678,N_14609);
and U16073 (N_16073,N_14777,N_14689);
nand U16074 (N_16074,N_14947,N_14509);
nor U16075 (N_16075,N_14267,N_14863);
or U16076 (N_16076,N_14603,N_14762);
nor U16077 (N_16077,N_14747,N_14215);
and U16078 (N_16078,N_13864,N_13733);
or U16079 (N_16079,N_14634,N_13626);
and U16080 (N_16080,N_14724,N_14856);
or U16081 (N_16081,N_14384,N_13857);
nor U16082 (N_16082,N_14712,N_14018);
and U16083 (N_16083,N_14788,N_14759);
and U16084 (N_16084,N_13750,N_14137);
xnor U16085 (N_16085,N_14874,N_13846);
nor U16086 (N_16086,N_14367,N_14044);
and U16087 (N_16087,N_14579,N_14951);
and U16088 (N_16088,N_13574,N_13620);
nand U16089 (N_16089,N_14887,N_14387);
xor U16090 (N_16090,N_14398,N_14657);
nor U16091 (N_16091,N_14259,N_13583);
and U16092 (N_16092,N_14663,N_13871);
or U16093 (N_16093,N_14685,N_13644);
and U16094 (N_16094,N_14065,N_14342);
xor U16095 (N_16095,N_14362,N_14299);
and U16096 (N_16096,N_14494,N_14583);
or U16097 (N_16097,N_14009,N_14519);
nor U16098 (N_16098,N_13744,N_14017);
nand U16099 (N_16099,N_14285,N_14990);
or U16100 (N_16100,N_13882,N_14478);
or U16101 (N_16101,N_13842,N_14810);
nand U16102 (N_16102,N_14612,N_13653);
nand U16103 (N_16103,N_14813,N_14233);
and U16104 (N_16104,N_14340,N_14357);
nand U16105 (N_16105,N_14849,N_14873);
or U16106 (N_16106,N_14854,N_14173);
xnor U16107 (N_16107,N_14122,N_14059);
nand U16108 (N_16108,N_14177,N_14861);
nor U16109 (N_16109,N_14399,N_14508);
xnor U16110 (N_16110,N_13653,N_13913);
nand U16111 (N_16111,N_13511,N_13734);
nand U16112 (N_16112,N_14758,N_14426);
nand U16113 (N_16113,N_13864,N_14442);
or U16114 (N_16114,N_13728,N_13540);
or U16115 (N_16115,N_14286,N_14904);
nand U16116 (N_16116,N_13513,N_13996);
nor U16117 (N_16117,N_14456,N_13811);
nor U16118 (N_16118,N_13544,N_14857);
and U16119 (N_16119,N_14109,N_14226);
nor U16120 (N_16120,N_14270,N_13792);
nor U16121 (N_16121,N_14388,N_14340);
nor U16122 (N_16122,N_14460,N_13705);
nand U16123 (N_16123,N_13843,N_13546);
and U16124 (N_16124,N_14798,N_14186);
nand U16125 (N_16125,N_14464,N_14100);
and U16126 (N_16126,N_14008,N_14239);
nor U16127 (N_16127,N_14500,N_14854);
and U16128 (N_16128,N_14585,N_14128);
and U16129 (N_16129,N_14396,N_14669);
or U16130 (N_16130,N_14966,N_14495);
nor U16131 (N_16131,N_14765,N_14696);
and U16132 (N_16132,N_13547,N_14782);
nor U16133 (N_16133,N_14070,N_14387);
and U16134 (N_16134,N_14773,N_14438);
or U16135 (N_16135,N_13840,N_14367);
nor U16136 (N_16136,N_14783,N_13608);
and U16137 (N_16137,N_14129,N_14404);
nor U16138 (N_16138,N_14786,N_14763);
or U16139 (N_16139,N_14933,N_13691);
nand U16140 (N_16140,N_14555,N_14495);
and U16141 (N_16141,N_13862,N_13683);
or U16142 (N_16142,N_14878,N_13953);
nand U16143 (N_16143,N_14939,N_13966);
xnor U16144 (N_16144,N_13554,N_14901);
nor U16145 (N_16145,N_13728,N_14885);
nor U16146 (N_16146,N_14909,N_14580);
xnor U16147 (N_16147,N_14380,N_13669);
or U16148 (N_16148,N_14960,N_13942);
nor U16149 (N_16149,N_14926,N_14311);
or U16150 (N_16150,N_13862,N_13743);
and U16151 (N_16151,N_13649,N_13701);
and U16152 (N_16152,N_13856,N_13768);
nor U16153 (N_16153,N_14587,N_13735);
nand U16154 (N_16154,N_14251,N_14787);
nand U16155 (N_16155,N_14153,N_14897);
nor U16156 (N_16156,N_13513,N_13854);
and U16157 (N_16157,N_13604,N_13992);
nor U16158 (N_16158,N_13831,N_14816);
or U16159 (N_16159,N_13817,N_14514);
nor U16160 (N_16160,N_13765,N_14292);
nand U16161 (N_16161,N_14780,N_14236);
or U16162 (N_16162,N_14693,N_14876);
or U16163 (N_16163,N_14353,N_13509);
xor U16164 (N_16164,N_14202,N_13518);
nor U16165 (N_16165,N_13986,N_14237);
nand U16166 (N_16166,N_14105,N_13859);
xnor U16167 (N_16167,N_14538,N_14417);
and U16168 (N_16168,N_13880,N_13887);
nor U16169 (N_16169,N_14319,N_14228);
xor U16170 (N_16170,N_13580,N_14798);
xor U16171 (N_16171,N_14106,N_14492);
or U16172 (N_16172,N_14184,N_13985);
xnor U16173 (N_16173,N_14697,N_14540);
xor U16174 (N_16174,N_14604,N_14808);
xnor U16175 (N_16175,N_13693,N_14088);
xnor U16176 (N_16176,N_14596,N_13638);
nand U16177 (N_16177,N_14605,N_14585);
and U16178 (N_16178,N_13535,N_13507);
or U16179 (N_16179,N_13828,N_14803);
or U16180 (N_16180,N_14192,N_13605);
nor U16181 (N_16181,N_14970,N_13909);
nor U16182 (N_16182,N_14150,N_14032);
and U16183 (N_16183,N_13922,N_14507);
nor U16184 (N_16184,N_14247,N_13847);
or U16185 (N_16185,N_14754,N_14048);
or U16186 (N_16186,N_14447,N_14952);
or U16187 (N_16187,N_14681,N_13721);
or U16188 (N_16188,N_14262,N_14169);
nand U16189 (N_16189,N_14909,N_14991);
xor U16190 (N_16190,N_14245,N_13947);
nor U16191 (N_16191,N_13844,N_13715);
nor U16192 (N_16192,N_13937,N_14889);
nor U16193 (N_16193,N_14743,N_13643);
xnor U16194 (N_16194,N_14061,N_14946);
or U16195 (N_16195,N_14476,N_14106);
nor U16196 (N_16196,N_14397,N_13792);
and U16197 (N_16197,N_14098,N_14120);
xor U16198 (N_16198,N_14745,N_13591);
and U16199 (N_16199,N_14776,N_14230);
nand U16200 (N_16200,N_14658,N_14871);
nand U16201 (N_16201,N_14847,N_14759);
xnor U16202 (N_16202,N_14184,N_13722);
xnor U16203 (N_16203,N_13688,N_14813);
or U16204 (N_16204,N_13770,N_14337);
nor U16205 (N_16205,N_13692,N_13702);
nand U16206 (N_16206,N_13670,N_14326);
nand U16207 (N_16207,N_13734,N_13665);
and U16208 (N_16208,N_14929,N_13510);
xor U16209 (N_16209,N_14493,N_14585);
or U16210 (N_16210,N_13543,N_13926);
nor U16211 (N_16211,N_14887,N_14556);
and U16212 (N_16212,N_13623,N_14558);
nor U16213 (N_16213,N_14700,N_14829);
and U16214 (N_16214,N_14259,N_14411);
and U16215 (N_16215,N_14054,N_13662);
xnor U16216 (N_16216,N_14498,N_13774);
nor U16217 (N_16217,N_13915,N_13727);
nand U16218 (N_16218,N_14158,N_14571);
nor U16219 (N_16219,N_14840,N_14497);
and U16220 (N_16220,N_14117,N_14036);
or U16221 (N_16221,N_14319,N_13676);
nand U16222 (N_16222,N_14562,N_13665);
xor U16223 (N_16223,N_14024,N_14469);
nand U16224 (N_16224,N_14470,N_14371);
and U16225 (N_16225,N_14523,N_14154);
nor U16226 (N_16226,N_14390,N_13590);
nor U16227 (N_16227,N_13919,N_13695);
nand U16228 (N_16228,N_14074,N_14761);
nand U16229 (N_16229,N_14627,N_14548);
nand U16230 (N_16230,N_13589,N_14766);
xnor U16231 (N_16231,N_13705,N_13808);
nor U16232 (N_16232,N_14248,N_14365);
nor U16233 (N_16233,N_14126,N_14099);
xnor U16234 (N_16234,N_14108,N_13594);
xnor U16235 (N_16235,N_13775,N_13818);
or U16236 (N_16236,N_14718,N_13688);
and U16237 (N_16237,N_13505,N_13759);
nand U16238 (N_16238,N_14333,N_14134);
xor U16239 (N_16239,N_14555,N_14171);
or U16240 (N_16240,N_13908,N_14296);
xor U16241 (N_16241,N_14592,N_13722);
nor U16242 (N_16242,N_14195,N_14168);
xnor U16243 (N_16243,N_14493,N_13695);
nand U16244 (N_16244,N_14887,N_13704);
nand U16245 (N_16245,N_13842,N_13727);
xor U16246 (N_16246,N_13814,N_14716);
nand U16247 (N_16247,N_13804,N_13762);
and U16248 (N_16248,N_14667,N_13790);
and U16249 (N_16249,N_14942,N_13713);
or U16250 (N_16250,N_14131,N_13555);
nor U16251 (N_16251,N_13846,N_14025);
nand U16252 (N_16252,N_14064,N_13714);
or U16253 (N_16253,N_13885,N_14691);
or U16254 (N_16254,N_14946,N_14623);
nor U16255 (N_16255,N_14379,N_14197);
nor U16256 (N_16256,N_14559,N_14869);
xnor U16257 (N_16257,N_13811,N_13803);
or U16258 (N_16258,N_14096,N_14126);
or U16259 (N_16259,N_13818,N_14170);
xnor U16260 (N_16260,N_14495,N_13775);
nand U16261 (N_16261,N_13595,N_13963);
and U16262 (N_16262,N_14753,N_14081);
or U16263 (N_16263,N_14412,N_13977);
nor U16264 (N_16264,N_14161,N_14753);
xnor U16265 (N_16265,N_13694,N_14349);
xnor U16266 (N_16266,N_14896,N_13646);
and U16267 (N_16267,N_13888,N_13880);
xor U16268 (N_16268,N_14461,N_14786);
nand U16269 (N_16269,N_14473,N_14353);
xnor U16270 (N_16270,N_14901,N_14729);
xnor U16271 (N_16271,N_13917,N_14469);
nor U16272 (N_16272,N_14906,N_14190);
nor U16273 (N_16273,N_14571,N_14640);
nor U16274 (N_16274,N_14327,N_14063);
nor U16275 (N_16275,N_14426,N_14350);
nor U16276 (N_16276,N_14384,N_14789);
nand U16277 (N_16277,N_13523,N_14164);
or U16278 (N_16278,N_14403,N_13623);
nand U16279 (N_16279,N_14581,N_13966);
nor U16280 (N_16280,N_13989,N_13878);
xnor U16281 (N_16281,N_13826,N_14302);
nand U16282 (N_16282,N_13851,N_13632);
or U16283 (N_16283,N_13592,N_14353);
and U16284 (N_16284,N_14318,N_14047);
xnor U16285 (N_16285,N_13692,N_13674);
xnor U16286 (N_16286,N_14219,N_14169);
and U16287 (N_16287,N_14641,N_14497);
and U16288 (N_16288,N_14219,N_14605);
xor U16289 (N_16289,N_14058,N_14862);
or U16290 (N_16290,N_14736,N_13728);
nor U16291 (N_16291,N_14678,N_14758);
nor U16292 (N_16292,N_14360,N_13584);
or U16293 (N_16293,N_14272,N_14749);
and U16294 (N_16294,N_14583,N_14434);
or U16295 (N_16295,N_14701,N_14199);
xnor U16296 (N_16296,N_13577,N_13507);
or U16297 (N_16297,N_13847,N_13571);
and U16298 (N_16298,N_13942,N_14250);
nand U16299 (N_16299,N_14265,N_13506);
nor U16300 (N_16300,N_13940,N_14503);
and U16301 (N_16301,N_14457,N_14145);
and U16302 (N_16302,N_13765,N_13610);
nand U16303 (N_16303,N_14927,N_13775);
and U16304 (N_16304,N_14524,N_13534);
and U16305 (N_16305,N_13541,N_14661);
nor U16306 (N_16306,N_14799,N_13736);
or U16307 (N_16307,N_14986,N_13996);
and U16308 (N_16308,N_14422,N_13994);
xor U16309 (N_16309,N_13948,N_13506);
xnor U16310 (N_16310,N_13840,N_14187);
and U16311 (N_16311,N_14544,N_14600);
nand U16312 (N_16312,N_14367,N_14739);
nand U16313 (N_16313,N_13639,N_13692);
and U16314 (N_16314,N_14180,N_14032);
nand U16315 (N_16315,N_14885,N_14928);
nor U16316 (N_16316,N_14688,N_14944);
nand U16317 (N_16317,N_14776,N_14063);
or U16318 (N_16318,N_14080,N_13859);
and U16319 (N_16319,N_14879,N_13814);
and U16320 (N_16320,N_14150,N_13559);
xnor U16321 (N_16321,N_14315,N_13702);
and U16322 (N_16322,N_14527,N_14432);
nor U16323 (N_16323,N_14727,N_13876);
and U16324 (N_16324,N_14203,N_13940);
xor U16325 (N_16325,N_14371,N_14513);
xor U16326 (N_16326,N_13558,N_14105);
nand U16327 (N_16327,N_14544,N_14248);
xnor U16328 (N_16328,N_14521,N_14127);
and U16329 (N_16329,N_13777,N_14488);
xor U16330 (N_16330,N_14511,N_13672);
nand U16331 (N_16331,N_14657,N_14283);
or U16332 (N_16332,N_14312,N_13669);
or U16333 (N_16333,N_14666,N_13784);
nand U16334 (N_16334,N_13940,N_13965);
or U16335 (N_16335,N_13517,N_14598);
nand U16336 (N_16336,N_14460,N_14954);
and U16337 (N_16337,N_14387,N_14718);
nor U16338 (N_16338,N_13524,N_13656);
nor U16339 (N_16339,N_14996,N_14223);
nor U16340 (N_16340,N_13788,N_14404);
nor U16341 (N_16341,N_14978,N_14033);
nor U16342 (N_16342,N_14501,N_14900);
xor U16343 (N_16343,N_13809,N_14839);
or U16344 (N_16344,N_14552,N_14525);
nor U16345 (N_16345,N_14146,N_14036);
nand U16346 (N_16346,N_14152,N_14637);
xnor U16347 (N_16347,N_14224,N_14822);
xnor U16348 (N_16348,N_13775,N_13508);
or U16349 (N_16349,N_14137,N_13564);
nand U16350 (N_16350,N_14756,N_14742);
and U16351 (N_16351,N_13589,N_13670);
nand U16352 (N_16352,N_14389,N_14693);
nand U16353 (N_16353,N_13758,N_14418);
and U16354 (N_16354,N_14692,N_14937);
nor U16355 (N_16355,N_13691,N_14123);
or U16356 (N_16356,N_14422,N_13658);
nor U16357 (N_16357,N_13761,N_14032);
or U16358 (N_16358,N_14358,N_13665);
and U16359 (N_16359,N_14084,N_14719);
xnor U16360 (N_16360,N_13897,N_14830);
or U16361 (N_16361,N_14453,N_13675);
and U16362 (N_16362,N_14555,N_13956);
and U16363 (N_16363,N_14703,N_13515);
nand U16364 (N_16364,N_14221,N_13984);
nor U16365 (N_16365,N_14780,N_14304);
and U16366 (N_16366,N_14270,N_14500);
nor U16367 (N_16367,N_14486,N_14102);
or U16368 (N_16368,N_14887,N_14365);
xor U16369 (N_16369,N_13835,N_14720);
nor U16370 (N_16370,N_14574,N_13780);
nor U16371 (N_16371,N_14130,N_14399);
or U16372 (N_16372,N_14504,N_14916);
nand U16373 (N_16373,N_13884,N_13933);
and U16374 (N_16374,N_14354,N_14498);
nand U16375 (N_16375,N_13856,N_14212);
xor U16376 (N_16376,N_13584,N_13782);
nor U16377 (N_16377,N_13864,N_14798);
and U16378 (N_16378,N_14787,N_14941);
nand U16379 (N_16379,N_14728,N_14104);
nor U16380 (N_16380,N_14541,N_13607);
nor U16381 (N_16381,N_14405,N_14480);
or U16382 (N_16382,N_14877,N_13686);
and U16383 (N_16383,N_14989,N_13723);
nor U16384 (N_16384,N_14016,N_14138);
or U16385 (N_16385,N_13878,N_14187);
or U16386 (N_16386,N_14062,N_14025);
xor U16387 (N_16387,N_14857,N_14359);
xnor U16388 (N_16388,N_14772,N_14288);
xnor U16389 (N_16389,N_14687,N_13529);
and U16390 (N_16390,N_13860,N_13621);
and U16391 (N_16391,N_14159,N_14390);
or U16392 (N_16392,N_14805,N_13612);
xnor U16393 (N_16393,N_14934,N_14288);
nor U16394 (N_16394,N_13523,N_14492);
and U16395 (N_16395,N_13559,N_13663);
or U16396 (N_16396,N_14564,N_14333);
nand U16397 (N_16397,N_13648,N_14306);
or U16398 (N_16398,N_13656,N_14643);
nor U16399 (N_16399,N_14252,N_13764);
nand U16400 (N_16400,N_14143,N_14957);
nor U16401 (N_16401,N_14120,N_14050);
nand U16402 (N_16402,N_13686,N_14858);
xor U16403 (N_16403,N_13664,N_14965);
nor U16404 (N_16404,N_14442,N_14312);
and U16405 (N_16405,N_14421,N_13935);
nor U16406 (N_16406,N_14322,N_14857);
nand U16407 (N_16407,N_13615,N_14806);
xnor U16408 (N_16408,N_14457,N_13754);
nor U16409 (N_16409,N_14175,N_14758);
nand U16410 (N_16410,N_14553,N_14514);
and U16411 (N_16411,N_13850,N_14953);
nand U16412 (N_16412,N_14011,N_14385);
and U16413 (N_16413,N_14728,N_13632);
xor U16414 (N_16414,N_13848,N_13509);
nand U16415 (N_16415,N_14052,N_14313);
and U16416 (N_16416,N_14526,N_13971);
or U16417 (N_16417,N_14457,N_13594);
xnor U16418 (N_16418,N_13841,N_14860);
xor U16419 (N_16419,N_13631,N_14914);
nor U16420 (N_16420,N_13854,N_14321);
and U16421 (N_16421,N_13962,N_14426);
xor U16422 (N_16422,N_14376,N_14991);
and U16423 (N_16423,N_14375,N_14228);
and U16424 (N_16424,N_14813,N_14247);
and U16425 (N_16425,N_13992,N_14187);
and U16426 (N_16426,N_13612,N_13674);
nor U16427 (N_16427,N_14473,N_13762);
nand U16428 (N_16428,N_14171,N_14342);
nor U16429 (N_16429,N_14331,N_13636);
and U16430 (N_16430,N_13616,N_14224);
nand U16431 (N_16431,N_13821,N_14559);
xor U16432 (N_16432,N_14638,N_14338);
nor U16433 (N_16433,N_14082,N_14677);
and U16434 (N_16434,N_14422,N_14669);
nand U16435 (N_16435,N_14604,N_13751);
and U16436 (N_16436,N_13988,N_13883);
and U16437 (N_16437,N_14132,N_14350);
nand U16438 (N_16438,N_14582,N_13809);
nor U16439 (N_16439,N_14864,N_13695);
or U16440 (N_16440,N_14013,N_13696);
xnor U16441 (N_16441,N_13562,N_14918);
and U16442 (N_16442,N_14130,N_14680);
nor U16443 (N_16443,N_14189,N_13707);
nand U16444 (N_16444,N_14422,N_13861);
or U16445 (N_16445,N_14564,N_13849);
nor U16446 (N_16446,N_14826,N_13914);
and U16447 (N_16447,N_13804,N_14784);
nor U16448 (N_16448,N_13985,N_14653);
xor U16449 (N_16449,N_13807,N_14618);
or U16450 (N_16450,N_14183,N_14706);
nor U16451 (N_16451,N_14927,N_14763);
and U16452 (N_16452,N_13575,N_13543);
and U16453 (N_16453,N_13702,N_14378);
xnor U16454 (N_16454,N_14811,N_13913);
and U16455 (N_16455,N_14729,N_14184);
xnor U16456 (N_16456,N_13877,N_14360);
or U16457 (N_16457,N_14730,N_14384);
xnor U16458 (N_16458,N_13839,N_13867);
nand U16459 (N_16459,N_13870,N_14083);
and U16460 (N_16460,N_14172,N_14300);
nor U16461 (N_16461,N_14955,N_14743);
and U16462 (N_16462,N_13779,N_14796);
or U16463 (N_16463,N_14340,N_14675);
or U16464 (N_16464,N_14697,N_13701);
and U16465 (N_16465,N_14136,N_14032);
and U16466 (N_16466,N_14453,N_14945);
or U16467 (N_16467,N_14596,N_14277);
xor U16468 (N_16468,N_14700,N_13709);
nor U16469 (N_16469,N_14373,N_13577);
nor U16470 (N_16470,N_14441,N_13897);
xnor U16471 (N_16471,N_13500,N_14598);
or U16472 (N_16472,N_14123,N_14731);
nor U16473 (N_16473,N_13976,N_14499);
and U16474 (N_16474,N_14117,N_14353);
and U16475 (N_16475,N_14506,N_13553);
nand U16476 (N_16476,N_14665,N_14568);
nand U16477 (N_16477,N_14374,N_14934);
xor U16478 (N_16478,N_14730,N_13548);
xor U16479 (N_16479,N_14846,N_14596);
nand U16480 (N_16480,N_14570,N_14860);
xor U16481 (N_16481,N_13696,N_14990);
nand U16482 (N_16482,N_13566,N_14422);
xnor U16483 (N_16483,N_14813,N_14495);
nand U16484 (N_16484,N_13850,N_14306);
or U16485 (N_16485,N_13932,N_14937);
or U16486 (N_16486,N_14948,N_14351);
nand U16487 (N_16487,N_14611,N_13856);
xor U16488 (N_16488,N_14791,N_13974);
or U16489 (N_16489,N_13861,N_14676);
xor U16490 (N_16490,N_13710,N_14886);
or U16491 (N_16491,N_14232,N_14177);
or U16492 (N_16492,N_14742,N_14312);
nand U16493 (N_16493,N_14859,N_14193);
and U16494 (N_16494,N_14415,N_14197);
xor U16495 (N_16495,N_14188,N_14662);
xnor U16496 (N_16496,N_14686,N_14310);
xor U16497 (N_16497,N_14780,N_14791);
nor U16498 (N_16498,N_13816,N_14096);
and U16499 (N_16499,N_14707,N_14713);
nor U16500 (N_16500,N_16295,N_16248);
and U16501 (N_16501,N_15681,N_16129);
nor U16502 (N_16502,N_15621,N_15310);
xor U16503 (N_16503,N_15434,N_16164);
or U16504 (N_16504,N_15123,N_15215);
or U16505 (N_16505,N_15097,N_15820);
or U16506 (N_16506,N_15529,N_16304);
nor U16507 (N_16507,N_15856,N_15865);
nor U16508 (N_16508,N_16134,N_15635);
xor U16509 (N_16509,N_16458,N_15027);
nand U16510 (N_16510,N_16039,N_16476);
and U16511 (N_16511,N_15589,N_15798);
xor U16512 (N_16512,N_16328,N_15707);
and U16513 (N_16513,N_15976,N_16418);
or U16514 (N_16514,N_15204,N_16029);
nor U16515 (N_16515,N_16474,N_15673);
xor U16516 (N_16516,N_15609,N_16341);
and U16517 (N_16517,N_16371,N_15172);
nor U16518 (N_16518,N_15700,N_16048);
and U16519 (N_16519,N_15535,N_16235);
xnor U16520 (N_16520,N_15365,N_16176);
nand U16521 (N_16521,N_15925,N_15230);
or U16522 (N_16522,N_16465,N_15427);
or U16523 (N_16523,N_16080,N_15489);
or U16524 (N_16524,N_15362,N_15000);
or U16525 (N_16525,N_15580,N_15004);
xor U16526 (N_16526,N_15800,N_16490);
xor U16527 (N_16527,N_15418,N_15463);
xor U16528 (N_16528,N_15471,N_16043);
or U16529 (N_16529,N_15792,N_16147);
nor U16530 (N_16530,N_15674,N_16415);
and U16531 (N_16531,N_15268,N_15703);
and U16532 (N_16532,N_15931,N_15823);
or U16533 (N_16533,N_16107,N_16018);
and U16534 (N_16534,N_15387,N_16197);
xnor U16535 (N_16535,N_15554,N_15914);
xor U16536 (N_16536,N_15450,N_16188);
or U16537 (N_16537,N_16177,N_16209);
xor U16538 (N_16538,N_15235,N_15223);
nand U16539 (N_16539,N_15182,N_15544);
xnor U16540 (N_16540,N_15668,N_16244);
and U16541 (N_16541,N_15275,N_16060);
nor U16542 (N_16542,N_16492,N_15484);
or U16543 (N_16543,N_15407,N_15338);
and U16544 (N_16544,N_16215,N_16464);
nor U16545 (N_16545,N_15558,N_15730);
or U16546 (N_16546,N_16286,N_15494);
or U16547 (N_16547,N_15905,N_16243);
xor U16548 (N_16548,N_15632,N_15079);
nand U16549 (N_16549,N_15939,N_15826);
or U16550 (N_16550,N_15393,N_15634);
and U16551 (N_16551,N_15591,N_15744);
and U16552 (N_16552,N_15133,N_16130);
nand U16553 (N_16553,N_15884,N_15442);
and U16554 (N_16554,N_15664,N_15750);
xor U16555 (N_16555,N_15847,N_16241);
or U16556 (N_16556,N_16128,N_15107);
nand U16557 (N_16557,N_15736,N_15919);
xor U16558 (N_16558,N_16360,N_16472);
nor U16559 (N_16559,N_15641,N_16375);
nor U16560 (N_16560,N_16477,N_16449);
and U16561 (N_16561,N_15036,N_15678);
and U16562 (N_16562,N_16253,N_15957);
and U16563 (N_16563,N_15451,N_15212);
and U16564 (N_16564,N_16370,N_15390);
nor U16565 (N_16565,N_15031,N_15189);
nand U16566 (N_16566,N_15026,N_15155);
and U16567 (N_16567,N_15907,N_16228);
xor U16568 (N_16568,N_15560,N_16262);
xor U16569 (N_16569,N_16263,N_15017);
xor U16570 (N_16570,N_15758,N_16156);
nand U16571 (N_16571,N_15572,N_16162);
or U16572 (N_16572,N_15254,N_15687);
xor U16573 (N_16573,N_15523,N_15252);
and U16574 (N_16574,N_15785,N_15422);
or U16575 (N_16575,N_15950,N_16310);
nand U16576 (N_16576,N_15721,N_16206);
or U16577 (N_16577,N_15153,N_16416);
and U16578 (N_16578,N_15814,N_15679);
xor U16579 (N_16579,N_15633,N_15654);
and U16580 (N_16580,N_15500,N_15717);
nand U16581 (N_16581,N_16182,N_15915);
nand U16582 (N_16582,N_15685,N_15374);
or U16583 (N_16583,N_15571,N_15049);
and U16584 (N_16584,N_16017,N_16136);
and U16585 (N_16585,N_15977,N_16424);
nand U16586 (N_16586,N_15184,N_15762);
nor U16587 (N_16587,N_15663,N_16426);
nand U16588 (N_16588,N_16079,N_16186);
xor U16589 (N_16589,N_15052,N_15935);
or U16590 (N_16590,N_16051,N_15209);
nand U16591 (N_16591,N_15456,N_15199);
xor U16592 (N_16592,N_16436,N_15350);
or U16593 (N_16593,N_15849,N_15394);
nand U16594 (N_16594,N_15039,N_15329);
nor U16595 (N_16595,N_15183,N_15249);
xor U16596 (N_16596,N_15605,N_16352);
or U16597 (N_16597,N_15819,N_16234);
xor U16598 (N_16598,N_16109,N_15872);
and U16599 (N_16599,N_15431,N_15071);
nor U16600 (N_16600,N_15552,N_15247);
and U16601 (N_16601,N_16346,N_15768);
nor U16602 (N_16602,N_15793,N_15995);
or U16603 (N_16603,N_15846,N_15131);
nor U16604 (N_16604,N_16379,N_15485);
nand U16605 (N_16605,N_15502,N_15594);
or U16606 (N_16606,N_15293,N_15253);
or U16607 (N_16607,N_15412,N_15741);
and U16608 (N_16608,N_16331,N_15218);
nand U16609 (N_16609,N_16444,N_16383);
nor U16610 (N_16610,N_15076,N_15568);
nand U16611 (N_16611,N_16067,N_16287);
and U16612 (N_16612,N_15445,N_15666);
nand U16613 (N_16613,N_15963,N_15972);
nor U16614 (N_16614,N_15263,N_16343);
and U16615 (N_16615,N_16101,N_15448);
nor U16616 (N_16616,N_15816,N_16045);
xnor U16617 (N_16617,N_15619,N_16170);
and U16618 (N_16618,N_15453,N_15459);
xor U16619 (N_16619,N_15234,N_15283);
xnor U16620 (N_16620,N_16337,N_15034);
xnor U16621 (N_16621,N_15755,N_16314);
or U16622 (N_16622,N_15145,N_15292);
xor U16623 (N_16623,N_15288,N_15642);
nand U16624 (N_16624,N_16272,N_15531);
xnor U16625 (N_16625,N_16261,N_15159);
nand U16626 (N_16626,N_15369,N_16457);
nand U16627 (N_16627,N_15074,N_15020);
xor U16628 (N_16628,N_16489,N_16448);
nand U16629 (N_16629,N_16283,N_16126);
and U16630 (N_16630,N_15910,N_15070);
nor U16631 (N_16631,N_16013,N_15379);
xor U16632 (N_16632,N_15831,N_16431);
and U16633 (N_16633,N_15607,N_15615);
or U16634 (N_16634,N_16306,N_15216);
nor U16635 (N_16635,N_15754,N_15801);
nor U16636 (N_16636,N_15201,N_15059);
or U16637 (N_16637,N_15037,N_15930);
nor U16638 (N_16638,N_15862,N_15655);
nor U16639 (N_16639,N_15937,N_16471);
nand U16640 (N_16640,N_16180,N_16240);
nand U16641 (N_16641,N_16044,N_15991);
xnor U16642 (N_16642,N_16120,N_15723);
nand U16643 (N_16643,N_15437,N_15091);
nor U16644 (N_16644,N_16399,N_15761);
or U16645 (N_16645,N_16117,N_15001);
and U16646 (N_16646,N_15922,N_16497);
and U16647 (N_16647,N_15547,N_15063);
and U16648 (N_16648,N_15380,N_15728);
nor U16649 (N_16649,N_15129,N_15999);
or U16650 (N_16650,N_15804,N_15978);
xor U16651 (N_16651,N_16000,N_16347);
nor U16652 (N_16652,N_15051,N_15698);
xnor U16653 (N_16653,N_16211,N_15898);
and U16654 (N_16654,N_15233,N_15349);
nand U16655 (N_16655,N_15467,N_16221);
or U16656 (N_16656,N_15699,N_15725);
nor U16657 (N_16657,N_15312,N_15186);
nor U16658 (N_16658,N_15836,N_16456);
and U16659 (N_16659,N_16031,N_16482);
nor U16660 (N_16660,N_16294,N_15714);
nor U16661 (N_16661,N_15114,N_15841);
nand U16662 (N_16662,N_16023,N_15130);
and U16663 (N_16663,N_15858,N_15592);
xnor U16664 (N_16664,N_15938,N_15008);
xnor U16665 (N_16665,N_15060,N_15083);
or U16666 (N_16666,N_15340,N_15259);
xor U16667 (N_16667,N_15576,N_16096);
nor U16668 (N_16668,N_16259,N_15828);
and U16669 (N_16669,N_15118,N_15273);
xor U16670 (N_16670,N_15108,N_15289);
nor U16671 (N_16671,N_15324,N_15524);
nand U16672 (N_16672,N_15990,N_15953);
xnor U16673 (N_16673,N_16100,N_15111);
nand U16674 (N_16674,N_15444,N_15706);
nand U16675 (N_16675,N_15688,N_16394);
nand U16676 (N_16676,N_15251,N_15169);
and U16677 (N_16677,N_15239,N_15277);
and U16678 (N_16678,N_15006,N_16406);
and U16679 (N_16679,N_15142,N_15158);
or U16680 (N_16680,N_15584,N_15557);
or U16681 (N_16681,N_15339,N_15299);
and U16682 (N_16682,N_15086,N_16053);
nand U16683 (N_16683,N_15889,N_15763);
nand U16684 (N_16684,N_15843,N_15261);
or U16685 (N_16685,N_15942,N_16203);
or U16686 (N_16686,N_15748,N_15177);
nor U16687 (N_16687,N_15505,N_16391);
or U16688 (N_16688,N_15737,N_15473);
nand U16689 (N_16689,N_15135,N_16099);
nand U16690 (N_16690,N_15784,N_16493);
or U16691 (N_16691,N_15848,N_16010);
and U16692 (N_16692,N_15775,N_16297);
nand U16693 (N_16693,N_15401,N_16007);
nand U16694 (N_16694,N_16168,N_16321);
xnor U16695 (N_16695,N_16196,N_15711);
xor U16696 (N_16696,N_16074,N_15503);
or U16697 (N_16697,N_15316,N_16305);
nor U16698 (N_16698,N_15481,N_15803);
and U16699 (N_16699,N_15466,N_15868);
or U16700 (N_16700,N_15890,N_15626);
nor U16701 (N_16701,N_15805,N_16423);
nor U16702 (N_16702,N_15024,N_15912);
and U16703 (N_16703,N_15886,N_15320);
and U16704 (N_16704,N_15274,N_16059);
nand U16705 (N_16705,N_15948,N_16325);
nor U16706 (N_16706,N_16082,N_15092);
xor U16707 (N_16707,N_15246,N_15656);
nand U16708 (N_16708,N_16288,N_15970);
nand U16709 (N_16709,N_16086,N_15945);
and U16710 (N_16710,N_16374,N_15636);
nor U16711 (N_16711,N_15331,N_16027);
nand U16712 (N_16712,N_15265,N_15009);
nor U16713 (N_16713,N_15840,N_15732);
nand U16714 (N_16714,N_15423,N_15867);
or U16715 (N_16715,N_15242,N_15810);
xnor U16716 (N_16716,N_16428,N_15787);
nor U16717 (N_16717,N_15593,N_15326);
and U16718 (N_16718,N_16293,N_15900);
or U16719 (N_16719,N_15478,N_16143);
nor U16720 (N_16720,N_15295,N_15376);
and U16721 (N_16721,N_15885,N_15993);
and U16722 (N_16722,N_15082,N_16388);
and U16723 (N_16723,N_16372,N_16118);
xnor U16724 (N_16724,N_15345,N_15157);
or U16725 (N_16725,N_15777,N_16189);
or U16726 (N_16726,N_16202,N_15967);
or U16727 (N_16727,N_16068,N_16403);
or U16728 (N_16728,N_16466,N_15852);
nand U16729 (N_16729,N_16145,N_15100);
nor U16730 (N_16730,N_15838,N_15837);
and U16731 (N_16731,N_16122,N_16105);
and U16732 (N_16732,N_15469,N_15802);
nor U16733 (N_16733,N_15460,N_15113);
nor U16734 (N_16734,N_15644,N_16382);
nand U16735 (N_16735,N_16095,N_15416);
and U16736 (N_16736,N_15257,N_15743);
nor U16737 (N_16737,N_15487,N_16098);
nor U16738 (N_16738,N_15400,N_16158);
or U16739 (N_16739,N_15417,N_16408);
nor U16740 (N_16740,N_15996,N_15014);
and U16741 (N_16741,N_16173,N_16378);
or U16742 (N_16742,N_16194,N_15109);
and U16743 (N_16743,N_15695,N_15294);
nor U16744 (N_16744,N_16016,N_15960);
xnor U16745 (N_16745,N_16455,N_16273);
xor U16746 (N_16746,N_15704,N_16227);
or U16747 (N_16747,N_15361,N_16055);
nand U16748 (N_16748,N_16367,N_16350);
xor U16749 (N_16749,N_15395,N_16160);
nand U16750 (N_16750,N_15906,N_15101);
xnor U16751 (N_16751,N_15335,N_15812);
and U16752 (N_16752,N_15541,N_15149);
or U16753 (N_16753,N_16470,N_15659);
xnor U16754 (N_16754,N_16069,N_15860);
xnor U16755 (N_16755,N_16121,N_16264);
or U16756 (N_16756,N_15224,N_15569);
nor U16757 (N_16757,N_16052,N_15264);
nand U16758 (N_16758,N_15982,N_15077);
nor U16759 (N_16759,N_15435,N_16387);
and U16760 (N_16760,N_15797,N_15389);
or U16761 (N_16761,N_15173,N_15047);
or U16762 (N_16762,N_15297,N_15165);
and U16763 (N_16763,N_15513,N_15064);
and U16764 (N_16764,N_15296,N_15864);
or U16765 (N_16765,N_16441,N_15232);
or U16766 (N_16766,N_16112,N_15778);
and U16767 (N_16767,N_16401,N_16094);
nor U16768 (N_16768,N_16024,N_15934);
xor U16769 (N_16769,N_16410,N_16038);
and U16770 (N_16770,N_15574,N_15432);
and U16771 (N_16771,N_16199,N_16004);
or U16772 (N_16772,N_16389,N_15764);
or U16773 (N_16773,N_15794,N_15044);
xor U16774 (N_16774,N_16340,N_16106);
xor U16775 (N_16775,N_15021,N_16002);
nand U16776 (N_16776,N_15282,N_15861);
or U16777 (N_16777,N_16127,N_15088);
or U16778 (N_16778,N_15065,N_15590);
nor U16779 (N_16779,N_15090,N_15166);
xnor U16780 (N_16780,N_15783,N_16278);
nand U16781 (N_16781,N_16056,N_16460);
or U16782 (N_16782,N_15197,N_15742);
and U16783 (N_16783,N_15105,N_15951);
nor U16784 (N_16784,N_16439,N_16047);
nor U16785 (N_16785,N_15933,N_16414);
and U16786 (N_16786,N_16015,N_15646);
xnor U16787 (N_16787,N_15038,N_16208);
xnor U16788 (N_16788,N_16386,N_15128);
xor U16789 (N_16789,N_15328,N_15344);
or U16790 (N_16790,N_15303,N_15112);
xnor U16791 (N_16791,N_16397,N_15102);
nand U16792 (N_16792,N_15306,N_16001);
and U16793 (N_16793,N_15276,N_16246);
nor U16794 (N_16794,N_15308,N_15458);
and U16795 (N_16795,N_15756,N_15504);
or U16796 (N_16796,N_15883,N_15206);
or U16797 (N_16797,N_15573,N_15551);
xnor U16798 (N_16798,N_15893,N_15488);
and U16799 (N_16799,N_15924,N_15392);
xor U16800 (N_16800,N_16192,N_15710);
nand U16801 (N_16801,N_15521,N_16054);
or U16802 (N_16802,N_15262,N_15989);
nand U16803 (N_16803,N_15103,N_16110);
nor U16804 (N_16804,N_15490,N_16220);
nand U16805 (N_16805,N_15538,N_15309);
xor U16806 (N_16806,N_15405,N_16300);
or U16807 (N_16807,N_16012,N_15733);
nand U16808 (N_16808,N_15355,N_15586);
or U16809 (N_16809,N_15583,N_16338);
nor U16810 (N_16810,N_16357,N_16429);
nor U16811 (N_16811,N_15588,N_15154);
nor U16812 (N_16812,N_15378,N_15319);
nor U16813 (N_16813,N_16213,N_15385);
and U16814 (N_16814,N_15360,N_15825);
and U16815 (N_16815,N_15645,N_15772);
and U16816 (N_16816,N_15542,N_15845);
xnor U16817 (N_16817,N_16050,N_16201);
and U16818 (N_16818,N_15483,N_16488);
and U16819 (N_16819,N_15667,N_15766);
nor U16820 (N_16820,N_16184,N_15622);
xor U16821 (N_16821,N_16361,N_15724);
nand U16822 (N_16822,N_15514,N_15480);
nand U16823 (N_16823,N_15256,N_15440);
nand U16824 (N_16824,N_15429,N_15002);
xnor U16825 (N_16825,N_16393,N_15863);
and U16826 (N_16826,N_16225,N_15353);
and U16827 (N_16827,N_15871,N_15409);
nor U16828 (N_16828,N_15833,N_16487);
or U16829 (N_16829,N_15318,N_15943);
xor U16830 (N_16830,N_15809,N_15124);
nand U16831 (N_16831,N_15786,N_15152);
nand U16832 (N_16832,N_15015,N_16046);
or U16833 (N_16833,N_15075,N_16285);
or U16834 (N_16834,N_15870,N_15979);
nand U16835 (N_16835,N_15835,N_15896);
nor U16836 (N_16836,N_15888,N_16445);
nand U16837 (N_16837,N_16422,N_15200);
nor U16838 (N_16838,N_15438,N_15348);
and U16839 (N_16839,N_15992,N_16237);
nand U16840 (N_16840,N_15769,N_15988);
xnor U16841 (N_16841,N_16485,N_15477);
and U16842 (N_16842,N_16443,N_15271);
nand U16843 (N_16843,N_16475,N_16042);
nand U16844 (N_16844,N_15507,N_15903);
nand U16845 (N_16845,N_15726,N_15962);
and U16846 (N_16846,N_15098,N_15985);
or U16847 (N_16847,N_15272,N_16159);
nand U16848 (N_16848,N_15528,N_16231);
or U16849 (N_16849,N_15419,N_15660);
xnor U16850 (N_16850,N_15791,N_15702);
xor U16851 (N_16851,N_16155,N_16473);
and U16852 (N_16852,N_15881,N_15045);
or U16853 (N_16853,N_15508,N_16033);
nor U16854 (N_16854,N_15649,N_15773);
xnor U16855 (N_16855,N_15258,N_15637);
xor U16856 (N_16856,N_15638,N_15604);
or U16857 (N_16857,N_15640,N_16268);
nand U16858 (N_16858,N_16185,N_15243);
nor U16859 (N_16859,N_15997,N_16179);
or U16860 (N_16860,N_15094,N_16413);
or U16861 (N_16861,N_15519,N_15482);
or U16862 (N_16862,N_16362,N_16355);
nand U16863 (N_16863,N_15747,N_16483);
nor U16864 (N_16864,N_15902,N_15661);
xnor U16865 (N_16865,N_15342,N_15601);
nand U16866 (N_16866,N_15869,N_15603);
and U16867 (N_16867,N_16409,N_15163);
nor U16868 (N_16868,N_16030,N_15449);
or U16869 (N_16869,N_15373,N_16430);
nand U16870 (N_16870,N_15366,N_15813);
and U16871 (N_16871,N_16486,N_15752);
xnor U16872 (N_16872,N_16142,N_16032);
or U16873 (N_16873,N_16022,N_15940);
nor U16874 (N_16874,N_16103,N_15399);
xnor U16875 (N_16875,N_15084,N_15596);
nand U16876 (N_16876,N_15713,N_15517);
nand U16877 (N_16877,N_15696,N_15620);
or U16878 (N_16878,N_16435,N_15248);
and U16879 (N_16879,N_15509,N_15032);
nand U16880 (N_16880,N_16267,N_15170);
or U16881 (N_16881,N_15069,N_16075);
nor U16882 (N_16882,N_15965,N_15187);
or U16883 (N_16883,N_16169,N_15443);
or U16884 (N_16884,N_16425,N_16006);
xnor U16885 (N_16885,N_15211,N_15479);
nand U16886 (N_16886,N_15190,N_16421);
xnor U16887 (N_16887,N_15375,N_15117);
xor U16888 (N_16888,N_15245,N_15739);
xnor U16889 (N_16889,N_15238,N_15352);
nand U16890 (N_16890,N_15959,N_15221);
and U16891 (N_16891,N_16276,N_15073);
nand U16892 (N_16892,N_16452,N_15096);
and U16893 (N_16893,N_16318,N_16195);
and U16894 (N_16894,N_15266,N_16308);
xnor U16895 (N_16895,N_15854,N_15857);
and U16896 (N_16896,N_15625,N_15624);
xnor U16897 (N_16897,N_15217,N_15746);
xnor U16898 (N_16898,N_15610,N_15735);
xor U16899 (N_16899,N_15617,N_15298);
xnor U16900 (N_16900,N_15677,N_15354);
nor U16901 (N_16901,N_15139,N_15827);
xor U16902 (N_16902,N_16411,N_16217);
xor U16903 (N_16903,N_16141,N_15821);
or U16904 (N_16904,N_16292,N_15194);
or U16905 (N_16905,N_15780,N_15291);
or U16906 (N_16906,N_16333,N_16066);
xor U16907 (N_16907,N_15424,N_16003);
nor U16908 (N_16908,N_16254,N_16041);
xnor U16909 (N_16909,N_16146,N_16214);
or U16910 (N_16910,N_15525,N_15562);
nand U16911 (N_16911,N_16467,N_15140);
or U16912 (N_16912,N_15359,N_15498);
xnor U16913 (N_16913,N_15347,N_15382);
or U16914 (N_16914,N_16124,N_16161);
nand U16915 (N_16915,N_16332,N_15612);
nor U16916 (N_16916,N_15964,N_15413);
xor U16917 (N_16917,N_16366,N_15279);
and U16918 (N_16918,N_15202,N_16395);
or U16919 (N_16919,N_15441,N_16137);
xnor U16920 (N_16920,N_16420,N_15048);
or U16921 (N_16921,N_15311,N_15122);
or U16922 (N_16922,N_16165,N_15408);
or U16923 (N_16923,N_15493,N_15824);
or U16924 (N_16924,N_16326,N_15404);
or U16925 (N_16925,N_15520,N_15333);
nor U16926 (N_16926,N_15901,N_15046);
nor U16927 (N_16927,N_15402,N_15946);
xor U16928 (N_16928,N_15533,N_15198);
and U16929 (N_16929,N_15410,N_16363);
and U16930 (N_16930,N_15949,N_16219);
nor U16931 (N_16931,N_16076,N_16365);
nor U16932 (N_16932,N_16200,N_16187);
nor U16933 (N_16933,N_16085,N_16178);
or U16934 (N_16934,N_16339,N_16174);
nand U16935 (N_16935,N_16083,N_16353);
xor U16936 (N_16936,N_16073,N_16139);
or U16937 (N_16937,N_16131,N_15127);
or U16938 (N_16938,N_15377,N_16284);
nor U16939 (N_16939,N_16432,N_16390);
or U16940 (N_16940,N_15120,N_15357);
nor U16941 (N_16941,N_15658,N_15231);
and U16942 (N_16942,N_16373,N_15143);
or U16943 (N_16943,N_15025,N_16437);
nor U16944 (N_16944,N_15151,N_15829);
nor U16945 (N_16945,N_15691,N_15952);
and U16946 (N_16946,N_15341,N_16020);
and U16947 (N_16947,N_15068,N_16057);
or U16948 (N_16948,N_15080,N_15403);
xor U16949 (N_16949,N_16229,N_15817);
and U16950 (N_16950,N_16058,N_16021);
or U16951 (N_16951,N_16070,N_15866);
xnor U16952 (N_16952,N_16205,N_15926);
nor U16953 (N_16953,N_16289,N_15629);
xor U16954 (N_16954,N_15581,N_15180);
or U16955 (N_16955,N_16078,N_15536);
or U16956 (N_16956,N_15358,N_16065);
nor U16957 (N_16957,N_16438,N_16291);
nor U16958 (N_16958,N_15219,N_15411);
nor U16959 (N_16959,N_15566,N_15555);
or U16960 (N_16960,N_16171,N_15757);
nand U16961 (N_16961,N_16125,N_15005);
xor U16962 (N_16962,N_15213,N_15731);
or U16963 (N_16963,N_16218,N_15530);
xor U16964 (N_16964,N_16089,N_16479);
nor U16965 (N_16965,N_16364,N_15899);
or U16966 (N_16966,N_16335,N_15892);
nand U16967 (N_16967,N_15878,N_15606);
nand U16968 (N_16968,N_15539,N_16062);
nand U16969 (N_16969,N_15278,N_15806);
nand U16970 (N_16970,N_15388,N_15011);
nor U16971 (N_16971,N_16299,N_15973);
nand U16972 (N_16972,N_15280,N_16025);
xnor U16973 (N_16973,N_15210,N_15880);
xor U16974 (N_16974,N_15381,N_15150);
or U16975 (N_16975,N_15672,N_15475);
xor U16976 (N_16976,N_16138,N_15121);
or U16977 (N_16977,N_15134,N_15771);
nor U16978 (N_16978,N_16064,N_16207);
nor U16979 (N_16979,N_15585,N_15690);
nand U16980 (N_16980,N_16320,N_15030);
and U16981 (N_16981,N_15904,N_15141);
xor U16982 (N_16982,N_16484,N_16348);
nand U16983 (N_16983,N_16434,N_15597);
nand U16984 (N_16984,N_15684,N_15176);
or U16985 (N_16985,N_15874,N_15174);
nand U16986 (N_16986,N_16344,N_15491);
xor U16987 (N_16987,N_15639,N_15708);
or U16988 (N_16988,N_16190,N_15987);
nand U16989 (N_16989,N_16412,N_15851);
nand U16990 (N_16990,N_15662,N_16226);
xor U16991 (N_16991,N_16359,N_16102);
xnor U16992 (N_16992,N_16249,N_15932);
nor U16993 (N_16993,N_15470,N_15089);
and U16994 (N_16994,N_15760,N_15877);
xor U16995 (N_16995,N_15225,N_15853);
xor U16996 (N_16996,N_16324,N_16036);
xor U16997 (N_16997,N_16149,N_15323);
or U16998 (N_16998,N_16097,N_15164);
and U16999 (N_16999,N_15226,N_15955);
xor U17000 (N_17000,N_15236,N_15168);
or U17001 (N_17001,N_16334,N_15830);
xnor U17002 (N_17002,N_15099,N_15729);
xnor U17003 (N_17003,N_16212,N_15058);
and U17004 (N_17004,N_16407,N_16459);
nor U17005 (N_17005,N_15879,N_16224);
nand U17006 (N_17006,N_15446,N_16404);
or U17007 (N_17007,N_15587,N_16302);
xor U17008 (N_17008,N_15921,N_15575);
xnor U17009 (N_17009,N_16108,N_16084);
nor U17010 (N_17010,N_16009,N_15119);
or U17011 (N_17011,N_16495,N_15284);
nand U17012 (N_17012,N_15414,N_16274);
nand U17013 (N_17013,N_15332,N_15969);
and U17014 (N_17014,N_15104,N_15720);
nor U17015 (N_17015,N_15767,N_16081);
xor U17016 (N_17016,N_15651,N_15795);
nand U17017 (N_17017,N_15087,N_15162);
xor U17018 (N_17018,N_15623,N_15185);
or U17019 (N_17019,N_16317,N_16153);
xor U17020 (N_17020,N_15260,N_16247);
nor U17021 (N_17021,N_16316,N_15671);
nor U17022 (N_17022,N_15630,N_15526);
nand U17023 (N_17023,N_15205,N_16035);
xnor U17024 (N_17024,N_15578,N_15454);
nand U17025 (N_17025,N_15281,N_16061);
and U17026 (N_17026,N_15913,N_15314);
xnor U17027 (N_17027,N_15023,N_16150);
xor U17028 (N_17028,N_15718,N_15304);
or U17029 (N_17029,N_15709,N_15582);
nor U17030 (N_17030,N_16133,N_15439);
xor U17031 (N_17031,N_15550,N_16392);
xnor U17032 (N_17032,N_15669,N_15193);
xnor U17033 (N_17033,N_15497,N_15895);
nor U17034 (N_17034,N_16400,N_15693);
xor U17035 (N_17035,N_15269,N_15776);
nor U17036 (N_17036,N_15749,N_16480);
and U17037 (N_17037,N_16315,N_15286);
nand U17038 (N_17038,N_15447,N_15564);
nand U17039 (N_17039,N_16468,N_15315);
and U17040 (N_17040,N_15191,N_15781);
xnor U17041 (N_17041,N_15697,N_16384);
and U17042 (N_17042,N_16376,N_16063);
nand U17043 (N_17043,N_15160,N_15181);
nor U17044 (N_17044,N_15897,N_15522);
and U17045 (N_17045,N_16323,N_16114);
or U17046 (N_17046,N_15822,N_15018);
nand U17047 (N_17047,N_15941,N_16269);
and U17048 (N_17048,N_15686,N_15106);
or U17049 (N_17049,N_15611,N_15613);
nor U17050 (N_17050,N_16322,N_15506);
nor U17051 (N_17051,N_15337,N_15370);
nand U17052 (N_17052,N_16183,N_15975);
or U17053 (N_17053,N_15873,N_15270);
nor U17054 (N_17054,N_16223,N_16026);
and U17055 (N_17055,N_15705,N_15543);
or U17056 (N_17056,N_15534,N_16312);
xor U17057 (N_17057,N_15753,N_16233);
nand U17058 (N_17058,N_15692,N_16256);
and U17059 (N_17059,N_16349,N_16311);
xnor U17060 (N_17060,N_16071,N_16402);
xnor U17061 (N_17061,N_16281,N_15476);
nor U17062 (N_17062,N_16282,N_15927);
or U17063 (N_17063,N_15330,N_15727);
nand U17064 (N_17064,N_15627,N_15518);
and U17065 (N_17065,N_15958,N_16451);
and U17066 (N_17066,N_15653,N_15715);
or U17067 (N_17067,N_16238,N_15192);
nand U17068 (N_17068,N_15834,N_16258);
or U17069 (N_17069,N_15909,N_16005);
nand U17070 (N_17070,N_15689,N_15042);
xor U17071 (N_17071,N_16087,N_15428);
or U17072 (N_17072,N_15003,N_15033);
nand U17073 (N_17073,N_15474,N_15516);
nor U17074 (N_17074,N_15559,N_15055);
nand U17075 (N_17075,N_15406,N_16446);
or U17076 (N_17076,N_16132,N_16191);
xor U17077 (N_17077,N_15894,N_16148);
and U17078 (N_17078,N_15712,N_16204);
and U17079 (N_17079,N_15928,N_15195);
and U17080 (N_17080,N_16330,N_15515);
nor U17081 (N_17081,N_15598,N_15436);
and U17082 (N_17082,N_16345,N_16239);
nand U17083 (N_17083,N_15455,N_15132);
nand U17084 (N_17084,N_16252,N_15188);
xor U17085 (N_17085,N_15178,N_15844);
nand U17086 (N_17086,N_15010,N_16427);
and U17087 (N_17087,N_15237,N_15062);
and U17088 (N_17088,N_16385,N_15167);
or U17089 (N_17089,N_15486,N_15998);
nor U17090 (N_17090,N_16037,N_15556);
nor U17091 (N_17091,N_16154,N_16469);
and U17092 (N_17092,N_15499,N_15567);
or U17093 (N_17093,N_16104,N_15956);
xor U17094 (N_17094,N_16313,N_16250);
or U17095 (N_17095,N_16419,N_15452);
and U17096 (N_17096,N_15790,N_16232);
or U17097 (N_17097,N_15954,N_15061);
nand U17098 (N_17098,N_15676,N_16336);
nand U17099 (N_17099,N_16478,N_15839);
xor U17100 (N_17100,N_15765,N_16144);
nor U17101 (N_17101,N_15057,N_15287);
or U17102 (N_17102,N_15983,N_15179);
nor U17103 (N_17103,N_15430,N_16222);
xor U17104 (N_17104,N_15631,N_15807);
nand U17105 (N_17105,N_15398,N_16461);
xor U17106 (N_17106,N_16275,N_16210);
nor U17107 (N_17107,N_16088,N_16091);
xor U17108 (N_17108,N_16491,N_16280);
and U17109 (N_17109,N_15019,N_15774);
nor U17110 (N_17110,N_16260,N_15643);
and U17111 (N_17111,N_15054,N_16111);
nor U17112 (N_17112,N_15918,N_15229);
nand U17113 (N_17113,N_15994,N_15012);
nand U17114 (N_17114,N_15250,N_16198);
nand U17115 (N_17115,N_15680,N_16040);
and U17116 (N_17116,N_15616,N_15433);
or U17117 (N_17117,N_15156,N_15072);
and U17118 (N_17118,N_15093,N_16296);
or U17119 (N_17119,N_15563,N_16354);
nand U17120 (N_17120,N_15396,N_16236);
xnor U17121 (N_17121,N_16307,N_16157);
xor U17122 (N_17122,N_16242,N_16442);
and U17123 (N_17123,N_15908,N_15734);
or U17124 (N_17124,N_16358,N_16279);
xnor U17125 (N_17125,N_16381,N_15196);
and U17126 (N_17126,N_15980,N_15115);
nor U17127 (N_17127,N_15788,N_15016);
or U17128 (N_17128,N_16277,N_15495);
or U17129 (N_17129,N_15136,N_15244);
nor U17130 (N_17130,N_16034,N_15468);
or U17131 (N_17131,N_15599,N_15968);
nor U17132 (N_17132,N_16123,N_16433);
and U17133 (N_17133,N_15028,N_15220);
nor U17134 (N_17134,N_16342,N_15947);
nor U17135 (N_17135,N_15929,N_15779);
nor U17136 (N_17136,N_15850,N_15035);
xor U17137 (N_17137,N_16166,N_15799);
nand U17138 (N_17138,N_15647,N_15738);
or U17139 (N_17139,N_15383,N_15618);
and U17140 (N_17140,N_16351,N_15040);
nand U17141 (N_17141,N_15501,N_15561);
or U17142 (N_17142,N_15138,N_15683);
or U17143 (N_17143,N_15759,N_15971);
nor U17144 (N_17144,N_15657,N_15511);
and U17145 (N_17145,N_15415,N_16216);
and U17146 (N_17146,N_16113,N_16140);
or U17147 (N_17147,N_16356,N_15214);
nand U17148 (N_17148,N_16405,N_16319);
xnor U17149 (N_17149,N_15917,N_16290);
nand U17150 (N_17150,N_15420,N_15161);
nor U17151 (N_17151,N_15981,N_16175);
nand U17152 (N_17152,N_16303,N_15148);
nand U17153 (N_17153,N_15371,N_15384);
nor U17154 (N_17154,N_15125,N_15363);
or U17155 (N_17155,N_15855,N_15175);
or U17156 (N_17156,N_15570,N_16049);
and U17157 (N_17157,N_16167,N_15670);
nor U17158 (N_17158,N_16301,N_15527);
nor U17159 (N_17159,N_15322,N_16019);
and U17160 (N_17160,N_15464,N_16008);
nor U17161 (N_17161,N_16135,N_16115);
nand U17162 (N_17162,N_15628,N_15078);
nand U17163 (N_17163,N_15789,N_15095);
nand U17164 (N_17164,N_15565,N_16257);
xor U17165 (N_17165,N_15984,N_15911);
or U17166 (N_17166,N_15346,N_15961);
or U17167 (N_17167,N_15832,N_15029);
and U17168 (N_17168,N_15462,N_15203);
xor U17169 (N_17169,N_15336,N_16152);
nor U17170 (N_17170,N_15545,N_15317);
or U17171 (N_17171,N_15540,N_15327);
xnor U17172 (N_17172,N_16417,N_15240);
nor U17173 (N_17173,N_15421,N_15325);
or U17174 (N_17174,N_16072,N_15472);
xor U17175 (N_17175,N_15465,N_15305);
and U17176 (N_17176,N_16309,N_16447);
nand U17177 (N_17177,N_16396,N_15056);
or U17178 (N_17178,N_16193,N_15842);
nand U17179 (N_17179,N_15875,N_15770);
nand U17180 (N_17180,N_15255,N_16454);
or U17181 (N_17181,N_16172,N_15923);
nor U17182 (N_17182,N_16251,N_15207);
nor U17183 (N_17183,N_16499,N_16092);
nand U17184 (N_17184,N_15652,N_15876);
nand U17185 (N_17185,N_15208,N_16453);
xor U17186 (N_17186,N_15887,N_15579);
nor U17187 (N_17187,N_15085,N_15300);
nand U17188 (N_17188,N_15313,N_15321);
nand U17189 (N_17189,N_15228,N_15936);
or U17190 (N_17190,N_16450,N_15882);
xor U17191 (N_17191,N_16028,N_15144);
nand U17192 (N_17192,N_15510,N_15457);
or U17193 (N_17193,N_15920,N_15859);
xnor U17194 (N_17194,N_15818,N_15351);
and U17195 (N_17195,N_15301,N_15577);
nand U17196 (N_17196,N_16496,N_16380);
and U17197 (N_17197,N_15966,N_15290);
or U17198 (N_17198,N_15307,N_15367);
nand U17199 (N_17199,N_16270,N_15595);
nand U17200 (N_17200,N_15368,N_15067);
or U17201 (N_17201,N_16265,N_16481);
or U17202 (N_17202,N_15302,N_15492);
nor U17203 (N_17203,N_15553,N_15682);
or U17204 (N_17204,N_15386,N_15397);
nand U17205 (N_17205,N_15512,N_16440);
and U17206 (N_17206,N_15648,N_15796);
or U17207 (N_17207,N_15461,N_15053);
xnor U17208 (N_17208,N_15222,N_15391);
or U17209 (N_17209,N_16151,N_15716);
nor U17210 (N_17210,N_15537,N_15372);
nand U17211 (N_17211,N_16093,N_15343);
nor U17212 (N_17212,N_15650,N_15126);
nand U17213 (N_17213,N_15891,N_16119);
nand U17214 (N_17214,N_15986,N_16011);
or U17215 (N_17215,N_15614,N_15608);
nand U17216 (N_17216,N_15974,N_15043);
nor U17217 (N_17217,N_16077,N_15600);
xor U17218 (N_17218,N_15694,N_15081);
nand U17219 (N_17219,N_16327,N_15701);
and U17220 (N_17220,N_15602,N_15425);
nand U17221 (N_17221,N_16245,N_15815);
xor U17222 (N_17222,N_15171,N_15285);
xnor U17223 (N_17223,N_15548,N_16462);
and U17224 (N_17224,N_16014,N_15782);
or U17225 (N_17225,N_15751,N_16255);
xor U17226 (N_17226,N_15007,N_15719);
nor U17227 (N_17227,N_15116,N_15137);
and U17228 (N_17228,N_16377,N_15808);
nand U17229 (N_17229,N_15146,N_15811);
xnor U17230 (N_17230,N_15334,N_15364);
nor U17231 (N_17231,N_16498,N_15041);
and U17232 (N_17232,N_15496,N_16230);
nor U17233 (N_17233,N_15241,N_15227);
nor U17234 (N_17234,N_15267,N_15426);
nor U17235 (N_17235,N_15944,N_15013);
nand U17236 (N_17236,N_16369,N_16329);
and U17237 (N_17237,N_15147,N_15665);
nand U17238 (N_17238,N_16494,N_15110);
nand U17239 (N_17239,N_16116,N_16090);
nor U17240 (N_17240,N_15740,N_15066);
nand U17241 (N_17241,N_16298,N_16398);
and U17242 (N_17242,N_16181,N_15050);
and U17243 (N_17243,N_16266,N_16463);
and U17244 (N_17244,N_15546,N_15916);
xor U17245 (N_17245,N_15549,N_15356);
nand U17246 (N_17246,N_15675,N_16271);
or U17247 (N_17247,N_16368,N_15745);
xnor U17248 (N_17248,N_16163,N_15722);
and U17249 (N_17249,N_15532,N_15022);
or U17250 (N_17250,N_16323,N_15907);
and U17251 (N_17251,N_15707,N_15692);
nand U17252 (N_17252,N_15757,N_15837);
or U17253 (N_17253,N_16062,N_16223);
nand U17254 (N_17254,N_16101,N_15428);
and U17255 (N_17255,N_15185,N_15186);
and U17256 (N_17256,N_15334,N_15902);
xor U17257 (N_17257,N_15514,N_15784);
xor U17258 (N_17258,N_15991,N_16100);
or U17259 (N_17259,N_15302,N_15548);
nand U17260 (N_17260,N_16029,N_15104);
and U17261 (N_17261,N_15524,N_15600);
nand U17262 (N_17262,N_16018,N_15080);
nand U17263 (N_17263,N_16015,N_15114);
and U17264 (N_17264,N_15522,N_15778);
xnor U17265 (N_17265,N_16206,N_16322);
or U17266 (N_17266,N_15289,N_16217);
or U17267 (N_17267,N_16079,N_15714);
nand U17268 (N_17268,N_15302,N_16220);
nor U17269 (N_17269,N_16354,N_16471);
and U17270 (N_17270,N_16193,N_15446);
and U17271 (N_17271,N_16378,N_16351);
xor U17272 (N_17272,N_15385,N_16233);
nor U17273 (N_17273,N_16103,N_15888);
nor U17274 (N_17274,N_15765,N_16409);
nand U17275 (N_17275,N_15955,N_16292);
and U17276 (N_17276,N_16463,N_15182);
nand U17277 (N_17277,N_15213,N_15967);
xor U17278 (N_17278,N_16014,N_16274);
nand U17279 (N_17279,N_16128,N_15390);
nand U17280 (N_17280,N_15444,N_15245);
or U17281 (N_17281,N_16105,N_15095);
and U17282 (N_17282,N_15305,N_15086);
nand U17283 (N_17283,N_15798,N_15710);
nor U17284 (N_17284,N_16448,N_15121);
or U17285 (N_17285,N_16411,N_15460);
and U17286 (N_17286,N_16186,N_15497);
and U17287 (N_17287,N_15071,N_15007);
and U17288 (N_17288,N_15830,N_15094);
or U17289 (N_17289,N_15227,N_15385);
nand U17290 (N_17290,N_16017,N_15506);
or U17291 (N_17291,N_15860,N_15272);
xnor U17292 (N_17292,N_15346,N_16429);
or U17293 (N_17293,N_15229,N_15721);
or U17294 (N_17294,N_16439,N_15442);
xor U17295 (N_17295,N_15065,N_16238);
or U17296 (N_17296,N_16499,N_15350);
xnor U17297 (N_17297,N_16128,N_16059);
xor U17298 (N_17298,N_15329,N_16361);
or U17299 (N_17299,N_16150,N_15328);
or U17300 (N_17300,N_15088,N_15577);
nor U17301 (N_17301,N_16470,N_16435);
xor U17302 (N_17302,N_16335,N_15006);
and U17303 (N_17303,N_15285,N_15617);
and U17304 (N_17304,N_16380,N_15349);
xor U17305 (N_17305,N_16457,N_16327);
or U17306 (N_17306,N_15253,N_16481);
or U17307 (N_17307,N_16096,N_16113);
nor U17308 (N_17308,N_15035,N_15986);
xnor U17309 (N_17309,N_15325,N_15794);
or U17310 (N_17310,N_15156,N_16319);
nor U17311 (N_17311,N_15910,N_15482);
and U17312 (N_17312,N_15520,N_15980);
nand U17313 (N_17313,N_16155,N_15864);
or U17314 (N_17314,N_15758,N_15383);
or U17315 (N_17315,N_15858,N_15941);
or U17316 (N_17316,N_15118,N_15733);
xor U17317 (N_17317,N_15433,N_15744);
nor U17318 (N_17318,N_15406,N_15436);
nand U17319 (N_17319,N_16325,N_15174);
nand U17320 (N_17320,N_16014,N_16087);
xnor U17321 (N_17321,N_15146,N_15822);
and U17322 (N_17322,N_15835,N_15396);
nand U17323 (N_17323,N_16262,N_15111);
nor U17324 (N_17324,N_16086,N_15034);
xnor U17325 (N_17325,N_15527,N_15578);
and U17326 (N_17326,N_15280,N_15457);
or U17327 (N_17327,N_15684,N_15842);
nor U17328 (N_17328,N_16458,N_15507);
nand U17329 (N_17329,N_15158,N_15467);
and U17330 (N_17330,N_15064,N_15309);
and U17331 (N_17331,N_16143,N_15937);
nand U17332 (N_17332,N_16045,N_15949);
nor U17333 (N_17333,N_16055,N_15404);
or U17334 (N_17334,N_15739,N_15918);
xor U17335 (N_17335,N_15176,N_16324);
or U17336 (N_17336,N_16177,N_15624);
xor U17337 (N_17337,N_15791,N_16361);
or U17338 (N_17338,N_15379,N_15421);
or U17339 (N_17339,N_16066,N_16496);
and U17340 (N_17340,N_16433,N_15739);
xnor U17341 (N_17341,N_16134,N_15080);
xor U17342 (N_17342,N_16473,N_15872);
and U17343 (N_17343,N_15197,N_15824);
nand U17344 (N_17344,N_16011,N_15786);
xor U17345 (N_17345,N_15365,N_16076);
nor U17346 (N_17346,N_15717,N_15179);
or U17347 (N_17347,N_15918,N_16014);
xnor U17348 (N_17348,N_16493,N_15802);
xnor U17349 (N_17349,N_15511,N_16492);
nor U17350 (N_17350,N_15720,N_16205);
and U17351 (N_17351,N_16440,N_15949);
or U17352 (N_17352,N_15237,N_15981);
xnor U17353 (N_17353,N_15862,N_15313);
nor U17354 (N_17354,N_16451,N_15762);
nand U17355 (N_17355,N_16167,N_16119);
nor U17356 (N_17356,N_15319,N_16336);
nor U17357 (N_17357,N_15516,N_16415);
nand U17358 (N_17358,N_15999,N_15280);
nand U17359 (N_17359,N_16397,N_16244);
nor U17360 (N_17360,N_16079,N_16258);
nand U17361 (N_17361,N_15423,N_15003);
nand U17362 (N_17362,N_15083,N_16061);
or U17363 (N_17363,N_15578,N_16290);
xor U17364 (N_17364,N_16015,N_16036);
or U17365 (N_17365,N_15364,N_15737);
and U17366 (N_17366,N_16006,N_16192);
and U17367 (N_17367,N_16290,N_15309);
and U17368 (N_17368,N_15781,N_16337);
or U17369 (N_17369,N_15784,N_16365);
or U17370 (N_17370,N_16194,N_15375);
nor U17371 (N_17371,N_16279,N_15352);
nand U17372 (N_17372,N_15253,N_15040);
nor U17373 (N_17373,N_16448,N_15404);
and U17374 (N_17374,N_16213,N_15388);
nand U17375 (N_17375,N_16313,N_15592);
nor U17376 (N_17376,N_15318,N_16296);
nand U17377 (N_17377,N_15365,N_15193);
or U17378 (N_17378,N_15732,N_16217);
xor U17379 (N_17379,N_15897,N_15495);
nor U17380 (N_17380,N_15792,N_15931);
xnor U17381 (N_17381,N_16238,N_15467);
or U17382 (N_17382,N_16141,N_16194);
or U17383 (N_17383,N_16373,N_16252);
or U17384 (N_17384,N_16074,N_16352);
nor U17385 (N_17385,N_15728,N_16225);
nand U17386 (N_17386,N_16311,N_16231);
nand U17387 (N_17387,N_16459,N_15334);
nor U17388 (N_17388,N_15793,N_15402);
xnor U17389 (N_17389,N_15476,N_15078);
or U17390 (N_17390,N_15225,N_15187);
and U17391 (N_17391,N_15901,N_15193);
or U17392 (N_17392,N_15950,N_15299);
nand U17393 (N_17393,N_15097,N_16157);
xor U17394 (N_17394,N_15754,N_15310);
nand U17395 (N_17395,N_15982,N_16362);
nor U17396 (N_17396,N_16159,N_16007);
xnor U17397 (N_17397,N_15935,N_15567);
nand U17398 (N_17398,N_15118,N_15049);
nor U17399 (N_17399,N_16221,N_15932);
xor U17400 (N_17400,N_15971,N_15602);
xnor U17401 (N_17401,N_16186,N_15396);
xnor U17402 (N_17402,N_15878,N_16282);
and U17403 (N_17403,N_15648,N_15571);
nor U17404 (N_17404,N_15466,N_15770);
or U17405 (N_17405,N_15225,N_15705);
nand U17406 (N_17406,N_16144,N_15676);
nand U17407 (N_17407,N_15920,N_15323);
nor U17408 (N_17408,N_15196,N_15166);
or U17409 (N_17409,N_15437,N_15670);
or U17410 (N_17410,N_16495,N_15919);
nor U17411 (N_17411,N_16080,N_16466);
nor U17412 (N_17412,N_16073,N_15092);
xnor U17413 (N_17413,N_15139,N_15849);
xnor U17414 (N_17414,N_15122,N_15024);
xor U17415 (N_17415,N_16427,N_15366);
or U17416 (N_17416,N_15369,N_15409);
nor U17417 (N_17417,N_15256,N_15919);
xor U17418 (N_17418,N_15684,N_15071);
and U17419 (N_17419,N_15886,N_15492);
or U17420 (N_17420,N_16149,N_15619);
nand U17421 (N_17421,N_15420,N_16028);
xor U17422 (N_17422,N_16421,N_16487);
or U17423 (N_17423,N_15691,N_15256);
nand U17424 (N_17424,N_16112,N_16097);
or U17425 (N_17425,N_15246,N_15564);
xor U17426 (N_17426,N_15122,N_15588);
nand U17427 (N_17427,N_16333,N_15278);
xnor U17428 (N_17428,N_16058,N_15080);
or U17429 (N_17429,N_16345,N_15855);
nand U17430 (N_17430,N_16066,N_16156);
and U17431 (N_17431,N_16217,N_15275);
nor U17432 (N_17432,N_16370,N_15349);
and U17433 (N_17433,N_16164,N_16280);
and U17434 (N_17434,N_15531,N_16113);
nand U17435 (N_17435,N_15401,N_15560);
nor U17436 (N_17436,N_15727,N_15439);
or U17437 (N_17437,N_15346,N_15370);
or U17438 (N_17438,N_15212,N_15342);
nor U17439 (N_17439,N_15351,N_15866);
or U17440 (N_17440,N_15557,N_16255);
xor U17441 (N_17441,N_15037,N_15910);
xnor U17442 (N_17442,N_16056,N_16278);
and U17443 (N_17443,N_15376,N_15145);
and U17444 (N_17444,N_16079,N_15307);
and U17445 (N_17445,N_16210,N_16005);
nor U17446 (N_17446,N_15138,N_15024);
nand U17447 (N_17447,N_16274,N_16104);
xnor U17448 (N_17448,N_15653,N_15827);
and U17449 (N_17449,N_15791,N_15814);
xor U17450 (N_17450,N_15279,N_15391);
or U17451 (N_17451,N_15719,N_15807);
nand U17452 (N_17452,N_16105,N_15237);
nand U17453 (N_17453,N_15118,N_15896);
xnor U17454 (N_17454,N_15359,N_16331);
xnor U17455 (N_17455,N_15567,N_16087);
or U17456 (N_17456,N_16234,N_15115);
or U17457 (N_17457,N_15440,N_15327);
or U17458 (N_17458,N_15744,N_15327);
nor U17459 (N_17459,N_15397,N_15062);
xnor U17460 (N_17460,N_15552,N_15073);
nor U17461 (N_17461,N_15071,N_16063);
and U17462 (N_17462,N_16137,N_16182);
nor U17463 (N_17463,N_15750,N_15192);
nand U17464 (N_17464,N_16359,N_16017);
xnor U17465 (N_17465,N_15959,N_15486);
xor U17466 (N_17466,N_16240,N_16145);
xnor U17467 (N_17467,N_15479,N_16230);
xor U17468 (N_17468,N_15549,N_16379);
nand U17469 (N_17469,N_15108,N_16038);
xnor U17470 (N_17470,N_16339,N_16041);
nand U17471 (N_17471,N_16020,N_16434);
nand U17472 (N_17472,N_15229,N_15551);
and U17473 (N_17473,N_15153,N_16018);
or U17474 (N_17474,N_15773,N_15132);
or U17475 (N_17475,N_16204,N_15914);
or U17476 (N_17476,N_16293,N_16057);
nor U17477 (N_17477,N_15860,N_15761);
or U17478 (N_17478,N_15882,N_16230);
nand U17479 (N_17479,N_15078,N_16288);
xnor U17480 (N_17480,N_15990,N_15529);
nand U17481 (N_17481,N_15414,N_16356);
or U17482 (N_17482,N_15917,N_16085);
xor U17483 (N_17483,N_15516,N_15645);
xor U17484 (N_17484,N_15518,N_15222);
or U17485 (N_17485,N_15809,N_15234);
xnor U17486 (N_17486,N_16395,N_15043);
nor U17487 (N_17487,N_15992,N_15559);
nor U17488 (N_17488,N_15660,N_16175);
nor U17489 (N_17489,N_15608,N_15173);
or U17490 (N_17490,N_15172,N_16027);
nor U17491 (N_17491,N_15674,N_15909);
and U17492 (N_17492,N_15962,N_16076);
nor U17493 (N_17493,N_15369,N_15395);
or U17494 (N_17494,N_16321,N_15093);
or U17495 (N_17495,N_15034,N_15001);
nor U17496 (N_17496,N_15697,N_15427);
xor U17497 (N_17497,N_16397,N_15853);
nor U17498 (N_17498,N_16473,N_15917);
nand U17499 (N_17499,N_15267,N_15779);
and U17500 (N_17500,N_15645,N_16266);
xnor U17501 (N_17501,N_15281,N_15792);
xor U17502 (N_17502,N_15917,N_15069);
or U17503 (N_17503,N_16093,N_15429);
nor U17504 (N_17504,N_15731,N_15333);
and U17505 (N_17505,N_15101,N_15307);
xor U17506 (N_17506,N_15268,N_16190);
or U17507 (N_17507,N_16362,N_15685);
and U17508 (N_17508,N_15121,N_16469);
nor U17509 (N_17509,N_15390,N_15594);
and U17510 (N_17510,N_15327,N_15296);
nor U17511 (N_17511,N_15918,N_15380);
or U17512 (N_17512,N_15098,N_16232);
xor U17513 (N_17513,N_16462,N_15334);
and U17514 (N_17514,N_15859,N_16161);
nor U17515 (N_17515,N_15710,N_16096);
nand U17516 (N_17516,N_16045,N_15304);
xnor U17517 (N_17517,N_15972,N_16277);
or U17518 (N_17518,N_16321,N_15553);
or U17519 (N_17519,N_15540,N_16335);
xor U17520 (N_17520,N_16010,N_15200);
nor U17521 (N_17521,N_15698,N_15323);
nand U17522 (N_17522,N_15057,N_16145);
or U17523 (N_17523,N_16411,N_15707);
and U17524 (N_17524,N_16339,N_15803);
nand U17525 (N_17525,N_15045,N_15666);
nand U17526 (N_17526,N_16006,N_16091);
nor U17527 (N_17527,N_16207,N_16112);
nand U17528 (N_17528,N_15755,N_15853);
xor U17529 (N_17529,N_15584,N_15429);
xor U17530 (N_17530,N_15251,N_16183);
nor U17531 (N_17531,N_16456,N_16068);
or U17532 (N_17532,N_15595,N_15629);
nand U17533 (N_17533,N_16256,N_15160);
or U17534 (N_17534,N_16425,N_15182);
xor U17535 (N_17535,N_15871,N_15039);
nor U17536 (N_17536,N_16307,N_16067);
nor U17537 (N_17537,N_16491,N_15426);
and U17538 (N_17538,N_16249,N_15473);
or U17539 (N_17539,N_16070,N_15496);
xor U17540 (N_17540,N_15157,N_16189);
and U17541 (N_17541,N_15411,N_16147);
or U17542 (N_17542,N_15948,N_15028);
or U17543 (N_17543,N_16446,N_15699);
and U17544 (N_17544,N_15658,N_16268);
nor U17545 (N_17545,N_15654,N_15518);
or U17546 (N_17546,N_15385,N_16013);
xnor U17547 (N_17547,N_16044,N_15189);
nor U17548 (N_17548,N_16289,N_16248);
nor U17549 (N_17549,N_15960,N_15028);
or U17550 (N_17550,N_16459,N_15179);
xor U17551 (N_17551,N_15782,N_15141);
xor U17552 (N_17552,N_16162,N_15471);
or U17553 (N_17553,N_15537,N_16411);
xor U17554 (N_17554,N_16013,N_15456);
and U17555 (N_17555,N_15808,N_16491);
nor U17556 (N_17556,N_15014,N_16193);
xnor U17557 (N_17557,N_15737,N_15397);
xor U17558 (N_17558,N_15727,N_15387);
and U17559 (N_17559,N_15820,N_15410);
or U17560 (N_17560,N_16036,N_16206);
and U17561 (N_17561,N_15606,N_15886);
nor U17562 (N_17562,N_16037,N_16170);
or U17563 (N_17563,N_15744,N_16418);
or U17564 (N_17564,N_15394,N_16003);
and U17565 (N_17565,N_15972,N_15950);
nand U17566 (N_17566,N_15353,N_15627);
and U17567 (N_17567,N_16445,N_16059);
or U17568 (N_17568,N_16343,N_16136);
nor U17569 (N_17569,N_15643,N_15625);
nor U17570 (N_17570,N_15166,N_15223);
and U17571 (N_17571,N_16331,N_16257);
and U17572 (N_17572,N_15887,N_15946);
nor U17573 (N_17573,N_15134,N_16270);
or U17574 (N_17574,N_16217,N_15368);
xnor U17575 (N_17575,N_16239,N_15796);
and U17576 (N_17576,N_15357,N_16473);
xnor U17577 (N_17577,N_15762,N_15816);
and U17578 (N_17578,N_15756,N_15495);
nand U17579 (N_17579,N_15938,N_15704);
xor U17580 (N_17580,N_15040,N_15802);
nand U17581 (N_17581,N_16005,N_15724);
nor U17582 (N_17582,N_15860,N_16490);
or U17583 (N_17583,N_16059,N_15705);
or U17584 (N_17584,N_15559,N_15642);
xor U17585 (N_17585,N_15921,N_15310);
nor U17586 (N_17586,N_15605,N_15583);
and U17587 (N_17587,N_15339,N_15349);
and U17588 (N_17588,N_16080,N_16054);
xor U17589 (N_17589,N_15570,N_16440);
nand U17590 (N_17590,N_15590,N_15388);
or U17591 (N_17591,N_16161,N_15202);
nor U17592 (N_17592,N_16083,N_16095);
nor U17593 (N_17593,N_16107,N_16209);
nor U17594 (N_17594,N_15817,N_15954);
or U17595 (N_17595,N_15407,N_15141);
nor U17596 (N_17596,N_16416,N_15996);
nand U17597 (N_17597,N_15222,N_16319);
or U17598 (N_17598,N_15280,N_16194);
nor U17599 (N_17599,N_16279,N_15673);
or U17600 (N_17600,N_15356,N_15441);
nor U17601 (N_17601,N_15358,N_15397);
or U17602 (N_17602,N_15438,N_15075);
xnor U17603 (N_17603,N_15735,N_15887);
xnor U17604 (N_17604,N_15090,N_16453);
nor U17605 (N_17605,N_15523,N_16307);
xor U17606 (N_17606,N_15953,N_16287);
nand U17607 (N_17607,N_15813,N_16027);
or U17608 (N_17608,N_15899,N_16487);
nor U17609 (N_17609,N_16256,N_16435);
nor U17610 (N_17610,N_16057,N_15273);
nor U17611 (N_17611,N_15485,N_15112);
or U17612 (N_17612,N_16126,N_15804);
nand U17613 (N_17613,N_16251,N_15195);
xnor U17614 (N_17614,N_16001,N_15293);
or U17615 (N_17615,N_15683,N_15361);
and U17616 (N_17616,N_15626,N_15294);
or U17617 (N_17617,N_16001,N_15577);
nand U17618 (N_17618,N_16441,N_15983);
or U17619 (N_17619,N_15654,N_16264);
and U17620 (N_17620,N_15589,N_15799);
nor U17621 (N_17621,N_15286,N_16084);
or U17622 (N_17622,N_16363,N_16181);
nand U17623 (N_17623,N_15213,N_15685);
and U17624 (N_17624,N_15598,N_16315);
or U17625 (N_17625,N_15713,N_16314);
or U17626 (N_17626,N_16491,N_15931);
nor U17627 (N_17627,N_15314,N_16283);
xor U17628 (N_17628,N_15649,N_15868);
or U17629 (N_17629,N_15996,N_15044);
nor U17630 (N_17630,N_15730,N_15834);
nor U17631 (N_17631,N_15931,N_15197);
or U17632 (N_17632,N_15967,N_16365);
xor U17633 (N_17633,N_15347,N_15168);
or U17634 (N_17634,N_16308,N_15981);
and U17635 (N_17635,N_15549,N_15149);
nor U17636 (N_17636,N_16098,N_15883);
and U17637 (N_17637,N_16119,N_16158);
and U17638 (N_17638,N_16403,N_16399);
or U17639 (N_17639,N_16385,N_16319);
and U17640 (N_17640,N_16429,N_15482);
or U17641 (N_17641,N_15720,N_15078);
nand U17642 (N_17642,N_15590,N_15612);
nor U17643 (N_17643,N_15286,N_15666);
and U17644 (N_17644,N_16243,N_15712);
nor U17645 (N_17645,N_15955,N_15250);
and U17646 (N_17646,N_15016,N_15514);
nand U17647 (N_17647,N_15123,N_16033);
xnor U17648 (N_17648,N_15182,N_15420);
xor U17649 (N_17649,N_15698,N_15724);
and U17650 (N_17650,N_15272,N_15810);
and U17651 (N_17651,N_16431,N_15219);
nand U17652 (N_17652,N_15619,N_15185);
or U17653 (N_17653,N_15851,N_15420);
xnor U17654 (N_17654,N_16427,N_16041);
nand U17655 (N_17655,N_15356,N_16104);
or U17656 (N_17656,N_15416,N_16006);
and U17657 (N_17657,N_15665,N_16066);
xor U17658 (N_17658,N_15476,N_15262);
nand U17659 (N_17659,N_16402,N_16293);
or U17660 (N_17660,N_15270,N_15946);
nand U17661 (N_17661,N_15767,N_15337);
xor U17662 (N_17662,N_15434,N_16077);
nand U17663 (N_17663,N_15449,N_16326);
and U17664 (N_17664,N_16479,N_15632);
nand U17665 (N_17665,N_15903,N_16331);
nor U17666 (N_17666,N_15526,N_16183);
nor U17667 (N_17667,N_15304,N_15762);
xnor U17668 (N_17668,N_15811,N_15265);
nand U17669 (N_17669,N_15078,N_15376);
nand U17670 (N_17670,N_15691,N_15727);
nor U17671 (N_17671,N_16014,N_16139);
nand U17672 (N_17672,N_15397,N_15661);
or U17673 (N_17673,N_16296,N_16045);
or U17674 (N_17674,N_16457,N_15646);
nand U17675 (N_17675,N_15684,N_15573);
and U17676 (N_17676,N_15774,N_16028);
or U17677 (N_17677,N_15635,N_15349);
or U17678 (N_17678,N_15594,N_15162);
or U17679 (N_17679,N_15996,N_15132);
and U17680 (N_17680,N_16375,N_15330);
and U17681 (N_17681,N_16426,N_16250);
xnor U17682 (N_17682,N_15621,N_16368);
nand U17683 (N_17683,N_15612,N_15103);
nand U17684 (N_17684,N_16206,N_15738);
nor U17685 (N_17685,N_16225,N_16412);
or U17686 (N_17686,N_16496,N_15371);
nand U17687 (N_17687,N_15615,N_15533);
nand U17688 (N_17688,N_15103,N_15016);
nand U17689 (N_17689,N_15110,N_15025);
or U17690 (N_17690,N_16471,N_15446);
xnor U17691 (N_17691,N_15526,N_15116);
and U17692 (N_17692,N_15952,N_15142);
and U17693 (N_17693,N_16161,N_15613);
nand U17694 (N_17694,N_16287,N_16384);
or U17695 (N_17695,N_15872,N_15484);
and U17696 (N_17696,N_16266,N_16098);
xnor U17697 (N_17697,N_15548,N_16242);
and U17698 (N_17698,N_16313,N_16218);
xnor U17699 (N_17699,N_15091,N_16022);
xnor U17700 (N_17700,N_15225,N_15252);
nand U17701 (N_17701,N_15202,N_15032);
xnor U17702 (N_17702,N_15357,N_15490);
or U17703 (N_17703,N_16244,N_15092);
or U17704 (N_17704,N_16058,N_15381);
nand U17705 (N_17705,N_15271,N_16410);
xor U17706 (N_17706,N_15499,N_15928);
or U17707 (N_17707,N_15490,N_15879);
nand U17708 (N_17708,N_16499,N_15549);
or U17709 (N_17709,N_15643,N_15960);
or U17710 (N_17710,N_16491,N_15839);
nand U17711 (N_17711,N_16134,N_15137);
nor U17712 (N_17712,N_15401,N_16300);
nand U17713 (N_17713,N_15565,N_16082);
nand U17714 (N_17714,N_15647,N_15842);
or U17715 (N_17715,N_16381,N_15968);
nor U17716 (N_17716,N_15849,N_15260);
xor U17717 (N_17717,N_15144,N_16453);
and U17718 (N_17718,N_15081,N_15844);
xor U17719 (N_17719,N_15129,N_16296);
xnor U17720 (N_17720,N_15246,N_15806);
nor U17721 (N_17721,N_15670,N_15886);
xnor U17722 (N_17722,N_16047,N_15141);
or U17723 (N_17723,N_16203,N_15143);
xnor U17724 (N_17724,N_15596,N_16231);
xor U17725 (N_17725,N_15515,N_16100);
or U17726 (N_17726,N_15299,N_15592);
or U17727 (N_17727,N_15654,N_16179);
and U17728 (N_17728,N_15126,N_16036);
xnor U17729 (N_17729,N_15545,N_16158);
nand U17730 (N_17730,N_16203,N_15434);
nand U17731 (N_17731,N_15111,N_16394);
or U17732 (N_17732,N_15353,N_15571);
xor U17733 (N_17733,N_16229,N_15727);
or U17734 (N_17734,N_15706,N_16385);
nand U17735 (N_17735,N_15048,N_15780);
nor U17736 (N_17736,N_15798,N_15516);
nor U17737 (N_17737,N_15797,N_15358);
or U17738 (N_17738,N_15863,N_15267);
or U17739 (N_17739,N_15985,N_15461);
or U17740 (N_17740,N_15838,N_16066);
xor U17741 (N_17741,N_15461,N_15328);
nand U17742 (N_17742,N_15084,N_16010);
xnor U17743 (N_17743,N_15692,N_16273);
nor U17744 (N_17744,N_15673,N_16039);
nor U17745 (N_17745,N_15814,N_16317);
nor U17746 (N_17746,N_16175,N_16034);
or U17747 (N_17747,N_16447,N_16390);
nand U17748 (N_17748,N_16026,N_15045);
nor U17749 (N_17749,N_15267,N_15448);
and U17750 (N_17750,N_16435,N_15597);
nor U17751 (N_17751,N_16113,N_15888);
nand U17752 (N_17752,N_16117,N_15884);
and U17753 (N_17753,N_15865,N_16264);
or U17754 (N_17754,N_15357,N_16389);
and U17755 (N_17755,N_16407,N_15868);
and U17756 (N_17756,N_16403,N_15436);
or U17757 (N_17757,N_16287,N_15733);
nand U17758 (N_17758,N_15172,N_16403);
or U17759 (N_17759,N_15483,N_15922);
or U17760 (N_17760,N_15022,N_15128);
xnor U17761 (N_17761,N_15312,N_16269);
nand U17762 (N_17762,N_16311,N_15739);
nand U17763 (N_17763,N_15109,N_15398);
or U17764 (N_17764,N_15038,N_16494);
nor U17765 (N_17765,N_15739,N_15478);
nand U17766 (N_17766,N_15977,N_15542);
xnor U17767 (N_17767,N_15664,N_15892);
xnor U17768 (N_17768,N_15748,N_15572);
or U17769 (N_17769,N_15003,N_15549);
or U17770 (N_17770,N_16301,N_15065);
xnor U17771 (N_17771,N_15608,N_15770);
xor U17772 (N_17772,N_15488,N_15484);
nor U17773 (N_17773,N_15069,N_15809);
nor U17774 (N_17774,N_15632,N_15511);
nor U17775 (N_17775,N_15205,N_15230);
nor U17776 (N_17776,N_15682,N_15303);
nand U17777 (N_17777,N_15857,N_16069);
and U17778 (N_17778,N_15577,N_15688);
and U17779 (N_17779,N_15811,N_15686);
nor U17780 (N_17780,N_16244,N_16231);
nor U17781 (N_17781,N_16012,N_16161);
and U17782 (N_17782,N_15139,N_16141);
nor U17783 (N_17783,N_15448,N_15067);
nand U17784 (N_17784,N_16451,N_15667);
or U17785 (N_17785,N_15945,N_15535);
or U17786 (N_17786,N_16352,N_15770);
or U17787 (N_17787,N_16228,N_16022);
or U17788 (N_17788,N_15130,N_15819);
nor U17789 (N_17789,N_15321,N_16375);
or U17790 (N_17790,N_15608,N_16239);
and U17791 (N_17791,N_16050,N_15608);
or U17792 (N_17792,N_15798,N_16141);
or U17793 (N_17793,N_15187,N_16177);
xor U17794 (N_17794,N_15495,N_16146);
nand U17795 (N_17795,N_15629,N_16409);
and U17796 (N_17796,N_15093,N_15968);
and U17797 (N_17797,N_15284,N_15076);
or U17798 (N_17798,N_15749,N_16322);
and U17799 (N_17799,N_15502,N_15642);
nand U17800 (N_17800,N_15245,N_15446);
and U17801 (N_17801,N_15968,N_15094);
nand U17802 (N_17802,N_16413,N_15283);
xnor U17803 (N_17803,N_15752,N_16071);
nand U17804 (N_17804,N_15608,N_15808);
or U17805 (N_17805,N_15904,N_16117);
nor U17806 (N_17806,N_15874,N_15484);
or U17807 (N_17807,N_16172,N_15569);
nand U17808 (N_17808,N_15933,N_15910);
and U17809 (N_17809,N_15569,N_15303);
and U17810 (N_17810,N_15449,N_16436);
nor U17811 (N_17811,N_15443,N_15565);
nor U17812 (N_17812,N_15263,N_15760);
and U17813 (N_17813,N_15963,N_15876);
nand U17814 (N_17814,N_15831,N_16182);
nor U17815 (N_17815,N_15951,N_16215);
nor U17816 (N_17816,N_15929,N_16382);
nor U17817 (N_17817,N_16068,N_15192);
or U17818 (N_17818,N_15979,N_16385);
nor U17819 (N_17819,N_15989,N_16210);
nor U17820 (N_17820,N_15945,N_16116);
xor U17821 (N_17821,N_16473,N_15680);
nor U17822 (N_17822,N_16411,N_15297);
or U17823 (N_17823,N_15152,N_16216);
nor U17824 (N_17824,N_15671,N_15819);
xnor U17825 (N_17825,N_16307,N_16469);
nand U17826 (N_17826,N_15407,N_15894);
nor U17827 (N_17827,N_15225,N_15375);
and U17828 (N_17828,N_15877,N_15513);
and U17829 (N_17829,N_15164,N_15138);
nor U17830 (N_17830,N_16083,N_15895);
and U17831 (N_17831,N_15687,N_15995);
nand U17832 (N_17832,N_16015,N_15010);
nor U17833 (N_17833,N_15135,N_15092);
xor U17834 (N_17834,N_16031,N_15532);
nand U17835 (N_17835,N_16005,N_15268);
xnor U17836 (N_17836,N_15065,N_16380);
nand U17837 (N_17837,N_15091,N_15427);
xnor U17838 (N_17838,N_15842,N_16142);
nor U17839 (N_17839,N_15963,N_16262);
xnor U17840 (N_17840,N_15773,N_16086);
nand U17841 (N_17841,N_15063,N_16411);
nand U17842 (N_17842,N_15145,N_15312);
nand U17843 (N_17843,N_15138,N_16142);
and U17844 (N_17844,N_15564,N_15183);
and U17845 (N_17845,N_15604,N_16369);
xnor U17846 (N_17846,N_16448,N_15653);
nand U17847 (N_17847,N_16300,N_15029);
xnor U17848 (N_17848,N_16215,N_15281);
nor U17849 (N_17849,N_16342,N_16084);
and U17850 (N_17850,N_15303,N_15691);
and U17851 (N_17851,N_15134,N_16328);
and U17852 (N_17852,N_15730,N_15581);
or U17853 (N_17853,N_15080,N_15092);
xor U17854 (N_17854,N_15165,N_15350);
nand U17855 (N_17855,N_15679,N_16426);
xnor U17856 (N_17856,N_15478,N_15651);
and U17857 (N_17857,N_15433,N_15381);
and U17858 (N_17858,N_16106,N_15295);
or U17859 (N_17859,N_15316,N_15271);
xor U17860 (N_17860,N_15918,N_15549);
nand U17861 (N_17861,N_15598,N_16360);
nand U17862 (N_17862,N_15498,N_15730);
nand U17863 (N_17863,N_16311,N_15665);
xor U17864 (N_17864,N_15023,N_15321);
and U17865 (N_17865,N_15105,N_15904);
and U17866 (N_17866,N_15581,N_16255);
and U17867 (N_17867,N_15807,N_15091);
and U17868 (N_17868,N_15715,N_15061);
nand U17869 (N_17869,N_16019,N_15250);
xor U17870 (N_17870,N_15091,N_15927);
nand U17871 (N_17871,N_16229,N_15968);
and U17872 (N_17872,N_15953,N_16102);
nor U17873 (N_17873,N_16106,N_15760);
nor U17874 (N_17874,N_15865,N_15050);
and U17875 (N_17875,N_15244,N_16018);
or U17876 (N_17876,N_15416,N_15385);
nand U17877 (N_17877,N_15627,N_15216);
and U17878 (N_17878,N_15600,N_15980);
nand U17879 (N_17879,N_15589,N_15190);
nor U17880 (N_17880,N_15599,N_15512);
nor U17881 (N_17881,N_15188,N_15624);
nand U17882 (N_17882,N_15379,N_15608);
or U17883 (N_17883,N_15399,N_16420);
xnor U17884 (N_17884,N_15842,N_15280);
xor U17885 (N_17885,N_15427,N_16206);
and U17886 (N_17886,N_15058,N_15540);
nand U17887 (N_17887,N_16235,N_15374);
nor U17888 (N_17888,N_16272,N_15103);
nor U17889 (N_17889,N_15382,N_16327);
and U17890 (N_17890,N_15730,N_15408);
nand U17891 (N_17891,N_15141,N_15000);
nand U17892 (N_17892,N_15789,N_15433);
nor U17893 (N_17893,N_15740,N_15264);
or U17894 (N_17894,N_15123,N_16403);
or U17895 (N_17895,N_15966,N_16179);
nand U17896 (N_17896,N_16391,N_15298);
nor U17897 (N_17897,N_15782,N_15891);
or U17898 (N_17898,N_16482,N_15981);
and U17899 (N_17899,N_15162,N_15109);
or U17900 (N_17900,N_15015,N_16247);
nor U17901 (N_17901,N_16011,N_15254);
nor U17902 (N_17902,N_16028,N_15394);
and U17903 (N_17903,N_15542,N_16301);
nor U17904 (N_17904,N_15137,N_15058);
nand U17905 (N_17905,N_15249,N_15445);
nor U17906 (N_17906,N_16378,N_15701);
nand U17907 (N_17907,N_15629,N_15687);
and U17908 (N_17908,N_15279,N_16160);
xor U17909 (N_17909,N_15376,N_16064);
nand U17910 (N_17910,N_15483,N_16154);
xnor U17911 (N_17911,N_16097,N_15878);
and U17912 (N_17912,N_15832,N_16255);
nand U17913 (N_17913,N_15185,N_16467);
nor U17914 (N_17914,N_16164,N_15032);
nand U17915 (N_17915,N_15031,N_15094);
and U17916 (N_17916,N_15958,N_16317);
xor U17917 (N_17917,N_15473,N_15191);
or U17918 (N_17918,N_16429,N_16433);
xnor U17919 (N_17919,N_15245,N_15232);
nand U17920 (N_17920,N_15745,N_16290);
nor U17921 (N_17921,N_16092,N_15607);
or U17922 (N_17922,N_15664,N_15235);
nand U17923 (N_17923,N_15806,N_16071);
and U17924 (N_17924,N_16262,N_15210);
or U17925 (N_17925,N_15492,N_16353);
and U17926 (N_17926,N_15174,N_16142);
and U17927 (N_17927,N_15260,N_15295);
or U17928 (N_17928,N_16298,N_16355);
nor U17929 (N_17929,N_15774,N_15183);
or U17930 (N_17930,N_16323,N_16456);
nand U17931 (N_17931,N_16201,N_16331);
or U17932 (N_17932,N_16379,N_15347);
xnor U17933 (N_17933,N_15403,N_15613);
nand U17934 (N_17934,N_15908,N_15818);
and U17935 (N_17935,N_15540,N_16004);
xor U17936 (N_17936,N_15350,N_15412);
nor U17937 (N_17937,N_15777,N_15789);
nand U17938 (N_17938,N_15484,N_15755);
nor U17939 (N_17939,N_15831,N_15651);
or U17940 (N_17940,N_16181,N_15341);
or U17941 (N_17941,N_16433,N_15113);
nand U17942 (N_17942,N_15033,N_16190);
and U17943 (N_17943,N_15416,N_15351);
nor U17944 (N_17944,N_15434,N_16263);
nor U17945 (N_17945,N_15726,N_16312);
nand U17946 (N_17946,N_15727,N_15115);
nor U17947 (N_17947,N_15352,N_15171);
or U17948 (N_17948,N_15596,N_15112);
and U17949 (N_17949,N_15252,N_15620);
xnor U17950 (N_17950,N_15562,N_15771);
and U17951 (N_17951,N_15354,N_15933);
and U17952 (N_17952,N_15233,N_15963);
and U17953 (N_17953,N_15326,N_16155);
nor U17954 (N_17954,N_16107,N_15746);
xnor U17955 (N_17955,N_15094,N_15577);
xor U17956 (N_17956,N_15724,N_15581);
nand U17957 (N_17957,N_16151,N_15820);
nand U17958 (N_17958,N_16199,N_15737);
nand U17959 (N_17959,N_16364,N_15267);
xnor U17960 (N_17960,N_15570,N_16493);
or U17961 (N_17961,N_16330,N_16022);
and U17962 (N_17962,N_15328,N_15520);
or U17963 (N_17963,N_15721,N_15889);
or U17964 (N_17964,N_15151,N_15673);
nor U17965 (N_17965,N_15593,N_15004);
or U17966 (N_17966,N_15026,N_15563);
nor U17967 (N_17967,N_16059,N_16000);
nand U17968 (N_17968,N_15747,N_15983);
xor U17969 (N_17969,N_15264,N_15473);
xnor U17970 (N_17970,N_15078,N_16175);
or U17971 (N_17971,N_15979,N_16441);
nand U17972 (N_17972,N_15900,N_15165);
nand U17973 (N_17973,N_16090,N_15390);
and U17974 (N_17974,N_15551,N_15564);
nand U17975 (N_17975,N_15569,N_15993);
or U17976 (N_17976,N_15074,N_16319);
nor U17977 (N_17977,N_16054,N_15668);
nand U17978 (N_17978,N_15690,N_16318);
and U17979 (N_17979,N_16267,N_15515);
or U17980 (N_17980,N_15450,N_16066);
or U17981 (N_17981,N_15457,N_15937);
or U17982 (N_17982,N_16173,N_15258);
nor U17983 (N_17983,N_16308,N_15067);
nor U17984 (N_17984,N_15113,N_16395);
nand U17985 (N_17985,N_15923,N_15150);
xor U17986 (N_17986,N_15125,N_15755);
nor U17987 (N_17987,N_16252,N_15626);
nand U17988 (N_17988,N_15117,N_15183);
nor U17989 (N_17989,N_16225,N_16058);
xnor U17990 (N_17990,N_15572,N_15220);
or U17991 (N_17991,N_15796,N_16381);
or U17992 (N_17992,N_15621,N_15453);
nor U17993 (N_17993,N_15060,N_15847);
xnor U17994 (N_17994,N_15630,N_15858);
and U17995 (N_17995,N_15900,N_16055);
and U17996 (N_17996,N_15062,N_15888);
nor U17997 (N_17997,N_15809,N_16401);
nand U17998 (N_17998,N_16061,N_16345);
nor U17999 (N_17999,N_16194,N_15281);
or U18000 (N_18000,N_17826,N_17361);
nor U18001 (N_18001,N_17027,N_17706);
and U18002 (N_18002,N_17930,N_16767);
and U18003 (N_18003,N_16563,N_17092);
nor U18004 (N_18004,N_17634,N_17152);
xor U18005 (N_18005,N_17228,N_17266);
and U18006 (N_18006,N_17920,N_17453);
xor U18007 (N_18007,N_17053,N_16517);
or U18008 (N_18008,N_17849,N_17049);
nor U18009 (N_18009,N_16590,N_16813);
or U18010 (N_18010,N_16540,N_17060);
or U18011 (N_18011,N_17752,N_17686);
or U18012 (N_18012,N_17010,N_16627);
nand U18013 (N_18013,N_16998,N_17946);
nor U18014 (N_18014,N_17513,N_17760);
nor U18015 (N_18015,N_17698,N_16888);
and U18016 (N_18016,N_17312,N_17810);
or U18017 (N_18017,N_17277,N_17133);
or U18018 (N_18018,N_17588,N_17790);
xor U18019 (N_18019,N_17523,N_17876);
nor U18020 (N_18020,N_16705,N_16957);
nand U18021 (N_18021,N_16656,N_16737);
or U18022 (N_18022,N_17116,N_17894);
nand U18023 (N_18023,N_17583,N_16732);
and U18024 (N_18024,N_17624,N_16869);
nand U18025 (N_18025,N_17573,N_17683);
xnor U18026 (N_18026,N_17633,N_17879);
and U18027 (N_18027,N_16582,N_17140);
and U18028 (N_18028,N_17471,N_17132);
xor U18029 (N_18029,N_17081,N_17380);
or U18030 (N_18030,N_17660,N_16778);
nor U18031 (N_18031,N_17337,N_16719);
xor U18032 (N_18032,N_17552,N_17891);
and U18033 (N_18033,N_16603,N_16789);
and U18034 (N_18034,N_17699,N_17550);
nand U18035 (N_18035,N_16626,N_16677);
xnor U18036 (N_18036,N_17271,N_16753);
nand U18037 (N_18037,N_16585,N_16931);
xor U18038 (N_18038,N_16623,N_17602);
nor U18039 (N_18039,N_17303,N_17368);
or U18040 (N_18040,N_16586,N_16845);
or U18041 (N_18041,N_16722,N_17911);
or U18042 (N_18042,N_17733,N_16924);
nor U18043 (N_18043,N_17632,N_16604);
nand U18044 (N_18044,N_16768,N_17926);
nor U18045 (N_18045,N_17396,N_16991);
nand U18046 (N_18046,N_16619,N_17286);
nor U18047 (N_18047,N_17122,N_16681);
or U18048 (N_18048,N_17666,N_17405);
nand U18049 (N_18049,N_16632,N_17769);
or U18050 (N_18050,N_17107,N_16673);
and U18051 (N_18051,N_16606,N_16579);
nor U18052 (N_18052,N_16727,N_17074);
xnor U18053 (N_18053,N_16791,N_17897);
nand U18054 (N_18054,N_17837,N_17594);
and U18055 (N_18055,N_17054,N_17886);
and U18056 (N_18056,N_16564,N_17157);
xnor U18057 (N_18057,N_17783,N_17064);
nor U18058 (N_18058,N_17969,N_17267);
nand U18059 (N_18059,N_17007,N_17576);
xnor U18060 (N_18060,N_16565,N_17324);
and U18061 (N_18061,N_17229,N_16983);
nand U18062 (N_18062,N_17527,N_17447);
nand U18063 (N_18063,N_17600,N_16600);
nor U18064 (N_18064,N_17689,N_17482);
nand U18065 (N_18065,N_16794,N_17457);
nor U18066 (N_18066,N_16618,N_17679);
nand U18067 (N_18067,N_17195,N_17118);
or U18068 (N_18068,N_17967,N_17547);
or U18069 (N_18069,N_16730,N_17807);
nor U18070 (N_18070,N_17412,N_16697);
nor U18071 (N_18071,N_17456,N_17024);
or U18072 (N_18072,N_17842,N_17665);
or U18073 (N_18073,N_16827,N_17892);
nand U18074 (N_18074,N_16850,N_17250);
nand U18075 (N_18075,N_17510,N_16928);
or U18076 (N_18076,N_16717,N_17598);
nor U18077 (N_18077,N_17794,N_17188);
xor U18078 (N_18078,N_17287,N_17243);
or U18079 (N_18079,N_17778,N_16916);
xnor U18080 (N_18080,N_16877,N_16823);
and U18081 (N_18081,N_17993,N_16855);
nor U18082 (N_18082,N_16833,N_17461);
xnor U18083 (N_18083,N_16873,N_17506);
and U18084 (N_18084,N_17675,N_17565);
or U18085 (N_18085,N_17785,N_17659);
or U18086 (N_18086,N_17497,N_17451);
and U18087 (N_18087,N_17454,N_16708);
xnor U18088 (N_18088,N_17311,N_16525);
xor U18089 (N_18089,N_16500,N_16748);
xor U18090 (N_18090,N_17742,N_16926);
nand U18091 (N_18091,N_17493,N_16639);
and U18092 (N_18092,N_16508,N_17559);
or U18093 (N_18093,N_17292,N_16786);
nand U18094 (N_18094,N_17623,N_17854);
xor U18095 (N_18095,N_16574,N_16883);
or U18096 (N_18096,N_17804,N_17525);
xnor U18097 (N_18097,N_17015,N_17128);
or U18098 (N_18098,N_17558,N_16758);
and U18099 (N_18099,N_17159,N_17431);
and U18100 (N_18100,N_17596,N_17065);
xnor U18101 (N_18101,N_16524,N_17342);
xor U18102 (N_18102,N_16890,N_17863);
and U18103 (N_18103,N_17982,N_17618);
nor U18104 (N_18104,N_17339,N_17922);
xor U18105 (N_18105,N_16909,N_17418);
nor U18106 (N_18106,N_17495,N_17714);
and U18107 (N_18107,N_16554,N_17925);
nand U18108 (N_18108,N_16974,N_17028);
xor U18109 (N_18109,N_16710,N_17035);
xnor U18110 (N_18110,N_16901,N_17958);
nand U18111 (N_18111,N_17984,N_17866);
xnor U18112 (N_18112,N_17590,N_16615);
or U18113 (N_18113,N_16930,N_17115);
nor U18114 (N_18114,N_17415,N_17038);
or U18115 (N_18115,N_17582,N_17455);
nor U18116 (N_18116,N_17387,N_16513);
xor U18117 (N_18117,N_17375,N_16964);
or U18118 (N_18118,N_16537,N_17649);
nor U18119 (N_18119,N_17927,N_16605);
nor U18120 (N_18120,N_16734,N_16746);
nor U18121 (N_18121,N_17275,N_17847);
and U18122 (N_18122,N_16569,N_16912);
and U18123 (N_18123,N_16642,N_16811);
xor U18124 (N_18124,N_17389,N_17123);
or U18125 (N_18125,N_16687,N_16820);
nand U18126 (N_18126,N_17094,N_16599);
or U18127 (N_18127,N_16933,N_17018);
nor U18128 (N_18128,N_17073,N_17715);
and U18129 (N_18129,N_16665,N_16976);
xor U18130 (N_18130,N_16509,N_17124);
nor U18131 (N_18131,N_16715,N_17829);
nor U18132 (N_18132,N_17856,N_17522);
nand U18133 (N_18133,N_16799,N_17254);
nor U18134 (N_18134,N_17792,N_17947);
nand U18135 (N_18135,N_17202,N_17592);
and U18136 (N_18136,N_17452,N_16830);
nor U18137 (N_18137,N_16894,N_17884);
and U18138 (N_18138,N_17986,N_17163);
xor U18139 (N_18139,N_16514,N_17627);
nand U18140 (N_18140,N_16714,N_16663);
or U18141 (N_18141,N_17750,N_17006);
and U18142 (N_18142,N_17002,N_17260);
xnor U18143 (N_18143,N_17043,N_17664);
nor U18144 (N_18144,N_16607,N_17083);
or U18145 (N_18145,N_17386,N_17318);
nand U18146 (N_18146,N_17687,N_17764);
nand U18147 (N_18147,N_16962,N_17612);
nor U18148 (N_18148,N_17647,N_17621);
or U18149 (N_18149,N_16515,N_17485);
and U18150 (N_18150,N_17727,N_17850);
and U18151 (N_18151,N_17668,N_16592);
and U18152 (N_18152,N_17808,N_16752);
nand U18153 (N_18153,N_17799,N_17104);
nand U18154 (N_18154,N_16690,N_17924);
nor U18155 (N_18155,N_16674,N_16906);
or U18156 (N_18156,N_17187,N_16760);
or U18157 (N_18157,N_16625,N_17688);
and U18158 (N_18158,N_17265,N_16939);
xnor U18159 (N_18159,N_16675,N_17761);
nor U18160 (N_18160,N_17992,N_17902);
or U18161 (N_18161,N_17258,N_16516);
and U18162 (N_18162,N_16634,N_16651);
or U18163 (N_18163,N_17816,N_17881);
nand U18164 (N_18164,N_17821,N_17432);
nor U18165 (N_18165,N_17516,N_17997);
or U18166 (N_18166,N_17721,N_16611);
nand U18167 (N_18167,N_17131,N_17540);
nand U18168 (N_18168,N_16836,N_17678);
xnor U18169 (N_18169,N_16751,N_16694);
nand U18170 (N_18170,N_16602,N_17971);
xor U18171 (N_18171,N_16958,N_16633);
xnor U18172 (N_18172,N_16560,N_17164);
xor U18173 (N_18173,N_16792,N_16724);
nor U18174 (N_18174,N_17383,N_16971);
nand U18175 (N_18175,N_17803,N_17204);
and U18176 (N_18176,N_17154,N_17753);
nand U18177 (N_18177,N_17746,N_17486);
nor U18178 (N_18178,N_17488,N_17839);
nor U18179 (N_18179,N_17631,N_16977);
or U18180 (N_18180,N_16763,N_16796);
xor U18181 (N_18181,N_17800,N_17641);
xnor U18182 (N_18182,N_16887,N_16650);
xnor U18183 (N_18183,N_17994,N_17817);
or U18184 (N_18184,N_17402,N_17409);
and U18185 (N_18185,N_17307,N_17620);
and U18186 (N_18186,N_16731,N_16821);
and U18187 (N_18187,N_17448,N_16631);
xor U18188 (N_18188,N_16718,N_17653);
xnor U18189 (N_18189,N_16812,N_17041);
xnor U18190 (N_18190,N_17009,N_16943);
and U18191 (N_18191,N_16709,N_16969);
nor U18192 (N_18192,N_17954,N_17741);
nand U18193 (N_18193,N_17102,N_16859);
and U18194 (N_18194,N_17904,N_17150);
and U18195 (N_18195,N_17419,N_17210);
nand U18196 (N_18196,N_16555,N_16698);
nand U18197 (N_18197,N_16583,N_17212);
and U18198 (N_18198,N_17692,N_17906);
or U18199 (N_18199,N_16503,N_16782);
and U18200 (N_18200,N_16502,N_17662);
nor U18201 (N_18201,N_16616,N_17185);
xnor U18202 (N_18202,N_17529,N_17572);
and U18203 (N_18203,N_17942,N_17232);
nand U18204 (N_18204,N_17321,N_17512);
nor U18205 (N_18205,N_17851,N_17609);
nand U18206 (N_18206,N_17438,N_17147);
or U18207 (N_18207,N_17076,N_17796);
or U18208 (N_18208,N_16646,N_16995);
xor U18209 (N_18209,N_17599,N_17352);
xnor U18210 (N_18210,N_17999,N_17606);
and U18211 (N_18211,N_16534,N_17445);
and U18212 (N_18212,N_17446,N_17069);
and U18213 (N_18213,N_17171,N_17155);
and U18214 (N_18214,N_16686,N_17240);
xnor U18215 (N_18215,N_17754,N_16580);
and U18216 (N_18216,N_17979,N_16562);
xor U18217 (N_18217,N_17033,N_17913);
nor U18218 (N_18218,N_16578,N_17005);
nand U18219 (N_18219,N_17838,N_17084);
nand U18220 (N_18220,N_16679,N_17531);
nor U18221 (N_18221,N_16941,N_16835);
and U18222 (N_18222,N_16934,N_17661);
and U18223 (N_18223,N_17444,N_17098);
nand U18224 (N_18224,N_16571,N_17639);
or U18225 (N_18225,N_17003,N_17196);
nand U18226 (N_18226,N_17019,N_17864);
and U18227 (N_18227,N_17561,N_17974);
nor U18228 (N_18228,N_17344,N_16601);
nor U18229 (N_18229,N_17422,N_17518);
xnor U18230 (N_18230,N_16527,N_16706);
nor U18231 (N_18231,N_17392,N_16842);
nand U18232 (N_18232,N_16536,N_17044);
or U18233 (N_18233,N_17694,N_17136);
nor U18234 (N_18234,N_17909,N_16922);
nand U18235 (N_18235,N_17358,N_16824);
or U18236 (N_18236,N_16925,N_16664);
or U18237 (N_18237,N_17809,N_17492);
nor U18238 (N_18238,N_17834,N_17549);
or U18239 (N_18239,N_17487,N_16567);
and U18240 (N_18240,N_17376,N_17981);
nor U18241 (N_18241,N_17371,N_17075);
and U18242 (N_18242,N_17093,N_17595);
and U18243 (N_18243,N_16817,N_17873);
nand U18244 (N_18244,N_17987,N_17734);
nand U18245 (N_18245,N_17551,N_16756);
nand U18246 (N_18246,N_17225,N_17840);
and U18247 (N_18247,N_17333,N_16692);
nor U18248 (N_18248,N_16549,N_17724);
nand U18249 (N_18249,N_16938,N_16612);
or U18250 (N_18250,N_17782,N_16541);
and U18251 (N_18251,N_16702,N_16902);
nor U18252 (N_18252,N_17468,N_17763);
nor U18253 (N_18253,N_17354,N_17604);
xor U18254 (N_18254,N_17231,N_17918);
nand U18255 (N_18255,N_17667,N_16860);
and U18256 (N_18256,N_17360,N_16595);
xor U18257 (N_18257,N_17233,N_17110);
and U18258 (N_18258,N_16653,N_16861);
nand U18259 (N_18259,N_17201,N_17190);
or U18260 (N_18260,N_17774,N_17941);
nand U18261 (N_18261,N_17732,N_17546);
nor U18262 (N_18262,N_17080,N_17217);
xnor U18263 (N_18263,N_16691,N_16846);
and U18264 (N_18264,N_17117,N_16935);
xor U18265 (N_18265,N_17428,N_16621);
or U18266 (N_18266,N_17670,N_17938);
or U18267 (N_18267,N_16893,N_17478);
nand U18268 (N_18268,N_17014,N_17086);
nand U18269 (N_18269,N_17385,N_17087);
or U18270 (N_18270,N_16764,N_16669);
nand U18271 (N_18271,N_17079,N_17168);
and U18272 (N_18272,N_16801,N_16986);
xor U18273 (N_18273,N_17335,N_16829);
nor U18274 (N_18274,N_17607,N_17174);
nor U18275 (N_18275,N_17937,N_17843);
xnor U18276 (N_18276,N_17962,N_16589);
and U18277 (N_18277,N_16946,N_17869);
nor U18278 (N_18278,N_17310,N_17637);
or U18279 (N_18279,N_16765,N_17973);
nor U18280 (N_18280,N_17626,N_17858);
or U18281 (N_18281,N_16963,N_16654);
nor U18282 (N_18282,N_16684,N_17744);
or U18283 (N_18283,N_17871,N_17343);
xnor U18284 (N_18284,N_17737,N_17226);
nor U18285 (N_18285,N_16886,N_17291);
and U18286 (N_18286,N_17305,N_17329);
xor U18287 (N_18287,N_17181,N_17956);
or U18288 (N_18288,N_17186,N_17972);
nor U18289 (N_18289,N_17533,N_16647);
nor U18290 (N_18290,N_17476,N_17730);
xor U18291 (N_18291,N_17710,N_17815);
or U18292 (N_18292,N_17297,N_17437);
and U18293 (N_18293,N_17121,N_17645);
and U18294 (N_18294,N_17762,N_17398);
nor U18295 (N_18295,N_16557,N_17931);
xor U18296 (N_18296,N_16573,N_17861);
nand U18297 (N_18297,N_17672,N_17078);
nor U18298 (N_18298,N_17504,N_17657);
and U18299 (N_18299,N_16501,N_16809);
or U18300 (N_18300,N_16908,N_16747);
and U18301 (N_18301,N_16804,N_16913);
or U18302 (N_18302,N_17224,N_17509);
nand U18303 (N_18303,N_16729,N_17601);
and U18304 (N_18304,N_17929,N_17655);
or U18305 (N_18305,N_17170,N_17877);
or U18306 (N_18306,N_17474,N_16519);
or U18307 (N_18307,N_17564,N_17613);
and U18308 (N_18308,N_16917,N_17740);
or U18309 (N_18309,N_16775,N_17544);
xor U18310 (N_18310,N_17872,N_17755);
xor U18311 (N_18311,N_17350,N_16529);
nand U18312 (N_18312,N_17591,N_17180);
xor U18313 (N_18313,N_16736,N_16783);
and U18314 (N_18314,N_17865,N_17268);
xnor U18315 (N_18315,N_17262,N_17642);
and U18316 (N_18316,N_16785,N_16858);
nand U18317 (N_18317,N_17247,N_16944);
nor U18318 (N_18318,N_16819,N_17220);
xor U18319 (N_18319,N_16826,N_17713);
and U18320 (N_18320,N_17109,N_17097);
nand U18321 (N_18321,N_17616,N_16570);
nand U18322 (N_18322,N_17161,N_17192);
nand U18323 (N_18323,N_17980,N_17052);
and U18324 (N_18324,N_16992,N_16982);
and U18325 (N_18325,N_17429,N_17111);
and U18326 (N_18326,N_16553,N_16629);
nor U18327 (N_18327,N_17103,N_17996);
and U18328 (N_18328,N_17968,N_16670);
nor U18329 (N_18329,N_17770,N_17126);
or U18330 (N_18330,N_16790,N_17481);
or U18331 (N_18331,N_17369,N_16787);
xnor U18332 (N_18332,N_17556,N_17197);
and U18333 (N_18333,N_17416,N_17055);
nor U18334 (N_18334,N_17537,N_17548);
and U18335 (N_18335,N_16568,N_16688);
or U18336 (N_18336,N_17189,N_16693);
and U18337 (N_18337,N_17646,N_16800);
or U18338 (N_18338,N_16994,N_16667);
or U18339 (N_18339,N_17914,N_17636);
xnor U18340 (N_18340,N_17503,N_17070);
nor U18341 (N_18341,N_16839,N_17313);
and U18342 (N_18342,N_17338,N_17151);
and U18343 (N_18343,N_17695,N_17793);
nor U18344 (N_18344,N_16637,N_17047);
and U18345 (N_18345,N_17833,N_17125);
nand U18346 (N_18346,N_17628,N_16788);
nand U18347 (N_18347,N_17805,N_16660);
xor U18348 (N_18348,N_17372,N_17205);
xnor U18349 (N_18349,N_17071,N_17820);
nor U18350 (N_18350,N_17953,N_17571);
nor U18351 (N_18351,N_17374,N_17883);
and U18352 (N_18352,N_17105,N_17857);
or U18353 (N_18353,N_17345,N_17697);
or U18354 (N_18354,N_17273,N_16659);
nor U18355 (N_18355,N_17085,N_17194);
or U18356 (N_18356,N_17421,N_17414);
or U18357 (N_18357,N_16520,N_16754);
and U18358 (N_18358,N_16889,N_17302);
nand U18359 (N_18359,N_17717,N_17290);
xnor U18360 (N_18360,N_16868,N_17890);
and U18361 (N_18361,N_17270,N_17399);
or U18362 (N_18362,N_17771,N_17542);
xor U18363 (N_18363,N_17108,N_16927);
and U18364 (N_18364,N_16620,N_16936);
and U18365 (N_18365,N_17269,N_16769);
nor U18366 (N_18366,N_16613,N_17766);
xor U18367 (N_18367,N_16539,N_17784);
xor U18368 (N_18368,N_17615,N_17395);
nor U18369 (N_18369,N_17703,N_17022);
nand U18370 (N_18370,N_17230,N_17200);
or U18371 (N_18371,N_17317,N_16643);
nor U18372 (N_18372,N_16648,N_17026);
and U18373 (N_18373,N_17176,N_16588);
xor U18374 (N_18374,N_17257,N_16733);
nand U18375 (N_18375,N_16506,N_17939);
and U18376 (N_18376,N_17878,N_16965);
nor U18377 (N_18377,N_17165,N_17406);
nor U18378 (N_18378,N_16852,N_17515);
nor U18379 (N_18379,N_17614,N_16511);
nor U18380 (N_18380,N_16635,N_17586);
xor U18381 (N_18381,N_17295,N_17720);
or U18382 (N_18382,N_16518,N_17353);
or U18383 (N_18383,N_16831,N_17397);
nor U18384 (N_18384,N_16896,N_17610);
xor U18385 (N_18385,N_16948,N_17394);
nor U18386 (N_18386,N_16556,N_17119);
and U18387 (N_18387,N_17908,N_17603);
xnor U18388 (N_18388,N_16981,N_17903);
xnor U18389 (N_18389,N_17617,N_17346);
xor U18390 (N_18390,N_16624,N_17252);
or U18391 (N_18391,N_17960,N_17553);
nand U18392 (N_18392,N_17327,N_17172);
nor U18393 (N_18393,N_17198,N_17282);
nand U18394 (N_18394,N_17806,N_16774);
and U18395 (N_18395,N_16728,N_17173);
and U18396 (N_18396,N_17036,N_17099);
or U18397 (N_18397,N_17722,N_17650);
and U18398 (N_18398,N_16810,N_17955);
xnor U18399 (N_18399,N_16742,N_17498);
nor U18400 (N_18400,N_17146,N_16857);
or U18401 (N_18401,N_17652,N_17673);
nand U18402 (N_18402,N_16895,N_17315);
or U18403 (N_18403,N_16707,N_17496);
and U18404 (N_18404,N_16853,N_16543);
xnor U18405 (N_18405,N_16640,N_16866);
nor U18406 (N_18406,N_17377,N_17061);
xnor U18407 (N_18407,N_17100,N_17408);
and U18408 (N_18408,N_16975,N_17932);
nand U18409 (N_18409,N_16780,N_17101);
nor U18410 (N_18410,N_17475,N_17751);
nor U18411 (N_18411,N_16773,N_16854);
nand U18412 (N_18412,N_16630,N_16990);
nand U18413 (N_18413,N_17177,N_17348);
nand U18414 (N_18414,N_17306,N_17963);
or U18415 (N_18415,N_16658,N_17207);
or U18416 (N_18416,N_16566,N_17985);
nor U18417 (N_18417,N_17434,N_17328);
nor U18418 (N_18418,N_17705,N_17952);
nor U18419 (N_18419,N_16777,N_16892);
or U18420 (N_18420,N_17656,N_16597);
or U18421 (N_18421,N_17625,N_17012);
xor U18422 (N_18422,N_16741,N_16735);
or U18423 (N_18423,N_16581,N_17729);
and U18424 (N_18424,N_17095,N_16870);
nand U18425 (N_18425,N_16900,N_17066);
nand U18426 (N_18426,N_16910,N_17417);
nand U18427 (N_18427,N_17709,N_16757);
xnor U18428 (N_18428,N_16701,N_17401);
nand U18429 (N_18429,N_17535,N_16644);
nor U18430 (N_18430,N_16776,N_16955);
xnor U18431 (N_18431,N_16802,N_17494);
nor U18432 (N_18432,N_17534,N_17370);
nand U18433 (N_18433,N_16551,N_17765);
nand U18434 (N_18434,N_16988,N_16972);
nand U18435 (N_18435,N_17088,N_17390);
or U18436 (N_18436,N_17211,N_17236);
nor U18437 (N_18437,N_17169,N_17917);
and U18438 (N_18438,N_16847,N_17427);
and U18439 (N_18439,N_16784,N_16825);
nor U18440 (N_18440,N_17309,N_17183);
or U18441 (N_18441,N_16849,N_16920);
nor U18442 (N_18442,N_16716,N_17251);
and U18443 (N_18443,N_17945,N_17234);
and U18444 (N_18444,N_16641,N_17823);
or U18445 (N_18445,N_17365,N_16512);
nor U18446 (N_18446,N_17577,N_17255);
nor U18447 (N_18447,N_17213,N_17473);
or U18448 (N_18448,N_17404,N_17316);
xnor U18449 (N_18449,N_17976,N_17669);
and U18450 (N_18450,N_17440,N_17378);
nand U18451 (N_18451,N_17597,N_17530);
nand U18452 (N_18452,N_17943,N_17491);
nand U18453 (N_18453,N_16671,N_17735);
nand U18454 (N_18454,N_16652,N_17680);
nand U18455 (N_18455,N_17517,N_17458);
or U18456 (N_18456,N_16984,N_17215);
and U18457 (N_18457,N_16711,N_17029);
or U18458 (N_18458,N_17222,N_17293);
or U18459 (N_18459,N_16918,N_17749);
nand U18460 (N_18460,N_16695,N_17701);
nand U18461 (N_18461,N_16546,N_17357);
xor U18462 (N_18462,N_17137,N_16956);
nand U18463 (N_18463,N_17663,N_17249);
or U18464 (N_18464,N_17145,N_17831);
nor U18465 (N_18465,N_16614,N_17852);
nand U18466 (N_18466,N_17322,N_17373);
or U18467 (N_18467,N_16951,N_17570);
xnor U18468 (N_18468,N_17300,N_17726);
nor U18469 (N_18469,N_17643,N_16528);
nor U18470 (N_18470,N_17813,N_17682);
or U18471 (N_18471,N_16960,N_16594);
or U18472 (N_18472,N_17812,N_17933);
nand U18473 (N_18473,N_17519,N_17023);
nand U18474 (N_18474,N_17638,N_17167);
or U18475 (N_18475,N_16805,N_17775);
nor U18476 (N_18476,N_17388,N_16657);
nand U18477 (N_18477,N_17400,N_16676);
xor U18478 (N_18478,N_16761,N_17998);
nor U18479 (N_18479,N_16884,N_16840);
nor U18480 (N_18480,N_17331,N_17334);
or U18481 (N_18481,N_17738,N_17031);
nor U18482 (N_18482,N_17355,N_17244);
nand U18483 (N_18483,N_17238,N_16841);
or U18484 (N_18484,N_16940,N_16772);
nor U18485 (N_18485,N_17538,N_16907);
and U18486 (N_18486,N_17961,N_17899);
nand U18487 (N_18487,N_16598,N_17772);
or U18488 (N_18488,N_17144,N_17801);
and U18489 (N_18489,N_17900,N_17153);
nor U18490 (N_18490,N_17777,N_17050);
nand U18491 (N_18491,N_17011,N_16575);
nand U18492 (N_18492,N_17261,N_16552);
or U18493 (N_18493,N_17578,N_17811);
or U18494 (N_18494,N_17629,N_16584);
or U18495 (N_18495,N_17209,N_17048);
nand U18496 (N_18496,N_17977,N_17622);
or U18497 (N_18497,N_17423,N_17511);
nor U18498 (N_18498,N_17214,N_16885);
or U18499 (N_18499,N_17725,N_16745);
nor U18500 (N_18500,N_16726,N_17676);
xnor U18501 (N_18501,N_17156,N_16510);
nor U18502 (N_18502,N_17435,N_17786);
xor U18503 (N_18503,N_17587,N_17868);
nand U18504 (N_18504,N_16921,N_17058);
nor U18505 (N_18505,N_17166,N_17221);
xor U18506 (N_18506,N_17948,N_16531);
or U18507 (N_18507,N_17797,N_17500);
or U18508 (N_18508,N_17480,N_16759);
and U18509 (N_18509,N_17096,N_17593);
xor U18510 (N_18510,N_17882,N_17301);
nand U18511 (N_18511,N_17279,N_17685);
nor U18512 (N_18512,N_17934,N_16749);
nand U18513 (N_18513,N_17462,N_17563);
nand U18514 (N_18514,N_17936,N_17193);
nand U18515 (N_18515,N_16904,N_16738);
nand U18516 (N_18516,N_17450,N_17460);
xnor U18517 (N_18517,N_17759,N_17289);
nand U18518 (N_18518,N_17366,N_17651);
and U18519 (N_18519,N_16587,N_16504);
xor U18520 (N_18520,N_17449,N_17067);
xor U18521 (N_18521,N_16689,N_17319);
nor U18522 (N_18522,N_17719,N_17179);
and U18523 (N_18523,N_17658,N_16915);
nor U18524 (N_18524,N_17885,N_16950);
or U18525 (N_18525,N_17818,N_17059);
or U18526 (N_18526,N_17000,N_17696);
and U18527 (N_18527,N_17787,N_17351);
or U18528 (N_18528,N_17135,N_17566);
and U18529 (N_18529,N_17030,N_17175);
or U18530 (N_18530,N_17367,N_17501);
nand U18531 (N_18531,N_17288,N_17507);
and U18532 (N_18532,N_17359,N_17139);
nor U18533 (N_18533,N_16999,N_17441);
and U18534 (N_18534,N_17781,N_17004);
nand U18535 (N_18535,N_17037,N_16834);
and U18536 (N_18536,N_17988,N_17524);
nor U18537 (N_18537,N_17827,N_17259);
xor U18538 (N_18538,N_16903,N_17983);
xnor U18539 (N_18539,N_17648,N_16744);
xnor U18540 (N_18540,N_16666,N_17206);
and U18541 (N_18541,N_16662,N_17426);
nor U18542 (N_18542,N_17867,N_17274);
xnor U18543 (N_18543,N_17424,N_16911);
and U18544 (N_18544,N_17470,N_17880);
xnor U18545 (N_18545,N_16876,N_16822);
and U18546 (N_18546,N_16523,N_16533);
and U18547 (N_18547,N_16797,N_17199);
xor U18548 (N_18548,N_16945,N_17089);
xnor U18549 (N_18549,N_17364,N_17870);
and U18550 (N_18550,N_16699,N_17248);
nor U18551 (N_18551,N_16720,N_17433);
nand U18552 (N_18552,N_17039,N_16865);
xor U18553 (N_18553,N_17285,N_16947);
and U18554 (N_18554,N_16532,N_16953);
and U18555 (N_18555,N_17020,N_17160);
nor U18556 (N_18556,N_17013,N_17825);
nor U18557 (N_18557,N_17284,N_17362);
or U18558 (N_18558,N_17472,N_17130);
or U18559 (N_18559,N_17340,N_17120);
nor U18560 (N_18560,N_17568,N_16771);
nor U18561 (N_18561,N_17802,N_17681);
and U18562 (N_18562,N_17995,N_16949);
xor U18563 (N_18563,N_17379,N_17691);
xnor U18564 (N_18564,N_16559,N_16808);
and U18565 (N_18565,N_16828,N_16668);
or U18566 (N_18566,N_17320,N_17743);
nand U18567 (N_18567,N_17605,N_17410);
nor U18568 (N_18568,N_16521,N_17436);
xnor U18569 (N_18569,N_17439,N_17846);
xnor U18570 (N_18570,N_16985,N_16550);
or U18571 (N_18571,N_17768,N_16703);
and U18572 (N_18572,N_17062,N_16793);
and U18573 (N_18573,N_17008,N_16937);
or U18574 (N_18574,N_17001,N_17555);
nor U18575 (N_18575,N_17674,N_17966);
nor U18576 (N_18576,N_17521,N_16596);
xnor U18577 (N_18577,N_17046,N_17443);
and U18578 (N_18578,N_17114,N_16961);
nor U18579 (N_18579,N_17855,N_17589);
nor U18580 (N_18580,N_17068,N_17218);
xor U18581 (N_18581,N_17580,N_17798);
xnor U18582 (N_18582,N_17935,N_16762);
nand U18583 (N_18583,N_17464,N_16704);
or U18584 (N_18584,N_17326,N_17748);
xor U18585 (N_18585,N_17554,N_17264);
and U18586 (N_18586,N_16872,N_17216);
and U18587 (N_18587,N_17528,N_17278);
and U18588 (N_18588,N_17585,N_17463);
xnor U18589 (N_18589,N_17112,N_16878);
and U18590 (N_18590,N_17245,N_17736);
xor U18591 (N_18591,N_17584,N_16959);
nor U18592 (N_18592,N_17063,N_17539);
nor U18593 (N_18593,N_16740,N_17017);
or U18594 (N_18594,N_16683,N_17718);
xor U18595 (N_18595,N_16803,N_17142);
or U18596 (N_18596,N_17241,N_17608);
nor U18597 (N_18597,N_17134,N_16997);
xnor U18598 (N_18598,N_16952,N_17949);
nand U18599 (N_18599,N_16544,N_16678);
nand U18600 (N_18600,N_17298,N_17887);
xor U18601 (N_18601,N_17990,N_17091);
and U18602 (N_18602,N_16542,N_17916);
or U18603 (N_18603,N_16548,N_16622);
nand U18604 (N_18604,N_17630,N_17219);
xor U18605 (N_18605,N_16954,N_17644);
nand U18606 (N_18606,N_17965,N_16680);
and U18607 (N_18607,N_17579,N_16807);
and U18608 (N_18608,N_17889,N_17557);
and U18609 (N_18609,N_17640,N_16871);
nor U18610 (N_18610,N_17567,N_17888);
nand U18611 (N_18611,N_17841,N_16875);
nor U18612 (N_18612,N_16505,N_17162);
nor U18613 (N_18613,N_16979,N_16881);
and U18614 (N_18614,N_16843,N_17635);
or U18615 (N_18615,N_17263,N_16867);
or U18616 (N_18616,N_16914,N_17928);
and U18617 (N_18617,N_17021,N_17532);
nand U18618 (N_18618,N_17700,N_16891);
or U18619 (N_18619,N_16609,N_17330);
or U18620 (N_18620,N_16725,N_17203);
nand U18621 (N_18621,N_17611,N_17970);
and U18622 (N_18622,N_17723,N_16770);
xnor U18623 (N_18623,N_17347,N_16779);
nand U18624 (N_18624,N_16848,N_17040);
xnor U18625 (N_18625,N_17502,N_17256);
or U18626 (N_18626,N_17693,N_16980);
nor U18627 (N_18627,N_17832,N_17581);
nand U18628 (N_18628,N_16572,N_17283);
nand U18629 (N_18629,N_16996,N_17989);
nor U18630 (N_18630,N_17828,N_16818);
or U18631 (N_18631,N_17702,N_17898);
and U18632 (N_18632,N_17341,N_17384);
nand U18633 (N_18633,N_16628,N_17325);
nand U18634 (N_18634,N_17057,N_17767);
nand U18635 (N_18635,N_17051,N_16661);
nand U18636 (N_18636,N_17756,N_16558);
and U18637 (N_18637,N_17032,N_17490);
and U18638 (N_18638,N_17964,N_16545);
and U18639 (N_18639,N_16970,N_17569);
xor U18640 (N_18640,N_17129,N_17747);
xor U18641 (N_18641,N_16816,N_16897);
nor U18642 (N_18642,N_16755,N_17141);
xor U18643 (N_18643,N_17975,N_17791);
nand U18644 (N_18644,N_17893,N_17505);
xnor U18645 (N_18645,N_17413,N_16766);
and U18646 (N_18646,N_17242,N_17138);
and U18647 (N_18647,N_16923,N_17148);
xor U18648 (N_18648,N_16526,N_16636);
xor U18649 (N_18649,N_16880,N_17848);
and U18650 (N_18650,N_16645,N_16987);
nor U18651 (N_18651,N_17844,N_17950);
nand U18652 (N_18652,N_17158,N_17127);
or U18653 (N_18653,N_17853,N_17711);
or U18654 (N_18654,N_16610,N_16750);
nand U18655 (N_18655,N_16973,N_17526);
nand U18656 (N_18656,N_17246,N_17757);
and U18657 (N_18657,N_17912,N_17910);
xnor U18658 (N_18658,N_17025,N_17391);
xnor U18659 (N_18659,N_17308,N_16576);
nor U18660 (N_18660,N_17356,N_17739);
and U18661 (N_18661,N_17381,N_17923);
xnor U18662 (N_18662,N_16814,N_17184);
or U18663 (N_18663,N_17845,N_16874);
and U18664 (N_18664,N_16593,N_16547);
nand U18665 (N_18665,N_16851,N_17959);
or U18666 (N_18666,N_17671,N_16863);
and U18667 (N_18667,N_17562,N_16781);
or U18668 (N_18668,N_16685,N_17280);
nor U18669 (N_18669,N_16942,N_17253);
nand U18670 (N_18670,N_16967,N_17411);
xnor U18671 (N_18671,N_17045,N_16672);
nand U18672 (N_18672,N_17077,N_16806);
nand U18673 (N_18673,N_17745,N_17716);
nor U18674 (N_18674,N_17951,N_17466);
nand U18675 (N_18675,N_16899,N_16856);
and U18676 (N_18676,N_17235,N_17363);
nand U18677 (N_18677,N_17819,N_16832);
or U18678 (N_18678,N_16617,N_17403);
xnor U18679 (N_18679,N_17469,N_17758);
nand U18680 (N_18680,N_17905,N_16898);
xor U18681 (N_18681,N_17545,N_17208);
or U18682 (N_18682,N_16743,N_17780);
or U18683 (N_18683,N_17814,N_17499);
and U18684 (N_18684,N_17895,N_17619);
or U18685 (N_18685,N_17575,N_17677);
nand U18686 (N_18686,N_17034,N_17874);
and U18687 (N_18687,N_16700,N_16932);
nor U18688 (N_18688,N_17237,N_17875);
nand U18689 (N_18689,N_17901,N_17281);
nor U18690 (N_18690,N_17223,N_16723);
or U18691 (N_18691,N_17541,N_17149);
nor U18692 (N_18692,N_16798,N_17182);
and U18693 (N_18693,N_17407,N_17191);
xor U18694 (N_18694,N_16739,N_17795);
or U18695 (N_18695,N_17072,N_16838);
nand U18696 (N_18696,N_17728,N_16608);
xnor U18697 (N_18697,N_17776,N_17042);
nand U18698 (N_18698,N_17896,N_17707);
nand U18699 (N_18699,N_16968,N_17106);
and U18700 (N_18700,N_17143,N_17690);
nor U18701 (N_18701,N_17276,N_16507);
xor U18702 (N_18702,N_17430,N_16712);
and U18703 (N_18703,N_17113,N_17830);
nor U18704 (N_18704,N_17919,N_17944);
nand U18705 (N_18705,N_17483,N_17477);
xnor U18706 (N_18706,N_17382,N_17299);
nor U18707 (N_18707,N_17304,N_17940);
or U18708 (N_18708,N_16882,N_16978);
and U18709 (N_18709,N_17978,N_17420);
nor U18710 (N_18710,N_17442,N_17425);
and U18711 (N_18711,N_17349,N_16721);
or U18712 (N_18712,N_16591,N_17479);
or U18713 (N_18713,N_17991,N_16815);
or U18714 (N_18714,N_17239,N_16561);
nand U18715 (N_18715,N_17332,N_17543);
nor U18716 (N_18716,N_17708,N_17859);
or U18717 (N_18717,N_17731,N_17227);
and U18718 (N_18718,N_17712,N_17836);
nor U18719 (N_18719,N_17684,N_17296);
or U18720 (N_18720,N_16522,N_17272);
nor U18721 (N_18721,N_17467,N_17336);
and U18722 (N_18722,N_17489,N_16795);
nand U18723 (N_18723,N_16966,N_16713);
nor U18724 (N_18724,N_17514,N_17484);
or U18725 (N_18725,N_17508,N_17824);
and U18726 (N_18726,N_16864,N_16862);
or U18727 (N_18727,N_17907,N_16993);
and U18728 (N_18728,N_16696,N_16879);
nand U18729 (N_18729,N_16538,N_16919);
xor U18730 (N_18730,N_17536,N_17393);
nor U18731 (N_18731,N_16989,N_17560);
nor U18732 (N_18732,N_17520,N_17788);
xnor U18733 (N_18733,N_17294,N_16844);
and U18734 (N_18734,N_16649,N_17654);
or U18735 (N_18735,N_17465,N_16535);
nor U18736 (N_18736,N_17178,N_17773);
nor U18737 (N_18737,N_17082,N_17459);
xnor U18738 (N_18738,N_17835,N_16837);
xnor U18739 (N_18739,N_17704,N_17779);
nand U18740 (N_18740,N_16929,N_17016);
xnor U18741 (N_18741,N_17921,N_17822);
and U18742 (N_18742,N_17314,N_17915);
nand U18743 (N_18743,N_17056,N_17957);
and U18744 (N_18744,N_16638,N_17789);
or U18745 (N_18745,N_17860,N_17090);
xnor U18746 (N_18746,N_17862,N_16577);
nand U18747 (N_18747,N_17323,N_16655);
xor U18748 (N_18748,N_16682,N_16530);
or U18749 (N_18749,N_17574,N_16905);
xnor U18750 (N_18750,N_17693,N_16994);
or U18751 (N_18751,N_16786,N_16847);
nor U18752 (N_18752,N_17711,N_17988);
nand U18753 (N_18753,N_16821,N_16666);
nor U18754 (N_18754,N_16833,N_17403);
nand U18755 (N_18755,N_16682,N_17332);
xnor U18756 (N_18756,N_17111,N_17953);
nor U18757 (N_18757,N_17464,N_17575);
xor U18758 (N_18758,N_17114,N_17935);
nor U18759 (N_18759,N_17296,N_17396);
or U18760 (N_18760,N_17041,N_17255);
nand U18761 (N_18761,N_16802,N_16750);
nand U18762 (N_18762,N_17325,N_16544);
nor U18763 (N_18763,N_17252,N_16746);
nand U18764 (N_18764,N_17195,N_17459);
nand U18765 (N_18765,N_16716,N_16753);
nand U18766 (N_18766,N_17206,N_16781);
nand U18767 (N_18767,N_17310,N_16662);
nor U18768 (N_18768,N_17190,N_17486);
nand U18769 (N_18769,N_16842,N_17595);
nand U18770 (N_18770,N_17616,N_16561);
nand U18771 (N_18771,N_17264,N_16819);
xor U18772 (N_18772,N_17792,N_16936);
nor U18773 (N_18773,N_17537,N_17415);
xor U18774 (N_18774,N_17699,N_17648);
nor U18775 (N_18775,N_17458,N_17173);
nor U18776 (N_18776,N_16764,N_17992);
and U18777 (N_18777,N_17967,N_17818);
xnor U18778 (N_18778,N_17735,N_17082);
xnor U18779 (N_18779,N_16928,N_17110);
nand U18780 (N_18780,N_16895,N_17520);
xor U18781 (N_18781,N_17771,N_17071);
and U18782 (N_18782,N_17586,N_16979);
or U18783 (N_18783,N_17362,N_17110);
nor U18784 (N_18784,N_17180,N_17854);
nand U18785 (N_18785,N_16863,N_16722);
nor U18786 (N_18786,N_17871,N_16679);
and U18787 (N_18787,N_16728,N_17345);
nand U18788 (N_18788,N_17805,N_17220);
nor U18789 (N_18789,N_17617,N_17892);
xnor U18790 (N_18790,N_17825,N_16624);
nor U18791 (N_18791,N_16719,N_17420);
xor U18792 (N_18792,N_17499,N_17285);
xnor U18793 (N_18793,N_16561,N_17773);
nor U18794 (N_18794,N_17824,N_17799);
nor U18795 (N_18795,N_17139,N_17659);
nand U18796 (N_18796,N_16626,N_17568);
nor U18797 (N_18797,N_16592,N_16671);
nor U18798 (N_18798,N_17559,N_17048);
nand U18799 (N_18799,N_16710,N_17691);
nor U18800 (N_18800,N_16805,N_17715);
nand U18801 (N_18801,N_17183,N_17600);
or U18802 (N_18802,N_17835,N_17060);
nand U18803 (N_18803,N_16581,N_17112);
and U18804 (N_18804,N_16805,N_17048);
xnor U18805 (N_18805,N_17149,N_17337);
xor U18806 (N_18806,N_17581,N_16664);
nand U18807 (N_18807,N_17164,N_16509);
and U18808 (N_18808,N_16666,N_17330);
nand U18809 (N_18809,N_16939,N_17663);
and U18810 (N_18810,N_16897,N_16618);
xor U18811 (N_18811,N_16886,N_17463);
nor U18812 (N_18812,N_16782,N_16520);
xnor U18813 (N_18813,N_17050,N_17311);
or U18814 (N_18814,N_17666,N_16714);
nand U18815 (N_18815,N_16932,N_17362);
and U18816 (N_18816,N_16516,N_17548);
nor U18817 (N_18817,N_17578,N_17488);
and U18818 (N_18818,N_16972,N_17323);
or U18819 (N_18819,N_16925,N_17624);
xor U18820 (N_18820,N_17861,N_17849);
nand U18821 (N_18821,N_17718,N_17028);
nand U18822 (N_18822,N_17465,N_17414);
or U18823 (N_18823,N_17129,N_16969);
and U18824 (N_18824,N_17273,N_17809);
xnor U18825 (N_18825,N_16936,N_16706);
or U18826 (N_18826,N_16961,N_16913);
nand U18827 (N_18827,N_16870,N_17057);
nand U18828 (N_18828,N_17942,N_17997);
xnor U18829 (N_18829,N_17164,N_17040);
xor U18830 (N_18830,N_16610,N_17058);
or U18831 (N_18831,N_16521,N_17326);
nand U18832 (N_18832,N_16726,N_16819);
nand U18833 (N_18833,N_17452,N_17477);
nor U18834 (N_18834,N_17207,N_17134);
and U18835 (N_18835,N_16639,N_17820);
or U18836 (N_18836,N_17379,N_17440);
nand U18837 (N_18837,N_17456,N_17096);
or U18838 (N_18838,N_17886,N_17360);
nand U18839 (N_18839,N_17638,N_17434);
and U18840 (N_18840,N_17758,N_17457);
or U18841 (N_18841,N_17726,N_17776);
xnor U18842 (N_18842,N_16902,N_16593);
and U18843 (N_18843,N_17323,N_17404);
nor U18844 (N_18844,N_17894,N_16601);
nor U18845 (N_18845,N_16580,N_17389);
nand U18846 (N_18846,N_17037,N_16956);
and U18847 (N_18847,N_16614,N_17000);
nor U18848 (N_18848,N_16779,N_16621);
xor U18849 (N_18849,N_16979,N_17050);
and U18850 (N_18850,N_17882,N_16986);
nand U18851 (N_18851,N_17538,N_17919);
nand U18852 (N_18852,N_16696,N_17845);
xor U18853 (N_18853,N_17739,N_17961);
xnor U18854 (N_18854,N_17851,N_16888);
or U18855 (N_18855,N_17753,N_17585);
nor U18856 (N_18856,N_16700,N_17497);
nor U18857 (N_18857,N_17187,N_17301);
and U18858 (N_18858,N_16525,N_17451);
nand U18859 (N_18859,N_16963,N_17498);
xor U18860 (N_18860,N_17286,N_17750);
nand U18861 (N_18861,N_17915,N_16941);
and U18862 (N_18862,N_17339,N_17996);
and U18863 (N_18863,N_17191,N_16610);
nor U18864 (N_18864,N_17502,N_16697);
nand U18865 (N_18865,N_17817,N_17054);
nor U18866 (N_18866,N_17450,N_16784);
and U18867 (N_18867,N_17735,N_17669);
xnor U18868 (N_18868,N_16526,N_16597);
nand U18869 (N_18869,N_16724,N_16873);
or U18870 (N_18870,N_16961,N_17756);
and U18871 (N_18871,N_16560,N_17543);
nand U18872 (N_18872,N_17043,N_16536);
nand U18873 (N_18873,N_16615,N_17623);
or U18874 (N_18874,N_16522,N_17970);
nand U18875 (N_18875,N_16895,N_16802);
and U18876 (N_18876,N_16901,N_16884);
xor U18877 (N_18877,N_17052,N_16921);
nor U18878 (N_18878,N_17035,N_17549);
nand U18879 (N_18879,N_17951,N_17520);
and U18880 (N_18880,N_17782,N_17094);
nor U18881 (N_18881,N_16749,N_16654);
or U18882 (N_18882,N_17844,N_17537);
and U18883 (N_18883,N_17787,N_17072);
and U18884 (N_18884,N_17228,N_16646);
nand U18885 (N_18885,N_17547,N_17640);
nor U18886 (N_18886,N_16798,N_17082);
nand U18887 (N_18887,N_17672,N_16820);
nor U18888 (N_18888,N_17688,N_16785);
xor U18889 (N_18889,N_17313,N_17573);
nor U18890 (N_18890,N_16722,N_17730);
xor U18891 (N_18891,N_16943,N_17278);
or U18892 (N_18892,N_17812,N_17652);
xnor U18893 (N_18893,N_16873,N_17314);
nand U18894 (N_18894,N_16793,N_17036);
nand U18895 (N_18895,N_17571,N_16822);
nor U18896 (N_18896,N_16666,N_17726);
xnor U18897 (N_18897,N_17725,N_17208);
nand U18898 (N_18898,N_17004,N_16856);
nand U18899 (N_18899,N_17658,N_17400);
or U18900 (N_18900,N_17562,N_17734);
or U18901 (N_18901,N_17053,N_16959);
xor U18902 (N_18902,N_17841,N_17254);
or U18903 (N_18903,N_17315,N_17382);
and U18904 (N_18904,N_17481,N_16586);
and U18905 (N_18905,N_17636,N_17595);
nand U18906 (N_18906,N_16593,N_17333);
and U18907 (N_18907,N_17872,N_16954);
or U18908 (N_18908,N_17507,N_17840);
or U18909 (N_18909,N_17031,N_16765);
nand U18910 (N_18910,N_17311,N_16800);
nor U18911 (N_18911,N_17811,N_17663);
or U18912 (N_18912,N_17214,N_17871);
xor U18913 (N_18913,N_16716,N_17881);
nand U18914 (N_18914,N_17972,N_16559);
nand U18915 (N_18915,N_17162,N_16887);
xnor U18916 (N_18916,N_17343,N_17360);
or U18917 (N_18917,N_16901,N_17003);
and U18918 (N_18918,N_16805,N_17211);
nor U18919 (N_18919,N_17545,N_17404);
nor U18920 (N_18920,N_17356,N_17878);
nand U18921 (N_18921,N_17233,N_17131);
nand U18922 (N_18922,N_16825,N_17851);
nand U18923 (N_18923,N_16650,N_17785);
xnor U18924 (N_18924,N_16769,N_17167);
or U18925 (N_18925,N_17276,N_16755);
nand U18926 (N_18926,N_17598,N_17706);
xnor U18927 (N_18927,N_17815,N_17724);
nand U18928 (N_18928,N_16885,N_16717);
and U18929 (N_18929,N_17401,N_17280);
nor U18930 (N_18930,N_17857,N_17617);
and U18931 (N_18931,N_16622,N_16637);
nand U18932 (N_18932,N_17293,N_17528);
or U18933 (N_18933,N_16933,N_17568);
xnor U18934 (N_18934,N_17352,N_17629);
xor U18935 (N_18935,N_17078,N_17068);
nand U18936 (N_18936,N_17373,N_16786);
or U18937 (N_18937,N_16917,N_16663);
and U18938 (N_18938,N_17793,N_17053);
nor U18939 (N_18939,N_17172,N_17522);
and U18940 (N_18940,N_16517,N_17816);
xnor U18941 (N_18941,N_17314,N_16840);
or U18942 (N_18942,N_17873,N_16962);
nor U18943 (N_18943,N_17768,N_16913);
nand U18944 (N_18944,N_17013,N_16853);
nand U18945 (N_18945,N_16814,N_17368);
nand U18946 (N_18946,N_16508,N_17606);
nand U18947 (N_18947,N_17662,N_17804);
xor U18948 (N_18948,N_17882,N_17905);
or U18949 (N_18949,N_17892,N_16539);
xnor U18950 (N_18950,N_17488,N_17191);
nand U18951 (N_18951,N_16542,N_17099);
and U18952 (N_18952,N_17934,N_17822);
xnor U18953 (N_18953,N_17993,N_17852);
and U18954 (N_18954,N_17412,N_16679);
nor U18955 (N_18955,N_17537,N_16701);
or U18956 (N_18956,N_17275,N_16891);
or U18957 (N_18957,N_17602,N_16633);
nand U18958 (N_18958,N_17892,N_17781);
nor U18959 (N_18959,N_17787,N_16949);
xor U18960 (N_18960,N_17828,N_17275);
nor U18961 (N_18961,N_17313,N_16550);
and U18962 (N_18962,N_17659,N_17327);
nand U18963 (N_18963,N_17665,N_17791);
xnor U18964 (N_18964,N_17149,N_16889);
or U18965 (N_18965,N_17073,N_16632);
xnor U18966 (N_18966,N_16661,N_16779);
nand U18967 (N_18967,N_16913,N_17086);
and U18968 (N_18968,N_17638,N_17619);
xnor U18969 (N_18969,N_17879,N_17994);
and U18970 (N_18970,N_17092,N_17604);
xnor U18971 (N_18971,N_17779,N_16831);
nor U18972 (N_18972,N_17142,N_16827);
nor U18973 (N_18973,N_16832,N_17459);
nand U18974 (N_18974,N_16557,N_17166);
nand U18975 (N_18975,N_17564,N_17659);
or U18976 (N_18976,N_17890,N_17913);
and U18977 (N_18977,N_17967,N_16726);
nand U18978 (N_18978,N_16678,N_17416);
nor U18979 (N_18979,N_17854,N_17666);
and U18980 (N_18980,N_16834,N_16520);
nor U18981 (N_18981,N_16599,N_16833);
nor U18982 (N_18982,N_17805,N_17605);
nand U18983 (N_18983,N_17612,N_17676);
nand U18984 (N_18984,N_17829,N_17627);
or U18985 (N_18985,N_17490,N_17600);
and U18986 (N_18986,N_17613,N_17711);
or U18987 (N_18987,N_16991,N_17769);
or U18988 (N_18988,N_17976,N_17702);
and U18989 (N_18989,N_17455,N_17827);
xnor U18990 (N_18990,N_16942,N_16706);
xnor U18991 (N_18991,N_17610,N_16754);
xor U18992 (N_18992,N_17869,N_16805);
nor U18993 (N_18993,N_17127,N_16993);
nor U18994 (N_18994,N_17112,N_16625);
nor U18995 (N_18995,N_17671,N_16857);
or U18996 (N_18996,N_17715,N_17538);
nor U18997 (N_18997,N_16504,N_16561);
and U18998 (N_18998,N_17387,N_17657);
nor U18999 (N_18999,N_16659,N_17702);
nor U19000 (N_19000,N_17760,N_16911);
and U19001 (N_19001,N_17796,N_17510);
xnor U19002 (N_19002,N_17264,N_17695);
nand U19003 (N_19003,N_16980,N_17131);
nand U19004 (N_19004,N_17882,N_17979);
or U19005 (N_19005,N_17156,N_17453);
and U19006 (N_19006,N_17582,N_16769);
xor U19007 (N_19007,N_17820,N_17275);
nor U19008 (N_19008,N_17002,N_16877);
nor U19009 (N_19009,N_17508,N_17846);
xor U19010 (N_19010,N_16557,N_17140);
xor U19011 (N_19011,N_17238,N_16812);
nor U19012 (N_19012,N_17950,N_16517);
or U19013 (N_19013,N_16556,N_17241);
nand U19014 (N_19014,N_17187,N_16632);
xor U19015 (N_19015,N_17027,N_17557);
and U19016 (N_19016,N_16923,N_17623);
nand U19017 (N_19017,N_16986,N_17894);
or U19018 (N_19018,N_16603,N_17948);
or U19019 (N_19019,N_17632,N_17002);
nand U19020 (N_19020,N_17756,N_17848);
or U19021 (N_19021,N_16814,N_17269);
and U19022 (N_19022,N_17072,N_17709);
or U19023 (N_19023,N_17053,N_16768);
or U19024 (N_19024,N_17262,N_17460);
nor U19025 (N_19025,N_17645,N_17776);
nand U19026 (N_19026,N_17372,N_16954);
xor U19027 (N_19027,N_17353,N_16981);
xor U19028 (N_19028,N_17746,N_17505);
and U19029 (N_19029,N_17219,N_16525);
or U19030 (N_19030,N_16955,N_17600);
nor U19031 (N_19031,N_16554,N_16995);
nor U19032 (N_19032,N_16894,N_17279);
or U19033 (N_19033,N_17114,N_17648);
xor U19034 (N_19034,N_17439,N_16531);
xor U19035 (N_19035,N_17443,N_16537);
nor U19036 (N_19036,N_17097,N_17526);
nor U19037 (N_19037,N_17829,N_17090);
and U19038 (N_19038,N_17821,N_17658);
or U19039 (N_19039,N_17397,N_16591);
or U19040 (N_19040,N_17579,N_17468);
nand U19041 (N_19041,N_17704,N_16842);
nand U19042 (N_19042,N_17063,N_16776);
and U19043 (N_19043,N_17164,N_17301);
nand U19044 (N_19044,N_17885,N_16755);
xor U19045 (N_19045,N_17802,N_16683);
and U19046 (N_19046,N_17309,N_17662);
nor U19047 (N_19047,N_17731,N_17875);
xor U19048 (N_19048,N_16518,N_16652);
or U19049 (N_19049,N_17151,N_16784);
nor U19050 (N_19050,N_17426,N_17767);
xor U19051 (N_19051,N_17033,N_17187);
and U19052 (N_19052,N_16836,N_16846);
xnor U19053 (N_19053,N_16886,N_17422);
xor U19054 (N_19054,N_16971,N_16984);
xnor U19055 (N_19055,N_17504,N_17043);
or U19056 (N_19056,N_17348,N_17295);
and U19057 (N_19057,N_17608,N_17429);
xnor U19058 (N_19058,N_16558,N_17868);
xnor U19059 (N_19059,N_16812,N_17743);
nand U19060 (N_19060,N_17435,N_16814);
xor U19061 (N_19061,N_17758,N_17190);
and U19062 (N_19062,N_17063,N_16919);
nor U19063 (N_19063,N_16652,N_16954);
or U19064 (N_19064,N_16521,N_17429);
and U19065 (N_19065,N_16716,N_16564);
nor U19066 (N_19066,N_17514,N_17471);
or U19067 (N_19067,N_17033,N_17951);
nor U19068 (N_19068,N_17433,N_16608);
nand U19069 (N_19069,N_17705,N_17583);
xor U19070 (N_19070,N_16555,N_16780);
and U19071 (N_19071,N_17869,N_17944);
or U19072 (N_19072,N_16891,N_17040);
or U19073 (N_19073,N_16694,N_17186);
or U19074 (N_19074,N_16536,N_16952);
nor U19075 (N_19075,N_17762,N_17697);
xor U19076 (N_19076,N_16996,N_16694);
nor U19077 (N_19077,N_17471,N_17972);
nor U19078 (N_19078,N_17199,N_16549);
xnor U19079 (N_19079,N_16667,N_17378);
nand U19080 (N_19080,N_17403,N_16845);
or U19081 (N_19081,N_16722,N_16529);
nand U19082 (N_19082,N_16794,N_17996);
xor U19083 (N_19083,N_16859,N_17708);
nor U19084 (N_19084,N_17545,N_17319);
or U19085 (N_19085,N_17017,N_17392);
or U19086 (N_19086,N_16563,N_16618);
xnor U19087 (N_19087,N_17103,N_17671);
or U19088 (N_19088,N_17072,N_17806);
and U19089 (N_19089,N_17073,N_17318);
xor U19090 (N_19090,N_17451,N_17726);
nand U19091 (N_19091,N_17281,N_17391);
xnor U19092 (N_19092,N_16996,N_17014);
nor U19093 (N_19093,N_16660,N_16706);
xnor U19094 (N_19094,N_17438,N_16813);
or U19095 (N_19095,N_17366,N_17168);
or U19096 (N_19096,N_17389,N_17155);
and U19097 (N_19097,N_17473,N_17240);
nand U19098 (N_19098,N_17319,N_17245);
nor U19099 (N_19099,N_16869,N_17459);
nand U19100 (N_19100,N_16797,N_17832);
xor U19101 (N_19101,N_17581,N_16885);
xor U19102 (N_19102,N_16622,N_17450);
and U19103 (N_19103,N_17044,N_17576);
and U19104 (N_19104,N_17041,N_17674);
or U19105 (N_19105,N_17404,N_17664);
and U19106 (N_19106,N_17963,N_17360);
or U19107 (N_19107,N_17413,N_17776);
nor U19108 (N_19108,N_17281,N_17318);
and U19109 (N_19109,N_17678,N_16797);
nand U19110 (N_19110,N_17509,N_16688);
and U19111 (N_19111,N_17255,N_17367);
xor U19112 (N_19112,N_16664,N_17243);
nor U19113 (N_19113,N_17396,N_17684);
xor U19114 (N_19114,N_17678,N_17081);
nand U19115 (N_19115,N_16672,N_17245);
xor U19116 (N_19116,N_16705,N_17931);
and U19117 (N_19117,N_17630,N_16750);
nor U19118 (N_19118,N_16548,N_17370);
and U19119 (N_19119,N_16904,N_16503);
and U19120 (N_19120,N_17030,N_17333);
and U19121 (N_19121,N_17401,N_17037);
nand U19122 (N_19122,N_16691,N_17939);
xnor U19123 (N_19123,N_16631,N_16863);
xnor U19124 (N_19124,N_16939,N_16843);
xnor U19125 (N_19125,N_16938,N_17826);
xnor U19126 (N_19126,N_17306,N_17856);
nand U19127 (N_19127,N_16581,N_16870);
or U19128 (N_19128,N_17304,N_17945);
and U19129 (N_19129,N_17004,N_17430);
or U19130 (N_19130,N_16533,N_17530);
and U19131 (N_19131,N_16585,N_16659);
nand U19132 (N_19132,N_16621,N_17613);
and U19133 (N_19133,N_17768,N_16628);
nand U19134 (N_19134,N_16590,N_16657);
nor U19135 (N_19135,N_16939,N_16944);
nand U19136 (N_19136,N_16995,N_16791);
nor U19137 (N_19137,N_16813,N_16733);
xnor U19138 (N_19138,N_16836,N_17862);
nor U19139 (N_19139,N_17930,N_16708);
nand U19140 (N_19140,N_16608,N_17156);
or U19141 (N_19141,N_16886,N_17261);
xor U19142 (N_19142,N_16832,N_17672);
or U19143 (N_19143,N_16576,N_17848);
nand U19144 (N_19144,N_16518,N_17930);
or U19145 (N_19145,N_17901,N_17313);
nor U19146 (N_19146,N_17215,N_17207);
xor U19147 (N_19147,N_17272,N_17646);
xor U19148 (N_19148,N_16594,N_17412);
xnor U19149 (N_19149,N_16944,N_17205);
xor U19150 (N_19150,N_16818,N_17824);
nand U19151 (N_19151,N_17931,N_17221);
nand U19152 (N_19152,N_17606,N_17425);
xnor U19153 (N_19153,N_17027,N_17752);
nor U19154 (N_19154,N_16658,N_16551);
or U19155 (N_19155,N_17671,N_17116);
nor U19156 (N_19156,N_17566,N_17728);
xor U19157 (N_19157,N_17687,N_17681);
or U19158 (N_19158,N_17840,N_17128);
and U19159 (N_19159,N_17431,N_17767);
nor U19160 (N_19160,N_17341,N_16997);
nand U19161 (N_19161,N_17798,N_16953);
and U19162 (N_19162,N_16652,N_17879);
nor U19163 (N_19163,N_16800,N_17432);
xor U19164 (N_19164,N_17146,N_17319);
nand U19165 (N_19165,N_16819,N_17523);
or U19166 (N_19166,N_16728,N_16617);
nor U19167 (N_19167,N_16746,N_17593);
xnor U19168 (N_19168,N_17163,N_17766);
xor U19169 (N_19169,N_16679,N_16621);
xor U19170 (N_19170,N_17818,N_17619);
nand U19171 (N_19171,N_17227,N_16620);
nor U19172 (N_19172,N_17113,N_17238);
nor U19173 (N_19173,N_16940,N_17086);
and U19174 (N_19174,N_17637,N_16535);
and U19175 (N_19175,N_17064,N_16623);
nor U19176 (N_19176,N_17643,N_17628);
nand U19177 (N_19177,N_16548,N_16592);
nand U19178 (N_19178,N_17395,N_16904);
xnor U19179 (N_19179,N_17644,N_17128);
or U19180 (N_19180,N_17237,N_16807);
xnor U19181 (N_19181,N_16797,N_16909);
nand U19182 (N_19182,N_17641,N_17830);
or U19183 (N_19183,N_17327,N_17885);
nand U19184 (N_19184,N_17360,N_17501);
nor U19185 (N_19185,N_17582,N_17740);
nor U19186 (N_19186,N_17362,N_16908);
xnor U19187 (N_19187,N_16881,N_17112);
and U19188 (N_19188,N_16973,N_16584);
nand U19189 (N_19189,N_16630,N_16678);
xnor U19190 (N_19190,N_17289,N_17548);
nand U19191 (N_19191,N_17505,N_17280);
xnor U19192 (N_19192,N_17856,N_16536);
xor U19193 (N_19193,N_16635,N_17420);
nand U19194 (N_19194,N_17643,N_17805);
nor U19195 (N_19195,N_17829,N_17764);
and U19196 (N_19196,N_17201,N_17375);
nand U19197 (N_19197,N_16809,N_17366);
and U19198 (N_19198,N_16753,N_16893);
and U19199 (N_19199,N_16821,N_17311);
nor U19200 (N_19200,N_17455,N_16826);
nor U19201 (N_19201,N_17779,N_17436);
or U19202 (N_19202,N_17905,N_16923);
nand U19203 (N_19203,N_17755,N_16609);
nand U19204 (N_19204,N_17913,N_16584);
and U19205 (N_19205,N_17817,N_17910);
or U19206 (N_19206,N_17029,N_16817);
and U19207 (N_19207,N_16743,N_17293);
xor U19208 (N_19208,N_16807,N_16993);
nor U19209 (N_19209,N_16788,N_17912);
or U19210 (N_19210,N_17673,N_17045);
and U19211 (N_19211,N_16801,N_17003);
nand U19212 (N_19212,N_17619,N_17041);
nor U19213 (N_19213,N_16909,N_17479);
nand U19214 (N_19214,N_17983,N_17670);
and U19215 (N_19215,N_17585,N_16739);
nor U19216 (N_19216,N_17207,N_17948);
or U19217 (N_19217,N_16972,N_17155);
nor U19218 (N_19218,N_17158,N_16733);
or U19219 (N_19219,N_17630,N_17056);
and U19220 (N_19220,N_17494,N_16627);
xor U19221 (N_19221,N_16558,N_17714);
nand U19222 (N_19222,N_17126,N_17378);
xor U19223 (N_19223,N_16783,N_16857);
or U19224 (N_19224,N_17203,N_17766);
xnor U19225 (N_19225,N_17254,N_17363);
xor U19226 (N_19226,N_16911,N_16699);
nor U19227 (N_19227,N_17667,N_16916);
nor U19228 (N_19228,N_17721,N_17773);
and U19229 (N_19229,N_17417,N_16893);
xor U19230 (N_19230,N_17823,N_17863);
and U19231 (N_19231,N_17425,N_17403);
xor U19232 (N_19232,N_17448,N_17249);
nand U19233 (N_19233,N_17490,N_17010);
nand U19234 (N_19234,N_17988,N_17149);
nor U19235 (N_19235,N_17176,N_17713);
nand U19236 (N_19236,N_17468,N_17661);
xor U19237 (N_19237,N_17950,N_17886);
nand U19238 (N_19238,N_17975,N_17969);
and U19239 (N_19239,N_16910,N_16935);
xor U19240 (N_19240,N_17656,N_17291);
and U19241 (N_19241,N_17504,N_16653);
or U19242 (N_19242,N_16605,N_17124);
nor U19243 (N_19243,N_16680,N_17253);
or U19244 (N_19244,N_16846,N_17673);
nor U19245 (N_19245,N_16845,N_17991);
nand U19246 (N_19246,N_17502,N_17328);
xnor U19247 (N_19247,N_17923,N_17960);
nand U19248 (N_19248,N_17023,N_16582);
xor U19249 (N_19249,N_17892,N_16890);
and U19250 (N_19250,N_17701,N_16693);
nand U19251 (N_19251,N_17995,N_16800);
xnor U19252 (N_19252,N_17758,N_16597);
xor U19253 (N_19253,N_17003,N_17036);
nor U19254 (N_19254,N_17804,N_16630);
or U19255 (N_19255,N_17990,N_17178);
nand U19256 (N_19256,N_16808,N_17926);
nor U19257 (N_19257,N_16736,N_17230);
and U19258 (N_19258,N_17281,N_17273);
or U19259 (N_19259,N_17949,N_16725);
or U19260 (N_19260,N_16886,N_16858);
xnor U19261 (N_19261,N_16601,N_17686);
nor U19262 (N_19262,N_17359,N_17809);
nor U19263 (N_19263,N_17108,N_17463);
nor U19264 (N_19264,N_17842,N_17368);
xor U19265 (N_19265,N_17792,N_17699);
nor U19266 (N_19266,N_17999,N_17563);
nor U19267 (N_19267,N_17066,N_17344);
xnor U19268 (N_19268,N_17134,N_17089);
nor U19269 (N_19269,N_17725,N_17235);
and U19270 (N_19270,N_17716,N_17751);
nor U19271 (N_19271,N_17809,N_16860);
or U19272 (N_19272,N_17289,N_16849);
or U19273 (N_19273,N_17753,N_16903);
and U19274 (N_19274,N_17237,N_17840);
xor U19275 (N_19275,N_17586,N_17545);
nor U19276 (N_19276,N_16759,N_17845);
or U19277 (N_19277,N_17954,N_16628);
or U19278 (N_19278,N_17278,N_17746);
nor U19279 (N_19279,N_16718,N_17697);
and U19280 (N_19280,N_16570,N_17426);
nand U19281 (N_19281,N_17463,N_17999);
nor U19282 (N_19282,N_16842,N_16901);
xor U19283 (N_19283,N_17044,N_17422);
xor U19284 (N_19284,N_16809,N_17428);
nor U19285 (N_19285,N_16851,N_17007);
and U19286 (N_19286,N_16906,N_16702);
nor U19287 (N_19287,N_17739,N_17900);
nand U19288 (N_19288,N_16750,N_17099);
nor U19289 (N_19289,N_17156,N_17516);
nor U19290 (N_19290,N_16752,N_17103);
or U19291 (N_19291,N_16816,N_16959);
nand U19292 (N_19292,N_17689,N_17812);
and U19293 (N_19293,N_17632,N_16975);
nor U19294 (N_19294,N_16567,N_16561);
and U19295 (N_19295,N_17877,N_16845);
and U19296 (N_19296,N_17978,N_17898);
nand U19297 (N_19297,N_17250,N_17594);
and U19298 (N_19298,N_17855,N_17463);
xnor U19299 (N_19299,N_17700,N_16712);
nor U19300 (N_19300,N_17026,N_17136);
nor U19301 (N_19301,N_16501,N_17370);
and U19302 (N_19302,N_17827,N_17716);
xnor U19303 (N_19303,N_17711,N_17977);
nor U19304 (N_19304,N_16630,N_17551);
and U19305 (N_19305,N_17633,N_17396);
xnor U19306 (N_19306,N_17100,N_17497);
xnor U19307 (N_19307,N_17810,N_16941);
xor U19308 (N_19308,N_17228,N_17148);
or U19309 (N_19309,N_17868,N_17395);
nor U19310 (N_19310,N_17943,N_16860);
xnor U19311 (N_19311,N_17809,N_17120);
or U19312 (N_19312,N_17855,N_17816);
xnor U19313 (N_19313,N_17566,N_16776);
and U19314 (N_19314,N_16540,N_17774);
xor U19315 (N_19315,N_17689,N_17969);
xnor U19316 (N_19316,N_16514,N_16561);
or U19317 (N_19317,N_17785,N_16549);
nor U19318 (N_19318,N_16565,N_17791);
nand U19319 (N_19319,N_17192,N_17039);
xor U19320 (N_19320,N_17425,N_17929);
nor U19321 (N_19321,N_16737,N_17157);
xnor U19322 (N_19322,N_17709,N_17053);
nand U19323 (N_19323,N_16501,N_17373);
nor U19324 (N_19324,N_17191,N_17958);
nor U19325 (N_19325,N_16939,N_17300);
nand U19326 (N_19326,N_17433,N_17991);
nor U19327 (N_19327,N_17380,N_17910);
and U19328 (N_19328,N_17057,N_17286);
nand U19329 (N_19329,N_17582,N_17243);
or U19330 (N_19330,N_17461,N_17942);
nor U19331 (N_19331,N_17316,N_17824);
xor U19332 (N_19332,N_17226,N_17254);
xor U19333 (N_19333,N_17091,N_16888);
or U19334 (N_19334,N_16999,N_17956);
or U19335 (N_19335,N_17022,N_17642);
nand U19336 (N_19336,N_16585,N_16945);
nor U19337 (N_19337,N_16661,N_16699);
or U19338 (N_19338,N_16978,N_17105);
or U19339 (N_19339,N_17149,N_17141);
or U19340 (N_19340,N_16879,N_16570);
and U19341 (N_19341,N_17585,N_17805);
and U19342 (N_19342,N_17341,N_17026);
nand U19343 (N_19343,N_17046,N_17259);
nand U19344 (N_19344,N_17746,N_17849);
nand U19345 (N_19345,N_17686,N_17493);
and U19346 (N_19346,N_17838,N_17373);
and U19347 (N_19347,N_16629,N_17891);
nor U19348 (N_19348,N_17320,N_17413);
xnor U19349 (N_19349,N_16612,N_16733);
xor U19350 (N_19350,N_17765,N_17338);
and U19351 (N_19351,N_17242,N_17889);
or U19352 (N_19352,N_17126,N_17688);
xnor U19353 (N_19353,N_17526,N_17825);
or U19354 (N_19354,N_17463,N_17336);
nand U19355 (N_19355,N_17036,N_17760);
nor U19356 (N_19356,N_17570,N_16561);
xor U19357 (N_19357,N_17122,N_16733);
nand U19358 (N_19358,N_17940,N_17145);
xor U19359 (N_19359,N_16659,N_17628);
xor U19360 (N_19360,N_17902,N_17577);
and U19361 (N_19361,N_17574,N_17942);
nand U19362 (N_19362,N_17736,N_17974);
nor U19363 (N_19363,N_16959,N_17610);
nor U19364 (N_19364,N_17779,N_17659);
nor U19365 (N_19365,N_16961,N_16845);
xnor U19366 (N_19366,N_17113,N_16981);
nand U19367 (N_19367,N_16615,N_17880);
nor U19368 (N_19368,N_16820,N_17735);
or U19369 (N_19369,N_16984,N_16844);
nand U19370 (N_19370,N_17495,N_17692);
nor U19371 (N_19371,N_17345,N_16747);
or U19372 (N_19372,N_17949,N_16963);
or U19373 (N_19373,N_17425,N_17877);
and U19374 (N_19374,N_17421,N_16807);
or U19375 (N_19375,N_17463,N_16990);
nor U19376 (N_19376,N_16568,N_16879);
and U19377 (N_19377,N_17606,N_17833);
nand U19378 (N_19378,N_16588,N_16786);
nor U19379 (N_19379,N_17081,N_17445);
xnor U19380 (N_19380,N_17931,N_17994);
or U19381 (N_19381,N_17914,N_17973);
or U19382 (N_19382,N_17529,N_17778);
or U19383 (N_19383,N_17141,N_16857);
or U19384 (N_19384,N_16706,N_16980);
nand U19385 (N_19385,N_17771,N_17851);
or U19386 (N_19386,N_17890,N_17355);
nand U19387 (N_19387,N_16593,N_16627);
or U19388 (N_19388,N_17260,N_17960);
xor U19389 (N_19389,N_17665,N_17583);
and U19390 (N_19390,N_17959,N_16677);
and U19391 (N_19391,N_17242,N_17548);
and U19392 (N_19392,N_16997,N_16505);
nor U19393 (N_19393,N_16536,N_17005);
xnor U19394 (N_19394,N_17892,N_16886);
nor U19395 (N_19395,N_16825,N_17642);
nand U19396 (N_19396,N_16501,N_16505);
nor U19397 (N_19397,N_17486,N_16795);
nand U19398 (N_19398,N_17186,N_17868);
and U19399 (N_19399,N_17972,N_17772);
nand U19400 (N_19400,N_16747,N_16799);
xor U19401 (N_19401,N_17560,N_17037);
nor U19402 (N_19402,N_17221,N_16500);
and U19403 (N_19403,N_16762,N_16953);
nand U19404 (N_19404,N_17742,N_17953);
and U19405 (N_19405,N_17741,N_17022);
or U19406 (N_19406,N_17735,N_17062);
xnor U19407 (N_19407,N_17218,N_17882);
or U19408 (N_19408,N_16623,N_17963);
and U19409 (N_19409,N_17670,N_17222);
or U19410 (N_19410,N_17896,N_17412);
xnor U19411 (N_19411,N_16700,N_16766);
and U19412 (N_19412,N_16518,N_17235);
nand U19413 (N_19413,N_17735,N_16502);
nor U19414 (N_19414,N_17411,N_16627);
nand U19415 (N_19415,N_17803,N_17543);
xor U19416 (N_19416,N_17402,N_17396);
nor U19417 (N_19417,N_17419,N_17877);
nor U19418 (N_19418,N_16783,N_17536);
xor U19419 (N_19419,N_17916,N_17773);
nor U19420 (N_19420,N_17462,N_17121);
or U19421 (N_19421,N_16805,N_16592);
nor U19422 (N_19422,N_17839,N_17022);
and U19423 (N_19423,N_17674,N_17256);
nand U19424 (N_19424,N_17993,N_17697);
and U19425 (N_19425,N_17751,N_17552);
nor U19426 (N_19426,N_17297,N_16516);
or U19427 (N_19427,N_16919,N_17339);
and U19428 (N_19428,N_17790,N_17581);
nand U19429 (N_19429,N_17206,N_17891);
or U19430 (N_19430,N_17880,N_17721);
nor U19431 (N_19431,N_17550,N_16533);
nor U19432 (N_19432,N_17789,N_16675);
nor U19433 (N_19433,N_17912,N_17221);
xnor U19434 (N_19434,N_16537,N_16811);
and U19435 (N_19435,N_17734,N_17488);
or U19436 (N_19436,N_17854,N_16606);
xnor U19437 (N_19437,N_17956,N_17039);
nor U19438 (N_19438,N_17286,N_17813);
and U19439 (N_19439,N_17421,N_17159);
and U19440 (N_19440,N_16624,N_16667);
nor U19441 (N_19441,N_17486,N_17979);
nand U19442 (N_19442,N_17957,N_16572);
nand U19443 (N_19443,N_17974,N_17211);
and U19444 (N_19444,N_16502,N_16589);
and U19445 (N_19445,N_17196,N_17318);
and U19446 (N_19446,N_16708,N_16566);
xnor U19447 (N_19447,N_17357,N_17046);
or U19448 (N_19448,N_16845,N_17589);
nand U19449 (N_19449,N_17772,N_16899);
and U19450 (N_19450,N_17373,N_17317);
and U19451 (N_19451,N_17514,N_17990);
and U19452 (N_19452,N_17244,N_16975);
nand U19453 (N_19453,N_16971,N_17375);
nand U19454 (N_19454,N_17481,N_17913);
or U19455 (N_19455,N_17991,N_17524);
or U19456 (N_19456,N_17984,N_16822);
nand U19457 (N_19457,N_16610,N_17644);
and U19458 (N_19458,N_16680,N_17838);
and U19459 (N_19459,N_16834,N_17944);
nor U19460 (N_19460,N_17053,N_17978);
nand U19461 (N_19461,N_17415,N_16609);
nor U19462 (N_19462,N_16907,N_16641);
or U19463 (N_19463,N_17900,N_17002);
nand U19464 (N_19464,N_17302,N_16545);
xnor U19465 (N_19465,N_16758,N_16862);
nor U19466 (N_19466,N_17341,N_17330);
xor U19467 (N_19467,N_17540,N_17174);
or U19468 (N_19468,N_17830,N_17411);
nor U19469 (N_19469,N_17786,N_16700);
nor U19470 (N_19470,N_16918,N_17476);
xor U19471 (N_19471,N_17961,N_16549);
or U19472 (N_19472,N_17557,N_16866);
nor U19473 (N_19473,N_17561,N_17293);
and U19474 (N_19474,N_17200,N_17918);
or U19475 (N_19475,N_17716,N_16776);
nand U19476 (N_19476,N_17260,N_16557);
and U19477 (N_19477,N_17836,N_17067);
nand U19478 (N_19478,N_17613,N_16711);
xor U19479 (N_19479,N_17882,N_17145);
nor U19480 (N_19480,N_17110,N_17328);
or U19481 (N_19481,N_16875,N_17916);
xor U19482 (N_19482,N_16823,N_16533);
nor U19483 (N_19483,N_17310,N_17793);
xnor U19484 (N_19484,N_16513,N_17483);
or U19485 (N_19485,N_16758,N_17111);
and U19486 (N_19486,N_16930,N_16901);
or U19487 (N_19487,N_17835,N_16886);
or U19488 (N_19488,N_17055,N_17709);
nand U19489 (N_19489,N_16905,N_17259);
and U19490 (N_19490,N_16630,N_17223);
xor U19491 (N_19491,N_17206,N_17551);
nand U19492 (N_19492,N_17173,N_17468);
and U19493 (N_19493,N_17232,N_17501);
nand U19494 (N_19494,N_16511,N_17848);
and U19495 (N_19495,N_16740,N_17546);
nand U19496 (N_19496,N_16797,N_16766);
or U19497 (N_19497,N_17253,N_17064);
nor U19498 (N_19498,N_17291,N_17812);
or U19499 (N_19499,N_17683,N_16631);
xor U19500 (N_19500,N_18139,N_18127);
or U19501 (N_19501,N_19131,N_18340);
nor U19502 (N_19502,N_18387,N_18291);
nand U19503 (N_19503,N_18839,N_18052);
xnor U19504 (N_19504,N_19300,N_19130);
and U19505 (N_19505,N_18475,N_18595);
nor U19506 (N_19506,N_18292,N_19105);
nor U19507 (N_19507,N_18159,N_18054);
xnor U19508 (N_19508,N_18241,N_18389);
or U19509 (N_19509,N_18437,N_18413);
or U19510 (N_19510,N_18145,N_19463);
nor U19511 (N_19511,N_19200,N_18277);
and U19512 (N_19512,N_18670,N_19398);
nor U19513 (N_19513,N_18360,N_18626);
and U19514 (N_19514,N_19447,N_18119);
or U19515 (N_19515,N_19012,N_19071);
or U19516 (N_19516,N_18644,N_18402);
and U19517 (N_19517,N_18819,N_18043);
nor U19518 (N_19518,N_18877,N_18947);
nor U19519 (N_19519,N_18272,N_18998);
and U19520 (N_19520,N_18608,N_19245);
xor U19521 (N_19521,N_19002,N_18632);
nor U19522 (N_19522,N_19124,N_19341);
xor U19523 (N_19523,N_18760,N_19191);
or U19524 (N_19524,N_18691,N_18612);
or U19525 (N_19525,N_18135,N_19125);
nor U19526 (N_19526,N_19466,N_18999);
nor U19527 (N_19527,N_18473,N_18955);
or U19528 (N_19528,N_18136,N_18414);
and U19529 (N_19529,N_18456,N_19255);
nand U19530 (N_19530,N_18216,N_19421);
and U19531 (N_19531,N_18111,N_18457);
and U19532 (N_19532,N_18311,N_19284);
nor U19533 (N_19533,N_18672,N_19244);
nor U19534 (N_19534,N_18396,N_18646);
and U19535 (N_19535,N_18502,N_19455);
or U19536 (N_19536,N_18912,N_18481);
nand U19537 (N_19537,N_18799,N_18783);
nor U19538 (N_19538,N_18914,N_18882);
and U19539 (N_19539,N_18883,N_19181);
nand U19540 (N_19540,N_18628,N_19231);
nand U19541 (N_19541,N_18880,N_18034);
xnor U19542 (N_19542,N_19456,N_19040);
or U19543 (N_19543,N_19265,N_19296);
and U19544 (N_19544,N_18070,N_19262);
nor U19545 (N_19545,N_18108,N_18723);
and U19546 (N_19546,N_19378,N_19415);
xor U19547 (N_19547,N_18784,N_18818);
or U19548 (N_19548,N_18341,N_18967);
and U19549 (N_19549,N_18253,N_18569);
xnor U19550 (N_19550,N_18012,N_18534);
or U19551 (N_19551,N_19473,N_18369);
nor U19552 (N_19552,N_18248,N_19392);
and U19553 (N_19553,N_19326,N_19268);
and U19554 (N_19554,N_18254,N_18333);
nor U19555 (N_19555,N_18422,N_19121);
and U19556 (N_19556,N_19331,N_18901);
and U19557 (N_19557,N_18150,N_19182);
nand U19558 (N_19558,N_18806,N_18170);
nand U19559 (N_19559,N_19008,N_18427);
nand U19560 (N_19560,N_18505,N_19282);
nand U19561 (N_19561,N_18313,N_19356);
nand U19562 (N_19562,N_18174,N_18721);
and U19563 (N_19563,N_18247,N_19285);
nand U19564 (N_19564,N_18220,N_18899);
and U19565 (N_19565,N_18500,N_18857);
nand U19566 (N_19566,N_19113,N_18467);
and U19567 (N_19567,N_18939,N_18529);
nand U19568 (N_19568,N_18197,N_18666);
xor U19569 (N_19569,N_19276,N_18526);
or U19570 (N_19570,N_19229,N_19334);
and U19571 (N_19571,N_18546,N_19007);
or U19572 (N_19572,N_18168,N_19153);
or U19573 (N_19573,N_18759,N_18874);
xor U19574 (N_19574,N_18544,N_19361);
and U19575 (N_19575,N_18162,N_19114);
nor U19576 (N_19576,N_19027,N_18611);
or U19577 (N_19577,N_18614,N_18957);
and U19578 (N_19578,N_19011,N_19358);
xnor U19579 (N_19579,N_18297,N_19157);
nor U19580 (N_19580,N_19496,N_18488);
nand U19581 (N_19581,N_18461,N_19189);
xnor U19582 (N_19582,N_18550,N_18978);
nand U19583 (N_19583,N_19050,N_18657);
nand U19584 (N_19584,N_18075,N_18835);
xnor U19585 (N_19585,N_18349,N_19281);
or U19586 (N_19586,N_18903,N_19333);
nand U19587 (N_19587,N_19150,N_18645);
nand U19588 (N_19588,N_18689,N_18151);
xnor U19589 (N_19589,N_19492,N_18714);
nand U19590 (N_19590,N_18794,N_18167);
or U19591 (N_19591,N_19485,N_19257);
xor U19592 (N_19592,N_18142,N_19058);
nor U19593 (N_19593,N_18838,N_18524);
nor U19594 (N_19594,N_18562,N_18022);
nand U19595 (N_19595,N_19236,N_18979);
nor U19596 (N_19596,N_18528,N_19348);
or U19597 (N_19597,N_18179,N_19029);
or U19598 (N_19598,N_18682,N_18314);
nor U19599 (N_19599,N_19448,N_18153);
and U19600 (N_19600,N_19070,N_18660);
xor U19601 (N_19601,N_18042,N_18888);
nor U19602 (N_19602,N_18002,N_18105);
xor U19603 (N_19603,N_18324,N_19039);
xor U19604 (N_19604,N_19472,N_18728);
or U19605 (N_19605,N_19446,N_19064);
nand U19606 (N_19606,N_18989,N_19406);
nand U19607 (N_19607,N_19022,N_18594);
and U19608 (N_19608,N_19045,N_19230);
nand U19609 (N_19609,N_19468,N_18952);
nand U19610 (N_19610,N_18230,N_18286);
xnor U19611 (N_19611,N_18050,N_18563);
nor U19612 (N_19612,N_18305,N_18264);
xnor U19613 (N_19613,N_19283,N_19261);
nor U19614 (N_19614,N_18683,N_19490);
or U19615 (N_19615,N_18918,N_18451);
nor U19616 (N_19616,N_18603,N_19227);
nor U19617 (N_19617,N_19266,N_18121);
and U19618 (N_19618,N_18074,N_18557);
and U19619 (N_19619,N_19216,N_19397);
nand U19620 (N_19620,N_18859,N_19219);
or U19621 (N_19621,N_19287,N_18803);
nor U19622 (N_19622,N_18251,N_18605);
nor U19623 (N_19623,N_18749,N_19366);
and U19624 (N_19624,N_18586,N_18415);
and U19625 (N_19625,N_19461,N_18056);
nand U19626 (N_19626,N_19363,N_18356);
nand U19627 (N_19627,N_18889,N_19400);
nor U19628 (N_19628,N_19053,N_18726);
nor U19629 (N_19629,N_19217,N_19260);
nand U19630 (N_19630,N_18780,N_18099);
and U19631 (N_19631,N_18280,N_19430);
nand U19632 (N_19632,N_19162,N_18198);
and U19633 (N_19633,N_18719,N_19041);
xnor U19634 (N_19634,N_19116,N_18161);
nand U19635 (N_19635,N_18897,N_18945);
and U19636 (N_19636,N_18828,N_19493);
nand U19637 (N_19637,N_18057,N_18982);
xor U19638 (N_19638,N_18662,N_19005);
nor U19639 (N_19639,N_18848,N_19286);
and U19640 (N_19640,N_18941,N_18447);
nor U19641 (N_19641,N_18066,N_18188);
or U19642 (N_19642,N_19313,N_19028);
xnor U19643 (N_19643,N_18047,N_18981);
and U19644 (N_19644,N_18064,N_18375);
and U19645 (N_19645,N_18191,N_19422);
or U19646 (N_19646,N_18992,N_19183);
xnor U19647 (N_19647,N_19104,N_18116);
or U19648 (N_19648,N_18364,N_18143);
xnor U19649 (N_19649,N_18570,N_18008);
nand U19650 (N_19650,N_18186,N_18913);
nor U19651 (N_19651,N_19478,N_18568);
nor U19652 (N_19652,N_18745,N_18246);
nand U19653 (N_19653,N_18923,N_18373);
and U19654 (N_19654,N_18394,N_18959);
xor U19655 (N_19655,N_18746,N_19139);
xnor U19656 (N_19656,N_18559,N_18538);
and U19657 (N_19657,N_18433,N_19140);
xor U19658 (N_19658,N_19156,N_18625);
nand U19659 (N_19659,N_19166,N_18518);
nor U19660 (N_19660,N_18958,N_18752);
and U19661 (N_19661,N_18761,N_18685);
nand U19662 (N_19662,N_18814,N_18381);
xor U19663 (N_19663,N_19048,N_18450);
or U19664 (N_19664,N_18269,N_18576);
and U19665 (N_19665,N_18738,N_18748);
nand U19666 (N_19666,N_18440,N_19207);
xnor U19667 (N_19667,N_18206,N_18204);
xnor U19668 (N_19668,N_19375,N_18320);
nor U19669 (N_19669,N_18511,N_18896);
nand U19670 (N_19670,N_18675,N_19129);
nor U19671 (N_19671,N_19147,N_18987);
nand U19672 (N_19672,N_18776,N_18290);
nor U19673 (N_19673,N_18696,N_18462);
nand U19674 (N_19674,N_19381,N_18885);
nand U19675 (N_19675,N_18325,N_18395);
or U19676 (N_19676,N_18956,N_18160);
xnor U19677 (N_19677,N_18508,N_19454);
nand U19678 (N_19678,N_18589,N_18668);
and U19679 (N_19679,N_18434,N_18652);
nor U19680 (N_19680,N_19362,N_18367);
nand U19681 (N_19681,N_18868,N_18821);
nand U19682 (N_19682,N_19187,N_19495);
xnor U19683 (N_19683,N_18149,N_18969);
xnor U19684 (N_19684,N_18489,N_18671);
nand U19685 (N_19685,N_19347,N_18736);
nand U19686 (N_19686,N_18937,N_18503);
nor U19687 (N_19687,N_18287,N_19310);
or U19688 (N_19688,N_18943,N_18622);
nand U19689 (N_19689,N_18083,N_19003);
and U19690 (N_19690,N_18158,N_18322);
or U19691 (N_19691,N_19394,N_18577);
nand U19692 (N_19692,N_18499,N_19133);
nand U19693 (N_19693,N_18732,N_18243);
nand U19694 (N_19694,N_19437,N_19094);
nor U19695 (N_19695,N_18970,N_18062);
and U19696 (N_19696,N_18497,N_19367);
or U19697 (N_19697,N_18094,N_18906);
nor U19698 (N_19698,N_18676,N_18275);
nand U19699 (N_19699,N_18229,N_18922);
and U19700 (N_19700,N_18713,N_19371);
or U19701 (N_19701,N_19308,N_18667);
and U19702 (N_19702,N_18853,N_18861);
or U19703 (N_19703,N_18694,N_19431);
xnor U19704 (N_19704,N_18417,N_18968);
xnor U19705 (N_19705,N_18664,N_18237);
nand U19706 (N_19706,N_18695,N_18207);
nand U19707 (N_19707,N_18040,N_18658);
nor U19708 (N_19708,N_18480,N_19086);
nor U19709 (N_19709,N_19004,N_18974);
nor U19710 (N_19710,N_19383,N_19254);
nand U19711 (N_19711,N_19401,N_18282);
xnor U19712 (N_19712,N_18581,N_18638);
or U19713 (N_19713,N_18724,N_19192);
or U19714 (N_19714,N_18444,N_19360);
and U19715 (N_19715,N_19160,N_19270);
nor U19716 (N_19716,N_18900,N_18512);
and U19717 (N_19717,N_19359,N_19280);
xnor U19718 (N_19718,N_19080,N_18084);
nand U19719 (N_19719,N_18323,N_18832);
or U19720 (N_19720,N_18257,N_18798);
nand U19721 (N_19721,N_18718,N_18202);
nor U19722 (N_19722,N_18984,N_18063);
nand U19723 (N_19723,N_19251,N_18080);
or U19724 (N_19724,N_18453,N_18782);
nor U19725 (N_19725,N_19488,N_18009);
nor U19726 (N_19726,N_19423,N_18400);
nor U19727 (N_19727,N_18565,N_19142);
nor U19728 (N_19728,N_18802,N_18843);
and U19729 (N_19729,N_18887,N_18796);
nor U19730 (N_19730,N_18750,N_18081);
xnor U19731 (N_19731,N_18866,N_18583);
xor U19732 (N_19732,N_18673,N_18331);
nand U19733 (N_19733,N_19317,N_19253);
xor U19734 (N_19734,N_18860,N_18114);
nand U19735 (N_19735,N_18102,N_18684);
nor U19736 (N_19736,N_18483,N_18731);
xor U19737 (N_19737,N_18758,N_19418);
or U19738 (N_19738,N_18920,N_18881);
nor U19739 (N_19739,N_18602,N_18370);
and U19740 (N_19740,N_19049,N_19063);
or U19741 (N_19741,N_18132,N_18771);
nand U19742 (N_19742,N_18397,N_18013);
xnor U19743 (N_19743,N_18869,N_19225);
and U19744 (N_19744,N_19357,N_18215);
xnor U19745 (N_19745,N_19190,N_18884);
xnor U19746 (N_19746,N_18729,N_18836);
nor U19747 (N_19747,N_18635,N_18663);
or U19748 (N_19748,N_18426,N_19099);
nor U19749 (N_19749,N_19117,N_18606);
nor U19750 (N_19750,N_18045,N_18232);
or U19751 (N_19751,N_18107,N_18295);
xnor U19752 (N_19752,N_18101,N_19148);
and U19753 (N_19753,N_19194,N_19228);
or U19754 (N_19754,N_18651,N_18337);
and U19755 (N_19755,N_18078,N_18768);
and U19756 (N_19756,N_18338,N_18224);
nand U19757 (N_19757,N_19293,N_18312);
xnor U19758 (N_19758,N_19449,N_19241);
and U19759 (N_19759,N_19055,N_18353);
nand U19760 (N_19760,N_18332,N_18643);
nor U19761 (N_19761,N_18919,N_19471);
nor U19762 (N_19762,N_18449,N_18309);
and U19763 (N_19763,N_18140,N_18468);
xnor U19764 (N_19764,N_18790,N_18712);
or U19765 (N_19765,N_19327,N_18983);
or U19766 (N_19766,N_18196,N_19209);
and U19767 (N_19767,N_18756,N_19025);
or U19768 (N_19768,N_18739,N_19032);
xor U19769 (N_19769,N_19416,N_18580);
xor U19770 (N_19770,N_18770,N_18376);
or U19771 (N_19771,N_19391,N_19035);
nand U19772 (N_19772,N_18878,N_18575);
xor U19773 (N_19773,N_18574,N_18420);
xnor U19774 (N_19774,N_18687,N_18813);
xnor U19775 (N_19775,N_19299,N_18495);
or U19776 (N_19776,N_18787,N_19298);
or U19777 (N_19777,N_18199,N_19073);
or U19778 (N_19778,N_18924,N_19062);
xnor U19779 (N_19779,N_18330,N_19453);
nor U19780 (N_19780,N_18408,N_18030);
nor U19781 (N_19781,N_18824,N_18742);
or U19782 (N_19782,N_18743,N_19204);
xor U19783 (N_19783,N_18192,N_18767);
nor U19784 (N_19784,N_18410,N_18104);
xnor U19785 (N_19785,N_18391,N_19015);
nor U19786 (N_19786,N_19373,N_18496);
xor U19787 (N_19787,N_18699,N_18336);
and U19788 (N_19788,N_18454,N_19179);
and U19789 (N_19789,N_19097,N_18035);
nand U19790 (N_19790,N_19013,N_18300);
nand U19791 (N_19791,N_19009,N_19354);
xnor U19792 (N_19792,N_18515,N_19295);
or U19793 (N_19793,N_19470,N_19305);
or U19794 (N_19794,N_19405,N_19374);
xnor U19795 (N_19795,N_18339,N_19324);
nor U19796 (N_19796,N_19314,N_18374);
or U19797 (N_19797,N_19078,N_19339);
xor U19798 (N_19798,N_18905,N_18494);
nor U19799 (N_19799,N_19038,N_18227);
and U19800 (N_19800,N_19123,N_19384);
nand U19801 (N_19801,N_19088,N_18807);
and U19802 (N_19802,N_18165,N_18704);
xnor U19803 (N_19803,N_18407,N_19091);
nor U19804 (N_19804,N_19108,N_18472);
and U19805 (N_19805,N_19074,N_18044);
nor U19806 (N_19806,N_18458,N_18334);
nand U19807 (N_19807,N_18553,N_18004);
or U19808 (N_19808,N_18128,N_18561);
nand U19809 (N_19809,N_19294,N_19102);
nor U19810 (N_19810,N_18328,N_18686);
and U19811 (N_19811,N_18182,N_18223);
or U19812 (N_19812,N_19076,N_18329);
xnor U19813 (N_19813,N_18493,N_18266);
nand U19814 (N_19814,N_18171,N_18637);
nor U19815 (N_19815,N_18741,N_18717);
nand U19816 (N_19816,N_19315,N_18636);
and U19817 (N_19817,N_18365,N_18973);
or U19818 (N_19818,N_18697,N_18304);
or U19819 (N_19819,N_18560,N_19480);
nand U19820 (N_19820,N_18951,N_19306);
nor U19821 (N_19821,N_18399,N_18928);
nor U19822 (N_19822,N_19047,N_18392);
or U19823 (N_19823,N_19438,N_18079);
nor U19824 (N_19824,N_19177,N_18733);
nor U19825 (N_19825,N_18210,N_18624);
xnor U19826 (N_19826,N_19134,N_18307);
xor U19827 (N_19827,N_18558,N_19250);
xor U19828 (N_19828,N_19126,N_19174);
or U19829 (N_19829,N_18347,N_18477);
nand U19830 (N_19830,N_18384,N_19467);
xor U19831 (N_19831,N_19095,N_18792);
nor U19832 (N_19832,N_19020,N_18778);
and U19833 (N_19833,N_18962,N_19197);
xor U19834 (N_19834,N_19389,N_18566);
nor U19835 (N_19835,N_18532,N_19386);
and U19836 (N_19836,N_18418,N_19399);
nand U19837 (N_19837,N_18706,N_18431);
nand U19838 (N_19838,N_19138,N_18630);
or U19839 (N_19839,N_19309,N_18772);
nand U19840 (N_19840,N_18716,N_18036);
and U19841 (N_19841,N_18465,N_19424);
nand U19842 (N_19842,N_18476,N_19412);
nand U19843 (N_19843,N_18598,N_18487);
nor U19844 (N_19844,N_18910,N_19272);
nand U19845 (N_19845,N_19106,N_18006);
or U19846 (N_19846,N_18255,N_18705);
or U19847 (N_19847,N_19052,N_18299);
and U19848 (N_19848,N_19497,N_19291);
and U19849 (N_19849,N_18076,N_19042);
xor U19850 (N_19850,N_19462,N_18540);
nor U19851 (N_19851,N_18423,N_18362);
or U19852 (N_19852,N_19180,N_19165);
nor U19853 (N_19853,N_18707,N_18944);
or U19854 (N_19854,N_18527,N_18293);
and U19855 (N_19855,N_18350,N_18517);
and U19856 (N_19856,N_18734,N_18591);
or U19857 (N_19857,N_18484,N_19376);
nand U19858 (N_19858,N_18491,N_18091);
or U19859 (N_19859,N_18001,N_19110);
nor U19860 (N_19860,N_19345,N_18530);
and U19861 (N_19861,N_19232,N_18619);
or U19862 (N_19862,N_19170,N_18366);
or U19863 (N_19863,N_19425,N_18985);
and U19864 (N_19864,N_18514,N_19368);
or U19865 (N_19865,N_18014,N_19037);
nand U19866 (N_19866,N_18823,N_18930);
or U19867 (N_19867,N_18003,N_18106);
nand U19868 (N_19868,N_19171,N_18708);
nand U19869 (N_19869,N_18157,N_19036);
nor U19870 (N_19870,N_19030,N_18909);
nor U19871 (N_19871,N_18634,N_19441);
and U19872 (N_19872,N_19172,N_18296);
nor U19873 (N_19873,N_19067,N_19307);
and U19874 (N_19874,N_19328,N_19304);
xor U19875 (N_19875,N_18315,N_18436);
or U19876 (N_19876,N_18873,N_18520);
nand U19877 (N_19877,N_18181,N_19079);
xnor U19878 (N_19878,N_18601,N_18507);
or U19879 (N_19879,N_19185,N_18986);
xor U19880 (N_19880,N_19066,N_18302);
and U19881 (N_19881,N_18267,N_19290);
nor U19882 (N_19882,N_18816,N_18378);
nand U19883 (N_19883,N_19264,N_18765);
nor U19884 (N_19884,N_18963,N_18876);
xor U19885 (N_19885,N_18343,N_18949);
nor U19886 (N_19886,N_19206,N_18425);
xnor U19887 (N_19887,N_18800,N_18825);
nor U19888 (N_19888,N_18361,N_19082);
and U19889 (N_19889,N_18274,N_18131);
xor U19890 (N_19890,N_18478,N_18310);
and U19891 (N_19891,N_18991,N_18582);
nand U19892 (N_19892,N_19319,N_18797);
or U19893 (N_19893,N_18112,N_18972);
nand U19894 (N_19894,N_18674,N_18442);
nor U19895 (N_19895,N_18964,N_19024);
nor U19896 (N_19896,N_18805,N_19128);
xnor U19897 (N_19897,N_19323,N_18416);
xor U19898 (N_19898,N_18163,N_18256);
nand U19899 (N_19899,N_19210,N_18096);
xnor U19900 (N_19900,N_19335,N_18217);
or U19901 (N_19901,N_18845,N_18954);
nor U19902 (N_19902,N_18189,N_18482);
or U19903 (N_19903,N_18085,N_18259);
and U19904 (N_19904,N_19426,N_18005);
nor U19905 (N_19905,N_18863,N_19469);
or U19906 (N_19906,N_18579,N_19479);
or U19907 (N_19907,N_18086,N_18895);
xnor U19908 (N_19908,N_18966,N_18915);
nand U19909 (N_19909,N_18020,N_18109);
and U19910 (N_19910,N_19188,N_18156);
nor U19911 (N_19911,N_19457,N_18463);
xnor U19912 (N_19912,N_18089,N_18543);
xnor U19913 (N_19913,N_19407,N_18211);
nor U19914 (N_19914,N_18278,N_18234);
xnor U19915 (N_19915,N_18406,N_18051);
xor U19916 (N_19916,N_18097,N_18424);
xor U19917 (N_19917,N_18698,N_18766);
or U19918 (N_19918,N_19084,N_18235);
or U19919 (N_19919,N_18026,N_18355);
or U19920 (N_19920,N_19444,N_19195);
nor U19921 (N_19921,N_18975,N_18940);
xor U19922 (N_19922,N_18735,N_18169);
or U19923 (N_19923,N_19202,N_18231);
xnor U19924 (N_19924,N_19186,N_19278);
or U19925 (N_19925,N_18931,N_19234);
nor U19926 (N_19926,N_18572,N_18715);
xor U19927 (N_19927,N_18492,N_19018);
and U19928 (N_19928,N_18093,N_19031);
xnor U19929 (N_19929,N_18599,N_18617);
nor U19930 (N_19930,N_19215,N_18757);
xnor U19931 (N_19931,N_19152,N_18471);
and U19932 (N_19932,N_18501,N_18172);
and U19933 (N_19933,N_18438,N_19096);
nor U19934 (N_19934,N_18710,N_19487);
nor U19935 (N_19935,N_18240,N_19111);
xnor U19936 (N_19936,N_19451,N_18830);
and U19937 (N_19937,N_18808,N_18409);
nand U19938 (N_19938,N_18702,N_18804);
and U19939 (N_19939,N_18867,N_18180);
or U19940 (N_19940,N_19297,N_18455);
or U19941 (N_19941,N_18125,N_18037);
nand U19942 (N_19942,N_19435,N_18545);
xnor U19943 (N_19943,N_18864,N_19379);
nor U19944 (N_19944,N_18849,N_19213);
and U19945 (N_19945,N_18464,N_18639);
or U19946 (N_19946,N_18996,N_19077);
nor U19947 (N_19947,N_19273,N_18610);
xor U19948 (N_19948,N_18469,N_18994);
nor U19949 (N_19949,N_18024,N_18072);
or U19950 (N_19950,N_19043,N_19087);
nand U19951 (N_19951,N_19151,N_18031);
nor U19952 (N_19952,N_18398,N_18788);
nand U19953 (N_19953,N_18067,N_18316);
nor U19954 (N_19954,N_18841,N_19101);
nor U19955 (N_19955,N_18680,N_19365);
nand U19956 (N_19956,N_18011,N_19271);
nor U19957 (N_19957,N_19289,N_18692);
nor U19958 (N_19958,N_18911,N_18276);
xor U19959 (N_19959,N_18669,N_19198);
or U19960 (N_19960,N_18175,N_19267);
nand U19961 (N_19961,N_19396,N_19075);
xnor U19962 (N_19962,N_18856,N_18294);
xnor U19963 (N_19963,N_19411,N_19127);
and U19964 (N_19964,N_18460,N_19006);
nand U19965 (N_19965,N_18926,N_18510);
xor U19966 (N_19966,N_18934,N_19342);
nand U19967 (N_19967,N_18596,N_18907);
or U19968 (N_19968,N_18352,N_19176);
and U19969 (N_19969,N_19428,N_19060);
nand U19970 (N_19970,N_19499,N_18871);
xor U19971 (N_19971,N_18590,N_19023);
nand U19972 (N_19972,N_18513,N_18221);
and U19973 (N_19973,N_19175,N_19145);
nand U19974 (N_19974,N_18242,N_18597);
xnor U19975 (N_19975,N_18244,N_18100);
or U19976 (N_19976,N_19352,N_18661);
and U19977 (N_19977,N_19442,N_18722);
xnor U19978 (N_19978,N_18383,N_18000);
nand U19979 (N_19979,N_18592,N_18516);
nand U19980 (N_19980,N_18405,N_19021);
xor U19981 (N_19981,N_18890,N_18725);
nand U19982 (N_19982,N_19222,N_19311);
nand U19983 (N_19983,N_18842,N_18164);
or U19984 (N_19984,N_18155,N_18386);
nor U19985 (N_19985,N_19256,N_18764);
and U19986 (N_19986,N_19051,N_18212);
or U19987 (N_19987,N_18303,N_18306);
and U19988 (N_19988,N_18146,N_19247);
or U19989 (N_19989,N_19380,N_18811);
xor U19990 (N_19990,N_18653,N_18858);
nand U19991 (N_19991,N_18781,N_18138);
and U19992 (N_19992,N_18088,N_19318);
nand U19993 (N_19993,N_18401,N_18372);
nor U19994 (N_19994,N_18377,N_18017);
nand U19995 (N_19995,N_19409,N_18194);
and U19996 (N_19996,N_18065,N_19385);
or U19997 (N_19997,N_19427,N_18609);
and U19998 (N_19998,N_18298,N_18284);
or U19999 (N_19999,N_18879,N_19489);
and U20000 (N_20000,N_18380,N_19477);
xor U20001 (N_20001,N_19034,N_18809);
and U20002 (N_20002,N_19016,N_19211);
xor U20003 (N_20003,N_18466,N_19010);
xor U20004 (N_20004,N_19393,N_18435);
or U20005 (N_20005,N_18388,N_18137);
or U20006 (N_20006,N_19118,N_19303);
and U20007 (N_20007,N_18321,N_18200);
nor U20008 (N_20008,N_18118,N_18317);
xnor U20009 (N_20009,N_18822,N_19372);
or U20010 (N_20010,N_18659,N_19321);
nor U20011 (N_20011,N_19208,N_19388);
and U20012 (N_20012,N_19445,N_18419);
nor U20013 (N_20013,N_18775,N_19173);
and U20014 (N_20014,N_18411,N_18263);
nand U20015 (N_20015,N_18587,N_18834);
or U20016 (N_20016,N_18486,N_18046);
xnor U20017 (N_20017,N_19103,N_19235);
nor U20018 (N_20018,N_19237,N_18938);
and U20019 (N_20019,N_19056,N_18631);
or U20020 (N_20020,N_18007,N_19404);
xor U20021 (N_20021,N_18519,N_18023);
and U20022 (N_20022,N_18700,N_18203);
or U20023 (N_20023,N_19269,N_18936);
nor U20024 (N_20024,N_18833,N_18016);
and U20025 (N_20025,N_19349,N_19484);
xor U20026 (N_20026,N_18327,N_19223);
xor U20027 (N_20027,N_18359,N_19112);
and U20028 (N_20028,N_18829,N_18850);
nor U20029 (N_20029,N_18567,N_18875);
nor U20030 (N_20030,N_18893,N_18649);
nand U20031 (N_20031,N_19212,N_19414);
nor U20032 (N_20032,N_19122,N_19350);
and U20033 (N_20033,N_18548,N_18665);
xor U20034 (N_20034,N_18837,N_18640);
xnor U20035 (N_20035,N_18785,N_19100);
nand U20036 (N_20036,N_19238,N_19370);
nor U20037 (N_20037,N_18921,N_18193);
or U20038 (N_20038,N_19252,N_19410);
and U20039 (N_20039,N_18747,N_18218);
xor U20040 (N_20040,N_19459,N_18647);
xnor U20041 (N_20041,N_18678,N_18260);
nor U20042 (N_20042,N_19109,N_19141);
nand U20043 (N_20043,N_18351,N_18412);
and U20044 (N_20044,N_18642,N_18953);
and U20045 (N_20045,N_19220,N_18249);
nor U20046 (N_20046,N_18618,N_19144);
xor U20047 (N_20047,N_18285,N_18820);
and U20048 (N_20048,N_18977,N_18531);
nand U20049 (N_20049,N_18048,N_18059);
nand U20050 (N_20050,N_18092,N_19336);
or U20051 (N_20051,N_19143,N_18152);
or U20052 (N_20052,N_19169,N_18250);
nor U20053 (N_20053,N_18993,N_19377);
nand U20054 (N_20054,N_18219,N_18961);
xor U20055 (N_20055,N_19119,N_19155);
nor U20056 (N_20056,N_19301,N_18069);
nor U20057 (N_20057,N_18301,N_19498);
nand U20058 (N_20058,N_19403,N_18916);
or U20059 (N_20059,N_18855,N_18021);
nor U20060 (N_20060,N_18509,N_19292);
nand U20061 (N_20061,N_18600,N_18268);
nand U20062 (N_20062,N_18041,N_19243);
or U20063 (N_20063,N_19093,N_18073);
nand U20064 (N_20064,N_18273,N_18363);
or U20065 (N_20065,N_18535,N_18061);
or U20066 (N_20066,N_18432,N_18225);
or U20067 (N_20067,N_18846,N_19044);
nand U20068 (N_20068,N_19054,N_18270);
or U20069 (N_20069,N_19316,N_18862);
or U20070 (N_20070,N_18459,N_19464);
xor U20071 (N_20071,N_19017,N_19387);
or U20072 (N_20072,N_18178,N_18446);
xor U20073 (N_20073,N_19344,N_18988);
or U20074 (N_20074,N_18345,N_18010);
or U20075 (N_20075,N_19115,N_18620);
and U20076 (N_20076,N_18727,N_19248);
or U20077 (N_20077,N_18390,N_18154);
or U20078 (N_20078,N_18892,N_18870);
nor U20079 (N_20079,N_18245,N_19098);
nand U20080 (N_20080,N_18421,N_18690);
nor U20081 (N_20081,N_18448,N_18942);
xor U20082 (N_20082,N_18443,N_19137);
or U20083 (N_20083,N_19475,N_18786);
and U20084 (N_20084,N_18655,N_19439);
nand U20085 (N_20085,N_18932,N_19458);
or U20086 (N_20086,N_18498,N_18965);
xor U20087 (N_20087,N_18755,N_18549);
nor U20088 (N_20088,N_18522,N_18288);
nor U20089 (N_20089,N_18654,N_18585);
nand U20090 (N_20090,N_19436,N_18904);
and U20091 (N_20091,N_18055,N_19178);
or U20092 (N_20092,N_18439,N_19332);
nand U20093 (N_20093,N_19199,N_19242);
or U20094 (N_20094,N_18371,N_18898);
nor U20095 (N_20095,N_19081,N_18238);
and U20096 (N_20096,N_18971,N_19072);
nor U20097 (N_20097,N_18817,N_18555);
or U20098 (N_20098,N_19205,N_18087);
xnor U20099 (N_20099,N_19274,N_18613);
and U20100 (N_20100,N_19136,N_19146);
nor U20101 (N_20101,N_18265,N_18851);
nand U20102 (N_20102,N_18205,N_18744);
nand U20103 (N_20103,N_18917,N_18688);
and U20104 (N_20104,N_18925,N_18847);
or U20105 (N_20105,N_19068,N_18902);
and U20106 (N_20106,N_18474,N_19408);
or U20107 (N_20107,N_19083,N_18740);
and U20108 (N_20108,N_18504,N_18679);
or U20109 (N_20109,N_18536,N_19330);
or U20110 (N_20110,N_18990,N_19059);
or U20111 (N_20111,N_18404,N_18049);
or U20112 (N_20112,N_18604,N_19014);
xnor U20113 (N_20113,N_18701,N_18382);
xor U20114 (N_20114,N_18252,N_19355);
nor U20115 (N_20115,N_18441,N_18730);
and U20116 (N_20116,N_18616,N_18946);
and U20117 (N_20117,N_19249,N_18720);
xor U20118 (N_20118,N_18428,N_18346);
or U20119 (N_20119,N_18815,N_19450);
or U20120 (N_20120,N_18533,N_18348);
nor U20121 (N_20121,N_18623,N_19218);
nand U20122 (N_20122,N_18261,N_18827);
xnor U20123 (N_20123,N_18190,N_19486);
nand U20124 (N_20124,N_19483,N_18693);
nand U20125 (N_20125,N_18490,N_18826);
or U20126 (N_20126,N_19279,N_19364);
xnor U20127 (N_20127,N_18077,N_18648);
nor U20128 (N_20128,N_19033,N_18239);
nor U20129 (N_20129,N_18038,N_18429);
and U20130 (N_20130,N_18886,N_18393);
nand U20131 (N_20131,N_19069,N_19168);
nand U20132 (N_20132,N_19320,N_18703);
and U20133 (N_20133,N_18523,N_18854);
xnor U20134 (N_20134,N_18681,N_19322);
xnor U20135 (N_20135,N_19346,N_18222);
nor U20136 (N_20136,N_19090,N_19258);
xnor U20137 (N_20137,N_18929,N_19000);
or U20138 (N_20138,N_19026,N_19132);
nor U20139 (N_20139,N_18506,N_18865);
nand U20140 (N_20140,N_18584,N_18058);
or U20141 (N_20141,N_19149,N_18115);
or U20142 (N_20142,N_19221,N_18015);
nor U20143 (N_20143,N_18053,N_19201);
xor U20144 (N_20144,N_19233,N_18777);
xnor U20145 (N_20145,N_18126,N_18271);
nor U20146 (N_20146,N_18995,N_19164);
nand U20147 (N_20147,N_18027,N_19351);
nor U20148 (N_20148,N_18556,N_18831);
and U20149 (N_20149,N_19154,N_18793);
nand U20150 (N_20150,N_19288,N_18185);
and U20151 (N_20151,N_18209,N_19491);
or U20152 (N_20152,N_18289,N_19061);
nor U20153 (N_20153,N_18120,N_19413);
and U20154 (N_20154,N_18773,N_18751);
xor U20155 (N_20155,N_18891,N_18445);
or U20156 (N_20156,N_19353,N_18573);
nand U20157 (N_20157,N_19390,N_18166);
xnor U20158 (N_20158,N_18173,N_18354);
nor U20159 (N_20159,N_18633,N_19433);
or U20160 (N_20160,N_18228,N_19302);
nor U20161 (N_20161,N_18233,N_18033);
xnor U20162 (N_20162,N_19312,N_18812);
nand U20163 (N_20163,N_18711,N_18213);
nor U20164 (N_20164,N_18090,N_19057);
xnor U20165 (N_20165,N_18539,N_19046);
nor U20166 (N_20166,N_18769,N_18113);
xnor U20167 (N_20167,N_19434,N_18187);
or U20168 (N_20168,N_19135,N_18148);
xor U20169 (N_20169,N_18385,N_18184);
nand U20170 (N_20170,N_18547,N_19246);
or U20171 (N_20171,N_18129,N_18130);
and U20172 (N_20172,N_18578,N_18335);
or U20173 (N_20173,N_18629,N_18357);
and U20174 (N_20174,N_18763,N_19474);
and U20175 (N_20175,N_18095,N_18779);
and U20176 (N_20176,N_18344,N_18283);
nand U20177 (N_20177,N_19338,N_18927);
and U20178 (N_20178,N_19167,N_19440);
and U20179 (N_20179,N_18872,N_18403);
or U20180 (N_20180,N_18933,N_18122);
nor U20181 (N_20181,N_18552,N_18110);
nor U20182 (N_20182,N_19214,N_19259);
nand U20183 (N_20183,N_19417,N_18258);
nor U20184 (N_20184,N_18039,N_18028);
nor U20185 (N_20185,N_19452,N_18279);
and U20186 (N_20186,N_18607,N_18791);
and U20187 (N_20187,N_19158,N_19482);
or U20188 (N_20188,N_18656,N_18542);
or U20189 (N_20189,N_18358,N_18281);
nor U20190 (N_20190,N_19107,N_19240);
nand U20191 (N_20191,N_19277,N_18019);
nand U20192 (N_20192,N_18123,N_18318);
nor U20193 (N_20193,N_19239,N_18935);
and U20194 (N_20194,N_18852,N_18521);
or U20195 (N_20195,N_18103,N_19460);
or U20196 (N_20196,N_19402,N_19226);
or U20197 (N_20197,N_19325,N_18226);
or U20198 (N_20198,N_18144,N_18479);
nand U20199 (N_20199,N_18709,N_18997);
nand U20200 (N_20200,N_18525,N_18147);
nand U20201 (N_20201,N_19019,N_19161);
nor U20202 (N_20202,N_19369,N_19275);
nor U20203 (N_20203,N_19382,N_19193);
xnor U20204 (N_20204,N_18071,N_19343);
xor U20205 (N_20205,N_18134,N_18236);
xnor U20206 (N_20206,N_18554,N_18018);
or U20207 (N_20207,N_18032,N_18262);
xor U20208 (N_20208,N_19196,N_18208);
nand U20209 (N_20209,N_18621,N_18762);
or U20210 (N_20210,N_18541,N_19224);
nand U20211 (N_20211,N_18588,N_18980);
nand U20212 (N_20212,N_19184,N_18840);
or U20213 (N_20213,N_19089,N_18342);
and U20214 (N_20214,N_19443,N_18117);
nor U20215 (N_20215,N_18641,N_19419);
and U20216 (N_20216,N_18737,N_18177);
nor U20217 (N_20217,N_18124,N_18537);
nand U20218 (N_20218,N_18029,N_19420);
or U20219 (N_20219,N_18308,N_18948);
xnor U20220 (N_20220,N_18753,N_18801);
nor U20221 (N_20221,N_19001,N_18183);
nand U20222 (N_20222,N_19429,N_18795);
and U20223 (N_20223,N_18810,N_18571);
nor U20224 (N_20224,N_18201,N_19340);
nor U20225 (N_20225,N_18615,N_19263);
nor U20226 (N_20226,N_19481,N_19476);
and U20227 (N_20227,N_18176,N_18060);
nor U20228 (N_20228,N_18551,N_18774);
nor U20229 (N_20229,N_19465,N_18650);
xor U20230 (N_20230,N_19329,N_18960);
nor U20231 (N_20231,N_18950,N_18564);
or U20232 (N_20232,N_18894,N_19065);
nand U20233 (N_20233,N_18470,N_18430);
and U20234 (N_20234,N_18485,N_18319);
or U20235 (N_20235,N_19163,N_18068);
or U20236 (N_20236,N_19337,N_18379);
nand U20237 (N_20237,N_18141,N_19159);
xor U20238 (N_20238,N_18789,N_18326);
nand U20239 (N_20239,N_18368,N_19085);
nor U20240 (N_20240,N_18082,N_18844);
nor U20241 (N_20241,N_18976,N_18025);
nand U20242 (N_20242,N_18098,N_19432);
xor U20243 (N_20243,N_18593,N_18908);
nor U20244 (N_20244,N_19395,N_18214);
nor U20245 (N_20245,N_18754,N_18195);
xnor U20246 (N_20246,N_18452,N_19494);
and U20247 (N_20247,N_19120,N_18133);
nand U20248 (N_20248,N_18677,N_19092);
and U20249 (N_20249,N_18627,N_19203);
nor U20250 (N_20250,N_18033,N_18688);
or U20251 (N_20251,N_19390,N_18051);
and U20252 (N_20252,N_19451,N_18970);
nor U20253 (N_20253,N_19003,N_18206);
and U20254 (N_20254,N_19074,N_18256);
and U20255 (N_20255,N_18564,N_18638);
xnor U20256 (N_20256,N_18418,N_18308);
xnor U20257 (N_20257,N_18608,N_18096);
nor U20258 (N_20258,N_18239,N_18779);
and U20259 (N_20259,N_19262,N_19396);
and U20260 (N_20260,N_18606,N_18899);
or U20261 (N_20261,N_18033,N_19432);
and U20262 (N_20262,N_18546,N_18944);
or U20263 (N_20263,N_18731,N_18205);
and U20264 (N_20264,N_19189,N_18834);
nor U20265 (N_20265,N_18148,N_18712);
or U20266 (N_20266,N_18002,N_18033);
nor U20267 (N_20267,N_19415,N_19377);
nand U20268 (N_20268,N_18680,N_18632);
or U20269 (N_20269,N_18255,N_18868);
xnor U20270 (N_20270,N_19034,N_18423);
nor U20271 (N_20271,N_19498,N_18567);
and U20272 (N_20272,N_19470,N_18533);
xnor U20273 (N_20273,N_18275,N_18452);
nand U20274 (N_20274,N_18729,N_19197);
or U20275 (N_20275,N_19262,N_18622);
or U20276 (N_20276,N_18789,N_18396);
xnor U20277 (N_20277,N_19003,N_19256);
and U20278 (N_20278,N_19160,N_19310);
xnor U20279 (N_20279,N_18875,N_19070);
or U20280 (N_20280,N_18635,N_19175);
xor U20281 (N_20281,N_18784,N_18720);
xnor U20282 (N_20282,N_19117,N_18952);
nor U20283 (N_20283,N_18654,N_18744);
xnor U20284 (N_20284,N_19315,N_18101);
or U20285 (N_20285,N_18600,N_18039);
and U20286 (N_20286,N_18830,N_18283);
nor U20287 (N_20287,N_18717,N_18768);
xor U20288 (N_20288,N_19151,N_18859);
xnor U20289 (N_20289,N_19003,N_18725);
nand U20290 (N_20290,N_18849,N_19462);
or U20291 (N_20291,N_19014,N_18402);
or U20292 (N_20292,N_19115,N_18451);
and U20293 (N_20293,N_18186,N_19284);
nand U20294 (N_20294,N_18801,N_19376);
and U20295 (N_20295,N_19456,N_18207);
xnor U20296 (N_20296,N_19456,N_19392);
nand U20297 (N_20297,N_18355,N_18015);
xor U20298 (N_20298,N_18740,N_19476);
and U20299 (N_20299,N_18394,N_18299);
nor U20300 (N_20300,N_18557,N_18463);
xnor U20301 (N_20301,N_19268,N_18979);
or U20302 (N_20302,N_18609,N_18183);
xor U20303 (N_20303,N_18648,N_19440);
and U20304 (N_20304,N_18026,N_19037);
or U20305 (N_20305,N_18649,N_19432);
nand U20306 (N_20306,N_18738,N_18969);
and U20307 (N_20307,N_19230,N_19416);
nor U20308 (N_20308,N_18321,N_18748);
and U20309 (N_20309,N_18108,N_19408);
nand U20310 (N_20310,N_19137,N_19356);
or U20311 (N_20311,N_19263,N_18953);
nand U20312 (N_20312,N_18819,N_18497);
nor U20313 (N_20313,N_19402,N_19376);
xor U20314 (N_20314,N_18129,N_18010);
and U20315 (N_20315,N_19354,N_19351);
or U20316 (N_20316,N_18221,N_19209);
nand U20317 (N_20317,N_19191,N_18306);
or U20318 (N_20318,N_18996,N_18183);
or U20319 (N_20319,N_18257,N_18522);
xnor U20320 (N_20320,N_18221,N_18485);
nand U20321 (N_20321,N_18693,N_18060);
or U20322 (N_20322,N_19474,N_18251);
xnor U20323 (N_20323,N_19429,N_18704);
nor U20324 (N_20324,N_19084,N_18038);
xnor U20325 (N_20325,N_19117,N_18844);
nor U20326 (N_20326,N_19050,N_19291);
nor U20327 (N_20327,N_18997,N_18548);
xnor U20328 (N_20328,N_19463,N_18578);
or U20329 (N_20329,N_18358,N_18900);
and U20330 (N_20330,N_18399,N_18644);
nor U20331 (N_20331,N_19105,N_19285);
nand U20332 (N_20332,N_18597,N_19014);
nor U20333 (N_20333,N_18111,N_19242);
nor U20334 (N_20334,N_18133,N_18076);
or U20335 (N_20335,N_19208,N_18610);
nand U20336 (N_20336,N_18516,N_19190);
and U20337 (N_20337,N_18063,N_19389);
nand U20338 (N_20338,N_19028,N_18975);
nand U20339 (N_20339,N_18008,N_18345);
or U20340 (N_20340,N_18046,N_18926);
or U20341 (N_20341,N_18859,N_19365);
and U20342 (N_20342,N_18209,N_18753);
nand U20343 (N_20343,N_18368,N_18139);
and U20344 (N_20344,N_19141,N_19095);
nor U20345 (N_20345,N_18625,N_18963);
nand U20346 (N_20346,N_18801,N_18374);
xnor U20347 (N_20347,N_18227,N_18117);
xor U20348 (N_20348,N_18441,N_18424);
nor U20349 (N_20349,N_18073,N_18861);
and U20350 (N_20350,N_18598,N_18837);
nand U20351 (N_20351,N_19228,N_19247);
or U20352 (N_20352,N_19068,N_18752);
nor U20353 (N_20353,N_18614,N_19240);
nor U20354 (N_20354,N_19274,N_18218);
or U20355 (N_20355,N_18330,N_19330);
and U20356 (N_20356,N_19321,N_19416);
xor U20357 (N_20357,N_18930,N_18746);
or U20358 (N_20358,N_18099,N_19388);
xnor U20359 (N_20359,N_18190,N_18640);
nand U20360 (N_20360,N_19050,N_18848);
xnor U20361 (N_20361,N_18068,N_18011);
xnor U20362 (N_20362,N_18756,N_19044);
or U20363 (N_20363,N_19439,N_18238);
nor U20364 (N_20364,N_19389,N_18338);
nor U20365 (N_20365,N_18208,N_18098);
nand U20366 (N_20366,N_19368,N_19209);
nand U20367 (N_20367,N_19436,N_18716);
or U20368 (N_20368,N_19302,N_18101);
nor U20369 (N_20369,N_18696,N_18080);
or U20370 (N_20370,N_18396,N_18895);
or U20371 (N_20371,N_18139,N_18596);
nand U20372 (N_20372,N_18348,N_18995);
nor U20373 (N_20373,N_18918,N_18037);
nor U20374 (N_20374,N_18762,N_18160);
nand U20375 (N_20375,N_18850,N_19175);
nand U20376 (N_20376,N_19125,N_18573);
xor U20377 (N_20377,N_19094,N_19372);
nand U20378 (N_20378,N_19174,N_19337);
nor U20379 (N_20379,N_18503,N_19163);
or U20380 (N_20380,N_18067,N_19071);
nor U20381 (N_20381,N_19107,N_18981);
nand U20382 (N_20382,N_18910,N_19468);
nand U20383 (N_20383,N_19492,N_19011);
xnor U20384 (N_20384,N_18360,N_19057);
nand U20385 (N_20385,N_18436,N_19428);
or U20386 (N_20386,N_19493,N_19269);
or U20387 (N_20387,N_19016,N_19042);
or U20388 (N_20388,N_18138,N_18810);
and U20389 (N_20389,N_19138,N_18390);
xor U20390 (N_20390,N_18982,N_18677);
or U20391 (N_20391,N_18423,N_19326);
nand U20392 (N_20392,N_18334,N_19287);
nor U20393 (N_20393,N_18125,N_19317);
or U20394 (N_20394,N_18173,N_18398);
nand U20395 (N_20395,N_18973,N_18681);
nor U20396 (N_20396,N_19457,N_18280);
and U20397 (N_20397,N_18104,N_19366);
nor U20398 (N_20398,N_18895,N_18513);
nand U20399 (N_20399,N_18170,N_18929);
xnor U20400 (N_20400,N_19366,N_19104);
xor U20401 (N_20401,N_19046,N_18584);
and U20402 (N_20402,N_18074,N_18392);
xnor U20403 (N_20403,N_18645,N_19312);
nor U20404 (N_20404,N_19418,N_18678);
xor U20405 (N_20405,N_19476,N_18244);
or U20406 (N_20406,N_18325,N_18322);
and U20407 (N_20407,N_19200,N_19479);
or U20408 (N_20408,N_18217,N_19095);
nor U20409 (N_20409,N_18666,N_18955);
and U20410 (N_20410,N_18618,N_19227);
or U20411 (N_20411,N_18902,N_18430);
or U20412 (N_20412,N_18689,N_18552);
nor U20413 (N_20413,N_18414,N_19210);
xnor U20414 (N_20414,N_18482,N_19436);
or U20415 (N_20415,N_19065,N_19035);
nor U20416 (N_20416,N_18947,N_18216);
nand U20417 (N_20417,N_18044,N_18761);
nor U20418 (N_20418,N_18024,N_18831);
nor U20419 (N_20419,N_19195,N_19428);
and U20420 (N_20420,N_18050,N_18071);
and U20421 (N_20421,N_18385,N_18278);
and U20422 (N_20422,N_19389,N_19042);
and U20423 (N_20423,N_19331,N_19406);
xnor U20424 (N_20424,N_18196,N_18720);
and U20425 (N_20425,N_18716,N_18675);
nand U20426 (N_20426,N_18701,N_18393);
xnor U20427 (N_20427,N_18343,N_18278);
nand U20428 (N_20428,N_19059,N_19102);
xnor U20429 (N_20429,N_19479,N_19107);
nand U20430 (N_20430,N_19359,N_18368);
and U20431 (N_20431,N_18410,N_19141);
nand U20432 (N_20432,N_18016,N_19336);
or U20433 (N_20433,N_18942,N_18441);
nand U20434 (N_20434,N_18947,N_18964);
or U20435 (N_20435,N_19199,N_18277);
xnor U20436 (N_20436,N_18397,N_19306);
nand U20437 (N_20437,N_19152,N_19080);
or U20438 (N_20438,N_18180,N_18410);
xor U20439 (N_20439,N_18023,N_19174);
xor U20440 (N_20440,N_19269,N_18250);
nand U20441 (N_20441,N_18249,N_19479);
and U20442 (N_20442,N_18648,N_18147);
and U20443 (N_20443,N_18693,N_19144);
nand U20444 (N_20444,N_19442,N_18210);
nor U20445 (N_20445,N_18929,N_19159);
or U20446 (N_20446,N_18951,N_18785);
or U20447 (N_20447,N_18821,N_18964);
nand U20448 (N_20448,N_18906,N_18002);
nor U20449 (N_20449,N_18479,N_18113);
and U20450 (N_20450,N_18811,N_18640);
xor U20451 (N_20451,N_19442,N_19256);
or U20452 (N_20452,N_18912,N_19137);
nor U20453 (N_20453,N_18060,N_18989);
or U20454 (N_20454,N_18499,N_19485);
nor U20455 (N_20455,N_18336,N_18618);
and U20456 (N_20456,N_19038,N_18529);
nand U20457 (N_20457,N_18789,N_19184);
or U20458 (N_20458,N_19191,N_18902);
or U20459 (N_20459,N_18986,N_18004);
nor U20460 (N_20460,N_18940,N_18132);
xor U20461 (N_20461,N_19236,N_19063);
and U20462 (N_20462,N_18489,N_19060);
and U20463 (N_20463,N_19457,N_19427);
nor U20464 (N_20464,N_18314,N_19243);
or U20465 (N_20465,N_19346,N_19438);
nand U20466 (N_20466,N_18636,N_18441);
and U20467 (N_20467,N_18583,N_19297);
xor U20468 (N_20468,N_19288,N_18274);
and U20469 (N_20469,N_18843,N_18448);
nand U20470 (N_20470,N_19298,N_18329);
nor U20471 (N_20471,N_19413,N_19220);
xnor U20472 (N_20472,N_18017,N_18505);
nor U20473 (N_20473,N_18557,N_18478);
nor U20474 (N_20474,N_18015,N_19074);
nand U20475 (N_20475,N_19053,N_19419);
nor U20476 (N_20476,N_18158,N_19141);
and U20477 (N_20477,N_18636,N_18656);
xnor U20478 (N_20478,N_19059,N_18731);
or U20479 (N_20479,N_18391,N_18747);
nor U20480 (N_20480,N_19201,N_19390);
nand U20481 (N_20481,N_18777,N_18429);
xor U20482 (N_20482,N_18153,N_18946);
nor U20483 (N_20483,N_18895,N_19114);
nor U20484 (N_20484,N_18896,N_18577);
xor U20485 (N_20485,N_18379,N_18110);
or U20486 (N_20486,N_18709,N_18035);
nor U20487 (N_20487,N_19319,N_18926);
and U20488 (N_20488,N_18373,N_18717);
or U20489 (N_20489,N_18553,N_18911);
or U20490 (N_20490,N_19137,N_18691);
xnor U20491 (N_20491,N_18079,N_18037);
and U20492 (N_20492,N_18951,N_18313);
xor U20493 (N_20493,N_18258,N_19019);
nor U20494 (N_20494,N_18043,N_19137);
and U20495 (N_20495,N_18854,N_18888);
or U20496 (N_20496,N_18575,N_18982);
xnor U20497 (N_20497,N_18279,N_18070);
nand U20498 (N_20498,N_18560,N_18237);
xnor U20499 (N_20499,N_19373,N_18040);
xor U20500 (N_20500,N_18266,N_19011);
xnor U20501 (N_20501,N_19077,N_19305);
or U20502 (N_20502,N_18972,N_18740);
nand U20503 (N_20503,N_18431,N_18159);
or U20504 (N_20504,N_19371,N_18627);
nor U20505 (N_20505,N_18566,N_18150);
xor U20506 (N_20506,N_18103,N_18143);
nor U20507 (N_20507,N_19477,N_18624);
or U20508 (N_20508,N_19019,N_18675);
and U20509 (N_20509,N_18852,N_19130);
and U20510 (N_20510,N_18298,N_18209);
xnor U20511 (N_20511,N_18361,N_19132);
nor U20512 (N_20512,N_19328,N_19405);
xor U20513 (N_20513,N_18301,N_19345);
xnor U20514 (N_20514,N_18808,N_19424);
and U20515 (N_20515,N_19232,N_19125);
nand U20516 (N_20516,N_19108,N_18596);
or U20517 (N_20517,N_18113,N_18741);
and U20518 (N_20518,N_18879,N_18412);
and U20519 (N_20519,N_18195,N_18129);
nor U20520 (N_20520,N_18891,N_18811);
xor U20521 (N_20521,N_18296,N_19490);
xor U20522 (N_20522,N_18926,N_18928);
nor U20523 (N_20523,N_18118,N_18382);
nor U20524 (N_20524,N_19475,N_19097);
nand U20525 (N_20525,N_18451,N_18016);
and U20526 (N_20526,N_18991,N_18537);
nand U20527 (N_20527,N_19198,N_18355);
xor U20528 (N_20528,N_18155,N_18054);
nand U20529 (N_20529,N_18049,N_19011);
nand U20530 (N_20530,N_19405,N_18633);
nor U20531 (N_20531,N_19281,N_18140);
xor U20532 (N_20532,N_19147,N_18267);
or U20533 (N_20533,N_18110,N_18301);
and U20534 (N_20534,N_18956,N_18779);
and U20535 (N_20535,N_19189,N_18849);
or U20536 (N_20536,N_19061,N_19278);
or U20537 (N_20537,N_19427,N_18590);
nor U20538 (N_20538,N_18210,N_18490);
or U20539 (N_20539,N_18031,N_18379);
nor U20540 (N_20540,N_18823,N_19143);
or U20541 (N_20541,N_18060,N_18823);
nor U20542 (N_20542,N_18749,N_18532);
or U20543 (N_20543,N_18778,N_19166);
nand U20544 (N_20544,N_19442,N_18939);
nand U20545 (N_20545,N_18047,N_18243);
xnor U20546 (N_20546,N_19143,N_18696);
or U20547 (N_20547,N_19468,N_19023);
and U20548 (N_20548,N_19198,N_18276);
nand U20549 (N_20549,N_18391,N_18562);
nor U20550 (N_20550,N_19103,N_18895);
xor U20551 (N_20551,N_19308,N_19454);
nor U20552 (N_20552,N_19429,N_18155);
or U20553 (N_20553,N_19222,N_18818);
nor U20554 (N_20554,N_18838,N_18857);
and U20555 (N_20555,N_19098,N_18306);
nor U20556 (N_20556,N_18270,N_19426);
nor U20557 (N_20557,N_18397,N_18521);
or U20558 (N_20558,N_18727,N_18171);
xor U20559 (N_20559,N_19401,N_18048);
and U20560 (N_20560,N_18564,N_19140);
nand U20561 (N_20561,N_19381,N_19104);
xor U20562 (N_20562,N_18344,N_18234);
nand U20563 (N_20563,N_18440,N_18706);
nor U20564 (N_20564,N_19332,N_19217);
or U20565 (N_20565,N_18259,N_19341);
nand U20566 (N_20566,N_18039,N_18236);
or U20567 (N_20567,N_19086,N_18362);
xnor U20568 (N_20568,N_19269,N_18566);
and U20569 (N_20569,N_19244,N_19092);
and U20570 (N_20570,N_18228,N_19460);
nand U20571 (N_20571,N_18475,N_18084);
or U20572 (N_20572,N_18061,N_18003);
xor U20573 (N_20573,N_18168,N_18796);
or U20574 (N_20574,N_18757,N_18065);
xor U20575 (N_20575,N_19181,N_18518);
nor U20576 (N_20576,N_18528,N_18981);
nand U20577 (N_20577,N_18364,N_19169);
and U20578 (N_20578,N_19356,N_19148);
and U20579 (N_20579,N_19062,N_18190);
and U20580 (N_20580,N_18430,N_18146);
nor U20581 (N_20581,N_18872,N_18751);
xor U20582 (N_20582,N_18302,N_18648);
xnor U20583 (N_20583,N_19487,N_18434);
nand U20584 (N_20584,N_18713,N_19050);
or U20585 (N_20585,N_18950,N_18302);
nand U20586 (N_20586,N_18179,N_18903);
nand U20587 (N_20587,N_18172,N_18620);
xnor U20588 (N_20588,N_18680,N_18887);
nand U20589 (N_20589,N_18823,N_18622);
nand U20590 (N_20590,N_18799,N_18477);
nor U20591 (N_20591,N_18293,N_18583);
xnor U20592 (N_20592,N_19333,N_19253);
or U20593 (N_20593,N_18149,N_18316);
xnor U20594 (N_20594,N_18420,N_19234);
nand U20595 (N_20595,N_19138,N_19139);
xor U20596 (N_20596,N_18311,N_19342);
nor U20597 (N_20597,N_18179,N_18152);
and U20598 (N_20598,N_19396,N_19241);
and U20599 (N_20599,N_18242,N_18748);
nor U20600 (N_20600,N_19436,N_19384);
nor U20601 (N_20601,N_18602,N_18982);
xnor U20602 (N_20602,N_19328,N_18839);
and U20603 (N_20603,N_18993,N_18831);
xnor U20604 (N_20604,N_19401,N_18305);
nor U20605 (N_20605,N_18500,N_18611);
and U20606 (N_20606,N_18154,N_18983);
nor U20607 (N_20607,N_18582,N_18597);
xor U20608 (N_20608,N_18022,N_18942);
nand U20609 (N_20609,N_18188,N_19489);
or U20610 (N_20610,N_18885,N_18296);
nand U20611 (N_20611,N_19235,N_19484);
or U20612 (N_20612,N_18533,N_18018);
nor U20613 (N_20613,N_18491,N_19001);
nor U20614 (N_20614,N_19105,N_18086);
nor U20615 (N_20615,N_19007,N_18262);
and U20616 (N_20616,N_18617,N_18369);
and U20617 (N_20617,N_18885,N_18830);
or U20618 (N_20618,N_18455,N_19323);
nor U20619 (N_20619,N_18788,N_19482);
or U20620 (N_20620,N_18628,N_19037);
nor U20621 (N_20621,N_18348,N_18746);
nor U20622 (N_20622,N_18278,N_18645);
and U20623 (N_20623,N_19046,N_19278);
nor U20624 (N_20624,N_19333,N_18663);
nand U20625 (N_20625,N_18793,N_18111);
and U20626 (N_20626,N_18452,N_18677);
nand U20627 (N_20627,N_18931,N_18669);
nand U20628 (N_20628,N_19209,N_18658);
nor U20629 (N_20629,N_19173,N_18533);
xor U20630 (N_20630,N_18086,N_19242);
xnor U20631 (N_20631,N_19132,N_18899);
nand U20632 (N_20632,N_19005,N_18975);
and U20633 (N_20633,N_19048,N_19289);
nand U20634 (N_20634,N_18360,N_18431);
nand U20635 (N_20635,N_18618,N_19287);
or U20636 (N_20636,N_18223,N_18850);
and U20637 (N_20637,N_18108,N_18822);
nand U20638 (N_20638,N_18951,N_19072);
xor U20639 (N_20639,N_18314,N_19406);
nand U20640 (N_20640,N_18989,N_18043);
or U20641 (N_20641,N_19381,N_18680);
or U20642 (N_20642,N_18370,N_18838);
and U20643 (N_20643,N_18146,N_19396);
nor U20644 (N_20644,N_18661,N_19245);
nand U20645 (N_20645,N_19087,N_18432);
nand U20646 (N_20646,N_18331,N_19215);
and U20647 (N_20647,N_18733,N_18520);
xnor U20648 (N_20648,N_18515,N_18999);
xnor U20649 (N_20649,N_18541,N_19387);
xnor U20650 (N_20650,N_18791,N_18610);
xor U20651 (N_20651,N_19159,N_18904);
nand U20652 (N_20652,N_18861,N_18044);
nor U20653 (N_20653,N_18139,N_19148);
nand U20654 (N_20654,N_19079,N_19443);
and U20655 (N_20655,N_19455,N_19020);
and U20656 (N_20656,N_19247,N_18965);
xnor U20657 (N_20657,N_18953,N_19244);
nand U20658 (N_20658,N_18134,N_18352);
nor U20659 (N_20659,N_18228,N_18696);
nand U20660 (N_20660,N_18437,N_18043);
or U20661 (N_20661,N_18991,N_19414);
xnor U20662 (N_20662,N_18869,N_18261);
nor U20663 (N_20663,N_18282,N_18080);
and U20664 (N_20664,N_18985,N_18044);
xnor U20665 (N_20665,N_18543,N_18281);
nand U20666 (N_20666,N_18406,N_19451);
xnor U20667 (N_20667,N_19157,N_18327);
xor U20668 (N_20668,N_18515,N_18425);
or U20669 (N_20669,N_18367,N_19452);
nor U20670 (N_20670,N_18843,N_19288);
nand U20671 (N_20671,N_19320,N_18022);
and U20672 (N_20672,N_18519,N_18112);
and U20673 (N_20673,N_19365,N_18360);
nand U20674 (N_20674,N_19165,N_18226);
nor U20675 (N_20675,N_18100,N_18517);
and U20676 (N_20676,N_18824,N_18977);
nor U20677 (N_20677,N_19446,N_19379);
xor U20678 (N_20678,N_18685,N_18123);
and U20679 (N_20679,N_18495,N_18588);
nor U20680 (N_20680,N_18566,N_18236);
nor U20681 (N_20681,N_18878,N_19436);
xnor U20682 (N_20682,N_19140,N_18589);
and U20683 (N_20683,N_18397,N_19328);
and U20684 (N_20684,N_18279,N_18956);
and U20685 (N_20685,N_18749,N_18975);
nor U20686 (N_20686,N_18485,N_18764);
and U20687 (N_20687,N_19386,N_18501);
nor U20688 (N_20688,N_19241,N_18111);
nand U20689 (N_20689,N_18669,N_18846);
and U20690 (N_20690,N_18578,N_18399);
or U20691 (N_20691,N_19422,N_18717);
or U20692 (N_20692,N_19000,N_18566);
xnor U20693 (N_20693,N_19316,N_19345);
nand U20694 (N_20694,N_18666,N_19317);
and U20695 (N_20695,N_18319,N_18986);
xnor U20696 (N_20696,N_18286,N_19288);
and U20697 (N_20697,N_18362,N_18779);
and U20698 (N_20698,N_18136,N_19350);
and U20699 (N_20699,N_18699,N_18176);
or U20700 (N_20700,N_18544,N_18927);
nand U20701 (N_20701,N_18238,N_18022);
xor U20702 (N_20702,N_19469,N_19011);
nor U20703 (N_20703,N_18996,N_18226);
nor U20704 (N_20704,N_19296,N_19218);
and U20705 (N_20705,N_18360,N_18114);
nor U20706 (N_20706,N_18782,N_19142);
or U20707 (N_20707,N_18578,N_18559);
xnor U20708 (N_20708,N_19321,N_18568);
and U20709 (N_20709,N_18633,N_19064);
nand U20710 (N_20710,N_18880,N_18429);
nor U20711 (N_20711,N_18524,N_19203);
nand U20712 (N_20712,N_18080,N_18474);
nor U20713 (N_20713,N_18838,N_19007);
nand U20714 (N_20714,N_18552,N_19073);
xnor U20715 (N_20715,N_19445,N_18843);
nand U20716 (N_20716,N_19370,N_19048);
and U20717 (N_20717,N_18559,N_18298);
or U20718 (N_20718,N_18425,N_19418);
nand U20719 (N_20719,N_18973,N_18772);
or U20720 (N_20720,N_19424,N_18415);
xor U20721 (N_20721,N_18213,N_18232);
and U20722 (N_20722,N_19074,N_18320);
and U20723 (N_20723,N_18877,N_18479);
nand U20724 (N_20724,N_18072,N_18627);
xnor U20725 (N_20725,N_18654,N_18134);
nand U20726 (N_20726,N_18996,N_18053);
nor U20727 (N_20727,N_19322,N_19224);
and U20728 (N_20728,N_18836,N_19214);
and U20729 (N_20729,N_18531,N_18566);
xor U20730 (N_20730,N_18654,N_18149);
xnor U20731 (N_20731,N_18054,N_18873);
and U20732 (N_20732,N_19216,N_19242);
nor U20733 (N_20733,N_18793,N_19466);
nor U20734 (N_20734,N_18022,N_19291);
nor U20735 (N_20735,N_18337,N_18116);
or U20736 (N_20736,N_18512,N_18550);
nor U20737 (N_20737,N_18410,N_19392);
nand U20738 (N_20738,N_18152,N_18031);
or U20739 (N_20739,N_18059,N_18292);
nor U20740 (N_20740,N_19029,N_19352);
or U20741 (N_20741,N_19079,N_19445);
xnor U20742 (N_20742,N_18279,N_18460);
or U20743 (N_20743,N_18036,N_18772);
xor U20744 (N_20744,N_18443,N_18330);
nand U20745 (N_20745,N_19448,N_19464);
nand U20746 (N_20746,N_18591,N_18318);
or U20747 (N_20747,N_19261,N_19332);
nand U20748 (N_20748,N_18065,N_18503);
xor U20749 (N_20749,N_19444,N_18876);
xnor U20750 (N_20750,N_18300,N_19054);
or U20751 (N_20751,N_18642,N_19337);
nand U20752 (N_20752,N_18135,N_18837);
and U20753 (N_20753,N_18522,N_18523);
xnor U20754 (N_20754,N_19173,N_18898);
or U20755 (N_20755,N_18265,N_19241);
or U20756 (N_20756,N_18623,N_18921);
nor U20757 (N_20757,N_19181,N_19437);
or U20758 (N_20758,N_18137,N_18460);
xor U20759 (N_20759,N_18141,N_18991);
and U20760 (N_20760,N_18634,N_18997);
nand U20761 (N_20761,N_19283,N_18801);
or U20762 (N_20762,N_18626,N_18714);
or U20763 (N_20763,N_19254,N_18174);
and U20764 (N_20764,N_19209,N_18477);
or U20765 (N_20765,N_19148,N_18165);
and U20766 (N_20766,N_19339,N_18180);
and U20767 (N_20767,N_18054,N_18118);
nor U20768 (N_20768,N_18644,N_18876);
nand U20769 (N_20769,N_18566,N_18738);
and U20770 (N_20770,N_19019,N_19318);
nand U20771 (N_20771,N_19446,N_18818);
nor U20772 (N_20772,N_18642,N_18590);
nand U20773 (N_20773,N_19070,N_19064);
or U20774 (N_20774,N_19487,N_18510);
nand U20775 (N_20775,N_18355,N_18159);
nand U20776 (N_20776,N_18655,N_19055);
xnor U20777 (N_20777,N_18176,N_18809);
or U20778 (N_20778,N_18139,N_18333);
and U20779 (N_20779,N_19161,N_18664);
xnor U20780 (N_20780,N_18434,N_18546);
nand U20781 (N_20781,N_18308,N_19011);
nor U20782 (N_20782,N_18459,N_18454);
or U20783 (N_20783,N_18421,N_18805);
nor U20784 (N_20784,N_19285,N_19136);
or U20785 (N_20785,N_18754,N_18873);
xnor U20786 (N_20786,N_18353,N_18511);
nand U20787 (N_20787,N_19000,N_18774);
nor U20788 (N_20788,N_19420,N_19232);
and U20789 (N_20789,N_18647,N_19277);
nand U20790 (N_20790,N_19409,N_18010);
nand U20791 (N_20791,N_19365,N_18593);
nor U20792 (N_20792,N_18001,N_19434);
nor U20793 (N_20793,N_19487,N_18408);
nand U20794 (N_20794,N_18156,N_18201);
nor U20795 (N_20795,N_19319,N_18529);
nor U20796 (N_20796,N_18487,N_18304);
nor U20797 (N_20797,N_18265,N_18238);
nand U20798 (N_20798,N_18097,N_18447);
nand U20799 (N_20799,N_18481,N_18438);
nor U20800 (N_20800,N_19406,N_18641);
nor U20801 (N_20801,N_18419,N_19463);
nand U20802 (N_20802,N_19098,N_18378);
nor U20803 (N_20803,N_19029,N_18957);
nand U20804 (N_20804,N_18496,N_19131);
or U20805 (N_20805,N_18123,N_18390);
nor U20806 (N_20806,N_18032,N_18658);
nand U20807 (N_20807,N_19447,N_18192);
nor U20808 (N_20808,N_18979,N_18353);
and U20809 (N_20809,N_18677,N_18555);
nand U20810 (N_20810,N_19149,N_18780);
or U20811 (N_20811,N_19385,N_19048);
or U20812 (N_20812,N_19310,N_18541);
or U20813 (N_20813,N_18035,N_18556);
or U20814 (N_20814,N_18607,N_18420);
xor U20815 (N_20815,N_18480,N_19114);
nor U20816 (N_20816,N_19407,N_19007);
xnor U20817 (N_20817,N_19152,N_18967);
and U20818 (N_20818,N_18874,N_18106);
nand U20819 (N_20819,N_19132,N_19259);
or U20820 (N_20820,N_19107,N_19418);
or U20821 (N_20821,N_18711,N_19479);
or U20822 (N_20822,N_19255,N_19257);
xnor U20823 (N_20823,N_18752,N_18003);
or U20824 (N_20824,N_18032,N_18363);
nor U20825 (N_20825,N_18087,N_19256);
nor U20826 (N_20826,N_18796,N_19201);
nand U20827 (N_20827,N_19088,N_18636);
and U20828 (N_20828,N_19039,N_19260);
nand U20829 (N_20829,N_19156,N_19287);
xnor U20830 (N_20830,N_18345,N_18216);
and U20831 (N_20831,N_18122,N_18920);
and U20832 (N_20832,N_19185,N_18729);
xnor U20833 (N_20833,N_18566,N_18594);
nor U20834 (N_20834,N_19292,N_19110);
nor U20835 (N_20835,N_19321,N_18428);
nand U20836 (N_20836,N_18351,N_18032);
nand U20837 (N_20837,N_18196,N_18893);
and U20838 (N_20838,N_19096,N_18373);
or U20839 (N_20839,N_18108,N_19187);
nand U20840 (N_20840,N_19291,N_19306);
or U20841 (N_20841,N_19201,N_18350);
xor U20842 (N_20842,N_18306,N_19210);
nor U20843 (N_20843,N_19202,N_18181);
and U20844 (N_20844,N_19216,N_18762);
xnor U20845 (N_20845,N_18023,N_18885);
nand U20846 (N_20846,N_18693,N_19299);
xnor U20847 (N_20847,N_18802,N_18956);
or U20848 (N_20848,N_18482,N_18248);
or U20849 (N_20849,N_18431,N_18781);
or U20850 (N_20850,N_18529,N_18323);
xnor U20851 (N_20851,N_19042,N_19049);
and U20852 (N_20852,N_18078,N_18682);
nor U20853 (N_20853,N_19438,N_18861);
nand U20854 (N_20854,N_18716,N_19495);
nor U20855 (N_20855,N_18153,N_18222);
xor U20856 (N_20856,N_18824,N_18097);
or U20857 (N_20857,N_18733,N_18522);
or U20858 (N_20858,N_18238,N_19408);
and U20859 (N_20859,N_18596,N_19206);
and U20860 (N_20860,N_18444,N_19152);
nand U20861 (N_20861,N_18393,N_18065);
or U20862 (N_20862,N_18330,N_18966);
xnor U20863 (N_20863,N_19353,N_18400);
or U20864 (N_20864,N_19194,N_18179);
xor U20865 (N_20865,N_19495,N_19127);
xnor U20866 (N_20866,N_19156,N_18739);
and U20867 (N_20867,N_18319,N_19442);
xnor U20868 (N_20868,N_19182,N_18837);
nor U20869 (N_20869,N_19495,N_18932);
nand U20870 (N_20870,N_19375,N_19450);
nor U20871 (N_20871,N_19003,N_19181);
or U20872 (N_20872,N_18175,N_19388);
nand U20873 (N_20873,N_19276,N_18361);
nand U20874 (N_20874,N_18802,N_19032);
or U20875 (N_20875,N_18910,N_19367);
nand U20876 (N_20876,N_19155,N_18252);
and U20877 (N_20877,N_18402,N_18127);
or U20878 (N_20878,N_19499,N_18083);
xor U20879 (N_20879,N_18073,N_19026);
and U20880 (N_20880,N_18981,N_18560);
xor U20881 (N_20881,N_18509,N_18949);
nand U20882 (N_20882,N_19427,N_18322);
and U20883 (N_20883,N_19371,N_18196);
nor U20884 (N_20884,N_19027,N_18803);
xnor U20885 (N_20885,N_18686,N_18544);
or U20886 (N_20886,N_19374,N_18027);
and U20887 (N_20887,N_18409,N_18536);
and U20888 (N_20888,N_18416,N_19287);
nand U20889 (N_20889,N_18749,N_18258);
nand U20890 (N_20890,N_18025,N_19302);
xnor U20891 (N_20891,N_18154,N_18176);
or U20892 (N_20892,N_19247,N_19266);
and U20893 (N_20893,N_18352,N_18899);
or U20894 (N_20894,N_18084,N_18516);
and U20895 (N_20895,N_19380,N_19128);
or U20896 (N_20896,N_18700,N_18515);
and U20897 (N_20897,N_19091,N_18433);
nor U20898 (N_20898,N_18977,N_18059);
and U20899 (N_20899,N_19224,N_18697);
or U20900 (N_20900,N_19494,N_18558);
and U20901 (N_20901,N_18480,N_18941);
or U20902 (N_20902,N_18976,N_18505);
or U20903 (N_20903,N_18923,N_18803);
and U20904 (N_20904,N_18285,N_18048);
or U20905 (N_20905,N_19231,N_19406);
nand U20906 (N_20906,N_18510,N_18994);
and U20907 (N_20907,N_18455,N_18318);
or U20908 (N_20908,N_18408,N_18582);
xor U20909 (N_20909,N_18074,N_18749);
nand U20910 (N_20910,N_19006,N_18982);
nand U20911 (N_20911,N_18777,N_18555);
and U20912 (N_20912,N_18120,N_18774);
nand U20913 (N_20913,N_18643,N_18272);
nor U20914 (N_20914,N_18793,N_18992);
and U20915 (N_20915,N_19424,N_18040);
or U20916 (N_20916,N_18612,N_19407);
or U20917 (N_20917,N_18310,N_19389);
or U20918 (N_20918,N_18111,N_19339);
and U20919 (N_20919,N_19390,N_18967);
nor U20920 (N_20920,N_18935,N_18263);
or U20921 (N_20921,N_19107,N_19069);
nor U20922 (N_20922,N_19246,N_19158);
nor U20923 (N_20923,N_18064,N_19049);
xnor U20924 (N_20924,N_19203,N_19457);
or U20925 (N_20925,N_18801,N_19205);
or U20926 (N_20926,N_18348,N_18452);
and U20927 (N_20927,N_18245,N_18259);
nor U20928 (N_20928,N_19262,N_19378);
nand U20929 (N_20929,N_18191,N_19402);
nor U20930 (N_20930,N_18130,N_19397);
and U20931 (N_20931,N_18193,N_18451);
and U20932 (N_20932,N_18490,N_18116);
nand U20933 (N_20933,N_19126,N_18213);
and U20934 (N_20934,N_18822,N_19187);
nand U20935 (N_20935,N_18466,N_18578);
and U20936 (N_20936,N_19346,N_18449);
or U20937 (N_20937,N_18346,N_18504);
and U20938 (N_20938,N_18195,N_19254);
nor U20939 (N_20939,N_18504,N_19267);
or U20940 (N_20940,N_18979,N_18558);
or U20941 (N_20941,N_19422,N_19325);
xor U20942 (N_20942,N_18076,N_18232);
xor U20943 (N_20943,N_18793,N_18014);
or U20944 (N_20944,N_18603,N_18756);
xor U20945 (N_20945,N_19373,N_19139);
or U20946 (N_20946,N_19305,N_19008);
nor U20947 (N_20947,N_18941,N_19325);
nor U20948 (N_20948,N_19158,N_19455);
xnor U20949 (N_20949,N_18276,N_19038);
and U20950 (N_20950,N_18556,N_19241);
and U20951 (N_20951,N_19446,N_18486);
nor U20952 (N_20952,N_18724,N_19265);
and U20953 (N_20953,N_18042,N_19476);
nor U20954 (N_20954,N_19293,N_18229);
xor U20955 (N_20955,N_18481,N_18024);
nand U20956 (N_20956,N_19442,N_19208);
and U20957 (N_20957,N_18443,N_18863);
or U20958 (N_20958,N_18508,N_18206);
xor U20959 (N_20959,N_18919,N_18009);
nand U20960 (N_20960,N_18500,N_18714);
and U20961 (N_20961,N_18798,N_18730);
or U20962 (N_20962,N_18030,N_18068);
or U20963 (N_20963,N_19253,N_19497);
nor U20964 (N_20964,N_19231,N_19215);
or U20965 (N_20965,N_18876,N_19465);
and U20966 (N_20966,N_18865,N_19366);
xor U20967 (N_20967,N_18595,N_19058);
xnor U20968 (N_20968,N_18401,N_19238);
and U20969 (N_20969,N_19161,N_19450);
nand U20970 (N_20970,N_19402,N_19458);
or U20971 (N_20971,N_19418,N_18612);
nand U20972 (N_20972,N_18631,N_18639);
nor U20973 (N_20973,N_18587,N_18701);
nand U20974 (N_20974,N_18097,N_19029);
xor U20975 (N_20975,N_19285,N_18332);
and U20976 (N_20976,N_18381,N_19085);
and U20977 (N_20977,N_19031,N_18789);
xnor U20978 (N_20978,N_18485,N_18005);
nand U20979 (N_20979,N_19373,N_19196);
nor U20980 (N_20980,N_18360,N_18660);
and U20981 (N_20981,N_18604,N_18511);
and U20982 (N_20982,N_18512,N_18910);
or U20983 (N_20983,N_18337,N_19238);
xnor U20984 (N_20984,N_18184,N_18537);
and U20985 (N_20985,N_19115,N_19274);
or U20986 (N_20986,N_19004,N_18012);
xnor U20987 (N_20987,N_18830,N_18394);
xor U20988 (N_20988,N_18331,N_19274);
or U20989 (N_20989,N_19263,N_18881);
nor U20990 (N_20990,N_18100,N_18393);
nor U20991 (N_20991,N_19161,N_18334);
or U20992 (N_20992,N_18980,N_18466);
or U20993 (N_20993,N_19068,N_18201);
or U20994 (N_20994,N_18512,N_19163);
nor U20995 (N_20995,N_18424,N_18476);
or U20996 (N_20996,N_18294,N_18610);
or U20997 (N_20997,N_18981,N_18770);
and U20998 (N_20998,N_18808,N_19223);
or U20999 (N_20999,N_19448,N_18329);
nor U21000 (N_21000,N_20147,N_20023);
or U21001 (N_21001,N_20884,N_20293);
nor U21002 (N_21002,N_19950,N_20094);
nand U21003 (N_21003,N_20126,N_19598);
nor U21004 (N_21004,N_20078,N_20607);
nand U21005 (N_21005,N_20201,N_20944);
xnor U21006 (N_21006,N_20509,N_20631);
nor U21007 (N_21007,N_20790,N_20617);
and U21008 (N_21008,N_20908,N_19707);
and U21009 (N_21009,N_20542,N_20350);
xor U21010 (N_21010,N_19640,N_20653);
nor U21011 (N_21011,N_19574,N_19838);
xor U21012 (N_21012,N_19505,N_20751);
xor U21013 (N_21013,N_20709,N_19647);
nand U21014 (N_21014,N_20981,N_20251);
nand U21015 (N_21015,N_20317,N_20222);
and U21016 (N_21016,N_20255,N_20046);
or U21017 (N_21017,N_20173,N_20907);
nand U21018 (N_21018,N_20633,N_20110);
or U21019 (N_21019,N_20732,N_20911);
xnor U21020 (N_21020,N_19846,N_20713);
or U21021 (N_21021,N_20168,N_20243);
xnor U21022 (N_21022,N_19655,N_20995);
and U21023 (N_21023,N_20053,N_20315);
and U21024 (N_21024,N_20465,N_20118);
or U21025 (N_21025,N_20368,N_20913);
or U21026 (N_21026,N_19861,N_19829);
nand U21027 (N_21027,N_20287,N_20540);
and U21028 (N_21028,N_20467,N_20754);
nor U21029 (N_21029,N_19924,N_20629);
or U21030 (N_21030,N_19964,N_20026);
nand U21031 (N_21031,N_20184,N_20331);
nand U21032 (N_21032,N_20226,N_20979);
nor U21033 (N_21033,N_19652,N_20820);
and U21034 (N_21034,N_20796,N_19600);
or U21035 (N_21035,N_20055,N_19824);
nand U21036 (N_21036,N_20530,N_20941);
nand U21037 (N_21037,N_19562,N_19943);
or U21038 (N_21038,N_20037,N_19526);
and U21039 (N_21039,N_20616,N_20558);
nand U21040 (N_21040,N_19591,N_20160);
and U21041 (N_21041,N_20186,N_20901);
nand U21042 (N_21042,N_19547,N_20143);
nor U21043 (N_21043,N_19587,N_20625);
xor U21044 (N_21044,N_20430,N_19999);
nand U21045 (N_21045,N_20389,N_20560);
or U21046 (N_21046,N_20415,N_20033);
and U21047 (N_21047,N_19650,N_20978);
nand U21048 (N_21048,N_20566,N_19544);
and U21049 (N_21049,N_19874,N_19528);
nor U21050 (N_21050,N_20440,N_20417);
or U21051 (N_21051,N_20262,N_20228);
nor U21052 (N_21052,N_20685,N_20497);
xnor U21053 (N_21053,N_20909,N_20066);
xor U21054 (N_21054,N_19963,N_20446);
nor U21055 (N_21055,N_19792,N_20920);
or U21056 (N_21056,N_20610,N_20730);
nor U21057 (N_21057,N_19810,N_20237);
xor U21058 (N_21058,N_20298,N_20710);
xnor U21059 (N_21059,N_20673,N_20665);
nand U21060 (N_21060,N_19847,N_20496);
xnor U21061 (N_21061,N_20933,N_20463);
xor U21062 (N_21062,N_20635,N_20883);
xor U21063 (N_21063,N_19932,N_19721);
xnor U21064 (N_21064,N_19651,N_19749);
nand U21065 (N_21065,N_20444,N_19850);
and U21066 (N_21066,N_19565,N_20830);
and U21067 (N_21067,N_20290,N_20586);
xor U21068 (N_21068,N_20271,N_20659);
nor U21069 (N_21069,N_20414,N_19585);
nor U21070 (N_21070,N_20547,N_20916);
nor U21071 (N_21071,N_20523,N_20829);
nand U21072 (N_21072,N_20443,N_20439);
or U21073 (N_21073,N_20205,N_19606);
xnor U21074 (N_21074,N_20674,N_20195);
nand U21075 (N_21075,N_19524,N_19772);
nor U21076 (N_21076,N_20000,N_20208);
nor U21077 (N_21077,N_20539,N_20162);
and U21078 (N_21078,N_20366,N_19513);
and U21079 (N_21079,N_19694,N_19763);
or U21080 (N_21080,N_20409,N_20548);
xnor U21081 (N_21081,N_20203,N_20488);
nand U21082 (N_21082,N_19614,N_20994);
nor U21083 (N_21083,N_20970,N_19827);
nor U21084 (N_21084,N_20087,N_20307);
and U21085 (N_21085,N_20371,N_19567);
and U21086 (N_21086,N_19835,N_19822);
xor U21087 (N_21087,N_20945,N_20434);
nand U21088 (N_21088,N_20642,N_20795);
nand U21089 (N_21089,N_20182,N_20137);
or U21090 (N_21090,N_20515,N_19560);
or U21091 (N_21091,N_20013,N_20257);
xor U21092 (N_21092,N_20050,N_20581);
nand U21093 (N_21093,N_20082,N_20282);
nor U21094 (N_21094,N_20520,N_20499);
nor U21095 (N_21095,N_19564,N_20999);
and U21096 (N_21096,N_19938,N_19746);
and U21097 (N_21097,N_20375,N_19751);
and U21098 (N_21098,N_20934,N_20516);
nand U21099 (N_21099,N_20645,N_20157);
nand U21100 (N_21100,N_20967,N_19823);
xor U21101 (N_21101,N_19788,N_20985);
nor U21102 (N_21102,N_20382,N_20454);
nand U21103 (N_21103,N_20461,N_19902);
or U21104 (N_21104,N_19516,N_20245);
nor U21105 (N_21105,N_19501,N_20860);
or U21106 (N_21106,N_20639,N_20272);
nand U21107 (N_21107,N_19580,N_20935);
or U21108 (N_21108,N_20025,N_20154);
xor U21109 (N_21109,N_20852,N_19919);
xor U21110 (N_21110,N_20242,N_19762);
xor U21111 (N_21111,N_19882,N_19812);
nor U21112 (N_21112,N_20622,N_20779);
nor U21113 (N_21113,N_20738,N_19977);
nand U21114 (N_21114,N_20127,N_19890);
xnor U21115 (N_21115,N_20768,N_20204);
or U21116 (N_21116,N_20445,N_20777);
and U21117 (N_21117,N_20554,N_19594);
or U21118 (N_21118,N_20717,N_20240);
xor U21119 (N_21119,N_20648,N_20517);
nor U21120 (N_21120,N_19857,N_19535);
nand U21121 (N_21121,N_19658,N_20506);
nand U21122 (N_21122,N_20274,N_19904);
nand U21123 (N_21123,N_19669,N_20169);
or U21124 (N_21124,N_20024,N_20672);
nand U21125 (N_21125,N_20976,N_20012);
nor U21126 (N_21126,N_20652,N_20453);
or U21127 (N_21127,N_20482,N_19660);
or U21128 (N_21128,N_19631,N_20031);
nand U21129 (N_21129,N_19778,N_20597);
and U21130 (N_21130,N_20585,N_19682);
nor U21131 (N_21131,N_20872,N_20239);
or U21132 (N_21132,N_20437,N_19512);
nor U21133 (N_21133,N_20474,N_20602);
xor U21134 (N_21134,N_19685,N_20011);
nand U21135 (N_21135,N_20227,N_20148);
nand U21136 (N_21136,N_20888,N_19733);
or U21137 (N_21137,N_20063,N_19803);
or U21138 (N_21138,N_20335,N_20057);
and U21139 (N_21139,N_20654,N_20526);
nor U21140 (N_21140,N_20265,N_20817);
and U21141 (N_21141,N_20327,N_19680);
nand U21142 (N_21142,N_19961,N_20522);
nor U21143 (N_21143,N_19716,N_20885);
xor U21144 (N_21144,N_20667,N_20952);
and U21145 (N_21145,N_20229,N_19538);
nor U21146 (N_21146,N_19825,N_19500);
or U21147 (N_21147,N_19689,N_20731);
nor U21148 (N_21148,N_20767,N_20197);
nor U21149 (N_21149,N_20662,N_19933);
nor U21150 (N_21150,N_19980,N_20305);
nand U21151 (N_21151,N_20707,N_20345);
nand U21152 (N_21152,N_20704,N_19880);
and U21153 (N_21153,N_20525,N_19639);
nor U21154 (N_21154,N_19706,N_20045);
xor U21155 (N_21155,N_20666,N_19627);
xnor U21156 (N_21156,N_20728,N_20249);
nand U21157 (N_21157,N_20743,N_20161);
and U21158 (N_21158,N_19947,N_19920);
or U21159 (N_21159,N_20093,N_19901);
nand U21160 (N_21160,N_20306,N_20775);
and U21161 (N_21161,N_19612,N_19998);
nor U21162 (N_21162,N_19917,N_20561);
nand U21163 (N_21163,N_20889,N_20988);
nand U21164 (N_21164,N_20246,N_20660);
or U21165 (N_21165,N_20125,N_19821);
or U21166 (N_21166,N_20951,N_20362);
xnor U21167 (N_21167,N_20213,N_20601);
nand U21168 (N_21168,N_20452,N_20179);
nor U21169 (N_21169,N_20144,N_19563);
xor U21170 (N_21170,N_20896,N_20181);
xor U21171 (N_21171,N_20798,N_20577);
or U21172 (N_21172,N_20176,N_20634);
and U21173 (N_21173,N_20878,N_20065);
or U21174 (N_21174,N_20569,N_20698);
nand U21175 (N_21175,N_19782,N_19724);
nor U21176 (N_21176,N_19806,N_19670);
or U21177 (N_21177,N_20359,N_19704);
xnor U21178 (N_21178,N_20841,N_19997);
xnor U21179 (N_21179,N_20259,N_19604);
or U21180 (N_21180,N_19845,N_19556);
and U21181 (N_21181,N_20591,N_19826);
nor U21182 (N_21182,N_20870,N_20688);
nand U21183 (N_21183,N_19542,N_19726);
xor U21184 (N_21184,N_20683,N_19653);
nor U21185 (N_21185,N_20675,N_20070);
nor U21186 (N_21186,N_20253,N_20756);
nand U21187 (N_21187,N_20328,N_20549);
or U21188 (N_21188,N_20962,N_19583);
xor U21189 (N_21189,N_20131,N_20394);
or U21190 (N_21190,N_19711,N_20048);
or U21191 (N_21191,N_19832,N_20734);
or U21192 (N_21192,N_19601,N_19520);
nor U21193 (N_21193,N_20799,N_19671);
xnor U21194 (N_21194,N_19799,N_19855);
and U21195 (N_21195,N_20122,N_19765);
xnor U21196 (N_21196,N_20408,N_19984);
nor U21197 (N_21197,N_20477,N_20291);
and U21198 (N_21198,N_20060,N_20977);
or U21199 (N_21199,N_19588,N_20469);
nand U21200 (N_21200,N_19602,N_20947);
or U21201 (N_21201,N_19797,N_19939);
and U21202 (N_21202,N_20599,N_20034);
and U21203 (N_21203,N_20297,N_19960);
nor U21204 (N_21204,N_19989,N_19703);
and U21205 (N_21205,N_19876,N_19622);
nand U21206 (N_21206,N_20397,N_20129);
nor U21207 (N_21207,N_20363,N_20062);
or U21208 (N_21208,N_20192,N_20369);
nand U21209 (N_21209,N_20355,N_19698);
and U21210 (N_21210,N_20442,N_20457);
xor U21211 (N_21211,N_19552,N_20395);
or U21212 (N_21212,N_20887,N_20924);
nand U21213 (N_21213,N_19905,N_20159);
nor U21214 (N_21214,N_20527,N_20493);
and U21215 (N_21215,N_19723,N_19931);
nand U21216 (N_21216,N_19854,N_20875);
nor U21217 (N_21217,N_20036,N_20391);
nor U21218 (N_21218,N_20280,N_19550);
nand U21219 (N_21219,N_20803,N_20460);
or U21220 (N_21220,N_20950,N_20998);
xnor U21221 (N_21221,N_19735,N_20720);
or U21222 (N_21222,N_20535,N_19828);
nor U21223 (N_21223,N_19579,N_20320);
nand U21224 (N_21224,N_20824,N_19713);
nor U21225 (N_21225,N_20559,N_20470);
and U21226 (N_21226,N_20780,N_20982);
or U21227 (N_21227,N_19586,N_19798);
nand U21228 (N_21228,N_20762,N_20725);
nand U21229 (N_21229,N_19523,N_20481);
or U21230 (N_21230,N_20845,N_19739);
nand U21231 (N_21231,N_20553,N_20658);
and U21232 (N_21232,N_19884,N_19618);
nand U21233 (N_21233,N_19915,N_20448);
nor U21234 (N_21234,N_20130,N_20876);
and U21235 (N_21235,N_20869,N_20124);
nor U21236 (N_21236,N_20311,N_20400);
or U21237 (N_21237,N_19804,N_20111);
nor U21238 (N_21238,N_20637,N_20727);
xnor U21239 (N_21239,N_20624,N_20270);
or U21240 (N_21240,N_19708,N_20628);
nand U21241 (N_21241,N_20149,N_19576);
and U21242 (N_21242,N_20574,N_19611);
nor U21243 (N_21243,N_20199,N_20302);
or U21244 (N_21244,N_19701,N_19796);
and U21245 (N_21245,N_20712,N_20260);
nor U21246 (N_21246,N_20578,N_20029);
xor U21247 (N_21247,N_20038,N_20552);
or U21248 (N_21248,N_20407,N_19819);
nand U21249 (N_21249,N_20505,N_20723);
and U21250 (N_21250,N_19949,N_19774);
nand U21251 (N_21251,N_20200,N_20073);
nand U21252 (N_21252,N_19510,N_19581);
or U21253 (N_21253,N_20922,N_20379);
and U21254 (N_21254,N_20840,N_20533);
xor U21255 (N_21255,N_20042,N_19787);
and U21256 (N_21256,N_20411,N_20806);
nand U21257 (N_21257,N_20353,N_20956);
and U21258 (N_21258,N_19750,N_19633);
nor U21259 (N_21259,N_20483,N_20356);
and U21260 (N_21260,N_20510,N_20096);
xnor U21261 (N_21261,N_20974,N_20823);
or U21262 (N_21262,N_19929,N_20172);
and U21263 (N_21263,N_19554,N_20690);
nand U21264 (N_21264,N_20039,N_20647);
or U21265 (N_21265,N_20833,N_19993);
nand U21266 (N_21266,N_19910,N_20451);
and U21267 (N_21267,N_20651,N_20447);
nand U21268 (N_21268,N_20233,N_19764);
nor U21269 (N_21269,N_20735,N_20296);
and U21270 (N_21270,N_20354,N_19789);
nand U21271 (N_21271,N_19599,N_20807);
and U21272 (N_21272,N_20582,N_20746);
nor U21273 (N_21273,N_19662,N_19519);
or U21274 (N_21274,N_19971,N_20018);
or U21275 (N_21275,N_20164,N_20134);
and U21276 (N_21276,N_19979,N_20749);
and U21277 (N_21277,N_20004,N_20808);
xor U21278 (N_21278,N_20183,N_20189);
and U21279 (N_21279,N_19504,N_20113);
nor U21280 (N_21280,N_20618,N_19946);
or U21281 (N_21281,N_20592,N_19521);
xor U21282 (N_21282,N_20401,N_20646);
and U21283 (N_21283,N_20322,N_19781);
nand U21284 (N_21284,N_19575,N_20514);
nor U21285 (N_21285,N_19957,N_20489);
and U21286 (N_21286,N_20670,N_20010);
nor U21287 (N_21287,N_20668,N_20859);
nand U21288 (N_21288,N_19690,N_19561);
and U21289 (N_21289,N_19678,N_20421);
or U21290 (N_21290,N_19934,N_19968);
nand U21291 (N_21291,N_20216,N_20902);
xor U21292 (N_21292,N_19955,N_20028);
xnor U21293 (N_21293,N_19952,N_19632);
nand U21294 (N_21294,N_20546,N_20219);
nor U21295 (N_21295,N_19744,N_20750);
xor U21296 (N_21296,N_20288,N_20825);
and U21297 (N_21297,N_20100,N_20404);
and U21298 (N_21298,N_19996,N_20276);
and U21299 (N_21299,N_20612,N_20759);
nor U21300 (N_21300,N_20891,N_20937);
or U21301 (N_21301,N_19784,N_20623);
nor U21302 (N_21302,N_19686,N_20881);
and U21303 (N_21303,N_19529,N_19783);
nand U21304 (N_21304,N_20615,N_20507);
or U21305 (N_21305,N_20300,N_20007);
or U21306 (N_21306,N_19770,N_20109);
nand U21307 (N_21307,N_20794,N_20816);
or U21308 (N_21308,N_19502,N_19696);
nor U21309 (N_21309,N_20171,N_20609);
nor U21310 (N_21310,N_19973,N_19986);
nor U21311 (N_21311,N_20850,N_19503);
and U21312 (N_21312,N_20049,N_20472);
nor U21313 (N_21313,N_20273,N_19755);
xor U21314 (N_21314,N_20563,N_20009);
xor U21315 (N_21315,N_19841,N_20386);
nand U21316 (N_21316,N_19815,N_19908);
nor U21317 (N_21317,N_20531,N_20696);
xor U21318 (N_21318,N_20008,N_20681);
and U21319 (N_21319,N_20016,N_20416);
nand U21320 (N_21320,N_20763,N_20103);
nor U21321 (N_21321,N_20487,N_20815);
nor U21322 (N_21322,N_19729,N_19687);
and U21323 (N_21323,N_19898,N_20158);
or U21324 (N_21324,N_19518,N_19572);
or U21325 (N_21325,N_20102,N_19752);
nand U21326 (N_21326,N_20855,N_20740);
or U21327 (N_21327,N_20502,N_20410);
or U21328 (N_21328,N_20556,N_20943);
xor U21329 (N_21329,N_20090,N_19509);
nand U21330 (N_21330,N_20792,N_20965);
or U21331 (N_21331,N_19665,N_20608);
xnor U21332 (N_21332,N_20001,N_20781);
and U21333 (N_21333,N_20972,N_20865);
nor U21334 (N_21334,N_20949,N_20248);
nor U21335 (N_21335,N_19941,N_20565);
nand U21336 (N_21336,N_20649,N_19754);
and U21337 (N_21337,N_19745,N_20211);
or U21338 (N_21338,N_20931,N_20996);
or U21339 (N_21339,N_19702,N_20479);
and U21340 (N_21340,N_19641,N_19531);
xnor U21341 (N_21341,N_20098,N_20364);
nand U21342 (N_21342,N_19864,N_20429);
or U21343 (N_21343,N_20402,N_19831);
xnor U21344 (N_21344,N_20374,N_20800);
nor U21345 (N_21345,N_19930,N_19892);
xor U21346 (N_21346,N_20333,N_19759);
xor U21347 (N_21347,N_20308,N_20705);
nand U21348 (N_21348,N_19753,N_19661);
nand U21349 (N_21349,N_20492,N_19870);
nor U21350 (N_21350,N_19860,N_19868);
or U21351 (N_21351,N_19843,N_20708);
and U21352 (N_21352,N_20106,N_20321);
or U21353 (N_21353,N_20420,N_20180);
nor U21354 (N_21354,N_20518,N_19568);
nand U21355 (N_21355,N_20721,N_20140);
or U21356 (N_21356,N_20084,N_20643);
and U21357 (N_21357,N_20729,N_19942);
xor U21358 (N_21358,N_20567,N_20471);
nor U21359 (N_21359,N_19863,N_20283);
or U21360 (N_21360,N_19675,N_20701);
or U21361 (N_21361,N_20726,N_19982);
nor U21362 (N_21362,N_19883,N_20174);
or U21363 (N_21363,N_20819,N_19922);
xor U21364 (N_21364,N_19710,N_20303);
and U21365 (N_21365,N_20692,N_20963);
and U21366 (N_21366,N_20689,N_20940);
xnor U21367 (N_21367,N_20209,N_20231);
nor U21368 (N_21368,N_20583,N_20543);
nand U21369 (N_21369,N_20564,N_20519);
and U21370 (N_21370,N_19899,N_19916);
and U21371 (N_21371,N_20459,N_20501);
nand U21372 (N_21372,N_20381,N_19911);
nand U21373 (N_21373,N_19985,N_20532);
xnor U21374 (N_21374,N_19515,N_20334);
and U21375 (N_21375,N_20880,N_20812);
nand U21376 (N_21376,N_19909,N_20809);
nand U21377 (N_21377,N_19715,N_20772);
or U21378 (N_21378,N_20292,N_20142);
nand U21379 (N_21379,N_19621,N_20105);
or U21380 (N_21380,N_20277,N_19914);
and U21381 (N_21381,N_19967,N_20206);
xnor U21382 (N_21382,N_19779,N_20663);
xnor U21383 (N_21383,N_20117,N_20352);
or U21384 (N_21384,N_19966,N_20244);
and U21385 (N_21385,N_19616,N_19743);
and U21386 (N_21386,N_20990,N_19780);
and U21387 (N_21387,N_20702,N_20221);
nand U21388 (N_21388,N_19557,N_19543);
or U21389 (N_21389,N_20571,N_20871);
nand U21390 (N_21390,N_20418,N_19673);
or U21391 (N_21391,N_20043,N_19748);
and U21392 (N_21392,N_20005,N_20851);
or U21393 (N_21393,N_20786,N_20827);
and U21394 (N_21394,N_20177,N_19906);
nor U21395 (N_21395,N_19813,N_20344);
nand U21396 (N_21396,N_19615,N_19642);
nand U21397 (N_21397,N_20771,N_20748);
or U21398 (N_21398,N_20324,N_19741);
and U21399 (N_21399,N_20022,N_20224);
nor U21400 (N_21400,N_20108,N_19805);
and U21401 (N_21401,N_20811,N_20831);
or U21402 (N_21402,N_19866,N_20006);
or U21403 (N_21403,N_20058,N_19873);
or U21404 (N_21404,N_19771,N_20165);
xnor U21405 (N_21405,N_19705,N_19730);
nand U21406 (N_21406,N_20266,N_19684);
xnor U21407 (N_21407,N_20684,N_19817);
or U21408 (N_21408,N_19717,N_19928);
and U21409 (N_21409,N_20114,N_19695);
and U21410 (N_21410,N_19649,N_20146);
xnor U21411 (N_21411,N_20150,N_20071);
xor U21412 (N_21412,N_19987,N_20484);
and U21413 (N_21413,N_20787,N_19636);
nor U21414 (N_21414,N_20938,N_19683);
xnor U21415 (N_21415,N_19619,N_19837);
xor U21416 (N_21416,N_20478,N_19786);
nand U21417 (N_21417,N_20644,N_20284);
nor U21418 (N_21418,N_19969,N_19912);
and U21419 (N_21419,N_19645,N_20846);
or U21420 (N_21420,N_19732,N_20893);
xnor U21421 (N_21421,N_20942,N_20264);
or U21422 (N_21422,N_19777,N_19761);
and U21423 (N_21423,N_20765,N_20318);
xor U21424 (N_21424,N_20905,N_20849);
nor U21425 (N_21425,N_19699,N_19918);
and U21426 (N_21426,N_20198,N_20661);
xor U21427 (N_21427,N_19954,N_20279);
nand U21428 (N_21428,N_20960,N_19545);
nand U21429 (N_21429,N_20217,N_20782);
nor U21430 (N_21430,N_20744,N_19959);
nand U21431 (N_21431,N_20312,N_20393);
or U21432 (N_21432,N_20691,N_20485);
nor U21433 (N_21433,N_20801,N_20955);
nor U21434 (N_21434,N_20632,N_19956);
or U21435 (N_21435,N_20433,N_20207);
nand U21436 (N_21436,N_20638,N_19718);
nand U21437 (N_21437,N_20676,N_19921);
nor U21438 (N_21438,N_20613,N_19700);
nand U21439 (N_21439,N_19527,N_20099);
nor U21440 (N_21440,N_19728,N_19532);
and U21441 (N_21441,N_20611,N_20475);
and U21442 (N_21442,N_20551,N_20858);
and U21443 (N_21443,N_20572,N_19584);
nand U21444 (N_21444,N_19852,N_20636);
and U21445 (N_21445,N_20462,N_20839);
and U21446 (N_21446,N_20722,N_20052);
and U21447 (N_21447,N_20399,N_20733);
and U21448 (N_21448,N_20241,N_19858);
or U21449 (N_21449,N_19625,N_20867);
nor U21450 (N_21450,N_20513,N_20576);
or U21451 (N_21451,N_20900,N_19807);
and U21452 (N_21452,N_20813,N_20267);
or U21453 (N_21453,N_20594,N_20897);
and U21454 (N_21454,N_20910,N_19893);
xor U21455 (N_21455,N_20873,N_19878);
and U21456 (N_21456,N_20258,N_20711);
and U21457 (N_21457,N_20640,N_20325);
nor U21458 (N_21458,N_20313,N_20538);
nor U21459 (N_21459,N_19768,N_20193);
or U21460 (N_21460,N_20456,N_20550);
and U21461 (N_21461,N_19676,N_20984);
xnor U21462 (N_21462,N_20092,N_19712);
xnor U21463 (N_21463,N_20120,N_19760);
nand U21464 (N_21464,N_20132,N_19551);
and U21465 (N_21465,N_20187,N_20650);
or U21466 (N_21466,N_20753,N_20657);
and U21467 (N_21467,N_20656,N_20387);
nand U21468 (N_21468,N_20679,N_19643);
nor U21469 (N_21469,N_19793,N_20853);
nand U21470 (N_21470,N_19975,N_19951);
nor U21471 (N_21471,N_20286,N_20573);
nand U21472 (N_21472,N_19927,N_20079);
and U21473 (N_21473,N_20992,N_19897);
xor U21474 (N_21474,N_20791,N_20329);
and U21475 (N_21475,N_20123,N_20600);
and U21476 (N_21476,N_19872,N_20139);
and U21477 (N_21477,N_20760,N_20191);
and U21478 (N_21478,N_20512,N_19573);
nand U21479 (N_21479,N_20089,N_20983);
xnor U21480 (N_21480,N_20220,N_19506);
and U21481 (N_21481,N_20504,N_20879);
and U21482 (N_21482,N_19811,N_20664);
nor U21483 (N_21483,N_19992,N_20868);
xnor U21484 (N_21484,N_19555,N_20714);
xnor U21485 (N_21485,N_20040,N_20215);
or U21486 (N_21486,N_20918,N_20426);
nor U21487 (N_21487,N_19571,N_20971);
nand U21488 (N_21488,N_19663,N_19525);
nand U21489 (N_21489,N_19508,N_19833);
or U21490 (N_21490,N_19981,N_20953);
and U21491 (N_21491,N_20719,N_19546);
nor U21492 (N_21492,N_20596,N_19900);
nor U21493 (N_21493,N_20570,N_19853);
or U21494 (N_21494,N_20699,N_19722);
nor U21495 (N_21495,N_20385,N_19867);
xnor U21496 (N_21496,N_19844,N_20834);
and U21497 (N_21497,N_19757,N_19709);
nand U21498 (N_21498,N_20991,N_20351);
and U21499 (N_21499,N_20051,N_20961);
or U21500 (N_21500,N_20521,N_20086);
xnor U21501 (N_21501,N_19697,N_20476);
xor U21502 (N_21502,N_19800,N_19818);
and U21503 (N_21503,N_20856,N_20061);
nand U21504 (N_21504,N_20068,N_20818);
nor U21505 (N_21505,N_20494,N_19983);
xnor U21506 (N_21506,N_19679,N_20370);
nor U21507 (N_21507,N_19638,N_20378);
or U21508 (N_21508,N_20458,N_20954);
or U21509 (N_21509,N_20196,N_20202);
nor U21510 (N_21510,N_20892,N_19558);
nand U21511 (N_21511,N_20138,N_19720);
nor U21512 (N_21512,N_19766,N_20682);
nand U21513 (N_21513,N_19648,N_20589);
and U21514 (N_21514,N_19756,N_20230);
nor U21515 (N_21515,N_20694,N_20390);
nand U21516 (N_21516,N_19888,N_20309);
nor U21517 (N_21517,N_19785,N_20715);
nor U21518 (N_21518,N_19540,N_20285);
or U21519 (N_21519,N_19923,N_20373);
and U21520 (N_21520,N_19668,N_19851);
or U21521 (N_21521,N_20376,N_20080);
and U21522 (N_21522,N_19895,N_20575);
and U21523 (N_21523,N_20508,N_20332);
nor U21524 (N_21524,N_20626,N_19767);
xnor U21525 (N_21525,N_20468,N_20104);
and U21526 (N_21526,N_19790,N_20555);
and U21527 (N_21527,N_19530,N_20789);
nand U21528 (N_21528,N_19537,N_20413);
nand U21529 (N_21529,N_20588,N_20141);
or U21530 (N_21530,N_20185,N_20361);
nand U21531 (N_21531,N_19609,N_20774);
nor U21532 (N_21532,N_20121,N_20966);
nand U21533 (N_21533,N_20557,N_20236);
or U21534 (N_21534,N_20337,N_19672);
xor U21535 (N_21535,N_19887,N_20349);
or U21536 (N_21536,N_20428,N_20278);
nor U21537 (N_21537,N_20528,N_20857);
and U21538 (N_21538,N_20848,N_20755);
and U21539 (N_21539,N_20975,N_19848);
and U21540 (N_21540,N_19667,N_19693);
and U21541 (N_21541,N_19582,N_19773);
and U21542 (N_21542,N_19628,N_19522);
nor U21543 (N_21543,N_19607,N_20926);
and U21544 (N_21544,N_20223,N_20805);
nand U21545 (N_21545,N_19577,N_19597);
and U21546 (N_21546,N_20997,N_20490);
nor U21547 (N_21547,N_20384,N_19885);
xnor U21548 (N_21548,N_20088,N_20832);
or U21549 (N_21549,N_19613,N_20968);
or U21550 (N_21550,N_20603,N_20680);
nor U21551 (N_21551,N_20059,N_20866);
or U21552 (N_21552,N_20380,N_20686);
or U21553 (N_21553,N_20838,N_19801);
nor U21554 (N_21554,N_20252,N_19935);
and U21555 (N_21555,N_19608,N_20403);
and U21556 (N_21556,N_20784,N_20190);
or U21557 (N_21557,N_20014,N_20747);
and U21558 (N_21558,N_19646,N_19948);
and U21559 (N_21559,N_20438,N_20742);
nor U21560 (N_21560,N_20614,N_20424);
and U21561 (N_21561,N_20116,N_20899);
and U21562 (N_21562,N_20678,N_20035);
nor U21563 (N_21563,N_19879,N_20330);
nand U21564 (N_21564,N_19995,N_19886);
and U21565 (N_21565,N_20405,N_20541);
or U21566 (N_21566,N_20341,N_20020);
nor U21567 (N_21567,N_20167,N_19791);
nor U21568 (N_21568,N_20986,N_20921);
nor U21569 (N_21569,N_19795,N_20269);
xnor U21570 (N_21570,N_19776,N_19978);
xnor U21571 (N_21571,N_20254,N_20814);
nor U21572 (N_21572,N_19592,N_19692);
or U21573 (N_21573,N_20419,N_20863);
or U21574 (N_21574,N_19875,N_20372);
nor U21575 (N_21575,N_20289,N_20605);
xor U21576 (N_21576,N_20641,N_20923);
nand U21577 (N_21577,N_20030,N_20895);
nand U21578 (N_21578,N_20388,N_20128);
and U21579 (N_21579,N_20178,N_19507);
nand U21580 (N_21580,N_20718,N_20987);
or U21581 (N_21581,N_20310,N_19589);
and U21582 (N_21582,N_19907,N_20135);
or U21583 (N_21583,N_20930,N_20238);
or U21584 (N_21584,N_19965,N_20339);
or U21585 (N_21585,N_20047,N_19962);
or U21586 (N_21586,N_20620,N_20151);
nand U21587 (N_21587,N_19727,N_20119);
xnor U21588 (N_21588,N_20281,N_20075);
nand U21589 (N_21589,N_20959,N_20822);
nand U21590 (N_21590,N_20980,N_19634);
and U21591 (N_21591,N_20511,N_20890);
xor U21592 (N_21592,N_20703,N_19856);
nor U21593 (N_21593,N_20783,N_20821);
nand U21594 (N_21594,N_19865,N_20545);
xor U21595 (N_21595,N_19566,N_20294);
or U21596 (N_21596,N_19871,N_19674);
nor U21597 (N_21597,N_20687,N_20969);
or U21598 (N_21598,N_20095,N_20724);
and U21599 (N_21599,N_20737,N_20455);
xnor U21600 (N_21600,N_20593,N_20894);
nor U21601 (N_21601,N_20946,N_20343);
or U21602 (N_21602,N_19725,N_19630);
xor U21603 (N_21603,N_19736,N_20568);
nor U21604 (N_21604,N_20925,N_20427);
xnor U21605 (N_21605,N_20348,N_20155);
nor U21606 (N_21606,N_20367,N_19610);
xnor U21607 (N_21607,N_20524,N_20973);
nand U21608 (N_21608,N_20097,N_20336);
nand U21609 (N_21609,N_20074,N_19991);
nor U21610 (N_21610,N_19994,N_20085);
and U21611 (N_21611,N_20773,N_20083);
nor U21612 (N_21612,N_20396,N_19889);
or U21613 (N_21613,N_19664,N_19775);
xnor U21614 (N_21614,N_20498,N_20915);
nor U21615 (N_21615,N_19626,N_20745);
xnor U21616 (N_21616,N_20425,N_19593);
and U21617 (N_21617,N_19620,N_19590);
or U21618 (N_21618,N_20136,N_20392);
or U21619 (N_21619,N_19937,N_19794);
and U21620 (N_21620,N_20788,N_20027);
or U21621 (N_21621,N_20797,N_19656);
nand U21622 (N_21622,N_20669,N_20347);
or U21623 (N_21623,N_19637,N_19990);
nor U21624 (N_21624,N_20948,N_20268);
nand U21625 (N_21625,N_20194,N_20766);
or U21626 (N_21626,N_20764,N_19734);
or U21627 (N_21627,N_20886,N_20579);
xor U21628 (N_21628,N_20235,N_20491);
nor U21629 (N_21629,N_20500,N_19970);
or U21630 (N_21630,N_20316,N_20655);
nor U21631 (N_21631,N_19836,N_20107);
nand U21632 (N_21632,N_20671,N_20133);
or U21633 (N_21633,N_20015,N_20112);
and U21634 (N_21634,N_19769,N_20793);
and U21635 (N_21635,N_19740,N_20919);
and U21636 (N_21636,N_20906,N_20166);
and U21637 (N_21637,N_19629,N_20041);
nor U21638 (N_21638,N_20412,N_20874);
or U21639 (N_21639,N_20342,N_20544);
xnor U21640 (N_21640,N_19869,N_20021);
nor U21641 (N_21641,N_20861,N_20032);
and U21642 (N_21642,N_20406,N_20338);
xnor U21643 (N_21643,N_20604,N_19840);
xor U21644 (N_21644,N_20101,N_20003);
xor U21645 (N_21645,N_20864,N_20769);
xor U21646 (N_21646,N_19603,N_20826);
nand U21647 (N_21647,N_20621,N_19849);
or U21648 (N_21648,N_19534,N_20449);
or U21649 (N_21649,N_20562,N_20153);
nor U21650 (N_21650,N_19541,N_19623);
nand U21651 (N_21651,N_20261,N_19681);
and U21652 (N_21652,N_20357,N_19834);
or U21653 (N_21653,N_20435,N_20828);
xnor U21654 (N_21654,N_19896,N_20904);
nor U21655 (N_21655,N_19953,N_20693);
nor U21656 (N_21656,N_20584,N_19644);
xor U21657 (N_21657,N_20067,N_20957);
xnor U21658 (N_21658,N_20064,N_20210);
and U21659 (N_21659,N_19596,N_20802);
nor U21660 (N_21660,N_20360,N_20993);
and U21661 (N_21661,N_20761,N_20700);
nor U21662 (N_21662,N_20473,N_20844);
or U21663 (N_21663,N_19731,N_19925);
and U21664 (N_21664,N_19659,N_19891);
nor U21665 (N_21665,N_20256,N_20002);
nand U21666 (N_21666,N_20537,N_19548);
and U21667 (N_21667,N_20019,N_20234);
nor U21668 (N_21668,N_19988,N_20928);
or U21669 (N_21669,N_20778,N_19859);
xor U21670 (N_21670,N_20752,N_20017);
and U21671 (N_21671,N_20319,N_20301);
nor U21672 (N_21672,N_19881,N_19737);
and U21673 (N_21673,N_20847,N_20358);
or U21674 (N_21674,N_20044,N_20214);
nand U21675 (N_21675,N_20398,N_19820);
xnor U21676 (N_21676,N_20441,N_19940);
nand U21677 (N_21677,N_19926,N_20077);
xnor U21678 (N_21678,N_20958,N_20072);
xnor U21679 (N_21679,N_20835,N_19657);
nor U21680 (N_21680,N_20436,N_20212);
or U21681 (N_21681,N_19972,N_19549);
or U21682 (N_21682,N_20340,N_20054);
nand U21683 (N_21683,N_20304,N_20706);
or U21684 (N_21684,N_20677,N_20152);
nand U21685 (N_21685,N_20056,N_19894);
and U21686 (N_21686,N_20423,N_20836);
or U21687 (N_21687,N_19842,N_20590);
and U21688 (N_21688,N_19605,N_20630);
nor U21689 (N_21689,N_20580,N_19877);
nor U21690 (N_21690,N_19514,N_20810);
and U21691 (N_21691,N_20076,N_20697);
or U21692 (N_21692,N_20188,N_19578);
xor U21693 (N_21693,N_19517,N_19738);
and U21694 (N_21694,N_20785,N_20346);
nand U21695 (N_21695,N_20480,N_19944);
or U21696 (N_21696,N_20383,N_19569);
nor U21697 (N_21697,N_20275,N_20365);
nand U21698 (N_21698,N_19742,N_20323);
or U21699 (N_21699,N_20917,N_20263);
or U21700 (N_21700,N_19758,N_19677);
xnor U21701 (N_21701,N_19654,N_19913);
and U21702 (N_21702,N_19862,N_20903);
xor U21703 (N_21703,N_20495,N_20770);
xor U21704 (N_21704,N_20529,N_20115);
or U21705 (N_21705,N_20536,N_20695);
nor U21706 (N_21706,N_20466,N_19945);
xor U21707 (N_21707,N_20862,N_20964);
nor U21708 (N_21708,N_20989,N_19719);
nand U21709 (N_21709,N_20170,N_19691);
xor U21710 (N_21710,N_20939,N_19802);
and U21711 (N_21711,N_20326,N_20912);
xnor U21712 (N_21712,N_19635,N_19559);
nand U21713 (N_21713,N_20619,N_20936);
or U21714 (N_21714,N_20431,N_20225);
and U21715 (N_21715,N_20587,N_20299);
nor U21716 (N_21716,N_20295,N_19539);
nor U21717 (N_21717,N_20156,N_19816);
or U21718 (N_21718,N_19536,N_20757);
and U21719 (N_21719,N_20854,N_20804);
and U21720 (N_21720,N_20898,N_20741);
nand U21721 (N_21721,N_20837,N_19814);
nand U21722 (N_21722,N_20432,N_20739);
nor U21723 (N_21723,N_19511,N_20877);
nand U21724 (N_21724,N_20716,N_19830);
nor U21725 (N_21725,N_19839,N_20534);
and U21726 (N_21726,N_20422,N_19624);
or U21727 (N_21727,N_20606,N_19958);
nor U21728 (N_21728,N_19570,N_20175);
xnor U21729 (N_21729,N_20932,N_19936);
nor U21730 (N_21730,N_19903,N_19666);
xnor U21731 (N_21731,N_19533,N_20914);
nand U21732 (N_21732,N_20486,N_20929);
and U21733 (N_21733,N_20464,N_20736);
and U21734 (N_21734,N_19688,N_19595);
nand U21735 (N_21735,N_20377,N_20247);
and U21736 (N_21736,N_20069,N_20232);
and U21737 (N_21737,N_20842,N_19809);
nand U21738 (N_21738,N_19714,N_20450);
or U21739 (N_21739,N_20882,N_19747);
and U21740 (N_21740,N_19974,N_19617);
or U21741 (N_21741,N_20163,N_20758);
xnor U21742 (N_21742,N_20081,N_19808);
nor U21743 (N_21743,N_20503,N_20927);
nor U21744 (N_21744,N_20598,N_20145);
xor U21745 (N_21745,N_20843,N_19553);
nand U21746 (N_21746,N_20091,N_20595);
or U21747 (N_21747,N_20314,N_19976);
nand U21748 (N_21748,N_20776,N_20250);
nor U21749 (N_21749,N_20627,N_20218);
or U21750 (N_21750,N_20579,N_20735);
and U21751 (N_21751,N_20393,N_20037);
xnor U21752 (N_21752,N_20833,N_19748);
nor U21753 (N_21753,N_20750,N_20504);
xor U21754 (N_21754,N_20406,N_20701);
nand U21755 (N_21755,N_20416,N_20618);
nor U21756 (N_21756,N_20159,N_20025);
and U21757 (N_21757,N_20904,N_19644);
xnor U21758 (N_21758,N_20471,N_20994);
xor U21759 (N_21759,N_20771,N_19909);
nor U21760 (N_21760,N_19899,N_19524);
xnor U21761 (N_21761,N_20542,N_20031);
and U21762 (N_21762,N_20002,N_20890);
xnor U21763 (N_21763,N_20200,N_19596);
xor U21764 (N_21764,N_20902,N_20462);
and U21765 (N_21765,N_20761,N_20638);
and U21766 (N_21766,N_19858,N_19586);
or U21767 (N_21767,N_20813,N_20793);
nor U21768 (N_21768,N_19745,N_20363);
or U21769 (N_21769,N_20628,N_20765);
and U21770 (N_21770,N_20231,N_20382);
nand U21771 (N_21771,N_20020,N_19877);
and U21772 (N_21772,N_19976,N_19571);
or U21773 (N_21773,N_20440,N_20394);
or U21774 (N_21774,N_20020,N_20975);
nor U21775 (N_21775,N_20150,N_20411);
and U21776 (N_21776,N_19960,N_20031);
xor U21777 (N_21777,N_20061,N_20755);
xnor U21778 (N_21778,N_19918,N_20091);
nand U21779 (N_21779,N_19717,N_20358);
nor U21780 (N_21780,N_20356,N_19718);
or U21781 (N_21781,N_20199,N_20482);
nor U21782 (N_21782,N_19796,N_20149);
nand U21783 (N_21783,N_20477,N_20803);
nand U21784 (N_21784,N_19918,N_20760);
nand U21785 (N_21785,N_20134,N_19801);
nor U21786 (N_21786,N_20682,N_19564);
xnor U21787 (N_21787,N_20559,N_20854);
nand U21788 (N_21788,N_19912,N_20888);
nand U21789 (N_21789,N_20290,N_20768);
nand U21790 (N_21790,N_20747,N_20977);
and U21791 (N_21791,N_20995,N_20804);
xnor U21792 (N_21792,N_19555,N_20934);
xnor U21793 (N_21793,N_20431,N_20678);
nor U21794 (N_21794,N_19852,N_20143);
or U21795 (N_21795,N_19533,N_20172);
nand U21796 (N_21796,N_20749,N_20813);
nand U21797 (N_21797,N_20371,N_19808);
and U21798 (N_21798,N_20728,N_19538);
nand U21799 (N_21799,N_19544,N_20982);
or U21800 (N_21800,N_20874,N_19536);
nor U21801 (N_21801,N_19778,N_19695);
nor U21802 (N_21802,N_20270,N_20380);
xnor U21803 (N_21803,N_20483,N_20935);
xor U21804 (N_21804,N_20415,N_20119);
nand U21805 (N_21805,N_20827,N_20044);
nand U21806 (N_21806,N_20585,N_20831);
xor U21807 (N_21807,N_20647,N_20755);
nand U21808 (N_21808,N_20832,N_19967);
and U21809 (N_21809,N_19672,N_19699);
and U21810 (N_21810,N_20861,N_19627);
nor U21811 (N_21811,N_19584,N_20006);
or U21812 (N_21812,N_19549,N_19504);
xor U21813 (N_21813,N_20649,N_20282);
and U21814 (N_21814,N_19524,N_20380);
nand U21815 (N_21815,N_20780,N_20715);
xor U21816 (N_21816,N_20807,N_20922);
or U21817 (N_21817,N_19762,N_20963);
nor U21818 (N_21818,N_20498,N_20962);
and U21819 (N_21819,N_20689,N_20247);
and U21820 (N_21820,N_20075,N_20772);
or U21821 (N_21821,N_20785,N_19786);
and U21822 (N_21822,N_19908,N_20901);
or U21823 (N_21823,N_20658,N_19944);
and U21824 (N_21824,N_20049,N_20855);
xor U21825 (N_21825,N_20275,N_20343);
nor U21826 (N_21826,N_20995,N_20381);
or U21827 (N_21827,N_19993,N_19773);
nand U21828 (N_21828,N_20829,N_20646);
xnor U21829 (N_21829,N_20717,N_19846);
and U21830 (N_21830,N_19598,N_19506);
nand U21831 (N_21831,N_19889,N_20434);
and U21832 (N_21832,N_19653,N_20512);
and U21833 (N_21833,N_19559,N_20869);
nor U21834 (N_21834,N_19969,N_20233);
or U21835 (N_21835,N_20597,N_19846);
xor U21836 (N_21836,N_20126,N_20585);
nand U21837 (N_21837,N_20463,N_20687);
xnor U21838 (N_21838,N_19569,N_20199);
nand U21839 (N_21839,N_20831,N_20187);
xnor U21840 (N_21840,N_19549,N_20846);
xnor U21841 (N_21841,N_19563,N_20214);
and U21842 (N_21842,N_20635,N_20312);
xor U21843 (N_21843,N_20724,N_19972);
nor U21844 (N_21844,N_20381,N_20405);
nand U21845 (N_21845,N_20058,N_19967);
and U21846 (N_21846,N_19824,N_19524);
nor U21847 (N_21847,N_20039,N_20364);
nand U21848 (N_21848,N_19805,N_20823);
or U21849 (N_21849,N_20423,N_20003);
xor U21850 (N_21850,N_20819,N_20051);
nand U21851 (N_21851,N_20997,N_20664);
xor U21852 (N_21852,N_20759,N_20662);
or U21853 (N_21853,N_19938,N_19618);
xnor U21854 (N_21854,N_20610,N_20992);
xor U21855 (N_21855,N_20624,N_19872);
xor U21856 (N_21856,N_20596,N_20013);
and U21857 (N_21857,N_20102,N_19527);
nor U21858 (N_21858,N_20556,N_19580);
xor U21859 (N_21859,N_20254,N_20986);
or U21860 (N_21860,N_19800,N_19833);
xor U21861 (N_21861,N_19947,N_20658);
xor U21862 (N_21862,N_20289,N_20580);
and U21863 (N_21863,N_20162,N_20803);
and U21864 (N_21864,N_20892,N_20121);
or U21865 (N_21865,N_20596,N_19656);
xnor U21866 (N_21866,N_19901,N_20735);
and U21867 (N_21867,N_19622,N_20898);
or U21868 (N_21868,N_20725,N_19559);
xor U21869 (N_21869,N_19783,N_19889);
xnor U21870 (N_21870,N_20250,N_20991);
and U21871 (N_21871,N_20819,N_19565);
nand U21872 (N_21872,N_20368,N_19612);
or U21873 (N_21873,N_20715,N_20250);
and U21874 (N_21874,N_19645,N_19657);
and U21875 (N_21875,N_19692,N_20470);
xnor U21876 (N_21876,N_20458,N_19726);
or U21877 (N_21877,N_20484,N_19841);
and U21878 (N_21878,N_20526,N_20904);
or U21879 (N_21879,N_19836,N_20716);
xor U21880 (N_21880,N_20198,N_19513);
nor U21881 (N_21881,N_20458,N_19866);
xor U21882 (N_21882,N_20818,N_20198);
nand U21883 (N_21883,N_19702,N_20091);
nor U21884 (N_21884,N_20992,N_19857);
nor U21885 (N_21885,N_19710,N_20051);
nor U21886 (N_21886,N_19887,N_19655);
and U21887 (N_21887,N_19506,N_19771);
and U21888 (N_21888,N_20688,N_20236);
nand U21889 (N_21889,N_20910,N_19756);
and U21890 (N_21890,N_20357,N_20607);
nor U21891 (N_21891,N_20256,N_20098);
or U21892 (N_21892,N_19797,N_20075);
nor U21893 (N_21893,N_20119,N_20942);
and U21894 (N_21894,N_20365,N_20732);
and U21895 (N_21895,N_20471,N_20669);
nand U21896 (N_21896,N_20679,N_20630);
xnor U21897 (N_21897,N_20224,N_19568);
xor U21898 (N_21898,N_19693,N_20731);
xor U21899 (N_21899,N_20422,N_19548);
nand U21900 (N_21900,N_20030,N_19896);
and U21901 (N_21901,N_20778,N_20100);
xor U21902 (N_21902,N_20490,N_20235);
nand U21903 (N_21903,N_19745,N_20048);
or U21904 (N_21904,N_19600,N_20508);
and U21905 (N_21905,N_20445,N_19561);
and U21906 (N_21906,N_19590,N_20840);
or U21907 (N_21907,N_20854,N_20565);
xor U21908 (N_21908,N_20545,N_20869);
nor U21909 (N_21909,N_19595,N_19836);
nand U21910 (N_21910,N_20786,N_20885);
nor U21911 (N_21911,N_20987,N_20287);
nor U21912 (N_21912,N_19711,N_20236);
nor U21913 (N_21913,N_20787,N_20973);
or U21914 (N_21914,N_19655,N_20049);
xnor U21915 (N_21915,N_19832,N_20771);
and U21916 (N_21916,N_20577,N_20551);
or U21917 (N_21917,N_19566,N_19920);
and U21918 (N_21918,N_20305,N_20427);
or U21919 (N_21919,N_20273,N_20780);
nand U21920 (N_21920,N_20474,N_20079);
and U21921 (N_21921,N_19635,N_19934);
and U21922 (N_21922,N_20747,N_20598);
or U21923 (N_21923,N_20418,N_20236);
nand U21924 (N_21924,N_20282,N_20075);
xor U21925 (N_21925,N_20192,N_20610);
or U21926 (N_21926,N_20312,N_20516);
and U21927 (N_21927,N_19860,N_19527);
or U21928 (N_21928,N_19852,N_20880);
and U21929 (N_21929,N_20676,N_20097);
xor U21930 (N_21930,N_20580,N_20933);
xor U21931 (N_21931,N_20611,N_19702);
and U21932 (N_21932,N_20054,N_20046);
nand U21933 (N_21933,N_20691,N_19966);
nand U21934 (N_21934,N_20904,N_20262);
nand U21935 (N_21935,N_20268,N_20551);
xnor U21936 (N_21936,N_20469,N_19644);
xor U21937 (N_21937,N_20690,N_19888);
nor U21938 (N_21938,N_19874,N_19683);
nand U21939 (N_21939,N_19555,N_19731);
nand U21940 (N_21940,N_19834,N_20556);
xor U21941 (N_21941,N_20516,N_20372);
and U21942 (N_21942,N_19663,N_20305);
and U21943 (N_21943,N_20032,N_19821);
xnor U21944 (N_21944,N_20294,N_19907);
nand U21945 (N_21945,N_20071,N_20231);
and U21946 (N_21946,N_20875,N_20398);
xnor U21947 (N_21947,N_20567,N_19820);
or U21948 (N_21948,N_20593,N_20356);
and U21949 (N_21949,N_20741,N_20924);
or U21950 (N_21950,N_20820,N_19786);
xnor U21951 (N_21951,N_20890,N_19697);
nor U21952 (N_21952,N_20039,N_19995);
nor U21953 (N_21953,N_20958,N_20723);
and U21954 (N_21954,N_19540,N_20737);
xnor U21955 (N_21955,N_19966,N_20154);
nand U21956 (N_21956,N_20113,N_20723);
nor U21957 (N_21957,N_20234,N_20938);
nor U21958 (N_21958,N_20789,N_19776);
or U21959 (N_21959,N_20438,N_20771);
and U21960 (N_21960,N_19902,N_20257);
nand U21961 (N_21961,N_20089,N_20535);
nor U21962 (N_21962,N_20311,N_19646);
or U21963 (N_21963,N_20110,N_20402);
nor U21964 (N_21964,N_20410,N_19991);
nand U21965 (N_21965,N_20851,N_19634);
and U21966 (N_21966,N_20569,N_19825);
xor U21967 (N_21967,N_20002,N_20857);
nand U21968 (N_21968,N_20721,N_19850);
and U21969 (N_21969,N_19965,N_20797);
or U21970 (N_21970,N_19901,N_20464);
nor U21971 (N_21971,N_20035,N_19641);
or U21972 (N_21972,N_20012,N_19837);
and U21973 (N_21973,N_20986,N_20683);
nand U21974 (N_21974,N_19621,N_20000);
nand U21975 (N_21975,N_20682,N_20300);
and U21976 (N_21976,N_20837,N_19720);
or U21977 (N_21977,N_19971,N_20442);
xor U21978 (N_21978,N_20024,N_20237);
nand U21979 (N_21979,N_19730,N_20540);
and U21980 (N_21980,N_20054,N_19774);
nand U21981 (N_21981,N_20378,N_20304);
nor U21982 (N_21982,N_19548,N_20800);
and U21983 (N_21983,N_20643,N_19639);
and U21984 (N_21984,N_20047,N_20303);
and U21985 (N_21985,N_20063,N_20424);
xnor U21986 (N_21986,N_20375,N_20317);
xor U21987 (N_21987,N_19670,N_20453);
nand U21988 (N_21988,N_19967,N_19842);
nand U21989 (N_21989,N_20049,N_19506);
nand U21990 (N_21990,N_20972,N_19883);
nand U21991 (N_21991,N_19700,N_20549);
or U21992 (N_21992,N_20019,N_19640);
and U21993 (N_21993,N_19929,N_20289);
and U21994 (N_21994,N_20059,N_19819);
and U21995 (N_21995,N_19947,N_20813);
nor U21996 (N_21996,N_19520,N_20655);
nand U21997 (N_21997,N_20109,N_20485);
nand U21998 (N_21998,N_20537,N_19877);
xnor U21999 (N_21999,N_20752,N_20456);
nor U22000 (N_22000,N_20723,N_19567);
xnor U22001 (N_22001,N_20210,N_20141);
nor U22002 (N_22002,N_20167,N_20279);
nor U22003 (N_22003,N_20523,N_20724);
or U22004 (N_22004,N_20985,N_20176);
nand U22005 (N_22005,N_19992,N_19602);
xor U22006 (N_22006,N_19705,N_20004);
nand U22007 (N_22007,N_19807,N_20042);
nor U22008 (N_22008,N_19622,N_19646);
or U22009 (N_22009,N_19897,N_20863);
or U22010 (N_22010,N_20741,N_20828);
or U22011 (N_22011,N_20816,N_19635);
nor U22012 (N_22012,N_20200,N_20039);
nor U22013 (N_22013,N_20981,N_20245);
and U22014 (N_22014,N_20555,N_20119);
xnor U22015 (N_22015,N_20894,N_20386);
nor U22016 (N_22016,N_20460,N_20513);
nor U22017 (N_22017,N_20306,N_19614);
xnor U22018 (N_22018,N_19919,N_19987);
or U22019 (N_22019,N_19864,N_20180);
nor U22020 (N_22020,N_20371,N_20239);
xnor U22021 (N_22021,N_19719,N_20513);
xnor U22022 (N_22022,N_20572,N_19885);
nand U22023 (N_22023,N_20891,N_20183);
and U22024 (N_22024,N_20115,N_19657);
or U22025 (N_22025,N_20424,N_20798);
xor U22026 (N_22026,N_20265,N_20098);
xnor U22027 (N_22027,N_20814,N_20299);
xnor U22028 (N_22028,N_20415,N_19836);
or U22029 (N_22029,N_20149,N_20421);
and U22030 (N_22030,N_20868,N_20728);
and U22031 (N_22031,N_20769,N_20393);
nand U22032 (N_22032,N_20442,N_20461);
or U22033 (N_22033,N_20624,N_19940);
nand U22034 (N_22034,N_20122,N_19866);
and U22035 (N_22035,N_20589,N_19558);
nand U22036 (N_22036,N_20895,N_19551);
nor U22037 (N_22037,N_20218,N_20114);
and U22038 (N_22038,N_20242,N_20396);
and U22039 (N_22039,N_20598,N_19829);
nor U22040 (N_22040,N_19682,N_20687);
xor U22041 (N_22041,N_19792,N_20704);
or U22042 (N_22042,N_20141,N_19678);
nor U22043 (N_22043,N_20097,N_20070);
or U22044 (N_22044,N_20982,N_19920);
nor U22045 (N_22045,N_19802,N_19545);
or U22046 (N_22046,N_20472,N_20352);
xnor U22047 (N_22047,N_19577,N_20379);
nor U22048 (N_22048,N_20062,N_19930);
nor U22049 (N_22049,N_20208,N_19774);
nand U22050 (N_22050,N_20116,N_20285);
or U22051 (N_22051,N_20999,N_20691);
xnor U22052 (N_22052,N_20378,N_19865);
and U22053 (N_22053,N_20860,N_20187);
or U22054 (N_22054,N_20728,N_20978);
nor U22055 (N_22055,N_19941,N_19696);
and U22056 (N_22056,N_20699,N_19584);
xor U22057 (N_22057,N_20585,N_19726);
nand U22058 (N_22058,N_20211,N_19995);
or U22059 (N_22059,N_20120,N_20876);
nand U22060 (N_22060,N_20277,N_19514);
nand U22061 (N_22061,N_19605,N_20359);
xnor U22062 (N_22062,N_20837,N_19554);
xnor U22063 (N_22063,N_20586,N_20202);
and U22064 (N_22064,N_20123,N_20811);
nor U22065 (N_22065,N_20690,N_19525);
or U22066 (N_22066,N_20095,N_20466);
xnor U22067 (N_22067,N_19994,N_20458);
or U22068 (N_22068,N_20502,N_20262);
nand U22069 (N_22069,N_20578,N_20329);
or U22070 (N_22070,N_20936,N_19778);
xor U22071 (N_22071,N_20029,N_19822);
or U22072 (N_22072,N_20232,N_20152);
or U22073 (N_22073,N_19791,N_19771);
xnor U22074 (N_22074,N_20626,N_20324);
and U22075 (N_22075,N_20105,N_20053);
nand U22076 (N_22076,N_20881,N_19634);
and U22077 (N_22077,N_20947,N_20877);
xnor U22078 (N_22078,N_19598,N_20008);
xor U22079 (N_22079,N_20818,N_20165);
or U22080 (N_22080,N_20150,N_20869);
and U22081 (N_22081,N_20158,N_20447);
nand U22082 (N_22082,N_19997,N_20185);
nor U22083 (N_22083,N_19900,N_20582);
and U22084 (N_22084,N_20450,N_20428);
and U22085 (N_22085,N_20860,N_20486);
nor U22086 (N_22086,N_19690,N_20752);
nand U22087 (N_22087,N_20844,N_20239);
nand U22088 (N_22088,N_20529,N_20960);
and U22089 (N_22089,N_19662,N_20048);
nand U22090 (N_22090,N_19583,N_20222);
xnor U22091 (N_22091,N_19992,N_20614);
or U22092 (N_22092,N_20185,N_20388);
and U22093 (N_22093,N_20526,N_19763);
or U22094 (N_22094,N_20774,N_20090);
nand U22095 (N_22095,N_19719,N_19635);
xor U22096 (N_22096,N_20683,N_20732);
or U22097 (N_22097,N_19594,N_20772);
and U22098 (N_22098,N_19724,N_20288);
xnor U22099 (N_22099,N_20796,N_19780);
and U22100 (N_22100,N_20790,N_20162);
or U22101 (N_22101,N_20123,N_20242);
or U22102 (N_22102,N_20207,N_20539);
nand U22103 (N_22103,N_20451,N_20110);
and U22104 (N_22104,N_19814,N_20522);
and U22105 (N_22105,N_19561,N_20550);
xor U22106 (N_22106,N_20601,N_19701);
xnor U22107 (N_22107,N_20309,N_20693);
or U22108 (N_22108,N_20510,N_20639);
nor U22109 (N_22109,N_20807,N_20717);
xor U22110 (N_22110,N_20418,N_19508);
xnor U22111 (N_22111,N_19703,N_19501);
or U22112 (N_22112,N_20461,N_19930);
xor U22113 (N_22113,N_19896,N_20354);
nor U22114 (N_22114,N_20941,N_20374);
or U22115 (N_22115,N_19753,N_19566);
xor U22116 (N_22116,N_20770,N_20834);
nand U22117 (N_22117,N_20350,N_20975);
and U22118 (N_22118,N_20031,N_19720);
or U22119 (N_22119,N_20027,N_20897);
or U22120 (N_22120,N_20536,N_19535);
nand U22121 (N_22121,N_20985,N_20635);
nand U22122 (N_22122,N_20783,N_19814);
nor U22123 (N_22123,N_20094,N_19570);
or U22124 (N_22124,N_19718,N_20121);
or U22125 (N_22125,N_20954,N_20049);
nand U22126 (N_22126,N_20300,N_20559);
or U22127 (N_22127,N_19651,N_19546);
nand U22128 (N_22128,N_19869,N_20517);
nand U22129 (N_22129,N_20647,N_19979);
xor U22130 (N_22130,N_20014,N_19935);
nor U22131 (N_22131,N_20536,N_19795);
nand U22132 (N_22132,N_20679,N_20293);
nand U22133 (N_22133,N_20650,N_20074);
nand U22134 (N_22134,N_19990,N_20688);
nor U22135 (N_22135,N_20790,N_20148);
nor U22136 (N_22136,N_20121,N_20076);
and U22137 (N_22137,N_20401,N_19523);
or U22138 (N_22138,N_19905,N_20502);
or U22139 (N_22139,N_20288,N_20773);
xor U22140 (N_22140,N_20627,N_19931);
nor U22141 (N_22141,N_20769,N_20541);
nand U22142 (N_22142,N_19867,N_20855);
nand U22143 (N_22143,N_20414,N_19513);
and U22144 (N_22144,N_19612,N_20780);
xnor U22145 (N_22145,N_20348,N_20744);
or U22146 (N_22146,N_20382,N_20618);
or U22147 (N_22147,N_19708,N_20364);
nor U22148 (N_22148,N_19880,N_19835);
or U22149 (N_22149,N_20582,N_20448);
and U22150 (N_22150,N_20575,N_19628);
nor U22151 (N_22151,N_19587,N_20254);
and U22152 (N_22152,N_20123,N_20553);
nor U22153 (N_22153,N_20579,N_19706);
xnor U22154 (N_22154,N_20156,N_19609);
xnor U22155 (N_22155,N_19715,N_20715);
nand U22156 (N_22156,N_19835,N_20851);
and U22157 (N_22157,N_20312,N_20964);
nor U22158 (N_22158,N_19942,N_19941);
nor U22159 (N_22159,N_20810,N_20731);
or U22160 (N_22160,N_20638,N_20350);
xor U22161 (N_22161,N_20854,N_20968);
xnor U22162 (N_22162,N_19552,N_19795);
nand U22163 (N_22163,N_20657,N_19710);
xnor U22164 (N_22164,N_20726,N_20638);
xnor U22165 (N_22165,N_19826,N_20558);
or U22166 (N_22166,N_20583,N_20438);
and U22167 (N_22167,N_20323,N_20095);
or U22168 (N_22168,N_20898,N_20639);
or U22169 (N_22169,N_20084,N_19601);
nand U22170 (N_22170,N_20433,N_19658);
nand U22171 (N_22171,N_20059,N_20936);
or U22172 (N_22172,N_20948,N_20352);
xor U22173 (N_22173,N_19528,N_19998);
and U22174 (N_22174,N_20392,N_20311);
nor U22175 (N_22175,N_20728,N_20270);
xnor U22176 (N_22176,N_19859,N_19745);
nand U22177 (N_22177,N_20239,N_20944);
xnor U22178 (N_22178,N_20638,N_19935);
nand U22179 (N_22179,N_20811,N_20075);
and U22180 (N_22180,N_20673,N_20293);
nor U22181 (N_22181,N_20516,N_20665);
nor U22182 (N_22182,N_20661,N_20671);
or U22183 (N_22183,N_20716,N_20953);
nor U22184 (N_22184,N_20844,N_20939);
xnor U22185 (N_22185,N_19926,N_19889);
nor U22186 (N_22186,N_19598,N_20905);
and U22187 (N_22187,N_19986,N_20826);
nor U22188 (N_22188,N_20460,N_20325);
nor U22189 (N_22189,N_20895,N_20170);
or U22190 (N_22190,N_19734,N_20470);
or U22191 (N_22191,N_20140,N_20124);
and U22192 (N_22192,N_20069,N_20490);
xnor U22193 (N_22193,N_19805,N_19905);
xnor U22194 (N_22194,N_20373,N_19604);
nor U22195 (N_22195,N_20079,N_20169);
and U22196 (N_22196,N_19750,N_20892);
nand U22197 (N_22197,N_19690,N_19835);
and U22198 (N_22198,N_20557,N_19527);
and U22199 (N_22199,N_20680,N_19819);
nand U22200 (N_22200,N_19568,N_20552);
nand U22201 (N_22201,N_20792,N_19962);
nand U22202 (N_22202,N_19964,N_19981);
nor U22203 (N_22203,N_19849,N_20400);
xnor U22204 (N_22204,N_20504,N_20820);
or U22205 (N_22205,N_20097,N_20040);
or U22206 (N_22206,N_20474,N_19934);
and U22207 (N_22207,N_19867,N_20839);
and U22208 (N_22208,N_19595,N_20033);
xnor U22209 (N_22209,N_19804,N_20910);
xnor U22210 (N_22210,N_20065,N_20818);
nand U22211 (N_22211,N_20210,N_20084);
xnor U22212 (N_22212,N_20016,N_20833);
nand U22213 (N_22213,N_20143,N_20724);
nor U22214 (N_22214,N_20376,N_20257);
or U22215 (N_22215,N_20403,N_20437);
nor U22216 (N_22216,N_20595,N_20925);
or U22217 (N_22217,N_20574,N_19618);
xnor U22218 (N_22218,N_19759,N_20662);
nor U22219 (N_22219,N_20160,N_20929);
xnor U22220 (N_22220,N_19988,N_20274);
nand U22221 (N_22221,N_20240,N_20540);
xnor U22222 (N_22222,N_20751,N_19964);
nor U22223 (N_22223,N_20088,N_20785);
nor U22224 (N_22224,N_19904,N_19735);
or U22225 (N_22225,N_20576,N_19927);
xor U22226 (N_22226,N_19905,N_20609);
nand U22227 (N_22227,N_19804,N_20621);
or U22228 (N_22228,N_20475,N_19854);
nor U22229 (N_22229,N_20767,N_20934);
nor U22230 (N_22230,N_20133,N_20009);
and U22231 (N_22231,N_19722,N_20857);
and U22232 (N_22232,N_20733,N_20661);
xor U22233 (N_22233,N_19902,N_20785);
xor U22234 (N_22234,N_20820,N_19969);
nor U22235 (N_22235,N_20522,N_20598);
nor U22236 (N_22236,N_20797,N_19629);
nand U22237 (N_22237,N_20590,N_20148);
or U22238 (N_22238,N_20001,N_20604);
or U22239 (N_22239,N_20674,N_20876);
and U22240 (N_22240,N_19813,N_20007);
xnor U22241 (N_22241,N_20101,N_20830);
or U22242 (N_22242,N_20260,N_20969);
nor U22243 (N_22243,N_20830,N_20121);
or U22244 (N_22244,N_20252,N_20837);
xnor U22245 (N_22245,N_19689,N_20904);
xnor U22246 (N_22246,N_20874,N_20171);
and U22247 (N_22247,N_19872,N_19648);
xor U22248 (N_22248,N_20103,N_20524);
and U22249 (N_22249,N_19687,N_20598);
and U22250 (N_22250,N_20380,N_20140);
nand U22251 (N_22251,N_19563,N_20027);
nand U22252 (N_22252,N_20160,N_19741);
xnor U22253 (N_22253,N_19823,N_20333);
or U22254 (N_22254,N_19769,N_19884);
xnor U22255 (N_22255,N_19611,N_19836);
nand U22256 (N_22256,N_19507,N_20096);
xor U22257 (N_22257,N_20698,N_20980);
or U22258 (N_22258,N_19739,N_20811);
and U22259 (N_22259,N_19763,N_20841);
nor U22260 (N_22260,N_20501,N_20289);
xor U22261 (N_22261,N_20098,N_19541);
nand U22262 (N_22262,N_20346,N_20550);
nor U22263 (N_22263,N_20641,N_20865);
or U22264 (N_22264,N_20214,N_20957);
xor U22265 (N_22265,N_20049,N_19885);
nor U22266 (N_22266,N_20559,N_20102);
nor U22267 (N_22267,N_20421,N_19698);
xor U22268 (N_22268,N_20528,N_19712);
and U22269 (N_22269,N_20148,N_20802);
or U22270 (N_22270,N_19656,N_20921);
nand U22271 (N_22271,N_20505,N_20519);
and U22272 (N_22272,N_20970,N_19705);
and U22273 (N_22273,N_19875,N_20152);
or U22274 (N_22274,N_19988,N_19962);
and U22275 (N_22275,N_19615,N_20860);
nand U22276 (N_22276,N_20609,N_19812);
nand U22277 (N_22277,N_19561,N_20980);
nand U22278 (N_22278,N_20245,N_20920);
nand U22279 (N_22279,N_20315,N_19848);
or U22280 (N_22280,N_20703,N_20720);
or U22281 (N_22281,N_19657,N_20227);
xnor U22282 (N_22282,N_19686,N_20869);
nor U22283 (N_22283,N_19635,N_20791);
and U22284 (N_22284,N_20426,N_20714);
nor U22285 (N_22285,N_20701,N_20061);
nor U22286 (N_22286,N_20053,N_20359);
xnor U22287 (N_22287,N_19827,N_20401);
nor U22288 (N_22288,N_19732,N_20442);
nor U22289 (N_22289,N_20931,N_20852);
and U22290 (N_22290,N_20214,N_20458);
and U22291 (N_22291,N_20744,N_20148);
or U22292 (N_22292,N_20712,N_20279);
and U22293 (N_22293,N_20657,N_19618);
nand U22294 (N_22294,N_20752,N_20723);
xor U22295 (N_22295,N_19796,N_20389);
nand U22296 (N_22296,N_20043,N_20044);
xor U22297 (N_22297,N_20677,N_20452);
or U22298 (N_22298,N_20218,N_20448);
or U22299 (N_22299,N_20767,N_19709);
xor U22300 (N_22300,N_19755,N_20753);
nand U22301 (N_22301,N_20651,N_19798);
nand U22302 (N_22302,N_20406,N_19988);
and U22303 (N_22303,N_20640,N_20487);
nor U22304 (N_22304,N_19889,N_20938);
nand U22305 (N_22305,N_20116,N_19926);
and U22306 (N_22306,N_20761,N_20121);
and U22307 (N_22307,N_20967,N_20397);
xor U22308 (N_22308,N_20136,N_20054);
nor U22309 (N_22309,N_20915,N_19582);
nand U22310 (N_22310,N_19778,N_20486);
xnor U22311 (N_22311,N_20373,N_19820);
nor U22312 (N_22312,N_20098,N_19811);
nand U22313 (N_22313,N_19855,N_20577);
xor U22314 (N_22314,N_20595,N_20568);
or U22315 (N_22315,N_20845,N_19760);
or U22316 (N_22316,N_20138,N_19995);
xor U22317 (N_22317,N_19573,N_20807);
or U22318 (N_22318,N_20294,N_19982);
and U22319 (N_22319,N_19605,N_20117);
and U22320 (N_22320,N_20720,N_19729);
xor U22321 (N_22321,N_20067,N_20821);
or U22322 (N_22322,N_20525,N_19796);
nand U22323 (N_22323,N_20196,N_19630);
xnor U22324 (N_22324,N_19910,N_19542);
and U22325 (N_22325,N_19923,N_20334);
xor U22326 (N_22326,N_20354,N_20641);
or U22327 (N_22327,N_20041,N_20951);
nor U22328 (N_22328,N_20101,N_20787);
or U22329 (N_22329,N_19730,N_19721);
nor U22330 (N_22330,N_19581,N_20834);
nor U22331 (N_22331,N_20730,N_20057);
nor U22332 (N_22332,N_20208,N_19678);
nor U22333 (N_22333,N_20535,N_19673);
nand U22334 (N_22334,N_19784,N_20965);
xor U22335 (N_22335,N_20861,N_20053);
xor U22336 (N_22336,N_20478,N_20569);
nor U22337 (N_22337,N_20891,N_20359);
and U22338 (N_22338,N_19891,N_20167);
nand U22339 (N_22339,N_20489,N_20013);
nor U22340 (N_22340,N_19775,N_19692);
nor U22341 (N_22341,N_20604,N_20148);
and U22342 (N_22342,N_20136,N_20315);
nor U22343 (N_22343,N_20483,N_19960);
xnor U22344 (N_22344,N_19511,N_20147);
and U22345 (N_22345,N_20683,N_20974);
xnor U22346 (N_22346,N_20316,N_20109);
nand U22347 (N_22347,N_20711,N_19758);
xor U22348 (N_22348,N_19634,N_20660);
and U22349 (N_22349,N_20066,N_20018);
xor U22350 (N_22350,N_20040,N_20037);
nor U22351 (N_22351,N_19942,N_19724);
or U22352 (N_22352,N_20746,N_19983);
xor U22353 (N_22353,N_20837,N_19931);
nand U22354 (N_22354,N_19737,N_19893);
and U22355 (N_22355,N_20165,N_20920);
xor U22356 (N_22356,N_19581,N_20343);
or U22357 (N_22357,N_20046,N_20471);
or U22358 (N_22358,N_20968,N_20824);
nand U22359 (N_22359,N_20455,N_20779);
nor U22360 (N_22360,N_20530,N_20573);
nand U22361 (N_22361,N_20595,N_20839);
or U22362 (N_22362,N_19660,N_20195);
and U22363 (N_22363,N_20216,N_20566);
and U22364 (N_22364,N_20655,N_20446);
or U22365 (N_22365,N_20725,N_19842);
and U22366 (N_22366,N_19957,N_20349);
or U22367 (N_22367,N_19533,N_19860);
nor U22368 (N_22368,N_20943,N_20867);
nor U22369 (N_22369,N_19971,N_20223);
or U22370 (N_22370,N_20823,N_19577);
nand U22371 (N_22371,N_20852,N_20374);
xnor U22372 (N_22372,N_20558,N_20079);
nand U22373 (N_22373,N_19627,N_19785);
nand U22374 (N_22374,N_20301,N_20124);
xor U22375 (N_22375,N_20477,N_20998);
nand U22376 (N_22376,N_20942,N_20806);
or U22377 (N_22377,N_20876,N_20534);
nor U22378 (N_22378,N_20413,N_20159);
nor U22379 (N_22379,N_19823,N_19583);
nand U22380 (N_22380,N_20549,N_20440);
or U22381 (N_22381,N_20774,N_20088);
nor U22382 (N_22382,N_20412,N_20925);
nand U22383 (N_22383,N_20558,N_19612);
or U22384 (N_22384,N_20973,N_20960);
nand U22385 (N_22385,N_19912,N_20384);
nor U22386 (N_22386,N_19660,N_20887);
nand U22387 (N_22387,N_20912,N_19591);
nor U22388 (N_22388,N_19570,N_19981);
nand U22389 (N_22389,N_20152,N_19980);
and U22390 (N_22390,N_20964,N_19985);
and U22391 (N_22391,N_20040,N_20776);
and U22392 (N_22392,N_19818,N_19847);
nand U22393 (N_22393,N_20310,N_20834);
and U22394 (N_22394,N_19883,N_20684);
nor U22395 (N_22395,N_19616,N_20559);
nor U22396 (N_22396,N_19964,N_20632);
and U22397 (N_22397,N_20864,N_20745);
nand U22398 (N_22398,N_20247,N_20485);
or U22399 (N_22399,N_19740,N_19917);
or U22400 (N_22400,N_20209,N_19676);
nand U22401 (N_22401,N_20684,N_20511);
or U22402 (N_22402,N_19857,N_20690);
and U22403 (N_22403,N_19586,N_19783);
nor U22404 (N_22404,N_19890,N_19543);
and U22405 (N_22405,N_20330,N_19693);
and U22406 (N_22406,N_20614,N_19714);
nand U22407 (N_22407,N_20437,N_19912);
nand U22408 (N_22408,N_20344,N_19926);
and U22409 (N_22409,N_20596,N_19608);
xor U22410 (N_22410,N_19929,N_20036);
nor U22411 (N_22411,N_19581,N_19555);
or U22412 (N_22412,N_20245,N_20086);
xnor U22413 (N_22413,N_20447,N_20267);
or U22414 (N_22414,N_20062,N_19740);
or U22415 (N_22415,N_19510,N_20587);
or U22416 (N_22416,N_19704,N_20296);
xor U22417 (N_22417,N_20229,N_20765);
xor U22418 (N_22418,N_20449,N_20443);
xnor U22419 (N_22419,N_20531,N_20639);
or U22420 (N_22420,N_19938,N_20547);
xor U22421 (N_22421,N_20259,N_20256);
nor U22422 (N_22422,N_19908,N_19842);
nor U22423 (N_22423,N_20877,N_20583);
nand U22424 (N_22424,N_20314,N_20107);
xor U22425 (N_22425,N_19634,N_20871);
or U22426 (N_22426,N_20294,N_20253);
xnor U22427 (N_22427,N_20688,N_19596);
or U22428 (N_22428,N_20741,N_20464);
and U22429 (N_22429,N_19550,N_20625);
xnor U22430 (N_22430,N_20868,N_20415);
and U22431 (N_22431,N_20755,N_20419);
or U22432 (N_22432,N_19874,N_19775);
xnor U22433 (N_22433,N_20522,N_20721);
and U22434 (N_22434,N_20000,N_19894);
or U22435 (N_22435,N_20484,N_20102);
and U22436 (N_22436,N_19836,N_20190);
nand U22437 (N_22437,N_20842,N_20349);
xor U22438 (N_22438,N_20301,N_19951);
or U22439 (N_22439,N_19589,N_20804);
and U22440 (N_22440,N_19551,N_19913);
and U22441 (N_22441,N_19661,N_20186);
and U22442 (N_22442,N_20563,N_20024);
and U22443 (N_22443,N_20672,N_20324);
nor U22444 (N_22444,N_19674,N_20030);
xor U22445 (N_22445,N_19622,N_20806);
or U22446 (N_22446,N_19550,N_19747);
and U22447 (N_22447,N_20925,N_20018);
xnor U22448 (N_22448,N_20623,N_20284);
or U22449 (N_22449,N_20368,N_20873);
nand U22450 (N_22450,N_19557,N_19752);
nor U22451 (N_22451,N_19930,N_20827);
or U22452 (N_22452,N_20410,N_20686);
and U22453 (N_22453,N_19719,N_19864);
and U22454 (N_22454,N_20108,N_19929);
nand U22455 (N_22455,N_20286,N_20009);
xor U22456 (N_22456,N_20428,N_20284);
nor U22457 (N_22457,N_20810,N_20940);
xor U22458 (N_22458,N_20535,N_19681);
or U22459 (N_22459,N_20277,N_20822);
xor U22460 (N_22460,N_19921,N_20783);
nand U22461 (N_22461,N_20875,N_19689);
and U22462 (N_22462,N_20798,N_20256);
and U22463 (N_22463,N_20115,N_20884);
nand U22464 (N_22464,N_19528,N_20940);
nor U22465 (N_22465,N_19642,N_20925);
nor U22466 (N_22466,N_19582,N_19879);
nand U22467 (N_22467,N_20093,N_20191);
or U22468 (N_22468,N_20618,N_19648);
and U22469 (N_22469,N_19868,N_20405);
nand U22470 (N_22470,N_20807,N_20177);
nand U22471 (N_22471,N_19756,N_20240);
nor U22472 (N_22472,N_20036,N_20853);
nor U22473 (N_22473,N_20928,N_19606);
nor U22474 (N_22474,N_20268,N_20487);
xor U22475 (N_22475,N_19927,N_19768);
nand U22476 (N_22476,N_20036,N_20570);
xor U22477 (N_22477,N_20063,N_20105);
nor U22478 (N_22478,N_19615,N_20143);
xnor U22479 (N_22479,N_19974,N_20683);
nor U22480 (N_22480,N_20504,N_20314);
nand U22481 (N_22481,N_20179,N_19580);
xnor U22482 (N_22482,N_19844,N_19945);
nand U22483 (N_22483,N_20126,N_19773);
or U22484 (N_22484,N_20753,N_20796);
or U22485 (N_22485,N_20755,N_20958);
xor U22486 (N_22486,N_20436,N_20257);
and U22487 (N_22487,N_20332,N_20609);
and U22488 (N_22488,N_20340,N_19693);
and U22489 (N_22489,N_20526,N_20837);
nand U22490 (N_22490,N_20345,N_19564);
nor U22491 (N_22491,N_20087,N_19804);
xor U22492 (N_22492,N_20018,N_20627);
nor U22493 (N_22493,N_20983,N_20066);
and U22494 (N_22494,N_19518,N_20235);
nand U22495 (N_22495,N_19732,N_20370);
nand U22496 (N_22496,N_20851,N_19547);
xnor U22497 (N_22497,N_20347,N_20438);
nor U22498 (N_22498,N_20940,N_20302);
xor U22499 (N_22499,N_19609,N_19926);
and U22500 (N_22500,N_22014,N_21945);
nand U22501 (N_22501,N_22084,N_21274);
xnor U22502 (N_22502,N_21229,N_21898);
and U22503 (N_22503,N_22331,N_21070);
or U22504 (N_22504,N_22309,N_21913);
and U22505 (N_22505,N_22289,N_21656);
or U22506 (N_22506,N_21414,N_21153);
or U22507 (N_22507,N_21046,N_21341);
and U22508 (N_22508,N_22157,N_22235);
nand U22509 (N_22509,N_22301,N_22418);
xnor U22510 (N_22510,N_21822,N_21935);
or U22511 (N_22511,N_21937,N_21757);
nor U22512 (N_22512,N_21402,N_21977);
xnor U22513 (N_22513,N_21396,N_21230);
nand U22514 (N_22514,N_21421,N_22112);
or U22515 (N_22515,N_22120,N_22404);
nor U22516 (N_22516,N_21487,N_21296);
nor U22517 (N_22517,N_21813,N_22079);
and U22518 (N_22518,N_21451,N_22060);
or U22519 (N_22519,N_21874,N_21731);
nand U22520 (N_22520,N_21654,N_21835);
nand U22521 (N_22521,N_22270,N_22127);
nand U22522 (N_22522,N_21009,N_22197);
nor U22523 (N_22523,N_22124,N_21792);
or U22524 (N_22524,N_22493,N_21307);
or U22525 (N_22525,N_21132,N_21083);
nand U22526 (N_22526,N_21418,N_22058);
xor U22527 (N_22527,N_21351,N_21071);
xnor U22528 (N_22528,N_21392,N_22129);
or U22529 (N_22529,N_21957,N_21056);
nor U22530 (N_22530,N_22241,N_21265);
or U22531 (N_22531,N_21773,N_21767);
nor U22532 (N_22532,N_21859,N_22009);
nand U22533 (N_22533,N_21380,N_22366);
nor U22534 (N_22534,N_22462,N_21171);
nor U22535 (N_22535,N_21799,N_21616);
and U22536 (N_22536,N_21725,N_21238);
nor U22537 (N_22537,N_21466,N_21002);
nor U22538 (N_22538,N_21247,N_21457);
xor U22539 (N_22539,N_22134,N_22170);
nor U22540 (N_22540,N_22487,N_21869);
xnor U22541 (N_22541,N_21320,N_22393);
and U22542 (N_22542,N_22162,N_22072);
xnor U22543 (N_22543,N_21377,N_21497);
nand U22544 (N_22544,N_22065,N_21409);
xnor U22545 (N_22545,N_22490,N_21806);
nand U22546 (N_22546,N_22022,N_21493);
xnor U22547 (N_22547,N_21729,N_21615);
xnor U22548 (N_22548,N_21355,N_21161);
or U22549 (N_22549,N_21867,N_21375);
or U22550 (N_22550,N_22423,N_22086);
xor U22551 (N_22551,N_21033,N_21860);
and U22552 (N_22552,N_22242,N_21478);
xor U22553 (N_22553,N_22210,N_22122);
xnor U22554 (N_22554,N_21820,N_21257);
xnor U22555 (N_22555,N_21653,N_21304);
and U22556 (N_22556,N_22095,N_21048);
nand U22557 (N_22557,N_22481,N_22427);
and U22558 (N_22558,N_22406,N_21105);
nand U22559 (N_22559,N_21743,N_21988);
or U22560 (N_22560,N_21079,N_21199);
xor U22561 (N_22561,N_21761,N_22254);
nor U22562 (N_22562,N_22051,N_21872);
and U22563 (N_22563,N_21469,N_22165);
xnor U22564 (N_22564,N_21192,N_21796);
nor U22565 (N_22565,N_22221,N_22004);
and U22566 (N_22566,N_21917,N_22128);
xor U22567 (N_22567,N_22078,N_22391);
or U22568 (N_22568,N_21410,N_22488);
and U22569 (N_22569,N_21144,N_21603);
nor U22570 (N_22570,N_22410,N_21017);
and U22571 (N_22571,N_21170,N_22377);
and U22572 (N_22572,N_21815,N_22230);
nand U22573 (N_22573,N_21186,N_22277);
nor U22574 (N_22574,N_21148,N_22327);
nand U22575 (N_22575,N_21805,N_21899);
xnor U22576 (N_22576,N_21774,N_22355);
nor U22577 (N_22577,N_21004,N_22190);
nor U22578 (N_22578,N_21811,N_21183);
nor U22579 (N_22579,N_22364,N_21962);
xnor U22580 (N_22580,N_22042,N_21188);
nor U22581 (N_22581,N_21042,N_21116);
xnor U22582 (N_22582,N_22397,N_21102);
nand U22583 (N_22583,N_22139,N_22275);
nand U22584 (N_22584,N_22040,N_21467);
and U22585 (N_22585,N_21456,N_22010);
nor U22586 (N_22586,N_22224,N_21007);
or U22587 (N_22587,N_21617,N_21034);
nor U22588 (N_22588,N_22117,N_21135);
xor U22589 (N_22589,N_22192,N_21736);
xnor U22590 (N_22590,N_22185,N_21700);
nand U22591 (N_22591,N_22193,N_21583);
xnor U22592 (N_22592,N_21692,N_21190);
and U22593 (N_22593,N_21018,N_21709);
nor U22594 (N_22594,N_22362,N_21400);
or U22595 (N_22595,N_21673,N_21342);
nor U22596 (N_22596,N_22181,N_21185);
and U22597 (N_22597,N_21240,N_22343);
nand U22598 (N_22598,N_22253,N_22283);
nor U22599 (N_22599,N_22274,N_22297);
xor U22600 (N_22600,N_21947,N_22325);
nor U22601 (N_22601,N_22153,N_21831);
or U22602 (N_22602,N_21424,N_21006);
or U22603 (N_22603,N_21726,N_21756);
nand U22604 (N_22604,N_22286,N_21950);
nand U22605 (N_22605,N_21152,N_21889);
and U22606 (N_22606,N_21722,N_21043);
nand U22607 (N_22607,N_21300,N_21140);
or U22608 (N_22608,N_21775,N_21597);
nor U22609 (N_22609,N_21781,N_22195);
xnor U22610 (N_22610,N_22482,N_21050);
nor U22611 (N_22611,N_21293,N_22172);
xnor U22612 (N_22612,N_21430,N_22345);
or U22613 (N_22613,N_21809,N_21463);
and U22614 (N_22614,N_22083,N_22308);
or U22615 (N_22615,N_21481,N_21302);
and U22616 (N_22616,N_21376,N_21718);
nor U22617 (N_22617,N_21339,N_21585);
and U22618 (N_22618,N_21398,N_22202);
or U22619 (N_22619,N_21219,N_22282);
and U22620 (N_22620,N_21028,N_21552);
nand U22621 (N_22621,N_22166,N_22432);
nor U22622 (N_22622,N_21504,N_21911);
or U22623 (N_22623,N_22233,N_21233);
and U22624 (N_22624,N_22350,N_21882);
xnor U22625 (N_22625,N_21411,N_22480);
nor U22626 (N_22626,N_22285,N_21172);
and U22627 (N_22627,N_22085,N_21836);
or U22628 (N_22628,N_21747,N_21139);
nand U22629 (N_22629,N_21429,N_21667);
or U22630 (N_22630,N_21470,N_22217);
or U22631 (N_22631,N_21156,N_22243);
nand U22632 (N_22632,N_21714,N_22461);
nand U22633 (N_22633,N_22413,N_22476);
and U22634 (N_22634,N_22104,N_22118);
or U22635 (N_22635,N_22305,N_21124);
or U22636 (N_22636,N_22464,N_21203);
xnor U22637 (N_22637,N_21143,N_21543);
xnor U22638 (N_22638,N_21989,N_22492);
nor U22639 (N_22639,N_22002,N_22215);
xor U22640 (N_22640,N_22407,N_21884);
nor U22641 (N_22641,N_22473,N_22451);
and U22642 (N_22642,N_22332,N_21569);
nor U22643 (N_22643,N_21561,N_22045);
xnor U22644 (N_22644,N_22211,N_21854);
nor U22645 (N_22645,N_21574,N_22069);
xnor U22646 (N_22646,N_21225,N_22005);
nand U22647 (N_22647,N_21605,N_22319);
and U22648 (N_22648,N_21448,N_22059);
nor U22649 (N_22649,N_22110,N_21657);
and U22650 (N_22650,N_21089,N_21178);
nand U22651 (N_22651,N_22115,N_22373);
nand U22652 (N_22652,N_21348,N_21968);
xnor U22653 (N_22653,N_21489,N_21754);
xnor U22654 (N_22654,N_22213,N_22191);
xnor U22655 (N_22655,N_22329,N_22357);
xor U22656 (N_22656,N_21146,N_22347);
xor U22657 (N_22657,N_22425,N_21189);
and U22658 (N_22658,N_21613,N_21983);
nand U22659 (N_22659,N_21092,N_21906);
nand U22660 (N_22660,N_21516,N_21534);
nand U22661 (N_22661,N_21630,N_22074);
and U22662 (N_22662,N_22416,N_21591);
xnor U22663 (N_22663,N_21313,N_21999);
nor U22664 (N_22664,N_21829,N_22394);
or U22665 (N_22665,N_21408,N_21084);
xnor U22666 (N_22666,N_21104,N_21220);
xnor U22667 (N_22667,N_22026,N_21498);
nor U22668 (N_22668,N_21059,N_21031);
nor U22669 (N_22669,N_22499,N_21024);
nor U22670 (N_22670,N_21310,N_22278);
or U22671 (N_22671,N_22483,N_22370);
and U22672 (N_22672,N_22453,N_22312);
and U22673 (N_22673,N_21912,N_21929);
and U22674 (N_22674,N_22189,N_21560);
or U22675 (N_22675,N_21519,N_21758);
nor U22676 (N_22676,N_22314,N_21741);
nor U22677 (N_22677,N_21705,N_22379);
and U22678 (N_22678,N_21938,N_21373);
xnor U22679 (N_22679,N_21579,N_22265);
and U22680 (N_22680,N_21287,N_22471);
nor U22681 (N_22681,N_22137,N_21795);
nand U22682 (N_22682,N_21788,N_21282);
or U22683 (N_22683,N_22175,N_22164);
or U22684 (N_22684,N_21998,N_21627);
and U22685 (N_22685,N_21057,N_22096);
nor U22686 (N_22686,N_21010,N_21475);
nor U22687 (N_22687,N_21520,N_22152);
xnor U22688 (N_22688,N_21594,N_21900);
nor U22689 (N_22689,N_21312,N_21821);
nand U22690 (N_22690,N_21800,N_22342);
or U22691 (N_22691,N_21191,N_22150);
nor U22692 (N_22692,N_21604,N_21733);
or U22693 (N_22693,N_21541,N_21096);
nor U22694 (N_22694,N_21039,N_21802);
xnor U22695 (N_22695,N_21350,N_21068);
and U22696 (N_22696,N_22489,N_22204);
or U22697 (N_22697,N_22234,N_21971);
or U22698 (N_22698,N_21555,N_21281);
and U22699 (N_22699,N_21345,N_21224);
and U22700 (N_22700,N_22299,N_22032);
nand U22701 (N_22701,N_22114,N_21868);
nand U22702 (N_22702,N_21887,N_21112);
and U22703 (N_22703,N_21445,N_21918);
nor U22704 (N_22704,N_21122,N_22087);
or U22705 (N_22705,N_21369,N_21526);
nand U22706 (N_22706,N_21215,N_22439);
or U22707 (N_22707,N_22417,N_21633);
and U22708 (N_22708,N_21846,N_21787);
xnor U22709 (N_22709,N_21259,N_21590);
nand U22710 (N_22710,N_21069,N_21683);
or U22711 (N_22711,N_21054,N_22419);
nand U22712 (N_22712,N_22392,N_22269);
xor U22713 (N_22713,N_22454,N_21194);
nor U22714 (N_22714,N_21058,N_21213);
nor U22715 (N_22715,N_22428,N_21208);
xnor U22716 (N_22716,N_21471,N_21209);
or U22717 (N_22717,N_22020,N_21063);
and U22718 (N_22718,N_21082,N_21405);
nand U22719 (N_22719,N_22006,N_21381);
and U22720 (N_22720,N_21299,N_21676);
and U22721 (N_22721,N_21542,N_21494);
and U22722 (N_22722,N_21367,N_21165);
or U22723 (N_22723,N_21349,N_21746);
or U22724 (N_22724,N_21027,N_22380);
or U22725 (N_22725,N_21234,N_21468);
xnor U22726 (N_22726,N_21385,N_22315);
nor U22727 (N_22727,N_21991,N_21511);
or U22728 (N_22728,N_21187,N_22238);
xor U22729 (N_22729,N_21557,N_21324);
or U22730 (N_22730,N_21528,N_21205);
and U22731 (N_22731,N_22361,N_22446);
and U22732 (N_22732,N_22207,N_22160);
nor U22733 (N_22733,N_21672,N_21707);
nor U22734 (N_22734,N_21765,N_21986);
nor U22735 (N_22735,N_21360,N_21883);
and U22736 (N_22736,N_21087,N_21180);
nand U22737 (N_22737,N_22280,N_21308);
xnor U22738 (N_22738,N_21588,N_22457);
and U22739 (N_22739,N_21567,N_22386);
xor U22740 (N_22740,N_22363,N_21828);
nand U22741 (N_22741,N_21173,N_21055);
nand U22742 (N_22742,N_22352,N_21242);
and U22743 (N_22743,N_21272,N_21825);
nand U22744 (N_22744,N_21982,N_21625);
or U22745 (N_22745,N_21618,N_21249);
xnor U22746 (N_22746,N_22307,N_21515);
and U22747 (N_22747,N_22222,N_22173);
xor U22748 (N_22748,N_21608,N_21704);
nor U22749 (N_22749,N_21842,N_21535);
nand U22750 (N_22750,N_22463,N_22216);
or U22751 (N_22751,N_21640,N_21362);
or U22752 (N_22752,N_22316,N_21159);
or U22753 (N_22753,N_21587,N_21479);
or U22754 (N_22754,N_22113,N_22030);
nor U22755 (N_22755,N_22293,N_21782);
nand U22756 (N_22756,N_21580,N_21446);
nand U22757 (N_22757,N_21064,N_21720);
xor U22758 (N_22758,N_21881,N_22247);
or U22759 (N_22759,N_21323,N_22376);
nand U22760 (N_22760,N_21931,N_22123);
nor U22761 (N_22761,N_21916,N_21995);
nor U22762 (N_22762,N_21202,N_21635);
nor U22763 (N_22763,N_21897,N_21217);
and U22764 (N_22764,N_21636,N_21706);
xnor U22765 (N_22765,N_21568,N_22318);
nand U22766 (N_22766,N_21357,N_21131);
or U22767 (N_22767,N_21563,N_21093);
xnor U22768 (N_22768,N_22107,N_21910);
nand U22769 (N_22769,N_22082,N_22437);
nor U22770 (N_22770,N_22184,N_21698);
nand U22771 (N_22771,N_22016,N_21125);
nor U22772 (N_22772,N_21067,N_21920);
nor U22773 (N_22773,N_21793,N_21334);
xnor U22774 (N_22774,N_22146,N_21877);
or U22775 (N_22775,N_22323,N_21227);
xor U22776 (N_22776,N_22449,N_21346);
nor U22777 (N_22777,N_22174,N_21168);
nand U22778 (N_22778,N_22047,N_22475);
nor U22779 (N_22779,N_21776,N_21008);
or U22780 (N_22780,N_21386,N_21699);
and U22781 (N_22781,N_21040,N_21644);
xnor U22782 (N_22782,N_21309,N_21892);
nor U22783 (N_22783,N_21110,N_21975);
or U22784 (N_22784,N_21888,N_21674);
nor U22785 (N_22785,N_21065,N_21849);
nor U22786 (N_22786,N_21974,N_21981);
or U22787 (N_22787,N_22106,N_21539);
or U22788 (N_22788,N_21517,N_21894);
or U22789 (N_22789,N_22205,N_21181);
and U22790 (N_22790,N_22132,N_21919);
xor U22791 (N_22791,N_21319,N_21701);
or U22792 (N_22792,N_21325,N_21129);
xnor U22793 (N_22793,N_22034,N_21136);
nor U22794 (N_22794,N_21669,N_21091);
xor U22795 (N_22795,N_21648,N_22149);
nand U22796 (N_22796,N_22039,N_21368);
nor U22797 (N_22797,N_21602,N_21160);
or U22798 (N_22798,N_21717,N_22264);
nand U22799 (N_22799,N_22321,N_21830);
nor U22800 (N_22800,N_21810,N_21435);
nor U22801 (N_22801,N_22103,N_21306);
xnor U22802 (N_22802,N_21374,N_21510);
xnor U22803 (N_22803,N_21314,N_21562);
and U22804 (N_22804,N_21531,N_22421);
nand U22805 (N_22805,N_21508,N_22431);
nand U22806 (N_22806,N_21730,N_22338);
nand U22807 (N_22807,N_22458,N_22187);
or U22808 (N_22808,N_21544,N_22249);
or U22809 (N_22809,N_21942,N_21291);
xnor U22810 (N_22810,N_21719,N_21123);
or U22811 (N_22811,N_21262,N_21907);
nand U22812 (N_22812,N_21275,N_21384);
nor U22813 (N_22813,N_21934,N_22186);
nand U22814 (N_22814,N_21958,N_21990);
nand U22815 (N_22815,N_21663,N_22426);
nand U22816 (N_22816,N_21575,N_21204);
xor U22817 (N_22817,N_21426,N_21780);
and U22818 (N_22818,N_22294,N_22262);
nand U22819 (N_22819,N_21394,N_21847);
nor U22820 (N_22820,N_22029,N_21823);
nor U22821 (N_22821,N_21915,N_21382);
and U22822 (N_22822,N_21465,N_22231);
nand U22823 (N_22823,N_21014,N_21485);
xnor U22824 (N_22824,N_22339,N_21791);
nand U22825 (N_22825,N_21764,N_21099);
nand U22826 (N_22826,N_21026,N_22024);
nor U22827 (N_22827,N_21826,N_22161);
xnor U22828 (N_22828,N_22050,N_21851);
or U22829 (N_22829,N_21570,N_22271);
nand U22830 (N_22830,N_22148,N_21151);
or U22831 (N_22831,N_21248,N_22220);
xor U22832 (N_22832,N_21413,N_21062);
nand U22833 (N_22833,N_22390,N_21984);
or U22834 (N_22834,N_21670,N_21537);
nor U22835 (N_22835,N_21979,N_21529);
and U22836 (N_22836,N_22344,N_21344);
and U22837 (N_22837,N_21378,N_21436);
or U22838 (N_22838,N_21101,N_21598);
or U22839 (N_22839,N_22227,N_21666);
or U22840 (N_22840,N_22182,N_22310);
xnor U22841 (N_22841,N_22300,N_21294);
xor U22842 (N_22842,N_22239,N_21556);
xnor U22843 (N_22843,N_22317,N_21253);
or U22844 (N_22844,N_21970,N_22424);
and U22845 (N_22845,N_22302,N_21558);
nand U22846 (N_22846,N_21843,N_21108);
and U22847 (N_22847,N_21525,N_22018);
or U22848 (N_22848,N_21121,N_22025);
or U22849 (N_22849,N_21861,N_21439);
and U22850 (N_22850,N_22011,N_21162);
nand U22851 (N_22851,N_22374,N_21922);
nand U22852 (N_22852,N_21474,N_21130);
or U22853 (N_22853,N_21280,N_22142);
or U22854 (N_22854,N_21629,N_21496);
xnor U22855 (N_22855,N_21295,N_22260);
or U22856 (N_22856,N_21075,N_22133);
xor U22857 (N_22857,N_21284,N_22469);
nor U22858 (N_22858,N_21154,N_21246);
or U22859 (N_22859,N_22441,N_21985);
xnor U22860 (N_22860,N_21315,N_21679);
or U22861 (N_22861,N_21438,N_22466);
and U22862 (N_22862,N_21174,N_22346);
nor U22863 (N_22863,N_22036,N_22281);
nand U22864 (N_22864,N_22007,N_22266);
nand U22865 (N_22865,N_21210,N_21878);
nor U22866 (N_22866,N_22445,N_21716);
xnor U22867 (N_22867,N_22093,N_22111);
and U22868 (N_22868,N_21255,N_22219);
nand U22869 (N_22869,N_21850,N_21972);
xor U22870 (N_22870,N_21682,N_21283);
xnor U22871 (N_22871,N_22395,N_22402);
or U22872 (N_22872,N_21524,N_21715);
and U22873 (N_22873,N_22396,N_21417);
or U22874 (N_22874,N_21459,N_21030);
and U22875 (N_22875,N_21997,N_21029);
nand U22876 (N_22876,N_21643,N_21862);
xor U22877 (N_22877,N_22015,N_21290);
xor U22878 (N_22878,N_22056,N_22420);
and U22879 (N_22879,N_21752,N_22077);
xor U22880 (N_22880,N_21880,N_21444);
xor U22881 (N_22881,N_22336,N_21383);
nand U22882 (N_22882,N_21514,N_21954);
nand U22883 (N_22883,N_22369,N_21814);
and U22884 (N_22884,N_22375,N_21966);
nand U22885 (N_22885,N_21532,N_21266);
nor U22886 (N_22886,N_22183,N_21708);
and U22887 (N_22887,N_21097,N_22066);
nand U22888 (N_22888,N_22470,N_22322);
or U22889 (N_22889,N_21100,N_21292);
and U22890 (N_22890,N_21777,N_21495);
or U22891 (N_22891,N_22141,N_22348);
nor U22892 (N_22892,N_22491,N_22102);
nor U22893 (N_22893,N_21818,N_21856);
or U22894 (N_22894,N_21755,N_21582);
xor U22895 (N_22895,N_21036,N_21372);
xnor U22896 (N_22896,N_22000,N_21166);
nand U22897 (N_22897,N_21371,N_22048);
or U22898 (N_22898,N_21354,N_21379);
nand U22899 (N_22899,N_21216,N_21571);
and U22900 (N_22900,N_22276,N_21025);
nor U22901 (N_22901,N_21370,N_21412);
and U22902 (N_22902,N_21335,N_22223);
xnor U22903 (N_22903,N_21019,N_22090);
xor U22904 (N_22904,N_22138,N_21576);
nor U22905 (N_22905,N_21994,N_21322);
and U22906 (N_22906,N_21020,N_21804);
xor U22907 (N_22907,N_21047,N_21142);
xor U22908 (N_22908,N_21505,N_21852);
or U22909 (N_22909,N_22163,N_21694);
nand U22910 (N_22910,N_21901,N_21232);
and U22911 (N_22911,N_22236,N_22267);
or U22912 (N_22912,N_21458,N_21509);
xnor U22913 (N_22913,N_21228,N_22468);
or U22914 (N_22914,N_21768,N_21483);
xor U22915 (N_22915,N_21035,N_21993);
nor U22916 (N_22916,N_21549,N_21401);
or U22917 (N_22917,N_22169,N_21518);
and U22918 (N_22918,N_21407,N_21477);
nor U22919 (N_22919,N_21023,N_22126);
nand U22920 (N_22920,N_22268,N_21462);
nor U22921 (N_22921,N_21267,N_21614);
xor U22922 (N_22922,N_22349,N_21326);
or U22923 (N_22923,N_21642,N_21158);
or U22924 (N_22924,N_21455,N_21737);
nor U22925 (N_22925,N_21713,N_22447);
nand U22926 (N_22926,N_22028,N_21789);
xor U22927 (N_22927,N_22038,N_22387);
nor U22928 (N_22928,N_21797,N_21858);
nor U22929 (N_22929,N_21432,N_21428);
and U22930 (N_22930,N_21661,N_22304);
and U22931 (N_22931,N_21236,N_21041);
nand U22932 (N_22932,N_22360,N_22388);
and U22933 (N_22933,N_21053,N_22245);
xnor U22934 (N_22934,N_21783,N_22291);
nor U22935 (N_22935,N_21573,N_22044);
xor U22936 (N_22936,N_21645,N_21660);
and U22937 (N_22937,N_21211,N_21536);
nand U22938 (N_22938,N_22201,N_21337);
nand U22939 (N_22939,N_21677,N_21359);
nor U22940 (N_22940,N_21179,N_21316);
nand U22941 (N_22941,N_21712,N_21786);
nor U22942 (N_22942,N_22237,N_21440);
and U22943 (N_22943,N_21288,N_21651);
nand U22944 (N_22944,N_22177,N_22131);
nand U22945 (N_22945,N_22119,N_22429);
nor U22946 (N_22946,N_21081,N_21925);
and U22947 (N_22947,N_22443,N_21620);
nor U22948 (N_22948,N_21052,N_21641);
xnor U22949 (N_22949,N_22405,N_21619);
and U22950 (N_22950,N_21329,N_21447);
xnor U22951 (N_22951,N_21689,N_21697);
or U22952 (N_22952,N_21460,N_21550);
nor U22953 (N_22953,N_22328,N_21927);
or U22954 (N_22954,N_21857,N_21032);
nand U22955 (N_22955,N_22013,N_21564);
and U22956 (N_22956,N_21269,N_22337);
nor U22957 (N_22957,N_21688,N_22168);
nor U22958 (N_22958,N_21317,N_21824);
or U22959 (N_22959,N_22228,N_21976);
nand U22960 (N_22960,N_21244,N_22214);
or U22961 (N_22961,N_21581,N_21512);
xor U22962 (N_22962,N_21655,N_21119);
nand U22963 (N_22963,N_21596,N_21749);
and U22964 (N_22964,N_22412,N_21461);
and U22965 (N_22965,N_21270,N_21578);
nand U22966 (N_22966,N_21903,N_22498);
and U22967 (N_22967,N_21453,N_21632);
nor U22968 (N_22968,N_21637,N_22340);
or U22969 (N_22969,N_21352,N_21926);
nand U22970 (N_22970,N_21303,N_21488);
and U22971 (N_22971,N_21013,N_21703);
xor U22972 (N_22972,N_22250,N_21696);
nand U22973 (N_22973,N_21239,N_21452);
nor U22974 (N_22974,N_22341,N_22415);
or U22975 (N_22975,N_22143,N_22444);
nor U22976 (N_22976,N_22023,N_22372);
nand U22977 (N_22977,N_22135,N_21671);
and U22978 (N_22978,N_21521,N_21431);
xnor U22979 (N_22979,N_21784,N_21340);
nor U22980 (N_22980,N_22151,N_22094);
nor U22981 (N_22981,N_22017,N_22306);
nor U22982 (N_22982,N_21120,N_21330);
xor U22983 (N_22983,N_21904,N_22144);
nor U22984 (N_22984,N_21527,N_21675);
nand U22985 (N_22985,N_22229,N_21951);
and U22986 (N_22986,N_21870,N_21328);
and U22987 (N_22987,N_22176,N_21338);
and U22988 (N_22988,N_21650,N_21134);
xor U22989 (N_22989,N_21473,N_22433);
nand U22990 (N_22990,N_22246,N_21164);
or U22991 (N_22991,N_21502,N_21252);
or U22992 (N_22992,N_21422,N_21658);
nor U22993 (N_22993,N_21946,N_22460);
and U22994 (N_22994,N_21114,N_22261);
or U22995 (N_22995,N_22455,N_21808);
xor U22996 (N_22996,N_21533,N_21647);
xor U22997 (N_22997,N_21996,N_22031);
or U22998 (N_22998,N_21623,N_22368);
nand U22999 (N_22999,N_21790,N_21949);
xnor U23000 (N_23000,N_21832,N_21289);
or U23001 (N_23001,N_21664,N_21197);
and U23002 (N_23002,N_21060,N_21298);
nand U23003 (N_23003,N_22465,N_21769);
nand U23004 (N_23004,N_21141,N_21837);
nand U23005 (N_23005,N_21223,N_21710);
and U23006 (N_23006,N_21522,N_21109);
xnor U23007 (N_23007,N_22244,N_22292);
or U23008 (N_23008,N_21163,N_22097);
nor U23009 (N_23009,N_21840,N_21546);
or U23010 (N_23010,N_21589,N_21798);
nor U23011 (N_23011,N_22452,N_21566);
nor U23012 (N_23012,N_22434,N_21763);
and U23013 (N_23013,N_21254,N_21639);
and U23014 (N_23014,N_21218,N_22259);
nor U23015 (N_23015,N_22384,N_22430);
nor U23016 (N_23016,N_21628,N_21005);
nand U23017 (N_23017,N_22442,N_22046);
xor U23018 (N_23018,N_22284,N_21921);
nor U23019 (N_23019,N_21003,N_21486);
and U23020 (N_23020,N_21437,N_22334);
xnor U23021 (N_23021,N_22288,N_22158);
nor U23022 (N_23022,N_21175,N_21049);
or U23023 (N_23023,N_21115,N_21772);
nor U23024 (N_23024,N_22440,N_21126);
or U23025 (N_23025,N_21871,N_22479);
or U23026 (N_23026,N_21690,N_21364);
or U23027 (N_23027,N_22061,N_21554);
nor U23028 (N_23028,N_21638,N_22062);
nor U23029 (N_23029,N_22092,N_22171);
nand U23030 (N_23030,N_22448,N_21356);
xnor U23031 (N_23031,N_22240,N_22188);
nand U23032 (N_23032,N_21169,N_22478);
nor U23033 (N_23033,N_22088,N_21149);
nor U23034 (N_23034,N_21212,N_22091);
or U23035 (N_23035,N_21095,N_21250);
nor U23036 (N_23036,N_22203,N_22212);
or U23037 (N_23037,N_21948,N_21037);
xor U23038 (N_23038,N_21078,N_22035);
nor U23039 (N_23039,N_22330,N_22287);
or U23040 (N_23040,N_21548,N_21622);
nand U23041 (N_23041,N_21779,N_21932);
nand U23042 (N_23042,N_21530,N_21610);
xnor U23043 (N_23043,N_21021,N_22037);
xor U23044 (N_23044,N_21200,N_21484);
or U23045 (N_23045,N_21902,N_21965);
nand U23046 (N_23046,N_21914,N_21875);
nand U23047 (N_23047,N_21001,N_22198);
nor U23048 (N_23048,N_22075,N_21363);
nor U23049 (N_23049,N_21311,N_22400);
and U23050 (N_23050,N_21702,N_21955);
or U23051 (N_23051,N_21941,N_22196);
nor U23052 (N_23052,N_22248,N_21404);
nand U23053 (N_23053,N_21833,N_22450);
nand U23054 (N_23054,N_22382,N_21523);
nor U23055 (N_23055,N_21397,N_22279);
nor U23056 (N_23056,N_21133,N_21973);
and U23057 (N_23057,N_21612,N_21157);
and U23058 (N_23058,N_21118,N_21321);
nor U23059 (N_23059,N_21624,N_21893);
and U23060 (N_23060,N_21506,N_21753);
nor U23061 (N_23061,N_21182,N_21358);
xor U23062 (N_23062,N_21540,N_21751);
xor U23063 (N_23063,N_21011,N_21442);
nor U23064 (N_23064,N_21454,N_21387);
xnor U23065 (N_23065,N_22383,N_21425);
xnor U23066 (N_23066,N_21685,N_22206);
or U23067 (N_23067,N_22226,N_21538);
or U23068 (N_23068,N_21305,N_21553);
nor U23069 (N_23069,N_22358,N_21198);
nand U23070 (N_23070,N_21665,N_21155);
or U23071 (N_23071,N_21953,N_21336);
nand U23072 (N_23072,N_22435,N_22414);
xnor U23073 (N_23073,N_21201,N_22258);
xnor U23074 (N_23074,N_21952,N_21406);
xnor U23075 (N_23075,N_21472,N_21176);
nor U23076 (N_23076,N_21727,N_22486);
and U23077 (N_23077,N_21268,N_22178);
and U23078 (N_23078,N_21419,N_21061);
nand U23079 (N_23079,N_21207,N_21853);
or U23080 (N_23080,N_21739,N_21278);
nor U23081 (N_23081,N_21251,N_21128);
nand U23082 (N_23082,N_21593,N_22365);
and U23083 (N_23083,N_21886,N_22167);
nor U23084 (N_23084,N_22313,N_22467);
or U23085 (N_23085,N_21841,N_22296);
nand U23086 (N_23086,N_21908,N_21361);
and U23087 (N_23087,N_21492,N_21817);
nor U23088 (N_23088,N_21490,N_21865);
nor U23089 (N_23089,N_21879,N_21801);
or U23090 (N_23090,N_22200,N_21332);
and U23091 (N_23091,N_21885,N_22012);
nand U23092 (N_23092,N_21891,N_22459);
xor U23093 (N_23093,N_21347,N_22477);
and U23094 (N_23094,N_22105,N_22008);
or U23095 (N_23095,N_21184,N_21681);
xor U23096 (N_23096,N_21264,N_22311);
nand U23097 (N_23097,N_21331,N_21662);
and U23098 (N_23098,N_21545,N_21038);
or U23099 (N_23099,N_21551,N_21678);
nand U23100 (N_23100,N_21606,N_22081);
and U23101 (N_23101,N_22257,N_21480);
xnor U23102 (N_23102,N_22218,N_21450);
or U23103 (N_23103,N_22073,N_22180);
xnor U23104 (N_23104,N_22411,N_22385);
xnor U23105 (N_23105,N_21415,N_21000);
xnor U23106 (N_23106,N_21770,N_22256);
nand U23107 (N_23107,N_22130,N_21735);
xnor U23108 (N_23108,N_21077,N_21167);
and U23109 (N_23109,N_21177,N_22080);
or U23110 (N_23110,N_21241,N_22495);
or U23111 (N_23111,N_21838,N_21482);
or U23112 (N_23112,N_21085,N_21195);
xnor U23113 (N_23113,N_22367,N_22147);
nand U23114 (N_23114,N_21012,N_21864);
xnor U23115 (N_23115,N_21193,N_22354);
and U23116 (N_23116,N_22389,N_22076);
nand U23117 (N_23117,N_21127,N_21206);
or U23118 (N_23118,N_22068,N_22089);
nand U23119 (N_23119,N_21066,N_21601);
and U23120 (N_23120,N_21956,N_21343);
nand U23121 (N_23121,N_21072,N_21626);
or U23122 (N_23122,N_22403,N_21819);
and U23123 (N_23123,N_21812,N_21734);
nor U23124 (N_23124,N_21592,N_21113);
nand U23125 (N_23125,N_22136,N_21609);
or U23126 (N_23126,N_22438,N_21992);
nor U23127 (N_23127,N_22033,N_21117);
nor U23128 (N_23128,N_21366,N_22179);
nand U23129 (N_23129,N_22101,N_21045);
or U23130 (N_23130,N_22108,N_22273);
or U23131 (N_23131,N_21258,N_21723);
and U23132 (N_23132,N_22409,N_22053);
xnor U23133 (N_23133,N_21607,N_21924);
xor U23134 (N_23134,N_21276,N_22326);
nor U23135 (N_23135,N_21427,N_22494);
and U23136 (N_23136,N_22333,N_22021);
and U23137 (N_23137,N_22335,N_21742);
and U23138 (N_23138,N_22067,N_22485);
nor U23139 (N_23139,N_22295,N_21214);
nor U23140 (N_23140,N_22496,N_22252);
nor U23141 (N_23141,N_22255,N_21231);
nand U23142 (N_23142,N_21353,N_22381);
nand U23143 (N_23143,N_22378,N_21221);
nor U23144 (N_23144,N_22027,N_21086);
nor U23145 (N_23145,N_21391,N_22140);
xor U23146 (N_23146,N_21740,N_21111);
and U23147 (N_23147,N_21476,N_21441);
xnor U23148 (N_23148,N_21297,N_21138);
nor U23149 (N_23149,N_21940,N_22063);
nand U23150 (N_23150,N_21855,N_22001);
or U23151 (N_23151,N_21235,N_21577);
xor U23152 (N_23152,N_21744,N_21695);
xor U23153 (N_23153,N_21711,N_21762);
or U23154 (N_23154,N_21978,N_21611);
and U23155 (N_23155,N_22057,N_21076);
nand U23156 (N_23156,N_21649,N_21277);
nor U23157 (N_23157,N_21245,N_22054);
xnor U23158 (N_23158,N_22194,N_22098);
nor U23159 (N_23159,N_21390,N_22351);
nor U23160 (N_23160,N_21987,N_22399);
nand U23161 (N_23161,N_21106,N_21260);
and U23162 (N_23162,N_22298,N_21261);
xor U23163 (N_23163,N_21890,N_21684);
nand U23164 (N_23164,N_21500,N_21016);
xnor U23165 (N_23165,N_21301,N_22070);
nand U23166 (N_23166,N_21074,N_21222);
nand U23167 (N_23167,N_21226,N_21073);
nor U23168 (N_23168,N_21286,N_21866);
xor U23169 (N_23169,N_22303,N_21848);
nor U23170 (N_23170,N_21909,N_22251);
xor U23171 (N_23171,N_21327,N_21631);
or U23172 (N_23172,N_21464,N_21333);
or U23173 (N_23173,N_22116,N_21963);
and U23174 (N_23174,N_21449,N_21961);
xnor U23175 (N_23175,N_21559,N_22422);
nor U23176 (N_23176,N_21403,N_21967);
nand U23177 (N_23177,N_21271,N_22125);
or U23178 (N_23178,N_21876,N_22272);
nand U23179 (N_23179,N_21724,N_21691);
xnor U23180 (N_23180,N_21565,N_21621);
and U23181 (N_23181,N_21423,N_21863);
nand U23182 (N_23182,N_22497,N_21845);
nor U23183 (N_23183,N_21807,N_21732);
and U23184 (N_23184,N_21959,N_22145);
nor U23185 (N_23185,N_21895,N_21365);
nor U23186 (N_23186,N_21745,N_21051);
xnor U23187 (N_23187,N_21771,N_21964);
and U23188 (N_23188,N_21513,N_21933);
nand U23189 (N_23189,N_21443,N_21243);
nand U23190 (N_23190,N_21196,N_21766);
and U23191 (N_23191,N_21094,N_22159);
and U23192 (N_23192,N_21547,N_22232);
and U23193 (N_23193,N_22019,N_22100);
xnor U23194 (N_23194,N_22154,N_22401);
or U23195 (N_23195,N_21399,N_22456);
nand U23196 (N_23196,N_21839,N_22208);
xor U23197 (N_23197,N_21044,N_21652);
nor U23198 (N_23198,N_21646,N_21750);
and U23199 (N_23199,N_22155,N_21090);
nor U23200 (N_23200,N_22225,N_21728);
and U23201 (N_23201,N_21969,N_22064);
nor U23202 (N_23202,N_21015,N_21939);
and U23203 (N_23203,N_22003,N_22041);
nor U23204 (N_23204,N_22290,N_21600);
and U23205 (N_23205,N_21668,N_21263);
nand U23206 (N_23206,N_21503,N_22356);
nor U23207 (N_23207,N_22209,N_21572);
xor U23208 (N_23208,N_21137,N_21107);
nor U23209 (N_23209,N_21905,N_21944);
nand U23210 (N_23210,N_22353,N_21103);
and U23211 (N_23211,N_22324,N_21395);
nand U23212 (N_23212,N_22052,N_22408);
or U23213 (N_23213,N_21686,N_22398);
xor U23214 (N_23214,N_21433,N_21960);
or U23215 (N_23215,N_21759,N_22320);
or U23216 (N_23216,N_21389,N_21586);
xnor U23217 (N_23217,N_21659,N_22121);
xor U23218 (N_23218,N_22199,N_21693);
nor U23219 (N_23219,N_21816,N_21595);
or U23220 (N_23220,N_21098,N_22055);
or U23221 (N_23221,N_21794,N_21022);
or U23222 (N_23222,N_21318,N_21584);
nand U23223 (N_23223,N_22109,N_22071);
nand U23224 (N_23224,N_22474,N_21420);
and U23225 (N_23225,N_21237,N_21980);
and U23226 (N_23226,N_22371,N_21634);
nand U23227 (N_23227,N_21680,N_22263);
and U23228 (N_23228,N_21803,N_21687);
xor U23229 (N_23229,N_21416,N_21088);
nand U23230 (N_23230,N_21491,N_21285);
nor U23231 (N_23231,N_21273,N_22049);
xnor U23232 (N_23232,N_22156,N_22359);
xor U23233 (N_23233,N_21279,N_21145);
nor U23234 (N_23234,N_22472,N_21501);
xnor U23235 (N_23235,N_21499,N_21507);
and U23236 (N_23236,N_22484,N_21748);
nor U23237 (N_23237,N_21393,N_21873);
nand U23238 (N_23238,N_21943,N_21827);
or U23239 (N_23239,N_21923,N_21896);
or U23240 (N_23240,N_21080,N_21150);
nand U23241 (N_23241,N_21738,N_21721);
nor U23242 (N_23242,N_21785,N_22043);
xor U23243 (N_23243,N_22436,N_21928);
xor U23244 (N_23244,N_21930,N_21599);
nor U23245 (N_23245,N_21388,N_21434);
or U23246 (N_23246,N_21778,N_21147);
and U23247 (N_23247,N_21834,N_22099);
and U23248 (N_23248,N_21936,N_21760);
or U23249 (N_23249,N_21844,N_21256);
and U23250 (N_23250,N_22398,N_22198);
or U23251 (N_23251,N_21358,N_22098);
xor U23252 (N_23252,N_22057,N_21629);
and U23253 (N_23253,N_22376,N_21577);
and U23254 (N_23254,N_22132,N_21377);
or U23255 (N_23255,N_21855,N_21334);
or U23256 (N_23256,N_22461,N_21081);
or U23257 (N_23257,N_22118,N_21234);
or U23258 (N_23258,N_21942,N_22330);
xor U23259 (N_23259,N_21420,N_22285);
nor U23260 (N_23260,N_22016,N_21842);
and U23261 (N_23261,N_22149,N_21491);
or U23262 (N_23262,N_22468,N_21252);
xor U23263 (N_23263,N_21192,N_21078);
and U23264 (N_23264,N_21896,N_21581);
or U23265 (N_23265,N_22497,N_21581);
xnor U23266 (N_23266,N_21322,N_21525);
xnor U23267 (N_23267,N_22175,N_21463);
nor U23268 (N_23268,N_21487,N_21705);
and U23269 (N_23269,N_21774,N_21068);
or U23270 (N_23270,N_21243,N_21368);
or U23271 (N_23271,N_21299,N_22112);
xor U23272 (N_23272,N_21307,N_21917);
xnor U23273 (N_23273,N_21400,N_21619);
nand U23274 (N_23274,N_21295,N_21200);
nor U23275 (N_23275,N_21206,N_22166);
xnor U23276 (N_23276,N_21504,N_21316);
nand U23277 (N_23277,N_21496,N_21941);
xnor U23278 (N_23278,N_21038,N_22164);
and U23279 (N_23279,N_21364,N_22212);
xnor U23280 (N_23280,N_22435,N_21273);
xnor U23281 (N_23281,N_21318,N_21930);
nand U23282 (N_23282,N_21145,N_22396);
nand U23283 (N_23283,N_22344,N_22280);
and U23284 (N_23284,N_22304,N_21261);
nand U23285 (N_23285,N_22355,N_22186);
nand U23286 (N_23286,N_21410,N_21692);
nor U23287 (N_23287,N_21760,N_22437);
nand U23288 (N_23288,N_21783,N_22031);
nand U23289 (N_23289,N_21691,N_21392);
nand U23290 (N_23290,N_22149,N_21745);
nor U23291 (N_23291,N_21574,N_22470);
or U23292 (N_23292,N_21427,N_22006);
and U23293 (N_23293,N_22199,N_21940);
nor U23294 (N_23294,N_21082,N_21732);
nor U23295 (N_23295,N_21167,N_22391);
xor U23296 (N_23296,N_21244,N_21893);
xnor U23297 (N_23297,N_21172,N_21037);
and U23298 (N_23298,N_22394,N_22408);
xnor U23299 (N_23299,N_21690,N_21904);
nand U23300 (N_23300,N_22352,N_22346);
or U23301 (N_23301,N_21597,N_21664);
xnor U23302 (N_23302,N_21744,N_21502);
and U23303 (N_23303,N_22280,N_21372);
nand U23304 (N_23304,N_22077,N_21695);
or U23305 (N_23305,N_21655,N_21039);
and U23306 (N_23306,N_22309,N_22154);
nand U23307 (N_23307,N_22119,N_21619);
nand U23308 (N_23308,N_21264,N_21479);
and U23309 (N_23309,N_21246,N_21810);
nor U23310 (N_23310,N_21251,N_21967);
nor U23311 (N_23311,N_21561,N_22017);
and U23312 (N_23312,N_22439,N_21608);
nor U23313 (N_23313,N_22342,N_22058);
nand U23314 (N_23314,N_21315,N_22267);
and U23315 (N_23315,N_21966,N_22075);
xnor U23316 (N_23316,N_21645,N_22341);
nand U23317 (N_23317,N_21831,N_21800);
nor U23318 (N_23318,N_21166,N_21075);
nor U23319 (N_23319,N_21753,N_21019);
nor U23320 (N_23320,N_21664,N_21356);
nor U23321 (N_23321,N_22487,N_21488);
xnor U23322 (N_23322,N_21339,N_22377);
nor U23323 (N_23323,N_21809,N_21603);
nor U23324 (N_23324,N_21752,N_21834);
nand U23325 (N_23325,N_22330,N_21647);
nand U23326 (N_23326,N_21098,N_22048);
xnor U23327 (N_23327,N_22471,N_21371);
nand U23328 (N_23328,N_21529,N_21539);
or U23329 (N_23329,N_21285,N_21471);
xor U23330 (N_23330,N_21690,N_21780);
or U23331 (N_23331,N_21777,N_21085);
or U23332 (N_23332,N_22496,N_22378);
nand U23333 (N_23333,N_22146,N_22057);
nor U23334 (N_23334,N_21413,N_22295);
or U23335 (N_23335,N_21575,N_22155);
nor U23336 (N_23336,N_21137,N_21402);
and U23337 (N_23337,N_22158,N_22304);
or U23338 (N_23338,N_21835,N_21349);
or U23339 (N_23339,N_21218,N_22364);
and U23340 (N_23340,N_21632,N_21627);
and U23341 (N_23341,N_21951,N_21139);
nor U23342 (N_23342,N_21375,N_21985);
nor U23343 (N_23343,N_21402,N_21327);
or U23344 (N_23344,N_21930,N_21465);
nor U23345 (N_23345,N_22040,N_21746);
and U23346 (N_23346,N_22324,N_21754);
xnor U23347 (N_23347,N_21811,N_22161);
or U23348 (N_23348,N_21434,N_22316);
nand U23349 (N_23349,N_21751,N_21961);
nand U23350 (N_23350,N_22186,N_21410);
xor U23351 (N_23351,N_22104,N_21453);
xnor U23352 (N_23352,N_21565,N_21081);
xor U23353 (N_23353,N_21883,N_21366);
xnor U23354 (N_23354,N_22067,N_21259);
or U23355 (N_23355,N_21987,N_21001);
xnor U23356 (N_23356,N_22150,N_21513);
nand U23357 (N_23357,N_21029,N_22249);
nor U23358 (N_23358,N_21566,N_21931);
or U23359 (N_23359,N_21597,N_21279);
nor U23360 (N_23360,N_21860,N_21906);
nor U23361 (N_23361,N_22395,N_22211);
and U23362 (N_23362,N_21850,N_22113);
xnor U23363 (N_23363,N_21310,N_21177);
nand U23364 (N_23364,N_21165,N_22415);
and U23365 (N_23365,N_21811,N_21911);
or U23366 (N_23366,N_21259,N_21011);
nor U23367 (N_23367,N_22425,N_21594);
and U23368 (N_23368,N_22439,N_22090);
nor U23369 (N_23369,N_21992,N_21291);
or U23370 (N_23370,N_22488,N_21807);
nor U23371 (N_23371,N_21946,N_21727);
nand U23372 (N_23372,N_22325,N_21591);
xnor U23373 (N_23373,N_21618,N_22034);
and U23374 (N_23374,N_22482,N_22057);
xor U23375 (N_23375,N_21298,N_21824);
or U23376 (N_23376,N_21265,N_22296);
and U23377 (N_23377,N_21700,N_21854);
nand U23378 (N_23378,N_21885,N_21749);
nand U23379 (N_23379,N_22354,N_22050);
and U23380 (N_23380,N_21308,N_21918);
or U23381 (N_23381,N_22247,N_22435);
or U23382 (N_23382,N_21099,N_21011);
and U23383 (N_23383,N_21900,N_21070);
xnor U23384 (N_23384,N_22202,N_22286);
or U23385 (N_23385,N_21952,N_21317);
nand U23386 (N_23386,N_22276,N_21632);
or U23387 (N_23387,N_22236,N_21528);
or U23388 (N_23388,N_21740,N_21718);
nand U23389 (N_23389,N_22343,N_22242);
or U23390 (N_23390,N_21323,N_22117);
nand U23391 (N_23391,N_22288,N_21471);
or U23392 (N_23392,N_21299,N_21086);
nor U23393 (N_23393,N_21685,N_21802);
xnor U23394 (N_23394,N_22210,N_21904);
xor U23395 (N_23395,N_21988,N_21303);
nand U23396 (N_23396,N_21470,N_21457);
and U23397 (N_23397,N_21521,N_22377);
or U23398 (N_23398,N_22365,N_21048);
or U23399 (N_23399,N_22400,N_21756);
nor U23400 (N_23400,N_22096,N_21255);
xnor U23401 (N_23401,N_22065,N_22075);
and U23402 (N_23402,N_22455,N_22218);
nand U23403 (N_23403,N_22122,N_21708);
xor U23404 (N_23404,N_22296,N_21031);
nor U23405 (N_23405,N_21699,N_21366);
xnor U23406 (N_23406,N_21744,N_21580);
nor U23407 (N_23407,N_21039,N_22168);
and U23408 (N_23408,N_22420,N_21249);
and U23409 (N_23409,N_21477,N_21453);
nand U23410 (N_23410,N_22195,N_21509);
or U23411 (N_23411,N_22477,N_21216);
nor U23412 (N_23412,N_21104,N_22133);
nor U23413 (N_23413,N_21707,N_21763);
nand U23414 (N_23414,N_21965,N_22177);
xor U23415 (N_23415,N_21670,N_21194);
and U23416 (N_23416,N_21888,N_21688);
nor U23417 (N_23417,N_22448,N_21476);
and U23418 (N_23418,N_22196,N_21827);
nor U23419 (N_23419,N_21209,N_21258);
and U23420 (N_23420,N_21336,N_21394);
xnor U23421 (N_23421,N_21574,N_22075);
and U23422 (N_23422,N_21053,N_21956);
and U23423 (N_23423,N_21449,N_22130);
xor U23424 (N_23424,N_21203,N_21126);
or U23425 (N_23425,N_21853,N_21688);
xnor U23426 (N_23426,N_21331,N_21566);
nor U23427 (N_23427,N_21671,N_22406);
xor U23428 (N_23428,N_21204,N_22257);
nor U23429 (N_23429,N_22413,N_21794);
and U23430 (N_23430,N_21949,N_21983);
or U23431 (N_23431,N_21486,N_22148);
nor U23432 (N_23432,N_21624,N_22248);
or U23433 (N_23433,N_22234,N_22118);
nand U23434 (N_23434,N_22348,N_22251);
and U23435 (N_23435,N_22299,N_21153);
nand U23436 (N_23436,N_22197,N_22362);
or U23437 (N_23437,N_21636,N_21953);
xor U23438 (N_23438,N_21814,N_22477);
or U23439 (N_23439,N_21237,N_21463);
nand U23440 (N_23440,N_22211,N_21595);
nor U23441 (N_23441,N_21182,N_22188);
xnor U23442 (N_23442,N_21404,N_21672);
xor U23443 (N_23443,N_22139,N_21588);
nor U23444 (N_23444,N_22480,N_21276);
nor U23445 (N_23445,N_22087,N_21795);
or U23446 (N_23446,N_22029,N_22290);
or U23447 (N_23447,N_21001,N_22059);
nand U23448 (N_23448,N_21503,N_21590);
nor U23449 (N_23449,N_22332,N_22006);
xnor U23450 (N_23450,N_21454,N_22397);
or U23451 (N_23451,N_22055,N_22382);
nor U23452 (N_23452,N_21525,N_22142);
xor U23453 (N_23453,N_21808,N_21519);
nand U23454 (N_23454,N_21893,N_21942);
or U23455 (N_23455,N_22190,N_21673);
nand U23456 (N_23456,N_22399,N_21473);
xnor U23457 (N_23457,N_21285,N_21899);
or U23458 (N_23458,N_21793,N_21630);
nand U23459 (N_23459,N_21286,N_21188);
xor U23460 (N_23460,N_22223,N_21939);
or U23461 (N_23461,N_22194,N_21101);
and U23462 (N_23462,N_21348,N_21740);
xor U23463 (N_23463,N_21918,N_21516);
or U23464 (N_23464,N_21732,N_22396);
or U23465 (N_23465,N_21269,N_22071);
nand U23466 (N_23466,N_21511,N_21160);
nand U23467 (N_23467,N_21934,N_21054);
nand U23468 (N_23468,N_21585,N_21827);
xor U23469 (N_23469,N_21674,N_21785);
or U23470 (N_23470,N_21934,N_21046);
nor U23471 (N_23471,N_21320,N_21790);
nand U23472 (N_23472,N_21455,N_21286);
nor U23473 (N_23473,N_21243,N_21056);
and U23474 (N_23474,N_22415,N_21999);
or U23475 (N_23475,N_21652,N_22178);
nor U23476 (N_23476,N_21757,N_22003);
nand U23477 (N_23477,N_21772,N_21639);
xnor U23478 (N_23478,N_21238,N_21599);
xor U23479 (N_23479,N_22398,N_21424);
xor U23480 (N_23480,N_21495,N_21903);
and U23481 (N_23481,N_21222,N_22372);
xor U23482 (N_23482,N_21515,N_21992);
nor U23483 (N_23483,N_21189,N_21482);
nor U23484 (N_23484,N_21038,N_21627);
nand U23485 (N_23485,N_21338,N_21031);
nor U23486 (N_23486,N_21591,N_21608);
nand U23487 (N_23487,N_21490,N_22271);
nand U23488 (N_23488,N_22330,N_22403);
xnor U23489 (N_23489,N_21050,N_22114);
xnor U23490 (N_23490,N_22362,N_21926);
and U23491 (N_23491,N_21032,N_21309);
and U23492 (N_23492,N_22120,N_21737);
xor U23493 (N_23493,N_21276,N_22095);
xor U23494 (N_23494,N_21602,N_21513);
nor U23495 (N_23495,N_21196,N_22095);
xor U23496 (N_23496,N_21420,N_21584);
or U23497 (N_23497,N_21203,N_22055);
or U23498 (N_23498,N_21220,N_21661);
nand U23499 (N_23499,N_21677,N_21982);
and U23500 (N_23500,N_21257,N_21346);
or U23501 (N_23501,N_22318,N_22402);
xnor U23502 (N_23502,N_21831,N_21648);
nand U23503 (N_23503,N_21164,N_22085);
and U23504 (N_23504,N_21852,N_21810);
and U23505 (N_23505,N_21119,N_21394);
and U23506 (N_23506,N_21105,N_21393);
and U23507 (N_23507,N_22159,N_21428);
and U23508 (N_23508,N_21886,N_21454);
nand U23509 (N_23509,N_21143,N_21085);
nor U23510 (N_23510,N_21211,N_21872);
nor U23511 (N_23511,N_22071,N_21794);
and U23512 (N_23512,N_21431,N_21044);
nor U23513 (N_23513,N_22391,N_21042);
xor U23514 (N_23514,N_21852,N_21088);
and U23515 (N_23515,N_21544,N_21310);
and U23516 (N_23516,N_21761,N_21489);
nand U23517 (N_23517,N_21643,N_21232);
nand U23518 (N_23518,N_21628,N_21356);
xnor U23519 (N_23519,N_21095,N_21361);
nor U23520 (N_23520,N_21307,N_21385);
or U23521 (N_23521,N_21015,N_21145);
and U23522 (N_23522,N_22015,N_21701);
nand U23523 (N_23523,N_22009,N_21470);
and U23524 (N_23524,N_22312,N_22215);
nor U23525 (N_23525,N_21797,N_21387);
or U23526 (N_23526,N_21443,N_22285);
nand U23527 (N_23527,N_22207,N_21424);
or U23528 (N_23528,N_21602,N_21642);
or U23529 (N_23529,N_21699,N_22073);
or U23530 (N_23530,N_21835,N_21770);
and U23531 (N_23531,N_21914,N_21923);
and U23532 (N_23532,N_21989,N_22165);
and U23533 (N_23533,N_22378,N_21267);
xor U23534 (N_23534,N_21759,N_21773);
or U23535 (N_23535,N_22137,N_22210);
nor U23536 (N_23536,N_21408,N_22393);
nor U23537 (N_23537,N_21986,N_21330);
and U23538 (N_23538,N_21679,N_22373);
nor U23539 (N_23539,N_21548,N_21504);
xnor U23540 (N_23540,N_21870,N_21214);
xor U23541 (N_23541,N_22240,N_22272);
nand U23542 (N_23542,N_22415,N_21798);
nor U23543 (N_23543,N_22292,N_21352);
nor U23544 (N_23544,N_21790,N_21328);
nor U23545 (N_23545,N_21528,N_22138);
nor U23546 (N_23546,N_21822,N_22434);
or U23547 (N_23547,N_22259,N_21710);
nand U23548 (N_23548,N_21436,N_21308);
or U23549 (N_23549,N_21804,N_21294);
nand U23550 (N_23550,N_21500,N_22244);
and U23551 (N_23551,N_22184,N_21523);
and U23552 (N_23552,N_22089,N_21743);
or U23553 (N_23553,N_21121,N_21319);
and U23554 (N_23554,N_21692,N_22406);
nor U23555 (N_23555,N_21609,N_22132);
xnor U23556 (N_23556,N_22241,N_21923);
and U23557 (N_23557,N_21087,N_21666);
and U23558 (N_23558,N_21252,N_21210);
or U23559 (N_23559,N_22104,N_21582);
and U23560 (N_23560,N_22433,N_22205);
or U23561 (N_23561,N_21291,N_22349);
or U23562 (N_23562,N_21104,N_21195);
nor U23563 (N_23563,N_21775,N_21831);
nor U23564 (N_23564,N_21336,N_21332);
xnor U23565 (N_23565,N_22200,N_21520);
xor U23566 (N_23566,N_22083,N_22213);
xnor U23567 (N_23567,N_21762,N_21991);
nor U23568 (N_23568,N_22267,N_21295);
nand U23569 (N_23569,N_21077,N_22172);
xor U23570 (N_23570,N_21508,N_22378);
nor U23571 (N_23571,N_22180,N_21893);
nor U23572 (N_23572,N_21968,N_21446);
xnor U23573 (N_23573,N_21450,N_21947);
nand U23574 (N_23574,N_21012,N_21817);
nand U23575 (N_23575,N_22327,N_21427);
nor U23576 (N_23576,N_21039,N_21903);
nor U23577 (N_23577,N_22292,N_22286);
xor U23578 (N_23578,N_21202,N_21742);
nor U23579 (N_23579,N_21585,N_21941);
nor U23580 (N_23580,N_22270,N_22404);
or U23581 (N_23581,N_22244,N_22257);
nor U23582 (N_23582,N_22380,N_21409);
xnor U23583 (N_23583,N_21164,N_21330);
xnor U23584 (N_23584,N_21600,N_21460);
nor U23585 (N_23585,N_21518,N_21130);
or U23586 (N_23586,N_21613,N_21402);
nor U23587 (N_23587,N_22274,N_22070);
nor U23588 (N_23588,N_21154,N_22038);
nor U23589 (N_23589,N_22167,N_21946);
nand U23590 (N_23590,N_22383,N_22433);
xor U23591 (N_23591,N_21309,N_21137);
and U23592 (N_23592,N_21285,N_21159);
nor U23593 (N_23593,N_21320,N_22313);
and U23594 (N_23594,N_22436,N_21911);
nand U23595 (N_23595,N_21530,N_21268);
nand U23596 (N_23596,N_22499,N_21573);
or U23597 (N_23597,N_22014,N_22418);
nand U23598 (N_23598,N_21480,N_21611);
xnor U23599 (N_23599,N_21591,N_22198);
or U23600 (N_23600,N_21794,N_21546);
or U23601 (N_23601,N_21322,N_21566);
or U23602 (N_23602,N_21733,N_22478);
nor U23603 (N_23603,N_22089,N_21464);
and U23604 (N_23604,N_22301,N_21185);
nor U23605 (N_23605,N_21501,N_21642);
or U23606 (N_23606,N_22156,N_22257);
xor U23607 (N_23607,N_21882,N_22367);
xor U23608 (N_23608,N_22166,N_21551);
nand U23609 (N_23609,N_22047,N_21706);
and U23610 (N_23610,N_21687,N_21748);
xnor U23611 (N_23611,N_21042,N_21673);
or U23612 (N_23612,N_22074,N_21316);
and U23613 (N_23613,N_22325,N_21607);
nand U23614 (N_23614,N_22297,N_21839);
nor U23615 (N_23615,N_21880,N_21663);
or U23616 (N_23616,N_22046,N_21679);
nand U23617 (N_23617,N_21956,N_22296);
or U23618 (N_23618,N_21306,N_21835);
and U23619 (N_23619,N_21432,N_21666);
or U23620 (N_23620,N_21860,N_21507);
nand U23621 (N_23621,N_21751,N_22473);
and U23622 (N_23622,N_21202,N_22068);
and U23623 (N_23623,N_21867,N_22470);
xor U23624 (N_23624,N_21355,N_22067);
and U23625 (N_23625,N_21681,N_21355);
nor U23626 (N_23626,N_22140,N_21987);
nor U23627 (N_23627,N_22255,N_22049);
nand U23628 (N_23628,N_21540,N_21228);
nor U23629 (N_23629,N_21513,N_21993);
nand U23630 (N_23630,N_21352,N_22140);
or U23631 (N_23631,N_22267,N_22201);
or U23632 (N_23632,N_22071,N_22405);
or U23633 (N_23633,N_22338,N_21869);
or U23634 (N_23634,N_21222,N_22293);
or U23635 (N_23635,N_22458,N_21826);
or U23636 (N_23636,N_21806,N_21062);
nand U23637 (N_23637,N_21520,N_21484);
or U23638 (N_23638,N_22144,N_22205);
xnor U23639 (N_23639,N_21816,N_21947);
nand U23640 (N_23640,N_22433,N_21551);
and U23641 (N_23641,N_21417,N_21335);
nand U23642 (N_23642,N_22270,N_21495);
nand U23643 (N_23643,N_21983,N_21652);
nor U23644 (N_23644,N_22329,N_22181);
xnor U23645 (N_23645,N_21456,N_22050);
nand U23646 (N_23646,N_21438,N_21528);
or U23647 (N_23647,N_22497,N_22188);
xnor U23648 (N_23648,N_21643,N_21033);
xor U23649 (N_23649,N_21571,N_21060);
or U23650 (N_23650,N_21440,N_21487);
and U23651 (N_23651,N_21274,N_21255);
and U23652 (N_23652,N_21561,N_21668);
and U23653 (N_23653,N_21095,N_21346);
xor U23654 (N_23654,N_21916,N_21814);
xor U23655 (N_23655,N_21068,N_21205);
nor U23656 (N_23656,N_21796,N_22260);
or U23657 (N_23657,N_21708,N_21249);
xor U23658 (N_23658,N_21339,N_22015);
nor U23659 (N_23659,N_22250,N_21625);
nand U23660 (N_23660,N_21034,N_22199);
nor U23661 (N_23661,N_21337,N_21041);
xor U23662 (N_23662,N_21216,N_22026);
xnor U23663 (N_23663,N_21569,N_21514);
and U23664 (N_23664,N_21106,N_21081);
nand U23665 (N_23665,N_21821,N_21997);
and U23666 (N_23666,N_21547,N_22268);
xnor U23667 (N_23667,N_21801,N_22023);
or U23668 (N_23668,N_21689,N_22398);
xor U23669 (N_23669,N_21581,N_21448);
nand U23670 (N_23670,N_21284,N_22239);
xor U23671 (N_23671,N_22195,N_21231);
xor U23672 (N_23672,N_21388,N_21179);
nor U23673 (N_23673,N_22134,N_21830);
xnor U23674 (N_23674,N_22039,N_21914);
or U23675 (N_23675,N_21984,N_22228);
xnor U23676 (N_23676,N_21033,N_21885);
nor U23677 (N_23677,N_21752,N_21395);
xor U23678 (N_23678,N_22469,N_21874);
nand U23679 (N_23679,N_21963,N_21855);
nand U23680 (N_23680,N_21212,N_22465);
nand U23681 (N_23681,N_21084,N_22190);
nand U23682 (N_23682,N_22050,N_22226);
or U23683 (N_23683,N_22047,N_21503);
nand U23684 (N_23684,N_21076,N_22136);
or U23685 (N_23685,N_22087,N_22271);
nor U23686 (N_23686,N_21043,N_22424);
and U23687 (N_23687,N_22333,N_21882);
and U23688 (N_23688,N_22044,N_21991);
or U23689 (N_23689,N_21269,N_21972);
xor U23690 (N_23690,N_21467,N_21415);
nor U23691 (N_23691,N_21418,N_21160);
nand U23692 (N_23692,N_21482,N_21008);
or U23693 (N_23693,N_21714,N_21813);
or U23694 (N_23694,N_21737,N_22275);
and U23695 (N_23695,N_21771,N_21266);
nand U23696 (N_23696,N_21239,N_21385);
xnor U23697 (N_23697,N_21818,N_21542);
nand U23698 (N_23698,N_21249,N_21589);
or U23699 (N_23699,N_22298,N_21967);
nor U23700 (N_23700,N_22308,N_21415);
nand U23701 (N_23701,N_21819,N_21612);
or U23702 (N_23702,N_21591,N_21895);
and U23703 (N_23703,N_21245,N_21153);
or U23704 (N_23704,N_21822,N_21632);
nor U23705 (N_23705,N_21184,N_21347);
nand U23706 (N_23706,N_21189,N_21876);
or U23707 (N_23707,N_21086,N_22148);
or U23708 (N_23708,N_21345,N_21557);
xor U23709 (N_23709,N_21055,N_21428);
xor U23710 (N_23710,N_22251,N_21302);
or U23711 (N_23711,N_22052,N_22447);
nand U23712 (N_23712,N_21948,N_21045);
or U23713 (N_23713,N_21062,N_21431);
nand U23714 (N_23714,N_21515,N_21780);
xnor U23715 (N_23715,N_21010,N_22022);
xor U23716 (N_23716,N_21600,N_22025);
nand U23717 (N_23717,N_22394,N_21119);
nand U23718 (N_23718,N_21992,N_21817);
nand U23719 (N_23719,N_22231,N_22171);
and U23720 (N_23720,N_22067,N_22035);
nand U23721 (N_23721,N_21810,N_21178);
xor U23722 (N_23722,N_21947,N_21959);
and U23723 (N_23723,N_21819,N_21698);
nand U23724 (N_23724,N_21902,N_21290);
nor U23725 (N_23725,N_21429,N_21271);
xnor U23726 (N_23726,N_22316,N_21645);
and U23727 (N_23727,N_21602,N_21941);
or U23728 (N_23728,N_21168,N_21131);
and U23729 (N_23729,N_21633,N_22379);
nand U23730 (N_23730,N_21087,N_22434);
or U23731 (N_23731,N_21218,N_22444);
and U23732 (N_23732,N_21491,N_21948);
xnor U23733 (N_23733,N_21433,N_22188);
or U23734 (N_23734,N_21642,N_22108);
and U23735 (N_23735,N_21839,N_21885);
xor U23736 (N_23736,N_21241,N_21686);
nand U23737 (N_23737,N_22102,N_22476);
nand U23738 (N_23738,N_21633,N_21241);
or U23739 (N_23739,N_21336,N_21821);
and U23740 (N_23740,N_22313,N_21896);
or U23741 (N_23741,N_21531,N_21577);
nor U23742 (N_23742,N_21472,N_21733);
nor U23743 (N_23743,N_21166,N_22112);
or U23744 (N_23744,N_21719,N_22404);
nor U23745 (N_23745,N_22061,N_21268);
and U23746 (N_23746,N_21528,N_21494);
nor U23747 (N_23747,N_21875,N_22064);
or U23748 (N_23748,N_21935,N_21275);
nand U23749 (N_23749,N_21033,N_21284);
nand U23750 (N_23750,N_21853,N_22137);
nor U23751 (N_23751,N_21558,N_22207);
nand U23752 (N_23752,N_21173,N_21127);
xor U23753 (N_23753,N_21967,N_22070);
and U23754 (N_23754,N_21654,N_22487);
and U23755 (N_23755,N_21803,N_21924);
or U23756 (N_23756,N_22347,N_21937);
and U23757 (N_23757,N_21196,N_22051);
nand U23758 (N_23758,N_21454,N_21511);
nor U23759 (N_23759,N_22454,N_22334);
or U23760 (N_23760,N_21098,N_21791);
xor U23761 (N_23761,N_22408,N_22170);
and U23762 (N_23762,N_21485,N_22094);
nor U23763 (N_23763,N_22312,N_21488);
xor U23764 (N_23764,N_22210,N_21391);
nor U23765 (N_23765,N_22329,N_21479);
nand U23766 (N_23766,N_22293,N_21895);
nand U23767 (N_23767,N_22374,N_22011);
xnor U23768 (N_23768,N_21503,N_21277);
nor U23769 (N_23769,N_22184,N_21248);
xor U23770 (N_23770,N_21662,N_22341);
xor U23771 (N_23771,N_22446,N_22369);
or U23772 (N_23772,N_21085,N_21791);
nand U23773 (N_23773,N_22300,N_21891);
nand U23774 (N_23774,N_21716,N_21511);
or U23775 (N_23775,N_21221,N_22422);
and U23776 (N_23776,N_21776,N_21072);
nand U23777 (N_23777,N_21359,N_22411);
nor U23778 (N_23778,N_21930,N_22122);
nand U23779 (N_23779,N_21798,N_21878);
and U23780 (N_23780,N_21056,N_21832);
or U23781 (N_23781,N_21418,N_21925);
nand U23782 (N_23782,N_22031,N_21369);
xnor U23783 (N_23783,N_22320,N_21625);
nor U23784 (N_23784,N_21427,N_21071);
nand U23785 (N_23785,N_21013,N_22423);
nor U23786 (N_23786,N_21016,N_21987);
or U23787 (N_23787,N_21670,N_22182);
nor U23788 (N_23788,N_21523,N_21640);
and U23789 (N_23789,N_21795,N_22228);
xnor U23790 (N_23790,N_21620,N_22351);
and U23791 (N_23791,N_21726,N_22009);
nor U23792 (N_23792,N_21343,N_22300);
and U23793 (N_23793,N_21054,N_22366);
and U23794 (N_23794,N_22003,N_21296);
or U23795 (N_23795,N_21999,N_22323);
or U23796 (N_23796,N_22153,N_21249);
nor U23797 (N_23797,N_21118,N_21544);
and U23798 (N_23798,N_21015,N_22308);
and U23799 (N_23799,N_22355,N_21458);
and U23800 (N_23800,N_21877,N_21794);
or U23801 (N_23801,N_21113,N_21136);
nor U23802 (N_23802,N_22151,N_21841);
and U23803 (N_23803,N_22377,N_21852);
and U23804 (N_23804,N_21862,N_22311);
and U23805 (N_23805,N_21213,N_21658);
and U23806 (N_23806,N_22491,N_21261);
and U23807 (N_23807,N_21117,N_21854);
nor U23808 (N_23808,N_21755,N_21798);
or U23809 (N_23809,N_22163,N_22256);
nor U23810 (N_23810,N_21317,N_21007);
and U23811 (N_23811,N_21225,N_21648);
nand U23812 (N_23812,N_22208,N_21496);
nor U23813 (N_23813,N_22042,N_21953);
nor U23814 (N_23814,N_22028,N_21550);
nand U23815 (N_23815,N_22010,N_21039);
and U23816 (N_23816,N_21698,N_21712);
or U23817 (N_23817,N_21167,N_22219);
nand U23818 (N_23818,N_22226,N_21308);
xnor U23819 (N_23819,N_21480,N_21614);
nor U23820 (N_23820,N_21381,N_21170);
nor U23821 (N_23821,N_22276,N_21805);
or U23822 (N_23822,N_22490,N_22299);
nor U23823 (N_23823,N_21424,N_22118);
and U23824 (N_23824,N_22329,N_22305);
and U23825 (N_23825,N_21960,N_21399);
nor U23826 (N_23826,N_21676,N_21182);
and U23827 (N_23827,N_21021,N_21909);
nor U23828 (N_23828,N_21541,N_22351);
and U23829 (N_23829,N_21990,N_22296);
nand U23830 (N_23830,N_22346,N_21613);
nor U23831 (N_23831,N_21256,N_21517);
xor U23832 (N_23832,N_22005,N_22423);
nand U23833 (N_23833,N_21048,N_22054);
or U23834 (N_23834,N_21678,N_21756);
nor U23835 (N_23835,N_21468,N_21122);
xnor U23836 (N_23836,N_21458,N_22253);
nand U23837 (N_23837,N_22167,N_22025);
or U23838 (N_23838,N_21463,N_22466);
and U23839 (N_23839,N_22147,N_21690);
and U23840 (N_23840,N_21758,N_21796);
nor U23841 (N_23841,N_22266,N_21736);
nor U23842 (N_23842,N_22422,N_21844);
nand U23843 (N_23843,N_22333,N_21255);
nor U23844 (N_23844,N_21419,N_21981);
or U23845 (N_23845,N_21616,N_22234);
and U23846 (N_23846,N_21703,N_22268);
nor U23847 (N_23847,N_22066,N_21853);
nor U23848 (N_23848,N_21241,N_21283);
and U23849 (N_23849,N_21959,N_21795);
xnor U23850 (N_23850,N_21046,N_21727);
nor U23851 (N_23851,N_21576,N_21206);
or U23852 (N_23852,N_21385,N_22395);
nor U23853 (N_23853,N_22248,N_21965);
nand U23854 (N_23854,N_21454,N_22414);
and U23855 (N_23855,N_21690,N_22318);
xnor U23856 (N_23856,N_21214,N_22058);
nand U23857 (N_23857,N_21447,N_22156);
nor U23858 (N_23858,N_21078,N_21978);
and U23859 (N_23859,N_21717,N_22103);
xnor U23860 (N_23860,N_21170,N_21438);
and U23861 (N_23861,N_21215,N_22477);
or U23862 (N_23862,N_21872,N_21885);
or U23863 (N_23863,N_22393,N_21523);
nand U23864 (N_23864,N_21876,N_21500);
and U23865 (N_23865,N_21810,N_22108);
nand U23866 (N_23866,N_22223,N_21306);
or U23867 (N_23867,N_21397,N_22120);
or U23868 (N_23868,N_21041,N_22154);
nor U23869 (N_23869,N_22368,N_22288);
xnor U23870 (N_23870,N_22024,N_21381);
nor U23871 (N_23871,N_22398,N_22258);
nor U23872 (N_23872,N_21816,N_21010);
nand U23873 (N_23873,N_21994,N_21730);
or U23874 (N_23874,N_22366,N_21733);
and U23875 (N_23875,N_21920,N_22364);
and U23876 (N_23876,N_21516,N_21569);
nand U23877 (N_23877,N_21019,N_21972);
nand U23878 (N_23878,N_21515,N_21673);
nand U23879 (N_23879,N_22101,N_22437);
or U23880 (N_23880,N_22134,N_22135);
xor U23881 (N_23881,N_21585,N_21917);
and U23882 (N_23882,N_21615,N_21983);
xor U23883 (N_23883,N_21961,N_21046);
nor U23884 (N_23884,N_21404,N_21893);
nand U23885 (N_23885,N_21685,N_21214);
nor U23886 (N_23886,N_21124,N_21686);
nand U23887 (N_23887,N_21048,N_21337);
xnor U23888 (N_23888,N_21562,N_21503);
nand U23889 (N_23889,N_22357,N_21362);
nor U23890 (N_23890,N_21666,N_21491);
nand U23891 (N_23891,N_21084,N_21518);
and U23892 (N_23892,N_22090,N_22288);
and U23893 (N_23893,N_21111,N_21888);
nor U23894 (N_23894,N_22431,N_21671);
and U23895 (N_23895,N_22349,N_21121);
and U23896 (N_23896,N_21369,N_21709);
or U23897 (N_23897,N_22126,N_22008);
and U23898 (N_23898,N_22263,N_22126);
nand U23899 (N_23899,N_22369,N_21308);
and U23900 (N_23900,N_21206,N_21542);
nor U23901 (N_23901,N_21085,N_21860);
nand U23902 (N_23902,N_22419,N_21573);
or U23903 (N_23903,N_22024,N_21403);
nor U23904 (N_23904,N_21782,N_21020);
nand U23905 (N_23905,N_22105,N_21984);
or U23906 (N_23906,N_22061,N_22047);
or U23907 (N_23907,N_22410,N_21636);
xor U23908 (N_23908,N_21591,N_21531);
or U23909 (N_23909,N_21951,N_21568);
nand U23910 (N_23910,N_21199,N_21702);
nor U23911 (N_23911,N_21008,N_21231);
or U23912 (N_23912,N_21556,N_21963);
and U23913 (N_23913,N_22050,N_22314);
or U23914 (N_23914,N_21192,N_21231);
and U23915 (N_23915,N_21602,N_21923);
or U23916 (N_23916,N_22419,N_21774);
xor U23917 (N_23917,N_21177,N_22391);
nand U23918 (N_23918,N_22037,N_21878);
nand U23919 (N_23919,N_21474,N_21771);
and U23920 (N_23920,N_21678,N_22022);
and U23921 (N_23921,N_21132,N_21240);
nand U23922 (N_23922,N_22289,N_22123);
and U23923 (N_23923,N_21904,N_22236);
or U23924 (N_23924,N_21191,N_21042);
and U23925 (N_23925,N_21624,N_21104);
and U23926 (N_23926,N_21765,N_21984);
xor U23927 (N_23927,N_21985,N_21829);
or U23928 (N_23928,N_21782,N_22363);
or U23929 (N_23929,N_21945,N_21846);
xor U23930 (N_23930,N_21973,N_22376);
xnor U23931 (N_23931,N_21266,N_21519);
or U23932 (N_23932,N_21003,N_21416);
nor U23933 (N_23933,N_22159,N_21552);
nor U23934 (N_23934,N_22481,N_21964);
xnor U23935 (N_23935,N_22251,N_21804);
nand U23936 (N_23936,N_21746,N_21327);
nor U23937 (N_23937,N_21516,N_21128);
and U23938 (N_23938,N_21645,N_21212);
nand U23939 (N_23939,N_21997,N_22054);
xor U23940 (N_23940,N_21270,N_21591);
xor U23941 (N_23941,N_21344,N_21632);
xor U23942 (N_23942,N_21809,N_21111);
xnor U23943 (N_23943,N_21929,N_22456);
xor U23944 (N_23944,N_22041,N_21053);
and U23945 (N_23945,N_21788,N_22064);
xor U23946 (N_23946,N_22168,N_22145);
xnor U23947 (N_23947,N_21272,N_21087);
and U23948 (N_23948,N_21511,N_21721);
xor U23949 (N_23949,N_21997,N_21382);
and U23950 (N_23950,N_21617,N_22384);
or U23951 (N_23951,N_21195,N_21987);
nor U23952 (N_23952,N_22014,N_21404);
nand U23953 (N_23953,N_21834,N_22024);
and U23954 (N_23954,N_22356,N_22159);
nor U23955 (N_23955,N_21250,N_21266);
nand U23956 (N_23956,N_21673,N_21221);
xor U23957 (N_23957,N_21090,N_21785);
nand U23958 (N_23958,N_22360,N_21360);
nor U23959 (N_23959,N_21163,N_22299);
xnor U23960 (N_23960,N_21777,N_21614);
and U23961 (N_23961,N_21532,N_21502);
and U23962 (N_23962,N_21297,N_21819);
and U23963 (N_23963,N_21418,N_22162);
nor U23964 (N_23964,N_21401,N_22006);
and U23965 (N_23965,N_21615,N_22047);
and U23966 (N_23966,N_22180,N_22228);
or U23967 (N_23967,N_21906,N_21076);
nor U23968 (N_23968,N_22146,N_21729);
or U23969 (N_23969,N_21001,N_21614);
nand U23970 (N_23970,N_21730,N_22164);
nand U23971 (N_23971,N_21307,N_21338);
xor U23972 (N_23972,N_21422,N_21477);
or U23973 (N_23973,N_21346,N_21222);
nor U23974 (N_23974,N_21902,N_22401);
and U23975 (N_23975,N_21993,N_21421);
nand U23976 (N_23976,N_22469,N_21906);
nor U23977 (N_23977,N_21171,N_22398);
or U23978 (N_23978,N_21578,N_21078);
or U23979 (N_23979,N_21935,N_22474);
nor U23980 (N_23980,N_22034,N_22489);
nand U23981 (N_23981,N_21591,N_21197);
xor U23982 (N_23982,N_22035,N_22413);
nand U23983 (N_23983,N_22139,N_21977);
xor U23984 (N_23984,N_21749,N_22079);
xnor U23985 (N_23985,N_21529,N_21582);
xnor U23986 (N_23986,N_21024,N_21415);
or U23987 (N_23987,N_21859,N_21209);
nor U23988 (N_23988,N_21091,N_21406);
and U23989 (N_23989,N_22008,N_21660);
or U23990 (N_23990,N_21600,N_22378);
or U23991 (N_23991,N_22084,N_22366);
xnor U23992 (N_23992,N_21339,N_21905);
xor U23993 (N_23993,N_22272,N_21709);
nor U23994 (N_23994,N_21448,N_22463);
xor U23995 (N_23995,N_22289,N_21905);
nand U23996 (N_23996,N_22248,N_22400);
xnor U23997 (N_23997,N_21862,N_21367);
and U23998 (N_23998,N_21404,N_21663);
or U23999 (N_23999,N_22191,N_21247);
nor U24000 (N_24000,N_23657,N_23432);
xnor U24001 (N_24001,N_23313,N_23211);
nor U24002 (N_24002,N_23884,N_23570);
nor U24003 (N_24003,N_23149,N_23721);
and U24004 (N_24004,N_23790,N_22720);
xor U24005 (N_24005,N_23034,N_23320);
nor U24006 (N_24006,N_23378,N_22662);
and U24007 (N_24007,N_22975,N_23163);
and U24008 (N_24008,N_23779,N_23515);
nor U24009 (N_24009,N_23248,N_23835);
or U24010 (N_24010,N_23323,N_22624);
xnor U24011 (N_24011,N_22997,N_23176);
and U24012 (N_24012,N_22703,N_23469);
and U24013 (N_24013,N_22695,N_22635);
xnor U24014 (N_24014,N_22972,N_23221);
or U24015 (N_24015,N_22774,N_23353);
or U24016 (N_24016,N_23670,N_22536);
xnor U24017 (N_24017,N_23077,N_23026);
xor U24018 (N_24018,N_23047,N_23068);
and U24019 (N_24019,N_23289,N_23634);
nor U24020 (N_24020,N_22967,N_22863);
xnor U24021 (N_24021,N_22823,N_22765);
xor U24022 (N_24022,N_22963,N_22831);
or U24023 (N_24023,N_23763,N_23167);
xor U24024 (N_24024,N_23510,N_23295);
xor U24025 (N_24025,N_22830,N_23494);
and U24026 (N_24026,N_23290,N_22818);
and U24027 (N_24027,N_23303,N_23562);
xor U24028 (N_24028,N_23777,N_22752);
or U24029 (N_24029,N_22746,N_22600);
or U24030 (N_24030,N_22648,N_23481);
or U24031 (N_24031,N_22591,N_23645);
nor U24032 (N_24032,N_22582,N_23193);
nor U24033 (N_24033,N_22702,N_23737);
nand U24034 (N_24034,N_23472,N_23132);
or U24035 (N_24035,N_23638,N_23943);
and U24036 (N_24036,N_23128,N_23946);
nand U24037 (N_24037,N_23924,N_23498);
or U24038 (N_24038,N_22503,N_23143);
or U24039 (N_24039,N_23403,N_23129);
nand U24040 (N_24040,N_23658,N_23892);
and U24041 (N_24041,N_22512,N_23118);
nand U24042 (N_24042,N_22849,N_23565);
xor U24043 (N_24043,N_23327,N_22511);
or U24044 (N_24044,N_22885,N_23233);
nor U24045 (N_24045,N_23591,N_23385);
nor U24046 (N_24046,N_23567,N_22527);
nor U24047 (N_24047,N_23896,N_23619);
nand U24048 (N_24048,N_23782,N_22881);
and U24049 (N_24049,N_23170,N_22783);
and U24050 (N_24050,N_23073,N_23535);
and U24051 (N_24051,N_23541,N_23746);
or U24052 (N_24052,N_23608,N_23144);
xor U24053 (N_24053,N_22739,N_23738);
nor U24054 (N_24054,N_23430,N_23933);
nor U24055 (N_24055,N_23484,N_22639);
xor U24056 (N_24056,N_23421,N_23610);
or U24057 (N_24057,N_23398,N_22510);
and U24058 (N_24058,N_22785,N_22854);
nand U24059 (N_24059,N_23775,N_23940);
or U24060 (N_24060,N_22688,N_22870);
xnor U24061 (N_24061,N_22607,N_22569);
xor U24062 (N_24062,N_23092,N_23527);
nand U24063 (N_24063,N_23112,N_23093);
nor U24064 (N_24064,N_23982,N_23711);
xnor U24065 (N_24065,N_22542,N_23257);
xor U24066 (N_24066,N_23100,N_23194);
and U24067 (N_24067,N_22508,N_23984);
and U24068 (N_24068,N_23250,N_23795);
xnor U24069 (N_24069,N_22796,N_23676);
xnor U24070 (N_24070,N_23949,N_23703);
or U24071 (N_24071,N_23369,N_22608);
and U24072 (N_24072,N_23329,N_23741);
or U24073 (N_24073,N_22782,N_23604);
nand U24074 (N_24074,N_23027,N_22916);
and U24075 (N_24075,N_23435,N_22737);
nor U24076 (N_24076,N_23715,N_23519);
and U24077 (N_24077,N_23865,N_23449);
nand U24078 (N_24078,N_22586,N_23319);
xor U24079 (N_24079,N_23989,N_23287);
and U24080 (N_24080,N_23564,N_23603);
nor U24081 (N_24081,N_23551,N_23104);
nand U24082 (N_24082,N_23954,N_23908);
xnor U24083 (N_24083,N_23044,N_23222);
or U24084 (N_24084,N_22731,N_22622);
nor U24085 (N_24085,N_23674,N_23810);
and U24086 (N_24086,N_23917,N_23899);
and U24087 (N_24087,N_23702,N_22883);
or U24088 (N_24088,N_23939,N_23124);
or U24089 (N_24089,N_23051,N_23596);
nor U24090 (N_24090,N_23103,N_22806);
nand U24091 (N_24091,N_22515,N_23723);
and U24092 (N_24092,N_23354,N_23069);
nor U24093 (N_24093,N_23190,N_23478);
xor U24094 (N_24094,N_22686,N_23483);
xnor U24095 (N_24095,N_23972,N_23107);
and U24096 (N_24096,N_23158,N_23082);
nor U24097 (N_24097,N_22659,N_23505);
and U24098 (N_24098,N_22960,N_22760);
or U24099 (N_24099,N_22875,N_23063);
nor U24100 (N_24100,N_23200,N_23004);
and U24101 (N_24101,N_23114,N_23245);
nand U24102 (N_24102,N_23117,N_22903);
and U24103 (N_24103,N_23827,N_22990);
or U24104 (N_24104,N_22947,N_23819);
xor U24105 (N_24105,N_23745,N_22565);
or U24106 (N_24106,N_22706,N_23601);
or U24107 (N_24107,N_23171,N_23631);
nor U24108 (N_24108,N_23405,N_23576);
or U24109 (N_24109,N_23188,N_23783);
nand U24110 (N_24110,N_23692,N_22729);
nand U24111 (N_24111,N_22541,N_22504);
nor U24112 (N_24112,N_22520,N_22502);
and U24113 (N_24113,N_22554,N_23504);
and U24114 (N_24114,N_22709,N_23440);
xor U24115 (N_24115,N_23719,N_23797);
or U24116 (N_24116,N_23014,N_23647);
or U24117 (N_24117,N_22721,N_23913);
nor U24118 (N_24118,N_22749,N_23849);
or U24119 (N_24119,N_22750,N_23363);
and U24120 (N_24120,N_22613,N_22692);
xor U24121 (N_24121,N_23197,N_23842);
or U24122 (N_24122,N_23108,N_23424);
and U24123 (N_24123,N_22681,N_22590);
nor U24124 (N_24124,N_22704,N_23630);
xnor U24125 (N_24125,N_22987,N_22759);
nand U24126 (N_24126,N_23729,N_22677);
xnor U24127 (N_24127,N_22812,N_23029);
nor U24128 (N_24128,N_22609,N_22905);
nor U24129 (N_24129,N_22955,N_22531);
and U24130 (N_24130,N_23667,N_23115);
nand U24131 (N_24131,N_23434,N_23411);
xor U24132 (N_24132,N_23249,N_23105);
and U24133 (N_24133,N_22580,N_23864);
xor U24134 (N_24134,N_23036,N_22816);
and U24135 (N_24135,N_23649,N_22650);
xnor U24136 (N_24136,N_23895,N_22566);
xor U24137 (N_24137,N_23888,N_23902);
xor U24138 (N_24138,N_22902,N_23276);
or U24139 (N_24139,N_22780,N_22835);
nor U24140 (N_24140,N_23686,N_22884);
or U24141 (N_24141,N_23852,N_23627);
or U24142 (N_24142,N_23488,N_22839);
nor U24143 (N_24143,N_23860,N_23552);
nand U24144 (N_24144,N_23655,N_23695);
nand U24145 (N_24145,N_22654,N_23714);
xnor U24146 (N_24146,N_22999,N_23404);
nand U24147 (N_24147,N_22507,N_23359);
and U24148 (N_24148,N_22973,N_23572);
nor U24149 (N_24149,N_23396,N_22957);
or U24150 (N_24150,N_22921,N_22755);
xor U24151 (N_24151,N_22841,N_23962);
nand U24152 (N_24152,N_23280,N_23212);
and U24153 (N_24153,N_23428,N_23662);
xor U24154 (N_24154,N_23208,N_23254);
xor U24155 (N_24155,N_23656,N_23644);
xor U24156 (N_24156,N_22573,N_22931);
or U24157 (N_24157,N_23735,N_23890);
or U24158 (N_24158,N_23928,N_23760);
nor U24159 (N_24159,N_23815,N_22584);
xnor U24160 (N_24160,N_23184,N_23925);
nand U24161 (N_24161,N_22917,N_23371);
and U24162 (N_24162,N_22705,N_23635);
xor U24163 (N_24163,N_22912,N_23583);
and U24164 (N_24164,N_23533,N_22714);
nor U24165 (N_24165,N_23712,N_22733);
and U24166 (N_24166,N_23102,N_23431);
xnor U24167 (N_24167,N_23322,N_23585);
nor U24168 (N_24168,N_22528,N_23672);
and U24169 (N_24169,N_23346,N_22778);
or U24170 (N_24170,N_23986,N_23773);
nor U24171 (N_24171,N_23389,N_22814);
and U24172 (N_24172,N_22718,N_22930);
nor U24173 (N_24173,N_23417,N_23834);
and U24174 (N_24174,N_23640,N_23531);
or U24175 (N_24175,N_23931,N_23343);
or U24176 (N_24176,N_23620,N_23569);
nor U24177 (N_24177,N_23001,N_23708);
or U24178 (N_24178,N_23750,N_23055);
or U24179 (N_24179,N_23707,N_22556);
xor U24180 (N_24180,N_23592,N_22577);
nor U24181 (N_24181,N_23938,N_22754);
xor U24182 (N_24182,N_22631,N_23406);
xor U24183 (N_24183,N_22652,N_23458);
nand U24184 (N_24184,N_22674,N_23263);
nand U24185 (N_24185,N_23206,N_23970);
nor U24186 (N_24186,N_23789,N_23127);
nand U24187 (N_24187,N_23755,N_22517);
nor U24188 (N_24188,N_22657,N_23305);
nand U24189 (N_24189,N_23247,N_22678);
nand U24190 (N_24190,N_23218,N_22651);
nor U24191 (N_24191,N_23372,N_23087);
or U24192 (N_24192,N_23258,N_22981);
nand U24193 (N_24193,N_22526,N_23936);
and U24194 (N_24194,N_23660,N_23455);
xnor U24195 (N_24195,N_23579,N_22633);
nor U24196 (N_24196,N_22988,N_23800);
and U24197 (N_24197,N_22642,N_23545);
nand U24198 (N_24198,N_22588,N_23781);
nand U24199 (N_24199,N_22529,N_23736);
or U24200 (N_24200,N_23784,N_23438);
and U24201 (N_24201,N_22667,N_23049);
or U24202 (N_24202,N_23877,N_22587);
nand U24203 (N_24203,N_23493,N_23198);
xnor U24204 (N_24204,N_23845,N_22521);
xnor U24205 (N_24205,N_23345,N_22575);
nand U24206 (N_24206,N_23952,N_23140);
nand U24207 (N_24207,N_23985,N_23556);
and U24208 (N_24208,N_22594,N_23587);
nand U24209 (N_24209,N_23005,N_22669);
nor U24210 (N_24210,N_23761,N_23123);
nand U24211 (N_24211,N_23806,N_22908);
and U24212 (N_24212,N_23187,N_23240);
or U24213 (N_24213,N_22799,N_22948);
nor U24214 (N_24214,N_23203,N_23872);
nand U24215 (N_24215,N_23452,N_23475);
nor U24216 (N_24216,N_23157,N_23612);
nand U24217 (N_24217,N_23487,N_23558);
and U24218 (N_24218,N_23397,N_23035);
nor U24219 (N_24219,N_22843,N_22898);
nand U24220 (N_24220,N_23568,N_22953);
nor U24221 (N_24221,N_23307,N_22661);
or U24222 (N_24222,N_23419,N_23024);
nor U24223 (N_24223,N_23727,N_23650);
xor U24224 (N_24224,N_22901,N_23999);
nor U24225 (N_24225,N_23122,N_23690);
and U24226 (N_24226,N_23529,N_23274);
nand U24227 (N_24227,N_23713,N_23709);
and U24228 (N_24228,N_23234,N_23915);
xor U24229 (N_24229,N_22880,N_22630);
and U24230 (N_24230,N_22819,N_23220);
and U24231 (N_24231,N_22810,N_22665);
and U24232 (N_24232,N_22712,N_23480);
or U24233 (N_24233,N_22506,N_23718);
and U24234 (N_24234,N_23532,N_23145);
or U24235 (N_24235,N_22864,N_23161);
or U24236 (N_24236,N_23751,N_22539);
nor U24237 (N_24237,N_22614,N_22919);
nor U24238 (N_24238,N_23930,N_23586);
nor U24239 (N_24239,N_22833,N_23770);
or U24240 (N_24240,N_23664,N_23056);
xnor U24241 (N_24241,N_23778,N_23978);
xnor U24242 (N_24242,N_23390,N_23409);
nor U24243 (N_24243,N_23683,N_23720);
nor U24244 (N_24244,N_23294,N_22699);
or U24245 (N_24245,N_22974,N_22598);
nand U24246 (N_24246,N_23859,N_23651);
nand U24247 (N_24247,N_23229,N_23089);
xor U24248 (N_24248,N_23801,N_23079);
xor U24249 (N_24249,N_23752,N_22548);
nor U24250 (N_24250,N_22562,N_23516);
xor U24251 (N_24251,N_23110,N_22940);
nor U24252 (N_24252,N_22860,N_23880);
or U24253 (N_24253,N_22932,N_23503);
nor U24254 (N_24254,N_23898,N_23698);
and U24255 (N_24255,N_22959,N_22578);
nor U24256 (N_24256,N_23688,N_23597);
xor U24257 (N_24257,N_22787,N_23018);
xnor U24258 (N_24258,N_22552,N_22592);
nor U24259 (N_24259,N_22942,N_23791);
nor U24260 (N_24260,N_22751,N_22876);
or U24261 (N_24261,N_23858,N_23066);
nand U24262 (N_24262,N_23669,N_22889);
nand U24263 (N_24263,N_22525,N_23909);
nand U24264 (N_24264,N_23975,N_22646);
xnor U24265 (N_24265,N_23052,N_23538);
and U24266 (N_24266,N_23547,N_23618);
or U24267 (N_24267,N_23734,N_22576);
nand U24268 (N_24268,N_22951,N_23401);
nor U24269 (N_24269,N_23701,N_23191);
nor U24270 (N_24270,N_22768,N_23410);
nor U24271 (N_24271,N_23617,N_22713);
or U24272 (N_24272,N_23526,N_22853);
xnor U24273 (N_24273,N_22716,N_23964);
and U24274 (N_24274,N_23942,N_22828);
xnor U24275 (N_24275,N_23091,N_23748);
and U24276 (N_24276,N_22732,N_23609);
and U24277 (N_24277,N_23111,N_23973);
or U24278 (N_24278,N_23282,N_23015);
and U24279 (N_24279,N_23341,N_23357);
xor U24280 (N_24280,N_23628,N_23654);
xor U24281 (N_24281,N_23181,N_23887);
xnor U24282 (N_24282,N_22914,N_23951);
nand U24283 (N_24283,N_22730,N_23134);
or U24284 (N_24284,N_22516,N_23333);
nand U24285 (N_24285,N_22952,N_22879);
nand U24286 (N_24286,N_23325,N_22866);
nand U24287 (N_24287,N_23444,N_23792);
and U24288 (N_24288,N_23347,N_23814);
or U24289 (N_24289,N_23956,N_23490);
or U24290 (N_24290,N_23622,N_23874);
nand U24291 (N_24291,N_22845,N_23934);
nor U24292 (N_24292,N_23607,N_23119);
nor U24293 (N_24293,N_23965,N_23577);
or U24294 (N_24294,N_23740,N_22763);
and U24295 (N_24295,N_22821,N_22567);
xor U24296 (N_24296,N_23360,N_22824);
xor U24297 (N_24297,N_22532,N_23159);
nand U24298 (N_24298,N_23809,N_23016);
nor U24299 (N_24299,N_23252,N_22557);
and U24300 (N_24300,N_23811,N_22872);
xnor U24301 (N_24301,N_23121,N_23590);
nand U24302 (N_24302,N_23230,N_23776);
xnor U24303 (N_24303,N_23853,N_23045);
or U24304 (N_24304,N_23967,N_23418);
or U24305 (N_24305,N_23626,N_23725);
and U24306 (N_24306,N_22615,N_22920);
or U24307 (N_24307,N_23213,N_23370);
xor U24308 (N_24308,N_23466,N_23958);
nor U24309 (N_24309,N_22789,N_23981);
nand U24310 (N_24310,N_22840,N_22900);
nand U24311 (N_24311,N_23316,N_23384);
or U24312 (N_24312,N_23020,N_23499);
or U24313 (N_24313,N_23297,N_23451);
xor U24314 (N_24314,N_23427,N_23283);
or U24315 (N_24315,N_22954,N_22777);
nand U24316 (N_24316,N_23846,N_23415);
nand U24317 (N_24317,N_23468,N_23095);
nor U24318 (N_24318,N_22968,N_23733);
nand U24319 (N_24319,N_23772,N_23335);
xnor U24320 (N_24320,N_22553,N_23030);
xnor U24321 (N_24321,N_23201,N_23543);
nand U24322 (N_24322,N_23796,N_22794);
and U24323 (N_24323,N_23994,N_22822);
xor U24324 (N_24324,N_23446,N_23106);
and U24325 (N_24325,N_22533,N_23947);
nand U24326 (N_24326,N_22804,N_22802);
nor U24327 (N_24327,N_23169,N_23367);
and U24328 (N_24328,N_23301,N_23813);
nor U24329 (N_24329,N_23511,N_23138);
xnor U24330 (N_24330,N_23017,N_23302);
or U24331 (N_24331,N_23050,N_23331);
xnor U24332 (N_24332,N_23224,N_22728);
xnor U24333 (N_24333,N_23697,N_22891);
nor U24334 (N_24334,N_23236,N_23793);
nand U24335 (N_24335,N_22998,N_23041);
nand U24336 (N_24336,N_22756,N_22523);
or U24337 (N_24337,N_23977,N_23255);
or U24338 (N_24338,N_23365,N_22513);
xor U24339 (N_24339,N_23416,N_23464);
nor U24340 (N_24340,N_23996,N_23262);
xor U24341 (N_24341,N_23172,N_22772);
nor U24342 (N_24342,N_23706,N_23207);
nor U24343 (N_24343,N_23120,N_23882);
and U24344 (N_24344,N_22623,N_23209);
nor U24345 (N_24345,N_22698,N_22869);
xnor U24346 (N_24346,N_23361,N_22585);
nor U24347 (N_24347,N_23682,N_22962);
nor U24348 (N_24348,N_22892,N_23855);
xor U24349 (N_24349,N_22753,N_23885);
and U24350 (N_24350,N_22805,N_23722);
or U24351 (N_24351,N_22736,N_23039);
nor U24352 (N_24352,N_22910,N_23328);
nand U24353 (N_24353,N_23461,N_23780);
nor U24354 (N_24354,N_22572,N_23728);
nand U24355 (N_24355,N_23086,N_23423);
nor U24356 (N_24356,N_23175,N_23643);
xnor U24357 (N_24357,N_23293,N_23270);
nand U24358 (N_24358,N_23223,N_23136);
nand U24359 (N_24359,N_23765,N_23351);
and U24360 (N_24360,N_22757,N_23724);
or U24361 (N_24361,N_23919,N_23555);
xor U24362 (N_24362,N_23009,N_23277);
nand U24363 (N_24363,N_22836,N_23154);
nand U24364 (N_24364,N_23021,N_22922);
xor U24365 (N_24365,N_22924,N_22538);
xnor U24366 (N_24366,N_22980,N_23495);
nor U24367 (N_24367,N_23311,N_23275);
or U24368 (N_24368,N_23377,N_23685);
and U24369 (N_24369,N_23987,N_23285);
xnor U24370 (N_24370,N_23716,N_23366);
nor U24371 (N_24371,N_23268,N_22882);
nor U24372 (N_24372,N_22738,N_23031);
or U24373 (N_24373,N_23893,N_22771);
xor U24374 (N_24374,N_23355,N_22670);
and U24375 (N_24375,N_23324,N_23309);
nand U24376 (N_24376,N_23349,N_22888);
and U24377 (N_24377,N_23876,N_22874);
and U24378 (N_24378,N_23040,N_22991);
xnor U24379 (N_24379,N_23334,N_22926);
or U24380 (N_24380,N_23704,N_22983);
nor U24381 (N_24381,N_23673,N_23629);
xnor U24382 (N_24382,N_22671,N_23147);
xor U24383 (N_24383,N_23457,N_23786);
nor U24384 (N_24384,N_23976,N_23391);
and U24385 (N_24385,N_23273,N_23929);
nand U24386 (N_24386,N_23336,N_23653);
xor U24387 (N_24387,N_22982,N_22627);
nand U24388 (N_24388,N_22899,N_22559);
and U24389 (N_24389,N_23348,N_23205);
xor U24390 (N_24390,N_23807,N_23957);
or U24391 (N_24391,N_23462,N_23665);
nor U24392 (N_24392,N_22871,N_22803);
or U24393 (N_24393,N_23173,N_22929);
and U24394 (N_24394,N_23575,N_23272);
or U24395 (N_24395,N_23094,N_22989);
or U24396 (N_24396,N_23375,N_23151);
or U24397 (N_24397,N_23439,N_23180);
xor U24398 (N_24398,N_23839,N_23983);
nand U24399 (N_24399,N_23910,N_22767);
and U24400 (N_24400,N_23788,N_23506);
xnor U24401 (N_24401,N_22769,N_23219);
nor U24402 (N_24402,N_23061,N_23589);
or U24403 (N_24403,N_23253,N_23148);
nor U24404 (N_24404,N_22658,N_23502);
or U24405 (N_24405,N_23083,N_22518);
xor U24406 (N_24406,N_23726,N_23314);
and U24407 (N_24407,N_23903,N_22643);
or U24408 (N_24408,N_22664,N_22690);
and U24409 (N_24409,N_22647,N_23216);
nand U24410 (N_24410,N_23474,N_23841);
nor U24411 (N_24411,N_23192,N_23296);
nor U24412 (N_24412,N_22687,N_22795);
nand U24413 (N_24413,N_22894,N_22602);
or U24414 (N_24414,N_23429,N_23991);
and U24415 (N_24415,N_23215,N_23267);
or U24416 (N_24416,N_22761,N_23879);
or U24417 (N_24417,N_23160,N_23559);
and U24418 (N_24418,N_23284,N_22612);
xor U24419 (N_24419,N_23997,N_23337);
xnor U24420 (N_24420,N_22873,N_22711);
nand U24421 (N_24421,N_23142,N_23768);
nor U24422 (N_24422,N_22744,N_22915);
nor U24423 (N_24423,N_22878,N_22640);
or U24424 (N_24424,N_23677,N_23412);
and U24425 (N_24425,N_22722,N_22621);
and U24426 (N_24426,N_22628,N_23130);
xor U24427 (N_24427,N_23269,N_23794);
nand U24428 (N_24428,N_23743,N_22918);
or U24429 (N_24429,N_23584,N_23072);
and U24430 (N_24430,N_23065,N_22969);
nor U24431 (N_24431,N_23243,N_22995);
and U24432 (N_24432,N_22897,N_23445);
nor U24433 (N_24433,N_23204,N_23854);
nor U24434 (N_24434,N_22797,N_23028);
nand U24435 (N_24435,N_23085,N_23742);
and U24436 (N_24436,N_23605,N_23186);
or U24437 (N_24437,N_23453,N_23485);
nand U24438 (N_24438,N_23174,N_22855);
or U24439 (N_24439,N_23561,N_22817);
nand U24440 (N_24440,N_22530,N_23600);
or U24441 (N_24441,N_23537,N_23812);
xnor U24442 (N_24442,N_22813,N_23033);
nor U24443 (N_24443,N_23637,N_23447);
xnor U24444 (N_24444,N_23486,N_23497);
xor U24445 (N_24445,N_23730,N_22636);
or U24446 (N_24446,N_22781,N_23615);
xnor U24447 (N_24447,N_22837,N_22597);
xnor U24448 (N_24448,N_23306,N_22945);
xor U24449 (N_24449,N_22534,N_22984);
or U24450 (N_24450,N_23580,N_22500);
or U24451 (N_24451,N_23832,N_23312);
xnor U24452 (N_24452,N_22555,N_22784);
nand U24453 (N_24453,N_22563,N_23010);
and U24454 (N_24454,N_22815,N_22685);
nor U24455 (N_24455,N_23442,N_23388);
nor U24456 (N_24456,N_23826,N_22847);
nor U24457 (N_24457,N_23407,N_22735);
nor U24458 (N_24458,N_23818,N_22857);
nor U24459 (N_24459,N_23489,N_23386);
or U24460 (N_24460,N_22606,N_23805);
and U24461 (N_24461,N_23179,N_22550);
and U24462 (N_24462,N_23847,N_23426);
or U24463 (N_24463,N_22682,N_23217);
nand U24464 (N_24464,N_22568,N_23006);
nor U24465 (N_24465,N_23993,N_23536);
xnor U24466 (N_24466,N_23582,N_23873);
or U24467 (N_24467,N_22571,N_23990);
or U24468 (N_24468,N_23661,N_22691);
nor U24469 (N_24469,N_23912,N_23566);
and U24470 (N_24470,N_23231,N_23691);
nor U24471 (N_24471,N_22514,N_23182);
xnor U24472 (N_24472,N_23731,N_22599);
or U24473 (N_24473,N_23945,N_23321);
or U24474 (N_24474,N_23666,N_23689);
xnor U24475 (N_24475,N_22747,N_23081);
nor U24476 (N_24476,N_23758,N_22694);
nand U24477 (N_24477,N_23802,N_22641);
or U24478 (N_24478,N_22680,N_22971);
nor U24479 (N_24479,N_22676,N_23808);
nor U24480 (N_24480,N_22776,N_23528);
or U24481 (N_24481,N_22724,N_22928);
nor U24482 (N_24482,N_22734,N_23969);
and U24483 (N_24483,N_23950,N_22977);
xor U24484 (N_24484,N_23995,N_23152);
xor U24485 (N_24485,N_22603,N_23693);
nand U24486 (N_24486,N_22710,N_23639);
nand U24487 (N_24487,N_23992,N_23869);
and U24488 (N_24488,N_22966,N_22993);
and U24489 (N_24489,N_22941,N_23459);
nor U24490 (N_24490,N_22509,N_23623);
xor U24491 (N_24491,N_23477,N_22540);
and U24492 (N_24492,N_23237,N_23739);
xor U24493 (N_24493,N_23828,N_23759);
xor U24494 (N_24494,N_23202,N_23299);
xnor U24495 (N_24495,N_22944,N_23042);
nand U24496 (N_24496,N_22766,N_23922);
and U24497 (N_24497,N_22637,N_22994);
nor U24498 (N_24498,N_22911,N_23680);
nor U24499 (N_24499,N_23684,N_23593);
nand U24500 (N_24500,N_23300,N_22549);
xor U24501 (N_24501,N_23594,N_22547);
and U24502 (N_24502,N_22848,N_23225);
nand U24503 (N_24503,N_23196,N_23141);
or U24504 (N_24504,N_23875,N_23941);
xor U24505 (N_24505,N_23659,N_23058);
xnor U24506 (N_24506,N_23113,N_23214);
nand U24507 (N_24507,N_23038,N_23646);
or U24508 (N_24508,N_22675,N_23133);
or U24509 (N_24509,N_23266,N_23553);
and U24510 (N_24510,N_23054,N_23076);
nor U24511 (N_24511,N_23563,N_22956);
or U24512 (N_24512,N_22865,N_22583);
nor U24513 (N_24513,N_23162,N_23395);
or U24514 (N_24514,N_23340,N_23126);
xor U24515 (N_24515,N_22519,N_23549);
and U24516 (N_24516,N_22727,N_23663);
or U24517 (N_24517,N_22779,N_22790);
nand U24518 (N_24518,N_23008,N_23292);
or U24519 (N_24519,N_22626,N_23901);
or U24520 (N_24520,N_23817,N_23338);
nand U24521 (N_24521,N_23053,N_22844);
and U24522 (N_24522,N_23671,N_22668);
xor U24523 (N_24523,N_23530,N_23747);
and U24524 (N_24524,N_23023,N_22801);
and U24525 (N_24525,N_22909,N_23642);
nor U24526 (N_24526,N_23342,N_23588);
nor U24527 (N_24527,N_23131,N_22505);
and U24528 (N_24528,N_22826,N_23920);
and U24529 (N_24529,N_23837,N_23139);
and U24530 (N_24530,N_22570,N_22773);
and U24531 (N_24531,N_23904,N_23769);
nor U24532 (N_24532,N_22775,N_23304);
or U24533 (N_24533,N_23150,N_22887);
nor U24534 (N_24534,N_23980,N_22545);
nand U24535 (N_24535,N_23916,N_22933);
nor U24536 (N_24536,N_23907,N_23521);
nand U24537 (N_24537,N_23932,N_23291);
nand U24538 (N_24538,N_23011,N_22673);
and U24539 (N_24539,N_22950,N_22632);
or U24540 (N_24540,N_23380,N_23862);
nand U24541 (N_24541,N_23829,N_22904);
and U24542 (N_24542,N_23402,N_22638);
xnor U24543 (N_24543,N_22958,N_23101);
xor U24544 (N_24544,N_23433,N_23096);
xnor U24545 (N_24545,N_23840,N_23279);
and U24546 (N_24546,N_23064,N_22745);
and U24547 (N_24547,N_22701,N_23652);
nand U24548 (N_24548,N_23544,N_22629);
or U24549 (N_24549,N_23060,N_23974);
xor U24550 (N_24550,N_23754,N_22937);
nand U24551 (N_24551,N_23998,N_22938);
nor U24552 (N_24552,N_23675,N_23062);
nor U24553 (N_24553,N_22617,N_23766);
or U24554 (N_24554,N_23878,N_23308);
nor U24555 (N_24555,N_23265,N_23851);
nand U24556 (N_24556,N_23955,N_23833);
nand U24557 (N_24557,N_22683,N_22707);
or U24558 (N_24558,N_23048,N_23641);
and U24559 (N_24559,N_22666,N_22820);
and U24560 (N_24560,N_22992,N_23344);
nor U24561 (N_24561,N_23413,N_22935);
nand U24562 (N_24562,N_22852,N_23534);
and U24563 (N_24563,N_23914,N_23135);
and U24564 (N_24564,N_22978,N_23948);
or U24565 (N_24565,N_22923,N_22717);
or U24566 (N_24566,N_22907,N_23244);
or U24567 (N_24567,N_23578,N_23678);
nor U24568 (N_24568,N_23979,N_23866);
xnor U24569 (N_24569,N_23116,N_22964);
and U24570 (N_24570,N_22850,N_23097);
and U24571 (N_24571,N_23330,N_22719);
or U24572 (N_24572,N_23926,N_23399);
or U24573 (N_24573,N_23025,N_23394);
xnor U24574 (N_24574,N_22579,N_23352);
or U24575 (N_24575,N_23003,N_23700);
nor U24576 (N_24576,N_23441,N_23239);
nor U24577 (N_24577,N_23476,N_23518);
nor U24578 (N_24578,N_22522,N_23844);
xor U24579 (N_24579,N_23821,N_23166);
and U24580 (N_24580,N_23906,N_23288);
xor U24581 (N_24581,N_22697,N_23032);
or U24582 (N_24582,N_22596,N_23961);
nand U24583 (N_24583,N_23492,N_23501);
nand U24584 (N_24584,N_23512,N_22792);
or U24585 (N_24585,N_23621,N_22842);
and U24586 (N_24586,N_23000,N_22660);
nor U24587 (N_24587,N_22961,N_22634);
nand U24588 (N_24588,N_22618,N_23900);
xor U24589 (N_24589,N_22560,N_23463);
or U24590 (N_24590,N_23425,N_22851);
nand U24591 (N_24591,N_23883,N_23816);
nor U24592 (N_24592,N_23271,N_23542);
and U24593 (N_24593,N_23507,N_23850);
nor U24594 (N_24594,N_22740,N_22581);
and U24595 (N_24595,N_23070,N_22610);
and U24596 (N_24596,N_23971,N_23326);
xor U24597 (N_24597,N_23408,N_23046);
xor U24598 (N_24598,N_22986,N_23632);
nor U24599 (N_24599,N_23927,N_23606);
nor U24600 (N_24600,N_23897,N_23546);
xnor U24601 (N_24601,N_23228,N_23803);
xor U24602 (N_24602,N_23717,N_23496);
xor U24603 (N_24603,N_23560,N_23548);
and U24604 (N_24604,N_22700,N_23679);
xor U24605 (N_24605,N_23364,N_23696);
and U24606 (N_24606,N_22743,N_23420);
nor U24607 (N_24607,N_23155,N_23164);
or U24608 (N_24608,N_23988,N_23798);
xor U24609 (N_24609,N_22524,N_22501);
nand U24610 (N_24610,N_22693,N_23373);
or U24611 (N_24611,N_22936,N_23473);
xnor U24612 (N_24612,N_22886,N_23358);
or U24613 (N_24613,N_23705,N_23256);
nand U24614 (N_24614,N_22537,N_23918);
and U24615 (N_24615,N_22798,N_23002);
and U24616 (N_24616,N_23226,N_23905);
or U24617 (N_24617,N_23339,N_23636);
and U24618 (N_24618,N_22546,N_22574);
nor U24619 (N_24619,N_22925,N_22825);
nor U24620 (N_24620,N_23830,N_23057);
and U24621 (N_24621,N_22645,N_23482);
nor U24622 (N_24622,N_22809,N_22970);
and U24623 (N_24623,N_22786,N_23687);
or U24624 (N_24624,N_23894,N_23251);
or U24625 (N_24625,N_23602,N_23785);
and U24626 (N_24626,N_23870,N_23350);
and U24627 (N_24627,N_23178,N_23241);
and U24628 (N_24628,N_23525,N_23822);
and U24629 (N_24629,N_23177,N_22949);
or U24630 (N_24630,N_23633,N_23012);
or U24631 (N_24631,N_22726,N_23935);
nor U24632 (N_24632,N_23467,N_22551);
nand U24633 (N_24633,N_22893,N_23465);
and U24634 (N_24634,N_23824,N_23080);
and U24635 (N_24635,N_23836,N_23820);
xor U24636 (N_24636,N_22943,N_22604);
and U24637 (N_24637,N_23613,N_23088);
nor U24638 (N_24638,N_23436,N_23007);
and U24639 (N_24639,N_22838,N_23109);
or U24640 (N_24640,N_23278,N_23937);
nand U24641 (N_24641,N_23831,N_22689);
nand U24642 (N_24642,N_23581,N_22861);
nand U24643 (N_24643,N_22811,N_23848);
nand U24644 (N_24644,N_23804,N_23749);
nor U24645 (N_24645,N_23614,N_23098);
nand U24646 (N_24646,N_23523,N_23210);
and U24647 (N_24647,N_22601,N_23078);
or U24648 (N_24648,N_23067,N_23557);
or U24649 (N_24649,N_22741,N_23823);
nand U24650 (N_24650,N_23911,N_23825);
nand U24651 (N_24651,N_22561,N_23881);
and U24652 (N_24652,N_22672,N_22625);
xor U24653 (N_24653,N_23799,N_22762);
or U24654 (N_24654,N_23315,N_22620);
and U24655 (N_24655,N_23383,N_23153);
nand U24656 (N_24656,N_23787,N_23857);
xor U24657 (N_24657,N_23889,N_23757);
nor U24658 (N_24658,N_22890,N_23125);
nand U24659 (N_24659,N_23393,N_23414);
or U24660 (N_24660,N_22846,N_23454);
nor U24661 (N_24661,N_23332,N_23891);
nand U24662 (N_24662,N_23767,N_22656);
nand U24663 (N_24663,N_23762,N_23470);
xnor U24664 (N_24664,N_22832,N_22856);
nor U24665 (N_24665,N_22644,N_23013);
nand U24666 (N_24666,N_22829,N_23382);
nand U24667 (N_24667,N_23242,N_23298);
nand U24668 (N_24668,N_23625,N_23137);
or U24669 (N_24669,N_22589,N_23422);
nor U24670 (N_24670,N_22939,N_23379);
xor U24671 (N_24671,N_23022,N_23448);
nor U24672 (N_24672,N_23550,N_23259);
nor U24673 (N_24673,N_23886,N_23571);
nand U24674 (N_24674,N_23168,N_23460);
nand U24675 (N_24675,N_23264,N_23868);
xnor U24676 (N_24676,N_23199,N_22595);
nor U24677 (N_24677,N_23246,N_23075);
xnor U24678 (N_24678,N_23071,N_23966);
xor U24679 (N_24679,N_23771,N_23376);
nand U24680 (N_24680,N_23554,N_23238);
or U24681 (N_24681,N_22791,N_23074);
and U24682 (N_24682,N_22896,N_23400);
nor U24683 (N_24683,N_23189,N_23710);
xor U24684 (N_24684,N_23479,N_22616);
nand U24685 (N_24685,N_23595,N_23732);
or U24686 (N_24686,N_22867,N_23863);
or U24687 (N_24687,N_22715,N_22663);
or U24688 (N_24688,N_22558,N_23084);
nor U24689 (N_24689,N_22535,N_23540);
nor U24690 (N_24690,N_23539,N_23099);
or U24691 (N_24691,N_22723,N_23921);
nor U24692 (N_24692,N_23232,N_23318);
nand U24693 (N_24693,N_23624,N_22927);
nand U24694 (N_24694,N_22564,N_23185);
xnor U24695 (N_24695,N_23387,N_23867);
and U24696 (N_24696,N_22611,N_23183);
nor U24697 (N_24697,N_22788,N_22800);
or U24698 (N_24698,N_23165,N_22679);
or U24699 (N_24699,N_23508,N_23694);
or U24700 (N_24700,N_23611,N_23443);
xnor U24701 (N_24701,N_23871,N_22758);
or U24702 (N_24702,N_23774,N_22868);
or U24703 (N_24703,N_23963,N_23699);
or U24704 (N_24704,N_22859,N_22655);
xor U24705 (N_24705,N_23019,N_23514);
nor U24706 (N_24706,N_22649,N_23317);
nand U24707 (N_24707,N_23450,N_22834);
and U24708 (N_24708,N_22544,N_23744);
xor U24709 (N_24709,N_23574,N_22807);
and U24710 (N_24710,N_23668,N_23524);
nand U24711 (N_24711,N_22877,N_23392);
and U24712 (N_24712,N_23368,N_22696);
and U24713 (N_24713,N_22605,N_23362);
and U24714 (N_24714,N_22858,N_23471);
nor U24715 (N_24715,N_22913,N_23953);
xor U24716 (N_24716,N_23227,N_22862);
or U24717 (N_24717,N_23090,N_23968);
nor U24718 (N_24718,N_23260,N_23598);
nor U24719 (N_24719,N_23356,N_23381);
xor U24720 (N_24720,N_23944,N_23838);
or U24721 (N_24721,N_23923,N_23616);
or U24722 (N_24722,N_22895,N_23491);
xnor U24723 (N_24723,N_22996,N_23517);
nor U24724 (N_24724,N_23195,N_22748);
nand U24725 (N_24725,N_22946,N_22770);
xnor U24726 (N_24726,N_23843,N_23960);
nand U24727 (N_24727,N_23437,N_22764);
xor U24728 (N_24728,N_23310,N_23522);
nor U24729 (N_24729,N_22979,N_23500);
nand U24730 (N_24730,N_22543,N_22985);
xor U24731 (N_24731,N_23573,N_22808);
xor U24732 (N_24732,N_23043,N_23146);
or U24733 (N_24733,N_22793,N_23599);
and U24734 (N_24734,N_22593,N_23235);
nor U24735 (N_24735,N_22976,N_23513);
nand U24736 (N_24736,N_22619,N_23261);
nor U24737 (N_24737,N_22965,N_23959);
xnor U24738 (N_24738,N_23756,N_23509);
and U24739 (N_24739,N_23156,N_22742);
xor U24740 (N_24740,N_22725,N_22934);
nand U24741 (N_24741,N_23059,N_23861);
and U24742 (N_24742,N_23374,N_22708);
nand U24743 (N_24743,N_23281,N_23753);
xor U24744 (N_24744,N_23286,N_23764);
xor U24745 (N_24745,N_23856,N_23648);
or U24746 (N_24746,N_23681,N_23037);
or U24747 (N_24747,N_23520,N_22684);
nand U24748 (N_24748,N_22653,N_22906);
or U24749 (N_24749,N_23456,N_22827);
xor U24750 (N_24750,N_22593,N_23443);
nand U24751 (N_24751,N_22885,N_23849);
nor U24752 (N_24752,N_23179,N_23127);
nor U24753 (N_24753,N_23843,N_22824);
nor U24754 (N_24754,N_22736,N_22716);
and U24755 (N_24755,N_23817,N_23688);
nand U24756 (N_24756,N_23136,N_23822);
nor U24757 (N_24757,N_23189,N_22726);
or U24758 (N_24758,N_22512,N_22675);
and U24759 (N_24759,N_23113,N_23418);
and U24760 (N_24760,N_22616,N_22899);
or U24761 (N_24761,N_22989,N_23689);
nand U24762 (N_24762,N_22563,N_23425);
xnor U24763 (N_24763,N_23465,N_22827);
nand U24764 (N_24764,N_22694,N_22869);
nand U24765 (N_24765,N_23138,N_23496);
xor U24766 (N_24766,N_23243,N_22970);
and U24767 (N_24767,N_23260,N_23360);
or U24768 (N_24768,N_23884,N_22587);
or U24769 (N_24769,N_23179,N_23944);
or U24770 (N_24770,N_22992,N_23213);
xor U24771 (N_24771,N_22914,N_23229);
nand U24772 (N_24772,N_23989,N_23742);
xnor U24773 (N_24773,N_23761,N_22861);
nand U24774 (N_24774,N_22878,N_22860);
and U24775 (N_24775,N_23555,N_22643);
or U24776 (N_24776,N_23558,N_23944);
nand U24777 (N_24777,N_23236,N_22682);
nor U24778 (N_24778,N_23566,N_23405);
nand U24779 (N_24779,N_23755,N_23215);
xor U24780 (N_24780,N_22973,N_23283);
or U24781 (N_24781,N_22794,N_23381);
nor U24782 (N_24782,N_22878,N_22976);
and U24783 (N_24783,N_22959,N_23942);
and U24784 (N_24784,N_23404,N_23793);
and U24785 (N_24785,N_22951,N_23254);
and U24786 (N_24786,N_22574,N_23416);
nor U24787 (N_24787,N_23902,N_23198);
or U24788 (N_24788,N_22526,N_23126);
or U24789 (N_24789,N_22653,N_23036);
nor U24790 (N_24790,N_23398,N_23454);
nand U24791 (N_24791,N_23456,N_22589);
or U24792 (N_24792,N_22974,N_22637);
xnor U24793 (N_24793,N_23377,N_23630);
xnor U24794 (N_24794,N_23894,N_22796);
or U24795 (N_24795,N_22650,N_23414);
nor U24796 (N_24796,N_23006,N_22506);
nor U24797 (N_24797,N_22734,N_23430);
and U24798 (N_24798,N_23136,N_23131);
nand U24799 (N_24799,N_23923,N_23873);
xnor U24800 (N_24800,N_23833,N_23491);
nand U24801 (N_24801,N_23819,N_23234);
and U24802 (N_24802,N_23304,N_23764);
nand U24803 (N_24803,N_23127,N_23690);
nand U24804 (N_24804,N_22824,N_22745);
and U24805 (N_24805,N_23780,N_23744);
xnor U24806 (N_24806,N_23841,N_22957);
and U24807 (N_24807,N_23977,N_23983);
or U24808 (N_24808,N_22516,N_22913);
nor U24809 (N_24809,N_23017,N_22917);
or U24810 (N_24810,N_23641,N_23980);
xnor U24811 (N_24811,N_23171,N_23077);
and U24812 (N_24812,N_22539,N_22826);
xnor U24813 (N_24813,N_23487,N_23793);
nor U24814 (N_24814,N_23004,N_23293);
nor U24815 (N_24815,N_23911,N_23190);
and U24816 (N_24816,N_22774,N_23293);
or U24817 (N_24817,N_23292,N_23478);
and U24818 (N_24818,N_23578,N_23715);
and U24819 (N_24819,N_23805,N_23098);
or U24820 (N_24820,N_22911,N_23964);
xnor U24821 (N_24821,N_22847,N_23270);
and U24822 (N_24822,N_23020,N_22932);
nor U24823 (N_24823,N_23610,N_22587);
xor U24824 (N_24824,N_23973,N_23985);
nor U24825 (N_24825,N_22547,N_22795);
nor U24826 (N_24826,N_23484,N_22849);
xor U24827 (N_24827,N_23334,N_23692);
nor U24828 (N_24828,N_23892,N_23045);
and U24829 (N_24829,N_22998,N_22884);
and U24830 (N_24830,N_22921,N_23873);
nand U24831 (N_24831,N_23826,N_23991);
nand U24832 (N_24832,N_22821,N_23175);
nand U24833 (N_24833,N_23265,N_23942);
nor U24834 (N_24834,N_23938,N_23950);
nor U24835 (N_24835,N_23048,N_23241);
and U24836 (N_24836,N_22525,N_23293);
xor U24837 (N_24837,N_23860,N_23144);
nand U24838 (N_24838,N_23466,N_23456);
and U24839 (N_24839,N_23979,N_23571);
and U24840 (N_24840,N_23790,N_23403);
nor U24841 (N_24841,N_22877,N_23481);
nand U24842 (N_24842,N_23748,N_23131);
nor U24843 (N_24843,N_23473,N_22817);
nor U24844 (N_24844,N_22540,N_23273);
xor U24845 (N_24845,N_22660,N_23521);
xnor U24846 (N_24846,N_22945,N_23098);
xnor U24847 (N_24847,N_23098,N_23915);
or U24848 (N_24848,N_22593,N_23897);
nand U24849 (N_24849,N_23927,N_23093);
xor U24850 (N_24850,N_23419,N_22628);
nor U24851 (N_24851,N_23596,N_22908);
and U24852 (N_24852,N_22965,N_23645);
and U24853 (N_24853,N_23555,N_23148);
nor U24854 (N_24854,N_23238,N_23142);
nor U24855 (N_24855,N_23107,N_23670);
and U24856 (N_24856,N_22558,N_23840);
xor U24857 (N_24857,N_23756,N_22882);
or U24858 (N_24858,N_23471,N_22924);
nor U24859 (N_24859,N_23788,N_23756);
nor U24860 (N_24860,N_22856,N_23099);
nor U24861 (N_24861,N_23662,N_23221);
or U24862 (N_24862,N_23482,N_23866);
or U24863 (N_24863,N_23028,N_23034);
nand U24864 (N_24864,N_23171,N_23954);
or U24865 (N_24865,N_23846,N_22859);
or U24866 (N_24866,N_23888,N_23097);
nor U24867 (N_24867,N_22777,N_23240);
xor U24868 (N_24868,N_23134,N_23878);
and U24869 (N_24869,N_22746,N_23946);
and U24870 (N_24870,N_23226,N_22709);
nand U24871 (N_24871,N_23571,N_22642);
or U24872 (N_24872,N_23069,N_23852);
xnor U24873 (N_24873,N_23908,N_23745);
and U24874 (N_24874,N_23339,N_23052);
and U24875 (N_24875,N_23721,N_22983);
xnor U24876 (N_24876,N_23692,N_23661);
xor U24877 (N_24877,N_23620,N_23173);
nor U24878 (N_24878,N_23297,N_22755);
or U24879 (N_24879,N_22961,N_23946);
or U24880 (N_24880,N_22723,N_22923);
xnor U24881 (N_24881,N_23582,N_23335);
nand U24882 (N_24882,N_23838,N_22883);
xnor U24883 (N_24883,N_22915,N_23620);
or U24884 (N_24884,N_23061,N_23253);
or U24885 (N_24885,N_23154,N_22714);
and U24886 (N_24886,N_23764,N_23330);
nand U24887 (N_24887,N_23222,N_23871);
xnor U24888 (N_24888,N_22537,N_22662);
and U24889 (N_24889,N_22586,N_23162);
xor U24890 (N_24890,N_23079,N_22741);
or U24891 (N_24891,N_23518,N_23746);
nor U24892 (N_24892,N_22928,N_23641);
xnor U24893 (N_24893,N_22763,N_23385);
and U24894 (N_24894,N_23748,N_22928);
nand U24895 (N_24895,N_22592,N_22598);
or U24896 (N_24896,N_23763,N_22689);
and U24897 (N_24897,N_22601,N_22649);
xor U24898 (N_24898,N_23106,N_22697);
xnor U24899 (N_24899,N_23875,N_23126);
xnor U24900 (N_24900,N_23182,N_23749);
and U24901 (N_24901,N_23845,N_22691);
nand U24902 (N_24902,N_23064,N_23003);
or U24903 (N_24903,N_23624,N_23433);
nand U24904 (N_24904,N_22863,N_23875);
and U24905 (N_24905,N_23524,N_22602);
nand U24906 (N_24906,N_22954,N_22640);
or U24907 (N_24907,N_22855,N_23898);
xnor U24908 (N_24908,N_22927,N_23646);
xor U24909 (N_24909,N_23750,N_22598);
and U24910 (N_24910,N_23996,N_22962);
nand U24911 (N_24911,N_23931,N_23600);
nor U24912 (N_24912,N_23331,N_22975);
or U24913 (N_24913,N_23463,N_23126);
nand U24914 (N_24914,N_23711,N_23196);
nor U24915 (N_24915,N_23785,N_22548);
xnor U24916 (N_24916,N_23698,N_23092);
nand U24917 (N_24917,N_23388,N_23100);
nor U24918 (N_24918,N_22944,N_23717);
xor U24919 (N_24919,N_23424,N_22710);
nor U24920 (N_24920,N_23018,N_23966);
and U24921 (N_24921,N_22587,N_22610);
and U24922 (N_24922,N_22651,N_23585);
nand U24923 (N_24923,N_23199,N_22696);
nor U24924 (N_24924,N_23246,N_22885);
nand U24925 (N_24925,N_22526,N_22576);
nor U24926 (N_24926,N_23763,N_23313);
or U24927 (N_24927,N_23341,N_23936);
xor U24928 (N_24928,N_22948,N_23332);
xnor U24929 (N_24929,N_22551,N_23915);
xor U24930 (N_24930,N_22997,N_23733);
and U24931 (N_24931,N_23744,N_22821);
xor U24932 (N_24932,N_22992,N_23820);
and U24933 (N_24933,N_23697,N_23070);
and U24934 (N_24934,N_23882,N_23457);
nand U24935 (N_24935,N_23969,N_23759);
or U24936 (N_24936,N_23761,N_22637);
and U24937 (N_24937,N_23236,N_22635);
xnor U24938 (N_24938,N_23649,N_23808);
nor U24939 (N_24939,N_23263,N_23699);
nand U24940 (N_24940,N_22849,N_22810);
and U24941 (N_24941,N_22540,N_22937);
xnor U24942 (N_24942,N_22864,N_22605);
nand U24943 (N_24943,N_22658,N_23927);
nand U24944 (N_24944,N_23958,N_23424);
or U24945 (N_24945,N_22701,N_23757);
xor U24946 (N_24946,N_22848,N_22970);
or U24947 (N_24947,N_22726,N_23270);
nand U24948 (N_24948,N_22569,N_22583);
or U24949 (N_24949,N_23881,N_22946);
nand U24950 (N_24950,N_23023,N_23425);
nor U24951 (N_24951,N_23297,N_23096);
xor U24952 (N_24952,N_23292,N_23796);
xnor U24953 (N_24953,N_23308,N_22954);
or U24954 (N_24954,N_23882,N_22943);
xnor U24955 (N_24955,N_22654,N_23957);
nand U24956 (N_24956,N_23220,N_23468);
or U24957 (N_24957,N_22561,N_22601);
or U24958 (N_24958,N_23655,N_23584);
or U24959 (N_24959,N_23452,N_23538);
xnor U24960 (N_24960,N_23092,N_23235);
nand U24961 (N_24961,N_23362,N_22572);
xnor U24962 (N_24962,N_22519,N_23490);
nand U24963 (N_24963,N_23269,N_22829);
nor U24964 (N_24964,N_23584,N_22729);
and U24965 (N_24965,N_23435,N_23456);
or U24966 (N_24966,N_23017,N_23115);
nor U24967 (N_24967,N_22553,N_22769);
xnor U24968 (N_24968,N_23804,N_23201);
nor U24969 (N_24969,N_23500,N_22912);
nor U24970 (N_24970,N_23173,N_23181);
nand U24971 (N_24971,N_22890,N_23917);
nand U24972 (N_24972,N_22928,N_22960);
xnor U24973 (N_24973,N_23671,N_22656);
and U24974 (N_24974,N_23996,N_23139);
nand U24975 (N_24975,N_23501,N_22579);
nor U24976 (N_24976,N_23865,N_23036);
nand U24977 (N_24977,N_23925,N_23018);
nand U24978 (N_24978,N_23071,N_22871);
nand U24979 (N_24979,N_22823,N_22831);
and U24980 (N_24980,N_23086,N_22642);
nand U24981 (N_24981,N_22768,N_23651);
and U24982 (N_24982,N_23822,N_23208);
or U24983 (N_24983,N_23961,N_23598);
nand U24984 (N_24984,N_22597,N_23526);
xor U24985 (N_24985,N_22740,N_22802);
nor U24986 (N_24986,N_23694,N_23384);
and U24987 (N_24987,N_22861,N_23302);
xor U24988 (N_24988,N_22747,N_23556);
or U24989 (N_24989,N_23923,N_22907);
nor U24990 (N_24990,N_22521,N_23578);
xor U24991 (N_24991,N_23684,N_22701);
xnor U24992 (N_24992,N_23981,N_22823);
xnor U24993 (N_24993,N_23482,N_23637);
nor U24994 (N_24994,N_23569,N_23101);
or U24995 (N_24995,N_23070,N_22579);
and U24996 (N_24996,N_23138,N_22732);
xnor U24997 (N_24997,N_22862,N_23338);
or U24998 (N_24998,N_22657,N_23478);
nor U24999 (N_24999,N_23782,N_23169);
nor U25000 (N_25000,N_23674,N_23012);
and U25001 (N_25001,N_22516,N_22546);
xor U25002 (N_25002,N_22678,N_22848);
or U25003 (N_25003,N_23348,N_22723);
nor U25004 (N_25004,N_22567,N_23913);
and U25005 (N_25005,N_23829,N_23621);
and U25006 (N_25006,N_22772,N_23546);
nor U25007 (N_25007,N_23364,N_22546);
nor U25008 (N_25008,N_23381,N_23035);
and U25009 (N_25009,N_23126,N_22923);
nor U25010 (N_25010,N_23034,N_23903);
and U25011 (N_25011,N_23842,N_23501);
nor U25012 (N_25012,N_23111,N_23665);
nor U25013 (N_25013,N_22517,N_23829);
nor U25014 (N_25014,N_22897,N_23914);
nand U25015 (N_25015,N_22994,N_23306);
and U25016 (N_25016,N_23844,N_22751);
and U25017 (N_25017,N_23772,N_23137);
and U25018 (N_25018,N_22806,N_23862);
or U25019 (N_25019,N_23753,N_23690);
xor U25020 (N_25020,N_23736,N_23162);
and U25021 (N_25021,N_22538,N_22801);
xor U25022 (N_25022,N_23394,N_23289);
xnor U25023 (N_25023,N_23711,N_23971);
xor U25024 (N_25024,N_23263,N_23777);
and U25025 (N_25025,N_22986,N_22505);
or U25026 (N_25026,N_22505,N_23441);
nand U25027 (N_25027,N_22859,N_22932);
or U25028 (N_25028,N_23593,N_23127);
xnor U25029 (N_25029,N_23024,N_23857);
and U25030 (N_25030,N_22722,N_22788);
or U25031 (N_25031,N_23747,N_22542);
or U25032 (N_25032,N_23901,N_22742);
or U25033 (N_25033,N_23365,N_22745);
xor U25034 (N_25034,N_23079,N_23930);
nor U25035 (N_25035,N_23158,N_23911);
nand U25036 (N_25036,N_22785,N_23280);
and U25037 (N_25037,N_23918,N_23543);
nor U25038 (N_25038,N_23057,N_23383);
and U25039 (N_25039,N_23314,N_23814);
or U25040 (N_25040,N_22622,N_22765);
or U25041 (N_25041,N_23536,N_23171);
and U25042 (N_25042,N_22565,N_23727);
xnor U25043 (N_25043,N_22744,N_23448);
nand U25044 (N_25044,N_23252,N_22835);
nand U25045 (N_25045,N_23453,N_23125);
nor U25046 (N_25046,N_23577,N_23979);
and U25047 (N_25047,N_23718,N_23723);
and U25048 (N_25048,N_23076,N_22705);
nand U25049 (N_25049,N_22946,N_22862);
nor U25050 (N_25050,N_23528,N_22877);
xnor U25051 (N_25051,N_23822,N_23620);
xor U25052 (N_25052,N_23974,N_23465);
or U25053 (N_25053,N_23256,N_23950);
nor U25054 (N_25054,N_23586,N_22836);
nor U25055 (N_25055,N_23401,N_23309);
nor U25056 (N_25056,N_23876,N_23991);
nor U25057 (N_25057,N_23455,N_23923);
nor U25058 (N_25058,N_23933,N_23453);
nor U25059 (N_25059,N_22625,N_23175);
nand U25060 (N_25060,N_23159,N_22702);
and U25061 (N_25061,N_23917,N_23970);
and U25062 (N_25062,N_22597,N_23801);
xnor U25063 (N_25063,N_22718,N_23737);
or U25064 (N_25064,N_23319,N_23450);
nor U25065 (N_25065,N_23102,N_23192);
and U25066 (N_25066,N_23440,N_23661);
and U25067 (N_25067,N_23817,N_23323);
nand U25068 (N_25068,N_23754,N_22511);
nand U25069 (N_25069,N_22843,N_22750);
or U25070 (N_25070,N_23429,N_23144);
nor U25071 (N_25071,N_22950,N_23249);
and U25072 (N_25072,N_23818,N_23587);
or U25073 (N_25073,N_23658,N_22968);
and U25074 (N_25074,N_23012,N_23913);
and U25075 (N_25075,N_23821,N_22819);
or U25076 (N_25076,N_23866,N_22639);
xnor U25077 (N_25077,N_23435,N_23501);
nand U25078 (N_25078,N_22829,N_23438);
or U25079 (N_25079,N_22853,N_23698);
or U25080 (N_25080,N_22995,N_23180);
or U25081 (N_25081,N_23848,N_22556);
or U25082 (N_25082,N_23948,N_23859);
and U25083 (N_25083,N_22972,N_23245);
or U25084 (N_25084,N_22553,N_23032);
or U25085 (N_25085,N_23581,N_23600);
xnor U25086 (N_25086,N_22757,N_23989);
nor U25087 (N_25087,N_23675,N_23205);
and U25088 (N_25088,N_23320,N_23822);
and U25089 (N_25089,N_22887,N_23738);
nor U25090 (N_25090,N_23273,N_23794);
nand U25091 (N_25091,N_23374,N_23059);
nor U25092 (N_25092,N_22934,N_23556);
or U25093 (N_25093,N_23953,N_23732);
and U25094 (N_25094,N_23191,N_23908);
nor U25095 (N_25095,N_23627,N_22979);
and U25096 (N_25096,N_23694,N_23726);
xnor U25097 (N_25097,N_22779,N_23053);
nor U25098 (N_25098,N_23250,N_22792);
xor U25099 (N_25099,N_23427,N_23165);
nor U25100 (N_25100,N_23090,N_23437);
nand U25101 (N_25101,N_23696,N_22541);
xor U25102 (N_25102,N_23359,N_23220);
nand U25103 (N_25103,N_23086,N_23952);
xnor U25104 (N_25104,N_23633,N_23612);
or U25105 (N_25105,N_22644,N_23245);
nand U25106 (N_25106,N_23990,N_23538);
nand U25107 (N_25107,N_23363,N_23139);
xor U25108 (N_25108,N_23270,N_23645);
and U25109 (N_25109,N_23786,N_23586);
nand U25110 (N_25110,N_23587,N_23747);
nand U25111 (N_25111,N_23887,N_23961);
nor U25112 (N_25112,N_23957,N_23834);
or U25113 (N_25113,N_23849,N_23895);
xnor U25114 (N_25114,N_23273,N_23718);
nand U25115 (N_25115,N_23418,N_23268);
nand U25116 (N_25116,N_23640,N_23449);
xnor U25117 (N_25117,N_23126,N_23754);
xor U25118 (N_25118,N_22551,N_22656);
or U25119 (N_25119,N_23307,N_22845);
xnor U25120 (N_25120,N_23985,N_22886);
xor U25121 (N_25121,N_23817,N_22592);
nand U25122 (N_25122,N_23099,N_23990);
nand U25123 (N_25123,N_23622,N_23922);
and U25124 (N_25124,N_22554,N_23221);
nor U25125 (N_25125,N_23670,N_22616);
nor U25126 (N_25126,N_23712,N_22606);
or U25127 (N_25127,N_22914,N_23064);
nand U25128 (N_25128,N_23165,N_23470);
and U25129 (N_25129,N_23044,N_23747);
xnor U25130 (N_25130,N_23355,N_23300);
nor U25131 (N_25131,N_23719,N_22850);
or U25132 (N_25132,N_23978,N_22582);
nor U25133 (N_25133,N_23856,N_22523);
nor U25134 (N_25134,N_23909,N_23564);
nand U25135 (N_25135,N_23506,N_22831);
nor U25136 (N_25136,N_23484,N_23153);
nor U25137 (N_25137,N_23163,N_23823);
or U25138 (N_25138,N_22579,N_23001);
nor U25139 (N_25139,N_22533,N_23741);
and U25140 (N_25140,N_22538,N_23082);
nor U25141 (N_25141,N_23694,N_23816);
or U25142 (N_25142,N_23926,N_23116);
nor U25143 (N_25143,N_23583,N_23236);
nor U25144 (N_25144,N_23753,N_23088);
nor U25145 (N_25145,N_22684,N_23580);
nor U25146 (N_25146,N_23721,N_22808);
nor U25147 (N_25147,N_23334,N_23740);
nor U25148 (N_25148,N_23942,N_22977);
xnor U25149 (N_25149,N_23545,N_23571);
nor U25150 (N_25150,N_23331,N_22686);
nand U25151 (N_25151,N_23677,N_23938);
xnor U25152 (N_25152,N_22563,N_22705);
nand U25153 (N_25153,N_22677,N_23242);
xor U25154 (N_25154,N_23658,N_23525);
xnor U25155 (N_25155,N_23128,N_23809);
xnor U25156 (N_25156,N_22589,N_23350);
or U25157 (N_25157,N_22575,N_22902);
nand U25158 (N_25158,N_22886,N_22717);
nand U25159 (N_25159,N_23200,N_23633);
and U25160 (N_25160,N_22678,N_22972);
and U25161 (N_25161,N_23468,N_22927);
or U25162 (N_25162,N_22987,N_23912);
nor U25163 (N_25163,N_23141,N_22882);
nand U25164 (N_25164,N_22910,N_22943);
nand U25165 (N_25165,N_22949,N_22609);
xor U25166 (N_25166,N_23735,N_23292);
nor U25167 (N_25167,N_23300,N_23874);
or U25168 (N_25168,N_23380,N_23068);
xor U25169 (N_25169,N_23276,N_23969);
or U25170 (N_25170,N_22893,N_22703);
and U25171 (N_25171,N_23053,N_23141);
xor U25172 (N_25172,N_23302,N_23126);
nor U25173 (N_25173,N_23657,N_22738);
xnor U25174 (N_25174,N_22776,N_23692);
or U25175 (N_25175,N_23353,N_23345);
or U25176 (N_25176,N_23663,N_23095);
nor U25177 (N_25177,N_22982,N_22723);
nand U25178 (N_25178,N_23568,N_23637);
or U25179 (N_25179,N_23266,N_23190);
xor U25180 (N_25180,N_23732,N_23341);
nand U25181 (N_25181,N_23591,N_23973);
or U25182 (N_25182,N_22641,N_23141);
xnor U25183 (N_25183,N_23638,N_23292);
nand U25184 (N_25184,N_23816,N_23565);
or U25185 (N_25185,N_23249,N_23647);
nor U25186 (N_25186,N_23319,N_23754);
nand U25187 (N_25187,N_22918,N_23511);
or U25188 (N_25188,N_23686,N_22662);
xnor U25189 (N_25189,N_23608,N_22876);
nor U25190 (N_25190,N_23542,N_23254);
nor U25191 (N_25191,N_22565,N_23685);
nand U25192 (N_25192,N_23752,N_22644);
and U25193 (N_25193,N_22601,N_22753);
or U25194 (N_25194,N_23327,N_23995);
or U25195 (N_25195,N_22694,N_22856);
xnor U25196 (N_25196,N_23912,N_22535);
nand U25197 (N_25197,N_23230,N_22600);
or U25198 (N_25198,N_23499,N_23465);
nor U25199 (N_25199,N_23765,N_22723);
and U25200 (N_25200,N_23495,N_22696);
or U25201 (N_25201,N_23344,N_23646);
or U25202 (N_25202,N_23533,N_23983);
and U25203 (N_25203,N_23423,N_23282);
nand U25204 (N_25204,N_23155,N_23067);
xnor U25205 (N_25205,N_23208,N_22948);
xor U25206 (N_25206,N_23691,N_23422);
or U25207 (N_25207,N_22927,N_22639);
nor U25208 (N_25208,N_23398,N_23773);
nor U25209 (N_25209,N_23758,N_22536);
nor U25210 (N_25210,N_22505,N_22995);
xor U25211 (N_25211,N_23411,N_23533);
nand U25212 (N_25212,N_23095,N_23001);
nand U25213 (N_25213,N_23623,N_22505);
or U25214 (N_25214,N_23956,N_23469);
xnor U25215 (N_25215,N_22689,N_23192);
nor U25216 (N_25216,N_22886,N_23045);
xor U25217 (N_25217,N_23115,N_23682);
nand U25218 (N_25218,N_23830,N_23374);
xor U25219 (N_25219,N_22922,N_22619);
nand U25220 (N_25220,N_23839,N_22911);
nor U25221 (N_25221,N_23990,N_23573);
xor U25222 (N_25222,N_23420,N_23236);
nor U25223 (N_25223,N_22558,N_23269);
nand U25224 (N_25224,N_23792,N_23750);
or U25225 (N_25225,N_23203,N_23765);
nor U25226 (N_25226,N_23105,N_23296);
or U25227 (N_25227,N_23716,N_22788);
and U25228 (N_25228,N_23932,N_22739);
and U25229 (N_25229,N_23839,N_22501);
nand U25230 (N_25230,N_22559,N_23750);
or U25231 (N_25231,N_22763,N_23843);
or U25232 (N_25232,N_23481,N_23340);
nor U25233 (N_25233,N_22876,N_22739);
nand U25234 (N_25234,N_23831,N_23240);
xnor U25235 (N_25235,N_22998,N_22653);
xor U25236 (N_25236,N_22897,N_23702);
nor U25237 (N_25237,N_23566,N_23337);
nor U25238 (N_25238,N_23025,N_22784);
and U25239 (N_25239,N_23248,N_23122);
or U25240 (N_25240,N_23610,N_22822);
nand U25241 (N_25241,N_22821,N_23323);
and U25242 (N_25242,N_23553,N_22875);
nand U25243 (N_25243,N_23547,N_22679);
xor U25244 (N_25244,N_23349,N_22744);
and U25245 (N_25245,N_22712,N_22529);
nor U25246 (N_25246,N_23968,N_22800);
nand U25247 (N_25247,N_23282,N_22596);
and U25248 (N_25248,N_22663,N_23655);
and U25249 (N_25249,N_23190,N_23740);
and U25250 (N_25250,N_23614,N_23921);
nand U25251 (N_25251,N_22803,N_23378);
nand U25252 (N_25252,N_22703,N_23059);
and U25253 (N_25253,N_23402,N_23319);
nor U25254 (N_25254,N_23434,N_23001);
or U25255 (N_25255,N_23486,N_22727);
or U25256 (N_25256,N_22720,N_23340);
nor U25257 (N_25257,N_23127,N_23097);
and U25258 (N_25258,N_23798,N_23569);
and U25259 (N_25259,N_23475,N_23105);
and U25260 (N_25260,N_23953,N_23357);
or U25261 (N_25261,N_23922,N_23071);
nor U25262 (N_25262,N_23172,N_23327);
and U25263 (N_25263,N_22538,N_23158);
or U25264 (N_25264,N_23117,N_23529);
nor U25265 (N_25265,N_23031,N_23102);
xor U25266 (N_25266,N_23523,N_23598);
xnor U25267 (N_25267,N_22942,N_23792);
or U25268 (N_25268,N_23501,N_23421);
nand U25269 (N_25269,N_23501,N_22855);
and U25270 (N_25270,N_23896,N_23385);
nand U25271 (N_25271,N_22873,N_22633);
and U25272 (N_25272,N_23086,N_23439);
or U25273 (N_25273,N_23512,N_23089);
nor U25274 (N_25274,N_22554,N_22601);
and U25275 (N_25275,N_22539,N_23499);
or U25276 (N_25276,N_22795,N_22996);
xor U25277 (N_25277,N_23814,N_23795);
nand U25278 (N_25278,N_23250,N_22850);
or U25279 (N_25279,N_23455,N_23199);
or U25280 (N_25280,N_22646,N_23544);
nand U25281 (N_25281,N_22517,N_23393);
nor U25282 (N_25282,N_23377,N_23178);
nand U25283 (N_25283,N_23923,N_23147);
xor U25284 (N_25284,N_23319,N_23583);
nand U25285 (N_25285,N_22968,N_23485);
xnor U25286 (N_25286,N_23713,N_22599);
xor U25287 (N_25287,N_22762,N_22594);
nand U25288 (N_25288,N_23712,N_23716);
and U25289 (N_25289,N_23353,N_23369);
or U25290 (N_25290,N_23828,N_23838);
and U25291 (N_25291,N_23735,N_22699);
nand U25292 (N_25292,N_22738,N_23109);
nand U25293 (N_25293,N_23045,N_23714);
and U25294 (N_25294,N_23690,N_23040);
and U25295 (N_25295,N_23424,N_23324);
and U25296 (N_25296,N_23698,N_23739);
or U25297 (N_25297,N_23629,N_23439);
or U25298 (N_25298,N_22963,N_23110);
nor U25299 (N_25299,N_22617,N_23542);
and U25300 (N_25300,N_22816,N_22849);
nor U25301 (N_25301,N_23908,N_23735);
xnor U25302 (N_25302,N_22994,N_23105);
and U25303 (N_25303,N_23119,N_23099);
and U25304 (N_25304,N_22827,N_22696);
nor U25305 (N_25305,N_22739,N_23539);
and U25306 (N_25306,N_23277,N_23842);
nor U25307 (N_25307,N_23305,N_23073);
nand U25308 (N_25308,N_22628,N_23378);
nor U25309 (N_25309,N_23069,N_22629);
xor U25310 (N_25310,N_22849,N_22876);
xor U25311 (N_25311,N_22766,N_22727);
or U25312 (N_25312,N_23190,N_23855);
nor U25313 (N_25313,N_22675,N_23297);
nand U25314 (N_25314,N_22836,N_23113);
or U25315 (N_25315,N_22995,N_23064);
and U25316 (N_25316,N_22825,N_23180);
and U25317 (N_25317,N_23301,N_23796);
or U25318 (N_25318,N_22966,N_23732);
nand U25319 (N_25319,N_23269,N_22694);
and U25320 (N_25320,N_23123,N_23052);
xnor U25321 (N_25321,N_23605,N_22922);
nand U25322 (N_25322,N_22506,N_23491);
nor U25323 (N_25323,N_23138,N_23046);
or U25324 (N_25324,N_22865,N_23548);
or U25325 (N_25325,N_22726,N_22811);
and U25326 (N_25326,N_23532,N_23770);
xor U25327 (N_25327,N_23611,N_22648);
or U25328 (N_25328,N_22604,N_23610);
nor U25329 (N_25329,N_23522,N_23091);
nand U25330 (N_25330,N_22732,N_22643);
xnor U25331 (N_25331,N_23528,N_23181);
nor U25332 (N_25332,N_23971,N_23941);
and U25333 (N_25333,N_22983,N_23616);
nor U25334 (N_25334,N_23215,N_22667);
or U25335 (N_25335,N_22890,N_22660);
or U25336 (N_25336,N_23300,N_23120);
nand U25337 (N_25337,N_23149,N_22826);
nand U25338 (N_25338,N_23785,N_22922);
nor U25339 (N_25339,N_22650,N_23961);
nand U25340 (N_25340,N_23376,N_23308);
nor U25341 (N_25341,N_23128,N_23905);
nand U25342 (N_25342,N_23300,N_23421);
nor U25343 (N_25343,N_23071,N_23537);
nor U25344 (N_25344,N_23777,N_22860);
and U25345 (N_25345,N_22945,N_22510);
nand U25346 (N_25346,N_23205,N_22538);
nand U25347 (N_25347,N_23636,N_23671);
or U25348 (N_25348,N_23783,N_23201);
and U25349 (N_25349,N_23526,N_22679);
nor U25350 (N_25350,N_23578,N_23123);
nand U25351 (N_25351,N_23962,N_23685);
xnor U25352 (N_25352,N_22576,N_23507);
and U25353 (N_25353,N_23284,N_22854);
and U25354 (N_25354,N_23285,N_22636);
or U25355 (N_25355,N_23429,N_23066);
and U25356 (N_25356,N_22973,N_22603);
nand U25357 (N_25357,N_22801,N_23412);
nor U25358 (N_25358,N_23778,N_22527);
xor U25359 (N_25359,N_23259,N_23505);
nor U25360 (N_25360,N_23287,N_23085);
nor U25361 (N_25361,N_23791,N_23084);
nand U25362 (N_25362,N_23010,N_22812);
xnor U25363 (N_25363,N_23320,N_23514);
xor U25364 (N_25364,N_23806,N_23781);
or U25365 (N_25365,N_22596,N_23916);
nand U25366 (N_25366,N_23840,N_22899);
xor U25367 (N_25367,N_23671,N_23745);
xnor U25368 (N_25368,N_23357,N_22673);
xor U25369 (N_25369,N_22890,N_23444);
or U25370 (N_25370,N_23764,N_22601);
xor U25371 (N_25371,N_22668,N_23717);
nand U25372 (N_25372,N_22753,N_23505);
nor U25373 (N_25373,N_23749,N_23652);
and U25374 (N_25374,N_23363,N_22942);
or U25375 (N_25375,N_23238,N_23177);
xnor U25376 (N_25376,N_22953,N_22902);
or U25377 (N_25377,N_23280,N_23491);
and U25378 (N_25378,N_23854,N_23778);
nand U25379 (N_25379,N_23816,N_23908);
nor U25380 (N_25380,N_22968,N_23279);
or U25381 (N_25381,N_23408,N_22732);
xnor U25382 (N_25382,N_22565,N_23638);
or U25383 (N_25383,N_23363,N_23159);
nor U25384 (N_25384,N_22965,N_23304);
nor U25385 (N_25385,N_23236,N_22804);
and U25386 (N_25386,N_22891,N_23632);
or U25387 (N_25387,N_23082,N_23330);
nor U25388 (N_25388,N_22862,N_23234);
nor U25389 (N_25389,N_22508,N_22544);
or U25390 (N_25390,N_23857,N_23622);
xnor U25391 (N_25391,N_23435,N_23805);
or U25392 (N_25392,N_23661,N_23932);
and U25393 (N_25393,N_22516,N_23358);
nand U25394 (N_25394,N_23798,N_23354);
and U25395 (N_25395,N_23720,N_23308);
or U25396 (N_25396,N_23739,N_23712);
nand U25397 (N_25397,N_22912,N_23598);
xor U25398 (N_25398,N_23228,N_23905);
nor U25399 (N_25399,N_22883,N_22680);
or U25400 (N_25400,N_23729,N_23591);
nor U25401 (N_25401,N_23018,N_23774);
xnor U25402 (N_25402,N_23885,N_23921);
xnor U25403 (N_25403,N_23695,N_23305);
and U25404 (N_25404,N_23867,N_23588);
or U25405 (N_25405,N_23869,N_23797);
nor U25406 (N_25406,N_23638,N_23834);
nand U25407 (N_25407,N_22769,N_23789);
and U25408 (N_25408,N_23268,N_23534);
nand U25409 (N_25409,N_22801,N_22751);
nor U25410 (N_25410,N_23125,N_23090);
and U25411 (N_25411,N_23860,N_22731);
xnor U25412 (N_25412,N_23886,N_23518);
and U25413 (N_25413,N_23797,N_22501);
or U25414 (N_25414,N_23889,N_22721);
or U25415 (N_25415,N_22635,N_23601);
nor U25416 (N_25416,N_23089,N_23927);
and U25417 (N_25417,N_23575,N_23954);
nor U25418 (N_25418,N_22884,N_23313);
or U25419 (N_25419,N_22991,N_22523);
and U25420 (N_25420,N_23048,N_22827);
and U25421 (N_25421,N_23794,N_23703);
nor U25422 (N_25422,N_23875,N_23371);
or U25423 (N_25423,N_22913,N_22774);
and U25424 (N_25424,N_23465,N_23387);
or U25425 (N_25425,N_22982,N_23410);
and U25426 (N_25426,N_23232,N_22952);
or U25427 (N_25427,N_23049,N_23760);
nor U25428 (N_25428,N_23532,N_23301);
and U25429 (N_25429,N_23799,N_22988);
nand U25430 (N_25430,N_22830,N_23312);
or U25431 (N_25431,N_23838,N_23712);
and U25432 (N_25432,N_23951,N_23263);
nand U25433 (N_25433,N_23680,N_22847);
nor U25434 (N_25434,N_23087,N_23837);
or U25435 (N_25435,N_23607,N_23246);
xor U25436 (N_25436,N_22670,N_23333);
xnor U25437 (N_25437,N_23257,N_23166);
xor U25438 (N_25438,N_23320,N_23353);
xor U25439 (N_25439,N_23822,N_22892);
and U25440 (N_25440,N_23763,N_22561);
nand U25441 (N_25441,N_23859,N_23657);
and U25442 (N_25442,N_22708,N_23729);
xor U25443 (N_25443,N_23108,N_23979);
and U25444 (N_25444,N_22556,N_22627);
nor U25445 (N_25445,N_23254,N_23629);
or U25446 (N_25446,N_23485,N_23909);
nand U25447 (N_25447,N_22567,N_23346);
xnor U25448 (N_25448,N_22655,N_23178);
or U25449 (N_25449,N_23602,N_23402);
and U25450 (N_25450,N_23574,N_23959);
or U25451 (N_25451,N_22698,N_22732);
nor U25452 (N_25452,N_23348,N_23962);
or U25453 (N_25453,N_23306,N_22778);
xnor U25454 (N_25454,N_23064,N_23741);
xnor U25455 (N_25455,N_23556,N_23916);
or U25456 (N_25456,N_23100,N_23271);
nand U25457 (N_25457,N_22801,N_23536);
nand U25458 (N_25458,N_23455,N_23154);
and U25459 (N_25459,N_23639,N_23395);
nand U25460 (N_25460,N_23479,N_23522);
nand U25461 (N_25461,N_23226,N_23538);
and U25462 (N_25462,N_23940,N_22828);
nor U25463 (N_25463,N_22857,N_23775);
nand U25464 (N_25464,N_23442,N_22514);
nand U25465 (N_25465,N_22837,N_22561);
nor U25466 (N_25466,N_23028,N_22824);
nor U25467 (N_25467,N_23070,N_22799);
nand U25468 (N_25468,N_23994,N_22814);
and U25469 (N_25469,N_23504,N_23562);
and U25470 (N_25470,N_23232,N_23113);
xnor U25471 (N_25471,N_23708,N_22568);
nand U25472 (N_25472,N_22616,N_23671);
and U25473 (N_25473,N_23801,N_22852);
nand U25474 (N_25474,N_23836,N_22683);
nand U25475 (N_25475,N_23598,N_23516);
and U25476 (N_25476,N_23896,N_23828);
xnor U25477 (N_25477,N_23946,N_22951);
nand U25478 (N_25478,N_23192,N_23554);
nand U25479 (N_25479,N_22585,N_23761);
nor U25480 (N_25480,N_23916,N_23041);
or U25481 (N_25481,N_23565,N_23140);
nand U25482 (N_25482,N_23968,N_23443);
or U25483 (N_25483,N_23835,N_23337);
nor U25484 (N_25484,N_22788,N_23569);
and U25485 (N_25485,N_22570,N_23664);
nor U25486 (N_25486,N_22928,N_23613);
nand U25487 (N_25487,N_23913,N_23103);
and U25488 (N_25488,N_22686,N_23060);
xnor U25489 (N_25489,N_23834,N_23678);
xor U25490 (N_25490,N_23959,N_23609);
nand U25491 (N_25491,N_23690,N_23632);
and U25492 (N_25492,N_22948,N_23740);
or U25493 (N_25493,N_23750,N_22764);
or U25494 (N_25494,N_23735,N_23368);
nor U25495 (N_25495,N_23676,N_23272);
or U25496 (N_25496,N_22674,N_23816);
or U25497 (N_25497,N_22857,N_22539);
and U25498 (N_25498,N_23288,N_23246);
or U25499 (N_25499,N_23759,N_22728);
or U25500 (N_25500,N_24746,N_24926);
xnor U25501 (N_25501,N_24732,N_25178);
nand U25502 (N_25502,N_24130,N_24395);
or U25503 (N_25503,N_25476,N_25429);
nand U25504 (N_25504,N_24463,N_24689);
nor U25505 (N_25505,N_24427,N_24382);
and U25506 (N_25506,N_24131,N_24919);
and U25507 (N_25507,N_25006,N_25408);
nand U25508 (N_25508,N_24243,N_24607);
and U25509 (N_25509,N_25356,N_24073);
or U25510 (N_25510,N_25053,N_24004);
and U25511 (N_25511,N_24883,N_25139);
nand U25512 (N_25512,N_24629,N_25270);
or U25513 (N_25513,N_25219,N_24314);
or U25514 (N_25514,N_25395,N_24474);
xnor U25515 (N_25515,N_24191,N_24356);
and U25516 (N_25516,N_24285,N_24050);
xor U25517 (N_25517,N_24547,N_25154);
or U25518 (N_25518,N_24240,N_25017);
xor U25519 (N_25519,N_24798,N_25252);
xnor U25520 (N_25520,N_25324,N_24394);
nor U25521 (N_25521,N_24107,N_25097);
and U25522 (N_25522,N_24118,N_24885);
xnor U25523 (N_25523,N_24495,N_24398);
xnor U25524 (N_25524,N_24003,N_24056);
or U25525 (N_25525,N_24088,N_24200);
nand U25526 (N_25526,N_24806,N_24620);
or U25527 (N_25527,N_24670,N_24138);
and U25528 (N_25528,N_24383,N_24949);
or U25529 (N_25529,N_24915,N_25454);
and U25530 (N_25530,N_24319,N_24340);
xor U25531 (N_25531,N_25110,N_24342);
and U25532 (N_25532,N_24709,N_24234);
and U25533 (N_25533,N_25211,N_24735);
and U25534 (N_25534,N_25049,N_24155);
nand U25535 (N_25535,N_24814,N_25182);
nand U25536 (N_25536,N_25285,N_24061);
or U25537 (N_25537,N_24054,N_24454);
xor U25538 (N_25538,N_24065,N_25209);
or U25539 (N_25539,N_24621,N_24533);
or U25540 (N_25540,N_24425,N_24786);
or U25541 (N_25541,N_24146,N_24119);
xnor U25542 (N_25542,N_25308,N_24112);
nand U25543 (N_25543,N_24040,N_25326);
nor U25544 (N_25544,N_24089,N_25045);
and U25545 (N_25545,N_25404,N_24163);
or U25546 (N_25546,N_25119,N_24460);
or U25547 (N_25547,N_24971,N_24470);
nor U25548 (N_25548,N_24106,N_24662);
xor U25549 (N_25549,N_24706,N_25185);
nand U25550 (N_25550,N_24743,N_25137);
nand U25551 (N_25551,N_24142,N_25384);
or U25552 (N_25552,N_24492,N_25321);
nand U25553 (N_25553,N_24766,N_24263);
nor U25554 (N_25554,N_25157,N_24210);
xor U25555 (N_25555,N_25187,N_24668);
nand U25556 (N_25556,N_24473,N_24120);
nand U25557 (N_25557,N_25072,N_24857);
and U25558 (N_25558,N_24811,N_24059);
nor U25559 (N_25559,N_24748,N_25066);
xnor U25560 (N_25560,N_24350,N_24975);
nor U25561 (N_25561,N_25405,N_24080);
nand U25562 (N_25562,N_24630,N_24432);
nor U25563 (N_25563,N_24140,N_24954);
nor U25564 (N_25564,N_24666,N_25189);
or U25565 (N_25565,N_25263,N_25392);
nand U25566 (N_25566,N_25329,N_24468);
nand U25567 (N_25567,N_24204,N_24172);
nand U25568 (N_25568,N_24891,N_24551);
nand U25569 (N_25569,N_24982,N_24197);
nor U25570 (N_25570,N_24440,N_24577);
xor U25571 (N_25571,N_24952,N_25150);
nor U25572 (N_25572,N_24249,N_24956);
nand U25573 (N_25573,N_25244,N_24377);
xnor U25574 (N_25574,N_25215,N_25122);
xor U25575 (N_25575,N_24181,N_25223);
xor U25576 (N_25576,N_24619,N_25192);
and U25577 (N_25577,N_24744,N_24353);
or U25578 (N_25578,N_24755,N_25320);
nor U25579 (N_25579,N_24058,N_24352);
nand U25580 (N_25580,N_25012,N_24438);
xor U25581 (N_25581,N_24888,N_24301);
xnor U25582 (N_25582,N_25010,N_25220);
or U25583 (N_25583,N_24611,N_24967);
and U25584 (N_25584,N_25453,N_24571);
and U25585 (N_25585,N_24946,N_24246);
nor U25586 (N_25586,N_25278,N_24115);
nand U25587 (N_25587,N_24113,N_24305);
nor U25588 (N_25588,N_25333,N_24722);
nand U25589 (N_25589,N_24400,N_25128);
and U25590 (N_25590,N_25355,N_24290);
nand U25591 (N_25591,N_24889,N_24288);
xor U25592 (N_25592,N_24716,N_24169);
xnor U25593 (N_25593,N_25251,N_24677);
nand U25594 (N_25594,N_25338,N_24762);
or U25595 (N_25595,N_25470,N_25120);
and U25596 (N_25596,N_25001,N_25257);
nand U25597 (N_25597,N_25058,N_25009);
xnor U25598 (N_25598,N_24166,N_25465);
nand U25599 (N_25599,N_25156,N_24209);
nor U25600 (N_25600,N_24333,N_24060);
and U25601 (N_25601,N_25485,N_24162);
or U25602 (N_25602,N_24160,N_24918);
xnor U25603 (N_25603,N_24657,N_25024);
xor U25604 (N_25604,N_24020,N_24974);
and U25605 (N_25605,N_24351,N_24963);
and U25606 (N_25606,N_24341,N_24417);
and U25607 (N_25607,N_25094,N_25037);
xnor U25608 (N_25608,N_24594,N_24944);
nand U25609 (N_25609,N_24121,N_25299);
nand U25610 (N_25610,N_24738,N_25241);
xnor U25611 (N_25611,N_24149,N_24126);
nand U25612 (N_25612,N_25048,N_24834);
or U25613 (N_25613,N_24573,N_24220);
and U25614 (N_25614,N_25193,N_25386);
nor U25615 (N_25615,N_25347,N_24075);
or U25616 (N_25616,N_24608,N_24632);
nand U25617 (N_25617,N_24028,N_24000);
nand U25618 (N_25618,N_25246,N_24507);
and U25619 (N_25619,N_24542,N_24094);
and U25620 (N_25620,N_24749,N_24456);
nand U25621 (N_25621,N_25224,N_25147);
or U25622 (N_25622,N_25346,N_25242);
nand U25623 (N_25623,N_24010,N_24252);
nor U25624 (N_25624,N_25231,N_25027);
nand U25625 (N_25625,N_24860,N_24179);
nand U25626 (N_25626,N_25226,N_24816);
or U25627 (N_25627,N_24877,N_24345);
and U25628 (N_25628,N_24895,N_25118);
nand U25629 (N_25629,N_24682,N_24792);
and U25630 (N_25630,N_24435,N_24408);
xor U25631 (N_25631,N_24313,N_25309);
nor U25632 (N_25632,N_24586,N_24973);
and U25633 (N_25633,N_25353,N_24307);
or U25634 (N_25634,N_25205,N_25460);
or U25635 (N_25635,N_25005,N_25172);
nor U25636 (N_25636,N_25445,N_24461);
nand U25637 (N_25637,N_25337,N_24256);
xor U25638 (N_25638,N_24494,N_25448);
nor U25639 (N_25639,N_25035,N_24866);
nand U25640 (N_25640,N_25265,N_24098);
and U25641 (N_25641,N_24157,N_24230);
xor U25642 (N_25642,N_24639,N_24457);
and U25643 (N_25643,N_24013,N_24569);
nor U25644 (N_25644,N_24083,N_24517);
xnor U25645 (N_25645,N_25365,N_24659);
or U25646 (N_25646,N_24580,N_24275);
nand U25647 (N_25647,N_25344,N_24136);
nor U25648 (N_25648,N_24585,N_24823);
nand U25649 (N_25649,N_24698,N_24316);
xnor U25650 (N_25650,N_24562,N_25440);
and U25651 (N_25651,N_24934,N_24153);
nand U25652 (N_25652,N_24487,N_25342);
xnor U25653 (N_25653,N_24264,N_25475);
nor U25654 (N_25654,N_25314,N_24912);
and U25655 (N_25655,N_24186,N_25116);
xnor U25656 (N_25656,N_24422,N_24654);
nor U25657 (N_25657,N_24265,N_24539);
xnor U25658 (N_25658,N_25415,N_24864);
or U25659 (N_25659,N_24530,N_24193);
nand U25660 (N_25660,N_24472,N_24201);
nor U25661 (N_25661,N_24647,N_25052);
or U25662 (N_25662,N_24795,N_25113);
nand U25663 (N_25663,N_24092,N_24183);
xor U25664 (N_25664,N_24424,N_24335);
nor U25665 (N_25665,N_24349,N_25032);
and U25666 (N_25666,N_25452,N_24582);
xor U25667 (N_25667,N_24773,N_25388);
and U25668 (N_25668,N_24851,N_24101);
and U25669 (N_25669,N_25435,N_24865);
and U25670 (N_25670,N_24522,N_24077);
nand U25671 (N_25671,N_24084,N_24688);
or U25672 (N_25672,N_24445,N_24600);
nor U25673 (N_25673,N_24134,N_24397);
or U25674 (N_25674,N_24712,N_24111);
nand U25675 (N_25675,N_24296,N_24320);
and U25676 (N_25676,N_24443,N_25311);
or U25677 (N_25677,N_24272,N_24991);
and U25678 (N_25678,N_24543,N_24635);
xnor U25679 (N_25679,N_24184,N_25450);
and U25680 (N_25680,N_24938,N_25466);
xnor U25681 (N_25681,N_25102,N_24886);
or U25682 (N_25682,N_24014,N_24298);
and U25683 (N_25683,N_24610,N_24525);
nor U25684 (N_25684,N_25130,N_24643);
and U25685 (N_25685,N_25140,N_24656);
nor U25686 (N_25686,N_24960,N_25385);
nand U25687 (N_25687,N_25334,N_24337);
nor U25688 (N_25688,N_24343,N_24399);
or U25689 (N_25689,N_24260,N_25283);
or U25690 (N_25690,N_25067,N_24675);
and U25691 (N_25691,N_25248,N_24133);
and U25692 (N_25692,N_24442,N_24125);
nor U25693 (N_25693,N_25196,N_25092);
xnor U25694 (N_25694,N_25389,N_24195);
nor U25695 (N_25695,N_25287,N_24791);
and U25696 (N_25696,N_25262,N_25437);
nor U25697 (N_25697,N_24318,N_24645);
or U25698 (N_25698,N_25480,N_24750);
nor U25699 (N_25699,N_24544,N_25461);
and U25700 (N_25700,N_25029,N_24008);
nor U25701 (N_25701,N_24510,N_25051);
xnor U25702 (N_25702,N_24038,N_24521);
or U25703 (N_25703,N_24637,N_24504);
nor U25704 (N_25704,N_25250,N_24541);
nor U25705 (N_25705,N_24784,N_25060);
nand U25706 (N_25706,N_24898,N_24616);
and U25707 (N_25707,N_24401,N_24489);
nor U25708 (N_25708,N_24797,N_24602);
nor U25709 (N_25709,N_24410,N_24211);
and U25710 (N_25710,N_24484,N_24909);
xnor U25711 (N_25711,N_24687,N_24943);
xor U25712 (N_25712,N_24788,N_25227);
and U25713 (N_25713,N_25259,N_24465);
xnor U25714 (N_25714,N_24601,N_24076);
and U25715 (N_25715,N_24344,N_25121);
xnor U25716 (N_25716,N_24807,N_24254);
or U25717 (N_25717,N_25125,N_24190);
nand U25718 (N_25718,N_24644,N_25015);
nor U25719 (N_25719,N_24966,N_24554);
nand U25720 (N_25720,N_24548,N_25063);
or U25721 (N_25721,N_24403,N_25247);
or U25722 (N_25722,N_24433,N_25163);
and U25723 (N_25723,N_25041,N_25095);
nor U25724 (N_25724,N_24365,N_25478);
nand U25725 (N_25725,N_24431,N_24853);
xnor U25726 (N_25726,N_25148,N_25368);
or U25727 (N_25727,N_24248,N_24292);
nand U25728 (N_25728,N_24836,N_24519);
nand U25729 (N_25729,N_24591,N_24595);
or U25730 (N_25730,N_24948,N_24763);
and U25731 (N_25731,N_24981,N_24317);
and U25732 (N_25732,N_25188,N_25394);
nor U25733 (N_25733,N_25016,N_25307);
nor U25734 (N_25734,N_25213,N_24518);
nor U25735 (N_25735,N_25494,N_24563);
or U25736 (N_25736,N_24032,N_25349);
xnor U25737 (N_25737,N_24226,N_24841);
xor U25738 (N_25738,N_25091,N_24994);
and U25739 (N_25739,N_24942,N_25362);
and U25740 (N_25740,N_24161,N_24035);
nor U25741 (N_25741,N_24920,N_24718);
and U25742 (N_25742,N_24587,N_24664);
nand U25743 (N_25743,N_25070,N_24513);
or U25744 (N_25744,N_24389,N_24202);
nor U25745 (N_25745,N_24947,N_24090);
xor U25746 (N_25746,N_25206,N_24052);
or U25747 (N_25747,N_25281,N_25499);
xor U25748 (N_25748,N_24801,N_24055);
or U25749 (N_25749,N_24158,N_24380);
nor U25750 (N_25750,N_24074,N_24289);
nor U25751 (N_25751,N_24110,N_25487);
and U25752 (N_25752,N_24143,N_24531);
xnor U25753 (N_25753,N_25151,N_24534);
nor U25754 (N_25754,N_25411,N_25431);
xor U25755 (N_25755,N_25434,N_24977);
or U25756 (N_25756,N_24280,N_24466);
nand U25757 (N_25757,N_24221,N_25175);
nand U25758 (N_25758,N_25239,N_24481);
nand U25759 (N_25759,N_24216,N_24810);
and U25760 (N_25760,N_24416,N_24141);
nand U25761 (N_25761,N_24705,N_25468);
nor U25762 (N_25762,N_24412,N_24419);
nand U25763 (N_25763,N_25038,N_25295);
nand U25764 (N_25764,N_24604,N_24612);
nor U25765 (N_25765,N_24219,N_25407);
nand U25766 (N_25766,N_25496,N_25360);
nor U25767 (N_25767,N_25033,N_24690);
xnor U25768 (N_25768,N_24414,N_25279);
xnor U25769 (N_25769,N_24714,N_24368);
and U25770 (N_25770,N_25133,N_24858);
nand U25771 (N_25771,N_25034,N_25275);
nor U25772 (N_25772,N_25336,N_24500);
or U25773 (N_25773,N_24295,N_24283);
xnor U25774 (N_25774,N_24132,N_24852);
and U25775 (N_25775,N_25216,N_24286);
nor U25776 (N_25776,N_25168,N_25317);
nand U25777 (N_25777,N_24578,N_25286);
and U25778 (N_25778,N_24993,N_24843);
or U25779 (N_25779,N_24135,N_25210);
and U25780 (N_25780,N_25218,N_25376);
and U25781 (N_25781,N_25026,N_25025);
and U25782 (N_25782,N_25000,N_25203);
xnor U25783 (N_25783,N_24482,N_24652);
nand U25784 (N_25784,N_25284,N_24067);
or U25785 (N_25785,N_25134,N_24557);
xnor U25786 (N_25786,N_25381,N_24123);
and U25787 (N_25787,N_24783,N_25018);
or U25788 (N_25788,N_24493,N_24062);
or U25789 (N_25789,N_24964,N_24925);
nand U25790 (N_25790,N_25078,N_25064);
nand U25791 (N_25791,N_24745,N_24180);
and U25792 (N_25792,N_24446,N_24998);
nor U25793 (N_25793,N_25442,N_24339);
and U25794 (N_25794,N_25331,N_24623);
nor U25795 (N_25795,N_24893,N_24238);
nor U25796 (N_25796,N_24294,N_25438);
and U25797 (N_25797,N_25080,N_24650);
nor U25798 (N_25798,N_24789,N_24034);
xnor U25799 (N_25799,N_25086,N_24485);
nor U25800 (N_25800,N_24139,N_24529);
xnor U25801 (N_25801,N_24820,N_24896);
nor U25802 (N_25802,N_24063,N_24561);
and U25803 (N_25803,N_24029,N_25042);
xor U25804 (N_25804,N_24672,N_24496);
or U25805 (N_25805,N_25387,N_25266);
and U25806 (N_25806,N_24660,N_24277);
and U25807 (N_25807,N_24808,N_24242);
nor U25808 (N_25808,N_24733,N_24802);
and U25809 (N_25809,N_24704,N_25028);
or U25810 (N_25810,N_24187,N_25361);
or U25811 (N_25811,N_24933,N_24764);
or U25812 (N_25812,N_25098,N_25129);
and U25813 (N_25813,N_24278,N_25249);
or U25814 (N_25814,N_25399,N_25303);
and U25815 (N_25815,N_25301,N_25426);
nor U25816 (N_25816,N_24369,N_24813);
nand U25817 (N_25817,N_24128,N_24894);
xor U25818 (N_25818,N_25100,N_24932);
or U25819 (N_25819,N_24108,N_24005);
xnor U25820 (N_25820,N_25031,N_24628);
and U25821 (N_25821,N_24636,N_25293);
nor U25822 (N_25822,N_25127,N_24734);
nor U25823 (N_25823,N_25439,N_24663);
or U25824 (N_25824,N_24250,N_25040);
nand U25825 (N_25825,N_24207,N_24208);
and U25826 (N_25826,N_24436,N_25477);
or U25827 (N_25827,N_25021,N_24825);
and U25828 (N_25828,N_24804,N_24581);
xor U25829 (N_25829,N_25483,N_25047);
and U25830 (N_25830,N_25327,N_24437);
and U25831 (N_25831,N_24961,N_24310);
xor U25832 (N_25832,N_25164,N_24887);
nand U25833 (N_25833,N_24729,N_24147);
nand U25834 (N_25834,N_24012,N_24086);
xor U25835 (N_25835,N_24879,N_25073);
and U25836 (N_25836,N_25222,N_24270);
xnor U25837 (N_25837,N_24568,N_25359);
and U25838 (N_25838,N_24775,N_25062);
nor U25839 (N_25839,N_25228,N_24194);
or U25840 (N_25840,N_25493,N_24081);
nor U25841 (N_25841,N_24429,N_24911);
and U25842 (N_25842,N_25370,N_24104);
or U25843 (N_25843,N_25152,N_24096);
or U25844 (N_25844,N_24378,N_24553);
or U25845 (N_25845,N_24646,N_24824);
nor U25846 (N_25846,N_25340,N_24990);
and U25847 (N_25847,N_25011,N_24405);
nor U25848 (N_25848,N_24838,N_24423);
and U25849 (N_25849,N_24781,N_24271);
and U25850 (N_25850,N_24701,N_25258);
xor U25851 (N_25851,N_24904,N_24379);
nor U25852 (N_25852,N_24821,N_24257);
and U25853 (N_25853,N_25003,N_24306);
nor U25854 (N_25854,N_24491,N_24253);
nand U25855 (N_25855,N_24418,N_24528);
xnor U25856 (N_25856,N_25300,N_24428);
nor U25857 (N_25857,N_24300,N_24988);
and U25858 (N_25858,N_24381,N_25479);
and U25859 (N_25859,N_24511,N_25104);
and U25860 (N_25860,N_24164,N_25079);
and U25861 (N_25861,N_25123,N_24840);
or U25862 (N_25862,N_25089,N_25162);
nor U25863 (N_25863,N_25305,N_24532);
xnor U25864 (N_25864,N_24178,N_25471);
xor U25865 (N_25865,N_25126,N_24527);
xor U25866 (N_25866,N_25106,N_24302);
nor U25867 (N_25867,N_25323,N_25298);
nor U25868 (N_25868,N_24550,N_24455);
xnor U25869 (N_25869,N_25111,N_24490);
nand U25870 (N_25870,N_24022,N_24899);
and U25871 (N_25871,N_25014,N_24346);
xnor U25872 (N_25872,N_24503,N_25357);
xnor U25873 (N_25873,N_25430,N_24631);
nand U25874 (N_25874,N_25418,N_25341);
nand U25875 (N_25875,N_24066,N_24269);
nand U25876 (N_25876,N_25190,N_24916);
nand U25877 (N_25877,N_25160,N_24373);
xor U25878 (N_25878,N_24793,N_24598);
nand U25879 (N_25879,N_24420,N_24276);
nor U25880 (N_25880,N_24930,N_24026);
nand U25881 (N_25881,N_24311,N_25383);
or U25882 (N_25882,N_24293,N_25061);
nand U25883 (N_25883,N_24707,N_24570);
or U25884 (N_25884,N_24069,N_24357);
and U25885 (N_25885,N_25225,N_25013);
or U25886 (N_25886,N_24622,N_24910);
and U25887 (N_25887,N_25161,N_24771);
nand U25888 (N_25888,N_25463,N_24721);
or U25889 (N_25889,N_24965,N_24176);
xor U25890 (N_25890,N_24393,N_24255);
nand U25891 (N_25891,N_25093,N_24430);
nand U25892 (N_25892,N_25312,N_25273);
xor U25893 (N_25893,N_24549,N_24606);
nor U25894 (N_25894,N_25456,N_24385);
xnor U25895 (N_25895,N_24592,N_24969);
nand U25896 (N_25896,N_24815,N_24363);
xor U25897 (N_25897,N_24177,N_25090);
xnor U25898 (N_25898,N_24777,N_25412);
nor U25899 (N_25899,N_25059,N_24359);
and U25900 (N_25900,N_24715,N_24599);
nor U25901 (N_25901,N_24448,N_24951);
nor U25902 (N_25902,N_24913,N_24374);
and U25903 (N_25903,N_24376,N_24693);
or U25904 (N_25904,N_24928,N_24002);
nor U25905 (N_25905,N_24935,N_25451);
xnor U25906 (N_25906,N_24325,N_24303);
nand U25907 (N_25907,N_24027,N_24679);
nor U25908 (N_25908,N_24057,N_24024);
and U25909 (N_25909,N_24859,N_25201);
xor U25910 (N_25910,N_25458,N_24170);
xor U25911 (N_25911,N_25083,N_24137);
and U25912 (N_25912,N_24236,N_24759);
xor U25913 (N_25913,N_24217,N_25417);
and U25914 (N_25914,N_24165,N_24985);
nor U25915 (N_25915,N_24720,N_25002);
xor U25916 (N_25916,N_24702,N_24787);
nand U25917 (N_25917,N_25269,N_24986);
or U25918 (N_25918,N_24968,N_24831);
or U25919 (N_25919,N_25413,N_24665);
xor U25920 (N_25920,N_25099,N_25069);
nor U25921 (N_25921,N_24741,N_24239);
xnor U25922 (N_25922,N_24618,N_24324);
or U25923 (N_25923,N_24970,N_24045);
xnor U25924 (N_25924,N_25158,N_24021);
nand U25925 (N_25925,N_25288,N_24790);
nor U25926 (N_25926,N_24923,N_24247);
xnor U25927 (N_25927,N_24869,N_24159);
xor U25928 (N_25928,N_24684,N_24772);
or U25929 (N_25929,N_24770,N_25108);
or U25930 (N_25930,N_25114,N_24651);
nand U25931 (N_25931,N_24148,N_24188);
nand U25932 (N_25932,N_24051,N_24742);
and U25933 (N_25933,N_25422,N_25304);
or U25934 (N_25934,N_24992,N_24962);
nand U25935 (N_25935,N_24728,N_24697);
nor U25936 (N_25936,N_24371,N_24471);
and U25937 (N_25937,N_25400,N_24361);
nor U25938 (N_25938,N_24655,N_24740);
or U25939 (N_25939,N_24614,N_24640);
nor U25940 (N_25940,N_25490,N_25195);
nand U25941 (N_25941,N_25217,N_24041);
and U25942 (N_25942,N_24453,N_24150);
and U25943 (N_25943,N_25351,N_24116);
or U25944 (N_25944,N_24850,N_25421);
and U25945 (N_25945,N_25358,N_24945);
xor U25946 (N_25946,N_25174,N_24044);
or U25947 (N_25947,N_24229,N_24304);
and U25948 (N_25948,N_24237,N_24244);
or U25949 (N_25949,N_24538,N_24873);
and U25950 (N_25950,N_24730,N_24641);
or U25951 (N_25951,N_24996,N_24819);
or U25952 (N_25952,N_25444,N_25377);
and U25953 (N_25953,N_25243,N_24151);
nand U25954 (N_25954,N_25176,N_24861);
nand U25955 (N_25955,N_25306,N_24856);
nand U25956 (N_25956,N_24737,N_25380);
nand U25957 (N_25957,N_24347,N_24117);
or U25958 (N_25958,N_24572,N_25443);
or U25959 (N_25959,N_25352,N_24072);
nand U25960 (N_25960,N_24958,N_24769);
nand U25961 (N_25961,N_24469,N_25354);
xor U25962 (N_25962,N_24145,N_25107);
nand U25963 (N_25963,N_24321,N_25419);
and U25964 (N_25964,N_24450,N_24036);
and U25965 (N_25965,N_24358,N_24071);
nor U25966 (N_25966,N_24800,N_24018);
nand U25967 (N_25967,N_24508,N_24322);
nor U25968 (N_25968,N_24579,N_24842);
nand U25969 (N_25969,N_24196,N_24761);
and U25970 (N_25970,N_24624,N_24782);
nor U25971 (N_25971,N_24863,N_24109);
and U25972 (N_25972,N_24227,N_25495);
nand U25973 (N_25973,N_25267,N_25020);
nor U25974 (N_25974,N_24648,N_24523);
or U25975 (N_25975,N_24514,N_24070);
xor U25976 (N_25976,N_24011,N_24833);
nand U25977 (N_25977,N_24683,N_24537);
nand U25978 (N_25978,N_24924,N_24681);
xnor U25979 (N_25979,N_24736,N_25101);
and U25980 (N_25980,N_24710,N_25330);
and U25981 (N_25981,N_24972,N_24099);
nand U25982 (N_25982,N_24042,N_24284);
and U25983 (N_25983,N_24922,N_24355);
or U25984 (N_25984,N_24520,N_24754);
nor U25985 (N_25985,N_25143,N_24025);
nand U25986 (N_25986,N_24223,N_25280);
xnor U25987 (N_25987,N_24174,N_24613);
nand U25988 (N_25988,N_25409,N_24512);
nand U25989 (N_25989,N_25153,N_24168);
and U25990 (N_25990,N_24902,N_24583);
or U25991 (N_25991,N_24847,N_24413);
nand U25992 (N_25992,N_25462,N_24871);
xnor U25993 (N_25993,N_24828,N_24082);
nor U25994 (N_25994,N_24282,N_25221);
or U25995 (N_25995,N_25207,N_24103);
xor U25996 (N_25996,N_24274,N_24906);
or U25997 (N_25997,N_24708,N_25112);
and U25998 (N_25998,N_25256,N_24392);
nor U25999 (N_25999,N_25171,N_24462);
nand U26000 (N_26000,N_24502,N_24692);
nor U26001 (N_26001,N_25369,N_24049);
nor U26002 (N_26002,N_24989,N_24524);
and U26003 (N_26003,N_24259,N_24780);
nor U26004 (N_26004,N_25482,N_24950);
xnor U26005 (N_26005,N_24867,N_24334);
nor U26006 (N_26006,N_25374,N_24979);
or U26007 (N_26007,N_24882,N_24905);
nor U26008 (N_26008,N_24189,N_24803);
or U26009 (N_26009,N_25166,N_24497);
xnor U26010 (N_26010,N_24279,N_24079);
nand U26011 (N_26011,N_24987,N_24603);
or U26012 (N_26012,N_24739,N_24214);
or U26013 (N_26013,N_24477,N_25366);
nand U26014 (N_26014,N_25497,N_24213);
and U26015 (N_26015,N_24669,N_24868);
nand U26016 (N_26016,N_25173,N_25325);
or U26017 (N_26017,N_25350,N_24827);
nand U26018 (N_26018,N_24609,N_25194);
nor U26019 (N_26019,N_24068,N_25277);
nor U26020 (N_26020,N_24362,N_25183);
and U26021 (N_26021,N_24329,N_25232);
nor U26022 (N_26022,N_24978,N_24390);
or U26023 (N_26023,N_24404,N_25459);
nor U26024 (N_26024,N_24372,N_24767);
nand U26025 (N_26025,N_24262,N_25428);
or U26026 (N_26026,N_24458,N_25274);
and U26027 (N_26027,N_25469,N_25484);
nor U26028 (N_26028,N_25289,N_24713);
xor U26029 (N_26029,N_24590,N_25492);
or U26030 (N_26030,N_25142,N_25328);
or U26031 (N_26031,N_24724,N_24953);
xnor U26032 (N_26032,N_25436,N_24367);
nand U26033 (N_26033,N_24326,N_25124);
nor U26034 (N_26034,N_24884,N_24768);
xor U26035 (N_26035,N_25030,N_24387);
nor U26036 (N_26036,N_24095,N_24386);
and U26037 (N_26037,N_24642,N_24917);
xnor U26038 (N_26038,N_25315,N_25393);
and U26039 (N_26039,N_25023,N_24501);
or U26040 (N_26040,N_24837,N_25074);
or U26041 (N_26041,N_24760,N_24627);
xnor U26042 (N_26042,N_24776,N_24939);
and U26043 (N_26043,N_25245,N_24829);
and U26044 (N_26044,N_24006,N_25199);
and U26045 (N_26045,N_24222,N_25202);
nor U26046 (N_26046,N_25022,N_24849);
nor U26047 (N_26047,N_24309,N_25375);
nand U26048 (N_26048,N_24114,N_24009);
nor U26049 (N_26049,N_25044,N_25132);
or U26050 (N_26050,N_25486,N_25416);
nor U26051 (N_26051,N_24822,N_24653);
nand U26052 (N_26052,N_25345,N_25424);
xnor U26053 (N_26053,N_24897,N_24396);
nand U26054 (N_26054,N_25177,N_24426);
and U26055 (N_26055,N_25464,N_24224);
or U26056 (N_26056,N_24475,N_24567);
nor U26057 (N_26057,N_24441,N_24555);
and U26058 (N_26058,N_25036,N_24699);
or U26059 (N_26059,N_24983,N_25170);
xnor U26060 (N_26060,N_25390,N_24731);
xor U26061 (N_26061,N_25198,N_24785);
and U26062 (N_26062,N_24559,N_24593);
nor U26063 (N_26063,N_25180,N_24596);
and U26064 (N_26064,N_24360,N_24199);
nand U26065 (N_26065,N_25076,N_24854);
nand U26066 (N_26066,N_24725,N_25082);
nand U26067 (N_26067,N_25240,N_24552);
and U26068 (N_26068,N_24848,N_24078);
xor U26069 (N_26069,N_24291,N_25008);
nor U26070 (N_26070,N_24509,N_24406);
nand U26071 (N_26071,N_24941,N_24407);
and U26072 (N_26072,N_25117,N_25473);
nor U26073 (N_26073,N_24617,N_24102);
or U26074 (N_26074,N_24862,N_25087);
and U26075 (N_26075,N_24031,N_24937);
nor U26076 (N_26076,N_25402,N_25410);
nand U26077 (N_26077,N_25004,N_24267);
xnor U26078 (N_26078,N_24658,N_25081);
or U26079 (N_26079,N_24625,N_25056);
xor U26080 (N_26080,N_24778,N_24232);
nand U26081 (N_26081,N_25253,N_24434);
nand U26082 (N_26082,N_25255,N_24774);
nand U26083 (N_26083,N_24415,N_24241);
xor U26084 (N_26084,N_25316,N_25237);
nand U26085 (N_26085,N_25367,N_25379);
nand U26086 (N_26086,N_25200,N_25472);
nand U26087 (N_26087,N_24402,N_25272);
xor U26088 (N_26088,N_24839,N_24674);
xnor U26089 (N_26089,N_24997,N_24676);
nand U26090 (N_26090,N_24999,N_24826);
xor U26091 (N_26091,N_25260,N_25068);
and U26092 (N_26092,N_25398,N_25149);
xnor U26093 (N_26093,N_24251,N_24881);
nand U26094 (N_26094,N_24799,N_24039);
or U26095 (N_26095,N_24931,N_24615);
xor U26096 (N_26096,N_24976,N_25291);
nor U26097 (N_26097,N_24691,N_25433);
xnor U26098 (N_26098,N_24556,N_25135);
and U26099 (N_26099,N_25096,N_25085);
nand U26100 (N_26100,N_24268,N_25467);
xor U26101 (N_26101,N_24929,N_24700);
nor U26102 (N_26102,N_24015,N_25179);
or U26103 (N_26103,N_24384,N_25276);
and U26104 (N_26104,N_24765,N_24696);
and U26105 (N_26105,N_24498,N_25449);
nor U26106 (N_26106,N_24375,N_24444);
xnor U26107 (N_26107,N_24726,N_25115);
nand U26108 (N_26108,N_24105,N_25208);
and U26109 (N_26109,N_24483,N_24124);
and U26110 (N_26110,N_25146,N_24752);
or U26111 (N_26111,N_25204,N_24185);
xor U26112 (N_26112,N_25318,N_25186);
nor U26113 (N_26113,N_24588,N_24233);
xnor U26114 (N_26114,N_25055,N_25414);
nor U26115 (N_26115,N_25212,N_25491);
nand U26116 (N_26116,N_24488,N_24830);
nand U26117 (N_26117,N_24087,N_25141);
or U26118 (N_26118,N_24794,N_24016);
xor U26119 (N_26119,N_24980,N_24001);
xor U26120 (N_26120,N_24452,N_24649);
or U26121 (N_26121,N_25498,N_25075);
or U26122 (N_26122,N_24940,N_24516);
nor U26123 (N_26123,N_24323,N_25077);
nor U26124 (N_26124,N_24175,N_25447);
nand U26125 (N_26125,N_24565,N_24315);
nor U26126 (N_26126,N_24855,N_24845);
nor U26127 (N_26127,N_25191,N_24205);
nand U26128 (N_26128,N_24908,N_24017);
nand U26129 (N_26129,N_24266,N_25457);
and U26130 (N_26130,N_24671,N_25294);
nor U26131 (N_26131,N_25363,N_24959);
or U26132 (N_26132,N_25310,N_24007);
or U26133 (N_26133,N_24936,N_25282);
nor U26134 (N_26134,N_24874,N_24245);
or U26135 (N_26135,N_24330,N_25169);
nand U26136 (N_26136,N_24100,N_24903);
xnor U26137 (N_26137,N_25382,N_24955);
nand U26138 (N_26138,N_25236,N_25488);
xnor U26139 (N_26139,N_24872,N_24900);
and U26140 (N_26140,N_25432,N_24479);
xor U26141 (N_26141,N_24818,N_24844);
nand U26142 (N_26142,N_24364,N_24817);
nand U26143 (N_26143,N_24575,N_24093);
nand U26144 (N_26144,N_24480,N_24685);
or U26145 (N_26145,N_25057,N_24907);
or U26146 (N_26146,N_24366,N_25313);
xor U26147 (N_26147,N_25425,N_25268);
xnor U26148 (N_26148,N_24661,N_25138);
xor U26149 (N_26149,N_25423,N_24144);
xor U26150 (N_26150,N_25302,N_24421);
xnor U26151 (N_26151,N_24756,N_24198);
nor U26152 (N_26152,N_24526,N_25364);
nand U26153 (N_26153,N_24171,N_24719);
and U26154 (N_26154,N_25290,N_24878);
nor U26155 (N_26155,N_24231,N_25420);
nand U26156 (N_26156,N_24037,N_25372);
nor U26157 (N_26157,N_24348,N_24129);
nor U26158 (N_26158,N_24812,N_24299);
xor U26159 (N_26159,N_24354,N_25455);
nand U26160 (N_26160,N_24717,N_25271);
and U26161 (N_26161,N_24880,N_25371);
and U26162 (N_26162,N_24667,N_25167);
xnor U26163 (N_26163,N_24753,N_24890);
nor U26164 (N_26164,N_25007,N_25292);
and U26165 (N_26165,N_25396,N_24558);
xnor U26166 (N_26166,N_24273,N_24439);
or U26167 (N_26167,N_25264,N_24182);
nor U26168 (N_26168,N_25234,N_24727);
nand U26169 (N_26169,N_24173,N_24576);
xnor U26170 (N_26170,N_24338,N_24589);
and U26171 (N_26171,N_25427,N_25233);
or U26172 (N_26172,N_25339,N_24711);
nor U26173 (N_26173,N_24957,N_24225);
or U26174 (N_26174,N_24626,N_24757);
and U26175 (N_26175,N_24499,N_24779);
and U26176 (N_26176,N_25165,N_24695);
nor U26177 (N_26177,N_25181,N_24703);
nand U26178 (N_26178,N_25197,N_25103);
nand U26179 (N_26179,N_25406,N_25071);
xor U26180 (N_26180,N_24995,N_24212);
and U26181 (N_26181,N_24927,N_24680);
nand U26182 (N_26182,N_24046,N_25019);
or U26183 (N_26183,N_24846,N_25229);
or U26184 (N_26184,N_24875,N_25144);
xnor U26185 (N_26185,N_24043,N_24694);
and U26186 (N_26186,N_24805,N_24486);
nand U26187 (N_26187,N_24634,N_25489);
or U26188 (N_26188,N_25054,N_25214);
nor U26189 (N_26189,N_25043,N_25474);
and U26190 (N_26190,N_25039,N_24030);
nor U26191 (N_26191,N_25235,N_24053);
nand U26192 (N_26192,N_24218,N_24048);
nand U26193 (N_26193,N_25159,N_24876);
nand U26194 (N_26194,N_25391,N_24287);
nor U26195 (N_26195,N_24566,N_24192);
or U26196 (N_26196,N_24156,N_24167);
xnor U26197 (N_26197,N_24064,N_24127);
and U26198 (N_26198,N_24447,N_25322);
nor U26199 (N_26199,N_25131,N_24228);
and U26200 (N_26200,N_24686,N_25481);
nand U26201 (N_26201,N_25155,N_24122);
nor U26202 (N_26202,N_24638,N_24584);
nand U26203 (N_26203,N_25319,N_24033);
or U26204 (N_26204,N_25238,N_25373);
and U26205 (N_26205,N_24464,N_24336);
and U26206 (N_26206,N_24409,N_25105);
nand U26207 (N_26207,N_24459,N_24914);
xnor U26208 (N_26208,N_24391,N_24870);
nor U26209 (N_26209,N_24540,N_24678);
or U26210 (N_26210,N_24747,N_24411);
and U26211 (N_26211,N_25378,N_25088);
xnor U26212 (N_26212,N_24545,N_24047);
or U26213 (N_26213,N_24297,N_24332);
nor U26214 (N_26214,N_24235,N_24085);
nor U26215 (N_26215,N_25335,N_24984);
xor U26216 (N_26216,N_24723,N_24597);
xor U26217 (N_26217,N_24203,N_24206);
or U26218 (N_26218,N_24633,N_24758);
nor U26219 (N_26219,N_25230,N_24535);
and U26220 (N_26220,N_25446,N_24835);
or U26221 (N_26221,N_25145,N_25136);
and U26222 (N_26222,N_24515,N_24832);
nand U26223 (N_26223,N_24506,N_24809);
nor U26224 (N_26224,N_25109,N_24327);
and U26225 (N_26225,N_24388,N_25254);
nor U26226 (N_26226,N_25348,N_24215);
and U26227 (N_26227,N_24449,N_25184);
xnor U26228 (N_26228,N_24536,N_24574);
xnor U26229 (N_26229,N_25441,N_24261);
and U26230 (N_26230,N_24505,N_24478);
xor U26231 (N_26231,N_24328,N_25343);
nand U26232 (N_26232,N_24097,N_24451);
nand U26233 (N_26233,N_24152,N_24921);
xor U26234 (N_26234,N_24023,N_25397);
or U26235 (N_26235,N_24091,N_24370);
xor U26236 (N_26236,N_24467,N_25046);
nand U26237 (N_26237,N_25261,N_24751);
nor U26238 (N_26238,N_24605,N_24331);
and U26239 (N_26239,N_24673,N_25297);
nor U26240 (N_26240,N_24796,N_24901);
xor U26241 (N_26241,N_24560,N_24312);
nand U26242 (N_26242,N_25296,N_25084);
xnor U26243 (N_26243,N_24546,N_25050);
xnor U26244 (N_26244,N_25403,N_24154);
xnor U26245 (N_26245,N_25332,N_24892);
and U26246 (N_26246,N_24281,N_24258);
nor U26247 (N_26247,N_24308,N_24476);
nand U26248 (N_26248,N_24019,N_25401);
or U26249 (N_26249,N_25065,N_24564);
and U26250 (N_26250,N_25323,N_25388);
nand U26251 (N_26251,N_24471,N_25321);
xor U26252 (N_26252,N_24560,N_24205);
nor U26253 (N_26253,N_24438,N_24870);
nor U26254 (N_26254,N_25218,N_25459);
and U26255 (N_26255,N_24342,N_25437);
and U26256 (N_26256,N_24246,N_24676);
nand U26257 (N_26257,N_24187,N_24806);
or U26258 (N_26258,N_24011,N_25012);
or U26259 (N_26259,N_25281,N_24677);
or U26260 (N_26260,N_24266,N_25192);
xnor U26261 (N_26261,N_24216,N_24283);
xor U26262 (N_26262,N_24643,N_25282);
xnor U26263 (N_26263,N_24268,N_24990);
or U26264 (N_26264,N_24595,N_24677);
nor U26265 (N_26265,N_25031,N_25398);
and U26266 (N_26266,N_24348,N_24976);
xor U26267 (N_26267,N_24313,N_24443);
nand U26268 (N_26268,N_25094,N_25009);
xor U26269 (N_26269,N_24104,N_24228);
or U26270 (N_26270,N_24914,N_24880);
nand U26271 (N_26271,N_24287,N_24282);
or U26272 (N_26272,N_24387,N_24514);
xor U26273 (N_26273,N_25002,N_24462);
xor U26274 (N_26274,N_24016,N_24871);
and U26275 (N_26275,N_25498,N_24348);
xor U26276 (N_26276,N_25340,N_24641);
and U26277 (N_26277,N_24376,N_24995);
nor U26278 (N_26278,N_24068,N_24566);
nand U26279 (N_26279,N_24380,N_24024);
nand U26280 (N_26280,N_24002,N_24622);
and U26281 (N_26281,N_24904,N_25277);
xor U26282 (N_26282,N_24347,N_25496);
or U26283 (N_26283,N_24812,N_24690);
xor U26284 (N_26284,N_24975,N_24467);
xor U26285 (N_26285,N_24700,N_24216);
and U26286 (N_26286,N_25220,N_25280);
nor U26287 (N_26287,N_24895,N_24862);
and U26288 (N_26288,N_25135,N_24104);
nand U26289 (N_26289,N_24689,N_24385);
or U26290 (N_26290,N_25495,N_24615);
xor U26291 (N_26291,N_24731,N_24908);
or U26292 (N_26292,N_24253,N_24383);
nor U26293 (N_26293,N_24059,N_24809);
nor U26294 (N_26294,N_24232,N_24448);
nand U26295 (N_26295,N_25118,N_24945);
and U26296 (N_26296,N_24056,N_24319);
xnor U26297 (N_26297,N_25336,N_24665);
nand U26298 (N_26298,N_24495,N_24457);
and U26299 (N_26299,N_24751,N_24563);
nand U26300 (N_26300,N_25127,N_25245);
and U26301 (N_26301,N_24826,N_25335);
and U26302 (N_26302,N_25119,N_24027);
nand U26303 (N_26303,N_24895,N_25245);
nand U26304 (N_26304,N_24745,N_24370);
and U26305 (N_26305,N_24872,N_24127);
nor U26306 (N_26306,N_24026,N_24954);
xor U26307 (N_26307,N_24684,N_25309);
nor U26308 (N_26308,N_24598,N_25093);
nand U26309 (N_26309,N_25122,N_24458);
nand U26310 (N_26310,N_24030,N_24568);
nor U26311 (N_26311,N_25349,N_24253);
and U26312 (N_26312,N_25405,N_25445);
and U26313 (N_26313,N_25392,N_24475);
nor U26314 (N_26314,N_25469,N_24943);
and U26315 (N_26315,N_24307,N_24469);
xor U26316 (N_26316,N_25073,N_25145);
xor U26317 (N_26317,N_24533,N_25458);
nor U26318 (N_26318,N_24039,N_24244);
xor U26319 (N_26319,N_24405,N_24388);
and U26320 (N_26320,N_25246,N_24677);
or U26321 (N_26321,N_24255,N_25170);
and U26322 (N_26322,N_24908,N_24497);
and U26323 (N_26323,N_25134,N_24009);
or U26324 (N_26324,N_25327,N_24172);
and U26325 (N_26325,N_25184,N_25195);
nor U26326 (N_26326,N_24413,N_24006);
nand U26327 (N_26327,N_24968,N_24687);
and U26328 (N_26328,N_24566,N_25145);
xnor U26329 (N_26329,N_24528,N_25117);
nor U26330 (N_26330,N_25011,N_25237);
and U26331 (N_26331,N_25022,N_24981);
nand U26332 (N_26332,N_24668,N_24572);
nand U26333 (N_26333,N_24803,N_24588);
nor U26334 (N_26334,N_24155,N_25217);
nor U26335 (N_26335,N_24069,N_25346);
and U26336 (N_26336,N_25313,N_25185);
and U26337 (N_26337,N_24188,N_24286);
and U26338 (N_26338,N_24478,N_25171);
or U26339 (N_26339,N_24469,N_25189);
and U26340 (N_26340,N_24900,N_24597);
and U26341 (N_26341,N_24632,N_24871);
and U26342 (N_26342,N_25288,N_24229);
nand U26343 (N_26343,N_24102,N_24730);
nand U26344 (N_26344,N_24247,N_24741);
nor U26345 (N_26345,N_24784,N_25326);
or U26346 (N_26346,N_24121,N_24137);
nor U26347 (N_26347,N_24024,N_24361);
nor U26348 (N_26348,N_24834,N_24471);
and U26349 (N_26349,N_24351,N_25147);
xnor U26350 (N_26350,N_24734,N_24953);
nor U26351 (N_26351,N_24243,N_24087);
nand U26352 (N_26352,N_24195,N_24409);
and U26353 (N_26353,N_24414,N_25214);
or U26354 (N_26354,N_24450,N_24528);
or U26355 (N_26355,N_24568,N_24831);
and U26356 (N_26356,N_25129,N_25421);
or U26357 (N_26357,N_25306,N_24055);
nand U26358 (N_26358,N_24525,N_25346);
xnor U26359 (N_26359,N_25468,N_24984);
xor U26360 (N_26360,N_24641,N_25264);
or U26361 (N_26361,N_24135,N_25362);
or U26362 (N_26362,N_24302,N_24861);
and U26363 (N_26363,N_24945,N_25029);
nor U26364 (N_26364,N_24999,N_24354);
and U26365 (N_26365,N_24950,N_25178);
xnor U26366 (N_26366,N_24606,N_24274);
or U26367 (N_26367,N_25306,N_24059);
or U26368 (N_26368,N_24397,N_24010);
or U26369 (N_26369,N_24491,N_24479);
or U26370 (N_26370,N_25459,N_24165);
xnor U26371 (N_26371,N_24602,N_24579);
and U26372 (N_26372,N_24658,N_24639);
or U26373 (N_26373,N_24984,N_24721);
or U26374 (N_26374,N_25093,N_25282);
xnor U26375 (N_26375,N_24023,N_24693);
nand U26376 (N_26376,N_24886,N_24283);
nor U26377 (N_26377,N_24942,N_24546);
nor U26378 (N_26378,N_25448,N_25238);
nand U26379 (N_26379,N_24288,N_25333);
xnor U26380 (N_26380,N_25109,N_25265);
nand U26381 (N_26381,N_24229,N_24757);
nand U26382 (N_26382,N_25393,N_24045);
nor U26383 (N_26383,N_24079,N_25388);
xnor U26384 (N_26384,N_24101,N_24015);
nor U26385 (N_26385,N_25474,N_24314);
or U26386 (N_26386,N_24052,N_25492);
and U26387 (N_26387,N_24644,N_24166);
or U26388 (N_26388,N_24882,N_24782);
nor U26389 (N_26389,N_24160,N_25094);
and U26390 (N_26390,N_24142,N_24405);
and U26391 (N_26391,N_24895,N_24247);
xnor U26392 (N_26392,N_24616,N_25168);
and U26393 (N_26393,N_24132,N_24407);
nor U26394 (N_26394,N_25227,N_24271);
and U26395 (N_26395,N_25184,N_25412);
and U26396 (N_26396,N_25082,N_24869);
nand U26397 (N_26397,N_24486,N_24099);
or U26398 (N_26398,N_24405,N_24133);
or U26399 (N_26399,N_24058,N_24394);
xor U26400 (N_26400,N_24117,N_24959);
or U26401 (N_26401,N_25253,N_24741);
xor U26402 (N_26402,N_25348,N_24420);
xnor U26403 (N_26403,N_24107,N_25484);
xor U26404 (N_26404,N_25458,N_25025);
or U26405 (N_26405,N_24665,N_24336);
nand U26406 (N_26406,N_25072,N_25013);
or U26407 (N_26407,N_25437,N_24405);
nor U26408 (N_26408,N_24829,N_24064);
and U26409 (N_26409,N_25055,N_24900);
nor U26410 (N_26410,N_24156,N_24432);
nand U26411 (N_26411,N_25297,N_25217);
and U26412 (N_26412,N_25461,N_24339);
xor U26413 (N_26413,N_24016,N_24405);
and U26414 (N_26414,N_24555,N_24851);
nand U26415 (N_26415,N_24268,N_24839);
and U26416 (N_26416,N_24050,N_25283);
nor U26417 (N_26417,N_24689,N_25227);
nand U26418 (N_26418,N_24063,N_24400);
xor U26419 (N_26419,N_24758,N_24183);
nand U26420 (N_26420,N_25424,N_24791);
or U26421 (N_26421,N_24872,N_24504);
nand U26422 (N_26422,N_25399,N_24234);
and U26423 (N_26423,N_25047,N_25374);
nor U26424 (N_26424,N_24660,N_24866);
xor U26425 (N_26425,N_25316,N_24644);
xnor U26426 (N_26426,N_24775,N_25210);
nor U26427 (N_26427,N_24701,N_24228);
or U26428 (N_26428,N_24190,N_24450);
and U26429 (N_26429,N_25123,N_25417);
or U26430 (N_26430,N_24594,N_25052);
or U26431 (N_26431,N_24687,N_24173);
xor U26432 (N_26432,N_25038,N_24406);
and U26433 (N_26433,N_25267,N_25296);
and U26434 (N_26434,N_24394,N_24448);
nor U26435 (N_26435,N_25346,N_25489);
and U26436 (N_26436,N_24673,N_25007);
or U26437 (N_26437,N_24720,N_24588);
and U26438 (N_26438,N_24997,N_25329);
and U26439 (N_26439,N_25029,N_24924);
nor U26440 (N_26440,N_25053,N_25495);
xnor U26441 (N_26441,N_25009,N_24904);
nand U26442 (N_26442,N_25326,N_25358);
nor U26443 (N_26443,N_24710,N_24364);
nand U26444 (N_26444,N_24639,N_24055);
xor U26445 (N_26445,N_25077,N_24569);
nand U26446 (N_26446,N_25275,N_24738);
or U26447 (N_26447,N_25484,N_24388);
or U26448 (N_26448,N_24938,N_25205);
nor U26449 (N_26449,N_24525,N_24714);
and U26450 (N_26450,N_24286,N_24528);
and U26451 (N_26451,N_24121,N_25105);
nor U26452 (N_26452,N_25237,N_24039);
xnor U26453 (N_26453,N_24728,N_24529);
nor U26454 (N_26454,N_25122,N_24762);
nor U26455 (N_26455,N_24049,N_25061);
nor U26456 (N_26456,N_24076,N_25166);
nand U26457 (N_26457,N_25083,N_24331);
xnor U26458 (N_26458,N_24963,N_25390);
xnor U26459 (N_26459,N_24338,N_24430);
nor U26460 (N_26460,N_24172,N_25111);
nor U26461 (N_26461,N_25347,N_24411);
xor U26462 (N_26462,N_25432,N_24939);
nand U26463 (N_26463,N_25156,N_24868);
or U26464 (N_26464,N_25171,N_24751);
and U26465 (N_26465,N_24443,N_24898);
nor U26466 (N_26466,N_25431,N_25360);
xor U26467 (N_26467,N_24014,N_24490);
xnor U26468 (N_26468,N_24074,N_24864);
xnor U26469 (N_26469,N_24201,N_25123);
and U26470 (N_26470,N_24089,N_24796);
nor U26471 (N_26471,N_24115,N_24370);
nor U26472 (N_26472,N_25128,N_25290);
and U26473 (N_26473,N_24832,N_25266);
and U26474 (N_26474,N_24218,N_25056);
xor U26475 (N_26475,N_24863,N_25280);
or U26476 (N_26476,N_24917,N_24935);
and U26477 (N_26477,N_24507,N_24840);
nor U26478 (N_26478,N_25384,N_24614);
and U26479 (N_26479,N_25480,N_24601);
and U26480 (N_26480,N_25280,N_25285);
and U26481 (N_26481,N_24424,N_25488);
nor U26482 (N_26482,N_25323,N_25127);
or U26483 (N_26483,N_24140,N_25441);
nor U26484 (N_26484,N_25019,N_25048);
or U26485 (N_26485,N_24232,N_24858);
nand U26486 (N_26486,N_25482,N_25029);
nor U26487 (N_26487,N_24182,N_24287);
or U26488 (N_26488,N_24382,N_25178);
or U26489 (N_26489,N_25378,N_25189);
or U26490 (N_26490,N_24391,N_24904);
or U26491 (N_26491,N_24598,N_24010);
and U26492 (N_26492,N_24375,N_24957);
nand U26493 (N_26493,N_25371,N_24727);
xnor U26494 (N_26494,N_24466,N_25093);
nand U26495 (N_26495,N_24266,N_24892);
nor U26496 (N_26496,N_25170,N_24038);
and U26497 (N_26497,N_25217,N_25444);
nor U26498 (N_26498,N_24557,N_24685);
nand U26499 (N_26499,N_25166,N_24301);
or U26500 (N_26500,N_25249,N_25006);
or U26501 (N_26501,N_25186,N_24245);
nor U26502 (N_26502,N_25247,N_24604);
or U26503 (N_26503,N_25078,N_24255);
xnor U26504 (N_26504,N_24601,N_24979);
nand U26505 (N_26505,N_25043,N_24453);
or U26506 (N_26506,N_24296,N_24099);
nor U26507 (N_26507,N_24553,N_24087);
nand U26508 (N_26508,N_25458,N_24224);
nand U26509 (N_26509,N_24620,N_25151);
nand U26510 (N_26510,N_24994,N_24526);
and U26511 (N_26511,N_24207,N_25415);
nand U26512 (N_26512,N_24371,N_25052);
and U26513 (N_26513,N_24480,N_24430);
nand U26514 (N_26514,N_24601,N_24834);
nand U26515 (N_26515,N_24442,N_25002);
xnor U26516 (N_26516,N_25057,N_25154);
xor U26517 (N_26517,N_24159,N_24311);
nand U26518 (N_26518,N_25109,N_25293);
nand U26519 (N_26519,N_25278,N_24898);
and U26520 (N_26520,N_25176,N_24155);
nand U26521 (N_26521,N_24033,N_25453);
or U26522 (N_26522,N_24629,N_24521);
and U26523 (N_26523,N_24109,N_24610);
xnor U26524 (N_26524,N_25431,N_25495);
nand U26525 (N_26525,N_24217,N_24429);
nor U26526 (N_26526,N_25420,N_25336);
nand U26527 (N_26527,N_24832,N_24024);
nor U26528 (N_26528,N_25483,N_25234);
xor U26529 (N_26529,N_24157,N_24194);
nor U26530 (N_26530,N_24575,N_24803);
nor U26531 (N_26531,N_24174,N_25364);
nand U26532 (N_26532,N_24570,N_24777);
nand U26533 (N_26533,N_24774,N_24086);
nor U26534 (N_26534,N_24527,N_25136);
nor U26535 (N_26535,N_25174,N_25307);
xnor U26536 (N_26536,N_24699,N_24486);
nand U26537 (N_26537,N_24176,N_24216);
or U26538 (N_26538,N_24426,N_24952);
and U26539 (N_26539,N_24835,N_24454);
and U26540 (N_26540,N_24137,N_24312);
and U26541 (N_26541,N_24654,N_25098);
xnor U26542 (N_26542,N_25164,N_24526);
nor U26543 (N_26543,N_24445,N_25333);
nor U26544 (N_26544,N_25262,N_24523);
and U26545 (N_26545,N_24763,N_25080);
xor U26546 (N_26546,N_25131,N_25156);
nand U26547 (N_26547,N_24986,N_25474);
xor U26548 (N_26548,N_25212,N_24233);
and U26549 (N_26549,N_24355,N_24019);
or U26550 (N_26550,N_24615,N_24992);
and U26551 (N_26551,N_24227,N_24052);
nand U26552 (N_26552,N_24844,N_24372);
xor U26553 (N_26553,N_24158,N_24009);
or U26554 (N_26554,N_24831,N_24154);
or U26555 (N_26555,N_24341,N_24129);
nor U26556 (N_26556,N_24962,N_24426);
and U26557 (N_26557,N_24689,N_24918);
xnor U26558 (N_26558,N_24654,N_25411);
nor U26559 (N_26559,N_25084,N_24535);
or U26560 (N_26560,N_24368,N_24506);
nor U26561 (N_26561,N_25422,N_24998);
nand U26562 (N_26562,N_25405,N_25098);
nor U26563 (N_26563,N_25109,N_24465);
or U26564 (N_26564,N_24255,N_24207);
nor U26565 (N_26565,N_25495,N_25369);
xnor U26566 (N_26566,N_25163,N_24198);
nor U26567 (N_26567,N_24552,N_25038);
or U26568 (N_26568,N_24592,N_24172);
and U26569 (N_26569,N_24199,N_24986);
and U26570 (N_26570,N_24248,N_24153);
or U26571 (N_26571,N_25310,N_24612);
nor U26572 (N_26572,N_24979,N_24820);
xor U26573 (N_26573,N_25477,N_24375);
nor U26574 (N_26574,N_25019,N_24912);
nor U26575 (N_26575,N_24989,N_24378);
and U26576 (N_26576,N_24235,N_25291);
xnor U26577 (N_26577,N_24043,N_25250);
xor U26578 (N_26578,N_25145,N_25384);
nor U26579 (N_26579,N_24378,N_24289);
and U26580 (N_26580,N_25287,N_24381);
nand U26581 (N_26581,N_24068,N_24176);
nor U26582 (N_26582,N_25256,N_24724);
nand U26583 (N_26583,N_25005,N_24818);
and U26584 (N_26584,N_24295,N_24452);
nand U26585 (N_26585,N_24953,N_24687);
or U26586 (N_26586,N_25216,N_24315);
nor U26587 (N_26587,N_24113,N_25039);
nand U26588 (N_26588,N_24520,N_25445);
nand U26589 (N_26589,N_25394,N_24742);
xnor U26590 (N_26590,N_24467,N_25409);
or U26591 (N_26591,N_24795,N_24655);
xor U26592 (N_26592,N_24213,N_24929);
or U26593 (N_26593,N_24252,N_25161);
nor U26594 (N_26594,N_25260,N_24645);
or U26595 (N_26595,N_24909,N_24750);
nor U26596 (N_26596,N_24663,N_24922);
xor U26597 (N_26597,N_25109,N_24813);
or U26598 (N_26598,N_24004,N_24490);
xnor U26599 (N_26599,N_24931,N_25096);
nor U26600 (N_26600,N_24081,N_25223);
xnor U26601 (N_26601,N_24145,N_25020);
xor U26602 (N_26602,N_24215,N_25037);
nor U26603 (N_26603,N_25095,N_25382);
and U26604 (N_26604,N_24784,N_24792);
xor U26605 (N_26605,N_24889,N_24862);
xor U26606 (N_26606,N_24210,N_24286);
nand U26607 (N_26607,N_24358,N_24749);
and U26608 (N_26608,N_25104,N_24272);
xnor U26609 (N_26609,N_24454,N_24627);
or U26610 (N_26610,N_24874,N_25259);
and U26611 (N_26611,N_25227,N_25389);
and U26612 (N_26612,N_24207,N_24437);
xor U26613 (N_26613,N_25416,N_24972);
nand U26614 (N_26614,N_24687,N_24918);
nand U26615 (N_26615,N_24895,N_25234);
xnor U26616 (N_26616,N_24015,N_24372);
nor U26617 (N_26617,N_24191,N_24283);
or U26618 (N_26618,N_24734,N_24467);
nor U26619 (N_26619,N_24909,N_24500);
xor U26620 (N_26620,N_25347,N_24913);
nor U26621 (N_26621,N_25167,N_24630);
nor U26622 (N_26622,N_24648,N_24278);
nand U26623 (N_26623,N_25436,N_24566);
xnor U26624 (N_26624,N_24922,N_24638);
nor U26625 (N_26625,N_24352,N_24915);
nand U26626 (N_26626,N_24011,N_24882);
or U26627 (N_26627,N_24764,N_25475);
nor U26628 (N_26628,N_24942,N_24979);
nor U26629 (N_26629,N_25227,N_25222);
and U26630 (N_26630,N_25315,N_25337);
nand U26631 (N_26631,N_24222,N_24794);
or U26632 (N_26632,N_24868,N_25116);
or U26633 (N_26633,N_25343,N_24220);
xnor U26634 (N_26634,N_25179,N_25273);
nand U26635 (N_26635,N_25119,N_24777);
nor U26636 (N_26636,N_25106,N_25026);
and U26637 (N_26637,N_24593,N_24911);
xor U26638 (N_26638,N_24722,N_25156);
nor U26639 (N_26639,N_25470,N_25406);
nand U26640 (N_26640,N_24236,N_24277);
nand U26641 (N_26641,N_24858,N_24822);
nand U26642 (N_26642,N_24800,N_24779);
xor U26643 (N_26643,N_24915,N_25326);
nor U26644 (N_26644,N_24697,N_24025);
and U26645 (N_26645,N_25301,N_24811);
nand U26646 (N_26646,N_25130,N_24895);
or U26647 (N_26647,N_24169,N_24783);
nand U26648 (N_26648,N_25369,N_25134);
and U26649 (N_26649,N_24595,N_24503);
and U26650 (N_26650,N_25016,N_25158);
xnor U26651 (N_26651,N_25138,N_25235);
and U26652 (N_26652,N_25377,N_24712);
nor U26653 (N_26653,N_24227,N_24156);
nor U26654 (N_26654,N_25157,N_24802);
xnor U26655 (N_26655,N_25449,N_24935);
or U26656 (N_26656,N_24211,N_24369);
or U26657 (N_26657,N_24041,N_24256);
nor U26658 (N_26658,N_24934,N_24206);
nand U26659 (N_26659,N_24291,N_24695);
xor U26660 (N_26660,N_24986,N_25204);
or U26661 (N_26661,N_24407,N_24665);
or U26662 (N_26662,N_25428,N_24570);
or U26663 (N_26663,N_24893,N_24163);
or U26664 (N_26664,N_24138,N_24836);
nand U26665 (N_26665,N_25469,N_24825);
xor U26666 (N_26666,N_24471,N_24734);
and U26667 (N_26667,N_24992,N_25158);
or U26668 (N_26668,N_25070,N_25455);
nor U26669 (N_26669,N_25193,N_24890);
or U26670 (N_26670,N_24803,N_24064);
and U26671 (N_26671,N_24192,N_25039);
nand U26672 (N_26672,N_24392,N_25395);
xnor U26673 (N_26673,N_24067,N_24565);
xnor U26674 (N_26674,N_24192,N_25470);
xor U26675 (N_26675,N_24534,N_24806);
and U26676 (N_26676,N_25113,N_24221);
and U26677 (N_26677,N_24877,N_24584);
nand U26678 (N_26678,N_25202,N_25115);
xor U26679 (N_26679,N_25337,N_24849);
xnor U26680 (N_26680,N_24925,N_24390);
nor U26681 (N_26681,N_25051,N_25133);
or U26682 (N_26682,N_24954,N_25100);
xnor U26683 (N_26683,N_24018,N_24686);
xor U26684 (N_26684,N_24763,N_24797);
nor U26685 (N_26685,N_25377,N_24571);
or U26686 (N_26686,N_25449,N_24448);
nor U26687 (N_26687,N_24774,N_24033);
or U26688 (N_26688,N_24987,N_24972);
xor U26689 (N_26689,N_24357,N_24588);
and U26690 (N_26690,N_25181,N_24734);
xor U26691 (N_26691,N_24051,N_24704);
nor U26692 (N_26692,N_25443,N_25231);
nand U26693 (N_26693,N_24333,N_24470);
and U26694 (N_26694,N_24066,N_25396);
nand U26695 (N_26695,N_25347,N_24455);
or U26696 (N_26696,N_24332,N_24193);
and U26697 (N_26697,N_24808,N_24215);
xnor U26698 (N_26698,N_24840,N_24532);
xnor U26699 (N_26699,N_24326,N_25092);
or U26700 (N_26700,N_24391,N_25498);
xor U26701 (N_26701,N_24284,N_24378);
and U26702 (N_26702,N_24803,N_24319);
and U26703 (N_26703,N_25342,N_25156);
and U26704 (N_26704,N_24555,N_25340);
nand U26705 (N_26705,N_24792,N_24370);
nand U26706 (N_26706,N_24635,N_25052);
and U26707 (N_26707,N_25347,N_25151);
nand U26708 (N_26708,N_25427,N_24946);
nor U26709 (N_26709,N_24049,N_25427);
nand U26710 (N_26710,N_24369,N_24996);
or U26711 (N_26711,N_24852,N_24698);
xor U26712 (N_26712,N_25323,N_24188);
nand U26713 (N_26713,N_25389,N_24460);
xnor U26714 (N_26714,N_24897,N_24801);
nand U26715 (N_26715,N_25071,N_24782);
nor U26716 (N_26716,N_24379,N_25026);
and U26717 (N_26717,N_24119,N_24091);
nor U26718 (N_26718,N_25310,N_24550);
or U26719 (N_26719,N_24686,N_24459);
and U26720 (N_26720,N_24304,N_24320);
and U26721 (N_26721,N_24859,N_24695);
nand U26722 (N_26722,N_25207,N_25123);
xnor U26723 (N_26723,N_24772,N_24716);
xor U26724 (N_26724,N_24483,N_24218);
nand U26725 (N_26725,N_24226,N_24757);
and U26726 (N_26726,N_24151,N_25281);
nand U26727 (N_26727,N_24267,N_24756);
and U26728 (N_26728,N_24143,N_25425);
xor U26729 (N_26729,N_24085,N_24197);
or U26730 (N_26730,N_24986,N_25252);
xor U26731 (N_26731,N_24122,N_24183);
or U26732 (N_26732,N_25033,N_24019);
and U26733 (N_26733,N_25236,N_24264);
nor U26734 (N_26734,N_24229,N_24528);
nand U26735 (N_26735,N_24121,N_24600);
xnor U26736 (N_26736,N_24260,N_25113);
nand U26737 (N_26737,N_25165,N_24391);
and U26738 (N_26738,N_25499,N_24666);
xor U26739 (N_26739,N_24267,N_24146);
nand U26740 (N_26740,N_24194,N_25322);
or U26741 (N_26741,N_24946,N_24977);
nor U26742 (N_26742,N_25452,N_24025);
nand U26743 (N_26743,N_24639,N_24420);
nand U26744 (N_26744,N_24110,N_25165);
nor U26745 (N_26745,N_24514,N_25040);
nand U26746 (N_26746,N_25243,N_25017);
and U26747 (N_26747,N_24053,N_24468);
or U26748 (N_26748,N_25171,N_24021);
xor U26749 (N_26749,N_24866,N_24810);
or U26750 (N_26750,N_25401,N_24610);
nor U26751 (N_26751,N_25479,N_25364);
or U26752 (N_26752,N_24676,N_24711);
or U26753 (N_26753,N_24949,N_24921);
nand U26754 (N_26754,N_24152,N_24572);
and U26755 (N_26755,N_24861,N_24063);
xor U26756 (N_26756,N_24183,N_24913);
and U26757 (N_26757,N_25467,N_25424);
or U26758 (N_26758,N_25323,N_24910);
nor U26759 (N_26759,N_24291,N_24396);
or U26760 (N_26760,N_25065,N_24856);
nand U26761 (N_26761,N_24511,N_24050);
nor U26762 (N_26762,N_24206,N_24432);
nand U26763 (N_26763,N_25452,N_25174);
or U26764 (N_26764,N_24869,N_24353);
nor U26765 (N_26765,N_24386,N_24985);
and U26766 (N_26766,N_24427,N_25132);
xnor U26767 (N_26767,N_25437,N_24412);
or U26768 (N_26768,N_24489,N_25280);
nor U26769 (N_26769,N_24310,N_24345);
xnor U26770 (N_26770,N_24582,N_24909);
or U26771 (N_26771,N_25493,N_24695);
xnor U26772 (N_26772,N_25135,N_25224);
and U26773 (N_26773,N_25059,N_25115);
or U26774 (N_26774,N_25070,N_24781);
and U26775 (N_26775,N_24227,N_25427);
nand U26776 (N_26776,N_24450,N_25072);
nor U26777 (N_26777,N_24222,N_24287);
nor U26778 (N_26778,N_25421,N_24055);
nor U26779 (N_26779,N_25283,N_24590);
nand U26780 (N_26780,N_25274,N_24103);
nor U26781 (N_26781,N_24345,N_24769);
and U26782 (N_26782,N_24120,N_24244);
nor U26783 (N_26783,N_24968,N_24029);
or U26784 (N_26784,N_25469,N_24916);
nand U26785 (N_26785,N_24044,N_25081);
and U26786 (N_26786,N_25361,N_25343);
or U26787 (N_26787,N_25401,N_25378);
nand U26788 (N_26788,N_24745,N_24175);
nand U26789 (N_26789,N_24916,N_24542);
and U26790 (N_26790,N_25151,N_24857);
or U26791 (N_26791,N_24832,N_24852);
xor U26792 (N_26792,N_24729,N_24748);
nor U26793 (N_26793,N_24700,N_24166);
or U26794 (N_26794,N_24575,N_24534);
nand U26795 (N_26795,N_24433,N_25047);
nor U26796 (N_26796,N_24206,N_24448);
nor U26797 (N_26797,N_25112,N_24194);
nor U26798 (N_26798,N_25059,N_24040);
or U26799 (N_26799,N_24869,N_24181);
nor U26800 (N_26800,N_24140,N_25021);
and U26801 (N_26801,N_24353,N_24432);
or U26802 (N_26802,N_24085,N_25103);
and U26803 (N_26803,N_24785,N_25012);
or U26804 (N_26804,N_24984,N_25303);
or U26805 (N_26805,N_25340,N_24374);
nand U26806 (N_26806,N_24883,N_24998);
nor U26807 (N_26807,N_24014,N_25324);
and U26808 (N_26808,N_24369,N_24057);
nor U26809 (N_26809,N_24712,N_24303);
xnor U26810 (N_26810,N_24216,N_24472);
xnor U26811 (N_26811,N_25020,N_24636);
or U26812 (N_26812,N_25178,N_24614);
xor U26813 (N_26813,N_24044,N_24804);
or U26814 (N_26814,N_24651,N_24388);
nand U26815 (N_26815,N_25102,N_24004);
or U26816 (N_26816,N_25427,N_25490);
nor U26817 (N_26817,N_24728,N_24860);
and U26818 (N_26818,N_24286,N_24237);
xor U26819 (N_26819,N_25196,N_24792);
or U26820 (N_26820,N_24913,N_24811);
and U26821 (N_26821,N_24069,N_24354);
nor U26822 (N_26822,N_25104,N_24750);
nand U26823 (N_26823,N_24754,N_24815);
nand U26824 (N_26824,N_24480,N_24869);
nand U26825 (N_26825,N_24150,N_24092);
xor U26826 (N_26826,N_24021,N_24324);
nand U26827 (N_26827,N_25007,N_24903);
xnor U26828 (N_26828,N_25416,N_25068);
nor U26829 (N_26829,N_25177,N_25116);
or U26830 (N_26830,N_24613,N_24641);
nand U26831 (N_26831,N_25446,N_24403);
nand U26832 (N_26832,N_24737,N_24834);
or U26833 (N_26833,N_24829,N_24485);
and U26834 (N_26834,N_24571,N_24650);
xnor U26835 (N_26835,N_24709,N_25415);
and U26836 (N_26836,N_24050,N_25434);
xor U26837 (N_26837,N_24351,N_25432);
or U26838 (N_26838,N_24783,N_24948);
and U26839 (N_26839,N_24290,N_24355);
xor U26840 (N_26840,N_24609,N_24598);
nand U26841 (N_26841,N_24992,N_24897);
or U26842 (N_26842,N_24591,N_25188);
nor U26843 (N_26843,N_24820,N_24684);
or U26844 (N_26844,N_24713,N_24418);
nor U26845 (N_26845,N_25413,N_25197);
xnor U26846 (N_26846,N_24259,N_25062);
or U26847 (N_26847,N_25095,N_24076);
nand U26848 (N_26848,N_24798,N_24157);
and U26849 (N_26849,N_24986,N_24289);
nand U26850 (N_26850,N_24369,N_25345);
nand U26851 (N_26851,N_25480,N_25034);
and U26852 (N_26852,N_24868,N_24542);
xnor U26853 (N_26853,N_25359,N_24923);
nor U26854 (N_26854,N_25367,N_24052);
nor U26855 (N_26855,N_24396,N_24419);
xnor U26856 (N_26856,N_24352,N_25376);
and U26857 (N_26857,N_25074,N_24300);
and U26858 (N_26858,N_25439,N_24743);
xor U26859 (N_26859,N_24313,N_24802);
nand U26860 (N_26860,N_24757,N_25324);
and U26861 (N_26861,N_24497,N_25268);
or U26862 (N_26862,N_24168,N_24431);
and U26863 (N_26863,N_25029,N_24458);
or U26864 (N_26864,N_25056,N_24254);
or U26865 (N_26865,N_24237,N_25365);
and U26866 (N_26866,N_24605,N_24912);
and U26867 (N_26867,N_24147,N_24646);
nor U26868 (N_26868,N_25129,N_24822);
nand U26869 (N_26869,N_24148,N_24139);
nand U26870 (N_26870,N_24852,N_25064);
xor U26871 (N_26871,N_25291,N_24375);
nor U26872 (N_26872,N_24434,N_24611);
nor U26873 (N_26873,N_24143,N_25054);
nor U26874 (N_26874,N_25306,N_24114);
nand U26875 (N_26875,N_24827,N_24383);
nor U26876 (N_26876,N_25395,N_24279);
or U26877 (N_26877,N_25077,N_24729);
nor U26878 (N_26878,N_25253,N_25035);
xor U26879 (N_26879,N_24050,N_24205);
and U26880 (N_26880,N_24806,N_24601);
or U26881 (N_26881,N_24916,N_24030);
or U26882 (N_26882,N_24115,N_24092);
or U26883 (N_26883,N_25082,N_24769);
and U26884 (N_26884,N_24726,N_24626);
and U26885 (N_26885,N_24969,N_25442);
nor U26886 (N_26886,N_25281,N_24879);
or U26887 (N_26887,N_24117,N_25488);
nor U26888 (N_26888,N_25279,N_24709);
nor U26889 (N_26889,N_24436,N_25177);
nor U26890 (N_26890,N_25384,N_25204);
nor U26891 (N_26891,N_24601,N_24966);
nor U26892 (N_26892,N_25207,N_25220);
nor U26893 (N_26893,N_24343,N_24903);
xor U26894 (N_26894,N_24642,N_24486);
nand U26895 (N_26895,N_24009,N_24278);
xnor U26896 (N_26896,N_25245,N_24836);
xnor U26897 (N_26897,N_25114,N_25493);
and U26898 (N_26898,N_25278,N_24111);
nor U26899 (N_26899,N_24778,N_25220);
nor U26900 (N_26900,N_25092,N_25182);
nand U26901 (N_26901,N_24847,N_25123);
nand U26902 (N_26902,N_24239,N_24583);
or U26903 (N_26903,N_24406,N_24925);
xor U26904 (N_26904,N_24658,N_24217);
xnor U26905 (N_26905,N_24590,N_25161);
nand U26906 (N_26906,N_25022,N_25069);
xnor U26907 (N_26907,N_25453,N_24851);
and U26908 (N_26908,N_24363,N_24567);
nand U26909 (N_26909,N_25229,N_25323);
xnor U26910 (N_26910,N_24942,N_24435);
nor U26911 (N_26911,N_25402,N_24486);
nor U26912 (N_26912,N_25129,N_25425);
or U26913 (N_26913,N_24355,N_24502);
nand U26914 (N_26914,N_25049,N_25052);
nor U26915 (N_26915,N_24788,N_24600);
and U26916 (N_26916,N_24484,N_25007);
xnor U26917 (N_26917,N_25300,N_24000);
and U26918 (N_26918,N_24229,N_24145);
nor U26919 (N_26919,N_24162,N_24646);
nor U26920 (N_26920,N_24489,N_25120);
xor U26921 (N_26921,N_24666,N_24037);
nand U26922 (N_26922,N_24783,N_25015);
nor U26923 (N_26923,N_25104,N_24030);
and U26924 (N_26924,N_24928,N_24315);
xor U26925 (N_26925,N_24368,N_25244);
or U26926 (N_26926,N_25227,N_24098);
xnor U26927 (N_26927,N_24860,N_24059);
and U26928 (N_26928,N_24960,N_24490);
xor U26929 (N_26929,N_24275,N_24873);
nand U26930 (N_26930,N_25490,N_24889);
and U26931 (N_26931,N_24084,N_24314);
and U26932 (N_26932,N_24799,N_25481);
xor U26933 (N_26933,N_25071,N_24137);
and U26934 (N_26934,N_24674,N_24212);
xnor U26935 (N_26935,N_25068,N_24231);
nand U26936 (N_26936,N_24952,N_24821);
nor U26937 (N_26937,N_24521,N_25175);
xor U26938 (N_26938,N_25333,N_25406);
or U26939 (N_26939,N_25243,N_24289);
nor U26940 (N_26940,N_25115,N_25462);
nand U26941 (N_26941,N_25070,N_25048);
and U26942 (N_26942,N_25195,N_25188);
nand U26943 (N_26943,N_25153,N_25190);
nor U26944 (N_26944,N_24069,N_24257);
and U26945 (N_26945,N_24435,N_25371);
and U26946 (N_26946,N_25320,N_25195);
or U26947 (N_26947,N_24623,N_24219);
and U26948 (N_26948,N_25006,N_25053);
or U26949 (N_26949,N_24781,N_24395);
nand U26950 (N_26950,N_24740,N_25241);
or U26951 (N_26951,N_25329,N_24417);
nor U26952 (N_26952,N_25100,N_24237);
or U26953 (N_26953,N_24429,N_25387);
nand U26954 (N_26954,N_24390,N_24794);
and U26955 (N_26955,N_25202,N_25447);
or U26956 (N_26956,N_24651,N_24669);
xnor U26957 (N_26957,N_24109,N_24633);
nand U26958 (N_26958,N_25065,N_25453);
and U26959 (N_26959,N_24949,N_25395);
or U26960 (N_26960,N_25207,N_25314);
nor U26961 (N_26961,N_24268,N_25306);
nor U26962 (N_26962,N_24075,N_24254);
xnor U26963 (N_26963,N_24887,N_24330);
nand U26964 (N_26964,N_24727,N_24019);
nor U26965 (N_26965,N_24654,N_25476);
nor U26966 (N_26966,N_24759,N_25310);
nor U26967 (N_26967,N_25480,N_24161);
and U26968 (N_26968,N_25219,N_24883);
nand U26969 (N_26969,N_24746,N_24742);
nor U26970 (N_26970,N_24379,N_24799);
nor U26971 (N_26971,N_25305,N_25486);
nand U26972 (N_26972,N_24358,N_25236);
nand U26973 (N_26973,N_24040,N_24194);
nand U26974 (N_26974,N_24141,N_24253);
or U26975 (N_26975,N_24950,N_24198);
or U26976 (N_26976,N_24313,N_24004);
or U26977 (N_26977,N_25225,N_25418);
xnor U26978 (N_26978,N_24679,N_25112);
nand U26979 (N_26979,N_25398,N_24373);
or U26980 (N_26980,N_24097,N_24421);
and U26981 (N_26981,N_24313,N_24905);
and U26982 (N_26982,N_25430,N_24197);
nor U26983 (N_26983,N_24907,N_24947);
nor U26984 (N_26984,N_24765,N_24772);
xor U26985 (N_26985,N_24456,N_24040);
nand U26986 (N_26986,N_24919,N_25260);
and U26987 (N_26987,N_25142,N_25436);
or U26988 (N_26988,N_24076,N_25218);
xor U26989 (N_26989,N_24775,N_24189);
and U26990 (N_26990,N_25495,N_24091);
and U26991 (N_26991,N_25228,N_24882);
nand U26992 (N_26992,N_25357,N_24288);
xor U26993 (N_26993,N_24659,N_24121);
and U26994 (N_26994,N_24670,N_24100);
nor U26995 (N_26995,N_24185,N_24639);
nor U26996 (N_26996,N_24918,N_24799);
or U26997 (N_26997,N_25119,N_25193);
or U26998 (N_26998,N_25388,N_24713);
nand U26999 (N_26999,N_25046,N_25420);
nand U27000 (N_27000,N_26393,N_25590);
nand U27001 (N_27001,N_26414,N_25545);
and U27002 (N_27002,N_26506,N_26047);
xor U27003 (N_27003,N_26424,N_25713);
nand U27004 (N_27004,N_26958,N_26824);
nor U27005 (N_27005,N_26591,N_26560);
or U27006 (N_27006,N_26607,N_26267);
xnor U27007 (N_27007,N_25555,N_25518);
xnor U27008 (N_27008,N_25591,N_25541);
nand U27009 (N_27009,N_25832,N_25919);
and U27010 (N_27010,N_26880,N_26777);
xor U27011 (N_27011,N_26054,N_26293);
and U27012 (N_27012,N_26355,N_25695);
xnor U27013 (N_27013,N_26905,N_26305);
and U27014 (N_27014,N_26222,N_26615);
xor U27015 (N_27015,N_26767,N_26096);
or U27016 (N_27016,N_26939,N_26733);
or U27017 (N_27017,N_26609,N_26704);
nor U27018 (N_27018,N_25965,N_25781);
and U27019 (N_27019,N_26045,N_26566);
nor U27020 (N_27020,N_26543,N_26041);
nor U27021 (N_27021,N_25831,N_25791);
nor U27022 (N_27022,N_26493,N_26116);
or U27023 (N_27023,N_25735,N_26515);
and U27024 (N_27024,N_26776,N_25905);
and U27025 (N_27025,N_26636,N_25893);
and U27026 (N_27026,N_26627,N_26429);
nor U27027 (N_27027,N_26729,N_25613);
or U27028 (N_27028,N_26849,N_26943);
and U27029 (N_27029,N_26915,N_25853);
and U27030 (N_27030,N_26783,N_26873);
and U27031 (N_27031,N_25951,N_26401);
xor U27032 (N_27032,N_25849,N_26082);
xor U27033 (N_27033,N_26223,N_26160);
and U27034 (N_27034,N_26086,N_26078);
and U27035 (N_27035,N_25921,N_26265);
or U27036 (N_27036,N_26145,N_26341);
nor U27037 (N_27037,N_26388,N_26790);
nand U27038 (N_27038,N_26641,N_25516);
nand U27039 (N_27039,N_26487,N_25614);
or U27040 (N_27040,N_26469,N_26765);
and U27041 (N_27041,N_26422,N_26276);
or U27042 (N_27042,N_26376,N_26108);
and U27043 (N_27043,N_26976,N_26471);
xnor U27044 (N_27044,N_26716,N_26978);
xor U27045 (N_27045,N_26373,N_26220);
or U27046 (N_27046,N_25856,N_26295);
or U27047 (N_27047,N_26121,N_26157);
nand U27048 (N_27048,N_26892,N_25773);
or U27049 (N_27049,N_25762,N_26021);
nor U27050 (N_27050,N_25631,N_25928);
nand U27051 (N_27051,N_26059,N_25754);
nor U27052 (N_27052,N_26044,N_26191);
or U27053 (N_27053,N_25747,N_25519);
nor U27054 (N_27054,N_26080,N_25764);
nor U27055 (N_27055,N_25912,N_26094);
and U27056 (N_27056,N_26536,N_26252);
and U27057 (N_27057,N_26372,N_25979);
or U27058 (N_27058,N_26707,N_26544);
and U27059 (N_27059,N_26375,N_25530);
xnor U27060 (N_27060,N_26092,N_25500);
nand U27061 (N_27061,N_26759,N_26511);
and U27062 (N_27062,N_25927,N_25734);
or U27063 (N_27063,N_26495,N_26194);
and U27064 (N_27064,N_26143,N_26822);
or U27065 (N_27065,N_26226,N_26365);
nor U27066 (N_27066,N_25971,N_26940);
or U27067 (N_27067,N_26137,N_25604);
nor U27068 (N_27068,N_25535,N_26533);
xnor U27069 (N_27069,N_25926,N_25743);
and U27070 (N_27070,N_25917,N_26012);
or U27071 (N_27071,N_25858,N_26296);
and U27072 (N_27072,N_25967,N_26903);
xor U27073 (N_27073,N_25878,N_25548);
xor U27074 (N_27074,N_26768,N_26735);
nor U27075 (N_27075,N_25969,N_26039);
and U27076 (N_27076,N_26348,N_25938);
nand U27077 (N_27077,N_26957,N_26250);
nand U27078 (N_27078,N_25987,N_25824);
nor U27079 (N_27079,N_25520,N_25793);
and U27080 (N_27080,N_26804,N_26952);
or U27081 (N_27081,N_25911,N_26407);
nor U27082 (N_27082,N_26269,N_25589);
or U27083 (N_27083,N_25801,N_25939);
or U27084 (N_27084,N_25780,N_25986);
nand U27085 (N_27085,N_25887,N_26251);
nor U27086 (N_27086,N_26572,N_25771);
or U27087 (N_27087,N_25746,N_26344);
nor U27088 (N_27088,N_26553,N_25855);
or U27089 (N_27089,N_26263,N_25636);
and U27090 (N_27090,N_26473,N_26899);
nor U27091 (N_27091,N_26842,N_25885);
or U27092 (N_27092,N_26606,N_26070);
nor U27093 (N_27093,N_26910,N_26608);
nand U27094 (N_27094,N_26749,N_26686);
nand U27095 (N_27095,N_25606,N_25852);
and U27096 (N_27096,N_25526,N_26925);
nand U27097 (N_27097,N_26254,N_25826);
and U27098 (N_27098,N_26245,N_26173);
xor U27099 (N_27099,N_25662,N_26256);
or U27100 (N_27100,N_26383,N_26288);
xor U27101 (N_27101,N_26156,N_26814);
nand U27102 (N_27102,N_25633,N_25661);
or U27103 (N_27103,N_26498,N_25597);
and U27104 (N_27104,N_25786,N_26834);
xor U27105 (N_27105,N_26603,N_26219);
and U27106 (N_27106,N_26400,N_26117);
or U27107 (N_27107,N_26638,N_25685);
nor U27108 (N_27108,N_26866,N_26587);
nand U27109 (N_27109,N_26539,N_25894);
or U27110 (N_27110,N_26022,N_26843);
nor U27111 (N_27111,N_26546,N_26404);
nand U27112 (N_27112,N_26476,N_26514);
nand U27113 (N_27113,N_25766,N_26505);
or U27114 (N_27114,N_26908,N_26653);
or U27115 (N_27115,N_26294,N_26530);
or U27116 (N_27116,N_26942,N_26218);
and U27117 (N_27117,N_26490,N_25991);
nor U27118 (N_27118,N_26684,N_25671);
and U27119 (N_27119,N_26483,N_26941);
nand U27120 (N_27120,N_26115,N_26929);
or U27121 (N_27121,N_25580,N_26172);
and U27122 (N_27122,N_25513,N_25783);
and U27123 (N_27123,N_25611,N_26797);
and U27124 (N_27124,N_26273,N_26153);
or U27125 (N_27125,N_25630,N_25770);
nand U27126 (N_27126,N_26053,N_26510);
nor U27127 (N_27127,N_25720,N_25542);
nand U27128 (N_27128,N_26077,N_25659);
or U27129 (N_27129,N_26324,N_25952);
and U27130 (N_27130,N_26014,N_25594);
or U27131 (N_27131,N_25554,N_26738);
nor U27132 (N_27132,N_26809,N_25994);
nand U27133 (N_27133,N_25634,N_26712);
nor U27134 (N_27134,N_26158,N_26730);
nor U27135 (N_27135,N_25515,N_25942);
xnor U27136 (N_27136,N_26060,N_25607);
and U27137 (N_27137,N_25930,N_26489);
nand U27138 (N_27138,N_26036,N_25903);
nand U27139 (N_27139,N_25523,N_26146);
xnor U27140 (N_27140,N_25683,N_26675);
nor U27141 (N_27141,N_26737,N_25948);
nor U27142 (N_27142,N_25829,N_25578);
xnor U27143 (N_27143,N_26188,N_26995);
xnor U27144 (N_27144,N_26678,N_26408);
xor U27145 (N_27145,N_25745,N_26631);
and U27146 (N_27146,N_25857,N_26329);
nand U27147 (N_27147,N_25937,N_26669);
and U27148 (N_27148,N_26437,N_25947);
nand U27149 (N_27149,N_26154,N_26075);
and U27150 (N_27150,N_25749,N_26823);
nand U27151 (N_27151,N_25755,N_26922);
xnor U27152 (N_27152,N_26171,N_26275);
xnor U27153 (N_27153,N_26272,N_25505);
nand U27154 (N_27154,N_26150,N_25510);
nor U27155 (N_27155,N_25645,N_25897);
or U27156 (N_27156,N_25813,N_26229);
xor U27157 (N_27157,N_25816,N_25815);
or U27158 (N_27158,N_26859,N_26991);
or U27159 (N_27159,N_26364,N_25504);
nand U27160 (N_27160,N_26628,N_26766);
nand U27161 (N_27161,N_26332,N_25776);
or U27162 (N_27162,N_25668,N_26479);
nor U27163 (N_27163,N_25888,N_26185);
xor U27164 (N_27164,N_26353,N_26527);
and U27165 (N_27165,N_26512,N_26984);
or U27166 (N_27166,N_25546,N_25559);
xnor U27167 (N_27167,N_26443,N_26581);
and U27168 (N_27168,N_26474,N_26019);
nand U27169 (N_27169,N_25709,N_26855);
and U27170 (N_27170,N_26719,N_26690);
or U27171 (N_27171,N_25981,N_26118);
or U27172 (N_27172,N_26284,N_26465);
nand U27173 (N_27173,N_25648,N_26649);
or U27174 (N_27174,N_25900,N_26655);
xor U27175 (N_27175,N_26755,N_25616);
and U27176 (N_27176,N_26240,N_26023);
or U27177 (N_27177,N_25737,N_25906);
xnor U27178 (N_27178,N_25875,N_26983);
or U27179 (N_27179,N_26061,N_26720);
and U27180 (N_27180,N_26805,N_26356);
nor U27181 (N_27181,N_26389,N_26379);
nor U27182 (N_27182,N_25644,N_25988);
or U27183 (N_27183,N_25689,N_25882);
xnor U27184 (N_27184,N_26852,N_26643);
xnor U27185 (N_27185,N_25723,N_26330);
and U27186 (N_27186,N_25717,N_25627);
nor U27187 (N_27187,N_26588,N_25797);
or U27188 (N_27188,N_26614,N_25840);
xor U27189 (N_27189,N_25909,N_26837);
nor U27190 (N_27190,N_26531,N_26415);
or U27191 (N_27191,N_26676,N_26613);
and U27192 (N_27192,N_26385,N_26697);
or U27193 (N_27193,N_26016,N_25638);
and U27194 (N_27194,N_25585,N_26111);
xor U27195 (N_27195,N_25821,N_26968);
nor U27196 (N_27196,N_26327,N_26017);
nor U27197 (N_27197,N_26625,N_25656);
or U27198 (N_27198,N_26782,N_26996);
xor U27199 (N_27199,N_25949,N_26889);
xor U27200 (N_27200,N_25890,N_26034);
and U27201 (N_27201,N_26828,N_26723);
and U27202 (N_27202,N_25836,N_26312);
and U27203 (N_27203,N_26442,N_26342);
and U27204 (N_27204,N_26419,N_26313);
xor U27205 (N_27205,N_26988,N_26985);
and U27206 (N_27206,N_26854,N_26516);
and U27207 (N_27207,N_25751,N_25758);
nor U27208 (N_27208,N_26541,N_25583);
xor U27209 (N_27209,N_25769,N_26593);
nand U27210 (N_27210,N_26763,N_25883);
xnor U27211 (N_27211,N_26425,N_25624);
nand U27212 (N_27212,N_26545,N_26128);
nor U27213 (N_27213,N_26197,N_25864);
or U27214 (N_27214,N_26569,N_25525);
nand U27215 (N_27215,N_26700,N_25936);
and U27216 (N_27216,N_26107,N_26326);
nor U27217 (N_27217,N_26243,N_25785);
nor U27218 (N_27218,N_26048,N_25778);
nor U27219 (N_27219,N_25753,N_26529);
and U27220 (N_27220,N_26278,N_25724);
xor U27221 (N_27221,N_25910,N_26001);
and U27222 (N_27222,N_26213,N_25881);
nor U27223 (N_27223,N_26024,N_26413);
nand U27224 (N_27224,N_25929,N_25584);
and U27225 (N_27225,N_25920,N_26167);
or U27226 (N_27226,N_26549,N_26580);
or U27227 (N_27227,N_26605,N_26785);
xor U27228 (N_27228,N_25649,N_26386);
and U27229 (N_27229,N_26253,N_26138);
xor U27230 (N_27230,N_25711,N_26203);
and U27231 (N_27231,N_26110,N_26890);
xor U27232 (N_27232,N_25923,N_25643);
xor U27233 (N_27233,N_26011,N_26321);
and U27234 (N_27234,N_26893,N_26930);
xor U27235 (N_27235,N_26722,N_25694);
or U27236 (N_27236,N_26277,N_26377);
or U27237 (N_27237,N_26395,N_25573);
nor U27238 (N_27238,N_26031,N_26444);
nand U27239 (N_27239,N_25845,N_25690);
or U27240 (N_27240,N_26283,N_26761);
nor U27241 (N_27241,N_26144,N_26583);
nor U27242 (N_27242,N_25602,N_26318);
and U27243 (N_27243,N_26225,N_25658);
xor U27244 (N_27244,N_25664,N_26242);
xor U27245 (N_27245,N_26702,N_26100);
nand U27246 (N_27246,N_25529,N_25763);
nand U27247 (N_27247,N_26463,N_26064);
xor U27248 (N_27248,N_26298,N_26708);
xor U27249 (N_27249,N_25802,N_26447);
xor U27250 (N_27250,N_26752,N_25731);
or U27251 (N_27251,N_26000,N_25739);
and U27252 (N_27252,N_26450,N_25729);
nand U27253 (N_27253,N_25847,N_25679);
nand U27254 (N_27254,N_25944,N_26207);
and U27255 (N_27255,N_26847,N_26066);
or U27256 (N_27256,N_26848,N_26973);
xnor U27257 (N_27257,N_26670,N_26799);
nand U27258 (N_27258,N_25830,N_26459);
and U27259 (N_27259,N_26956,N_26148);
nor U27260 (N_27260,N_25953,N_26087);
nand U27261 (N_27261,N_25972,N_25677);
or U27262 (N_27262,N_26586,N_25886);
xnor U27263 (N_27263,N_26548,N_25703);
nand U27264 (N_27264,N_25581,N_26946);
and U27265 (N_27265,N_26637,N_26891);
or U27266 (N_27266,N_25609,N_25788);
xor U27267 (N_27267,N_26113,N_26647);
and U27268 (N_27268,N_26705,N_26757);
nand U27269 (N_27269,N_26525,N_26951);
or U27270 (N_27270,N_25637,N_26507);
xor U27271 (N_27271,N_26482,N_26975);
nor U27272 (N_27272,N_26102,N_25619);
and U27273 (N_27273,N_26683,N_26534);
xnor U27274 (N_27274,N_26500,N_26551);
or U27275 (N_27275,N_26056,N_26879);
nor U27276 (N_27276,N_26709,N_26181);
and U27277 (N_27277,N_25667,N_26909);
or U27278 (N_27278,N_26468,N_25896);
or U27279 (N_27279,N_26745,N_25895);
nand U27280 (N_27280,N_26556,N_26165);
nor U27281 (N_27281,N_26202,N_25588);
xnor U27282 (N_27282,N_26212,N_26331);
and U27283 (N_27283,N_26695,N_26867);
and U27284 (N_27284,N_26953,N_25511);
xor U27285 (N_27285,N_26004,N_25782);
or U27286 (N_27286,N_26542,N_25865);
and U27287 (N_27287,N_25652,N_25579);
nand U27288 (N_27288,N_26597,N_25543);
or U27289 (N_27289,N_25742,N_25876);
or U27290 (N_27290,N_25880,N_26950);
nor U27291 (N_27291,N_25684,N_26561);
xnor U27292 (N_27292,N_26792,N_26055);
nand U27293 (N_27293,N_26285,N_26453);
and U27294 (N_27294,N_26457,N_25859);
nor U27295 (N_27295,N_25531,N_26679);
and U27296 (N_27296,N_26199,N_26441);
nor U27297 (N_27297,N_26876,N_26345);
or U27298 (N_27298,N_26451,N_26945);
nor U27299 (N_27299,N_25725,N_25941);
xnor U27300 (N_27300,N_25985,N_26472);
xor U27301 (N_27301,N_26926,N_26521);
and U27302 (N_27302,N_26504,N_25809);
and U27303 (N_27303,N_25561,N_26286);
or U27304 (N_27304,N_25733,N_26035);
nand U27305 (N_27305,N_26937,N_26622);
xnor U27306 (N_27306,N_26431,N_26200);
or U27307 (N_27307,N_25973,N_25521);
or U27308 (N_27308,N_25657,N_25784);
nor U27309 (N_27309,N_25592,N_26274);
or U27310 (N_27310,N_26193,N_25756);
and U27311 (N_27311,N_25870,N_25873);
nor U27312 (N_27312,N_26582,N_25595);
xor U27313 (N_27313,N_26865,N_25915);
xor U27314 (N_27314,N_26570,N_26858);
and U27315 (N_27315,N_26142,N_25699);
nor U27316 (N_27316,N_26399,N_26833);
nand U27317 (N_27317,N_26180,N_26994);
and U27318 (N_27318,N_25946,N_25945);
and U27319 (N_27319,N_25999,N_26680);
nand U27320 (N_27320,N_26906,N_26006);
nand U27321 (N_27321,N_26503,N_26300);
nor U27322 (N_27322,N_26965,N_25673);
xor U27323 (N_27323,N_26619,N_26772);
and U27324 (N_27324,N_25736,N_25572);
xor U27325 (N_27325,N_26693,N_25678);
nand U27326 (N_27326,N_26677,N_26452);
xor U27327 (N_27327,N_26519,N_26791);
nand U27328 (N_27328,N_26416,N_26800);
xnor U27329 (N_27329,N_25995,N_26911);
nand U27330 (N_27330,N_26186,N_26499);
nand U27331 (N_27331,N_26887,N_26992);
xor U27332 (N_27332,N_26576,N_26462);
nand U27333 (N_27333,N_26596,N_26961);
or U27334 (N_27334,N_26163,N_26161);
nand U27335 (N_27335,N_26125,N_26747);
xor U27336 (N_27336,N_26317,N_26552);
nor U27337 (N_27337,N_26717,N_25696);
or U27338 (N_27338,N_25715,N_26362);
nor U27339 (N_27339,N_26394,N_26564);
xnor U27340 (N_27340,N_26592,N_26756);
or U27341 (N_27341,N_26106,N_26502);
or U27342 (N_27342,N_26139,N_26827);
nor U27343 (N_27343,N_25931,N_26105);
and U27344 (N_27344,N_25646,N_25688);
nand U27345 (N_27345,N_26657,N_26518);
nand U27346 (N_27346,N_26338,N_26853);
and U27347 (N_27347,N_25804,N_25760);
nand U27348 (N_27348,N_25807,N_25538);
and U27349 (N_27349,N_25798,N_26897);
nor U27350 (N_27350,N_25838,N_25502);
nand U27351 (N_27351,N_26179,N_25655);
nor U27352 (N_27352,N_25547,N_26538);
xnor U27353 (N_27353,N_26497,N_26812);
xor U27354 (N_27354,N_25539,N_26248);
nand U27355 (N_27355,N_25997,N_26685);
nor U27356 (N_27356,N_26184,N_26058);
or U27357 (N_27357,N_26175,N_26639);
nand U27358 (N_27358,N_26434,N_26878);
xnor U27359 (N_27359,N_25514,N_26771);
and U27360 (N_27360,N_26802,N_26754);
xnor U27361 (N_27361,N_26018,N_25775);
nor U27362 (N_27362,N_25962,N_26780);
nand U27363 (N_27363,N_26646,N_26980);
nor U27364 (N_27364,N_26857,N_26005);
nand U27365 (N_27365,N_26346,N_26862);
and U27366 (N_27366,N_26602,N_26632);
nand U27367 (N_27367,N_25833,N_26454);
or U27368 (N_27368,N_25978,N_26931);
nor U27369 (N_27369,N_26691,N_26666);
nand U27370 (N_27370,N_25586,N_26319);
nor U27371 (N_27371,N_26601,N_26798);
nand U27372 (N_27372,N_25846,N_26303);
nand U27373 (N_27373,N_25794,N_26784);
and U27374 (N_27374,N_26938,N_26470);
or U27375 (N_27375,N_26164,N_26692);
or U27376 (N_27376,N_26336,N_26239);
and U27377 (N_27377,N_26289,N_26508);
nor U27378 (N_27378,N_25792,N_25869);
xor U27379 (N_27379,N_26612,N_26032);
or U27380 (N_27380,N_25839,N_26883);
nand U27381 (N_27381,N_25710,N_25692);
nand U27382 (N_27382,N_26370,N_26458);
and U27383 (N_27383,N_25593,N_26266);
or U27384 (N_27384,N_26645,N_26122);
xnor U27385 (N_27385,N_26020,N_26725);
nand U27386 (N_27386,N_26829,N_26037);
nor U27387 (N_27387,N_26013,N_26562);
and U27388 (N_27388,N_26083,N_26900);
and U27389 (N_27389,N_25556,N_26871);
xnor U27390 (N_27390,N_25621,N_25551);
nor U27391 (N_27391,N_25669,N_25680);
and U27392 (N_27392,N_26119,N_26159);
nor U27393 (N_27393,N_26682,N_26896);
and U27394 (N_27394,N_26744,N_26532);
nand U27395 (N_27395,N_26262,N_26674);
xnor U27396 (N_27396,N_26933,N_26196);
or U27397 (N_27397,N_26721,N_25603);
xor U27398 (N_27398,N_26381,N_26921);
nor U27399 (N_27399,N_26368,N_26071);
xor U27400 (N_27400,N_26033,N_25601);
and U27401 (N_27401,N_25706,N_25716);
and U27402 (N_27402,N_26412,N_26466);
and U27403 (N_27403,N_25557,N_26478);
nor U27404 (N_27404,N_26127,N_25777);
nor U27405 (N_27405,N_26971,N_25512);
nor U27406 (N_27406,N_26281,N_26358);
xnor U27407 (N_27407,N_25629,N_25626);
nor U27408 (N_27408,N_25767,N_26072);
and U27409 (N_27409,N_25740,N_26270);
xor U27410 (N_27410,N_25732,N_25622);
xnor U27411 (N_27411,N_26189,N_26810);
or U27412 (N_27412,N_26448,N_26480);
and U27413 (N_27413,N_26114,N_26435);
xnor U27414 (N_27414,N_26818,N_26673);
and U27415 (N_27415,N_26563,N_25922);
nand U27416 (N_27416,N_26732,N_25958);
nand U27417 (N_27417,N_26820,N_26559);
xnor U27418 (N_27418,N_25811,N_26815);
xnor U27419 (N_27419,N_25899,N_26947);
nor U27420 (N_27420,N_26109,N_26291);
or U27421 (N_27421,N_26367,N_25765);
xnor U27422 (N_27422,N_26015,N_26456);
nand U27423 (N_27423,N_26714,N_26651);
xor U27424 (N_27424,N_25774,N_26069);
and U27425 (N_27425,N_25641,N_26467);
nand U27426 (N_27426,N_26860,N_26042);
xor U27427 (N_27427,N_25814,N_26793);
xnor U27428 (N_27428,N_25730,N_26540);
xnor U27429 (N_27429,N_25748,N_26773);
xor U27430 (N_27430,N_26287,N_26085);
and U27431 (N_27431,N_26183,N_25674);
nor U27432 (N_27432,N_26875,N_26152);
xor U27433 (N_27433,N_26134,N_26417);
and U27434 (N_27434,N_25924,N_26369);
or U27435 (N_27435,N_26192,N_25795);
nand U27436 (N_27436,N_26919,N_26650);
nor U27437 (N_27437,N_26681,N_26936);
nand U27438 (N_27438,N_26104,N_26492);
or U27439 (N_27439,N_26314,N_26120);
and U27440 (N_27440,N_26758,N_25620);
xor U27441 (N_27441,N_26297,N_26170);
nor U27442 (N_27442,N_25600,N_26839);
and U27443 (N_27443,N_26124,N_25835);
nor U27444 (N_27444,N_25841,N_25983);
or U27445 (N_27445,N_26352,N_25956);
xor U27446 (N_27446,N_25892,N_25570);
xnor U27447 (N_27447,N_25898,N_25761);
nor U27448 (N_27448,N_26611,N_26520);
xor U27449 (N_27449,N_26049,N_26604);
xor U27450 (N_27450,N_25722,N_26308);
xnor U27451 (N_27451,N_25618,N_26881);
or U27452 (N_27452,N_25850,N_26050);
nor U27453 (N_27453,N_26347,N_26418);
xnor U27454 (N_27454,N_25560,N_25860);
xnor U27455 (N_27455,N_25822,N_26660);
nand U27456 (N_27456,N_26236,N_26509);
nand U27457 (N_27457,N_26140,N_25540);
nand U27458 (N_27458,N_26201,N_26863);
xnor U27459 (N_27459,N_25503,N_25727);
nor U27460 (N_27460,N_26391,N_26969);
xnor U27461 (N_27461,N_26221,N_26535);
nand U27462 (N_27462,N_26885,N_25827);
nand U27463 (N_27463,N_25960,N_26097);
xor U27464 (N_27464,N_26359,N_26571);
and U27465 (N_27465,N_25779,N_26962);
or U27466 (N_27466,N_26232,N_26960);
nand U27467 (N_27467,N_26068,N_26496);
nor U27468 (N_27468,N_26486,N_25536);
or U27469 (N_27469,N_26403,N_26234);
or U27470 (N_27470,N_26652,N_26598);
and U27471 (N_27471,N_26568,N_26501);
nor U27472 (N_27472,N_25741,N_26577);
nand U27473 (N_27473,N_26028,N_25702);
nor U27474 (N_27474,N_25863,N_26112);
xnor U27475 (N_27475,N_25562,N_26565);
and U27476 (N_27476,N_26610,N_25553);
and U27477 (N_27477,N_26662,N_26898);
nor U27478 (N_27478,N_26811,N_26384);
nand U27479 (N_27479,N_26816,N_26629);
xnor U27480 (N_27480,N_26029,N_26715);
xnor U27481 (N_27481,N_26279,N_25625);
nor U27482 (N_27482,N_26131,N_26846);
and U27483 (N_27483,N_26233,N_25612);
and U27484 (N_27484,N_26009,N_26406);
and U27485 (N_27485,N_25916,N_25744);
or U27486 (N_27486,N_26409,N_26932);
xor U27487 (N_27487,N_26410,N_26257);
xnor U27488 (N_27488,N_25955,N_25508);
nand U27489 (N_27489,N_25660,N_25700);
or U27490 (N_27490,N_26485,N_26067);
nor U27491 (N_27491,N_26522,N_25918);
and U27492 (N_27492,N_26205,N_26076);
nor U27493 (N_27493,N_25635,N_25992);
and U27494 (N_27494,N_26882,N_25989);
and U27495 (N_27495,N_26917,N_26363);
and U27496 (N_27496,N_26040,N_26579);
nor U27497 (N_27497,N_26654,N_25817);
nor U27498 (N_27498,N_26557,N_26706);
nor U27499 (N_27499,N_26360,N_25799);
nor U27500 (N_27500,N_25834,N_26944);
or U27501 (N_27501,N_25707,N_26149);
and U27502 (N_27502,N_26635,N_26282);
or U27503 (N_27503,N_26043,N_26206);
nor U27504 (N_27504,N_26840,N_25963);
or U27505 (N_27505,N_26803,N_26710);
and U27506 (N_27506,N_25933,N_26091);
xor U27507 (N_27507,N_26090,N_25615);
or U27508 (N_27508,N_26268,N_26982);
and U27509 (N_27509,N_26558,N_25522);
xor U27510 (N_27510,N_26132,N_26258);
or U27511 (N_27511,N_25726,N_25577);
or U27512 (N_27512,N_26130,N_26786);
xor U27513 (N_27513,N_25768,N_25819);
or U27514 (N_27514,N_26698,N_26665);
xnor U27515 (N_27515,N_26624,N_26238);
and U27516 (N_27516,N_26081,N_26585);
and U27517 (N_27517,N_25701,N_26806);
nor U27518 (N_27518,N_26309,N_25718);
xor U27519 (N_27519,N_25848,N_26063);
nand U27520 (N_27520,N_26057,N_26868);
and U27521 (N_27521,N_25823,N_26301);
xnor U27522 (N_27522,N_26169,N_26764);
nand U27523 (N_27523,N_26623,N_26151);
or U27524 (N_27524,N_26398,N_26819);
xnor U27525 (N_27525,N_26328,N_26007);
nor U27526 (N_27526,N_26433,N_26870);
nor U27527 (N_27527,N_26633,N_25872);
nand U27528 (N_27528,N_26280,N_26397);
nand U27529 (N_27529,N_25549,N_26010);
xnor U27530 (N_27530,N_25705,N_26966);
or U27531 (N_27531,N_25566,N_26038);
nor U27532 (N_27532,N_26230,N_26550);
nor U27533 (N_27533,N_26382,N_25984);
xnor U27534 (N_27534,N_26977,N_25708);
nand U27535 (N_27535,N_25750,N_25837);
xor U27536 (N_27536,N_25582,N_25576);
xor U27537 (N_27537,N_25874,N_26974);
nor U27538 (N_27538,N_25868,N_26775);
nand U27539 (N_27539,N_26689,N_26748);
nor U27540 (N_27540,N_25796,N_26209);
xor U27541 (N_27541,N_26361,N_26640);
or U27542 (N_27542,N_26322,N_25975);
or U27543 (N_27543,N_25805,N_25563);
or U27544 (N_27544,N_26850,N_26595);
or U27545 (N_27545,N_25528,N_26888);
nor U27546 (N_27546,N_26333,N_26260);
nand U27547 (N_27547,N_26794,N_26074);
and U27548 (N_27548,N_25574,N_26307);
and U27549 (N_27549,N_26224,N_26003);
xor U27550 (N_27550,N_26584,N_25532);
xnor U27551 (N_27551,N_26101,N_26664);
nor U27552 (N_27552,N_25666,N_26573);
and U27553 (N_27553,N_25907,N_26030);
nand U27554 (N_27554,N_26455,N_26065);
xor U27555 (N_27555,N_26726,N_26445);
nand U27556 (N_27556,N_26026,N_26769);
or U27557 (N_27557,N_26575,N_25617);
nand U27558 (N_27558,N_26554,N_26098);
xnor U27559 (N_27559,N_26343,N_26851);
xnor U27560 (N_27560,N_26694,N_26727);
and U27561 (N_27561,N_25552,N_25914);
xnor U27562 (N_27562,N_26599,N_25569);
nor U27563 (N_27563,N_25810,N_26902);
or U27564 (N_27564,N_26845,N_25966);
and U27565 (N_27565,N_25990,N_26736);
xnor U27566 (N_27566,N_26162,N_26350);
or U27567 (N_27567,N_26084,N_25908);
xnor U27568 (N_27568,N_25654,N_26970);
nor U27569 (N_27569,N_25861,N_26427);
or U27570 (N_27570,N_26449,N_25934);
nor U27571 (N_27571,N_26830,N_26241);
nand U27572 (N_27572,N_25501,N_26133);
nor U27573 (N_27573,N_26177,N_25940);
or U27574 (N_27574,N_26366,N_26796);
nand U27575 (N_27575,N_26195,N_26739);
nand U27576 (N_27576,N_25558,N_26340);
xnor U27577 (N_27577,N_26841,N_26877);
nor U27578 (N_27578,N_26430,N_26711);
or U27579 (N_27579,N_26831,N_26774);
nand U27580 (N_27580,N_26832,N_26299);
xor U27581 (N_27581,N_26825,N_26630);
nand U27582 (N_27582,N_26949,N_26923);
nor U27583 (N_27583,N_26204,N_26616);
nor U27584 (N_27584,N_25672,N_26967);
and U27585 (N_27585,N_26661,N_25675);
or U27586 (N_27586,N_26523,N_26642);
and U27587 (N_27587,N_25653,N_26316);
and U27588 (N_27588,N_26981,N_26948);
or U27589 (N_27589,N_25623,N_26964);
and U27590 (N_27590,N_26237,N_26126);
xnor U27591 (N_27591,N_26390,N_25676);
or U27592 (N_27592,N_26979,N_25698);
or U27593 (N_27593,N_25803,N_25533);
and U27594 (N_27594,N_25943,N_26537);
nand U27595 (N_27595,N_26713,N_25728);
and U27596 (N_27596,N_25565,N_25998);
and U27597 (N_27597,N_26198,N_25681);
or U27598 (N_27598,N_26380,N_26872);
nand U27599 (N_27599,N_25902,N_26339);
xnor U27600 (N_27600,N_25808,N_26208);
and U27601 (N_27601,N_25599,N_26216);
nor U27602 (N_27602,N_26993,N_26954);
and U27603 (N_27603,N_26920,N_26856);
and U27604 (N_27604,N_26261,N_26864);
xor U27605 (N_27605,N_26411,N_26290);
nor U27606 (N_27606,N_26741,N_26826);
nor U27607 (N_27607,N_26594,N_25639);
nand U27608 (N_27608,N_26762,N_26168);
xnor U27609 (N_27609,N_25691,N_26306);
xnor U27610 (N_27610,N_26073,N_26817);
nor U27611 (N_27611,N_25632,N_26740);
or U27612 (N_27612,N_26928,N_26432);
nand U27613 (N_27613,N_26869,N_25812);
and U27614 (N_27614,N_25567,N_26176);
xnor U27615 (N_27615,N_26292,N_25534);
nand U27616 (N_27616,N_25820,N_25647);
and U27617 (N_27617,N_26123,N_25884);
xnor U27618 (N_27618,N_25961,N_26325);
nand U27619 (N_27619,N_25640,N_25806);
xor U27620 (N_27620,N_26918,N_26526);
or U27621 (N_27621,N_26095,N_26392);
and U27622 (N_27622,N_25904,N_26513);
and U27623 (N_27623,N_25550,N_25704);
or U27624 (N_27624,N_26807,N_26079);
xor U27625 (N_27625,N_26396,N_26227);
and U27626 (N_27626,N_25871,N_26371);
nand U27627 (N_27627,N_26590,N_25650);
nand U27628 (N_27628,N_25993,N_26002);
nor U27629 (N_27629,N_25605,N_26935);
and U27630 (N_27630,N_26672,N_26484);
nand U27631 (N_27631,N_26600,N_25738);
nor U27632 (N_27632,N_25670,N_26027);
and U27633 (N_27633,N_26440,N_26916);
nor U27634 (N_27634,N_26436,N_26770);
or U27635 (N_27635,N_26904,N_26997);
nand U27636 (N_27636,N_25527,N_26524);
or U27637 (N_27637,N_26813,N_25901);
nor U27638 (N_27638,N_26808,N_26703);
or U27639 (N_27639,N_26987,N_25977);
and U27640 (N_27640,N_26235,N_26190);
or U27641 (N_27641,N_26335,N_26246);
or U27642 (N_27642,N_26753,N_26088);
nand U27643 (N_27643,N_26093,N_26894);
and U27644 (N_27644,N_26963,N_26617);
nor U27645 (N_27645,N_26658,N_26998);
or U27646 (N_27646,N_26701,N_25959);
xnor U27647 (N_27647,N_25517,N_26687);
nor U27648 (N_27648,N_26835,N_26310);
nand U27649 (N_27649,N_26421,N_26099);
nand U27650 (N_27650,N_26402,N_26574);
nand U27651 (N_27651,N_25524,N_26136);
and U27652 (N_27652,N_25935,N_26787);
nand U27653 (N_27653,N_25996,N_26420);
nand U27654 (N_27654,N_26438,N_26217);
nand U27655 (N_27655,N_25571,N_26844);
xor U27656 (N_27656,N_26255,N_26446);
nor U27657 (N_27657,N_26886,N_26731);
or U27658 (N_27658,N_26046,N_25537);
or U27659 (N_27659,N_26423,N_26838);
or U27660 (N_27660,N_26907,N_26634);
nand U27661 (N_27661,N_25932,N_26724);
or U27662 (N_27662,N_25964,N_25721);
or U27663 (N_27663,N_26728,N_26323);
nor U27664 (N_27664,N_25844,N_26589);
xor U27665 (N_27665,N_26999,N_26912);
xnor U27666 (N_27666,N_26688,N_25866);
xnor U27667 (N_27667,N_26746,N_26751);
nor U27668 (N_27668,N_26354,N_26460);
nor U27669 (N_27669,N_26174,N_26405);
xor U27670 (N_27670,N_26517,N_26668);
nand U27671 (N_27671,N_25854,N_25568);
nor U27672 (N_27672,N_26567,N_26491);
nand U27673 (N_27673,N_26228,N_25828);
or U27674 (N_27674,N_26315,N_26439);
xor U27675 (N_27675,N_26972,N_25889);
nand U27676 (N_27676,N_26989,N_26264);
nand U27677 (N_27677,N_25772,N_26914);
and U27678 (N_27678,N_26337,N_26062);
xnor U27679 (N_27679,N_26349,N_25687);
nor U27680 (N_27680,N_25575,N_26779);
nand U27681 (N_27681,N_25789,N_26555);
xnor U27682 (N_27682,N_26990,N_26461);
nand U27683 (N_27683,N_26211,N_25867);
nor U27684 (N_27684,N_26924,N_26426);
and U27685 (N_27685,N_25651,N_26788);
nor U27686 (N_27686,N_26821,N_25891);
nand U27687 (N_27687,N_26718,N_26663);
and U27688 (N_27688,N_25950,N_26626);
xnor U27689 (N_27689,N_25982,N_26750);
or U27690 (N_27690,N_25970,N_26351);
nand U27691 (N_27691,N_26699,N_26025);
nand U27692 (N_27692,N_26155,N_26141);
nand U27693 (N_27693,N_26374,N_25825);
xor U27694 (N_27694,N_26789,N_25507);
nand U27695 (N_27695,N_25843,N_26781);
nor U27696 (N_27696,N_26166,N_25752);
xnor U27697 (N_27697,N_26302,N_26667);
nand U27698 (N_27698,N_25564,N_25879);
nor U27699 (N_27699,N_25954,N_26147);
nor U27700 (N_27700,N_26959,N_25598);
xnor U27701 (N_27701,N_26304,N_26008);
or U27702 (N_27702,N_25980,N_26578);
nor U27703 (N_27703,N_26378,N_26214);
nor U27704 (N_27704,N_26178,N_26311);
and U27705 (N_27705,N_25974,N_25925);
nor U27706 (N_27706,N_26743,N_26884);
or U27707 (N_27707,N_26052,N_26742);
nor U27708 (N_27708,N_26051,N_25757);
or U27709 (N_27709,N_26760,N_26901);
or U27710 (N_27710,N_26247,N_26671);
or U27711 (N_27711,N_26187,N_26528);
xnor U27712 (N_27712,N_25976,N_25608);
nor U27713 (N_27713,N_26387,N_25968);
or U27714 (N_27714,N_26927,N_26620);
nor U27715 (N_27715,N_26836,N_26475);
nor U27716 (N_27716,N_25862,N_26734);
or U27717 (N_27717,N_26801,N_25642);
or U27718 (N_27718,N_25610,N_26481);
nand U27719 (N_27719,N_25787,N_26103);
xnor U27720 (N_27720,N_26955,N_26874);
xor U27721 (N_27721,N_25790,N_25913);
xnor U27722 (N_27722,N_25877,N_26986);
nor U27723 (N_27723,N_25851,N_26259);
xor U27724 (N_27724,N_26861,N_26648);
nand U27725 (N_27725,N_26895,N_25697);
nor U27726 (N_27726,N_25509,N_26618);
or U27727 (N_27727,N_26231,N_25665);
nor U27728 (N_27728,N_26659,N_26320);
or U27729 (N_27729,N_26129,N_26271);
nor U27730 (N_27730,N_25628,N_26644);
xnor U27731 (N_27731,N_25759,N_25506);
xnor U27732 (N_27732,N_26249,N_25682);
nand U27733 (N_27733,N_26210,N_25957);
xor U27734 (N_27734,N_26795,N_25714);
or U27735 (N_27735,N_26477,N_25663);
nand U27736 (N_27736,N_26778,N_26656);
xnor U27737 (N_27737,N_26494,N_25587);
or U27738 (N_27738,N_26696,N_26357);
nand U27739 (N_27739,N_26428,N_26244);
and U27740 (N_27740,N_26182,N_26464);
nand U27741 (N_27741,N_26334,N_26135);
or U27742 (N_27742,N_25712,N_26913);
nor U27743 (N_27743,N_25818,N_25686);
or U27744 (N_27744,N_25800,N_26621);
xnor U27745 (N_27745,N_25544,N_25719);
nand U27746 (N_27746,N_26488,N_26547);
or U27747 (N_27747,N_25842,N_26089);
nand U27748 (N_27748,N_25596,N_26934);
or U27749 (N_27749,N_25693,N_26215);
nand U27750 (N_27750,N_25611,N_25795);
nand U27751 (N_27751,N_25607,N_25782);
and U27752 (N_27752,N_26686,N_26255);
nor U27753 (N_27753,N_26043,N_25595);
or U27754 (N_27754,N_26923,N_25558);
and U27755 (N_27755,N_25633,N_26409);
or U27756 (N_27756,N_26300,N_26165);
xnor U27757 (N_27757,N_26075,N_26628);
nand U27758 (N_27758,N_26259,N_26958);
or U27759 (N_27759,N_26036,N_26891);
nand U27760 (N_27760,N_26875,N_26222);
nor U27761 (N_27761,N_26836,N_26564);
and U27762 (N_27762,N_25805,N_26068);
nor U27763 (N_27763,N_26860,N_26358);
or U27764 (N_27764,N_26405,N_25919);
nor U27765 (N_27765,N_26398,N_26952);
xor U27766 (N_27766,N_26031,N_26790);
or U27767 (N_27767,N_26159,N_26991);
nor U27768 (N_27768,N_26571,N_26164);
nand U27769 (N_27769,N_26471,N_25966);
and U27770 (N_27770,N_25666,N_26458);
xnor U27771 (N_27771,N_26827,N_26610);
or U27772 (N_27772,N_26632,N_26917);
nand U27773 (N_27773,N_26446,N_26385);
nand U27774 (N_27774,N_25637,N_26304);
and U27775 (N_27775,N_26418,N_26913);
and U27776 (N_27776,N_26771,N_26276);
or U27777 (N_27777,N_26883,N_26130);
or U27778 (N_27778,N_25746,N_26242);
nand U27779 (N_27779,N_26768,N_25793);
or U27780 (N_27780,N_25862,N_26357);
or U27781 (N_27781,N_26383,N_26412);
nor U27782 (N_27782,N_25932,N_26175);
nand U27783 (N_27783,N_26702,N_26797);
nor U27784 (N_27784,N_26880,N_26399);
and U27785 (N_27785,N_25708,N_26343);
nor U27786 (N_27786,N_26986,N_25960);
xnor U27787 (N_27787,N_26827,N_26537);
nor U27788 (N_27788,N_25557,N_25576);
xor U27789 (N_27789,N_25957,N_26540);
xor U27790 (N_27790,N_25855,N_25611);
and U27791 (N_27791,N_26438,N_26732);
or U27792 (N_27792,N_26951,N_25638);
and U27793 (N_27793,N_26436,N_26184);
nor U27794 (N_27794,N_26830,N_26727);
nor U27795 (N_27795,N_26525,N_26008);
nand U27796 (N_27796,N_26835,N_26999);
and U27797 (N_27797,N_26963,N_26032);
nand U27798 (N_27798,N_25516,N_26037);
nand U27799 (N_27799,N_25959,N_25869);
nand U27800 (N_27800,N_26379,N_25841);
and U27801 (N_27801,N_26957,N_25543);
nand U27802 (N_27802,N_26880,N_26970);
nor U27803 (N_27803,N_25576,N_25721);
nand U27804 (N_27804,N_26152,N_25616);
nor U27805 (N_27805,N_25924,N_26165);
and U27806 (N_27806,N_26905,N_26531);
or U27807 (N_27807,N_25976,N_26870);
and U27808 (N_27808,N_25815,N_26610);
nor U27809 (N_27809,N_26025,N_25827);
xnor U27810 (N_27810,N_26800,N_26482);
nand U27811 (N_27811,N_26682,N_26010);
and U27812 (N_27812,N_25812,N_26541);
nor U27813 (N_27813,N_25817,N_25819);
or U27814 (N_27814,N_25630,N_25986);
xor U27815 (N_27815,N_26414,N_26980);
and U27816 (N_27816,N_26471,N_25916);
or U27817 (N_27817,N_26886,N_26807);
xor U27818 (N_27818,N_26684,N_26000);
or U27819 (N_27819,N_26631,N_26956);
and U27820 (N_27820,N_26859,N_25846);
and U27821 (N_27821,N_25971,N_26195);
nand U27822 (N_27822,N_26358,N_26379);
or U27823 (N_27823,N_25773,N_26459);
and U27824 (N_27824,N_26607,N_26309);
xnor U27825 (N_27825,N_25724,N_26596);
or U27826 (N_27826,N_26142,N_25849);
nand U27827 (N_27827,N_26849,N_26608);
or U27828 (N_27828,N_26943,N_26040);
xor U27829 (N_27829,N_26855,N_26927);
xnor U27830 (N_27830,N_26475,N_25532);
nand U27831 (N_27831,N_25885,N_26733);
or U27832 (N_27832,N_26691,N_26397);
xnor U27833 (N_27833,N_26781,N_26517);
nand U27834 (N_27834,N_26938,N_25582);
nor U27835 (N_27835,N_25938,N_25874);
nand U27836 (N_27836,N_26297,N_26747);
nor U27837 (N_27837,N_26033,N_26122);
xor U27838 (N_27838,N_26937,N_26275);
xnor U27839 (N_27839,N_26815,N_26079);
nand U27840 (N_27840,N_26544,N_25597);
or U27841 (N_27841,N_26187,N_26118);
nand U27842 (N_27842,N_26678,N_25604);
nor U27843 (N_27843,N_26832,N_26770);
xor U27844 (N_27844,N_26558,N_25976);
or U27845 (N_27845,N_25757,N_26327);
nand U27846 (N_27846,N_26996,N_26299);
xnor U27847 (N_27847,N_26813,N_26781);
nand U27848 (N_27848,N_26526,N_25669);
nor U27849 (N_27849,N_25897,N_26764);
nand U27850 (N_27850,N_25784,N_25819);
nor U27851 (N_27851,N_26423,N_26168);
nand U27852 (N_27852,N_26138,N_25516);
nor U27853 (N_27853,N_26952,N_25938);
xor U27854 (N_27854,N_25546,N_26228);
xor U27855 (N_27855,N_26381,N_26056);
or U27856 (N_27856,N_26759,N_25875);
and U27857 (N_27857,N_26721,N_26738);
nand U27858 (N_27858,N_25897,N_26834);
nand U27859 (N_27859,N_26108,N_26146);
and U27860 (N_27860,N_26901,N_26876);
nor U27861 (N_27861,N_25564,N_26681);
nor U27862 (N_27862,N_26380,N_25993);
or U27863 (N_27863,N_26386,N_25656);
nand U27864 (N_27864,N_26561,N_25945);
xor U27865 (N_27865,N_26001,N_26216);
and U27866 (N_27866,N_26287,N_25614);
nand U27867 (N_27867,N_26563,N_26853);
or U27868 (N_27868,N_26439,N_26184);
nor U27869 (N_27869,N_25507,N_25963);
xor U27870 (N_27870,N_26156,N_26685);
and U27871 (N_27871,N_25989,N_25592);
xnor U27872 (N_27872,N_26379,N_26121);
or U27873 (N_27873,N_26688,N_26534);
nand U27874 (N_27874,N_25526,N_26018);
nor U27875 (N_27875,N_26204,N_26803);
nor U27876 (N_27876,N_26546,N_26951);
or U27877 (N_27877,N_26582,N_25692);
nand U27878 (N_27878,N_26891,N_25539);
and U27879 (N_27879,N_25641,N_25628);
nand U27880 (N_27880,N_25557,N_26231);
nor U27881 (N_27881,N_26185,N_25857);
or U27882 (N_27882,N_26340,N_25703);
nor U27883 (N_27883,N_26079,N_26995);
and U27884 (N_27884,N_25851,N_26927);
or U27885 (N_27885,N_26016,N_25725);
or U27886 (N_27886,N_25998,N_26425);
and U27887 (N_27887,N_26534,N_26353);
nor U27888 (N_27888,N_25959,N_26245);
nor U27889 (N_27889,N_26241,N_25891);
and U27890 (N_27890,N_26114,N_26025);
or U27891 (N_27891,N_26440,N_25657);
xnor U27892 (N_27892,N_26040,N_26035);
xnor U27893 (N_27893,N_26762,N_25780);
xor U27894 (N_27894,N_25859,N_25951);
and U27895 (N_27895,N_26036,N_26988);
xor U27896 (N_27896,N_26376,N_26551);
nor U27897 (N_27897,N_26288,N_25523);
nor U27898 (N_27898,N_26528,N_25771);
and U27899 (N_27899,N_26420,N_25887);
and U27900 (N_27900,N_26769,N_26270);
or U27901 (N_27901,N_26158,N_26268);
nand U27902 (N_27902,N_26472,N_25686);
or U27903 (N_27903,N_25518,N_26023);
xnor U27904 (N_27904,N_25523,N_26455);
xor U27905 (N_27905,N_26142,N_26764);
nand U27906 (N_27906,N_26343,N_25832);
xnor U27907 (N_27907,N_26684,N_26483);
and U27908 (N_27908,N_26144,N_25570);
or U27909 (N_27909,N_26905,N_25627);
nand U27910 (N_27910,N_26074,N_26874);
nor U27911 (N_27911,N_26787,N_26142);
nand U27912 (N_27912,N_26272,N_25619);
or U27913 (N_27913,N_26167,N_25843);
nand U27914 (N_27914,N_26261,N_25865);
nor U27915 (N_27915,N_26934,N_26379);
nand U27916 (N_27916,N_26429,N_26017);
and U27917 (N_27917,N_26556,N_26410);
nand U27918 (N_27918,N_26543,N_25949);
and U27919 (N_27919,N_26013,N_26155);
xor U27920 (N_27920,N_26977,N_25881);
nor U27921 (N_27921,N_26859,N_26097);
xnor U27922 (N_27922,N_25882,N_26728);
and U27923 (N_27923,N_26325,N_26365);
xor U27924 (N_27924,N_25634,N_25796);
or U27925 (N_27925,N_25619,N_26091);
and U27926 (N_27926,N_26501,N_26707);
nand U27927 (N_27927,N_26278,N_26506);
nand U27928 (N_27928,N_26380,N_26226);
and U27929 (N_27929,N_25883,N_26131);
nor U27930 (N_27930,N_26964,N_26805);
or U27931 (N_27931,N_26559,N_26400);
nand U27932 (N_27932,N_26462,N_26955);
nor U27933 (N_27933,N_26759,N_26787);
nand U27934 (N_27934,N_26066,N_26014);
nand U27935 (N_27935,N_26680,N_26044);
nor U27936 (N_27936,N_25538,N_26325);
nor U27937 (N_27937,N_26645,N_26867);
or U27938 (N_27938,N_26669,N_26181);
nor U27939 (N_27939,N_26240,N_26904);
nor U27940 (N_27940,N_25867,N_26543);
or U27941 (N_27941,N_25504,N_25963);
xnor U27942 (N_27942,N_26931,N_25517);
nand U27943 (N_27943,N_26085,N_26585);
or U27944 (N_27944,N_26100,N_25644);
or U27945 (N_27945,N_26428,N_26976);
and U27946 (N_27946,N_26446,N_26640);
nor U27947 (N_27947,N_26426,N_26013);
xnor U27948 (N_27948,N_25720,N_26186);
or U27949 (N_27949,N_25500,N_25635);
and U27950 (N_27950,N_25660,N_25506);
nand U27951 (N_27951,N_26916,N_26914);
nor U27952 (N_27952,N_26398,N_26107);
or U27953 (N_27953,N_26970,N_26927);
or U27954 (N_27954,N_26881,N_25592);
and U27955 (N_27955,N_26137,N_25959);
nand U27956 (N_27956,N_25933,N_25725);
and U27957 (N_27957,N_25769,N_26572);
or U27958 (N_27958,N_26878,N_25580);
nand U27959 (N_27959,N_25788,N_26148);
xnor U27960 (N_27960,N_26587,N_26904);
nor U27961 (N_27961,N_25929,N_26185);
or U27962 (N_27962,N_26191,N_25715);
and U27963 (N_27963,N_26775,N_25761);
or U27964 (N_27964,N_26343,N_25507);
nand U27965 (N_27965,N_25805,N_26932);
and U27966 (N_27966,N_26557,N_26529);
or U27967 (N_27967,N_26246,N_25911);
nand U27968 (N_27968,N_25845,N_26540);
nor U27969 (N_27969,N_26206,N_26649);
and U27970 (N_27970,N_26581,N_25707);
nor U27971 (N_27971,N_25968,N_26248);
and U27972 (N_27972,N_26222,N_25656);
nor U27973 (N_27973,N_26937,N_25501);
nor U27974 (N_27974,N_25822,N_25754);
xor U27975 (N_27975,N_26549,N_26633);
and U27976 (N_27976,N_26435,N_26189);
nor U27977 (N_27977,N_26087,N_26985);
nand U27978 (N_27978,N_26298,N_26455);
nand U27979 (N_27979,N_25553,N_25789);
nor U27980 (N_27980,N_25953,N_26356);
nor U27981 (N_27981,N_26625,N_25694);
or U27982 (N_27982,N_26071,N_26597);
and U27983 (N_27983,N_26247,N_26609);
and U27984 (N_27984,N_25698,N_26433);
or U27985 (N_27985,N_26381,N_25991);
or U27986 (N_27986,N_25735,N_26812);
nor U27987 (N_27987,N_26466,N_25989);
or U27988 (N_27988,N_25963,N_26061);
or U27989 (N_27989,N_26435,N_26380);
nor U27990 (N_27990,N_26481,N_26424);
or U27991 (N_27991,N_25722,N_26765);
or U27992 (N_27992,N_26926,N_26150);
or U27993 (N_27993,N_26406,N_26467);
nand U27994 (N_27994,N_26246,N_26749);
nor U27995 (N_27995,N_26438,N_26460);
or U27996 (N_27996,N_26100,N_26755);
xor U27997 (N_27997,N_26700,N_25555);
nor U27998 (N_27998,N_26135,N_26677);
xnor U27999 (N_27999,N_26252,N_26760);
or U28000 (N_28000,N_25972,N_26765);
and U28001 (N_28001,N_26241,N_26188);
xor U28002 (N_28002,N_26931,N_25971);
xor U28003 (N_28003,N_26716,N_26298);
or U28004 (N_28004,N_25833,N_25992);
nor U28005 (N_28005,N_26081,N_26241);
nand U28006 (N_28006,N_25770,N_25559);
nand U28007 (N_28007,N_25817,N_25619);
or U28008 (N_28008,N_26787,N_26322);
xnor U28009 (N_28009,N_25556,N_25969);
or U28010 (N_28010,N_26269,N_25997);
xnor U28011 (N_28011,N_26493,N_26739);
or U28012 (N_28012,N_25943,N_25825);
xnor U28013 (N_28013,N_25864,N_26885);
nand U28014 (N_28014,N_25774,N_26983);
or U28015 (N_28015,N_26845,N_26532);
or U28016 (N_28016,N_25812,N_26982);
nand U28017 (N_28017,N_26582,N_26250);
nor U28018 (N_28018,N_25751,N_26118);
and U28019 (N_28019,N_25665,N_26305);
nand U28020 (N_28020,N_26777,N_25876);
nand U28021 (N_28021,N_25934,N_25718);
or U28022 (N_28022,N_25618,N_26949);
xnor U28023 (N_28023,N_26192,N_26899);
or U28024 (N_28024,N_26762,N_26530);
or U28025 (N_28025,N_26621,N_26863);
xnor U28026 (N_28026,N_26817,N_25747);
and U28027 (N_28027,N_26609,N_26719);
nor U28028 (N_28028,N_25900,N_26082);
and U28029 (N_28029,N_26394,N_26126);
xnor U28030 (N_28030,N_25674,N_25560);
and U28031 (N_28031,N_26076,N_26624);
or U28032 (N_28032,N_26374,N_26095);
nand U28033 (N_28033,N_26982,N_26537);
nand U28034 (N_28034,N_26857,N_26535);
nor U28035 (N_28035,N_25597,N_26213);
nand U28036 (N_28036,N_25945,N_25907);
nand U28037 (N_28037,N_26826,N_25972);
xor U28038 (N_28038,N_26548,N_25609);
nand U28039 (N_28039,N_26630,N_25616);
xor U28040 (N_28040,N_26349,N_25820);
or U28041 (N_28041,N_26944,N_26176);
nand U28042 (N_28042,N_26746,N_26500);
and U28043 (N_28043,N_26329,N_26722);
xnor U28044 (N_28044,N_26527,N_25998);
nor U28045 (N_28045,N_26202,N_26715);
xor U28046 (N_28046,N_26811,N_26845);
and U28047 (N_28047,N_26768,N_26484);
xor U28048 (N_28048,N_26241,N_26866);
nor U28049 (N_28049,N_26554,N_26877);
xnor U28050 (N_28050,N_26496,N_26403);
nor U28051 (N_28051,N_25735,N_25945);
nand U28052 (N_28052,N_26863,N_26149);
nand U28053 (N_28053,N_26280,N_26464);
xnor U28054 (N_28054,N_26845,N_25929);
nand U28055 (N_28055,N_26999,N_26952);
nand U28056 (N_28056,N_26238,N_25550);
and U28057 (N_28057,N_26774,N_26361);
nand U28058 (N_28058,N_26590,N_26971);
nor U28059 (N_28059,N_25954,N_26474);
or U28060 (N_28060,N_25619,N_25689);
or U28061 (N_28061,N_26505,N_25895);
nand U28062 (N_28062,N_25592,N_25569);
nand U28063 (N_28063,N_26022,N_25557);
nor U28064 (N_28064,N_25954,N_26324);
nor U28065 (N_28065,N_25940,N_25849);
nand U28066 (N_28066,N_26551,N_26563);
and U28067 (N_28067,N_26185,N_26599);
nand U28068 (N_28068,N_26641,N_25760);
xnor U28069 (N_28069,N_26518,N_26424);
or U28070 (N_28070,N_25675,N_25527);
nor U28071 (N_28071,N_26533,N_26009);
or U28072 (N_28072,N_25979,N_25706);
nand U28073 (N_28073,N_26680,N_26767);
xnor U28074 (N_28074,N_26523,N_26497);
or U28075 (N_28075,N_25593,N_26204);
and U28076 (N_28076,N_26431,N_25633);
nor U28077 (N_28077,N_26918,N_26806);
or U28078 (N_28078,N_26773,N_25887);
and U28079 (N_28079,N_25585,N_26182);
xnor U28080 (N_28080,N_26285,N_25852);
xnor U28081 (N_28081,N_26505,N_26738);
or U28082 (N_28082,N_25898,N_26566);
nor U28083 (N_28083,N_26428,N_25773);
nand U28084 (N_28084,N_26590,N_25894);
xnor U28085 (N_28085,N_26447,N_26940);
nor U28086 (N_28086,N_26590,N_25934);
nand U28087 (N_28087,N_26268,N_26362);
or U28088 (N_28088,N_25959,N_26024);
and U28089 (N_28089,N_25937,N_26879);
and U28090 (N_28090,N_25792,N_26123);
xor U28091 (N_28091,N_26758,N_26249);
nand U28092 (N_28092,N_25925,N_25747);
nand U28093 (N_28093,N_26499,N_25653);
xnor U28094 (N_28094,N_25927,N_26009);
or U28095 (N_28095,N_26188,N_25546);
or U28096 (N_28096,N_26564,N_25780);
and U28097 (N_28097,N_26013,N_26716);
or U28098 (N_28098,N_26355,N_26641);
and U28099 (N_28099,N_26294,N_26133);
and U28100 (N_28100,N_26423,N_25768);
and U28101 (N_28101,N_26888,N_26439);
nand U28102 (N_28102,N_26428,N_26594);
or U28103 (N_28103,N_25563,N_26144);
xor U28104 (N_28104,N_26038,N_26563);
xor U28105 (N_28105,N_25692,N_25852);
and U28106 (N_28106,N_26419,N_26897);
nand U28107 (N_28107,N_26040,N_25909);
or U28108 (N_28108,N_26192,N_25510);
nand U28109 (N_28109,N_26251,N_26785);
or U28110 (N_28110,N_26753,N_25670);
nand U28111 (N_28111,N_26111,N_26546);
nand U28112 (N_28112,N_26740,N_25690);
nand U28113 (N_28113,N_26949,N_25553);
or U28114 (N_28114,N_25610,N_26288);
and U28115 (N_28115,N_25744,N_26220);
xor U28116 (N_28116,N_26550,N_25888);
and U28117 (N_28117,N_26786,N_25560);
or U28118 (N_28118,N_26262,N_26729);
and U28119 (N_28119,N_26640,N_25875);
nor U28120 (N_28120,N_25709,N_26644);
or U28121 (N_28121,N_25692,N_26065);
nor U28122 (N_28122,N_25808,N_26607);
or U28123 (N_28123,N_26979,N_26499);
nand U28124 (N_28124,N_25621,N_25843);
nor U28125 (N_28125,N_26381,N_26323);
or U28126 (N_28126,N_26608,N_25790);
nand U28127 (N_28127,N_25722,N_26529);
or U28128 (N_28128,N_26365,N_26059);
xor U28129 (N_28129,N_26937,N_26237);
and U28130 (N_28130,N_26140,N_26143);
and U28131 (N_28131,N_26809,N_26520);
xor U28132 (N_28132,N_25692,N_26578);
and U28133 (N_28133,N_26664,N_26113);
and U28134 (N_28134,N_26436,N_25690);
nand U28135 (N_28135,N_26578,N_25565);
nand U28136 (N_28136,N_25858,N_26482);
nand U28137 (N_28137,N_26660,N_25729);
and U28138 (N_28138,N_25590,N_26994);
or U28139 (N_28139,N_25721,N_26404);
nand U28140 (N_28140,N_26555,N_26544);
xnor U28141 (N_28141,N_26626,N_26048);
or U28142 (N_28142,N_26811,N_26705);
and U28143 (N_28143,N_26657,N_26053);
nand U28144 (N_28144,N_26591,N_25656);
or U28145 (N_28145,N_25818,N_25977);
or U28146 (N_28146,N_26005,N_26022);
or U28147 (N_28147,N_26433,N_26461);
xnor U28148 (N_28148,N_25763,N_25968);
nand U28149 (N_28149,N_26708,N_25621);
xor U28150 (N_28150,N_26877,N_25916);
and U28151 (N_28151,N_26713,N_26215);
xnor U28152 (N_28152,N_26129,N_25614);
nor U28153 (N_28153,N_25530,N_25763);
and U28154 (N_28154,N_26224,N_25727);
xnor U28155 (N_28155,N_26225,N_26332);
xnor U28156 (N_28156,N_26064,N_26776);
and U28157 (N_28157,N_25706,N_26602);
nand U28158 (N_28158,N_26069,N_25725);
nand U28159 (N_28159,N_26906,N_26969);
nor U28160 (N_28160,N_25597,N_26194);
xnor U28161 (N_28161,N_26564,N_26136);
xnor U28162 (N_28162,N_26673,N_26654);
or U28163 (N_28163,N_26443,N_26860);
nand U28164 (N_28164,N_26986,N_25676);
nand U28165 (N_28165,N_26079,N_26764);
or U28166 (N_28166,N_26103,N_26741);
nand U28167 (N_28167,N_26500,N_26708);
nand U28168 (N_28168,N_25633,N_25993);
or U28169 (N_28169,N_25784,N_26948);
and U28170 (N_28170,N_26904,N_25640);
nand U28171 (N_28171,N_26347,N_25561);
or U28172 (N_28172,N_26454,N_26400);
nand U28173 (N_28173,N_26579,N_26078);
or U28174 (N_28174,N_25685,N_26894);
and U28175 (N_28175,N_26531,N_26273);
nand U28176 (N_28176,N_25752,N_26860);
and U28177 (N_28177,N_26828,N_26268);
and U28178 (N_28178,N_26713,N_26532);
and U28179 (N_28179,N_26648,N_25862);
and U28180 (N_28180,N_26844,N_26636);
nand U28181 (N_28181,N_26700,N_26650);
xnor U28182 (N_28182,N_26987,N_26686);
or U28183 (N_28183,N_26096,N_26920);
nor U28184 (N_28184,N_26551,N_25572);
and U28185 (N_28185,N_26605,N_25500);
xnor U28186 (N_28186,N_26845,N_25987);
nor U28187 (N_28187,N_26118,N_26255);
nor U28188 (N_28188,N_26637,N_26634);
nand U28189 (N_28189,N_26725,N_26422);
xnor U28190 (N_28190,N_26435,N_26952);
nor U28191 (N_28191,N_26856,N_26809);
or U28192 (N_28192,N_26472,N_26714);
xnor U28193 (N_28193,N_25969,N_25850);
nor U28194 (N_28194,N_26542,N_26886);
and U28195 (N_28195,N_26330,N_26890);
or U28196 (N_28196,N_26889,N_26268);
xnor U28197 (N_28197,N_26285,N_25605);
nor U28198 (N_28198,N_25982,N_26686);
xor U28199 (N_28199,N_25588,N_26686);
and U28200 (N_28200,N_26307,N_26777);
or U28201 (N_28201,N_26932,N_26304);
xnor U28202 (N_28202,N_26378,N_26353);
nand U28203 (N_28203,N_26825,N_26204);
nand U28204 (N_28204,N_26306,N_25992);
nand U28205 (N_28205,N_26193,N_26332);
xor U28206 (N_28206,N_26867,N_26008);
nor U28207 (N_28207,N_26896,N_25936);
nand U28208 (N_28208,N_25666,N_26645);
nand U28209 (N_28209,N_26660,N_26741);
nor U28210 (N_28210,N_25640,N_26467);
nor U28211 (N_28211,N_26332,N_26512);
or U28212 (N_28212,N_25645,N_26176);
or U28213 (N_28213,N_26294,N_25624);
or U28214 (N_28214,N_26990,N_26218);
nand U28215 (N_28215,N_25765,N_26642);
or U28216 (N_28216,N_26096,N_26152);
nor U28217 (N_28217,N_26668,N_26340);
nand U28218 (N_28218,N_26220,N_25916);
xnor U28219 (N_28219,N_25544,N_25702);
or U28220 (N_28220,N_26544,N_26129);
nand U28221 (N_28221,N_26902,N_26347);
or U28222 (N_28222,N_25852,N_26665);
nor U28223 (N_28223,N_26965,N_25630);
nor U28224 (N_28224,N_26212,N_26107);
nor U28225 (N_28225,N_26443,N_26712);
nor U28226 (N_28226,N_26516,N_26617);
or U28227 (N_28227,N_25530,N_25972);
or U28228 (N_28228,N_26689,N_26772);
xnor U28229 (N_28229,N_26824,N_25792);
nor U28230 (N_28230,N_26476,N_26313);
nor U28231 (N_28231,N_26777,N_26068);
and U28232 (N_28232,N_26997,N_25766);
or U28233 (N_28233,N_25639,N_26270);
xor U28234 (N_28234,N_26990,N_26565);
nand U28235 (N_28235,N_26824,N_26092);
nor U28236 (N_28236,N_26836,N_26248);
nor U28237 (N_28237,N_25573,N_26657);
nor U28238 (N_28238,N_26025,N_25713);
xnor U28239 (N_28239,N_26895,N_25866);
nand U28240 (N_28240,N_26964,N_26761);
or U28241 (N_28241,N_25883,N_26624);
xnor U28242 (N_28242,N_26548,N_26270);
nand U28243 (N_28243,N_26121,N_25590);
nand U28244 (N_28244,N_25805,N_26082);
and U28245 (N_28245,N_26363,N_26694);
and U28246 (N_28246,N_25974,N_26159);
and U28247 (N_28247,N_26091,N_26478);
and U28248 (N_28248,N_26637,N_26965);
nor U28249 (N_28249,N_26765,N_26327);
nand U28250 (N_28250,N_26108,N_25978);
nor U28251 (N_28251,N_26483,N_26416);
or U28252 (N_28252,N_25722,N_26399);
nand U28253 (N_28253,N_26225,N_26255);
and U28254 (N_28254,N_25514,N_26580);
nand U28255 (N_28255,N_26012,N_25609);
and U28256 (N_28256,N_25989,N_26881);
and U28257 (N_28257,N_26416,N_26371);
and U28258 (N_28258,N_26629,N_25776);
xnor U28259 (N_28259,N_26904,N_26395);
nand U28260 (N_28260,N_25848,N_25737);
and U28261 (N_28261,N_25860,N_26504);
nand U28262 (N_28262,N_26653,N_26619);
nand U28263 (N_28263,N_25834,N_25925);
xor U28264 (N_28264,N_26515,N_26292);
or U28265 (N_28265,N_25822,N_26067);
or U28266 (N_28266,N_26241,N_26079);
or U28267 (N_28267,N_26439,N_25627);
nor U28268 (N_28268,N_26156,N_26061);
xnor U28269 (N_28269,N_26400,N_26605);
nand U28270 (N_28270,N_25702,N_26677);
nor U28271 (N_28271,N_26686,N_26446);
nand U28272 (N_28272,N_26048,N_25997);
and U28273 (N_28273,N_26488,N_26112);
and U28274 (N_28274,N_25559,N_25632);
xor U28275 (N_28275,N_26195,N_25988);
nor U28276 (N_28276,N_26429,N_26315);
nand U28277 (N_28277,N_26757,N_26427);
xor U28278 (N_28278,N_25966,N_25565);
and U28279 (N_28279,N_25623,N_26035);
and U28280 (N_28280,N_26225,N_26004);
and U28281 (N_28281,N_26354,N_26739);
nand U28282 (N_28282,N_26616,N_26037);
or U28283 (N_28283,N_26412,N_26349);
or U28284 (N_28284,N_26420,N_26579);
nor U28285 (N_28285,N_26394,N_26371);
and U28286 (N_28286,N_26742,N_26804);
or U28287 (N_28287,N_25968,N_26349);
and U28288 (N_28288,N_25854,N_26792);
or U28289 (N_28289,N_26852,N_25755);
xor U28290 (N_28290,N_26087,N_25668);
nand U28291 (N_28291,N_25825,N_26471);
xnor U28292 (N_28292,N_26944,N_25923);
xnor U28293 (N_28293,N_26183,N_25572);
and U28294 (N_28294,N_26276,N_25639);
or U28295 (N_28295,N_25640,N_25860);
xnor U28296 (N_28296,N_26124,N_25615);
or U28297 (N_28297,N_26615,N_26369);
xor U28298 (N_28298,N_26821,N_25806);
and U28299 (N_28299,N_26990,N_26655);
xnor U28300 (N_28300,N_25660,N_26758);
xnor U28301 (N_28301,N_26703,N_26322);
or U28302 (N_28302,N_25921,N_26159);
and U28303 (N_28303,N_26459,N_26947);
or U28304 (N_28304,N_25658,N_26895);
or U28305 (N_28305,N_26878,N_26143);
or U28306 (N_28306,N_26655,N_26387);
xor U28307 (N_28307,N_25658,N_26985);
or U28308 (N_28308,N_26635,N_26853);
nand U28309 (N_28309,N_25802,N_25666);
nor U28310 (N_28310,N_26773,N_25717);
or U28311 (N_28311,N_26381,N_26098);
nor U28312 (N_28312,N_26570,N_25818);
and U28313 (N_28313,N_26880,N_25586);
nand U28314 (N_28314,N_26273,N_26893);
xnor U28315 (N_28315,N_25691,N_25538);
xor U28316 (N_28316,N_25730,N_25926);
xnor U28317 (N_28317,N_25655,N_25751);
xnor U28318 (N_28318,N_26901,N_25729);
nor U28319 (N_28319,N_26300,N_26298);
and U28320 (N_28320,N_26254,N_25976);
nand U28321 (N_28321,N_25521,N_26930);
or U28322 (N_28322,N_26581,N_26889);
or U28323 (N_28323,N_26732,N_26566);
nand U28324 (N_28324,N_26859,N_26101);
nor U28325 (N_28325,N_26048,N_26922);
nand U28326 (N_28326,N_26806,N_26881);
or U28327 (N_28327,N_26075,N_25677);
nor U28328 (N_28328,N_26260,N_26806);
nand U28329 (N_28329,N_26241,N_25743);
nor U28330 (N_28330,N_26621,N_25633);
and U28331 (N_28331,N_26152,N_26409);
or U28332 (N_28332,N_25988,N_26840);
xor U28333 (N_28333,N_26402,N_26620);
nand U28334 (N_28334,N_25933,N_26497);
nor U28335 (N_28335,N_26906,N_26346);
nor U28336 (N_28336,N_26299,N_26509);
nand U28337 (N_28337,N_26357,N_26811);
nor U28338 (N_28338,N_25855,N_26185);
nor U28339 (N_28339,N_26019,N_26667);
nor U28340 (N_28340,N_25680,N_25659);
nor U28341 (N_28341,N_25585,N_26814);
nor U28342 (N_28342,N_26495,N_26744);
and U28343 (N_28343,N_26685,N_25842);
or U28344 (N_28344,N_25824,N_26426);
or U28345 (N_28345,N_26723,N_25675);
nand U28346 (N_28346,N_26792,N_26234);
nand U28347 (N_28347,N_26470,N_26907);
nor U28348 (N_28348,N_26956,N_25564);
nor U28349 (N_28349,N_26228,N_25924);
nor U28350 (N_28350,N_25682,N_26449);
or U28351 (N_28351,N_26054,N_25974);
nor U28352 (N_28352,N_26877,N_25986);
and U28353 (N_28353,N_26492,N_26735);
xor U28354 (N_28354,N_26770,N_26743);
xnor U28355 (N_28355,N_25754,N_25690);
or U28356 (N_28356,N_26882,N_26513);
or U28357 (N_28357,N_25755,N_26854);
or U28358 (N_28358,N_25770,N_25614);
and U28359 (N_28359,N_26074,N_25919);
xnor U28360 (N_28360,N_26221,N_26582);
nand U28361 (N_28361,N_26924,N_26918);
nor U28362 (N_28362,N_25536,N_26627);
and U28363 (N_28363,N_25795,N_25520);
xor U28364 (N_28364,N_26838,N_26363);
and U28365 (N_28365,N_26874,N_25879);
or U28366 (N_28366,N_26006,N_25543);
or U28367 (N_28367,N_25940,N_26603);
and U28368 (N_28368,N_25790,N_25836);
or U28369 (N_28369,N_26255,N_25950);
nor U28370 (N_28370,N_26568,N_25801);
xnor U28371 (N_28371,N_26371,N_26081);
nor U28372 (N_28372,N_26697,N_25814);
nor U28373 (N_28373,N_26807,N_26831);
xnor U28374 (N_28374,N_25822,N_26673);
nor U28375 (N_28375,N_25824,N_26760);
xnor U28376 (N_28376,N_26801,N_26474);
or U28377 (N_28377,N_26081,N_26874);
or U28378 (N_28378,N_25921,N_25789);
nand U28379 (N_28379,N_26771,N_26425);
or U28380 (N_28380,N_25502,N_25929);
nor U28381 (N_28381,N_26408,N_25758);
or U28382 (N_28382,N_26207,N_26224);
and U28383 (N_28383,N_25936,N_26388);
nor U28384 (N_28384,N_26280,N_26273);
nor U28385 (N_28385,N_26482,N_26246);
nor U28386 (N_28386,N_26271,N_25661);
nor U28387 (N_28387,N_26233,N_26097);
nor U28388 (N_28388,N_25688,N_26285);
and U28389 (N_28389,N_26268,N_26038);
xnor U28390 (N_28390,N_26834,N_25966);
and U28391 (N_28391,N_26082,N_25906);
xnor U28392 (N_28392,N_26260,N_25816);
or U28393 (N_28393,N_25841,N_26540);
and U28394 (N_28394,N_26334,N_26855);
xnor U28395 (N_28395,N_25607,N_26846);
or U28396 (N_28396,N_26962,N_26482);
nor U28397 (N_28397,N_26295,N_26829);
nor U28398 (N_28398,N_26974,N_25785);
and U28399 (N_28399,N_26922,N_26705);
and U28400 (N_28400,N_25890,N_26952);
or U28401 (N_28401,N_25669,N_26632);
and U28402 (N_28402,N_25890,N_26436);
nor U28403 (N_28403,N_25712,N_26867);
nand U28404 (N_28404,N_26872,N_26666);
nand U28405 (N_28405,N_26234,N_25859);
nand U28406 (N_28406,N_26515,N_26618);
nand U28407 (N_28407,N_25997,N_25957);
or U28408 (N_28408,N_25707,N_25978);
nand U28409 (N_28409,N_25883,N_26065);
or U28410 (N_28410,N_26733,N_25998);
and U28411 (N_28411,N_25998,N_26624);
and U28412 (N_28412,N_25727,N_26181);
or U28413 (N_28413,N_26443,N_25687);
xnor U28414 (N_28414,N_26602,N_26124);
xnor U28415 (N_28415,N_26297,N_26979);
and U28416 (N_28416,N_25760,N_26811);
xnor U28417 (N_28417,N_26463,N_26343);
or U28418 (N_28418,N_25671,N_25554);
and U28419 (N_28419,N_26851,N_25569);
nand U28420 (N_28420,N_26588,N_26720);
xnor U28421 (N_28421,N_25936,N_26680);
nor U28422 (N_28422,N_26299,N_26279);
nand U28423 (N_28423,N_25517,N_25635);
nor U28424 (N_28424,N_26390,N_26177);
nor U28425 (N_28425,N_26922,N_26853);
and U28426 (N_28426,N_26634,N_26991);
nand U28427 (N_28427,N_26948,N_25923);
and U28428 (N_28428,N_25820,N_26618);
or U28429 (N_28429,N_25837,N_25532);
nand U28430 (N_28430,N_26210,N_26889);
xor U28431 (N_28431,N_26226,N_25758);
and U28432 (N_28432,N_26149,N_26134);
xnor U28433 (N_28433,N_26055,N_26245);
nor U28434 (N_28434,N_26969,N_26137);
and U28435 (N_28435,N_25897,N_25511);
nand U28436 (N_28436,N_25717,N_26827);
nor U28437 (N_28437,N_26129,N_25779);
xnor U28438 (N_28438,N_26155,N_25922);
and U28439 (N_28439,N_26673,N_26676);
or U28440 (N_28440,N_26032,N_25637);
and U28441 (N_28441,N_26383,N_26212);
xor U28442 (N_28442,N_26721,N_26238);
and U28443 (N_28443,N_25904,N_26229);
and U28444 (N_28444,N_26843,N_25978);
xnor U28445 (N_28445,N_25999,N_26754);
or U28446 (N_28446,N_25928,N_25593);
or U28447 (N_28447,N_25929,N_26069);
nand U28448 (N_28448,N_26057,N_26993);
or U28449 (N_28449,N_26109,N_26410);
and U28450 (N_28450,N_26901,N_26106);
nor U28451 (N_28451,N_26017,N_26836);
xnor U28452 (N_28452,N_26166,N_26834);
nor U28453 (N_28453,N_26475,N_26739);
or U28454 (N_28454,N_26600,N_26189);
nor U28455 (N_28455,N_26552,N_26522);
xnor U28456 (N_28456,N_26825,N_26081);
nand U28457 (N_28457,N_26481,N_25726);
xor U28458 (N_28458,N_26356,N_25800);
or U28459 (N_28459,N_25526,N_25631);
xnor U28460 (N_28460,N_25961,N_25867);
and U28461 (N_28461,N_26818,N_25702);
or U28462 (N_28462,N_26122,N_26548);
and U28463 (N_28463,N_25844,N_26873);
and U28464 (N_28464,N_26202,N_25627);
and U28465 (N_28465,N_25585,N_26239);
or U28466 (N_28466,N_25513,N_25692);
or U28467 (N_28467,N_26988,N_25521);
nand U28468 (N_28468,N_25624,N_25874);
nand U28469 (N_28469,N_26413,N_26959);
xnor U28470 (N_28470,N_26446,N_25882);
or U28471 (N_28471,N_26232,N_26929);
and U28472 (N_28472,N_26451,N_25658);
xor U28473 (N_28473,N_25798,N_26204);
xnor U28474 (N_28474,N_26615,N_26743);
xnor U28475 (N_28475,N_26380,N_26445);
nand U28476 (N_28476,N_26868,N_26201);
nand U28477 (N_28477,N_25569,N_26988);
xnor U28478 (N_28478,N_25902,N_26364);
or U28479 (N_28479,N_26109,N_25541);
nor U28480 (N_28480,N_26553,N_25678);
and U28481 (N_28481,N_26763,N_25604);
and U28482 (N_28482,N_26348,N_25797);
nor U28483 (N_28483,N_25955,N_26452);
and U28484 (N_28484,N_26327,N_26998);
and U28485 (N_28485,N_25745,N_26538);
xnor U28486 (N_28486,N_25665,N_26385);
xor U28487 (N_28487,N_26481,N_26566);
nand U28488 (N_28488,N_25873,N_26876);
nor U28489 (N_28489,N_25659,N_25932);
and U28490 (N_28490,N_26801,N_25976);
nand U28491 (N_28491,N_25897,N_25578);
nand U28492 (N_28492,N_26816,N_26041);
xor U28493 (N_28493,N_26449,N_26405);
and U28494 (N_28494,N_26997,N_26524);
xnor U28495 (N_28495,N_25687,N_26555);
nand U28496 (N_28496,N_26406,N_26681);
and U28497 (N_28497,N_25654,N_26460);
nor U28498 (N_28498,N_26338,N_25720);
xor U28499 (N_28499,N_26017,N_26559);
nand U28500 (N_28500,N_28421,N_28007);
nand U28501 (N_28501,N_27852,N_28152);
nor U28502 (N_28502,N_28077,N_28447);
or U28503 (N_28503,N_27468,N_27223);
nand U28504 (N_28504,N_27447,N_28094);
nand U28505 (N_28505,N_28497,N_27199);
nand U28506 (N_28506,N_28203,N_27779);
nand U28507 (N_28507,N_27641,N_28170);
and U28508 (N_28508,N_28245,N_27542);
nor U28509 (N_28509,N_27697,N_27178);
or U28510 (N_28510,N_27898,N_27407);
and U28511 (N_28511,N_27343,N_27258);
or U28512 (N_28512,N_27410,N_27083);
and U28513 (N_28513,N_27392,N_27785);
xnor U28514 (N_28514,N_28195,N_27008);
or U28515 (N_28515,N_27401,N_28361);
xnor U28516 (N_28516,N_27572,N_27602);
and U28517 (N_28517,N_27707,N_27648);
xnor U28518 (N_28518,N_28256,N_28453);
nor U28519 (N_28519,N_27453,N_27679);
or U28520 (N_28520,N_28327,N_27222);
xnor U28521 (N_28521,N_27563,N_27022);
and U28522 (N_28522,N_27352,N_27505);
nor U28523 (N_28523,N_27794,N_27026);
xnor U28524 (N_28524,N_27763,N_27769);
nor U28525 (N_28525,N_27093,N_27620);
nor U28526 (N_28526,N_27860,N_27825);
nand U28527 (N_28527,N_27100,N_28084);
xor U28528 (N_28528,N_28221,N_28124);
or U28529 (N_28529,N_28012,N_27454);
nand U28530 (N_28530,N_27206,N_28038);
xor U28531 (N_28531,N_28458,N_27722);
xor U28532 (N_28532,N_27378,N_28248);
and U28533 (N_28533,N_27612,N_27025);
and U28534 (N_28534,N_28252,N_27465);
or U28535 (N_28535,N_28401,N_27265);
and U28536 (N_28536,N_28039,N_28489);
nor U28537 (N_28537,N_27740,N_27293);
and U28538 (N_28538,N_28455,N_28352);
nor U28539 (N_28539,N_28157,N_28377);
nand U28540 (N_28540,N_27932,N_27901);
or U28541 (N_28541,N_27342,N_27607);
nor U28542 (N_28542,N_27067,N_27221);
xnor U28543 (N_28543,N_27528,N_28459);
nand U28544 (N_28544,N_28285,N_27382);
xor U28545 (N_28545,N_28277,N_28190);
nor U28546 (N_28546,N_27765,N_28389);
xnor U28547 (N_28547,N_28136,N_28499);
nand U28548 (N_28548,N_28165,N_27208);
or U28549 (N_28549,N_28130,N_28063);
xnor U28550 (N_28550,N_28200,N_27942);
and U28551 (N_28551,N_28046,N_28324);
xor U28552 (N_28552,N_28099,N_28270);
and U28553 (N_28553,N_28049,N_28028);
nand U28554 (N_28554,N_27294,N_27623);
and U28555 (N_28555,N_28359,N_28255);
nand U28556 (N_28556,N_27063,N_27192);
nand U28557 (N_28557,N_27667,N_27492);
nand U28558 (N_28558,N_27303,N_27347);
nand U28559 (N_28559,N_28120,N_27739);
nor U28560 (N_28560,N_27913,N_27155);
and U28561 (N_28561,N_27263,N_27460);
nor U28562 (N_28562,N_27012,N_27538);
xor U28563 (N_28563,N_27649,N_27243);
nor U28564 (N_28564,N_28131,N_28280);
nand U28565 (N_28565,N_27500,N_28238);
xnor U28566 (N_28566,N_27949,N_27712);
xor U28567 (N_28567,N_27481,N_27182);
xnor U28568 (N_28568,N_28479,N_27130);
nor U28569 (N_28569,N_27409,N_27872);
nand U28570 (N_28570,N_27080,N_27736);
or U28571 (N_28571,N_28316,N_28054);
nor U28572 (N_28572,N_27502,N_28303);
and U28573 (N_28573,N_27205,N_27828);
or U28574 (N_28574,N_27190,N_28178);
or U28575 (N_28575,N_28350,N_28486);
nand U28576 (N_28576,N_28430,N_28261);
nand U28577 (N_28577,N_28317,N_27189);
and U28578 (N_28578,N_28269,N_27473);
nand U28579 (N_28579,N_27692,N_28388);
and U28580 (N_28580,N_27362,N_27903);
nand U28581 (N_28581,N_27630,N_27742);
and U28582 (N_28582,N_27506,N_27933);
xor U28583 (N_28583,N_27940,N_27833);
xor U28584 (N_28584,N_27319,N_28167);
and U28585 (N_28585,N_27467,N_27116);
and U28586 (N_28586,N_27137,N_27590);
or U28587 (N_28587,N_27445,N_27286);
nor U28588 (N_28588,N_27776,N_27651);
or U28589 (N_28589,N_27511,N_27879);
nor U28590 (N_28590,N_27694,N_28073);
xnor U28591 (N_28591,N_27826,N_28408);
or U28592 (N_28592,N_27513,N_27162);
and U28593 (N_28593,N_27832,N_28246);
nand U28594 (N_28594,N_28493,N_28475);
xor U28595 (N_28595,N_27323,N_27062);
nor U28596 (N_28596,N_27811,N_27863);
or U28597 (N_28597,N_27016,N_27536);
and U28598 (N_28598,N_28417,N_28380);
xnor U28599 (N_28599,N_28158,N_27868);
and U28600 (N_28600,N_27298,N_27227);
xor U28601 (N_28601,N_28217,N_27814);
nor U28602 (N_28602,N_27708,N_27615);
and U28603 (N_28603,N_28125,N_27916);
xor U28604 (N_28604,N_27504,N_27474);
nor U28605 (N_28605,N_27802,N_27895);
and U28606 (N_28606,N_27246,N_27803);
nor U28607 (N_28607,N_28212,N_27558);
or U28608 (N_28608,N_27232,N_27226);
or U28609 (N_28609,N_28266,N_27735);
xnor U28610 (N_28610,N_27021,N_28045);
xnor U28611 (N_28611,N_27011,N_28069);
nand U28612 (N_28612,N_27480,N_27818);
or U28613 (N_28613,N_27254,N_27234);
xnor U28614 (N_28614,N_27730,N_27124);
nor U28615 (N_28615,N_28101,N_27096);
nand U28616 (N_28616,N_28473,N_27775);
or U28617 (N_28617,N_28498,N_27476);
xnor U28618 (N_28618,N_28095,N_27095);
or U28619 (N_28619,N_28376,N_27876);
or U28620 (N_28620,N_27867,N_27924);
nor U28621 (N_28621,N_28367,N_27645);
nor U28622 (N_28622,N_27132,N_28188);
nor U28623 (N_28623,N_27691,N_28406);
nor U28624 (N_28624,N_27372,N_28199);
nor U28625 (N_28625,N_28399,N_27585);
nand U28626 (N_28626,N_27703,N_28283);
xnor U28627 (N_28627,N_27812,N_27908);
nand U28628 (N_28628,N_27220,N_27522);
and U28629 (N_28629,N_27201,N_27902);
nor U28630 (N_28630,N_27592,N_27282);
and U28631 (N_28631,N_28305,N_28434);
nand U28632 (N_28632,N_27526,N_27040);
or U28633 (N_28633,N_28348,N_28098);
and U28634 (N_28634,N_27161,N_28278);
and U28635 (N_28635,N_27449,N_27517);
and U28636 (N_28636,N_27984,N_27520);
and U28637 (N_28637,N_27020,N_27972);
and U28638 (N_28638,N_27399,N_27823);
xor U28639 (N_28639,N_27798,N_28088);
nor U28640 (N_28640,N_28308,N_27665);
xnor U28641 (N_28641,N_27397,N_28228);
nor U28642 (N_28642,N_28233,N_27793);
nand U28643 (N_28643,N_27421,N_27570);
and U28644 (N_28644,N_28263,N_27405);
xor U28645 (N_28645,N_27479,N_27927);
or U28646 (N_28646,N_27121,N_27324);
and U28647 (N_28647,N_28426,N_27287);
nor U28648 (N_28648,N_28171,N_27035);
nor U28649 (N_28649,N_27332,N_27256);
nand U28650 (N_28650,N_28139,N_27678);
nand U28651 (N_28651,N_27531,N_28370);
nor U28652 (N_28652,N_28240,N_27569);
nand U28653 (N_28653,N_27849,N_28145);
or U28654 (N_28654,N_27819,N_27325);
and U28655 (N_28655,N_27231,N_28214);
nand U28656 (N_28656,N_27261,N_28378);
xor U28657 (N_28657,N_27726,N_27669);
and U28658 (N_28658,N_27809,N_28379);
nor U28659 (N_28659,N_27230,N_27269);
xnor U28660 (N_28660,N_28336,N_27448);
and U28661 (N_28661,N_27180,N_27524);
or U28662 (N_28662,N_27787,N_27052);
nor U28663 (N_28663,N_27990,N_28047);
nor U28664 (N_28664,N_27112,N_27183);
nor U28665 (N_28665,N_28396,N_27334);
or U28666 (N_28666,N_27551,N_27338);
or U28667 (N_28667,N_28268,N_27488);
or U28668 (N_28668,N_27545,N_28474);
and U28669 (N_28669,N_27611,N_27001);
xnor U28670 (N_28670,N_28340,N_27235);
and U28671 (N_28671,N_28106,N_27154);
or U28672 (N_28672,N_27875,N_28064);
nor U28673 (N_28673,N_28452,N_27946);
nand U28674 (N_28674,N_27519,N_27601);
nand U28675 (N_28675,N_28097,N_27786);
xor U28676 (N_28676,N_27143,N_27591);
nand U28677 (N_28677,N_28351,N_27416);
xor U28678 (N_28678,N_27682,N_27166);
nor U28679 (N_28679,N_27967,N_27631);
nand U28680 (N_28680,N_27218,N_27829);
or U28681 (N_28681,N_27037,N_28232);
nand U28682 (N_28682,N_28250,N_27835);
and U28683 (N_28683,N_27259,N_28224);
xor U28684 (N_28684,N_28437,N_27851);
or U28685 (N_28685,N_27584,N_27482);
xnor U28686 (N_28686,N_28074,N_27887);
nand U28687 (N_28687,N_27613,N_27894);
nor U28688 (N_28688,N_27370,N_27075);
and U28689 (N_28689,N_27329,N_27676);
nor U28690 (N_28690,N_28031,N_27573);
nor U28691 (N_28691,N_27574,N_27437);
xor U28692 (N_28692,N_27483,N_27024);
nand U28693 (N_28693,N_28247,N_28309);
or U28694 (N_28694,N_27518,N_27109);
and U28695 (N_28695,N_27310,N_27748);
or U28696 (N_28696,N_27088,N_27800);
nor U28697 (N_28697,N_27501,N_27097);
nor U28698 (N_28698,N_27577,N_28290);
and U28699 (N_28699,N_28024,N_28287);
xnor U28700 (N_28700,N_28339,N_27149);
nor U28701 (N_28701,N_27698,N_27306);
xnor U28702 (N_28702,N_28194,N_27113);
or U28703 (N_28703,N_28107,N_27374);
and U28704 (N_28704,N_27530,N_27050);
xnor U28705 (N_28705,N_27733,N_28008);
xnor U28706 (N_28706,N_28411,N_28119);
or U28707 (N_28707,N_28148,N_27215);
and U28708 (N_28708,N_27301,N_27181);
nand U28709 (N_28709,N_28410,N_27440);
or U28710 (N_28710,N_28092,N_27163);
nand U28711 (N_28711,N_28419,N_27159);
or U28712 (N_28712,N_27595,N_28236);
nor U28713 (N_28713,N_27042,N_27821);
nand U28714 (N_28714,N_27945,N_28333);
nor U28715 (N_28715,N_28402,N_28225);
nand U28716 (N_28716,N_28456,N_28164);
or U28717 (N_28717,N_27516,N_27644);
xnor U28718 (N_28718,N_28035,N_27827);
nor U28719 (N_28719,N_27015,N_27552);
nor U28720 (N_28720,N_27187,N_27690);
nand U28721 (N_28721,N_28496,N_28442);
or U28722 (N_28722,N_27890,N_27627);
and U28723 (N_28723,N_28113,N_27571);
nand U28724 (N_28724,N_28363,N_27795);
xor U28725 (N_28725,N_27652,N_27813);
or U28726 (N_28726,N_27788,N_28320);
xnor U28727 (N_28727,N_27033,N_28307);
or U28728 (N_28728,N_27317,N_27139);
xor U28729 (N_28729,N_27906,N_27443);
nor U28730 (N_28730,N_27731,N_27559);
xnor U28731 (N_28731,N_28090,N_27418);
nor U28732 (N_28732,N_27843,N_27593);
nor U28733 (N_28733,N_28267,N_27308);
xor U28734 (N_28734,N_28160,N_28487);
nand U28735 (N_28735,N_28279,N_27245);
nor U28736 (N_28736,N_27262,N_27878);
xor U28737 (N_28737,N_28142,N_27348);
nand U28738 (N_28738,N_28443,N_27715);
nor U28739 (N_28739,N_27486,N_28414);
nand U28740 (N_28740,N_27944,N_27955);
and U28741 (N_28741,N_27820,N_27283);
and U28742 (N_28742,N_27081,N_28286);
and U28743 (N_28743,N_27117,N_28302);
nand U28744 (N_28744,N_28126,N_27700);
and U28745 (N_28745,N_27302,N_27133);
or U28746 (N_28746,N_28323,N_27060);
nor U28747 (N_28747,N_28067,N_28226);
nand U28748 (N_28748,N_28362,N_27704);
nor U28749 (N_28749,N_27764,N_27998);
nor U28750 (N_28750,N_27989,N_27791);
xor U28751 (N_28751,N_27281,N_28050);
or U28752 (N_28752,N_28193,N_27251);
and U28753 (N_28753,N_27300,N_27351);
xor U28754 (N_28754,N_27533,N_27606);
nor U28755 (N_28755,N_27805,N_27197);
nand U28756 (N_28756,N_27555,N_27781);
and U28757 (N_28757,N_27158,N_27871);
xor U28758 (N_28758,N_27434,N_28253);
nor U28759 (N_28759,N_27078,N_27084);
xnor U28760 (N_28760,N_28464,N_28326);
xor U28761 (N_28761,N_28281,N_27295);
xor U28762 (N_28762,N_28040,N_28328);
and U28763 (N_28763,N_27017,N_28304);
xnor U28764 (N_28764,N_27253,N_28470);
and U28765 (N_28765,N_28017,N_28072);
or U28766 (N_28766,N_27054,N_27224);
xnor U28767 (N_28767,N_28070,N_28030);
nor U28768 (N_28768,N_27959,N_27387);
xor U28769 (N_28769,N_27801,N_27321);
nand U28770 (N_28770,N_28461,N_27846);
nor U28771 (N_28771,N_28284,N_28445);
and U28772 (N_28772,N_28349,N_27364);
nor U28773 (N_28773,N_28183,N_28000);
and U28774 (N_28774,N_27762,N_27587);
or U28775 (N_28775,N_28471,N_27036);
nand U28776 (N_28776,N_27755,N_27431);
or U28777 (N_28777,N_27966,N_27371);
nand U28778 (N_28778,N_28089,N_27249);
or U28779 (N_28779,N_28211,N_27562);
or U28780 (N_28780,N_27009,N_27091);
nor U28781 (N_28781,N_27633,N_27315);
nand U28782 (N_28782,N_27101,N_27424);
xnor U28783 (N_28783,N_28483,N_28229);
nor U28784 (N_28784,N_27489,N_27244);
xor U28785 (N_28785,N_27128,N_28325);
nand U28786 (N_28786,N_27209,N_27535);
or U28787 (N_28787,N_28372,N_27977);
nor U28788 (N_28788,N_27041,N_28365);
nand U28789 (N_28789,N_28026,N_28260);
or U28790 (N_28790,N_27272,N_28395);
nand U28791 (N_28791,N_27344,N_27389);
or U28792 (N_28792,N_27156,N_28301);
xor U28793 (N_28793,N_27670,N_27757);
and U28794 (N_28794,N_27750,N_28086);
xor U28795 (N_28795,N_28288,N_27919);
nor U28796 (N_28796,N_27929,N_28173);
xor U28797 (N_28797,N_27999,N_27507);
xor U28798 (N_28798,N_27186,N_28132);
or U28799 (N_28799,N_28344,N_27127);
nand U28800 (N_28800,N_27268,N_28181);
xor U28801 (N_28801,N_28207,N_28314);
nor U28802 (N_28802,N_28150,N_27953);
or U28803 (N_28803,N_27292,N_27403);
xnor U28804 (N_28804,N_27194,N_27285);
nand U28805 (N_28805,N_27576,N_27568);
nand U28806 (N_28806,N_27636,N_27979);
and U28807 (N_28807,N_28293,N_28368);
nor U28808 (N_28808,N_27674,N_28202);
nor U28809 (N_28809,N_27337,N_27836);
xor U28810 (N_28810,N_27188,N_27019);
or U28811 (N_28811,N_27807,N_28011);
or U28812 (N_28812,N_28206,N_27006);
or U28813 (N_28813,N_27521,N_27353);
nor U28814 (N_28814,N_28387,N_27493);
and U28815 (N_28815,N_28213,N_28121);
nand U28816 (N_28816,N_27861,N_28257);
nand U28817 (N_28817,N_28300,N_28400);
nor U28818 (N_28818,N_27043,N_28179);
nor U28819 (N_28819,N_27655,N_27614);
nor U28820 (N_28820,N_27824,N_27915);
nand U28821 (N_28821,N_27381,N_28373);
nand U28822 (N_28822,N_27886,N_27543);
xnor U28823 (N_28823,N_27564,N_28205);
nor U28824 (N_28824,N_28112,N_28296);
xnor U28825 (N_28825,N_27525,N_28085);
or U28826 (N_28826,N_28490,N_27164);
nand U28827 (N_28827,N_28423,N_28264);
nor U28828 (N_28828,N_28066,N_27610);
xor U28829 (N_28829,N_27425,N_27055);
and U28830 (N_28830,N_27892,N_28025);
xnor U28831 (N_28831,N_28422,N_27257);
nand U28832 (N_28832,N_27074,N_27202);
nor U28833 (N_28833,N_28115,N_28295);
nand U28834 (N_28834,N_28358,N_28436);
or U28835 (N_28835,N_27135,N_27609);
or U28836 (N_28836,N_28058,N_27115);
xnor U28837 (N_28837,N_27904,N_28243);
or U28838 (N_28838,N_27047,N_27938);
or U28839 (N_28839,N_28018,N_27756);
or U28840 (N_28840,N_27219,N_27312);
or U28841 (N_28841,N_28154,N_27335);
or U28842 (N_28842,N_27920,N_27331);
and U28843 (N_28843,N_27626,N_27656);
and U28844 (N_28844,N_27588,N_28111);
nor U28845 (N_28845,N_27893,N_27647);
nor U28846 (N_28846,N_27107,N_27575);
nor U28847 (N_28847,N_28397,N_28016);
or U28848 (N_28848,N_28371,N_27921);
nand U28849 (N_28849,N_27304,N_27491);
and U28850 (N_28850,N_27496,N_27777);
xor U28851 (N_28851,N_28209,N_27854);
nor U28852 (N_28852,N_27841,N_27071);
nand U28853 (N_28853,N_27138,N_27087);
or U28854 (N_28854,N_28201,N_27724);
or U28855 (N_28855,N_27316,N_27737);
and U28856 (N_28856,N_27267,N_27023);
xnor U28857 (N_28857,N_28390,N_28078);
or U28858 (N_28858,N_27086,N_27677);
xnor U28859 (N_28859,N_27956,N_27470);
nand U28860 (N_28860,N_27553,N_28166);
nor U28861 (N_28861,N_28075,N_28032);
nor U28862 (N_28862,N_27650,N_28187);
xor U28863 (N_28863,N_28055,N_28392);
xor U28864 (N_28864,N_28335,N_27550);
or U28865 (N_28865,N_27108,N_28109);
and U28866 (N_28866,N_27617,N_28042);
nand U28867 (N_28867,N_27239,N_27848);
nor U28868 (N_28868,N_28022,N_28198);
xor U28869 (N_28869,N_28374,N_27621);
nor U28870 (N_28870,N_27983,N_27356);
nor U28871 (N_28871,N_27689,N_27427);
nor U28872 (N_28872,N_27605,N_28439);
nand U28873 (N_28873,N_28494,N_27658);
nand U28874 (N_28874,N_27436,N_27110);
nor U28875 (N_28875,N_28116,N_28093);
xnor U28876 (N_28876,N_27069,N_28440);
and U28877 (N_28877,N_27770,N_28292);
or U28878 (N_28878,N_27705,N_28415);
and U28879 (N_28879,N_28080,N_27973);
nand U28880 (N_28880,N_28197,N_27049);
or U28881 (N_28881,N_28386,N_28182);
nor U28882 (N_28882,N_27873,N_27532);
nand U28883 (N_28883,N_27394,N_27547);
or U28884 (N_28884,N_27745,N_28061);
xor U28885 (N_28885,N_28208,N_28424);
xor U28886 (N_28886,N_27299,N_27907);
xnor U28887 (N_28887,N_28021,N_27544);
xor U28888 (N_28888,N_27327,N_27179);
and U28889 (N_28889,N_27625,N_27284);
xor U28890 (N_28890,N_28403,N_27792);
xor U28891 (N_28891,N_27277,N_27497);
or U28892 (N_28892,N_28027,N_28052);
xor U28893 (N_28893,N_28343,N_28172);
and U28894 (N_28894,N_27373,N_27589);
nand U28895 (N_28895,N_28068,N_27982);
xnor U28896 (N_28896,N_28407,N_28416);
nor U28897 (N_28897,N_27950,N_27064);
nand U28898 (N_28898,N_27126,N_27475);
xor U28899 (N_28899,N_28156,N_27350);
nor U28900 (N_28900,N_27296,N_28015);
nand U28901 (N_28901,N_27732,N_27478);
nand U28902 (N_28902,N_27171,N_27495);
xnor U28903 (N_28903,N_27808,N_27540);
and U28904 (N_28904,N_28176,N_27305);
nand U28905 (N_28905,N_27217,N_28135);
and U28906 (N_28906,N_27952,N_27581);
nand U28907 (N_28907,N_27203,N_27672);
nor U28908 (N_28908,N_27815,N_27870);
nor U28909 (N_28909,N_27599,N_27375);
xnor U28910 (N_28910,N_28029,N_27681);
nor U28911 (N_28911,N_28180,N_27406);
xor U28912 (N_28912,N_28044,N_27992);
xor U28913 (N_28913,N_27830,N_27376);
nand U28914 (N_28914,N_27790,N_27388);
or U28915 (N_28915,N_27600,N_27198);
nor U28916 (N_28916,N_27214,N_27313);
xnor U28917 (N_28917,N_28128,N_27092);
nor U28918 (N_28918,N_27673,N_27419);
nand U28919 (N_28919,N_27297,N_28251);
nand U28920 (N_28920,N_27918,N_27508);
and U28921 (N_28921,N_27582,N_27141);
nand U28922 (N_28922,N_27877,N_27954);
nor U28923 (N_28923,N_27837,N_27354);
nor U28924 (N_28924,N_28353,N_28398);
nand U28925 (N_28925,N_27002,N_27099);
or U28926 (N_28926,N_27789,N_27856);
nor U28927 (N_28927,N_27193,N_28241);
xor U28928 (N_28928,N_28420,N_28048);
and U28929 (N_28929,N_28169,N_27628);
and U28930 (N_28930,N_27216,N_27509);
or U28931 (N_28931,N_28451,N_27196);
nand U28932 (N_28932,N_28043,N_27291);
nor U28933 (N_28933,N_28282,N_28299);
and U28934 (N_28934,N_27146,N_28298);
xnor U28935 (N_28935,N_27048,N_27646);
or U28936 (N_28936,N_28001,N_27958);
nor U28937 (N_28937,N_27774,N_27204);
nor U28938 (N_28938,N_27874,N_28364);
xnor U28939 (N_28939,N_27900,N_28330);
nand U28940 (N_28940,N_27385,N_27438);
xnor U28941 (N_28941,N_27452,N_27784);
xnor U28942 (N_28942,N_28062,N_28056);
xor U28943 (N_28943,N_27464,N_27840);
nand U28944 (N_28944,N_27991,N_28272);
or U28945 (N_28945,N_27663,N_27345);
xnor U28946 (N_28946,N_28219,N_28341);
xnor U28947 (N_28947,N_28168,N_27122);
and U28948 (N_28948,N_27653,N_28432);
xnor U28949 (N_28949,N_28249,N_27537);
xnor U28950 (N_28950,N_27384,N_27152);
xor U28951 (N_28951,N_27914,N_28191);
or U28952 (N_28952,N_27939,N_27273);
xor U28953 (N_28953,N_27328,N_27118);
xnor U28954 (N_28954,N_28467,N_28412);
and U28955 (N_28955,N_27666,N_27469);
nand U28956 (N_28956,N_27668,N_27675);
and U28957 (N_28957,N_28104,N_27367);
nor U28958 (N_28958,N_27961,N_27106);
and U28959 (N_28959,N_27266,N_28123);
xnor U28960 (N_28960,N_27242,N_27632);
nand U28961 (N_28961,N_28337,N_27432);
xnor U28962 (N_28962,N_27619,N_27346);
or U28963 (N_28963,N_27422,N_27685);
nor U28964 (N_28964,N_27637,N_27714);
and U28965 (N_28965,N_27541,N_28134);
or U28966 (N_28966,N_28019,N_28034);
nor U28967 (N_28967,N_27855,N_27869);
nor U28968 (N_28968,N_27260,N_27608);
and U28969 (N_28969,N_27911,N_27276);
nor U28970 (N_28970,N_27170,N_27881);
nand U28971 (N_28971,N_27160,N_27527);
and U28972 (N_28972,N_27971,N_28375);
nor U28973 (N_28973,N_28311,N_28102);
or U28974 (N_28974,N_27566,N_27228);
xor U28975 (N_28975,N_27693,N_27494);
nand U28976 (N_28976,N_28186,N_27360);
xnor U28977 (N_28977,N_27909,N_28433);
and U28978 (N_28978,N_27839,N_27398);
nor U28979 (N_28979,N_28342,N_27629);
xor U28980 (N_28980,N_27834,N_28014);
nand U28981 (N_28981,N_27831,N_27318);
nand U28982 (N_28982,N_28331,N_28258);
and U28983 (N_28983,N_28053,N_27512);
nand U28984 (N_28984,N_27862,N_28332);
nor U28985 (N_28985,N_27484,N_27144);
or U28986 (N_28986,N_27937,N_27899);
or U28987 (N_28987,N_27073,N_27307);
or U28988 (N_28988,N_27275,N_28175);
nor U28989 (N_28989,N_28492,N_28122);
nand U28990 (N_28990,N_27290,N_27185);
nor U28991 (N_28991,N_27046,N_28174);
and U28992 (N_28992,N_28425,N_27103);
and U28993 (N_28993,N_27150,N_27211);
or U28994 (N_28994,N_27680,N_27167);
and U28995 (N_28995,N_27905,N_27030);
nand U28996 (N_28996,N_28005,N_28041);
and U28997 (N_28997,N_27980,N_27782);
nor U28998 (N_28998,N_27487,N_27710);
xor U28999 (N_28999,N_28431,N_27754);
nor U29000 (N_29000,N_28141,N_27413);
nor U29001 (N_29001,N_28329,N_27365);
or U29002 (N_29002,N_27357,N_27695);
or U29003 (N_29003,N_27173,N_28216);
or U29004 (N_29004,N_27457,N_27255);
xor U29005 (N_29005,N_27604,N_27120);
or U29006 (N_29006,N_28313,N_28108);
nor U29007 (N_29007,N_27773,N_28448);
and U29008 (N_29008,N_28485,N_28177);
nand U29009 (N_29009,N_28262,N_27114);
nand U29010 (N_29010,N_27278,N_27270);
nor U29011 (N_29011,N_27549,N_28488);
nor U29012 (N_29012,N_27412,N_27148);
xor U29013 (N_29013,N_27897,N_27408);
xor U29014 (N_29014,N_28091,N_27664);
nand U29015 (N_29015,N_27738,N_27688);
nor U29016 (N_29016,N_28105,N_27061);
or U29017 (N_29017,N_27965,N_28274);
xor U29018 (N_29018,N_28321,N_28117);
nand U29019 (N_29019,N_28338,N_27729);
and U29020 (N_29020,N_28319,N_27274);
and U29021 (N_29021,N_27810,N_27884);
nand U29022 (N_29022,N_27719,N_28450);
xnor U29023 (N_29023,N_28480,N_27386);
nor U29024 (N_29024,N_27417,N_27994);
nor U29025 (N_29025,N_28444,N_27711);
or U29026 (N_29026,N_28355,N_28138);
and U29027 (N_29027,N_28393,N_27654);
or U29028 (N_29028,N_27896,N_27169);
and U29029 (N_29029,N_27010,N_27420);
xor U29030 (N_29030,N_28144,N_28204);
and U29031 (N_29031,N_28133,N_28465);
and U29032 (N_29032,N_27922,N_27366);
nand U29033 (N_29033,N_28149,N_27948);
nor U29034 (N_29034,N_28143,N_27435);
or U29035 (N_29035,N_27414,N_27288);
or U29036 (N_29036,N_28297,N_27175);
or U29037 (N_29037,N_27411,N_27583);
nand U29038 (N_29038,N_28462,N_27014);
nand U29039 (N_29039,N_28306,N_27320);
nor U29040 (N_29040,N_27717,N_27058);
xnor U29041 (N_29041,N_28100,N_28155);
or U29042 (N_29042,N_27066,N_28059);
nor U29043 (N_29043,N_28477,N_27622);
nor U29044 (N_29044,N_27923,N_27032);
nor U29045 (N_29045,N_27758,N_27134);
xor U29046 (N_29046,N_28404,N_27451);
nor U29047 (N_29047,N_27477,N_27076);
xnor U29048 (N_29048,N_27951,N_27462);
and U29049 (N_29049,N_27168,N_28162);
xor U29050 (N_29050,N_27236,N_27368);
xor U29051 (N_29051,N_27102,N_27341);
nand U29052 (N_29052,N_27027,N_28231);
xor U29053 (N_29053,N_27891,N_27195);
or U29054 (N_29054,N_27034,N_27885);
nand U29055 (N_29055,N_28118,N_28446);
nor U29056 (N_29056,N_27850,N_27962);
nor U29057 (N_29057,N_28391,N_27842);
and U29058 (N_29058,N_27634,N_28129);
nor U29059 (N_29059,N_27988,N_28222);
or U29060 (N_29060,N_27985,N_27174);
and U29061 (N_29061,N_27548,N_27806);
or U29062 (N_29062,N_27603,N_27838);
and U29063 (N_29063,N_28322,N_27031);
xor U29064 (N_29064,N_27051,N_28242);
nor U29065 (N_29065,N_27402,N_27642);
nand U29066 (N_29066,N_28254,N_27311);
or U29067 (N_29067,N_27747,N_27463);
and U29068 (N_29068,N_27941,N_28495);
nor U29069 (N_29069,N_27390,N_27799);
or U29070 (N_29070,N_28369,N_28354);
and U29071 (N_29071,N_27005,N_27252);
nor U29072 (N_29072,N_28037,N_27696);
nand U29073 (N_29073,N_27018,N_27429);
nor U29074 (N_29074,N_28227,N_27702);
nand U29075 (N_29075,N_27771,N_28275);
or U29076 (N_29076,N_27229,N_27529);
nor U29077 (N_29077,N_27423,N_28429);
nor U29078 (N_29078,N_27845,N_27727);
and U29079 (N_29079,N_28033,N_27662);
or U29080 (N_29080,N_27142,N_28147);
or U29081 (N_29081,N_28020,N_27804);
nor U29082 (N_29082,N_27485,N_27780);
or U29083 (N_29083,N_27864,N_28273);
nor U29084 (N_29084,N_27716,N_27749);
and U29085 (N_29085,N_28312,N_27326);
or U29086 (N_29086,N_27172,N_28215);
nand U29087 (N_29087,N_27461,N_27094);
nor U29088 (N_29088,N_27661,N_27210);
nand U29089 (N_29089,N_27442,N_28081);
nor U29090 (N_29090,N_27241,N_27640);
nor U29091 (N_29091,N_27271,N_27131);
xor U29092 (N_29092,N_27340,N_28096);
or U29093 (N_29093,N_27865,N_27969);
or U29094 (N_29094,N_27056,N_28010);
xnor U29095 (N_29095,N_27383,N_27858);
nand U29096 (N_29096,N_28394,N_27355);
and U29097 (N_29097,N_27721,N_28484);
nor U29098 (N_29098,N_27145,N_27358);
xnor U29099 (N_29099,N_27446,N_28009);
xnor U29100 (N_29100,N_28163,N_27960);
and U29101 (N_29101,N_27459,N_27709);
nor U29102 (N_29102,N_28289,N_28076);
xnor U29103 (N_29103,N_27237,N_28469);
xor U29104 (N_29104,N_27746,N_28137);
xor U29105 (N_29105,N_27225,N_27013);
nand U29106 (N_29106,N_27766,N_27987);
or U29107 (N_29107,N_28383,N_27718);
xnor U29108 (N_29108,N_27104,N_28476);
or U29109 (N_29109,N_27503,N_28237);
xnor U29110 (N_29110,N_27706,N_27761);
nor U29111 (N_29111,N_27515,N_27686);
xnor U29112 (N_29112,N_27751,N_28409);
nor U29113 (N_29113,N_27560,N_27510);
nor U29114 (N_29114,N_27523,N_28381);
xnor U29115 (N_29115,N_27930,N_27065);
and U29116 (N_29116,N_28196,N_27772);
xnor U29117 (N_29117,N_27123,N_28472);
xor U29118 (N_29118,N_27534,N_27847);
and U29119 (N_29119,N_27441,N_27391);
and U29120 (N_29120,N_27359,N_27671);
and U29121 (N_29121,N_27044,N_28146);
or U29122 (N_29122,N_27561,N_28051);
or U29123 (N_29123,N_27111,N_27098);
xor U29124 (N_29124,N_27090,N_28127);
nand U29125 (N_29125,N_27028,N_27882);
and U29126 (N_29126,N_27796,N_27638);
or U29127 (N_29127,N_27546,N_28438);
nand U29128 (N_29128,N_27888,N_27598);
or U29129 (N_29129,N_28482,N_28294);
and U29130 (N_29130,N_27567,N_27039);
nand U29131 (N_29131,N_28184,N_28003);
nand U29132 (N_29132,N_28079,N_27280);
xor U29133 (N_29133,N_27498,N_28223);
or U29134 (N_29134,N_27085,N_27105);
or U29135 (N_29135,N_27997,N_28457);
xnor U29136 (N_29136,N_27597,N_27377);
and U29137 (N_29137,N_27743,N_28036);
or U29138 (N_29138,N_28454,N_28478);
nand U29139 (N_29139,N_27539,N_27596);
or U29140 (N_29140,N_27683,N_28244);
and U29141 (N_29141,N_27247,N_28346);
and U29142 (N_29142,N_28153,N_27844);
xnor U29143 (N_29143,N_27499,N_27594);
nor U29144 (N_29144,N_27322,N_27029);
xor U29145 (N_29145,N_28413,N_27556);
xor U29146 (N_29146,N_27165,N_28345);
nor U29147 (N_29147,N_27565,N_28082);
xnor U29148 (N_29148,N_27045,N_28234);
xor U29149 (N_29149,N_27760,N_27635);
and U29150 (N_29150,N_27200,N_27136);
or U29151 (N_29151,N_27995,N_27713);
or U29152 (N_29152,N_27734,N_27400);
nor U29153 (N_29153,N_28463,N_27912);
nand U29154 (N_29154,N_28140,N_28210);
or U29155 (N_29155,N_28491,N_27191);
and U29156 (N_29156,N_27240,N_27931);
and U29157 (N_29157,N_27176,N_28189);
nand U29158 (N_29158,N_27889,N_28418);
and U29159 (N_29159,N_27057,N_27993);
and U29160 (N_29160,N_27177,N_27395);
or U29161 (N_29161,N_27428,N_28318);
xor U29162 (N_29162,N_27430,N_27974);
nor U29163 (N_29163,N_27767,N_28449);
nand U29164 (N_29164,N_28265,N_27783);
xor U29165 (N_29165,N_27184,N_27444);
nor U29166 (N_29166,N_27580,N_27639);
nor U29167 (N_29167,N_27004,N_28006);
nor U29168 (N_29168,N_27554,N_27964);
xnor U29169 (N_29169,N_27433,N_27079);
or U29170 (N_29170,N_28235,N_27349);
nand U29171 (N_29171,N_27934,N_28427);
nor U29172 (N_29172,N_28271,N_27264);
nand U29173 (N_29173,N_27557,N_27968);
nor U29174 (N_29174,N_27925,N_28159);
nor U29175 (N_29175,N_27778,N_27309);
xor U29176 (N_29176,N_27947,N_28083);
nand U29177 (N_29177,N_27657,N_27687);
xnor U29178 (N_29178,N_27883,N_27720);
nand U29179 (N_29179,N_28435,N_27089);
nor U29180 (N_29180,N_28347,N_27404);
or U29181 (N_29181,N_27279,N_28023);
nor U29182 (N_29182,N_28468,N_28405);
xnor U29183 (N_29183,N_27943,N_28315);
nor U29184 (N_29184,N_27238,N_27917);
nand U29185 (N_29185,N_28185,N_27970);
and U29186 (N_29186,N_27471,N_28002);
nand U29187 (N_29187,N_28110,N_28460);
xnor U29188 (N_29188,N_27859,N_27643);
nand U29189 (N_29189,N_27578,N_28218);
and U29190 (N_29190,N_27426,N_27618);
nand U29191 (N_29191,N_27975,N_27976);
or U29192 (N_29192,N_28310,N_27853);
or U29193 (N_29193,N_27744,N_27822);
nor U29194 (N_29194,N_28441,N_27147);
nand U29195 (N_29195,N_27072,N_28360);
nand U29196 (N_29196,N_27456,N_27741);
nand U29197 (N_29197,N_28239,N_28428);
nor U29198 (N_29198,N_27880,N_28013);
or U29199 (N_29199,N_27978,N_27725);
and U29200 (N_29200,N_28065,N_27957);
xor U29201 (N_29201,N_27996,N_28161);
nor U29202 (N_29202,N_28103,N_27624);
and U29203 (N_29203,N_27857,N_27935);
nor U29204 (N_29204,N_27816,N_27339);
and U29205 (N_29205,N_27212,N_27986);
or U29206 (N_29206,N_27207,N_27458);
and U29207 (N_29207,N_27415,N_28384);
nor U29208 (N_29208,N_27514,N_28382);
and U29209 (N_29209,N_27866,N_28114);
nor U29210 (N_29210,N_27233,N_27797);
and U29211 (N_29211,N_27450,N_27759);
and U29212 (N_29212,N_27003,N_28291);
nor U29213 (N_29213,N_27659,N_27380);
xnor U29214 (N_29214,N_28259,N_27153);
and U29215 (N_29215,N_27926,N_28357);
or U29216 (N_29216,N_27077,N_28385);
xnor U29217 (N_29217,N_27723,N_27038);
nand U29218 (N_29218,N_27817,N_27363);
and U29219 (N_29219,N_27981,N_27314);
nand U29220 (N_29220,N_27963,N_28230);
and U29221 (N_29221,N_27213,N_27157);
and U29222 (N_29222,N_27752,N_28087);
nor U29223 (N_29223,N_27684,N_28334);
nand U29224 (N_29224,N_28481,N_27070);
xnor U29225 (N_29225,N_28356,N_27393);
nand U29226 (N_29226,N_27140,N_27616);
xor U29227 (N_29227,N_27119,N_27289);
nand U29228 (N_29228,N_27439,N_27250);
and U29229 (N_29229,N_27928,N_27472);
nand U29230 (N_29230,N_27248,N_27379);
nand U29231 (N_29231,N_28276,N_27369);
xor U29232 (N_29232,N_27082,N_27753);
nor U29233 (N_29233,N_28366,N_27129);
xnor U29234 (N_29234,N_27361,N_28192);
and U29235 (N_29235,N_27333,N_27701);
or U29236 (N_29236,N_27579,N_27699);
nor U29237 (N_29237,N_27455,N_27490);
xnor U29238 (N_29238,N_27910,N_27000);
and U29239 (N_29239,N_28220,N_27336);
or U29240 (N_29240,N_28151,N_27768);
and U29241 (N_29241,N_28466,N_27151);
and U29242 (N_29242,N_28071,N_28060);
or U29243 (N_29243,N_27125,N_27007);
xnor U29244 (N_29244,N_27330,N_28057);
nor U29245 (N_29245,N_27936,N_27466);
nand U29246 (N_29246,N_27586,N_27053);
xor U29247 (N_29247,N_27396,N_28004);
nor U29248 (N_29248,N_27068,N_27059);
nand U29249 (N_29249,N_27728,N_27660);
nand U29250 (N_29250,N_27547,N_27958);
nand U29251 (N_29251,N_28408,N_27438);
xnor U29252 (N_29252,N_27436,N_28458);
and U29253 (N_29253,N_28032,N_27252);
xnor U29254 (N_29254,N_27205,N_28123);
and U29255 (N_29255,N_28214,N_28489);
or U29256 (N_29256,N_27053,N_27976);
and U29257 (N_29257,N_27802,N_28179);
nand U29258 (N_29258,N_27163,N_28465);
xor U29259 (N_29259,N_28478,N_27831);
nor U29260 (N_29260,N_28478,N_27143);
and U29261 (N_29261,N_27120,N_27885);
nor U29262 (N_29262,N_27868,N_27410);
or U29263 (N_29263,N_27582,N_28266);
nor U29264 (N_29264,N_27403,N_28186);
nand U29265 (N_29265,N_27949,N_28254);
and U29266 (N_29266,N_27628,N_28440);
and U29267 (N_29267,N_27984,N_27312);
xnor U29268 (N_29268,N_27306,N_28419);
or U29269 (N_29269,N_27415,N_27827);
and U29270 (N_29270,N_27759,N_27517);
and U29271 (N_29271,N_28051,N_28249);
or U29272 (N_29272,N_28228,N_28336);
and U29273 (N_29273,N_27461,N_28027);
or U29274 (N_29274,N_27994,N_27109);
or U29275 (N_29275,N_27751,N_28348);
nor U29276 (N_29276,N_28432,N_28498);
nand U29277 (N_29277,N_27883,N_27422);
nor U29278 (N_29278,N_27846,N_27638);
nand U29279 (N_29279,N_28318,N_27622);
or U29280 (N_29280,N_27852,N_27866);
or U29281 (N_29281,N_27436,N_28127);
and U29282 (N_29282,N_27216,N_28150);
and U29283 (N_29283,N_27933,N_27257);
xor U29284 (N_29284,N_27501,N_28040);
nor U29285 (N_29285,N_27193,N_27391);
or U29286 (N_29286,N_28189,N_27548);
and U29287 (N_29287,N_27115,N_27827);
nand U29288 (N_29288,N_27067,N_27137);
xnor U29289 (N_29289,N_28331,N_28177);
and U29290 (N_29290,N_27954,N_27447);
xor U29291 (N_29291,N_28164,N_28033);
nor U29292 (N_29292,N_27734,N_28491);
and U29293 (N_29293,N_28301,N_27866);
and U29294 (N_29294,N_28075,N_27602);
and U29295 (N_29295,N_27714,N_27246);
and U29296 (N_29296,N_28329,N_28158);
nand U29297 (N_29297,N_28325,N_28037);
and U29298 (N_29298,N_28184,N_27472);
or U29299 (N_29299,N_27458,N_28260);
nand U29300 (N_29300,N_27729,N_27803);
xor U29301 (N_29301,N_27732,N_27489);
or U29302 (N_29302,N_27370,N_27303);
nor U29303 (N_29303,N_27751,N_27316);
nor U29304 (N_29304,N_28369,N_27421);
or U29305 (N_29305,N_27731,N_28384);
xor U29306 (N_29306,N_27895,N_27015);
or U29307 (N_29307,N_27110,N_27038);
nand U29308 (N_29308,N_27456,N_28374);
xnor U29309 (N_29309,N_27793,N_27329);
and U29310 (N_29310,N_27182,N_28436);
nand U29311 (N_29311,N_27665,N_27107);
and U29312 (N_29312,N_28279,N_27494);
and U29313 (N_29313,N_27348,N_28021);
nand U29314 (N_29314,N_27379,N_28109);
xor U29315 (N_29315,N_27567,N_27473);
nor U29316 (N_29316,N_27233,N_28204);
xor U29317 (N_29317,N_27055,N_28447);
and U29318 (N_29318,N_28060,N_27050);
and U29319 (N_29319,N_28228,N_28173);
and U29320 (N_29320,N_27436,N_28331);
or U29321 (N_29321,N_27409,N_28118);
nor U29322 (N_29322,N_27024,N_28225);
nand U29323 (N_29323,N_27014,N_28417);
xnor U29324 (N_29324,N_27729,N_28391);
xnor U29325 (N_29325,N_28030,N_27420);
or U29326 (N_29326,N_28471,N_28106);
and U29327 (N_29327,N_27079,N_28145);
xnor U29328 (N_29328,N_27934,N_27437);
xnor U29329 (N_29329,N_28292,N_27135);
nor U29330 (N_29330,N_27110,N_28474);
or U29331 (N_29331,N_27832,N_27890);
nor U29332 (N_29332,N_27116,N_27516);
or U29333 (N_29333,N_27919,N_27875);
and U29334 (N_29334,N_27668,N_28330);
xor U29335 (N_29335,N_27891,N_28498);
xnor U29336 (N_29336,N_27638,N_28215);
nand U29337 (N_29337,N_27871,N_28074);
nor U29338 (N_29338,N_27768,N_28402);
and U29339 (N_29339,N_27222,N_28487);
xor U29340 (N_29340,N_28442,N_27439);
xnor U29341 (N_29341,N_27729,N_28003);
nand U29342 (N_29342,N_27147,N_27258);
and U29343 (N_29343,N_27845,N_28132);
and U29344 (N_29344,N_27957,N_27410);
or U29345 (N_29345,N_28396,N_27618);
nand U29346 (N_29346,N_27732,N_27875);
nand U29347 (N_29347,N_27069,N_27079);
or U29348 (N_29348,N_27504,N_27702);
and U29349 (N_29349,N_28265,N_27999);
xnor U29350 (N_29350,N_27352,N_27307);
nor U29351 (N_29351,N_28052,N_27989);
nand U29352 (N_29352,N_28442,N_27609);
and U29353 (N_29353,N_28278,N_28333);
and U29354 (N_29354,N_27674,N_28119);
nand U29355 (N_29355,N_27826,N_27046);
or U29356 (N_29356,N_28042,N_27745);
nand U29357 (N_29357,N_28399,N_27871);
and U29358 (N_29358,N_27042,N_27056);
nand U29359 (N_29359,N_28155,N_28327);
or U29360 (N_29360,N_27463,N_27127);
or U29361 (N_29361,N_27899,N_27728);
and U29362 (N_29362,N_28141,N_27885);
nor U29363 (N_29363,N_27366,N_27566);
and U29364 (N_29364,N_27007,N_28476);
nor U29365 (N_29365,N_27291,N_28459);
and U29366 (N_29366,N_27130,N_27648);
nor U29367 (N_29367,N_27728,N_28105);
or U29368 (N_29368,N_27054,N_27167);
nor U29369 (N_29369,N_28453,N_27358);
xor U29370 (N_29370,N_28246,N_28209);
and U29371 (N_29371,N_27756,N_28357);
nor U29372 (N_29372,N_28033,N_27401);
or U29373 (N_29373,N_28440,N_28296);
and U29374 (N_29374,N_28372,N_28201);
nand U29375 (N_29375,N_28474,N_27535);
and U29376 (N_29376,N_27711,N_28345);
nor U29377 (N_29377,N_28478,N_27432);
or U29378 (N_29378,N_27844,N_27219);
nand U29379 (N_29379,N_27043,N_27817);
nor U29380 (N_29380,N_27907,N_27009);
or U29381 (N_29381,N_28451,N_28366);
and U29382 (N_29382,N_28089,N_27306);
nand U29383 (N_29383,N_27180,N_28404);
nand U29384 (N_29384,N_27005,N_27976);
nand U29385 (N_29385,N_28072,N_27073);
nand U29386 (N_29386,N_27660,N_27845);
nand U29387 (N_29387,N_27891,N_27506);
nor U29388 (N_29388,N_27199,N_28481);
xor U29389 (N_29389,N_27100,N_28290);
xnor U29390 (N_29390,N_27953,N_27186);
xnor U29391 (N_29391,N_27152,N_27405);
xnor U29392 (N_29392,N_28123,N_27281);
or U29393 (N_29393,N_27401,N_27303);
nand U29394 (N_29394,N_27247,N_28322);
xor U29395 (N_29395,N_27312,N_28150);
or U29396 (N_29396,N_27943,N_27886);
and U29397 (N_29397,N_28161,N_27835);
nor U29398 (N_29398,N_28414,N_28123);
nor U29399 (N_29399,N_28462,N_28220);
or U29400 (N_29400,N_28478,N_28451);
or U29401 (N_29401,N_27491,N_28024);
xnor U29402 (N_29402,N_27134,N_28472);
or U29403 (N_29403,N_28036,N_27513);
or U29404 (N_29404,N_28310,N_27556);
nor U29405 (N_29405,N_28293,N_27292);
nand U29406 (N_29406,N_27634,N_27125);
nor U29407 (N_29407,N_28460,N_27545);
or U29408 (N_29408,N_27480,N_27948);
and U29409 (N_29409,N_27358,N_27489);
nand U29410 (N_29410,N_27028,N_27872);
nor U29411 (N_29411,N_27493,N_27942);
xor U29412 (N_29412,N_27742,N_28141);
or U29413 (N_29413,N_28010,N_27693);
xnor U29414 (N_29414,N_27093,N_28324);
nand U29415 (N_29415,N_27311,N_27426);
xor U29416 (N_29416,N_27731,N_27812);
or U29417 (N_29417,N_27547,N_27671);
nor U29418 (N_29418,N_27913,N_27636);
nor U29419 (N_29419,N_28407,N_27933);
and U29420 (N_29420,N_28125,N_27514);
nand U29421 (N_29421,N_27515,N_28003);
or U29422 (N_29422,N_27696,N_27377);
or U29423 (N_29423,N_27525,N_27681);
nor U29424 (N_29424,N_27379,N_27307);
or U29425 (N_29425,N_27772,N_27234);
nor U29426 (N_29426,N_27415,N_27034);
or U29427 (N_29427,N_28235,N_27121);
nand U29428 (N_29428,N_27222,N_28225);
and U29429 (N_29429,N_27536,N_27287);
or U29430 (N_29430,N_28174,N_27649);
and U29431 (N_29431,N_27834,N_27850);
nand U29432 (N_29432,N_28401,N_28306);
or U29433 (N_29433,N_27768,N_27626);
nand U29434 (N_29434,N_28492,N_27719);
and U29435 (N_29435,N_27406,N_28412);
nand U29436 (N_29436,N_27304,N_27006);
nand U29437 (N_29437,N_28113,N_28217);
or U29438 (N_29438,N_27766,N_27095);
or U29439 (N_29439,N_27111,N_27310);
or U29440 (N_29440,N_28324,N_27438);
and U29441 (N_29441,N_27149,N_27994);
xor U29442 (N_29442,N_27912,N_28461);
nor U29443 (N_29443,N_27283,N_27725);
and U29444 (N_29444,N_27533,N_28041);
or U29445 (N_29445,N_27998,N_28351);
nor U29446 (N_29446,N_27143,N_28197);
or U29447 (N_29447,N_28379,N_27556);
nand U29448 (N_29448,N_28320,N_28469);
and U29449 (N_29449,N_27725,N_27254);
nand U29450 (N_29450,N_28273,N_27787);
nor U29451 (N_29451,N_27890,N_27448);
nor U29452 (N_29452,N_27759,N_27617);
xor U29453 (N_29453,N_27371,N_27177);
xnor U29454 (N_29454,N_27275,N_28242);
nor U29455 (N_29455,N_28400,N_28439);
xor U29456 (N_29456,N_28497,N_27861);
and U29457 (N_29457,N_27388,N_27137);
nand U29458 (N_29458,N_27312,N_28260);
and U29459 (N_29459,N_27071,N_27712);
or U29460 (N_29460,N_27779,N_28346);
nor U29461 (N_29461,N_27414,N_27530);
nor U29462 (N_29462,N_27496,N_28481);
nor U29463 (N_29463,N_28313,N_27195);
and U29464 (N_29464,N_27255,N_27913);
and U29465 (N_29465,N_27651,N_27454);
nand U29466 (N_29466,N_27021,N_27636);
and U29467 (N_29467,N_27371,N_28241);
and U29468 (N_29468,N_27300,N_28029);
nor U29469 (N_29469,N_27264,N_27494);
xnor U29470 (N_29470,N_27452,N_27331);
nand U29471 (N_29471,N_27550,N_27047);
xor U29472 (N_29472,N_28094,N_27984);
and U29473 (N_29473,N_27873,N_28482);
nor U29474 (N_29474,N_27236,N_28091);
or U29475 (N_29475,N_27047,N_28456);
or U29476 (N_29476,N_27676,N_27128);
xnor U29477 (N_29477,N_28325,N_27719);
nand U29478 (N_29478,N_27719,N_27861);
nand U29479 (N_29479,N_27224,N_27783);
nor U29480 (N_29480,N_28244,N_27481);
nand U29481 (N_29481,N_28311,N_28418);
xor U29482 (N_29482,N_28030,N_27331);
nor U29483 (N_29483,N_27760,N_27213);
and U29484 (N_29484,N_27155,N_28281);
nor U29485 (N_29485,N_27297,N_27058);
nor U29486 (N_29486,N_28396,N_28276);
nand U29487 (N_29487,N_28372,N_27189);
nand U29488 (N_29488,N_27121,N_28231);
xor U29489 (N_29489,N_27597,N_27115);
or U29490 (N_29490,N_27489,N_28307);
nor U29491 (N_29491,N_27095,N_27786);
or U29492 (N_29492,N_27674,N_27368);
nand U29493 (N_29493,N_27163,N_27490);
or U29494 (N_29494,N_27164,N_27498);
nand U29495 (N_29495,N_27698,N_27239);
nand U29496 (N_29496,N_27417,N_27912);
nor U29497 (N_29497,N_27221,N_28061);
xor U29498 (N_29498,N_27967,N_27999);
nand U29499 (N_29499,N_28229,N_27420);
or U29500 (N_29500,N_27575,N_27118);
nor U29501 (N_29501,N_27732,N_27944);
xor U29502 (N_29502,N_28107,N_28447);
xnor U29503 (N_29503,N_28493,N_28461);
xor U29504 (N_29504,N_27469,N_28069);
nand U29505 (N_29505,N_28152,N_27222);
and U29506 (N_29506,N_28492,N_27920);
xnor U29507 (N_29507,N_27815,N_27600);
and U29508 (N_29508,N_27147,N_27747);
xor U29509 (N_29509,N_27155,N_28475);
nand U29510 (N_29510,N_27191,N_27860);
and U29511 (N_29511,N_28317,N_28044);
or U29512 (N_29512,N_27138,N_27029);
or U29513 (N_29513,N_27435,N_27150);
xor U29514 (N_29514,N_27566,N_27092);
xnor U29515 (N_29515,N_28169,N_28414);
nor U29516 (N_29516,N_28490,N_28388);
xnor U29517 (N_29517,N_27912,N_27593);
nor U29518 (N_29518,N_27055,N_27381);
xor U29519 (N_29519,N_27270,N_27261);
and U29520 (N_29520,N_27331,N_27461);
xor U29521 (N_29521,N_28453,N_27881);
or U29522 (N_29522,N_27250,N_27652);
nand U29523 (N_29523,N_27287,N_28331);
nand U29524 (N_29524,N_27321,N_27653);
xor U29525 (N_29525,N_27227,N_28119);
nand U29526 (N_29526,N_28495,N_27988);
xor U29527 (N_29527,N_27780,N_28199);
nor U29528 (N_29528,N_28078,N_28141);
and U29529 (N_29529,N_28052,N_27414);
nor U29530 (N_29530,N_28489,N_27195);
nor U29531 (N_29531,N_27556,N_28366);
or U29532 (N_29532,N_28386,N_27853);
xnor U29533 (N_29533,N_27172,N_27123);
xor U29534 (N_29534,N_27455,N_27235);
and U29535 (N_29535,N_27417,N_28061);
xnor U29536 (N_29536,N_27741,N_28210);
xnor U29537 (N_29537,N_28236,N_27845);
nor U29538 (N_29538,N_27171,N_27263);
and U29539 (N_29539,N_27450,N_27376);
or U29540 (N_29540,N_27410,N_28069);
nand U29541 (N_29541,N_28289,N_27116);
or U29542 (N_29542,N_27987,N_28024);
xnor U29543 (N_29543,N_28386,N_27929);
xor U29544 (N_29544,N_27757,N_28303);
and U29545 (N_29545,N_27551,N_27788);
nor U29546 (N_29546,N_27393,N_27561);
nand U29547 (N_29547,N_27224,N_27585);
and U29548 (N_29548,N_27703,N_28495);
nand U29549 (N_29549,N_27973,N_27438);
nor U29550 (N_29550,N_28035,N_27381);
nor U29551 (N_29551,N_28190,N_28460);
or U29552 (N_29552,N_27754,N_27243);
or U29553 (N_29553,N_27241,N_27372);
or U29554 (N_29554,N_28354,N_28387);
nand U29555 (N_29555,N_27910,N_27176);
and U29556 (N_29556,N_27748,N_28282);
or U29557 (N_29557,N_27986,N_27939);
nor U29558 (N_29558,N_27740,N_28239);
or U29559 (N_29559,N_28243,N_28321);
nand U29560 (N_29560,N_27782,N_27493);
and U29561 (N_29561,N_28239,N_27469);
xnor U29562 (N_29562,N_27327,N_27406);
nand U29563 (N_29563,N_27068,N_27395);
and U29564 (N_29564,N_27571,N_27567);
or U29565 (N_29565,N_28130,N_27858);
or U29566 (N_29566,N_27491,N_28262);
nand U29567 (N_29567,N_27824,N_27885);
and U29568 (N_29568,N_27798,N_28374);
nor U29569 (N_29569,N_27564,N_28216);
nor U29570 (N_29570,N_28271,N_28302);
xor U29571 (N_29571,N_28495,N_27070);
and U29572 (N_29572,N_28444,N_27587);
nand U29573 (N_29573,N_27744,N_27635);
nand U29574 (N_29574,N_28438,N_28057);
or U29575 (N_29575,N_27439,N_28342);
nand U29576 (N_29576,N_27489,N_27600);
or U29577 (N_29577,N_27547,N_27333);
xor U29578 (N_29578,N_28413,N_28425);
nand U29579 (N_29579,N_27384,N_28395);
or U29580 (N_29580,N_28280,N_28282);
or U29581 (N_29581,N_27871,N_27532);
nor U29582 (N_29582,N_27298,N_28092);
or U29583 (N_29583,N_27713,N_27972);
xnor U29584 (N_29584,N_27255,N_28151);
xor U29585 (N_29585,N_27136,N_28267);
nor U29586 (N_29586,N_27724,N_27283);
nand U29587 (N_29587,N_27497,N_27904);
or U29588 (N_29588,N_28209,N_27797);
nand U29589 (N_29589,N_27758,N_27311);
and U29590 (N_29590,N_27839,N_28351);
nand U29591 (N_29591,N_27165,N_28335);
nand U29592 (N_29592,N_27058,N_27873);
or U29593 (N_29593,N_28187,N_27787);
nor U29594 (N_29594,N_27064,N_27440);
or U29595 (N_29595,N_27305,N_27842);
nand U29596 (N_29596,N_27270,N_28124);
nor U29597 (N_29597,N_27683,N_28367);
nor U29598 (N_29598,N_27762,N_27858);
or U29599 (N_29599,N_27434,N_27069);
or U29600 (N_29600,N_27401,N_27829);
and U29601 (N_29601,N_27477,N_27540);
and U29602 (N_29602,N_27233,N_28202);
or U29603 (N_29603,N_27103,N_28264);
nor U29604 (N_29604,N_27496,N_28174);
or U29605 (N_29605,N_27506,N_27397);
nand U29606 (N_29606,N_27720,N_27948);
nand U29607 (N_29607,N_27367,N_28329);
nand U29608 (N_29608,N_28117,N_27232);
nor U29609 (N_29609,N_27089,N_27490);
or U29610 (N_29610,N_28142,N_27996);
nor U29611 (N_29611,N_28055,N_28210);
nor U29612 (N_29612,N_27945,N_27195);
nand U29613 (N_29613,N_27447,N_27354);
nor U29614 (N_29614,N_27018,N_28142);
xor U29615 (N_29615,N_28228,N_27387);
and U29616 (N_29616,N_27558,N_27954);
or U29617 (N_29617,N_28489,N_28302);
and U29618 (N_29618,N_27299,N_28262);
nand U29619 (N_29619,N_27562,N_27786);
and U29620 (N_29620,N_27741,N_28283);
and U29621 (N_29621,N_28430,N_28184);
xor U29622 (N_29622,N_27335,N_27561);
xnor U29623 (N_29623,N_27919,N_27326);
and U29624 (N_29624,N_27619,N_27070);
nor U29625 (N_29625,N_28250,N_27176);
and U29626 (N_29626,N_27919,N_28477);
nor U29627 (N_29627,N_27949,N_27409);
xor U29628 (N_29628,N_28136,N_28133);
xor U29629 (N_29629,N_27418,N_28224);
xor U29630 (N_29630,N_28300,N_27541);
xnor U29631 (N_29631,N_27343,N_27899);
or U29632 (N_29632,N_27712,N_27126);
and U29633 (N_29633,N_28429,N_27226);
and U29634 (N_29634,N_28260,N_27167);
and U29635 (N_29635,N_28107,N_27549);
nor U29636 (N_29636,N_27396,N_27797);
or U29637 (N_29637,N_27416,N_27572);
nand U29638 (N_29638,N_28155,N_28325);
and U29639 (N_29639,N_28297,N_28034);
xnor U29640 (N_29640,N_28366,N_28347);
or U29641 (N_29641,N_28023,N_27552);
and U29642 (N_29642,N_27494,N_27021);
nor U29643 (N_29643,N_28175,N_27102);
and U29644 (N_29644,N_27719,N_27644);
or U29645 (N_29645,N_27386,N_27841);
nor U29646 (N_29646,N_27523,N_27950);
xor U29647 (N_29647,N_27129,N_28449);
nor U29648 (N_29648,N_28150,N_28174);
xnor U29649 (N_29649,N_28430,N_27507);
nand U29650 (N_29650,N_27832,N_28403);
and U29651 (N_29651,N_27094,N_28122);
xor U29652 (N_29652,N_27756,N_27249);
and U29653 (N_29653,N_27285,N_28469);
or U29654 (N_29654,N_27923,N_28321);
or U29655 (N_29655,N_28278,N_27308);
and U29656 (N_29656,N_27940,N_27845);
or U29657 (N_29657,N_28438,N_27484);
or U29658 (N_29658,N_27923,N_27547);
nor U29659 (N_29659,N_27328,N_27890);
and U29660 (N_29660,N_27966,N_27982);
nand U29661 (N_29661,N_27874,N_27409);
nor U29662 (N_29662,N_28414,N_28387);
nand U29663 (N_29663,N_27123,N_27788);
and U29664 (N_29664,N_27791,N_27657);
or U29665 (N_29665,N_27937,N_28371);
xnor U29666 (N_29666,N_27319,N_27104);
nor U29667 (N_29667,N_27746,N_28311);
nor U29668 (N_29668,N_27347,N_27379);
nand U29669 (N_29669,N_28212,N_27824);
or U29670 (N_29670,N_27513,N_27552);
xnor U29671 (N_29671,N_27491,N_28274);
and U29672 (N_29672,N_27325,N_27127);
or U29673 (N_29673,N_28416,N_27866);
xnor U29674 (N_29674,N_27590,N_27221);
or U29675 (N_29675,N_28440,N_27312);
or U29676 (N_29676,N_27703,N_28392);
nand U29677 (N_29677,N_28228,N_27234);
or U29678 (N_29678,N_28466,N_28295);
or U29679 (N_29679,N_27913,N_28198);
nand U29680 (N_29680,N_27071,N_28036);
or U29681 (N_29681,N_27065,N_27371);
nor U29682 (N_29682,N_27056,N_27494);
and U29683 (N_29683,N_27697,N_27323);
and U29684 (N_29684,N_27160,N_27403);
and U29685 (N_29685,N_27791,N_27252);
or U29686 (N_29686,N_28425,N_27613);
xnor U29687 (N_29687,N_28077,N_28017);
nor U29688 (N_29688,N_27192,N_27725);
nand U29689 (N_29689,N_28324,N_27193);
and U29690 (N_29690,N_27997,N_27259);
xnor U29691 (N_29691,N_27351,N_27781);
and U29692 (N_29692,N_27601,N_27119);
xnor U29693 (N_29693,N_28225,N_28240);
and U29694 (N_29694,N_27815,N_28083);
nor U29695 (N_29695,N_27976,N_28073);
and U29696 (N_29696,N_28460,N_28050);
nor U29697 (N_29697,N_28183,N_27997);
or U29698 (N_29698,N_28231,N_28318);
nor U29699 (N_29699,N_27529,N_28362);
and U29700 (N_29700,N_27661,N_28028);
nand U29701 (N_29701,N_27340,N_27502);
and U29702 (N_29702,N_27154,N_28251);
or U29703 (N_29703,N_27370,N_27236);
and U29704 (N_29704,N_27071,N_28139);
and U29705 (N_29705,N_27725,N_27879);
xnor U29706 (N_29706,N_28070,N_28025);
and U29707 (N_29707,N_28245,N_27371);
nand U29708 (N_29708,N_27202,N_28138);
and U29709 (N_29709,N_27577,N_27303);
or U29710 (N_29710,N_27963,N_28311);
xnor U29711 (N_29711,N_28034,N_28291);
and U29712 (N_29712,N_27364,N_27263);
xor U29713 (N_29713,N_27638,N_27666);
nand U29714 (N_29714,N_27859,N_27750);
nand U29715 (N_29715,N_28057,N_27550);
and U29716 (N_29716,N_28115,N_28357);
or U29717 (N_29717,N_27464,N_27946);
xor U29718 (N_29718,N_27488,N_27995);
or U29719 (N_29719,N_27548,N_27634);
nor U29720 (N_29720,N_27386,N_28350);
or U29721 (N_29721,N_27858,N_28273);
and U29722 (N_29722,N_27026,N_28456);
and U29723 (N_29723,N_27155,N_27146);
and U29724 (N_29724,N_27013,N_28409);
nand U29725 (N_29725,N_27004,N_27457);
and U29726 (N_29726,N_27229,N_27651);
and U29727 (N_29727,N_28199,N_28149);
and U29728 (N_29728,N_27543,N_27854);
and U29729 (N_29729,N_27870,N_27909);
and U29730 (N_29730,N_27533,N_27988);
or U29731 (N_29731,N_27800,N_27664);
xor U29732 (N_29732,N_28485,N_28411);
nand U29733 (N_29733,N_27556,N_27590);
xor U29734 (N_29734,N_27920,N_27162);
xnor U29735 (N_29735,N_27373,N_27443);
and U29736 (N_29736,N_27753,N_28430);
or U29737 (N_29737,N_27784,N_27034);
or U29738 (N_29738,N_28287,N_27560);
and U29739 (N_29739,N_27974,N_28121);
and U29740 (N_29740,N_28375,N_27271);
nor U29741 (N_29741,N_28357,N_28079);
and U29742 (N_29742,N_28212,N_27001);
nand U29743 (N_29743,N_27430,N_27051);
nor U29744 (N_29744,N_28109,N_28449);
nor U29745 (N_29745,N_27084,N_27603);
nor U29746 (N_29746,N_27512,N_27082);
nor U29747 (N_29747,N_27863,N_27776);
or U29748 (N_29748,N_27432,N_28384);
or U29749 (N_29749,N_27254,N_28211);
and U29750 (N_29750,N_27910,N_27306);
or U29751 (N_29751,N_27462,N_27494);
nor U29752 (N_29752,N_27713,N_27567);
and U29753 (N_29753,N_27925,N_27848);
nand U29754 (N_29754,N_28174,N_27812);
nor U29755 (N_29755,N_27047,N_27565);
nor U29756 (N_29756,N_27264,N_27702);
xor U29757 (N_29757,N_27723,N_27534);
and U29758 (N_29758,N_27807,N_27029);
xor U29759 (N_29759,N_27060,N_27010);
nor U29760 (N_29760,N_27877,N_28223);
nand U29761 (N_29761,N_27294,N_27449);
xnor U29762 (N_29762,N_27989,N_27034);
nor U29763 (N_29763,N_28266,N_28215);
xor U29764 (N_29764,N_27626,N_27118);
and U29765 (N_29765,N_28154,N_28102);
xor U29766 (N_29766,N_28016,N_28464);
nand U29767 (N_29767,N_28494,N_27346);
or U29768 (N_29768,N_28265,N_27996);
nor U29769 (N_29769,N_27965,N_28308);
and U29770 (N_29770,N_27638,N_27696);
or U29771 (N_29771,N_27937,N_27889);
nand U29772 (N_29772,N_28307,N_27031);
nand U29773 (N_29773,N_27785,N_28068);
nand U29774 (N_29774,N_27351,N_27399);
nor U29775 (N_29775,N_27286,N_27066);
xor U29776 (N_29776,N_27237,N_27012);
and U29777 (N_29777,N_27994,N_27043);
and U29778 (N_29778,N_27971,N_27389);
xor U29779 (N_29779,N_27246,N_27347);
and U29780 (N_29780,N_27761,N_27863);
and U29781 (N_29781,N_27377,N_28257);
and U29782 (N_29782,N_28375,N_27388);
and U29783 (N_29783,N_27222,N_27485);
nand U29784 (N_29784,N_28426,N_28453);
xor U29785 (N_29785,N_27836,N_27723);
or U29786 (N_29786,N_28200,N_27960);
nor U29787 (N_29787,N_27189,N_28353);
and U29788 (N_29788,N_27103,N_28223);
nand U29789 (N_29789,N_27708,N_28100);
and U29790 (N_29790,N_27543,N_27249);
nor U29791 (N_29791,N_27007,N_27508);
nor U29792 (N_29792,N_27366,N_27623);
nand U29793 (N_29793,N_27125,N_27432);
and U29794 (N_29794,N_27886,N_28147);
nand U29795 (N_29795,N_27516,N_27634);
nand U29796 (N_29796,N_27666,N_27653);
and U29797 (N_29797,N_27285,N_27289);
nand U29798 (N_29798,N_28153,N_28186);
xor U29799 (N_29799,N_27490,N_28125);
nor U29800 (N_29800,N_27459,N_27644);
or U29801 (N_29801,N_27356,N_28029);
and U29802 (N_29802,N_27408,N_28284);
nand U29803 (N_29803,N_28028,N_27622);
and U29804 (N_29804,N_27586,N_27921);
xnor U29805 (N_29805,N_28325,N_28271);
or U29806 (N_29806,N_27044,N_27560);
or U29807 (N_29807,N_28217,N_27526);
or U29808 (N_29808,N_27682,N_28140);
nand U29809 (N_29809,N_28264,N_27764);
and U29810 (N_29810,N_27277,N_28199);
xnor U29811 (N_29811,N_27421,N_27452);
xnor U29812 (N_29812,N_27823,N_27034);
or U29813 (N_29813,N_27221,N_27098);
or U29814 (N_29814,N_28133,N_28319);
or U29815 (N_29815,N_27861,N_27688);
and U29816 (N_29816,N_28072,N_28428);
nand U29817 (N_29817,N_28084,N_28207);
and U29818 (N_29818,N_27003,N_28050);
nand U29819 (N_29819,N_28099,N_27420);
xor U29820 (N_29820,N_27687,N_27331);
and U29821 (N_29821,N_27068,N_27524);
xor U29822 (N_29822,N_28361,N_27197);
and U29823 (N_29823,N_27046,N_27422);
or U29824 (N_29824,N_27577,N_27725);
and U29825 (N_29825,N_28328,N_28305);
xnor U29826 (N_29826,N_28297,N_28176);
nor U29827 (N_29827,N_28366,N_28257);
xnor U29828 (N_29828,N_27313,N_27456);
nand U29829 (N_29829,N_28325,N_27068);
and U29830 (N_29830,N_27325,N_28440);
or U29831 (N_29831,N_27155,N_28132);
xor U29832 (N_29832,N_27726,N_27864);
and U29833 (N_29833,N_27291,N_28389);
or U29834 (N_29834,N_28366,N_27541);
and U29835 (N_29835,N_27466,N_27052);
xnor U29836 (N_29836,N_27137,N_27784);
xnor U29837 (N_29837,N_28123,N_28229);
xnor U29838 (N_29838,N_27726,N_28339);
nor U29839 (N_29839,N_27625,N_27502);
nor U29840 (N_29840,N_28113,N_28441);
xnor U29841 (N_29841,N_27672,N_27584);
xnor U29842 (N_29842,N_28231,N_27120);
xor U29843 (N_29843,N_28256,N_28162);
and U29844 (N_29844,N_27220,N_27982);
or U29845 (N_29845,N_27870,N_27803);
xnor U29846 (N_29846,N_27779,N_28247);
nor U29847 (N_29847,N_28109,N_28338);
nand U29848 (N_29848,N_27639,N_27801);
xor U29849 (N_29849,N_27046,N_28136);
xnor U29850 (N_29850,N_27001,N_27788);
nand U29851 (N_29851,N_27767,N_27819);
nand U29852 (N_29852,N_27125,N_28132);
xor U29853 (N_29853,N_28127,N_27416);
or U29854 (N_29854,N_27417,N_27830);
xnor U29855 (N_29855,N_27852,N_28100);
nor U29856 (N_29856,N_27819,N_28161);
nand U29857 (N_29857,N_27921,N_28073);
nor U29858 (N_29858,N_27629,N_28384);
xor U29859 (N_29859,N_28237,N_27088);
xor U29860 (N_29860,N_27361,N_27610);
nand U29861 (N_29861,N_27026,N_27536);
and U29862 (N_29862,N_28010,N_27062);
and U29863 (N_29863,N_27918,N_27292);
or U29864 (N_29864,N_28263,N_27642);
xor U29865 (N_29865,N_28466,N_27702);
and U29866 (N_29866,N_28159,N_27215);
nor U29867 (N_29867,N_28141,N_27149);
nor U29868 (N_29868,N_27496,N_27637);
and U29869 (N_29869,N_27908,N_28082);
or U29870 (N_29870,N_27428,N_27148);
nor U29871 (N_29871,N_28120,N_27848);
nand U29872 (N_29872,N_28425,N_27576);
xnor U29873 (N_29873,N_27505,N_27406);
nand U29874 (N_29874,N_28274,N_27122);
or U29875 (N_29875,N_27337,N_27778);
xnor U29876 (N_29876,N_27392,N_28155);
nor U29877 (N_29877,N_27858,N_28193);
nand U29878 (N_29878,N_27521,N_27007);
nand U29879 (N_29879,N_28078,N_28256);
xor U29880 (N_29880,N_28248,N_27189);
nand U29881 (N_29881,N_28027,N_27671);
and U29882 (N_29882,N_27198,N_27965);
nor U29883 (N_29883,N_27493,N_27852);
nor U29884 (N_29884,N_28168,N_27363);
or U29885 (N_29885,N_27788,N_28133);
or U29886 (N_29886,N_27082,N_28031);
nor U29887 (N_29887,N_27251,N_27101);
and U29888 (N_29888,N_27591,N_28008);
or U29889 (N_29889,N_28304,N_27671);
and U29890 (N_29890,N_27245,N_27962);
xor U29891 (N_29891,N_27241,N_27982);
nor U29892 (N_29892,N_28487,N_28071);
nor U29893 (N_29893,N_28045,N_28114);
nand U29894 (N_29894,N_27895,N_27765);
nand U29895 (N_29895,N_28421,N_28449);
and U29896 (N_29896,N_28234,N_28094);
and U29897 (N_29897,N_28369,N_27845);
or U29898 (N_29898,N_27537,N_27071);
or U29899 (N_29899,N_28163,N_28348);
or U29900 (N_29900,N_27763,N_28462);
nor U29901 (N_29901,N_27312,N_27059);
nor U29902 (N_29902,N_28043,N_28342);
and U29903 (N_29903,N_27959,N_28315);
or U29904 (N_29904,N_28078,N_28185);
xnor U29905 (N_29905,N_27300,N_27140);
xnor U29906 (N_29906,N_27099,N_27861);
nor U29907 (N_29907,N_28384,N_27730);
xor U29908 (N_29908,N_27046,N_27361);
or U29909 (N_29909,N_27190,N_28435);
or U29910 (N_29910,N_28345,N_28359);
and U29911 (N_29911,N_27662,N_27964);
xor U29912 (N_29912,N_28168,N_27826);
xnor U29913 (N_29913,N_27800,N_28195);
nor U29914 (N_29914,N_28014,N_27726);
or U29915 (N_29915,N_27654,N_28206);
nand U29916 (N_29916,N_28340,N_27715);
nand U29917 (N_29917,N_27622,N_27164);
nor U29918 (N_29918,N_28223,N_27863);
xor U29919 (N_29919,N_27091,N_27718);
xor U29920 (N_29920,N_27377,N_27263);
and U29921 (N_29921,N_28233,N_27425);
or U29922 (N_29922,N_27093,N_27432);
nor U29923 (N_29923,N_27249,N_27090);
xor U29924 (N_29924,N_27263,N_27984);
and U29925 (N_29925,N_28079,N_27433);
and U29926 (N_29926,N_28435,N_28235);
xnor U29927 (N_29927,N_28019,N_27341);
or U29928 (N_29928,N_27804,N_28482);
xnor U29929 (N_29929,N_27154,N_27954);
and U29930 (N_29930,N_27874,N_27336);
nand U29931 (N_29931,N_28157,N_27265);
xor U29932 (N_29932,N_27579,N_28200);
and U29933 (N_29933,N_27783,N_28330);
nor U29934 (N_29934,N_27123,N_27812);
xnor U29935 (N_29935,N_27435,N_27594);
and U29936 (N_29936,N_27906,N_27814);
and U29937 (N_29937,N_27858,N_28222);
or U29938 (N_29938,N_28256,N_27728);
and U29939 (N_29939,N_27488,N_27704);
nand U29940 (N_29940,N_27551,N_27101);
nand U29941 (N_29941,N_28448,N_27713);
nand U29942 (N_29942,N_27630,N_28092);
xor U29943 (N_29943,N_27855,N_27847);
nor U29944 (N_29944,N_27425,N_28450);
nor U29945 (N_29945,N_28041,N_27065);
and U29946 (N_29946,N_28249,N_28204);
and U29947 (N_29947,N_28427,N_28439);
nand U29948 (N_29948,N_28078,N_27592);
nor U29949 (N_29949,N_27930,N_27103);
and U29950 (N_29950,N_28461,N_27360);
or U29951 (N_29951,N_28066,N_27451);
nor U29952 (N_29952,N_27211,N_27160);
nand U29953 (N_29953,N_27498,N_27709);
nand U29954 (N_29954,N_27121,N_28145);
nor U29955 (N_29955,N_27379,N_27796);
and U29956 (N_29956,N_27222,N_28484);
nor U29957 (N_29957,N_28391,N_27313);
xor U29958 (N_29958,N_27899,N_28059);
xnor U29959 (N_29959,N_28400,N_27140);
nand U29960 (N_29960,N_27996,N_27250);
nor U29961 (N_29961,N_27945,N_27751);
nand U29962 (N_29962,N_27170,N_28008);
and U29963 (N_29963,N_28097,N_27626);
nor U29964 (N_29964,N_27888,N_27901);
and U29965 (N_29965,N_27792,N_27913);
nor U29966 (N_29966,N_27363,N_27456);
nand U29967 (N_29967,N_27024,N_27248);
xor U29968 (N_29968,N_27737,N_27466);
and U29969 (N_29969,N_27144,N_27283);
nor U29970 (N_29970,N_27374,N_28277);
xor U29971 (N_29971,N_27811,N_27098);
or U29972 (N_29972,N_27020,N_28283);
or U29973 (N_29973,N_27305,N_27769);
nor U29974 (N_29974,N_27617,N_27517);
nand U29975 (N_29975,N_27970,N_28494);
or U29976 (N_29976,N_27871,N_28369);
or U29977 (N_29977,N_28164,N_27681);
nand U29978 (N_29978,N_28063,N_27378);
nand U29979 (N_29979,N_28101,N_27978);
nand U29980 (N_29980,N_28414,N_27375);
xor U29981 (N_29981,N_28307,N_27359);
xnor U29982 (N_29982,N_28102,N_28124);
nor U29983 (N_29983,N_28306,N_28433);
nand U29984 (N_29984,N_27782,N_27498);
nor U29985 (N_29985,N_27550,N_27756);
or U29986 (N_29986,N_28020,N_27383);
and U29987 (N_29987,N_27140,N_27476);
or U29988 (N_29988,N_27151,N_27825);
nand U29989 (N_29989,N_28085,N_28499);
xnor U29990 (N_29990,N_28456,N_27895);
xor U29991 (N_29991,N_28358,N_27899);
or U29992 (N_29992,N_27811,N_27394);
xor U29993 (N_29993,N_28232,N_28329);
or U29994 (N_29994,N_27463,N_28450);
nor U29995 (N_29995,N_27329,N_27629);
and U29996 (N_29996,N_28314,N_27393);
nor U29997 (N_29997,N_27026,N_27654);
nor U29998 (N_29998,N_28235,N_28401);
xnor U29999 (N_29999,N_28343,N_28412);
and UO_0 (O_0,N_29197,N_29287);
or UO_1 (O_1,N_29955,N_28677);
nor UO_2 (O_2,N_29905,N_29186);
xnor UO_3 (O_3,N_29342,N_29031);
nand UO_4 (O_4,N_29935,N_29801);
nor UO_5 (O_5,N_28706,N_29367);
xnor UO_6 (O_6,N_29244,N_29979);
and UO_7 (O_7,N_29793,N_29318);
and UO_8 (O_8,N_29510,N_29994);
nor UO_9 (O_9,N_28550,N_29782);
nand UO_10 (O_10,N_29308,N_29634);
xor UO_11 (O_11,N_29565,N_28880);
nand UO_12 (O_12,N_28508,N_29242);
or UO_13 (O_13,N_29571,N_28609);
xnor UO_14 (O_14,N_29427,N_28997);
and UO_15 (O_15,N_29037,N_29878);
nand UO_16 (O_16,N_29666,N_29005);
nand UO_17 (O_17,N_29806,N_29385);
xnor UO_18 (O_18,N_29193,N_28962);
nand UO_19 (O_19,N_29681,N_28852);
xor UO_20 (O_20,N_28972,N_28794);
or UO_21 (O_21,N_28988,N_28515);
nor UO_22 (O_22,N_28790,N_28657);
xor UO_23 (O_23,N_29757,N_28637);
or UO_24 (O_24,N_29047,N_29977);
and UO_25 (O_25,N_29265,N_29992);
nand UO_26 (O_26,N_29383,N_29475);
nor UO_27 (O_27,N_29876,N_29426);
nor UO_28 (O_28,N_28853,N_28712);
xnor UO_29 (O_29,N_28773,N_29463);
xnor UO_30 (O_30,N_29141,N_29187);
xor UO_31 (O_31,N_28930,N_29457);
nor UO_32 (O_32,N_29100,N_29888);
xor UO_33 (O_33,N_29201,N_28691);
nand UO_34 (O_34,N_29202,N_28513);
nor UO_35 (O_35,N_29021,N_29550);
and UO_36 (O_36,N_29792,N_28592);
xnor UO_37 (O_37,N_29957,N_28888);
nor UO_38 (O_38,N_29313,N_29337);
and UO_39 (O_39,N_29259,N_29543);
nor UO_40 (O_40,N_29508,N_28617);
and UO_41 (O_41,N_28814,N_29401);
and UO_42 (O_42,N_29079,N_28524);
nor UO_43 (O_43,N_29150,N_29040);
nor UO_44 (O_44,N_29767,N_29591);
and UO_45 (O_45,N_29573,N_29518);
and UO_46 (O_46,N_29737,N_29618);
and UO_47 (O_47,N_29178,N_29814);
xor UO_48 (O_48,N_28537,N_29903);
nor UO_49 (O_49,N_28650,N_29617);
nand UO_50 (O_50,N_29430,N_28805);
nor UO_51 (O_51,N_28571,N_29722);
or UO_52 (O_52,N_29524,N_29700);
nor UO_53 (O_53,N_29820,N_28865);
nor UO_54 (O_54,N_29651,N_29413);
and UO_55 (O_55,N_29760,N_29717);
nand UO_56 (O_56,N_29723,N_29061);
or UO_57 (O_57,N_29776,N_29323);
xor UO_58 (O_58,N_29827,N_29583);
nand UO_59 (O_59,N_29500,N_28858);
and UO_60 (O_60,N_29721,N_29248);
and UO_61 (O_61,N_29212,N_29387);
nand UO_62 (O_62,N_29262,N_29836);
xnor UO_63 (O_63,N_28569,N_29729);
nor UO_64 (O_64,N_28742,N_28829);
or UO_65 (O_65,N_29111,N_29215);
nand UO_66 (O_66,N_29185,N_28683);
nor UO_67 (O_67,N_28655,N_29319);
nand UO_68 (O_68,N_28785,N_28968);
nand UO_69 (O_69,N_29764,N_29177);
and UO_70 (O_70,N_29606,N_28931);
and UO_71 (O_71,N_28594,N_28799);
nand UO_72 (O_72,N_29143,N_28653);
nor UO_73 (O_73,N_29740,N_28603);
or UO_74 (O_74,N_29848,N_29235);
xor UO_75 (O_75,N_28900,N_29639);
and UO_76 (O_76,N_29445,N_29514);
nand UO_77 (O_77,N_29902,N_28539);
and UO_78 (O_78,N_29347,N_29364);
nor UO_79 (O_79,N_28574,N_29277);
nor UO_80 (O_80,N_29861,N_29266);
xnor UO_81 (O_81,N_28693,N_29419);
nor UO_82 (O_82,N_29522,N_29412);
or UO_83 (O_83,N_29844,N_28516);
or UO_84 (O_84,N_28743,N_28694);
or UO_85 (O_85,N_29123,N_28964);
and UO_86 (O_86,N_29440,N_29691);
nor UO_87 (O_87,N_29711,N_28656);
nand UO_88 (O_88,N_28620,N_29492);
nand UO_89 (O_89,N_29439,N_29746);
nor UO_90 (O_90,N_28784,N_29136);
and UO_91 (O_91,N_28767,N_29483);
xor UO_92 (O_92,N_29520,N_29288);
or UO_93 (O_93,N_29054,N_29164);
nand UO_94 (O_94,N_29211,N_28837);
nor UO_95 (O_95,N_28555,N_28976);
nor UO_96 (O_96,N_29709,N_29418);
nand UO_97 (O_97,N_28764,N_29554);
xnor UO_98 (O_98,N_29636,N_29166);
nand UO_99 (O_99,N_28669,N_29728);
xnor UO_100 (O_100,N_29829,N_29513);
and UO_101 (O_101,N_29042,N_29547);
and UO_102 (O_102,N_29001,N_29415);
xnor UO_103 (O_103,N_29218,N_28591);
or UO_104 (O_104,N_28749,N_29798);
nand UO_105 (O_105,N_29952,N_29605);
nand UO_106 (O_106,N_28720,N_29112);
or UO_107 (O_107,N_29945,N_29727);
nand UO_108 (O_108,N_28943,N_28827);
nand UO_109 (O_109,N_29470,N_29188);
nor UO_110 (O_110,N_28938,N_28604);
and UO_111 (O_111,N_29135,N_29803);
nand UO_112 (O_112,N_29568,N_29104);
nor UO_113 (O_113,N_29595,N_29494);
and UO_114 (O_114,N_29748,N_29693);
or UO_115 (O_115,N_29102,N_29255);
nor UO_116 (O_116,N_29015,N_29065);
nor UO_117 (O_117,N_29237,N_29134);
xnor UO_118 (O_118,N_29147,N_29264);
and UO_119 (O_119,N_28692,N_29207);
and UO_120 (O_120,N_29790,N_29738);
or UO_121 (O_121,N_29481,N_29159);
and UO_122 (O_122,N_29250,N_29390);
xnor UO_123 (O_123,N_28768,N_29022);
or UO_124 (O_124,N_29537,N_29299);
and UO_125 (O_125,N_29535,N_28697);
nand UO_126 (O_126,N_29630,N_29460);
nor UO_127 (O_127,N_28601,N_29400);
or UO_128 (O_128,N_28662,N_28889);
nor UO_129 (O_129,N_28946,N_29261);
xor UO_130 (O_130,N_29485,N_29742);
nand UO_131 (O_131,N_29502,N_29446);
and UO_132 (O_132,N_29824,N_28651);
and UO_133 (O_133,N_29466,N_29916);
nor UO_134 (O_134,N_28917,N_28748);
xor UO_135 (O_135,N_28899,N_28991);
nand UO_136 (O_136,N_29257,N_29887);
nand UO_137 (O_137,N_28675,N_29296);
nor UO_138 (O_138,N_29167,N_29113);
nand UO_139 (O_139,N_29358,N_28965);
nor UO_140 (O_140,N_28845,N_28672);
xor UO_141 (O_141,N_29090,N_29582);
or UO_142 (O_142,N_29231,N_28873);
nand UO_143 (O_143,N_28618,N_29733);
and UO_144 (O_144,N_29956,N_28772);
or UO_145 (O_145,N_29091,N_28820);
nor UO_146 (O_146,N_29777,N_29804);
xnor UO_147 (O_147,N_29025,N_29766);
nand UO_148 (O_148,N_29105,N_29063);
or UO_149 (O_149,N_28998,N_28685);
nor UO_150 (O_150,N_29145,N_28817);
nand UO_151 (O_151,N_28607,N_29971);
xor UO_152 (O_152,N_29856,N_29851);
nor UO_153 (O_153,N_29119,N_28734);
xnor UO_154 (O_154,N_29769,N_28925);
or UO_155 (O_155,N_29469,N_28831);
and UO_156 (O_156,N_29074,N_29673);
nand UO_157 (O_157,N_29230,N_28560);
and UO_158 (O_158,N_29566,N_29454);
and UO_159 (O_159,N_29110,N_28735);
or UO_160 (O_160,N_28954,N_29768);
nor UO_161 (O_161,N_29894,N_29677);
nor UO_162 (O_162,N_29515,N_28568);
nor UO_163 (O_163,N_29155,N_28680);
or UO_164 (O_164,N_28690,N_28652);
nand UO_165 (O_165,N_28920,N_29208);
or UO_166 (O_166,N_29689,N_29871);
xnor UO_167 (O_167,N_29072,N_29997);
nand UO_168 (O_168,N_29930,N_29396);
nor UO_169 (O_169,N_29958,N_29819);
or UO_170 (O_170,N_28544,N_29149);
nand UO_171 (O_171,N_29509,N_29756);
and UO_172 (O_172,N_29101,N_28564);
or UO_173 (O_173,N_29172,N_29785);
xor UO_174 (O_174,N_28957,N_29256);
or UO_175 (O_175,N_29254,N_28895);
and UO_176 (O_176,N_29642,N_29908);
xnor UO_177 (O_177,N_29650,N_29459);
xor UO_178 (O_178,N_29750,N_28953);
nand UO_179 (O_179,N_29708,N_28987);
xnor UO_180 (O_180,N_29374,N_29596);
or UO_181 (O_181,N_29986,N_28638);
nand UO_182 (O_182,N_28950,N_28769);
nand UO_183 (O_183,N_29773,N_29089);
nand UO_184 (O_184,N_28534,N_29562);
or UO_185 (O_185,N_29245,N_28870);
nand UO_186 (O_186,N_29555,N_29823);
nor UO_187 (O_187,N_29234,N_28684);
nor UO_188 (O_188,N_29778,N_29095);
xor UO_189 (O_189,N_29238,N_29758);
nand UO_190 (O_190,N_29783,N_28891);
or UO_191 (O_191,N_29282,N_28632);
nor UO_192 (O_192,N_28924,N_28506);
or UO_193 (O_193,N_28867,N_29954);
xnor UO_194 (O_194,N_28762,N_29306);
or UO_195 (O_195,N_29205,N_29959);
and UO_196 (O_196,N_29420,N_28782);
xor UO_197 (O_197,N_29716,N_29525);
nand UO_198 (O_198,N_29909,N_29027);
nand UO_199 (O_199,N_29923,N_28802);
and UO_200 (O_200,N_29637,N_29870);
or UO_201 (O_201,N_29246,N_28885);
and UO_202 (O_202,N_29668,N_29542);
nor UO_203 (O_203,N_29911,N_29927);
xnor UO_204 (O_204,N_29682,N_28877);
nand UO_205 (O_205,N_29796,N_29528);
nor UO_206 (O_206,N_28812,N_28741);
and UO_207 (O_207,N_29098,N_28583);
nand UO_208 (O_208,N_29322,N_28951);
and UO_209 (O_209,N_28630,N_29532);
and UO_210 (O_210,N_29627,N_29654);
nand UO_211 (O_211,N_29278,N_29204);
nor UO_212 (O_212,N_29477,N_29701);
nor UO_213 (O_213,N_29375,N_29464);
xor UO_214 (O_214,N_29395,N_29991);
or UO_215 (O_215,N_29842,N_29519);
nor UO_216 (O_216,N_29381,N_29160);
xnor UO_217 (O_217,N_29125,N_29441);
nor UO_218 (O_218,N_28860,N_28597);
or UO_219 (O_219,N_29036,N_29132);
and UO_220 (O_220,N_28578,N_29697);
and UO_221 (O_221,N_29601,N_29372);
nand UO_222 (O_222,N_29191,N_29094);
nor UO_223 (O_223,N_29226,N_29540);
nand UO_224 (O_224,N_28966,N_28708);
nor UO_225 (O_225,N_29023,N_28822);
nand UO_226 (O_226,N_29996,N_29116);
nand UO_227 (O_227,N_29019,N_29696);
or UO_228 (O_228,N_29153,N_29608);
xor UO_229 (O_229,N_28626,N_29781);
nand UO_230 (O_230,N_28777,N_29807);
nand UO_231 (O_231,N_28908,N_29498);
nand UO_232 (O_232,N_28786,N_29588);
nand UO_233 (O_233,N_28557,N_28766);
nor UO_234 (O_234,N_29391,N_29165);
xor UO_235 (O_235,N_29359,N_29484);
or UO_236 (O_236,N_29973,N_28960);
nor UO_237 (O_237,N_29070,N_29735);
and UO_238 (O_238,N_29180,N_29526);
or UO_239 (O_239,N_29895,N_29942);
or UO_240 (O_240,N_28902,N_28509);
or UO_241 (O_241,N_29886,N_29676);
xnor UO_242 (O_242,N_29915,N_29645);
nor UO_243 (O_243,N_29698,N_28781);
nand UO_244 (O_244,N_29142,N_29013);
and UO_245 (O_245,N_29144,N_29099);
nor UO_246 (O_246,N_29043,N_28973);
nor UO_247 (O_247,N_29718,N_28566);
or UO_248 (O_248,N_28824,N_28956);
and UO_249 (O_249,N_29813,N_28575);
xnor UO_250 (O_250,N_28756,N_29663);
nand UO_251 (O_251,N_28563,N_28737);
and UO_252 (O_252,N_29799,N_28505);
and UO_253 (O_253,N_29397,N_29613);
nand UO_254 (O_254,N_28722,N_29073);
nor UO_255 (O_255,N_28702,N_28818);
nand UO_256 (O_256,N_29633,N_29967);
nand UO_257 (O_257,N_28989,N_29569);
or UO_258 (O_258,N_29103,N_29703);
and UO_259 (O_259,N_28811,N_29152);
or UO_260 (O_260,N_28542,N_29731);
and UO_261 (O_261,N_29068,N_28726);
nand UO_262 (O_262,N_28587,N_28979);
or UO_263 (O_263,N_28934,N_28952);
and UO_264 (O_264,N_29066,N_28647);
xnor UO_265 (O_265,N_29978,N_29239);
nor UO_266 (O_266,N_29563,N_29121);
xor UO_267 (O_267,N_29117,N_29922);
xor UO_268 (O_268,N_28990,N_29310);
nor UO_269 (O_269,N_28501,N_29548);
nand UO_270 (O_270,N_29897,N_29406);
xnor UO_271 (O_271,N_28992,N_28752);
nand UO_272 (O_272,N_29096,N_28840);
nand UO_273 (O_273,N_28945,N_28670);
nand UO_274 (O_274,N_29051,N_28668);
xnor UO_275 (O_275,N_29744,N_29329);
nor UO_276 (O_276,N_29516,N_29821);
nor UO_277 (O_277,N_28919,N_29879);
nand UO_278 (O_278,N_29539,N_28775);
or UO_279 (O_279,N_29402,N_29864);
xnor UO_280 (O_280,N_29362,N_28529);
and UO_281 (O_281,N_28518,N_29085);
and UO_282 (O_282,N_29683,N_29182);
nand UO_283 (O_283,N_29295,N_28793);
xnor UO_284 (O_284,N_28703,N_29724);
or UO_285 (O_285,N_29369,N_28755);
and UO_286 (O_286,N_29770,N_29702);
xnor UO_287 (O_287,N_28549,N_29884);
nor UO_288 (O_288,N_29904,N_28798);
nand UO_289 (O_289,N_29765,N_28730);
nand UO_290 (O_290,N_28881,N_29268);
and UO_291 (O_291,N_29292,N_29126);
or UO_292 (O_292,N_29855,N_28526);
and UO_293 (O_293,N_28532,N_29062);
nor UO_294 (O_294,N_29340,N_28654);
nor UO_295 (O_295,N_28584,N_29538);
xnor UO_296 (O_296,N_28646,N_29416);
or UO_297 (O_297,N_29789,N_29473);
nand UO_298 (O_298,N_29055,N_29148);
xor UO_299 (O_299,N_29567,N_29564);
and UO_300 (O_300,N_28796,N_28678);
xor UO_301 (O_301,N_28875,N_29603);
or UO_302 (O_302,N_29199,N_29384);
nand UO_303 (O_303,N_29556,N_29679);
xnor UO_304 (O_304,N_29108,N_29623);
and UO_305 (O_305,N_29086,N_29328);
nand UO_306 (O_306,N_29106,N_29124);
and UO_307 (O_307,N_28771,N_28750);
xnor UO_308 (O_308,N_29570,N_28792);
nor UO_309 (O_309,N_28510,N_28579);
nor UO_310 (O_310,N_29410,N_29671);
and UO_311 (O_311,N_28589,N_28971);
nand UO_312 (O_312,N_29414,N_29423);
nand UO_313 (O_313,N_29726,N_28547);
nand UO_314 (O_314,N_29429,N_29417);
nand UO_315 (O_315,N_28746,N_28927);
xnor UO_316 (O_316,N_28665,N_29482);
nor UO_317 (O_317,N_28800,N_28942);
nand UO_318 (O_318,N_29133,N_28779);
xor UO_319 (O_319,N_29961,N_29840);
nand UO_320 (O_320,N_29236,N_29808);
or UO_321 (O_321,N_29694,N_28522);
nand UO_322 (O_322,N_29326,N_29946);
and UO_323 (O_323,N_29593,N_29011);
nor UO_324 (O_324,N_29780,N_28580);
or UO_325 (O_325,N_29962,N_29646);
and UO_326 (O_326,N_28525,N_29734);
and UO_327 (O_327,N_29291,N_29267);
nor UO_328 (O_328,N_29438,N_28819);
xor UO_329 (O_329,N_29233,N_29880);
xor UO_330 (O_330,N_29488,N_29467);
nand UO_331 (O_331,N_28562,N_29343);
and UO_332 (O_332,N_28548,N_29975);
xnor UO_333 (O_333,N_28770,N_28725);
and UO_334 (O_334,N_29404,N_28641);
or UO_335 (O_335,N_28883,N_29589);
xor UO_336 (O_336,N_28958,N_29604);
nor UO_337 (O_337,N_28649,N_28761);
and UO_338 (O_338,N_29157,N_29658);
and UO_339 (O_339,N_29356,N_29759);
or UO_340 (O_340,N_28713,N_28842);
nor UO_341 (O_341,N_29951,N_29355);
nor UO_342 (O_342,N_29752,N_29209);
nand UO_343 (O_343,N_28520,N_29293);
xor UO_344 (O_344,N_28633,N_29028);
or UO_345 (O_345,N_29504,N_29629);
nand UO_346 (O_346,N_28984,N_29704);
or UO_347 (O_347,N_29219,N_28558);
xnor UO_348 (O_348,N_28606,N_29656);
nand UO_349 (O_349,N_28612,N_29719);
or UO_350 (O_350,N_29932,N_29712);
nand UO_351 (O_351,N_29580,N_29558);
or UO_352 (O_352,N_29998,N_28795);
nor UO_353 (O_353,N_29379,N_29739);
nor UO_354 (O_354,N_28705,N_29680);
nor UO_355 (O_355,N_29076,N_28977);
nand UO_356 (O_356,N_28622,N_29016);
or UO_357 (O_357,N_29316,N_28826);
xnor UO_358 (O_358,N_29869,N_29812);
and UO_359 (O_359,N_28839,N_28538);
and UO_360 (O_360,N_29003,N_29393);
or UO_361 (O_361,N_28789,N_29139);
nand UO_362 (O_362,N_29811,N_28573);
nand UO_363 (O_363,N_29317,N_28724);
nand UO_364 (O_364,N_28944,N_29619);
xnor UO_365 (O_365,N_29411,N_29649);
or UO_366 (O_366,N_29044,N_28871);
xor UO_367 (O_367,N_28545,N_29963);
nand UO_368 (O_368,N_29553,N_28846);
and UO_369 (O_369,N_28745,N_29622);
xor UO_370 (O_370,N_29499,N_29928);
nand UO_371 (O_371,N_28928,N_28704);
and UO_372 (O_372,N_29640,N_29859);
nand UO_373 (O_373,N_29747,N_29779);
and UO_374 (O_374,N_29156,N_28914);
nor UO_375 (O_375,N_28503,N_28980);
and UO_376 (O_376,N_28803,N_28936);
nand UO_377 (O_377,N_29109,N_28540);
xor UO_378 (O_378,N_28611,N_28648);
xor UO_379 (O_379,N_29787,N_29331);
nor UO_380 (O_380,N_28816,N_28874);
nand UO_381 (O_381,N_29286,N_28898);
or UO_382 (O_382,N_29632,N_29217);
xor UO_383 (O_383,N_29660,N_28915);
or UO_384 (O_384,N_29223,N_29349);
and UO_385 (O_385,N_29966,N_29900);
nand UO_386 (O_386,N_28869,N_28729);
nand UO_387 (O_387,N_29453,N_29269);
or UO_388 (O_388,N_29800,N_29877);
and UO_389 (O_389,N_29652,N_29885);
xor UO_390 (O_390,N_29339,N_29363);
xor UO_391 (O_391,N_29577,N_29382);
nor UO_392 (O_392,N_28955,N_28774);
or UO_393 (O_393,N_29635,N_29491);
or UO_394 (O_394,N_29969,N_28906);
nand UO_395 (O_395,N_29449,N_29373);
and UO_396 (O_396,N_28535,N_29127);
nor UO_397 (O_397,N_29592,N_29093);
xnor UO_398 (O_398,N_29872,N_29881);
and UO_399 (O_399,N_28500,N_28602);
nand UO_400 (O_400,N_29817,N_29594);
or UO_401 (O_401,N_29533,N_28610);
or UO_402 (O_402,N_28504,N_29692);
nand UO_403 (O_403,N_28507,N_29118);
or UO_404 (O_404,N_29444,N_28673);
or UO_405 (O_405,N_29487,N_29545);
xor UO_406 (O_406,N_29490,N_28689);
nand UO_407 (O_407,N_29338,N_28577);
or UO_408 (O_408,N_28760,N_29838);
xor UO_409 (O_409,N_29621,N_28905);
xor UO_410 (O_410,N_28517,N_28614);
or UO_411 (O_411,N_28896,N_29049);
or UO_412 (O_412,N_29981,N_28797);
or UO_413 (O_413,N_29984,N_28975);
or UO_414 (O_414,N_29544,N_29270);
and UO_415 (O_415,N_28808,N_29541);
or UO_416 (O_416,N_28884,N_28996);
nand UO_417 (O_417,N_29882,N_29301);
xnor UO_418 (O_418,N_29643,N_29140);
or UO_419 (O_419,N_29610,N_28995);
and UO_420 (O_420,N_29120,N_28961);
xnor UO_421 (O_421,N_29240,N_29834);
nor UO_422 (O_422,N_28728,N_28894);
and UO_423 (O_423,N_28595,N_29321);
xor UO_424 (O_424,N_29875,N_29324);
nand UO_425 (O_425,N_29989,N_29389);
and UO_426 (O_426,N_29297,N_28857);
and UO_427 (O_427,N_28864,N_28872);
xor UO_428 (O_428,N_29392,N_29368);
nor UO_429 (O_429,N_29950,N_29122);
or UO_430 (O_430,N_29581,N_29910);
xor UO_431 (O_431,N_28994,N_29181);
and UO_432 (O_432,N_29598,N_29536);
or UO_433 (O_433,N_29653,N_29081);
nor UO_434 (O_434,N_28901,N_29276);
and UO_435 (O_435,N_29354,N_28736);
xor UO_436 (O_436,N_29987,N_29751);
or UO_437 (O_437,N_29468,N_29826);
or UO_438 (O_438,N_28682,N_29743);
and UO_439 (O_439,N_28974,N_29931);
and UO_440 (O_440,N_28791,N_28834);
xor UO_441 (O_441,N_29786,N_29380);
nor UO_442 (O_442,N_28727,N_28658);
xor UO_443 (O_443,N_29560,N_29071);
or UO_444 (O_444,N_29847,N_28776);
nor UO_445 (O_445,N_28502,N_28939);
nor UO_446 (O_446,N_28629,N_29045);
xnor UO_447 (O_447,N_29559,N_29995);
xor UO_448 (O_448,N_29920,N_28903);
nand UO_449 (O_449,N_29284,N_28986);
and UO_450 (O_450,N_29912,N_29549);
nor UO_451 (O_451,N_29597,N_29599);
and UO_452 (O_452,N_28838,N_28861);
nand UO_453 (O_453,N_29833,N_29398);
nor UO_454 (O_454,N_29082,N_29529);
xnor UO_455 (O_455,N_29273,N_28759);
and UO_456 (O_456,N_29422,N_29341);
nor UO_457 (O_457,N_29213,N_28556);
nor UO_458 (O_458,N_29575,N_29059);
xnor UO_459 (O_459,N_29281,N_29868);
nor UO_460 (O_460,N_29784,N_28941);
nor UO_461 (O_461,N_29258,N_28581);
or UO_462 (O_462,N_28847,N_29046);
or UO_463 (O_463,N_29190,N_29788);
and UO_464 (O_464,N_29131,N_28598);
or UO_465 (O_465,N_29688,N_29590);
nor UO_466 (O_466,N_29456,N_29452);
and UO_467 (O_467,N_29004,N_29020);
xnor UO_468 (O_468,N_29512,N_29993);
or UO_469 (O_469,N_29644,N_28600);
nand UO_470 (O_470,N_29587,N_29706);
nor UO_471 (O_471,N_29137,N_28863);
xor UO_472 (O_472,N_29741,N_28893);
and UO_473 (O_473,N_28747,N_28681);
and UO_474 (O_474,N_29304,N_29705);
or UO_475 (O_475,N_28830,N_29053);
and UO_476 (O_476,N_29489,N_28688);
or UO_477 (O_477,N_29667,N_29432);
nand UO_478 (O_478,N_28911,N_29818);
and UO_479 (O_479,N_28859,N_29243);
xor UO_480 (O_480,N_28644,N_29290);
nand UO_481 (O_481,N_29092,N_29849);
nor UO_482 (O_482,N_28699,N_29229);
or UO_483 (O_483,N_28719,N_29831);
nor UO_484 (O_484,N_28572,N_29203);
xnor UO_485 (O_485,N_29707,N_29616);
and UO_486 (O_486,N_28621,N_29303);
or UO_487 (O_487,N_29315,N_28530);
nand UO_488 (O_488,N_29858,N_29405);
xnor UO_489 (O_489,N_29039,N_29307);
and UO_490 (O_490,N_28854,N_29365);
nor UO_491 (O_491,N_28868,N_28666);
nand UO_492 (O_492,N_29947,N_28567);
xnor UO_493 (O_493,N_28663,N_28970);
or UO_494 (O_494,N_29672,N_29274);
or UO_495 (O_495,N_29018,N_29351);
xnor UO_496 (O_496,N_29346,N_28778);
and UO_497 (O_497,N_29797,N_29574);
xnor UO_498 (O_498,N_28753,N_28616);
and UO_499 (O_499,N_29161,N_28821);
nor UO_500 (O_500,N_28848,N_29360);
nand UO_501 (O_501,N_29129,N_29761);
nor UO_502 (O_502,N_28922,N_28907);
xnor UO_503 (O_503,N_28933,N_28586);
or UO_504 (O_504,N_28686,N_29496);
and UO_505 (O_505,N_29480,N_29227);
and UO_506 (O_506,N_29087,N_29710);
nand UO_507 (O_507,N_28721,N_29151);
or UO_508 (O_508,N_28765,N_29546);
or UO_509 (O_509,N_28758,N_29745);
xor UO_510 (O_510,N_29699,N_29377);
nor UO_511 (O_511,N_29486,N_28851);
nor UO_512 (O_512,N_28751,N_29447);
nand UO_513 (O_513,N_28576,N_28718);
xnor UO_514 (O_514,N_29352,N_28552);
nor UO_515 (O_515,N_29980,N_29195);
nor UO_516 (O_516,N_29925,N_29376);
xnor UO_517 (O_517,N_29919,N_28615);
nand UO_518 (O_518,N_28605,N_29999);
nor UO_519 (O_519,N_29763,N_29000);
and UO_520 (O_520,N_28613,N_28862);
xnor UO_521 (O_521,N_29057,N_29625);
nand UO_522 (O_522,N_29853,N_29584);
nand UO_523 (O_523,N_28643,N_29732);
nor UO_524 (O_524,N_28850,N_29184);
or UO_525 (O_525,N_29241,N_29953);
or UO_526 (O_526,N_29175,N_29918);
nand UO_527 (O_527,N_29200,N_29448);
or UO_528 (O_528,N_29664,N_29899);
nand UO_529 (O_529,N_29399,N_28921);
and UO_530 (O_530,N_29451,N_28588);
xor UO_531 (O_531,N_28533,N_29041);
nand UO_532 (O_532,N_28787,N_29913);
nor UO_533 (O_533,N_29822,N_29442);
xnor UO_534 (O_534,N_29576,N_28809);
and UO_535 (O_535,N_29662,N_29348);
and UO_536 (O_536,N_29865,N_29366);
and UO_537 (O_537,N_29736,N_28948);
xor UO_538 (O_538,N_29852,N_29158);
and UO_539 (O_539,N_29408,N_28739);
or UO_540 (O_540,N_29435,N_29183);
or UO_541 (O_541,N_29551,N_28892);
xor UO_542 (O_542,N_28886,N_29948);
and UO_543 (O_543,N_29907,N_28959);
or UO_544 (O_544,N_29050,N_29631);
or UO_545 (O_545,N_29607,N_28937);
nor UO_546 (O_546,N_29163,N_28590);
or UO_547 (O_547,N_28897,N_29114);
or UO_548 (O_548,N_28608,N_29171);
nor UO_549 (O_549,N_29421,N_29225);
nor UO_550 (O_550,N_29138,N_29889);
xnor UO_551 (O_551,N_28570,N_29353);
nor UO_552 (O_552,N_29837,N_29505);
or UO_553 (O_553,N_29774,N_29394);
nor UO_554 (O_554,N_29517,N_29600);
nand UO_555 (O_555,N_29146,N_29333);
nor UO_556 (O_556,N_29320,N_29507);
xor UO_557 (O_557,N_28660,N_28625);
xor UO_558 (O_558,N_29810,N_29674);
xnor UO_559 (O_559,N_29263,N_29921);
nor UO_560 (O_560,N_28536,N_28833);
xnor UO_561 (O_561,N_29906,N_29450);
xnor UO_562 (O_562,N_28940,N_29370);
nand UO_563 (O_563,N_29965,N_29988);
and UO_564 (O_564,N_29495,N_29194);
and UO_565 (O_565,N_29431,N_29771);
nand UO_566 (O_566,N_29843,N_28754);
nand UO_567 (O_567,N_29222,N_29893);
and UO_568 (O_568,N_29655,N_28947);
or UO_569 (O_569,N_29403,N_28910);
nand UO_570 (O_570,N_29060,N_28828);
xnor UO_571 (O_571,N_28543,N_29534);
xnor UO_572 (O_572,N_28631,N_29816);
nor UO_573 (O_573,N_28963,N_29472);
or UO_574 (O_574,N_28904,N_28981);
nand UO_575 (O_575,N_28627,N_28807);
nand UO_576 (O_576,N_29300,N_29247);
nor UO_577 (O_577,N_29260,N_29192);
nor UO_578 (O_578,N_29064,N_29294);
xnor UO_579 (O_579,N_29898,N_28935);
xnor UO_580 (O_580,N_29944,N_28671);
xor UO_581 (O_581,N_29896,N_29943);
and UO_582 (O_582,N_29857,N_29221);
nand UO_583 (O_583,N_29762,N_28523);
nand UO_584 (O_584,N_29309,N_28551);
and UO_585 (O_585,N_29078,N_28528);
or UO_586 (O_586,N_29579,N_29198);
nor UO_587 (O_587,N_28582,N_29657);
nand UO_588 (O_588,N_28593,N_28836);
nand UO_589 (O_589,N_29361,N_28855);
nand UO_590 (O_590,N_29176,N_28744);
nand UO_591 (O_591,N_28926,N_28823);
and UO_592 (O_592,N_29791,N_29461);
nand UO_593 (O_593,N_28710,N_28674);
xor UO_594 (O_594,N_29478,N_29990);
nor UO_595 (O_595,N_28695,N_29252);
xnor UO_596 (O_596,N_29424,N_28890);
nand UO_597 (O_597,N_28932,N_29835);
nand UO_598 (O_598,N_29285,N_29845);
or UO_599 (O_599,N_29873,N_29690);
nand UO_600 (O_600,N_28554,N_29012);
or UO_601 (O_601,N_29620,N_29612);
nor UO_602 (O_602,N_29860,N_28740);
nand UO_603 (O_603,N_29002,N_29433);
xor UO_604 (O_604,N_28978,N_29941);
nand UO_605 (O_605,N_29029,N_28561);
nor UO_606 (O_606,N_29960,N_29034);
xor UO_607 (O_607,N_28531,N_29890);
nor UO_608 (O_608,N_29327,N_28715);
xor UO_609 (O_609,N_29686,N_29305);
nor UO_610 (O_610,N_28806,N_29010);
or UO_611 (O_611,N_28599,N_29052);
xor UO_612 (O_612,N_29527,N_29815);
or UO_613 (O_613,N_28882,N_29170);
or UO_614 (O_614,N_29972,N_29224);
nor UO_615 (O_615,N_29196,N_29867);
xnor UO_616 (O_616,N_29249,N_29455);
xor UO_617 (O_617,N_29841,N_28832);
or UO_618 (O_618,N_29883,N_29775);
nor UO_619 (O_619,N_29901,N_29030);
or UO_620 (O_620,N_29929,N_28804);
and UO_621 (O_621,N_29314,N_29611);
nand UO_622 (O_622,N_29964,N_29854);
nor UO_623 (O_623,N_28923,N_29067);
and UO_624 (O_624,N_28733,N_29024);
nor UO_625 (O_625,N_29189,N_29298);
or UO_626 (O_626,N_28519,N_28701);
nor UO_627 (O_627,N_29056,N_29275);
or UO_628 (O_628,N_29279,N_29939);
nor UO_629 (O_629,N_28619,N_29795);
or UO_630 (O_630,N_28844,N_29714);
nand UO_631 (O_631,N_28912,N_29678);
xor UO_632 (O_632,N_28596,N_29008);
xor UO_633 (O_633,N_29685,N_29128);
and UO_634 (O_634,N_28559,N_29130);
or UO_635 (O_635,N_29378,N_28514);
xor UO_636 (O_636,N_28635,N_29609);
nand UO_637 (O_637,N_29497,N_29586);
xor UO_638 (O_638,N_29006,N_28876);
xor UO_639 (O_639,N_29501,N_28661);
nand UO_640 (O_640,N_29940,N_29557);
and UO_641 (O_641,N_28763,N_29026);
xor UO_642 (O_642,N_29465,N_29511);
and UO_643 (O_643,N_28546,N_29007);
or UO_644 (O_644,N_29471,N_29214);
or UO_645 (O_645,N_29210,N_29443);
xnor UO_646 (O_646,N_28717,N_28879);
xnor UO_647 (O_647,N_28640,N_29830);
or UO_648 (O_648,N_29713,N_29661);
nor UO_649 (O_649,N_28801,N_29179);
or UO_650 (O_650,N_28636,N_28856);
nor UO_651 (O_651,N_29968,N_29794);
nand UO_652 (O_652,N_29174,N_29107);
xor UO_653 (O_653,N_29648,N_29335);
nor UO_654 (O_654,N_29615,N_29846);
xnor UO_655 (O_655,N_29917,N_29017);
nand UO_656 (O_656,N_28985,N_29162);
xnor UO_657 (O_657,N_29069,N_29436);
nand UO_658 (O_658,N_29659,N_28841);
or UO_659 (O_659,N_29572,N_28679);
nand UO_660 (O_660,N_29531,N_28993);
and UO_661 (O_661,N_28813,N_29585);
xnor UO_662 (O_662,N_28788,N_29949);
nor UO_663 (O_663,N_29924,N_29173);
nor UO_664 (O_664,N_29216,N_29985);
xnor UO_665 (O_665,N_29206,N_29749);
nand UO_666 (O_666,N_29628,N_29220);
or UO_667 (O_667,N_29311,N_28709);
nand UO_668 (O_668,N_29937,N_28512);
and UO_669 (O_669,N_28949,N_29232);
nor UO_670 (O_670,N_28916,N_29325);
and UO_671 (O_671,N_29251,N_28810);
or UO_672 (O_672,N_29983,N_29825);
or UO_673 (O_673,N_29641,N_29345);
or UO_674 (O_674,N_29832,N_28553);
xor UO_675 (O_675,N_29334,N_28815);
xnor UO_676 (O_676,N_29115,N_28835);
xnor UO_677 (O_677,N_29048,N_29938);
nor UO_678 (O_678,N_28659,N_29350);
and UO_679 (O_679,N_29506,N_29695);
or UO_680 (O_680,N_28967,N_28711);
or UO_681 (O_681,N_28624,N_28918);
nand UO_682 (O_682,N_28723,N_28639);
or UO_683 (O_683,N_29982,N_29458);
and UO_684 (O_684,N_28999,N_29754);
and UO_685 (O_685,N_28527,N_29552);
xor UO_686 (O_686,N_29675,N_29753);
and UO_687 (O_687,N_28707,N_29970);
nor UO_688 (O_688,N_29272,N_29687);
or UO_689 (O_689,N_28645,N_29154);
or UO_690 (O_690,N_29386,N_29462);
and UO_691 (O_691,N_28700,N_29388);
nor UO_692 (O_692,N_29614,N_29271);
and UO_693 (O_693,N_29084,N_29228);
or UO_694 (O_694,N_28780,N_29805);
nor UO_695 (O_695,N_29523,N_29344);
nor UO_696 (O_696,N_29097,N_28738);
xnor UO_697 (O_697,N_29669,N_28843);
and UO_698 (O_698,N_29866,N_29638);
xor UO_699 (O_699,N_29715,N_28887);
nand UO_700 (O_700,N_28982,N_28878);
or UO_701 (O_701,N_29493,N_29926);
xnor UO_702 (O_702,N_28585,N_29088);
nand UO_703 (O_703,N_29009,N_29730);
nand UO_704 (O_704,N_29755,N_29933);
nand UO_705 (O_705,N_29169,N_28731);
nor UO_706 (O_706,N_28714,N_28783);
nand UO_707 (O_707,N_29014,N_29578);
nor UO_708 (O_708,N_29892,N_29077);
and UO_709 (O_709,N_29647,N_29503);
xor UO_710 (O_710,N_29626,N_29530);
nor UO_711 (O_711,N_29974,N_29602);
and UO_712 (O_712,N_28541,N_29561);
nor UO_713 (O_713,N_28969,N_28521);
nor UO_714 (O_714,N_29425,N_29357);
xor UO_715 (O_715,N_29850,N_29725);
nor UO_716 (O_716,N_29684,N_29168);
nor UO_717 (O_717,N_28849,N_29934);
and UO_718 (O_718,N_29670,N_29914);
nand UO_719 (O_719,N_29474,N_29253);
or UO_720 (O_720,N_29828,N_29874);
xnor UO_721 (O_721,N_28667,N_28676);
or UO_722 (O_722,N_28634,N_29437);
or UO_723 (O_723,N_29032,N_28511);
nand UO_724 (O_724,N_28757,N_28698);
nand UO_725 (O_725,N_29772,N_28642);
or UO_726 (O_726,N_29976,N_28732);
nor UO_727 (O_727,N_29521,N_29809);
and UO_728 (O_728,N_29280,N_29863);
and UO_729 (O_729,N_29083,N_29936);
and UO_730 (O_730,N_28866,N_29434);
or UO_731 (O_731,N_29409,N_28929);
xnor UO_732 (O_732,N_29289,N_29839);
or UO_733 (O_733,N_29624,N_29038);
xor UO_734 (O_734,N_29665,N_28623);
or UO_735 (O_735,N_29720,N_29330);
or UO_736 (O_736,N_29080,N_29283);
nand UO_737 (O_737,N_29075,N_29035);
and UO_738 (O_738,N_28909,N_29332);
or UO_739 (O_739,N_29802,N_28628);
and UO_740 (O_740,N_29479,N_29302);
and UO_741 (O_741,N_28696,N_29476);
nand UO_742 (O_742,N_29862,N_28913);
nor UO_743 (O_743,N_28687,N_29336);
nand UO_744 (O_744,N_28825,N_29058);
nand UO_745 (O_745,N_29428,N_29033);
or UO_746 (O_746,N_29371,N_28565);
nand UO_747 (O_747,N_28983,N_29312);
and UO_748 (O_748,N_29407,N_28716);
nor UO_749 (O_749,N_28664,N_29891);
nor UO_750 (O_750,N_28829,N_29813);
nand UO_751 (O_751,N_29237,N_29882);
nand UO_752 (O_752,N_29831,N_29858);
xnor UO_753 (O_753,N_28984,N_29396);
nor UO_754 (O_754,N_29344,N_29911);
nor UO_755 (O_755,N_29416,N_29994);
and UO_756 (O_756,N_29002,N_28509);
and UO_757 (O_757,N_29667,N_28988);
nor UO_758 (O_758,N_28914,N_29516);
and UO_759 (O_759,N_29090,N_29332);
nand UO_760 (O_760,N_29741,N_29306);
or UO_761 (O_761,N_29629,N_29897);
nor UO_762 (O_762,N_29456,N_28960);
nor UO_763 (O_763,N_29732,N_29365);
and UO_764 (O_764,N_28630,N_29554);
nor UO_765 (O_765,N_28841,N_29692);
and UO_766 (O_766,N_29945,N_29157);
nand UO_767 (O_767,N_29555,N_29860);
nand UO_768 (O_768,N_29830,N_29106);
nand UO_769 (O_769,N_29056,N_29379);
xnor UO_770 (O_770,N_29886,N_29049);
or UO_771 (O_771,N_29162,N_29584);
nor UO_772 (O_772,N_29090,N_29652);
nor UO_773 (O_773,N_29689,N_29856);
or UO_774 (O_774,N_29526,N_28565);
xnor UO_775 (O_775,N_29325,N_29822);
xor UO_776 (O_776,N_29097,N_29922);
xor UO_777 (O_777,N_29721,N_29937);
or UO_778 (O_778,N_28789,N_29650);
nor UO_779 (O_779,N_29985,N_29313);
xnor UO_780 (O_780,N_28857,N_28728);
xnor UO_781 (O_781,N_29083,N_29571);
nand UO_782 (O_782,N_28529,N_29929);
or UO_783 (O_783,N_29016,N_29753);
xor UO_784 (O_784,N_29017,N_29279);
or UO_785 (O_785,N_28889,N_28519);
or UO_786 (O_786,N_28736,N_29848);
and UO_787 (O_787,N_28889,N_29390);
and UO_788 (O_788,N_29006,N_29236);
xnor UO_789 (O_789,N_28673,N_29377);
xnor UO_790 (O_790,N_29783,N_28843);
xor UO_791 (O_791,N_29645,N_28784);
nor UO_792 (O_792,N_29505,N_28597);
and UO_793 (O_793,N_29700,N_28688);
or UO_794 (O_794,N_29024,N_29502);
or UO_795 (O_795,N_28658,N_29511);
or UO_796 (O_796,N_29825,N_28542);
nor UO_797 (O_797,N_28695,N_28902);
or UO_798 (O_798,N_29849,N_29848);
nand UO_799 (O_799,N_29837,N_29653);
xnor UO_800 (O_800,N_28795,N_29121);
nand UO_801 (O_801,N_29032,N_29425);
nor UO_802 (O_802,N_28890,N_29294);
nand UO_803 (O_803,N_29860,N_29499);
or UO_804 (O_804,N_29196,N_29131);
and UO_805 (O_805,N_28583,N_28708);
nand UO_806 (O_806,N_28819,N_29565);
nand UO_807 (O_807,N_28925,N_29677);
nor UO_808 (O_808,N_29000,N_29372);
nor UO_809 (O_809,N_29534,N_29775);
nand UO_810 (O_810,N_29672,N_29269);
nand UO_811 (O_811,N_28938,N_29016);
or UO_812 (O_812,N_29035,N_29572);
xor UO_813 (O_813,N_28966,N_29391);
and UO_814 (O_814,N_29062,N_29119);
nand UO_815 (O_815,N_28915,N_28815);
nand UO_816 (O_816,N_29459,N_29161);
or UO_817 (O_817,N_29589,N_29428);
nor UO_818 (O_818,N_29229,N_29700);
nor UO_819 (O_819,N_29075,N_29896);
nor UO_820 (O_820,N_29584,N_29108);
nand UO_821 (O_821,N_28783,N_29747);
or UO_822 (O_822,N_28858,N_28566);
xnor UO_823 (O_823,N_29477,N_29913);
or UO_824 (O_824,N_29327,N_29387);
and UO_825 (O_825,N_29170,N_28616);
or UO_826 (O_826,N_28933,N_28581);
nand UO_827 (O_827,N_28516,N_29397);
and UO_828 (O_828,N_28671,N_29683);
nor UO_829 (O_829,N_28571,N_29226);
and UO_830 (O_830,N_28567,N_28953);
xor UO_831 (O_831,N_29259,N_29330);
xnor UO_832 (O_832,N_28727,N_29637);
and UO_833 (O_833,N_29602,N_29176);
nand UO_834 (O_834,N_29206,N_28547);
nand UO_835 (O_835,N_29981,N_28617);
and UO_836 (O_836,N_29444,N_29293);
xor UO_837 (O_837,N_29285,N_29167);
or UO_838 (O_838,N_28661,N_29726);
nand UO_839 (O_839,N_29365,N_29121);
or UO_840 (O_840,N_29798,N_29194);
nand UO_841 (O_841,N_28558,N_29018);
or UO_842 (O_842,N_28558,N_29311);
nand UO_843 (O_843,N_29938,N_29956);
xnor UO_844 (O_844,N_29767,N_29470);
nand UO_845 (O_845,N_28919,N_29722);
nand UO_846 (O_846,N_29648,N_29263);
and UO_847 (O_847,N_29160,N_29309);
nand UO_848 (O_848,N_28874,N_29411);
and UO_849 (O_849,N_29722,N_29078);
xor UO_850 (O_850,N_29800,N_28546);
xor UO_851 (O_851,N_29772,N_29340);
nor UO_852 (O_852,N_29026,N_29545);
nand UO_853 (O_853,N_29265,N_28737);
nor UO_854 (O_854,N_29516,N_29780);
or UO_855 (O_855,N_29065,N_28966);
nor UO_856 (O_856,N_29638,N_29803);
nand UO_857 (O_857,N_28704,N_28804);
nor UO_858 (O_858,N_28627,N_28590);
nor UO_859 (O_859,N_29044,N_29902);
and UO_860 (O_860,N_29088,N_29469);
nand UO_861 (O_861,N_29142,N_29682);
and UO_862 (O_862,N_29428,N_29104);
nor UO_863 (O_863,N_29784,N_29241);
or UO_864 (O_864,N_28633,N_29538);
xor UO_865 (O_865,N_29577,N_28522);
xnor UO_866 (O_866,N_28652,N_29234);
nand UO_867 (O_867,N_28604,N_29061);
and UO_868 (O_868,N_28500,N_29314);
nor UO_869 (O_869,N_28573,N_29398);
nand UO_870 (O_870,N_29402,N_28836);
nor UO_871 (O_871,N_28589,N_28948);
and UO_872 (O_872,N_28656,N_28881);
or UO_873 (O_873,N_28634,N_28968);
nor UO_874 (O_874,N_29054,N_29407);
xor UO_875 (O_875,N_29498,N_29527);
or UO_876 (O_876,N_29165,N_29328);
nor UO_877 (O_877,N_28761,N_28825);
nor UO_878 (O_878,N_29083,N_28575);
xor UO_879 (O_879,N_29350,N_29487);
nor UO_880 (O_880,N_29565,N_28885);
and UO_881 (O_881,N_28676,N_28897);
nor UO_882 (O_882,N_29623,N_29500);
xnor UO_883 (O_883,N_29886,N_29974);
or UO_884 (O_884,N_29258,N_29403);
nand UO_885 (O_885,N_29769,N_29677);
nand UO_886 (O_886,N_28557,N_28954);
nand UO_887 (O_887,N_29804,N_29166);
or UO_888 (O_888,N_29854,N_28728);
and UO_889 (O_889,N_29296,N_29083);
and UO_890 (O_890,N_29432,N_28719);
nand UO_891 (O_891,N_29496,N_29712);
or UO_892 (O_892,N_28913,N_28732);
and UO_893 (O_893,N_28581,N_29614);
and UO_894 (O_894,N_28651,N_29191);
nor UO_895 (O_895,N_29204,N_29993);
xnor UO_896 (O_896,N_29936,N_29846);
xnor UO_897 (O_897,N_29690,N_29364);
nand UO_898 (O_898,N_29300,N_28836);
xnor UO_899 (O_899,N_29256,N_29082);
xor UO_900 (O_900,N_29493,N_29337);
nand UO_901 (O_901,N_28744,N_29810);
or UO_902 (O_902,N_29215,N_29440);
nor UO_903 (O_903,N_29141,N_28841);
nand UO_904 (O_904,N_29110,N_28993);
or UO_905 (O_905,N_28989,N_29477);
and UO_906 (O_906,N_28941,N_29589);
nand UO_907 (O_907,N_29511,N_29328);
or UO_908 (O_908,N_29661,N_29796);
xnor UO_909 (O_909,N_29739,N_29557);
nor UO_910 (O_910,N_28687,N_28964);
xor UO_911 (O_911,N_29740,N_29197);
nor UO_912 (O_912,N_29416,N_29963);
or UO_913 (O_913,N_29284,N_29675);
nor UO_914 (O_914,N_29617,N_28984);
or UO_915 (O_915,N_28916,N_28660);
nor UO_916 (O_916,N_29586,N_29082);
and UO_917 (O_917,N_29746,N_28687);
or UO_918 (O_918,N_28792,N_28785);
nand UO_919 (O_919,N_28777,N_29544);
or UO_920 (O_920,N_29623,N_29874);
and UO_921 (O_921,N_28698,N_29003);
or UO_922 (O_922,N_28813,N_29488);
and UO_923 (O_923,N_28533,N_29515);
xnor UO_924 (O_924,N_29398,N_29055);
and UO_925 (O_925,N_28741,N_29897);
or UO_926 (O_926,N_29060,N_29466);
xnor UO_927 (O_927,N_29624,N_29254);
xor UO_928 (O_928,N_29160,N_29414);
xor UO_929 (O_929,N_29779,N_29357);
and UO_930 (O_930,N_29361,N_28572);
or UO_931 (O_931,N_29291,N_29168);
xnor UO_932 (O_932,N_29201,N_29464);
nand UO_933 (O_933,N_29429,N_29630);
nor UO_934 (O_934,N_29529,N_29370);
xnor UO_935 (O_935,N_29716,N_29647);
or UO_936 (O_936,N_29441,N_28565);
or UO_937 (O_937,N_28842,N_28867);
or UO_938 (O_938,N_28523,N_29062);
or UO_939 (O_939,N_28913,N_29207);
and UO_940 (O_940,N_28799,N_29615);
or UO_941 (O_941,N_29740,N_29257);
nor UO_942 (O_942,N_29380,N_29710);
nand UO_943 (O_943,N_29092,N_29338);
nand UO_944 (O_944,N_29739,N_29650);
nand UO_945 (O_945,N_28573,N_28805);
nor UO_946 (O_946,N_29728,N_29528);
nand UO_947 (O_947,N_29836,N_29947);
nor UO_948 (O_948,N_28655,N_29337);
nand UO_949 (O_949,N_29342,N_29001);
and UO_950 (O_950,N_29862,N_29186);
and UO_951 (O_951,N_28885,N_28983);
or UO_952 (O_952,N_29344,N_28932);
and UO_953 (O_953,N_29032,N_29583);
and UO_954 (O_954,N_29601,N_28663);
nor UO_955 (O_955,N_29968,N_29253);
nand UO_956 (O_956,N_29423,N_29017);
and UO_957 (O_957,N_29286,N_29217);
and UO_958 (O_958,N_29924,N_29390);
and UO_959 (O_959,N_29003,N_29811);
xnor UO_960 (O_960,N_29743,N_29146);
xor UO_961 (O_961,N_29443,N_29411);
xor UO_962 (O_962,N_29727,N_29664);
or UO_963 (O_963,N_28876,N_29654);
nor UO_964 (O_964,N_28931,N_29628);
xor UO_965 (O_965,N_28895,N_28879);
and UO_966 (O_966,N_29022,N_29056);
nor UO_967 (O_967,N_28909,N_29508);
or UO_968 (O_968,N_28966,N_28653);
xor UO_969 (O_969,N_28680,N_29574);
nor UO_970 (O_970,N_28838,N_28616);
nand UO_971 (O_971,N_29247,N_29771);
nor UO_972 (O_972,N_28859,N_28665);
nor UO_973 (O_973,N_29068,N_28629);
or UO_974 (O_974,N_29795,N_29728);
xor UO_975 (O_975,N_28520,N_29100);
xnor UO_976 (O_976,N_28869,N_28616);
or UO_977 (O_977,N_28935,N_28904);
xor UO_978 (O_978,N_29386,N_28990);
nor UO_979 (O_979,N_29764,N_29842);
xor UO_980 (O_980,N_29502,N_29688);
or UO_981 (O_981,N_29715,N_29520);
nor UO_982 (O_982,N_28706,N_29950);
nor UO_983 (O_983,N_29033,N_29582);
and UO_984 (O_984,N_29458,N_29159);
or UO_985 (O_985,N_29388,N_28531);
nand UO_986 (O_986,N_29669,N_29825);
nor UO_987 (O_987,N_29997,N_29338);
or UO_988 (O_988,N_29328,N_29383);
nand UO_989 (O_989,N_28983,N_29464);
and UO_990 (O_990,N_29479,N_29824);
and UO_991 (O_991,N_29853,N_28925);
nand UO_992 (O_992,N_29985,N_28838);
nor UO_993 (O_993,N_28537,N_29828);
or UO_994 (O_994,N_29366,N_29165);
nor UO_995 (O_995,N_28775,N_29521);
xnor UO_996 (O_996,N_29990,N_28586);
xor UO_997 (O_997,N_29498,N_29412);
nor UO_998 (O_998,N_29747,N_29713);
or UO_999 (O_999,N_29263,N_28851);
nand UO_1000 (O_1000,N_29327,N_29050);
nand UO_1001 (O_1001,N_29054,N_28925);
xor UO_1002 (O_1002,N_29078,N_28878);
or UO_1003 (O_1003,N_29518,N_28867);
or UO_1004 (O_1004,N_28682,N_28875);
nand UO_1005 (O_1005,N_28747,N_29413);
nand UO_1006 (O_1006,N_29457,N_28690);
nor UO_1007 (O_1007,N_29030,N_28537);
nor UO_1008 (O_1008,N_28748,N_29796);
xor UO_1009 (O_1009,N_29892,N_29572);
nand UO_1010 (O_1010,N_28660,N_29987);
and UO_1011 (O_1011,N_29673,N_29593);
or UO_1012 (O_1012,N_28793,N_29189);
nor UO_1013 (O_1013,N_28671,N_29742);
xnor UO_1014 (O_1014,N_29017,N_28619);
or UO_1015 (O_1015,N_29937,N_28597);
nand UO_1016 (O_1016,N_28521,N_29351);
or UO_1017 (O_1017,N_29727,N_28814);
and UO_1018 (O_1018,N_28986,N_29337);
and UO_1019 (O_1019,N_28900,N_29348);
and UO_1020 (O_1020,N_29851,N_29981);
and UO_1021 (O_1021,N_29518,N_29160);
xnor UO_1022 (O_1022,N_29043,N_29833);
nand UO_1023 (O_1023,N_28648,N_28831);
xor UO_1024 (O_1024,N_29260,N_28691);
nand UO_1025 (O_1025,N_29747,N_28894);
and UO_1026 (O_1026,N_28637,N_28890);
nor UO_1027 (O_1027,N_28598,N_29823);
and UO_1028 (O_1028,N_28591,N_29494);
xor UO_1029 (O_1029,N_29126,N_28690);
and UO_1030 (O_1030,N_28586,N_28877);
nand UO_1031 (O_1031,N_29775,N_28603);
xnor UO_1032 (O_1032,N_29620,N_28925);
and UO_1033 (O_1033,N_28611,N_28641);
and UO_1034 (O_1034,N_29327,N_29673);
and UO_1035 (O_1035,N_28926,N_28557);
xor UO_1036 (O_1036,N_29097,N_29939);
or UO_1037 (O_1037,N_28935,N_28691);
xor UO_1038 (O_1038,N_28838,N_29068);
and UO_1039 (O_1039,N_28703,N_29322);
and UO_1040 (O_1040,N_29752,N_29742);
and UO_1041 (O_1041,N_29129,N_28779);
xnor UO_1042 (O_1042,N_28866,N_28839);
nor UO_1043 (O_1043,N_29391,N_29171);
xor UO_1044 (O_1044,N_28926,N_29723);
nor UO_1045 (O_1045,N_28598,N_29391);
xnor UO_1046 (O_1046,N_28514,N_29926);
or UO_1047 (O_1047,N_29281,N_29130);
or UO_1048 (O_1048,N_29352,N_28854);
xor UO_1049 (O_1049,N_28827,N_28867);
and UO_1050 (O_1050,N_29567,N_29643);
and UO_1051 (O_1051,N_28507,N_29691);
nor UO_1052 (O_1052,N_29050,N_29256);
nand UO_1053 (O_1053,N_29185,N_29804);
xor UO_1054 (O_1054,N_29501,N_28527);
nand UO_1055 (O_1055,N_29342,N_29783);
and UO_1056 (O_1056,N_29934,N_29942);
nand UO_1057 (O_1057,N_28918,N_29798);
nand UO_1058 (O_1058,N_29254,N_29936);
nor UO_1059 (O_1059,N_29519,N_29429);
nand UO_1060 (O_1060,N_29679,N_29082);
nand UO_1061 (O_1061,N_28896,N_28684);
nand UO_1062 (O_1062,N_29193,N_29873);
nand UO_1063 (O_1063,N_29441,N_29457);
nand UO_1064 (O_1064,N_28688,N_28576);
and UO_1065 (O_1065,N_29768,N_29582);
xnor UO_1066 (O_1066,N_28500,N_29376);
nor UO_1067 (O_1067,N_29228,N_28855);
or UO_1068 (O_1068,N_28828,N_29014);
xnor UO_1069 (O_1069,N_29812,N_28645);
nor UO_1070 (O_1070,N_28598,N_29170);
or UO_1071 (O_1071,N_29930,N_29015);
nand UO_1072 (O_1072,N_28650,N_28967);
nor UO_1073 (O_1073,N_29477,N_28858);
xnor UO_1074 (O_1074,N_29603,N_29050);
or UO_1075 (O_1075,N_29730,N_29195);
xor UO_1076 (O_1076,N_28615,N_28860);
and UO_1077 (O_1077,N_28938,N_29079);
nand UO_1078 (O_1078,N_29471,N_29763);
nand UO_1079 (O_1079,N_28629,N_28546);
xor UO_1080 (O_1080,N_28922,N_29663);
nand UO_1081 (O_1081,N_28541,N_29630);
nand UO_1082 (O_1082,N_28532,N_29283);
nor UO_1083 (O_1083,N_29272,N_28901);
nor UO_1084 (O_1084,N_28842,N_29869);
or UO_1085 (O_1085,N_29900,N_29448);
xnor UO_1086 (O_1086,N_28975,N_28994);
nor UO_1087 (O_1087,N_28900,N_28955);
nor UO_1088 (O_1088,N_29023,N_29907);
nor UO_1089 (O_1089,N_29758,N_29980);
xor UO_1090 (O_1090,N_28587,N_28711);
and UO_1091 (O_1091,N_29330,N_28937);
nor UO_1092 (O_1092,N_29947,N_28754);
xor UO_1093 (O_1093,N_29720,N_29269);
nand UO_1094 (O_1094,N_29629,N_29631);
and UO_1095 (O_1095,N_29996,N_29348);
nand UO_1096 (O_1096,N_29614,N_29434);
nand UO_1097 (O_1097,N_29012,N_29597);
nand UO_1098 (O_1098,N_28740,N_29875);
nand UO_1099 (O_1099,N_29218,N_28734);
xor UO_1100 (O_1100,N_28833,N_29198);
or UO_1101 (O_1101,N_29789,N_29687);
or UO_1102 (O_1102,N_28914,N_29159);
or UO_1103 (O_1103,N_28960,N_28727);
nor UO_1104 (O_1104,N_29511,N_29991);
nand UO_1105 (O_1105,N_28716,N_29419);
nand UO_1106 (O_1106,N_28632,N_28675);
nor UO_1107 (O_1107,N_28822,N_28600);
nand UO_1108 (O_1108,N_29427,N_28525);
xnor UO_1109 (O_1109,N_28543,N_29566);
and UO_1110 (O_1110,N_29524,N_29689);
and UO_1111 (O_1111,N_28622,N_29878);
xor UO_1112 (O_1112,N_28928,N_28655);
xnor UO_1113 (O_1113,N_29640,N_29627);
nand UO_1114 (O_1114,N_28789,N_28905);
or UO_1115 (O_1115,N_29250,N_28580);
nand UO_1116 (O_1116,N_29409,N_29137);
or UO_1117 (O_1117,N_29832,N_29825);
or UO_1118 (O_1118,N_29319,N_29621);
nand UO_1119 (O_1119,N_29076,N_29880);
nand UO_1120 (O_1120,N_29872,N_29602);
nor UO_1121 (O_1121,N_29138,N_29218);
and UO_1122 (O_1122,N_29849,N_29134);
or UO_1123 (O_1123,N_29763,N_28626);
xor UO_1124 (O_1124,N_29070,N_29481);
or UO_1125 (O_1125,N_29277,N_29244);
nand UO_1126 (O_1126,N_29104,N_29723);
or UO_1127 (O_1127,N_29558,N_29694);
or UO_1128 (O_1128,N_28528,N_29018);
xor UO_1129 (O_1129,N_28504,N_29260);
nand UO_1130 (O_1130,N_28633,N_28914);
xor UO_1131 (O_1131,N_29752,N_28599);
xnor UO_1132 (O_1132,N_29112,N_29887);
or UO_1133 (O_1133,N_29290,N_28670);
and UO_1134 (O_1134,N_28532,N_29954);
or UO_1135 (O_1135,N_29359,N_28649);
nand UO_1136 (O_1136,N_28797,N_29777);
nor UO_1137 (O_1137,N_29241,N_29337);
xnor UO_1138 (O_1138,N_29229,N_29933);
or UO_1139 (O_1139,N_28799,N_29503);
nand UO_1140 (O_1140,N_29102,N_28823);
nand UO_1141 (O_1141,N_29504,N_28819);
xnor UO_1142 (O_1142,N_29785,N_29360);
nand UO_1143 (O_1143,N_29918,N_29415);
and UO_1144 (O_1144,N_29598,N_29925);
nor UO_1145 (O_1145,N_29278,N_28582);
or UO_1146 (O_1146,N_29875,N_29231);
and UO_1147 (O_1147,N_29725,N_28957);
nand UO_1148 (O_1148,N_28993,N_29678);
nor UO_1149 (O_1149,N_29836,N_29326);
xnor UO_1150 (O_1150,N_28675,N_28996);
or UO_1151 (O_1151,N_28876,N_28937);
xor UO_1152 (O_1152,N_28693,N_29438);
nand UO_1153 (O_1153,N_29844,N_28937);
nor UO_1154 (O_1154,N_29164,N_29926);
or UO_1155 (O_1155,N_29213,N_28642);
xnor UO_1156 (O_1156,N_28817,N_29015);
or UO_1157 (O_1157,N_28779,N_28726);
and UO_1158 (O_1158,N_28566,N_29284);
nor UO_1159 (O_1159,N_29001,N_28943);
xor UO_1160 (O_1160,N_28919,N_28658);
nand UO_1161 (O_1161,N_29672,N_29608);
nand UO_1162 (O_1162,N_29599,N_28746);
nor UO_1163 (O_1163,N_28955,N_29171);
or UO_1164 (O_1164,N_28505,N_29451);
xnor UO_1165 (O_1165,N_28653,N_28606);
nand UO_1166 (O_1166,N_28769,N_29564);
nor UO_1167 (O_1167,N_29568,N_29875);
nor UO_1168 (O_1168,N_29237,N_29959);
nand UO_1169 (O_1169,N_29837,N_29420);
nand UO_1170 (O_1170,N_29784,N_29812);
or UO_1171 (O_1171,N_29951,N_29914);
nor UO_1172 (O_1172,N_29982,N_29843);
xor UO_1173 (O_1173,N_29969,N_29200);
nand UO_1174 (O_1174,N_29558,N_29185);
and UO_1175 (O_1175,N_28841,N_29465);
nor UO_1176 (O_1176,N_29581,N_29923);
nor UO_1177 (O_1177,N_29617,N_29626);
or UO_1178 (O_1178,N_29452,N_28855);
xnor UO_1179 (O_1179,N_28815,N_28559);
xor UO_1180 (O_1180,N_29248,N_29578);
nor UO_1181 (O_1181,N_29483,N_29256);
or UO_1182 (O_1182,N_29928,N_29802);
and UO_1183 (O_1183,N_28771,N_28685);
and UO_1184 (O_1184,N_29779,N_29037);
xnor UO_1185 (O_1185,N_29469,N_29211);
xor UO_1186 (O_1186,N_28957,N_29630);
nor UO_1187 (O_1187,N_29854,N_29204);
xnor UO_1188 (O_1188,N_28607,N_29562);
and UO_1189 (O_1189,N_28760,N_29418);
or UO_1190 (O_1190,N_29319,N_29804);
xnor UO_1191 (O_1191,N_28921,N_28754);
nor UO_1192 (O_1192,N_28920,N_28905);
nor UO_1193 (O_1193,N_28823,N_29860);
nor UO_1194 (O_1194,N_28930,N_29687);
nand UO_1195 (O_1195,N_29419,N_28522);
and UO_1196 (O_1196,N_29053,N_28611);
nor UO_1197 (O_1197,N_29412,N_29949);
or UO_1198 (O_1198,N_29016,N_28701);
xnor UO_1199 (O_1199,N_28784,N_29516);
xor UO_1200 (O_1200,N_29000,N_28985);
nor UO_1201 (O_1201,N_29139,N_29462);
nand UO_1202 (O_1202,N_28811,N_28604);
xor UO_1203 (O_1203,N_28515,N_29241);
and UO_1204 (O_1204,N_29518,N_29558);
nand UO_1205 (O_1205,N_28757,N_29895);
nor UO_1206 (O_1206,N_29420,N_29818);
or UO_1207 (O_1207,N_29750,N_29511);
and UO_1208 (O_1208,N_28761,N_28635);
nor UO_1209 (O_1209,N_29359,N_29335);
xnor UO_1210 (O_1210,N_28708,N_29110);
xor UO_1211 (O_1211,N_29022,N_28812);
xor UO_1212 (O_1212,N_28631,N_28885);
or UO_1213 (O_1213,N_28909,N_29448);
xor UO_1214 (O_1214,N_29589,N_29980);
and UO_1215 (O_1215,N_29745,N_29893);
nor UO_1216 (O_1216,N_29222,N_28709);
or UO_1217 (O_1217,N_29377,N_29410);
nand UO_1218 (O_1218,N_29229,N_29560);
or UO_1219 (O_1219,N_29489,N_29547);
nor UO_1220 (O_1220,N_28544,N_29888);
or UO_1221 (O_1221,N_29877,N_29461);
or UO_1222 (O_1222,N_28609,N_29132);
nand UO_1223 (O_1223,N_29387,N_29262);
nand UO_1224 (O_1224,N_29265,N_29630);
nor UO_1225 (O_1225,N_29802,N_28948);
nor UO_1226 (O_1226,N_29140,N_29156);
xnor UO_1227 (O_1227,N_29743,N_29048);
nand UO_1228 (O_1228,N_29006,N_28618);
nand UO_1229 (O_1229,N_29875,N_29474);
nor UO_1230 (O_1230,N_29165,N_29037);
xnor UO_1231 (O_1231,N_29196,N_28541);
nor UO_1232 (O_1232,N_28795,N_29636);
or UO_1233 (O_1233,N_29149,N_29861);
or UO_1234 (O_1234,N_29894,N_29389);
or UO_1235 (O_1235,N_28728,N_29678);
xnor UO_1236 (O_1236,N_29727,N_29540);
nor UO_1237 (O_1237,N_28816,N_29348);
and UO_1238 (O_1238,N_28638,N_29544);
or UO_1239 (O_1239,N_29504,N_29385);
or UO_1240 (O_1240,N_29895,N_29364);
xnor UO_1241 (O_1241,N_29945,N_29749);
xor UO_1242 (O_1242,N_28931,N_29228);
xnor UO_1243 (O_1243,N_29245,N_29675);
and UO_1244 (O_1244,N_29437,N_29956);
nor UO_1245 (O_1245,N_29499,N_29859);
xnor UO_1246 (O_1246,N_29974,N_29946);
xnor UO_1247 (O_1247,N_29464,N_29070);
and UO_1248 (O_1248,N_29891,N_29178);
nor UO_1249 (O_1249,N_29021,N_28849);
xor UO_1250 (O_1250,N_28868,N_29891);
xnor UO_1251 (O_1251,N_28906,N_29417);
and UO_1252 (O_1252,N_29193,N_28615);
nand UO_1253 (O_1253,N_29466,N_29631);
nand UO_1254 (O_1254,N_29288,N_28509);
nor UO_1255 (O_1255,N_28596,N_29600);
xnor UO_1256 (O_1256,N_29162,N_29801);
nand UO_1257 (O_1257,N_28560,N_29795);
xor UO_1258 (O_1258,N_29894,N_29635);
xnor UO_1259 (O_1259,N_29589,N_29039);
nand UO_1260 (O_1260,N_28844,N_29130);
and UO_1261 (O_1261,N_29202,N_29439);
xnor UO_1262 (O_1262,N_29863,N_29014);
nand UO_1263 (O_1263,N_29758,N_28574);
nand UO_1264 (O_1264,N_29173,N_29887);
nand UO_1265 (O_1265,N_29277,N_29726);
nand UO_1266 (O_1266,N_28819,N_29248);
and UO_1267 (O_1267,N_29969,N_28678);
or UO_1268 (O_1268,N_29486,N_29235);
nand UO_1269 (O_1269,N_29865,N_29975);
nor UO_1270 (O_1270,N_28883,N_29729);
nor UO_1271 (O_1271,N_29999,N_29606);
or UO_1272 (O_1272,N_29524,N_29312);
nand UO_1273 (O_1273,N_29613,N_29594);
and UO_1274 (O_1274,N_28638,N_28933);
and UO_1275 (O_1275,N_29928,N_29962);
or UO_1276 (O_1276,N_29390,N_28535);
xor UO_1277 (O_1277,N_29474,N_28875);
nand UO_1278 (O_1278,N_29769,N_28575);
xnor UO_1279 (O_1279,N_29624,N_29426);
nor UO_1280 (O_1280,N_28537,N_28805);
xor UO_1281 (O_1281,N_29693,N_29005);
xor UO_1282 (O_1282,N_29636,N_29616);
xnor UO_1283 (O_1283,N_29926,N_29368);
and UO_1284 (O_1284,N_28739,N_29357);
and UO_1285 (O_1285,N_29175,N_29712);
or UO_1286 (O_1286,N_29272,N_28858);
and UO_1287 (O_1287,N_28946,N_28620);
nand UO_1288 (O_1288,N_29223,N_28655);
xnor UO_1289 (O_1289,N_29392,N_29757);
or UO_1290 (O_1290,N_28866,N_29192);
nor UO_1291 (O_1291,N_28808,N_29396);
xnor UO_1292 (O_1292,N_28509,N_29904);
xor UO_1293 (O_1293,N_28531,N_28931);
nor UO_1294 (O_1294,N_29969,N_29085);
and UO_1295 (O_1295,N_28909,N_29641);
nand UO_1296 (O_1296,N_28865,N_29238);
nand UO_1297 (O_1297,N_29345,N_28833);
nor UO_1298 (O_1298,N_29230,N_28645);
or UO_1299 (O_1299,N_28982,N_29107);
xnor UO_1300 (O_1300,N_29356,N_29725);
xor UO_1301 (O_1301,N_28629,N_28599);
and UO_1302 (O_1302,N_28511,N_29008);
and UO_1303 (O_1303,N_29648,N_29902);
nand UO_1304 (O_1304,N_29367,N_29865);
nand UO_1305 (O_1305,N_29635,N_28615);
and UO_1306 (O_1306,N_29693,N_29730);
and UO_1307 (O_1307,N_29122,N_29011);
or UO_1308 (O_1308,N_29163,N_29886);
nor UO_1309 (O_1309,N_29775,N_28999);
nand UO_1310 (O_1310,N_28714,N_29820);
and UO_1311 (O_1311,N_28768,N_29179);
xor UO_1312 (O_1312,N_29765,N_29903);
nor UO_1313 (O_1313,N_29174,N_29526);
nand UO_1314 (O_1314,N_29316,N_28916);
and UO_1315 (O_1315,N_29872,N_29019);
and UO_1316 (O_1316,N_29977,N_28784);
nand UO_1317 (O_1317,N_29023,N_28759);
nor UO_1318 (O_1318,N_28894,N_29889);
nand UO_1319 (O_1319,N_28978,N_28913);
xor UO_1320 (O_1320,N_28980,N_28593);
nand UO_1321 (O_1321,N_29661,N_29608);
or UO_1322 (O_1322,N_29522,N_29662);
or UO_1323 (O_1323,N_29041,N_28778);
and UO_1324 (O_1324,N_29313,N_28811);
nand UO_1325 (O_1325,N_29038,N_29798);
and UO_1326 (O_1326,N_29589,N_29186);
nor UO_1327 (O_1327,N_29019,N_29415);
xor UO_1328 (O_1328,N_29364,N_29088);
xor UO_1329 (O_1329,N_29879,N_29604);
xor UO_1330 (O_1330,N_29187,N_29869);
and UO_1331 (O_1331,N_29674,N_29426);
or UO_1332 (O_1332,N_29120,N_29188);
or UO_1333 (O_1333,N_29368,N_29606);
nor UO_1334 (O_1334,N_29571,N_29947);
or UO_1335 (O_1335,N_29065,N_28850);
nor UO_1336 (O_1336,N_29489,N_28880);
or UO_1337 (O_1337,N_29770,N_29779);
xnor UO_1338 (O_1338,N_29850,N_29997);
or UO_1339 (O_1339,N_28838,N_29069);
and UO_1340 (O_1340,N_29345,N_29296);
or UO_1341 (O_1341,N_29925,N_29451);
xnor UO_1342 (O_1342,N_29757,N_29981);
nand UO_1343 (O_1343,N_29578,N_28965);
nand UO_1344 (O_1344,N_29681,N_28814);
nor UO_1345 (O_1345,N_28781,N_29401);
or UO_1346 (O_1346,N_29015,N_29926);
and UO_1347 (O_1347,N_28601,N_29224);
xnor UO_1348 (O_1348,N_28765,N_29991);
or UO_1349 (O_1349,N_29871,N_29137);
xor UO_1350 (O_1350,N_28743,N_29810);
nand UO_1351 (O_1351,N_29149,N_29410);
and UO_1352 (O_1352,N_28934,N_29366);
nor UO_1353 (O_1353,N_29460,N_28799);
or UO_1354 (O_1354,N_28821,N_28874);
and UO_1355 (O_1355,N_29496,N_29007);
and UO_1356 (O_1356,N_29213,N_29449);
nand UO_1357 (O_1357,N_28584,N_28635);
and UO_1358 (O_1358,N_28965,N_28688);
nor UO_1359 (O_1359,N_28675,N_28956);
and UO_1360 (O_1360,N_29544,N_29829);
nand UO_1361 (O_1361,N_29651,N_29024);
or UO_1362 (O_1362,N_29070,N_29157);
nor UO_1363 (O_1363,N_29825,N_28568);
or UO_1364 (O_1364,N_29856,N_28862);
nor UO_1365 (O_1365,N_29259,N_28542);
xnor UO_1366 (O_1366,N_29500,N_28747);
and UO_1367 (O_1367,N_28586,N_29821);
xor UO_1368 (O_1368,N_29987,N_29065);
nor UO_1369 (O_1369,N_28856,N_28693);
nand UO_1370 (O_1370,N_29639,N_28771);
nand UO_1371 (O_1371,N_29902,N_28641);
xor UO_1372 (O_1372,N_29056,N_29883);
xnor UO_1373 (O_1373,N_29153,N_29525);
and UO_1374 (O_1374,N_29112,N_29414);
or UO_1375 (O_1375,N_28794,N_29137);
xnor UO_1376 (O_1376,N_29698,N_28888);
xor UO_1377 (O_1377,N_29426,N_29793);
or UO_1378 (O_1378,N_29973,N_29159);
and UO_1379 (O_1379,N_28828,N_29156);
and UO_1380 (O_1380,N_29811,N_28804);
and UO_1381 (O_1381,N_29663,N_29793);
nor UO_1382 (O_1382,N_28785,N_28658);
and UO_1383 (O_1383,N_29234,N_29003);
or UO_1384 (O_1384,N_29993,N_29920);
or UO_1385 (O_1385,N_28616,N_28792);
or UO_1386 (O_1386,N_29639,N_28784);
nand UO_1387 (O_1387,N_29201,N_29810);
xnor UO_1388 (O_1388,N_29394,N_29459);
and UO_1389 (O_1389,N_29080,N_29747);
nand UO_1390 (O_1390,N_29094,N_29727);
and UO_1391 (O_1391,N_29088,N_28852);
nand UO_1392 (O_1392,N_29830,N_29453);
nor UO_1393 (O_1393,N_29505,N_28726);
nor UO_1394 (O_1394,N_29624,N_29858);
or UO_1395 (O_1395,N_29962,N_29332);
nor UO_1396 (O_1396,N_29923,N_29123);
and UO_1397 (O_1397,N_28974,N_28987);
and UO_1398 (O_1398,N_28902,N_29303);
nor UO_1399 (O_1399,N_29111,N_29470);
nor UO_1400 (O_1400,N_28979,N_28636);
nand UO_1401 (O_1401,N_29893,N_28996);
and UO_1402 (O_1402,N_28508,N_28752);
nand UO_1403 (O_1403,N_29173,N_29454);
or UO_1404 (O_1404,N_29274,N_29643);
nor UO_1405 (O_1405,N_29346,N_29066);
nand UO_1406 (O_1406,N_29351,N_29763);
or UO_1407 (O_1407,N_28635,N_28594);
or UO_1408 (O_1408,N_29879,N_28843);
nor UO_1409 (O_1409,N_29072,N_29750);
nor UO_1410 (O_1410,N_28807,N_29358);
nor UO_1411 (O_1411,N_29902,N_28849);
or UO_1412 (O_1412,N_29390,N_28681);
and UO_1413 (O_1413,N_29867,N_29145);
or UO_1414 (O_1414,N_28713,N_28666);
nor UO_1415 (O_1415,N_28510,N_29924);
and UO_1416 (O_1416,N_28794,N_28624);
nand UO_1417 (O_1417,N_29016,N_29238);
and UO_1418 (O_1418,N_29622,N_29405);
and UO_1419 (O_1419,N_28868,N_29878);
or UO_1420 (O_1420,N_28784,N_29912);
or UO_1421 (O_1421,N_29867,N_29590);
xor UO_1422 (O_1422,N_28966,N_29559);
and UO_1423 (O_1423,N_29130,N_29238);
or UO_1424 (O_1424,N_29436,N_28554);
and UO_1425 (O_1425,N_29494,N_29194);
nor UO_1426 (O_1426,N_29492,N_28837);
nand UO_1427 (O_1427,N_29237,N_29615);
or UO_1428 (O_1428,N_29725,N_29712);
nor UO_1429 (O_1429,N_29647,N_29336);
nor UO_1430 (O_1430,N_29611,N_29885);
nand UO_1431 (O_1431,N_29388,N_29265);
xor UO_1432 (O_1432,N_28912,N_29560);
xor UO_1433 (O_1433,N_28542,N_29572);
nand UO_1434 (O_1434,N_29033,N_29264);
nand UO_1435 (O_1435,N_28785,N_28850);
nand UO_1436 (O_1436,N_28519,N_28624);
nand UO_1437 (O_1437,N_29052,N_29821);
or UO_1438 (O_1438,N_29213,N_29050);
nor UO_1439 (O_1439,N_29773,N_29411);
or UO_1440 (O_1440,N_29439,N_28952);
xnor UO_1441 (O_1441,N_29519,N_29197);
nor UO_1442 (O_1442,N_28890,N_28669);
nand UO_1443 (O_1443,N_29432,N_29325);
or UO_1444 (O_1444,N_29877,N_28971);
xor UO_1445 (O_1445,N_28502,N_29524);
nor UO_1446 (O_1446,N_29084,N_28510);
and UO_1447 (O_1447,N_29193,N_29628);
and UO_1448 (O_1448,N_29625,N_28782);
or UO_1449 (O_1449,N_29001,N_28687);
and UO_1450 (O_1450,N_29881,N_29026);
xnor UO_1451 (O_1451,N_28862,N_28527);
or UO_1452 (O_1452,N_29999,N_29859);
xor UO_1453 (O_1453,N_28971,N_28748);
and UO_1454 (O_1454,N_28723,N_29678);
or UO_1455 (O_1455,N_28967,N_29110);
xor UO_1456 (O_1456,N_29154,N_28925);
or UO_1457 (O_1457,N_28889,N_29943);
or UO_1458 (O_1458,N_28678,N_29414);
xnor UO_1459 (O_1459,N_29288,N_29218);
nand UO_1460 (O_1460,N_28894,N_29371);
nor UO_1461 (O_1461,N_29132,N_29024);
xor UO_1462 (O_1462,N_29671,N_28757);
and UO_1463 (O_1463,N_28537,N_28713);
and UO_1464 (O_1464,N_29835,N_29143);
and UO_1465 (O_1465,N_28941,N_29606);
nor UO_1466 (O_1466,N_28992,N_29478);
or UO_1467 (O_1467,N_29434,N_28795);
nor UO_1468 (O_1468,N_29683,N_29847);
nor UO_1469 (O_1469,N_29332,N_29877);
xor UO_1470 (O_1470,N_28539,N_28985);
nor UO_1471 (O_1471,N_28954,N_29232);
xor UO_1472 (O_1472,N_29738,N_28626);
nor UO_1473 (O_1473,N_29831,N_29938);
or UO_1474 (O_1474,N_28743,N_29904);
nor UO_1475 (O_1475,N_29821,N_29400);
nand UO_1476 (O_1476,N_28644,N_28993);
nor UO_1477 (O_1477,N_29680,N_29781);
or UO_1478 (O_1478,N_29445,N_29803);
xnor UO_1479 (O_1479,N_29299,N_28817);
or UO_1480 (O_1480,N_28769,N_28666);
or UO_1481 (O_1481,N_29435,N_29166);
nor UO_1482 (O_1482,N_29679,N_29023);
nor UO_1483 (O_1483,N_29257,N_28654);
xnor UO_1484 (O_1484,N_28519,N_29366);
nor UO_1485 (O_1485,N_29777,N_29909);
nor UO_1486 (O_1486,N_28693,N_29529);
or UO_1487 (O_1487,N_29596,N_29701);
xor UO_1488 (O_1488,N_29259,N_29484);
and UO_1489 (O_1489,N_29229,N_29161);
and UO_1490 (O_1490,N_29742,N_28943);
and UO_1491 (O_1491,N_29432,N_29289);
and UO_1492 (O_1492,N_28910,N_29054);
nor UO_1493 (O_1493,N_28963,N_28862);
nand UO_1494 (O_1494,N_29938,N_29560);
nor UO_1495 (O_1495,N_29856,N_29243);
or UO_1496 (O_1496,N_29570,N_29701);
nand UO_1497 (O_1497,N_29543,N_29653);
or UO_1498 (O_1498,N_29217,N_29274);
and UO_1499 (O_1499,N_28512,N_28757);
xor UO_1500 (O_1500,N_28727,N_29874);
nand UO_1501 (O_1501,N_28813,N_29243);
nor UO_1502 (O_1502,N_28540,N_28690);
xor UO_1503 (O_1503,N_29762,N_29764);
nor UO_1504 (O_1504,N_29045,N_29169);
xor UO_1505 (O_1505,N_29373,N_29336);
or UO_1506 (O_1506,N_29739,N_28688);
xor UO_1507 (O_1507,N_28734,N_28601);
and UO_1508 (O_1508,N_29347,N_28696);
and UO_1509 (O_1509,N_29094,N_29216);
and UO_1510 (O_1510,N_28546,N_29152);
nor UO_1511 (O_1511,N_29770,N_29524);
xnor UO_1512 (O_1512,N_28995,N_29512);
or UO_1513 (O_1513,N_28963,N_29831);
or UO_1514 (O_1514,N_29687,N_29323);
and UO_1515 (O_1515,N_29046,N_29075);
xor UO_1516 (O_1516,N_28899,N_28648);
xor UO_1517 (O_1517,N_29027,N_29905);
or UO_1518 (O_1518,N_28747,N_29869);
or UO_1519 (O_1519,N_29646,N_28746);
nor UO_1520 (O_1520,N_29414,N_29335);
nor UO_1521 (O_1521,N_29729,N_29464);
nor UO_1522 (O_1522,N_28877,N_28643);
nor UO_1523 (O_1523,N_29608,N_28819);
nand UO_1524 (O_1524,N_28989,N_28602);
and UO_1525 (O_1525,N_29759,N_29511);
xnor UO_1526 (O_1526,N_28621,N_29772);
xor UO_1527 (O_1527,N_29306,N_29343);
or UO_1528 (O_1528,N_29188,N_29786);
or UO_1529 (O_1529,N_28717,N_29834);
and UO_1530 (O_1530,N_29484,N_29867);
nor UO_1531 (O_1531,N_28764,N_28630);
or UO_1532 (O_1532,N_29754,N_28864);
xnor UO_1533 (O_1533,N_28956,N_29213);
xnor UO_1534 (O_1534,N_29312,N_29711);
and UO_1535 (O_1535,N_29390,N_29027);
nand UO_1536 (O_1536,N_29509,N_28867);
xor UO_1537 (O_1537,N_29346,N_28881);
and UO_1538 (O_1538,N_29779,N_28616);
and UO_1539 (O_1539,N_29260,N_29189);
nand UO_1540 (O_1540,N_28666,N_29120);
and UO_1541 (O_1541,N_29034,N_29508);
and UO_1542 (O_1542,N_29870,N_29416);
xor UO_1543 (O_1543,N_29970,N_29450);
or UO_1544 (O_1544,N_29890,N_29057);
nor UO_1545 (O_1545,N_28549,N_28948);
xnor UO_1546 (O_1546,N_29431,N_28743);
nand UO_1547 (O_1547,N_29606,N_29809);
xnor UO_1548 (O_1548,N_29189,N_28672);
and UO_1549 (O_1549,N_29837,N_29716);
and UO_1550 (O_1550,N_28815,N_29148);
and UO_1551 (O_1551,N_28554,N_29593);
xor UO_1552 (O_1552,N_29463,N_29879);
and UO_1553 (O_1553,N_29477,N_29350);
xnor UO_1554 (O_1554,N_28925,N_28731);
or UO_1555 (O_1555,N_29668,N_29568);
nor UO_1556 (O_1556,N_29599,N_29108);
xor UO_1557 (O_1557,N_28571,N_29535);
xor UO_1558 (O_1558,N_29229,N_29676);
and UO_1559 (O_1559,N_29268,N_29376);
nand UO_1560 (O_1560,N_28702,N_29096);
and UO_1561 (O_1561,N_29925,N_29288);
or UO_1562 (O_1562,N_29470,N_29679);
xnor UO_1563 (O_1563,N_29839,N_28877);
or UO_1564 (O_1564,N_28647,N_29428);
xor UO_1565 (O_1565,N_29155,N_28852);
and UO_1566 (O_1566,N_29495,N_29446);
nor UO_1567 (O_1567,N_29121,N_29778);
and UO_1568 (O_1568,N_28700,N_29217);
or UO_1569 (O_1569,N_28770,N_28533);
and UO_1570 (O_1570,N_29931,N_29799);
nor UO_1571 (O_1571,N_29135,N_29398);
xor UO_1572 (O_1572,N_29127,N_28663);
and UO_1573 (O_1573,N_29200,N_29478);
xnor UO_1574 (O_1574,N_29316,N_29138);
and UO_1575 (O_1575,N_29893,N_29913);
nor UO_1576 (O_1576,N_29531,N_28994);
xor UO_1577 (O_1577,N_29347,N_28658);
nor UO_1578 (O_1578,N_29416,N_29812);
or UO_1579 (O_1579,N_29641,N_28739);
nor UO_1580 (O_1580,N_29081,N_29242);
nor UO_1581 (O_1581,N_29130,N_29910);
nand UO_1582 (O_1582,N_28993,N_28640);
and UO_1583 (O_1583,N_29597,N_29302);
and UO_1584 (O_1584,N_29751,N_29596);
xor UO_1585 (O_1585,N_29330,N_29432);
nand UO_1586 (O_1586,N_29383,N_29030);
nor UO_1587 (O_1587,N_28564,N_29883);
and UO_1588 (O_1588,N_28674,N_28619);
xnor UO_1589 (O_1589,N_29064,N_28712);
or UO_1590 (O_1590,N_28559,N_29654);
xnor UO_1591 (O_1591,N_29918,N_28627);
or UO_1592 (O_1592,N_29702,N_28701);
and UO_1593 (O_1593,N_29244,N_29415);
nand UO_1594 (O_1594,N_28771,N_29968);
or UO_1595 (O_1595,N_29946,N_29058);
xor UO_1596 (O_1596,N_29902,N_28828);
nand UO_1597 (O_1597,N_29059,N_28797);
and UO_1598 (O_1598,N_29123,N_29031);
xnor UO_1599 (O_1599,N_28649,N_29807);
nor UO_1600 (O_1600,N_28688,N_29430);
nand UO_1601 (O_1601,N_29823,N_28806);
nor UO_1602 (O_1602,N_29433,N_29901);
nor UO_1603 (O_1603,N_29189,N_28819);
xor UO_1604 (O_1604,N_29640,N_29593);
and UO_1605 (O_1605,N_29795,N_29166);
xor UO_1606 (O_1606,N_28739,N_28609);
nor UO_1607 (O_1607,N_28973,N_29263);
and UO_1608 (O_1608,N_29113,N_28554);
nand UO_1609 (O_1609,N_28606,N_29558);
nor UO_1610 (O_1610,N_28788,N_29863);
nor UO_1611 (O_1611,N_29568,N_29258);
xor UO_1612 (O_1612,N_29714,N_29182);
or UO_1613 (O_1613,N_29903,N_29367);
xnor UO_1614 (O_1614,N_28955,N_29929);
nor UO_1615 (O_1615,N_29235,N_29713);
nand UO_1616 (O_1616,N_29201,N_29430);
nand UO_1617 (O_1617,N_29638,N_28927);
and UO_1618 (O_1618,N_29118,N_29958);
or UO_1619 (O_1619,N_29278,N_29877);
nand UO_1620 (O_1620,N_29461,N_29288);
xor UO_1621 (O_1621,N_28769,N_28584);
or UO_1622 (O_1622,N_28988,N_28923);
nand UO_1623 (O_1623,N_29768,N_29935);
and UO_1624 (O_1624,N_29865,N_28634);
or UO_1625 (O_1625,N_29169,N_28665);
nand UO_1626 (O_1626,N_29151,N_29925);
and UO_1627 (O_1627,N_29692,N_29740);
nor UO_1628 (O_1628,N_29651,N_29759);
nand UO_1629 (O_1629,N_28652,N_29309);
xnor UO_1630 (O_1630,N_28984,N_29862);
nor UO_1631 (O_1631,N_29895,N_29270);
xnor UO_1632 (O_1632,N_28664,N_28529);
or UO_1633 (O_1633,N_29660,N_28642);
and UO_1634 (O_1634,N_28881,N_29111);
and UO_1635 (O_1635,N_29774,N_28963);
or UO_1636 (O_1636,N_29810,N_28987);
and UO_1637 (O_1637,N_28974,N_29875);
nand UO_1638 (O_1638,N_29262,N_29414);
nor UO_1639 (O_1639,N_28879,N_29506);
nor UO_1640 (O_1640,N_29532,N_28624);
and UO_1641 (O_1641,N_29518,N_29844);
nor UO_1642 (O_1642,N_29191,N_28749);
nand UO_1643 (O_1643,N_29842,N_29883);
xnor UO_1644 (O_1644,N_29022,N_28631);
nand UO_1645 (O_1645,N_29675,N_29663);
nand UO_1646 (O_1646,N_29410,N_28652);
and UO_1647 (O_1647,N_29894,N_28810);
or UO_1648 (O_1648,N_29893,N_29204);
or UO_1649 (O_1649,N_28680,N_29854);
nor UO_1650 (O_1650,N_28664,N_29175);
xnor UO_1651 (O_1651,N_28863,N_28667);
xor UO_1652 (O_1652,N_29544,N_28817);
xnor UO_1653 (O_1653,N_29360,N_29569);
xnor UO_1654 (O_1654,N_28545,N_28639);
nand UO_1655 (O_1655,N_28752,N_28516);
nand UO_1656 (O_1656,N_29521,N_29957);
nand UO_1657 (O_1657,N_29495,N_29230);
xnor UO_1658 (O_1658,N_29453,N_29414);
and UO_1659 (O_1659,N_29870,N_28733);
nand UO_1660 (O_1660,N_29964,N_28702);
and UO_1661 (O_1661,N_29884,N_28539);
nand UO_1662 (O_1662,N_28656,N_28867);
or UO_1663 (O_1663,N_29715,N_28973);
nand UO_1664 (O_1664,N_28755,N_29036);
and UO_1665 (O_1665,N_29655,N_28896);
nand UO_1666 (O_1666,N_29493,N_29187);
nand UO_1667 (O_1667,N_29638,N_28753);
nand UO_1668 (O_1668,N_29397,N_29601);
nand UO_1669 (O_1669,N_29669,N_29896);
and UO_1670 (O_1670,N_29277,N_29843);
and UO_1671 (O_1671,N_28742,N_29783);
and UO_1672 (O_1672,N_29745,N_28553);
or UO_1673 (O_1673,N_29780,N_29648);
nor UO_1674 (O_1674,N_29947,N_29289);
or UO_1675 (O_1675,N_29773,N_29884);
nor UO_1676 (O_1676,N_29034,N_29144);
nand UO_1677 (O_1677,N_28752,N_28989);
xor UO_1678 (O_1678,N_29020,N_28622);
nor UO_1679 (O_1679,N_29173,N_28764);
xnor UO_1680 (O_1680,N_29062,N_29037);
or UO_1681 (O_1681,N_29937,N_29662);
and UO_1682 (O_1682,N_29154,N_29547);
nand UO_1683 (O_1683,N_29451,N_29906);
xor UO_1684 (O_1684,N_28503,N_28967);
xor UO_1685 (O_1685,N_28675,N_29535);
nor UO_1686 (O_1686,N_28647,N_29535);
or UO_1687 (O_1687,N_29226,N_29244);
nand UO_1688 (O_1688,N_29761,N_29477);
nor UO_1689 (O_1689,N_29788,N_28829);
or UO_1690 (O_1690,N_29492,N_29529);
nor UO_1691 (O_1691,N_28619,N_29183);
and UO_1692 (O_1692,N_29725,N_29585);
nand UO_1693 (O_1693,N_29927,N_29820);
or UO_1694 (O_1694,N_29282,N_29917);
nand UO_1695 (O_1695,N_29945,N_28702);
and UO_1696 (O_1696,N_29319,N_29134);
and UO_1697 (O_1697,N_29913,N_28868);
nor UO_1698 (O_1698,N_28645,N_29238);
or UO_1699 (O_1699,N_29680,N_29705);
xor UO_1700 (O_1700,N_28787,N_28879);
xor UO_1701 (O_1701,N_29728,N_28999);
and UO_1702 (O_1702,N_29047,N_29925);
xnor UO_1703 (O_1703,N_29088,N_29078);
and UO_1704 (O_1704,N_28787,N_28594);
nand UO_1705 (O_1705,N_28534,N_29036);
xnor UO_1706 (O_1706,N_29710,N_29913);
and UO_1707 (O_1707,N_28631,N_28896);
and UO_1708 (O_1708,N_29553,N_28894);
nor UO_1709 (O_1709,N_29077,N_29484);
nand UO_1710 (O_1710,N_29256,N_29153);
nor UO_1711 (O_1711,N_29974,N_29125);
and UO_1712 (O_1712,N_29131,N_28670);
xor UO_1713 (O_1713,N_29297,N_29491);
and UO_1714 (O_1714,N_29422,N_29882);
nor UO_1715 (O_1715,N_29540,N_29861);
and UO_1716 (O_1716,N_28621,N_28971);
nor UO_1717 (O_1717,N_28869,N_29313);
and UO_1718 (O_1718,N_28763,N_29162);
nand UO_1719 (O_1719,N_28845,N_28756);
nand UO_1720 (O_1720,N_29150,N_29906);
or UO_1721 (O_1721,N_29770,N_28658);
nand UO_1722 (O_1722,N_29971,N_28820);
and UO_1723 (O_1723,N_29009,N_28924);
or UO_1724 (O_1724,N_29073,N_29124);
nand UO_1725 (O_1725,N_29760,N_28744);
nor UO_1726 (O_1726,N_29754,N_29282);
or UO_1727 (O_1727,N_29599,N_29123);
nand UO_1728 (O_1728,N_29110,N_29746);
xor UO_1729 (O_1729,N_28621,N_29530);
nor UO_1730 (O_1730,N_29089,N_28516);
or UO_1731 (O_1731,N_28839,N_29200);
and UO_1732 (O_1732,N_28942,N_29549);
or UO_1733 (O_1733,N_29190,N_28786);
xnor UO_1734 (O_1734,N_28608,N_29398);
or UO_1735 (O_1735,N_29042,N_29906);
and UO_1736 (O_1736,N_29091,N_28838);
and UO_1737 (O_1737,N_28733,N_29680);
nor UO_1738 (O_1738,N_29357,N_28850);
nand UO_1739 (O_1739,N_28756,N_28830);
xnor UO_1740 (O_1740,N_29160,N_28559);
nor UO_1741 (O_1741,N_28560,N_29865);
nor UO_1742 (O_1742,N_29101,N_29587);
nor UO_1743 (O_1743,N_29045,N_29753);
xor UO_1744 (O_1744,N_29066,N_29336);
xnor UO_1745 (O_1745,N_29566,N_29726);
or UO_1746 (O_1746,N_29493,N_29462);
nand UO_1747 (O_1747,N_29662,N_28939);
nor UO_1748 (O_1748,N_29957,N_28845);
and UO_1749 (O_1749,N_29219,N_28975);
or UO_1750 (O_1750,N_29081,N_29538);
nor UO_1751 (O_1751,N_29783,N_29612);
and UO_1752 (O_1752,N_29697,N_29324);
and UO_1753 (O_1753,N_29188,N_29743);
or UO_1754 (O_1754,N_29878,N_28765);
and UO_1755 (O_1755,N_29436,N_29844);
xnor UO_1756 (O_1756,N_29146,N_29222);
or UO_1757 (O_1757,N_28826,N_29146);
and UO_1758 (O_1758,N_29614,N_28640);
and UO_1759 (O_1759,N_29107,N_29264);
and UO_1760 (O_1760,N_29264,N_28752);
nor UO_1761 (O_1761,N_28502,N_29971);
or UO_1762 (O_1762,N_29422,N_28984);
xnor UO_1763 (O_1763,N_28652,N_29153);
and UO_1764 (O_1764,N_28699,N_28948);
and UO_1765 (O_1765,N_28821,N_29735);
or UO_1766 (O_1766,N_29445,N_28733);
nor UO_1767 (O_1767,N_28799,N_29668);
nor UO_1768 (O_1768,N_28739,N_29478);
and UO_1769 (O_1769,N_28802,N_28588);
nand UO_1770 (O_1770,N_29566,N_29623);
and UO_1771 (O_1771,N_29443,N_29701);
and UO_1772 (O_1772,N_29611,N_29483);
nand UO_1773 (O_1773,N_29576,N_29391);
nand UO_1774 (O_1774,N_28663,N_29681);
nor UO_1775 (O_1775,N_28619,N_29628);
or UO_1776 (O_1776,N_28929,N_28555);
and UO_1777 (O_1777,N_28865,N_29639);
nor UO_1778 (O_1778,N_29035,N_29944);
nand UO_1779 (O_1779,N_29602,N_29651);
nor UO_1780 (O_1780,N_29486,N_29844);
and UO_1781 (O_1781,N_29165,N_29344);
and UO_1782 (O_1782,N_29461,N_29761);
nor UO_1783 (O_1783,N_29312,N_28726);
and UO_1784 (O_1784,N_29703,N_29200);
xor UO_1785 (O_1785,N_28915,N_29414);
nor UO_1786 (O_1786,N_29536,N_29361);
nand UO_1787 (O_1787,N_28771,N_29939);
and UO_1788 (O_1788,N_28905,N_29633);
nor UO_1789 (O_1789,N_29983,N_28952);
xor UO_1790 (O_1790,N_29382,N_29875);
or UO_1791 (O_1791,N_29041,N_29292);
nor UO_1792 (O_1792,N_29755,N_29663);
nand UO_1793 (O_1793,N_29945,N_29086);
xnor UO_1794 (O_1794,N_28741,N_28607);
xor UO_1795 (O_1795,N_29401,N_29857);
nand UO_1796 (O_1796,N_28751,N_29602);
and UO_1797 (O_1797,N_28984,N_29096);
nor UO_1798 (O_1798,N_29136,N_28652);
nand UO_1799 (O_1799,N_29969,N_29933);
and UO_1800 (O_1800,N_29617,N_29274);
xor UO_1801 (O_1801,N_29820,N_28514);
xor UO_1802 (O_1802,N_29241,N_29445);
xor UO_1803 (O_1803,N_29496,N_28527);
or UO_1804 (O_1804,N_29911,N_29980);
and UO_1805 (O_1805,N_29603,N_28724);
nand UO_1806 (O_1806,N_29869,N_29357);
nor UO_1807 (O_1807,N_28841,N_28826);
or UO_1808 (O_1808,N_29009,N_29424);
or UO_1809 (O_1809,N_28560,N_29552);
and UO_1810 (O_1810,N_29756,N_28529);
nor UO_1811 (O_1811,N_29122,N_29074);
and UO_1812 (O_1812,N_28822,N_29286);
and UO_1813 (O_1813,N_29620,N_28547);
or UO_1814 (O_1814,N_28502,N_29886);
nor UO_1815 (O_1815,N_28781,N_29674);
and UO_1816 (O_1816,N_28502,N_29530);
and UO_1817 (O_1817,N_29711,N_29431);
nor UO_1818 (O_1818,N_29863,N_29419);
xnor UO_1819 (O_1819,N_29288,N_29506);
xnor UO_1820 (O_1820,N_28583,N_29052);
xor UO_1821 (O_1821,N_29776,N_28819);
nor UO_1822 (O_1822,N_29554,N_29796);
nor UO_1823 (O_1823,N_28563,N_29103);
xor UO_1824 (O_1824,N_29132,N_29035);
nor UO_1825 (O_1825,N_29380,N_29754);
xor UO_1826 (O_1826,N_29027,N_29654);
and UO_1827 (O_1827,N_29433,N_28579);
nor UO_1828 (O_1828,N_28981,N_29426);
nand UO_1829 (O_1829,N_28502,N_29924);
and UO_1830 (O_1830,N_29400,N_29828);
nand UO_1831 (O_1831,N_29657,N_28946);
nor UO_1832 (O_1832,N_29649,N_28842);
nor UO_1833 (O_1833,N_28856,N_29041);
nand UO_1834 (O_1834,N_28535,N_28995);
xnor UO_1835 (O_1835,N_29731,N_28619);
xor UO_1836 (O_1836,N_28589,N_29426);
or UO_1837 (O_1837,N_29759,N_28505);
nand UO_1838 (O_1838,N_28949,N_29141);
or UO_1839 (O_1839,N_28627,N_29542);
and UO_1840 (O_1840,N_29154,N_28538);
nand UO_1841 (O_1841,N_29571,N_28871);
or UO_1842 (O_1842,N_28833,N_29043);
nand UO_1843 (O_1843,N_28774,N_29004);
nand UO_1844 (O_1844,N_29981,N_28581);
nor UO_1845 (O_1845,N_28608,N_28849);
and UO_1846 (O_1846,N_28647,N_28634);
and UO_1847 (O_1847,N_29392,N_29965);
xor UO_1848 (O_1848,N_29938,N_28787);
or UO_1849 (O_1849,N_29334,N_29643);
nor UO_1850 (O_1850,N_28931,N_29043);
or UO_1851 (O_1851,N_29140,N_28982);
nand UO_1852 (O_1852,N_28870,N_28854);
and UO_1853 (O_1853,N_29591,N_29590);
xor UO_1854 (O_1854,N_28630,N_29163);
nand UO_1855 (O_1855,N_28532,N_28718);
and UO_1856 (O_1856,N_29236,N_28526);
and UO_1857 (O_1857,N_29548,N_28590);
xnor UO_1858 (O_1858,N_29703,N_28821);
and UO_1859 (O_1859,N_29194,N_29335);
xnor UO_1860 (O_1860,N_29441,N_28879);
or UO_1861 (O_1861,N_29860,N_29525);
nand UO_1862 (O_1862,N_29983,N_29341);
nand UO_1863 (O_1863,N_28895,N_29528);
nand UO_1864 (O_1864,N_29533,N_28968);
nand UO_1865 (O_1865,N_29221,N_28864);
nor UO_1866 (O_1866,N_29657,N_29416);
nand UO_1867 (O_1867,N_29859,N_29377);
and UO_1868 (O_1868,N_29153,N_29798);
xnor UO_1869 (O_1869,N_28817,N_29992);
and UO_1870 (O_1870,N_28956,N_28900);
and UO_1871 (O_1871,N_28721,N_29193);
xor UO_1872 (O_1872,N_29386,N_28523);
nor UO_1873 (O_1873,N_29449,N_29361);
nand UO_1874 (O_1874,N_29103,N_28825);
or UO_1875 (O_1875,N_29244,N_28509);
nor UO_1876 (O_1876,N_29882,N_29982);
nor UO_1877 (O_1877,N_29218,N_29921);
or UO_1878 (O_1878,N_29619,N_29953);
and UO_1879 (O_1879,N_29038,N_29291);
xnor UO_1880 (O_1880,N_29880,N_29970);
nand UO_1881 (O_1881,N_29386,N_29893);
xor UO_1882 (O_1882,N_29222,N_29899);
or UO_1883 (O_1883,N_29586,N_29199);
nor UO_1884 (O_1884,N_28618,N_28627);
xor UO_1885 (O_1885,N_29721,N_28741);
nand UO_1886 (O_1886,N_28889,N_29840);
nand UO_1887 (O_1887,N_29832,N_29844);
or UO_1888 (O_1888,N_29223,N_28912);
nand UO_1889 (O_1889,N_28629,N_29508);
and UO_1890 (O_1890,N_29746,N_28830);
nor UO_1891 (O_1891,N_28770,N_29698);
xnor UO_1892 (O_1892,N_29812,N_28984);
and UO_1893 (O_1893,N_28559,N_28611);
or UO_1894 (O_1894,N_29815,N_28963);
nand UO_1895 (O_1895,N_28971,N_28764);
and UO_1896 (O_1896,N_29641,N_29243);
and UO_1897 (O_1897,N_28771,N_29781);
xor UO_1898 (O_1898,N_28711,N_29286);
nor UO_1899 (O_1899,N_29916,N_29790);
nor UO_1900 (O_1900,N_29139,N_29734);
nor UO_1901 (O_1901,N_29070,N_28582);
or UO_1902 (O_1902,N_28516,N_29697);
xnor UO_1903 (O_1903,N_28544,N_29318);
and UO_1904 (O_1904,N_28793,N_29671);
or UO_1905 (O_1905,N_29087,N_28908);
nor UO_1906 (O_1906,N_29773,N_29126);
nand UO_1907 (O_1907,N_28725,N_29733);
and UO_1908 (O_1908,N_29097,N_29364);
nor UO_1909 (O_1909,N_29408,N_28631);
and UO_1910 (O_1910,N_28714,N_29703);
xnor UO_1911 (O_1911,N_28952,N_29114);
nor UO_1912 (O_1912,N_29252,N_28853);
or UO_1913 (O_1913,N_29011,N_29852);
xnor UO_1914 (O_1914,N_29408,N_29541);
and UO_1915 (O_1915,N_29469,N_28717);
nor UO_1916 (O_1916,N_28790,N_29090);
xnor UO_1917 (O_1917,N_29368,N_29278);
xor UO_1918 (O_1918,N_29168,N_29495);
nor UO_1919 (O_1919,N_29443,N_29541);
nor UO_1920 (O_1920,N_29876,N_28876);
or UO_1921 (O_1921,N_29445,N_29207);
nand UO_1922 (O_1922,N_29734,N_29706);
nand UO_1923 (O_1923,N_29078,N_28796);
and UO_1924 (O_1924,N_29419,N_28525);
or UO_1925 (O_1925,N_29763,N_29310);
nand UO_1926 (O_1926,N_29711,N_29732);
nor UO_1927 (O_1927,N_29186,N_29967);
nand UO_1928 (O_1928,N_29481,N_29483);
and UO_1929 (O_1929,N_29005,N_29051);
nor UO_1930 (O_1930,N_29272,N_29449);
nor UO_1931 (O_1931,N_29131,N_28938);
nor UO_1932 (O_1932,N_28509,N_29192);
xnor UO_1933 (O_1933,N_29801,N_29175);
xor UO_1934 (O_1934,N_28874,N_28637);
nor UO_1935 (O_1935,N_29322,N_28929);
or UO_1936 (O_1936,N_28693,N_29573);
or UO_1937 (O_1937,N_29076,N_28504);
nor UO_1938 (O_1938,N_29252,N_29251);
xor UO_1939 (O_1939,N_29095,N_28633);
and UO_1940 (O_1940,N_29951,N_29672);
nor UO_1941 (O_1941,N_29136,N_29711);
nor UO_1942 (O_1942,N_28595,N_29716);
nor UO_1943 (O_1943,N_29167,N_29481);
or UO_1944 (O_1944,N_28876,N_28717);
nor UO_1945 (O_1945,N_28722,N_28962);
xnor UO_1946 (O_1946,N_28720,N_28545);
or UO_1947 (O_1947,N_28843,N_28799);
xnor UO_1948 (O_1948,N_29862,N_29831);
nand UO_1949 (O_1949,N_29981,N_29475);
and UO_1950 (O_1950,N_28773,N_29340);
xor UO_1951 (O_1951,N_29328,N_29246);
nor UO_1952 (O_1952,N_29898,N_29000);
or UO_1953 (O_1953,N_28520,N_28719);
or UO_1954 (O_1954,N_29731,N_29095);
nand UO_1955 (O_1955,N_29214,N_29057);
or UO_1956 (O_1956,N_29100,N_29982);
nand UO_1957 (O_1957,N_29593,N_28709);
and UO_1958 (O_1958,N_29271,N_29060);
and UO_1959 (O_1959,N_29664,N_29139);
xnor UO_1960 (O_1960,N_28776,N_29710);
nand UO_1961 (O_1961,N_28623,N_28836);
nor UO_1962 (O_1962,N_28565,N_29733);
nor UO_1963 (O_1963,N_29401,N_29035);
nor UO_1964 (O_1964,N_28526,N_29265);
nand UO_1965 (O_1965,N_29569,N_29247);
nand UO_1966 (O_1966,N_29838,N_29221);
and UO_1967 (O_1967,N_28783,N_29447);
or UO_1968 (O_1968,N_29280,N_28728);
and UO_1969 (O_1969,N_28772,N_29351);
and UO_1970 (O_1970,N_28836,N_28850);
nand UO_1971 (O_1971,N_29309,N_28541);
nand UO_1972 (O_1972,N_29967,N_29299);
and UO_1973 (O_1973,N_28534,N_29441);
nor UO_1974 (O_1974,N_29149,N_29444);
nor UO_1975 (O_1975,N_29068,N_29478);
and UO_1976 (O_1976,N_29118,N_28555);
nor UO_1977 (O_1977,N_29550,N_29204);
or UO_1978 (O_1978,N_29558,N_29965);
nor UO_1979 (O_1979,N_29555,N_29812);
or UO_1980 (O_1980,N_29874,N_29279);
nand UO_1981 (O_1981,N_29995,N_29882);
or UO_1982 (O_1982,N_29130,N_29651);
or UO_1983 (O_1983,N_29951,N_29594);
xor UO_1984 (O_1984,N_29674,N_29097);
xor UO_1985 (O_1985,N_29077,N_29368);
nand UO_1986 (O_1986,N_28792,N_29975);
nor UO_1987 (O_1987,N_28500,N_29414);
and UO_1988 (O_1988,N_28518,N_29003);
nor UO_1989 (O_1989,N_28910,N_29627);
and UO_1990 (O_1990,N_29969,N_28850);
nand UO_1991 (O_1991,N_29050,N_28715);
and UO_1992 (O_1992,N_29385,N_29139);
and UO_1993 (O_1993,N_29316,N_29066);
or UO_1994 (O_1994,N_28683,N_29480);
or UO_1995 (O_1995,N_28622,N_29364);
nor UO_1996 (O_1996,N_28644,N_29784);
and UO_1997 (O_1997,N_29085,N_29529);
or UO_1998 (O_1998,N_29993,N_28910);
nand UO_1999 (O_1999,N_29161,N_29598);
nand UO_2000 (O_2000,N_29581,N_28578);
xor UO_2001 (O_2001,N_28511,N_29701);
nand UO_2002 (O_2002,N_28934,N_29591);
and UO_2003 (O_2003,N_29822,N_28614);
xor UO_2004 (O_2004,N_29511,N_29178);
nand UO_2005 (O_2005,N_29526,N_29247);
nor UO_2006 (O_2006,N_29150,N_29846);
or UO_2007 (O_2007,N_28758,N_29154);
nor UO_2008 (O_2008,N_29110,N_28644);
nor UO_2009 (O_2009,N_28975,N_28935);
xor UO_2010 (O_2010,N_28928,N_28960);
nand UO_2011 (O_2011,N_29928,N_29057);
or UO_2012 (O_2012,N_29578,N_29492);
xnor UO_2013 (O_2013,N_29292,N_29982);
nand UO_2014 (O_2014,N_28664,N_29396);
or UO_2015 (O_2015,N_29796,N_28671);
xor UO_2016 (O_2016,N_28857,N_28866);
xnor UO_2017 (O_2017,N_29298,N_29346);
xnor UO_2018 (O_2018,N_29168,N_29372);
nand UO_2019 (O_2019,N_29142,N_29692);
or UO_2020 (O_2020,N_29649,N_29570);
nor UO_2021 (O_2021,N_29064,N_29493);
and UO_2022 (O_2022,N_29171,N_29020);
nand UO_2023 (O_2023,N_29763,N_28566);
or UO_2024 (O_2024,N_28544,N_29803);
or UO_2025 (O_2025,N_29525,N_29389);
and UO_2026 (O_2026,N_29361,N_29091);
and UO_2027 (O_2027,N_28946,N_29109);
xnor UO_2028 (O_2028,N_29004,N_28847);
and UO_2029 (O_2029,N_29451,N_28808);
or UO_2030 (O_2030,N_28530,N_28825);
or UO_2031 (O_2031,N_29155,N_29273);
or UO_2032 (O_2032,N_29116,N_28749);
xnor UO_2033 (O_2033,N_28833,N_28983);
and UO_2034 (O_2034,N_28861,N_29281);
or UO_2035 (O_2035,N_29050,N_29740);
or UO_2036 (O_2036,N_29625,N_28715);
xor UO_2037 (O_2037,N_28881,N_28625);
nand UO_2038 (O_2038,N_28944,N_28890);
and UO_2039 (O_2039,N_29656,N_29858);
xor UO_2040 (O_2040,N_29835,N_29576);
xor UO_2041 (O_2041,N_29436,N_28723);
nor UO_2042 (O_2042,N_29545,N_29287);
nor UO_2043 (O_2043,N_29410,N_29498);
nor UO_2044 (O_2044,N_29869,N_28799);
nor UO_2045 (O_2045,N_29147,N_28819);
and UO_2046 (O_2046,N_28804,N_29414);
xnor UO_2047 (O_2047,N_28585,N_29584);
nand UO_2048 (O_2048,N_29303,N_29085);
or UO_2049 (O_2049,N_29118,N_29105);
nand UO_2050 (O_2050,N_29776,N_28809);
and UO_2051 (O_2051,N_29252,N_29163);
and UO_2052 (O_2052,N_29225,N_29333);
and UO_2053 (O_2053,N_28996,N_28781);
nor UO_2054 (O_2054,N_29072,N_29320);
xor UO_2055 (O_2055,N_29085,N_29733);
or UO_2056 (O_2056,N_28943,N_29075);
or UO_2057 (O_2057,N_29392,N_29080);
or UO_2058 (O_2058,N_29429,N_28942);
nor UO_2059 (O_2059,N_29579,N_29484);
xnor UO_2060 (O_2060,N_29639,N_29057);
or UO_2061 (O_2061,N_29416,N_29114);
nand UO_2062 (O_2062,N_29762,N_29754);
or UO_2063 (O_2063,N_29116,N_29405);
nand UO_2064 (O_2064,N_29576,N_29642);
nand UO_2065 (O_2065,N_29817,N_29075);
xnor UO_2066 (O_2066,N_29726,N_28566);
nand UO_2067 (O_2067,N_29944,N_28663);
nor UO_2068 (O_2068,N_28962,N_29269);
and UO_2069 (O_2069,N_29478,N_28594);
nor UO_2070 (O_2070,N_29724,N_28580);
and UO_2071 (O_2071,N_29213,N_29979);
nor UO_2072 (O_2072,N_29018,N_28814);
nor UO_2073 (O_2073,N_28554,N_29039);
nor UO_2074 (O_2074,N_29017,N_29846);
nor UO_2075 (O_2075,N_29346,N_28906);
or UO_2076 (O_2076,N_29087,N_29899);
nand UO_2077 (O_2077,N_28970,N_28560);
and UO_2078 (O_2078,N_28847,N_28616);
nand UO_2079 (O_2079,N_29561,N_28507);
or UO_2080 (O_2080,N_29148,N_29123);
nand UO_2081 (O_2081,N_28913,N_29209);
nand UO_2082 (O_2082,N_29000,N_29790);
nor UO_2083 (O_2083,N_29392,N_29516);
and UO_2084 (O_2084,N_29299,N_29715);
and UO_2085 (O_2085,N_28650,N_29087);
and UO_2086 (O_2086,N_28562,N_29376);
nand UO_2087 (O_2087,N_29003,N_29442);
or UO_2088 (O_2088,N_28823,N_28881);
nor UO_2089 (O_2089,N_29216,N_28576);
nand UO_2090 (O_2090,N_29148,N_28601);
nor UO_2091 (O_2091,N_29839,N_28911);
xor UO_2092 (O_2092,N_28733,N_28791);
xor UO_2093 (O_2093,N_28980,N_28651);
nor UO_2094 (O_2094,N_28698,N_29964);
nand UO_2095 (O_2095,N_29256,N_28596);
and UO_2096 (O_2096,N_29711,N_28736);
and UO_2097 (O_2097,N_28712,N_28801);
nor UO_2098 (O_2098,N_29436,N_29589);
nor UO_2099 (O_2099,N_29174,N_29166);
nand UO_2100 (O_2100,N_28748,N_28675);
nor UO_2101 (O_2101,N_28704,N_29671);
xor UO_2102 (O_2102,N_29341,N_28631);
or UO_2103 (O_2103,N_29835,N_29541);
nor UO_2104 (O_2104,N_29797,N_29697);
nand UO_2105 (O_2105,N_28596,N_29162);
or UO_2106 (O_2106,N_29934,N_29430);
or UO_2107 (O_2107,N_29468,N_29269);
xor UO_2108 (O_2108,N_28598,N_29625);
nand UO_2109 (O_2109,N_28923,N_28905);
xnor UO_2110 (O_2110,N_29979,N_28517);
and UO_2111 (O_2111,N_29532,N_29988);
nor UO_2112 (O_2112,N_29747,N_29325);
nand UO_2113 (O_2113,N_29951,N_29688);
and UO_2114 (O_2114,N_29326,N_28702);
nor UO_2115 (O_2115,N_29314,N_29071);
nand UO_2116 (O_2116,N_29673,N_28688);
or UO_2117 (O_2117,N_28800,N_29295);
nand UO_2118 (O_2118,N_29147,N_29444);
nor UO_2119 (O_2119,N_28862,N_29002);
xnor UO_2120 (O_2120,N_29950,N_28503);
and UO_2121 (O_2121,N_29592,N_29431);
nand UO_2122 (O_2122,N_29288,N_28713);
xor UO_2123 (O_2123,N_29099,N_29181);
xor UO_2124 (O_2124,N_29634,N_29909);
xor UO_2125 (O_2125,N_29543,N_29510);
xor UO_2126 (O_2126,N_29039,N_29711);
nor UO_2127 (O_2127,N_28938,N_29650);
nor UO_2128 (O_2128,N_29448,N_29820);
xor UO_2129 (O_2129,N_29055,N_29149);
nor UO_2130 (O_2130,N_29639,N_29928);
xor UO_2131 (O_2131,N_28970,N_28968);
nand UO_2132 (O_2132,N_29506,N_29898);
nor UO_2133 (O_2133,N_28509,N_29603);
xor UO_2134 (O_2134,N_29015,N_29204);
and UO_2135 (O_2135,N_29257,N_29368);
nor UO_2136 (O_2136,N_28824,N_29456);
nand UO_2137 (O_2137,N_29812,N_29349);
xnor UO_2138 (O_2138,N_29745,N_29985);
or UO_2139 (O_2139,N_28676,N_28926);
and UO_2140 (O_2140,N_28648,N_29495);
or UO_2141 (O_2141,N_28506,N_29971);
nor UO_2142 (O_2142,N_29430,N_28806);
xnor UO_2143 (O_2143,N_29121,N_28999);
nand UO_2144 (O_2144,N_29864,N_29376);
xnor UO_2145 (O_2145,N_28885,N_29922);
and UO_2146 (O_2146,N_29574,N_29566);
and UO_2147 (O_2147,N_28791,N_29296);
and UO_2148 (O_2148,N_28987,N_29765);
nand UO_2149 (O_2149,N_28795,N_29568);
nor UO_2150 (O_2150,N_29712,N_28748);
nor UO_2151 (O_2151,N_29582,N_29479);
or UO_2152 (O_2152,N_28551,N_29450);
nand UO_2153 (O_2153,N_29858,N_29690);
xor UO_2154 (O_2154,N_29198,N_28929);
nor UO_2155 (O_2155,N_29190,N_29036);
and UO_2156 (O_2156,N_28741,N_28815);
nand UO_2157 (O_2157,N_29444,N_28872);
or UO_2158 (O_2158,N_29668,N_29487);
nand UO_2159 (O_2159,N_29788,N_29687);
or UO_2160 (O_2160,N_28610,N_29741);
nand UO_2161 (O_2161,N_29862,N_28739);
and UO_2162 (O_2162,N_29079,N_29542);
xor UO_2163 (O_2163,N_29762,N_29889);
nor UO_2164 (O_2164,N_29532,N_29862);
or UO_2165 (O_2165,N_29196,N_29405);
nand UO_2166 (O_2166,N_29064,N_28580);
and UO_2167 (O_2167,N_28843,N_29661);
nor UO_2168 (O_2168,N_29023,N_29027);
nor UO_2169 (O_2169,N_29002,N_28857);
and UO_2170 (O_2170,N_29663,N_29613);
or UO_2171 (O_2171,N_29677,N_29781);
or UO_2172 (O_2172,N_28707,N_28814);
nor UO_2173 (O_2173,N_29604,N_28829);
xnor UO_2174 (O_2174,N_28597,N_29016);
nor UO_2175 (O_2175,N_28884,N_29587);
xor UO_2176 (O_2176,N_29454,N_29094);
xnor UO_2177 (O_2177,N_29523,N_28812);
and UO_2178 (O_2178,N_29162,N_28771);
or UO_2179 (O_2179,N_28879,N_28698);
nor UO_2180 (O_2180,N_29877,N_29175);
nor UO_2181 (O_2181,N_29069,N_29090);
nor UO_2182 (O_2182,N_29600,N_28570);
xnor UO_2183 (O_2183,N_29134,N_29081);
nor UO_2184 (O_2184,N_28518,N_29817);
xnor UO_2185 (O_2185,N_29935,N_28537);
nand UO_2186 (O_2186,N_29434,N_29757);
nand UO_2187 (O_2187,N_29505,N_29707);
xnor UO_2188 (O_2188,N_28666,N_29020);
nand UO_2189 (O_2189,N_28620,N_29132);
nor UO_2190 (O_2190,N_29370,N_29827);
and UO_2191 (O_2191,N_28819,N_29788);
or UO_2192 (O_2192,N_29248,N_29239);
nand UO_2193 (O_2193,N_28815,N_28600);
xor UO_2194 (O_2194,N_28986,N_28893);
nor UO_2195 (O_2195,N_29207,N_28565);
nor UO_2196 (O_2196,N_29111,N_29534);
nor UO_2197 (O_2197,N_29966,N_29469);
or UO_2198 (O_2198,N_29536,N_29795);
or UO_2199 (O_2199,N_29392,N_29172);
and UO_2200 (O_2200,N_29840,N_28534);
nand UO_2201 (O_2201,N_29468,N_28983);
nand UO_2202 (O_2202,N_29429,N_29070);
or UO_2203 (O_2203,N_29960,N_29646);
or UO_2204 (O_2204,N_28820,N_29248);
nor UO_2205 (O_2205,N_28620,N_28595);
nor UO_2206 (O_2206,N_28873,N_29891);
xnor UO_2207 (O_2207,N_29365,N_28587);
nor UO_2208 (O_2208,N_28652,N_29654);
and UO_2209 (O_2209,N_28500,N_29233);
and UO_2210 (O_2210,N_29346,N_28511);
nand UO_2211 (O_2211,N_29113,N_28776);
xor UO_2212 (O_2212,N_29268,N_29794);
or UO_2213 (O_2213,N_29292,N_29101);
nor UO_2214 (O_2214,N_28766,N_29795);
or UO_2215 (O_2215,N_28640,N_29645);
xnor UO_2216 (O_2216,N_29477,N_29287);
and UO_2217 (O_2217,N_28758,N_29207);
xor UO_2218 (O_2218,N_28841,N_29093);
or UO_2219 (O_2219,N_29986,N_29368);
nand UO_2220 (O_2220,N_28860,N_29790);
nand UO_2221 (O_2221,N_29317,N_29517);
nor UO_2222 (O_2222,N_29506,N_29698);
xnor UO_2223 (O_2223,N_28634,N_28733);
or UO_2224 (O_2224,N_28587,N_28507);
nand UO_2225 (O_2225,N_29252,N_29325);
and UO_2226 (O_2226,N_28730,N_29055);
nand UO_2227 (O_2227,N_29031,N_28580);
xor UO_2228 (O_2228,N_29026,N_29113);
or UO_2229 (O_2229,N_29578,N_29387);
nand UO_2230 (O_2230,N_29366,N_28602);
xnor UO_2231 (O_2231,N_28594,N_29464);
and UO_2232 (O_2232,N_28551,N_29323);
nand UO_2233 (O_2233,N_29921,N_28736);
xnor UO_2234 (O_2234,N_29878,N_29599);
and UO_2235 (O_2235,N_28514,N_29517);
nand UO_2236 (O_2236,N_28860,N_29293);
nand UO_2237 (O_2237,N_29181,N_29535);
or UO_2238 (O_2238,N_29779,N_29348);
xor UO_2239 (O_2239,N_29510,N_29236);
or UO_2240 (O_2240,N_28555,N_29648);
or UO_2241 (O_2241,N_28650,N_28588);
nor UO_2242 (O_2242,N_28652,N_29583);
xnor UO_2243 (O_2243,N_29576,N_29962);
nand UO_2244 (O_2244,N_28864,N_28626);
nor UO_2245 (O_2245,N_29314,N_29166);
nor UO_2246 (O_2246,N_29315,N_29773);
or UO_2247 (O_2247,N_29492,N_29021);
nand UO_2248 (O_2248,N_28947,N_29067);
or UO_2249 (O_2249,N_29313,N_29501);
or UO_2250 (O_2250,N_28893,N_29826);
nand UO_2251 (O_2251,N_28750,N_29965);
or UO_2252 (O_2252,N_29847,N_29598);
xnor UO_2253 (O_2253,N_29536,N_28826);
or UO_2254 (O_2254,N_29966,N_29255);
nor UO_2255 (O_2255,N_29706,N_28770);
or UO_2256 (O_2256,N_28582,N_29602);
and UO_2257 (O_2257,N_29192,N_29265);
nor UO_2258 (O_2258,N_29028,N_29068);
or UO_2259 (O_2259,N_29192,N_28996);
nor UO_2260 (O_2260,N_29274,N_28837);
and UO_2261 (O_2261,N_29104,N_29560);
nor UO_2262 (O_2262,N_29948,N_29626);
and UO_2263 (O_2263,N_29707,N_29182);
and UO_2264 (O_2264,N_29831,N_29931);
or UO_2265 (O_2265,N_29671,N_28735);
nor UO_2266 (O_2266,N_29889,N_28909);
nor UO_2267 (O_2267,N_29441,N_28569);
nand UO_2268 (O_2268,N_29915,N_28817);
and UO_2269 (O_2269,N_29092,N_29810);
nand UO_2270 (O_2270,N_29457,N_29583);
xor UO_2271 (O_2271,N_28747,N_29682);
and UO_2272 (O_2272,N_29489,N_29653);
nor UO_2273 (O_2273,N_28775,N_28916);
nand UO_2274 (O_2274,N_29125,N_29848);
or UO_2275 (O_2275,N_28758,N_29643);
and UO_2276 (O_2276,N_28865,N_29542);
nand UO_2277 (O_2277,N_28517,N_29209);
nand UO_2278 (O_2278,N_29029,N_28542);
xnor UO_2279 (O_2279,N_28977,N_29067);
xor UO_2280 (O_2280,N_29929,N_28502);
and UO_2281 (O_2281,N_29894,N_29982);
nand UO_2282 (O_2282,N_29576,N_29488);
xor UO_2283 (O_2283,N_29161,N_28870);
nor UO_2284 (O_2284,N_29699,N_29357);
and UO_2285 (O_2285,N_28883,N_29228);
xnor UO_2286 (O_2286,N_29262,N_29263);
nor UO_2287 (O_2287,N_29256,N_29818);
nor UO_2288 (O_2288,N_28629,N_29567);
nor UO_2289 (O_2289,N_28850,N_29340);
nor UO_2290 (O_2290,N_29382,N_28825);
or UO_2291 (O_2291,N_29839,N_29220);
xor UO_2292 (O_2292,N_28807,N_29206);
nand UO_2293 (O_2293,N_29920,N_29402);
and UO_2294 (O_2294,N_29175,N_28877);
and UO_2295 (O_2295,N_28602,N_29959);
nor UO_2296 (O_2296,N_29132,N_29684);
or UO_2297 (O_2297,N_28608,N_29488);
or UO_2298 (O_2298,N_29470,N_29935);
xnor UO_2299 (O_2299,N_29961,N_29386);
or UO_2300 (O_2300,N_29414,N_29933);
nor UO_2301 (O_2301,N_29794,N_28842);
nor UO_2302 (O_2302,N_29068,N_29636);
xor UO_2303 (O_2303,N_29708,N_28852);
or UO_2304 (O_2304,N_29742,N_29655);
nand UO_2305 (O_2305,N_29604,N_29579);
and UO_2306 (O_2306,N_28642,N_28769);
nand UO_2307 (O_2307,N_29678,N_28606);
and UO_2308 (O_2308,N_28726,N_29543);
nand UO_2309 (O_2309,N_28530,N_29031);
xnor UO_2310 (O_2310,N_28593,N_29695);
or UO_2311 (O_2311,N_29687,N_29333);
nor UO_2312 (O_2312,N_29611,N_28671);
xnor UO_2313 (O_2313,N_29856,N_29066);
xor UO_2314 (O_2314,N_28753,N_28877);
nand UO_2315 (O_2315,N_29490,N_29508);
nand UO_2316 (O_2316,N_29487,N_29844);
xor UO_2317 (O_2317,N_29329,N_28825);
and UO_2318 (O_2318,N_29712,N_29045);
xor UO_2319 (O_2319,N_28905,N_29261);
xnor UO_2320 (O_2320,N_28895,N_29699);
and UO_2321 (O_2321,N_28692,N_29519);
nor UO_2322 (O_2322,N_28993,N_29758);
xor UO_2323 (O_2323,N_29551,N_28581);
nand UO_2324 (O_2324,N_29838,N_29114);
nor UO_2325 (O_2325,N_29545,N_29181);
nand UO_2326 (O_2326,N_29645,N_28917);
nand UO_2327 (O_2327,N_29969,N_29417);
xor UO_2328 (O_2328,N_29603,N_29888);
or UO_2329 (O_2329,N_29565,N_28765);
nor UO_2330 (O_2330,N_29126,N_29184);
and UO_2331 (O_2331,N_29501,N_29490);
and UO_2332 (O_2332,N_28952,N_29438);
and UO_2333 (O_2333,N_29345,N_28772);
nor UO_2334 (O_2334,N_29447,N_29762);
nor UO_2335 (O_2335,N_29183,N_28949);
or UO_2336 (O_2336,N_29655,N_28699);
xor UO_2337 (O_2337,N_28920,N_29185);
or UO_2338 (O_2338,N_28626,N_29310);
and UO_2339 (O_2339,N_28574,N_29478);
and UO_2340 (O_2340,N_28907,N_29216);
nand UO_2341 (O_2341,N_29502,N_28712);
and UO_2342 (O_2342,N_29335,N_29635);
nor UO_2343 (O_2343,N_29784,N_29956);
nor UO_2344 (O_2344,N_29746,N_29229);
xnor UO_2345 (O_2345,N_28955,N_28718);
nor UO_2346 (O_2346,N_28525,N_29868);
nand UO_2347 (O_2347,N_28601,N_29150);
nand UO_2348 (O_2348,N_28716,N_29972);
nand UO_2349 (O_2349,N_29730,N_29448);
or UO_2350 (O_2350,N_29462,N_28551);
and UO_2351 (O_2351,N_29498,N_28655);
xor UO_2352 (O_2352,N_29211,N_29069);
or UO_2353 (O_2353,N_29404,N_29889);
and UO_2354 (O_2354,N_29439,N_29860);
or UO_2355 (O_2355,N_29284,N_29738);
nand UO_2356 (O_2356,N_29506,N_29172);
and UO_2357 (O_2357,N_28555,N_29477);
nand UO_2358 (O_2358,N_29429,N_28827);
and UO_2359 (O_2359,N_29518,N_29770);
nor UO_2360 (O_2360,N_28758,N_29935);
nand UO_2361 (O_2361,N_29558,N_28837);
xnor UO_2362 (O_2362,N_28756,N_29256);
and UO_2363 (O_2363,N_29784,N_28578);
nor UO_2364 (O_2364,N_29362,N_29665);
nor UO_2365 (O_2365,N_29575,N_29042);
or UO_2366 (O_2366,N_28562,N_29224);
or UO_2367 (O_2367,N_28904,N_29380);
nand UO_2368 (O_2368,N_29680,N_29018);
or UO_2369 (O_2369,N_29288,N_29611);
and UO_2370 (O_2370,N_29481,N_29064);
nand UO_2371 (O_2371,N_28666,N_29242);
nor UO_2372 (O_2372,N_28726,N_29688);
nor UO_2373 (O_2373,N_28742,N_28754);
nor UO_2374 (O_2374,N_29778,N_29883);
nand UO_2375 (O_2375,N_29250,N_29426);
or UO_2376 (O_2376,N_29290,N_28788);
nor UO_2377 (O_2377,N_29066,N_29972);
xor UO_2378 (O_2378,N_29254,N_29256);
nand UO_2379 (O_2379,N_29574,N_29041);
nand UO_2380 (O_2380,N_29061,N_29228);
nor UO_2381 (O_2381,N_28508,N_29477);
nand UO_2382 (O_2382,N_29830,N_28748);
nand UO_2383 (O_2383,N_29223,N_29440);
nor UO_2384 (O_2384,N_29119,N_29591);
and UO_2385 (O_2385,N_29320,N_28703);
and UO_2386 (O_2386,N_28730,N_29332);
nor UO_2387 (O_2387,N_29818,N_29793);
xnor UO_2388 (O_2388,N_28774,N_29235);
xnor UO_2389 (O_2389,N_28598,N_29085);
xnor UO_2390 (O_2390,N_29101,N_28993);
nand UO_2391 (O_2391,N_29121,N_29544);
and UO_2392 (O_2392,N_28836,N_29157);
nor UO_2393 (O_2393,N_29927,N_29118);
nor UO_2394 (O_2394,N_28614,N_28964);
and UO_2395 (O_2395,N_29967,N_28736);
xor UO_2396 (O_2396,N_29336,N_29307);
nand UO_2397 (O_2397,N_29743,N_29948);
xnor UO_2398 (O_2398,N_28563,N_29500);
nor UO_2399 (O_2399,N_28528,N_28935);
nand UO_2400 (O_2400,N_28785,N_29423);
or UO_2401 (O_2401,N_29324,N_29813);
nor UO_2402 (O_2402,N_29255,N_29917);
and UO_2403 (O_2403,N_29706,N_29575);
xor UO_2404 (O_2404,N_29760,N_29148);
xnor UO_2405 (O_2405,N_29372,N_29265);
or UO_2406 (O_2406,N_28983,N_29460);
nand UO_2407 (O_2407,N_29614,N_29989);
and UO_2408 (O_2408,N_28937,N_29811);
nand UO_2409 (O_2409,N_29067,N_29540);
nor UO_2410 (O_2410,N_28996,N_29366);
nor UO_2411 (O_2411,N_28978,N_29081);
and UO_2412 (O_2412,N_29616,N_28625);
xor UO_2413 (O_2413,N_29718,N_28839);
nand UO_2414 (O_2414,N_29627,N_28671);
and UO_2415 (O_2415,N_29002,N_29460);
xnor UO_2416 (O_2416,N_29740,N_29216);
nand UO_2417 (O_2417,N_28534,N_29555);
xor UO_2418 (O_2418,N_29063,N_28698);
nor UO_2419 (O_2419,N_28946,N_28622);
and UO_2420 (O_2420,N_28917,N_29361);
or UO_2421 (O_2421,N_29884,N_29938);
nor UO_2422 (O_2422,N_29087,N_29600);
xnor UO_2423 (O_2423,N_29727,N_29958);
and UO_2424 (O_2424,N_29839,N_29528);
or UO_2425 (O_2425,N_29889,N_28601);
or UO_2426 (O_2426,N_29910,N_29601);
xor UO_2427 (O_2427,N_28594,N_29418);
and UO_2428 (O_2428,N_29415,N_29180);
nor UO_2429 (O_2429,N_29607,N_28761);
nand UO_2430 (O_2430,N_28529,N_29802);
nor UO_2431 (O_2431,N_29436,N_29780);
and UO_2432 (O_2432,N_28778,N_28696);
nand UO_2433 (O_2433,N_29228,N_29079);
xor UO_2434 (O_2434,N_28771,N_28910);
xor UO_2435 (O_2435,N_28732,N_29381);
or UO_2436 (O_2436,N_28555,N_28514);
and UO_2437 (O_2437,N_28781,N_28853);
nand UO_2438 (O_2438,N_29808,N_29455);
nor UO_2439 (O_2439,N_29528,N_28970);
nor UO_2440 (O_2440,N_29095,N_29872);
nand UO_2441 (O_2441,N_29090,N_29990);
xnor UO_2442 (O_2442,N_29410,N_29809);
nor UO_2443 (O_2443,N_29233,N_29558);
nand UO_2444 (O_2444,N_29022,N_28741);
or UO_2445 (O_2445,N_28676,N_28713);
nor UO_2446 (O_2446,N_29478,N_29186);
xnor UO_2447 (O_2447,N_28511,N_29160);
nor UO_2448 (O_2448,N_29305,N_28605);
nand UO_2449 (O_2449,N_29323,N_29968);
nor UO_2450 (O_2450,N_28781,N_28573);
nor UO_2451 (O_2451,N_28786,N_28773);
or UO_2452 (O_2452,N_28890,N_29089);
and UO_2453 (O_2453,N_28693,N_28889);
xnor UO_2454 (O_2454,N_29641,N_28529);
nand UO_2455 (O_2455,N_29876,N_29221);
and UO_2456 (O_2456,N_29772,N_29126);
xnor UO_2457 (O_2457,N_29254,N_29940);
nor UO_2458 (O_2458,N_28708,N_29763);
or UO_2459 (O_2459,N_28882,N_29128);
and UO_2460 (O_2460,N_29084,N_28583);
or UO_2461 (O_2461,N_29408,N_29274);
and UO_2462 (O_2462,N_29865,N_29589);
and UO_2463 (O_2463,N_29785,N_29893);
nor UO_2464 (O_2464,N_29825,N_28829);
xnor UO_2465 (O_2465,N_29393,N_28843);
nand UO_2466 (O_2466,N_29734,N_29071);
xor UO_2467 (O_2467,N_29804,N_29657);
nor UO_2468 (O_2468,N_29966,N_29919);
and UO_2469 (O_2469,N_28859,N_29416);
nor UO_2470 (O_2470,N_29749,N_29818);
xor UO_2471 (O_2471,N_28900,N_29038);
nor UO_2472 (O_2472,N_29970,N_29431);
xor UO_2473 (O_2473,N_29239,N_29985);
nor UO_2474 (O_2474,N_29215,N_29759);
nand UO_2475 (O_2475,N_29556,N_29358);
nor UO_2476 (O_2476,N_29851,N_28824);
and UO_2477 (O_2477,N_29014,N_28540);
xnor UO_2478 (O_2478,N_28724,N_29399);
nand UO_2479 (O_2479,N_28869,N_29036);
nand UO_2480 (O_2480,N_28600,N_28990);
and UO_2481 (O_2481,N_29775,N_29646);
or UO_2482 (O_2482,N_29871,N_28725);
and UO_2483 (O_2483,N_29223,N_28778);
nor UO_2484 (O_2484,N_29340,N_28611);
nor UO_2485 (O_2485,N_28833,N_29851);
nor UO_2486 (O_2486,N_29949,N_29603);
and UO_2487 (O_2487,N_29442,N_29959);
and UO_2488 (O_2488,N_29418,N_29423);
and UO_2489 (O_2489,N_29371,N_29387);
xor UO_2490 (O_2490,N_29575,N_28773);
nand UO_2491 (O_2491,N_29177,N_29084);
nor UO_2492 (O_2492,N_29422,N_29999);
xor UO_2493 (O_2493,N_29729,N_29831);
nor UO_2494 (O_2494,N_29945,N_29454);
or UO_2495 (O_2495,N_29268,N_29505);
xnor UO_2496 (O_2496,N_28816,N_29879);
nand UO_2497 (O_2497,N_29565,N_29863);
or UO_2498 (O_2498,N_28764,N_29289);
nor UO_2499 (O_2499,N_28820,N_29524);
nand UO_2500 (O_2500,N_29046,N_28594);
or UO_2501 (O_2501,N_29957,N_28602);
xnor UO_2502 (O_2502,N_29753,N_29170);
nand UO_2503 (O_2503,N_29419,N_28768);
or UO_2504 (O_2504,N_29908,N_28617);
and UO_2505 (O_2505,N_28969,N_29274);
or UO_2506 (O_2506,N_29467,N_29615);
or UO_2507 (O_2507,N_29976,N_29430);
nand UO_2508 (O_2508,N_29003,N_29731);
nand UO_2509 (O_2509,N_28862,N_29802);
xnor UO_2510 (O_2510,N_29810,N_29095);
nor UO_2511 (O_2511,N_29845,N_29510);
and UO_2512 (O_2512,N_29509,N_29956);
or UO_2513 (O_2513,N_29295,N_29860);
nand UO_2514 (O_2514,N_29738,N_29657);
nand UO_2515 (O_2515,N_29907,N_28891);
nor UO_2516 (O_2516,N_28649,N_28898);
or UO_2517 (O_2517,N_29203,N_28534);
xnor UO_2518 (O_2518,N_29578,N_28529);
or UO_2519 (O_2519,N_29211,N_29230);
or UO_2520 (O_2520,N_29282,N_29458);
or UO_2521 (O_2521,N_29885,N_29282);
xnor UO_2522 (O_2522,N_29475,N_28745);
xnor UO_2523 (O_2523,N_29658,N_29074);
xor UO_2524 (O_2524,N_29040,N_29952);
or UO_2525 (O_2525,N_29540,N_29718);
xor UO_2526 (O_2526,N_29312,N_29731);
nand UO_2527 (O_2527,N_29567,N_29187);
nand UO_2528 (O_2528,N_28828,N_29194);
xnor UO_2529 (O_2529,N_28527,N_28510);
or UO_2530 (O_2530,N_29332,N_29338);
or UO_2531 (O_2531,N_29883,N_29954);
and UO_2532 (O_2532,N_29997,N_28720);
xor UO_2533 (O_2533,N_29996,N_29860);
or UO_2534 (O_2534,N_29971,N_29062);
xnor UO_2535 (O_2535,N_28594,N_29121);
or UO_2536 (O_2536,N_29864,N_28850);
nor UO_2537 (O_2537,N_28736,N_29493);
nor UO_2538 (O_2538,N_29718,N_29238);
nor UO_2539 (O_2539,N_29976,N_29830);
nor UO_2540 (O_2540,N_29155,N_29412);
and UO_2541 (O_2541,N_29249,N_29214);
nor UO_2542 (O_2542,N_29425,N_28992);
and UO_2543 (O_2543,N_29035,N_28991);
and UO_2544 (O_2544,N_29406,N_29214);
or UO_2545 (O_2545,N_28750,N_29223);
nor UO_2546 (O_2546,N_28645,N_28780);
nor UO_2547 (O_2547,N_28902,N_29361);
nand UO_2548 (O_2548,N_28825,N_29350);
or UO_2549 (O_2549,N_29921,N_28791);
and UO_2550 (O_2550,N_29224,N_29767);
nor UO_2551 (O_2551,N_29466,N_29893);
nor UO_2552 (O_2552,N_29542,N_29919);
nor UO_2553 (O_2553,N_28553,N_29366);
or UO_2554 (O_2554,N_29466,N_29080);
and UO_2555 (O_2555,N_28950,N_29755);
nand UO_2556 (O_2556,N_29449,N_29334);
or UO_2557 (O_2557,N_29207,N_28705);
and UO_2558 (O_2558,N_29034,N_29171);
xnor UO_2559 (O_2559,N_29343,N_29805);
and UO_2560 (O_2560,N_28963,N_29424);
nand UO_2561 (O_2561,N_29316,N_28720);
or UO_2562 (O_2562,N_28666,N_29768);
or UO_2563 (O_2563,N_28975,N_29950);
nor UO_2564 (O_2564,N_29088,N_28546);
or UO_2565 (O_2565,N_29390,N_28503);
nand UO_2566 (O_2566,N_29204,N_28679);
or UO_2567 (O_2567,N_29111,N_29130);
and UO_2568 (O_2568,N_28886,N_29023);
xnor UO_2569 (O_2569,N_29805,N_29344);
xor UO_2570 (O_2570,N_29188,N_29591);
xnor UO_2571 (O_2571,N_29480,N_29654);
nand UO_2572 (O_2572,N_29434,N_29844);
nor UO_2573 (O_2573,N_29231,N_29977);
nand UO_2574 (O_2574,N_29272,N_29044);
or UO_2575 (O_2575,N_29991,N_28785);
nand UO_2576 (O_2576,N_29096,N_29408);
and UO_2577 (O_2577,N_28709,N_28648);
or UO_2578 (O_2578,N_29980,N_29959);
nor UO_2579 (O_2579,N_29305,N_28622);
nor UO_2580 (O_2580,N_28992,N_29875);
and UO_2581 (O_2581,N_29641,N_29262);
nand UO_2582 (O_2582,N_28539,N_29657);
or UO_2583 (O_2583,N_28802,N_29289);
and UO_2584 (O_2584,N_28934,N_29451);
nand UO_2585 (O_2585,N_29530,N_29449);
xnor UO_2586 (O_2586,N_29013,N_29757);
and UO_2587 (O_2587,N_29225,N_28671);
nor UO_2588 (O_2588,N_28689,N_28589);
nor UO_2589 (O_2589,N_29499,N_29264);
or UO_2590 (O_2590,N_28947,N_29472);
xnor UO_2591 (O_2591,N_29522,N_29253);
nor UO_2592 (O_2592,N_28623,N_29927);
xor UO_2593 (O_2593,N_29173,N_28661);
or UO_2594 (O_2594,N_29876,N_29510);
or UO_2595 (O_2595,N_29789,N_29084);
or UO_2596 (O_2596,N_28603,N_29609);
and UO_2597 (O_2597,N_29722,N_29677);
or UO_2598 (O_2598,N_28555,N_28834);
nor UO_2599 (O_2599,N_29506,N_29027);
xnor UO_2600 (O_2600,N_28758,N_28536);
nor UO_2601 (O_2601,N_29535,N_28553);
nand UO_2602 (O_2602,N_28501,N_28508);
and UO_2603 (O_2603,N_29536,N_28838);
nor UO_2604 (O_2604,N_29987,N_29896);
or UO_2605 (O_2605,N_28826,N_28666);
nand UO_2606 (O_2606,N_29686,N_29700);
xnor UO_2607 (O_2607,N_29337,N_29297);
nand UO_2608 (O_2608,N_28762,N_29716);
or UO_2609 (O_2609,N_29729,N_28548);
or UO_2610 (O_2610,N_29332,N_28578);
or UO_2611 (O_2611,N_29904,N_29274);
and UO_2612 (O_2612,N_28521,N_29697);
and UO_2613 (O_2613,N_28840,N_29491);
nand UO_2614 (O_2614,N_29202,N_29569);
or UO_2615 (O_2615,N_29424,N_29967);
nor UO_2616 (O_2616,N_28840,N_29650);
and UO_2617 (O_2617,N_28549,N_29503);
xor UO_2618 (O_2618,N_29811,N_29216);
or UO_2619 (O_2619,N_29061,N_29430);
nor UO_2620 (O_2620,N_28673,N_29304);
and UO_2621 (O_2621,N_29220,N_29042);
or UO_2622 (O_2622,N_29170,N_29124);
xor UO_2623 (O_2623,N_29762,N_28784);
nor UO_2624 (O_2624,N_28686,N_29147);
xnor UO_2625 (O_2625,N_29786,N_29047);
or UO_2626 (O_2626,N_29013,N_28889);
nor UO_2627 (O_2627,N_28707,N_29808);
nand UO_2628 (O_2628,N_28893,N_29432);
nand UO_2629 (O_2629,N_29609,N_29650);
and UO_2630 (O_2630,N_29534,N_28834);
or UO_2631 (O_2631,N_29588,N_29751);
and UO_2632 (O_2632,N_29089,N_29290);
nand UO_2633 (O_2633,N_28757,N_29195);
nand UO_2634 (O_2634,N_28873,N_28840);
xnor UO_2635 (O_2635,N_29959,N_29755);
nand UO_2636 (O_2636,N_28756,N_29514);
xnor UO_2637 (O_2637,N_29773,N_29573);
xor UO_2638 (O_2638,N_29801,N_29537);
xor UO_2639 (O_2639,N_29772,N_29530);
and UO_2640 (O_2640,N_29888,N_28813);
nand UO_2641 (O_2641,N_28780,N_29298);
and UO_2642 (O_2642,N_28665,N_29309);
or UO_2643 (O_2643,N_28838,N_29351);
or UO_2644 (O_2644,N_28813,N_28987);
nand UO_2645 (O_2645,N_29883,N_29904);
or UO_2646 (O_2646,N_29706,N_29390);
xnor UO_2647 (O_2647,N_28649,N_28904);
and UO_2648 (O_2648,N_28827,N_29752);
nor UO_2649 (O_2649,N_29407,N_28756);
nand UO_2650 (O_2650,N_28796,N_29999);
xnor UO_2651 (O_2651,N_28801,N_29534);
or UO_2652 (O_2652,N_29727,N_29175);
and UO_2653 (O_2653,N_29794,N_29653);
and UO_2654 (O_2654,N_29752,N_28773);
and UO_2655 (O_2655,N_28507,N_28756);
xor UO_2656 (O_2656,N_29585,N_29664);
xnor UO_2657 (O_2657,N_29747,N_28833);
nand UO_2658 (O_2658,N_28662,N_29548);
nor UO_2659 (O_2659,N_28543,N_28830);
and UO_2660 (O_2660,N_29144,N_29981);
xnor UO_2661 (O_2661,N_29397,N_29654);
nand UO_2662 (O_2662,N_29818,N_28918);
xor UO_2663 (O_2663,N_29494,N_29382);
nor UO_2664 (O_2664,N_29371,N_29944);
nor UO_2665 (O_2665,N_28686,N_29488);
xor UO_2666 (O_2666,N_29406,N_29241);
nor UO_2667 (O_2667,N_28843,N_28533);
nand UO_2668 (O_2668,N_28966,N_29026);
or UO_2669 (O_2669,N_29486,N_28921);
xor UO_2670 (O_2670,N_29075,N_29326);
nor UO_2671 (O_2671,N_28768,N_28806);
xor UO_2672 (O_2672,N_29000,N_29715);
nand UO_2673 (O_2673,N_29246,N_29141);
and UO_2674 (O_2674,N_29095,N_28621);
nand UO_2675 (O_2675,N_28837,N_28884);
or UO_2676 (O_2676,N_29851,N_28874);
or UO_2677 (O_2677,N_28753,N_29853);
nor UO_2678 (O_2678,N_29941,N_29675);
or UO_2679 (O_2679,N_29696,N_29449);
nor UO_2680 (O_2680,N_28558,N_28942);
or UO_2681 (O_2681,N_29351,N_29938);
xnor UO_2682 (O_2682,N_29831,N_28657);
nand UO_2683 (O_2683,N_28658,N_28675);
nand UO_2684 (O_2684,N_29703,N_29677);
or UO_2685 (O_2685,N_29915,N_29752);
nor UO_2686 (O_2686,N_29318,N_28502);
or UO_2687 (O_2687,N_29016,N_28900);
and UO_2688 (O_2688,N_29851,N_29874);
or UO_2689 (O_2689,N_28877,N_29793);
or UO_2690 (O_2690,N_29391,N_28928);
or UO_2691 (O_2691,N_29368,N_29939);
xor UO_2692 (O_2692,N_28572,N_29400);
or UO_2693 (O_2693,N_28875,N_29104);
xor UO_2694 (O_2694,N_29758,N_28603);
xor UO_2695 (O_2695,N_29477,N_28631);
xor UO_2696 (O_2696,N_29116,N_29576);
xor UO_2697 (O_2697,N_28734,N_29907);
nand UO_2698 (O_2698,N_28851,N_28670);
nor UO_2699 (O_2699,N_29489,N_29499);
and UO_2700 (O_2700,N_29410,N_28812);
xor UO_2701 (O_2701,N_29531,N_29080);
nor UO_2702 (O_2702,N_28860,N_29863);
xor UO_2703 (O_2703,N_28812,N_28977);
nor UO_2704 (O_2704,N_29756,N_29053);
nor UO_2705 (O_2705,N_29419,N_29474);
xor UO_2706 (O_2706,N_29759,N_28920);
xor UO_2707 (O_2707,N_29251,N_29185);
nand UO_2708 (O_2708,N_29426,N_29324);
xnor UO_2709 (O_2709,N_29926,N_29000);
or UO_2710 (O_2710,N_29500,N_28871);
nor UO_2711 (O_2711,N_29638,N_29073);
nor UO_2712 (O_2712,N_28791,N_28559);
nand UO_2713 (O_2713,N_29110,N_28798);
xor UO_2714 (O_2714,N_28894,N_28736);
or UO_2715 (O_2715,N_29126,N_29906);
nand UO_2716 (O_2716,N_29666,N_28841);
nand UO_2717 (O_2717,N_28858,N_28821);
nand UO_2718 (O_2718,N_28697,N_29243);
xnor UO_2719 (O_2719,N_29488,N_29562);
nor UO_2720 (O_2720,N_29914,N_29924);
or UO_2721 (O_2721,N_29263,N_29752);
nor UO_2722 (O_2722,N_29536,N_28828);
xor UO_2723 (O_2723,N_28687,N_29611);
or UO_2724 (O_2724,N_29484,N_28696);
and UO_2725 (O_2725,N_29822,N_29878);
nor UO_2726 (O_2726,N_29579,N_28628);
nand UO_2727 (O_2727,N_28815,N_28594);
nor UO_2728 (O_2728,N_29321,N_29730);
and UO_2729 (O_2729,N_29674,N_28697);
xnor UO_2730 (O_2730,N_28927,N_29603);
nor UO_2731 (O_2731,N_29085,N_29040);
xor UO_2732 (O_2732,N_29153,N_29556);
and UO_2733 (O_2733,N_29083,N_28891);
nor UO_2734 (O_2734,N_28591,N_29451);
nor UO_2735 (O_2735,N_29564,N_29464);
xnor UO_2736 (O_2736,N_29441,N_28884);
nand UO_2737 (O_2737,N_29136,N_28927);
xor UO_2738 (O_2738,N_29049,N_29544);
nor UO_2739 (O_2739,N_29147,N_28611);
and UO_2740 (O_2740,N_29261,N_28561);
or UO_2741 (O_2741,N_29365,N_28518);
or UO_2742 (O_2742,N_29390,N_29473);
or UO_2743 (O_2743,N_28550,N_29417);
xnor UO_2744 (O_2744,N_29096,N_29845);
or UO_2745 (O_2745,N_29552,N_29158);
and UO_2746 (O_2746,N_29802,N_29976);
and UO_2747 (O_2747,N_29783,N_29116);
nand UO_2748 (O_2748,N_29879,N_29315);
xnor UO_2749 (O_2749,N_29342,N_28791);
nor UO_2750 (O_2750,N_29679,N_29585);
nand UO_2751 (O_2751,N_29157,N_28843);
xor UO_2752 (O_2752,N_28556,N_28695);
nor UO_2753 (O_2753,N_29700,N_28556);
and UO_2754 (O_2754,N_29802,N_29993);
xnor UO_2755 (O_2755,N_29450,N_28902);
nor UO_2756 (O_2756,N_29071,N_29310);
or UO_2757 (O_2757,N_28612,N_29798);
nand UO_2758 (O_2758,N_29139,N_28688);
and UO_2759 (O_2759,N_29814,N_28775);
and UO_2760 (O_2760,N_29871,N_28787);
and UO_2761 (O_2761,N_28574,N_29337);
or UO_2762 (O_2762,N_29822,N_29556);
and UO_2763 (O_2763,N_29769,N_28591);
nor UO_2764 (O_2764,N_29028,N_29319);
or UO_2765 (O_2765,N_28612,N_28777);
nor UO_2766 (O_2766,N_29312,N_29946);
or UO_2767 (O_2767,N_28836,N_29851);
nor UO_2768 (O_2768,N_28819,N_29987);
or UO_2769 (O_2769,N_29478,N_29008);
xor UO_2770 (O_2770,N_28889,N_29889);
nor UO_2771 (O_2771,N_28978,N_29133);
or UO_2772 (O_2772,N_29026,N_28505);
nand UO_2773 (O_2773,N_29854,N_29395);
and UO_2774 (O_2774,N_29094,N_28974);
or UO_2775 (O_2775,N_29808,N_29092);
nor UO_2776 (O_2776,N_29184,N_29364);
and UO_2777 (O_2777,N_29129,N_29682);
nor UO_2778 (O_2778,N_28697,N_29732);
and UO_2779 (O_2779,N_28816,N_29481);
nor UO_2780 (O_2780,N_29392,N_29945);
nand UO_2781 (O_2781,N_29923,N_28935);
and UO_2782 (O_2782,N_28783,N_29366);
nor UO_2783 (O_2783,N_29223,N_28715);
nor UO_2784 (O_2784,N_29560,N_29093);
and UO_2785 (O_2785,N_28901,N_28754);
xor UO_2786 (O_2786,N_29031,N_29677);
or UO_2787 (O_2787,N_28562,N_29564);
nor UO_2788 (O_2788,N_29247,N_29695);
xnor UO_2789 (O_2789,N_28942,N_29147);
or UO_2790 (O_2790,N_29587,N_29963);
or UO_2791 (O_2791,N_29695,N_29719);
nand UO_2792 (O_2792,N_29913,N_29933);
nand UO_2793 (O_2793,N_29539,N_28979);
nand UO_2794 (O_2794,N_29905,N_29796);
and UO_2795 (O_2795,N_29922,N_29237);
and UO_2796 (O_2796,N_28840,N_29888);
nor UO_2797 (O_2797,N_29621,N_29180);
or UO_2798 (O_2798,N_28513,N_29681);
nand UO_2799 (O_2799,N_28588,N_29706);
xor UO_2800 (O_2800,N_29660,N_29121);
nor UO_2801 (O_2801,N_28649,N_29038);
and UO_2802 (O_2802,N_29897,N_29902);
and UO_2803 (O_2803,N_28532,N_29862);
nor UO_2804 (O_2804,N_29972,N_29803);
nor UO_2805 (O_2805,N_29028,N_29862);
nor UO_2806 (O_2806,N_29974,N_29388);
xnor UO_2807 (O_2807,N_29039,N_29409);
nand UO_2808 (O_2808,N_29197,N_29300);
xor UO_2809 (O_2809,N_29013,N_29035);
or UO_2810 (O_2810,N_28684,N_28634);
xnor UO_2811 (O_2811,N_28957,N_29295);
nand UO_2812 (O_2812,N_29906,N_28944);
nand UO_2813 (O_2813,N_29080,N_29526);
nand UO_2814 (O_2814,N_28880,N_29429);
or UO_2815 (O_2815,N_28753,N_29622);
and UO_2816 (O_2816,N_28742,N_29474);
nor UO_2817 (O_2817,N_29821,N_28800);
xnor UO_2818 (O_2818,N_29355,N_29385);
or UO_2819 (O_2819,N_29491,N_29709);
nor UO_2820 (O_2820,N_28808,N_29469);
xnor UO_2821 (O_2821,N_28899,N_28805);
nand UO_2822 (O_2822,N_29344,N_29679);
and UO_2823 (O_2823,N_29890,N_29566);
nor UO_2824 (O_2824,N_28511,N_28811);
xor UO_2825 (O_2825,N_29573,N_28721);
nand UO_2826 (O_2826,N_29568,N_28789);
and UO_2827 (O_2827,N_28720,N_28921);
nor UO_2828 (O_2828,N_29280,N_28540);
nand UO_2829 (O_2829,N_28532,N_29342);
nor UO_2830 (O_2830,N_29948,N_29186);
and UO_2831 (O_2831,N_28776,N_28870);
nand UO_2832 (O_2832,N_29369,N_29327);
nand UO_2833 (O_2833,N_29855,N_28514);
xnor UO_2834 (O_2834,N_29219,N_29886);
nand UO_2835 (O_2835,N_29894,N_29864);
and UO_2836 (O_2836,N_29254,N_28599);
xnor UO_2837 (O_2837,N_28712,N_29681);
xnor UO_2838 (O_2838,N_28773,N_29942);
nor UO_2839 (O_2839,N_29546,N_29878);
nand UO_2840 (O_2840,N_28763,N_28618);
nor UO_2841 (O_2841,N_28756,N_29021);
or UO_2842 (O_2842,N_29901,N_29190);
nor UO_2843 (O_2843,N_28559,N_29193);
nand UO_2844 (O_2844,N_28675,N_28933);
or UO_2845 (O_2845,N_29306,N_28651);
nor UO_2846 (O_2846,N_29613,N_28761);
xor UO_2847 (O_2847,N_28965,N_29316);
or UO_2848 (O_2848,N_28707,N_29996);
and UO_2849 (O_2849,N_29946,N_28846);
nor UO_2850 (O_2850,N_28747,N_29955);
and UO_2851 (O_2851,N_29330,N_28591);
nand UO_2852 (O_2852,N_28990,N_29480);
or UO_2853 (O_2853,N_29009,N_29709);
xnor UO_2854 (O_2854,N_29701,N_29608);
xnor UO_2855 (O_2855,N_28839,N_29467);
nor UO_2856 (O_2856,N_28889,N_29189);
xor UO_2857 (O_2857,N_29978,N_29124);
or UO_2858 (O_2858,N_29294,N_28551);
nor UO_2859 (O_2859,N_28900,N_29478);
and UO_2860 (O_2860,N_28655,N_29390);
nor UO_2861 (O_2861,N_29504,N_29524);
xor UO_2862 (O_2862,N_29628,N_28640);
nand UO_2863 (O_2863,N_29260,N_29654);
and UO_2864 (O_2864,N_29317,N_28579);
nand UO_2865 (O_2865,N_29432,N_29406);
nor UO_2866 (O_2866,N_29245,N_29732);
and UO_2867 (O_2867,N_28534,N_29740);
nand UO_2868 (O_2868,N_29128,N_28596);
xnor UO_2869 (O_2869,N_29089,N_29535);
or UO_2870 (O_2870,N_29116,N_28951);
xor UO_2871 (O_2871,N_28800,N_28884);
xnor UO_2872 (O_2872,N_29757,N_28675);
xnor UO_2873 (O_2873,N_29219,N_29547);
or UO_2874 (O_2874,N_28741,N_28692);
xnor UO_2875 (O_2875,N_28777,N_28657);
nor UO_2876 (O_2876,N_29027,N_29702);
and UO_2877 (O_2877,N_29391,N_29452);
and UO_2878 (O_2878,N_29308,N_29266);
and UO_2879 (O_2879,N_29355,N_29695);
and UO_2880 (O_2880,N_29679,N_29598);
nor UO_2881 (O_2881,N_29862,N_29907);
or UO_2882 (O_2882,N_29973,N_29683);
and UO_2883 (O_2883,N_29138,N_29147);
xnor UO_2884 (O_2884,N_28895,N_28792);
nand UO_2885 (O_2885,N_29071,N_29473);
xor UO_2886 (O_2886,N_29195,N_28969);
nand UO_2887 (O_2887,N_29439,N_28809);
nor UO_2888 (O_2888,N_29929,N_29407);
nor UO_2889 (O_2889,N_28919,N_29844);
nand UO_2890 (O_2890,N_28755,N_29748);
or UO_2891 (O_2891,N_29517,N_28976);
and UO_2892 (O_2892,N_29196,N_29563);
and UO_2893 (O_2893,N_29893,N_29155);
and UO_2894 (O_2894,N_29653,N_28971);
nand UO_2895 (O_2895,N_29093,N_29498);
nand UO_2896 (O_2896,N_29238,N_28773);
and UO_2897 (O_2897,N_29106,N_29945);
nand UO_2898 (O_2898,N_28701,N_28730);
and UO_2899 (O_2899,N_29089,N_29403);
and UO_2900 (O_2900,N_28602,N_29097);
or UO_2901 (O_2901,N_29715,N_29974);
or UO_2902 (O_2902,N_29465,N_28628);
xor UO_2903 (O_2903,N_29958,N_28674);
or UO_2904 (O_2904,N_29140,N_28940);
and UO_2905 (O_2905,N_29201,N_28938);
or UO_2906 (O_2906,N_29591,N_28583);
or UO_2907 (O_2907,N_29337,N_29990);
nand UO_2908 (O_2908,N_29454,N_29896);
and UO_2909 (O_2909,N_29581,N_28777);
nor UO_2910 (O_2910,N_28582,N_29787);
or UO_2911 (O_2911,N_29311,N_29485);
nand UO_2912 (O_2912,N_29685,N_29336);
nor UO_2913 (O_2913,N_29669,N_29409);
nand UO_2914 (O_2914,N_29891,N_29403);
xnor UO_2915 (O_2915,N_29465,N_29193);
nor UO_2916 (O_2916,N_28747,N_29030);
and UO_2917 (O_2917,N_29368,N_29573);
or UO_2918 (O_2918,N_28914,N_28901);
nor UO_2919 (O_2919,N_29896,N_28717);
and UO_2920 (O_2920,N_28804,N_29392);
nand UO_2921 (O_2921,N_29488,N_28680);
nor UO_2922 (O_2922,N_28633,N_29401);
and UO_2923 (O_2923,N_28538,N_29850);
or UO_2924 (O_2924,N_29984,N_28827);
nand UO_2925 (O_2925,N_29267,N_29581);
xnor UO_2926 (O_2926,N_28898,N_29737);
xor UO_2927 (O_2927,N_28797,N_29280);
nand UO_2928 (O_2928,N_29181,N_29420);
xnor UO_2929 (O_2929,N_28933,N_29422);
nand UO_2930 (O_2930,N_29963,N_28938);
or UO_2931 (O_2931,N_29948,N_28541);
nor UO_2932 (O_2932,N_29551,N_28811);
nor UO_2933 (O_2933,N_28807,N_28518);
or UO_2934 (O_2934,N_29012,N_28534);
xor UO_2935 (O_2935,N_28798,N_28687);
xor UO_2936 (O_2936,N_29336,N_29097);
xor UO_2937 (O_2937,N_28524,N_29521);
xor UO_2938 (O_2938,N_29402,N_29870);
xnor UO_2939 (O_2939,N_28552,N_29530);
nand UO_2940 (O_2940,N_28961,N_29079);
nand UO_2941 (O_2941,N_29770,N_29542);
and UO_2942 (O_2942,N_29126,N_28669);
and UO_2943 (O_2943,N_29006,N_29622);
and UO_2944 (O_2944,N_29576,N_28749);
xnor UO_2945 (O_2945,N_28537,N_28785);
or UO_2946 (O_2946,N_29838,N_29550);
nand UO_2947 (O_2947,N_29114,N_28953);
xor UO_2948 (O_2948,N_29292,N_28771);
xor UO_2949 (O_2949,N_29592,N_29591);
or UO_2950 (O_2950,N_29332,N_29140);
or UO_2951 (O_2951,N_29025,N_29037);
xor UO_2952 (O_2952,N_29828,N_29324);
or UO_2953 (O_2953,N_28518,N_28848);
and UO_2954 (O_2954,N_29852,N_29515);
or UO_2955 (O_2955,N_28675,N_29997);
xnor UO_2956 (O_2956,N_29291,N_29351);
nand UO_2957 (O_2957,N_29589,N_28676);
or UO_2958 (O_2958,N_29946,N_28685);
xor UO_2959 (O_2959,N_29137,N_28855);
nand UO_2960 (O_2960,N_28670,N_29324);
xor UO_2961 (O_2961,N_28836,N_28642);
or UO_2962 (O_2962,N_28818,N_28778);
xor UO_2963 (O_2963,N_29208,N_29473);
nand UO_2964 (O_2964,N_29055,N_29519);
xnor UO_2965 (O_2965,N_29421,N_29269);
and UO_2966 (O_2966,N_29530,N_29152);
or UO_2967 (O_2967,N_29393,N_29047);
or UO_2968 (O_2968,N_29402,N_29321);
nand UO_2969 (O_2969,N_28654,N_29136);
nand UO_2970 (O_2970,N_28760,N_28557);
nor UO_2971 (O_2971,N_28965,N_29487);
or UO_2972 (O_2972,N_28635,N_29108);
and UO_2973 (O_2973,N_29190,N_29777);
or UO_2974 (O_2974,N_28892,N_29188);
or UO_2975 (O_2975,N_29942,N_29425);
nor UO_2976 (O_2976,N_28713,N_29652);
or UO_2977 (O_2977,N_29343,N_29783);
xnor UO_2978 (O_2978,N_29655,N_28766);
and UO_2979 (O_2979,N_29930,N_29640);
xnor UO_2980 (O_2980,N_29237,N_28660);
and UO_2981 (O_2981,N_29233,N_29547);
or UO_2982 (O_2982,N_29599,N_28942);
nor UO_2983 (O_2983,N_28851,N_28759);
nor UO_2984 (O_2984,N_29044,N_29991);
and UO_2985 (O_2985,N_29956,N_29783);
and UO_2986 (O_2986,N_29316,N_29577);
or UO_2987 (O_2987,N_29216,N_29861);
nor UO_2988 (O_2988,N_29018,N_28953);
or UO_2989 (O_2989,N_29792,N_29286);
nand UO_2990 (O_2990,N_28976,N_29993);
nand UO_2991 (O_2991,N_29866,N_29260);
nor UO_2992 (O_2992,N_28611,N_29226);
or UO_2993 (O_2993,N_29394,N_28790);
xor UO_2994 (O_2994,N_28680,N_29341);
nand UO_2995 (O_2995,N_29016,N_29191);
or UO_2996 (O_2996,N_28502,N_29141);
nand UO_2997 (O_2997,N_29868,N_29562);
xor UO_2998 (O_2998,N_29625,N_28958);
xor UO_2999 (O_2999,N_28633,N_29913);
xnor UO_3000 (O_3000,N_29801,N_29447);
and UO_3001 (O_3001,N_28551,N_29030);
and UO_3002 (O_3002,N_29575,N_29770);
xnor UO_3003 (O_3003,N_28690,N_29722);
and UO_3004 (O_3004,N_29244,N_29693);
xor UO_3005 (O_3005,N_28928,N_28729);
nor UO_3006 (O_3006,N_29886,N_28544);
xnor UO_3007 (O_3007,N_28726,N_29110);
nand UO_3008 (O_3008,N_29965,N_28538);
nand UO_3009 (O_3009,N_29751,N_29142);
and UO_3010 (O_3010,N_28871,N_28827);
nor UO_3011 (O_3011,N_29619,N_28627);
nand UO_3012 (O_3012,N_29121,N_29962);
and UO_3013 (O_3013,N_29835,N_28943);
xor UO_3014 (O_3014,N_28674,N_28647);
xnor UO_3015 (O_3015,N_29026,N_29364);
nand UO_3016 (O_3016,N_29046,N_29548);
xor UO_3017 (O_3017,N_29791,N_28517);
nor UO_3018 (O_3018,N_29773,N_29686);
nand UO_3019 (O_3019,N_29224,N_28612);
nand UO_3020 (O_3020,N_28749,N_28976);
or UO_3021 (O_3021,N_28879,N_29943);
xnor UO_3022 (O_3022,N_29353,N_29611);
xor UO_3023 (O_3023,N_29591,N_29951);
or UO_3024 (O_3024,N_29979,N_28650);
nor UO_3025 (O_3025,N_28655,N_29885);
or UO_3026 (O_3026,N_29558,N_28793);
xor UO_3027 (O_3027,N_28784,N_28711);
nand UO_3028 (O_3028,N_29433,N_29477);
nor UO_3029 (O_3029,N_29196,N_28898);
xor UO_3030 (O_3030,N_29302,N_28713);
nand UO_3031 (O_3031,N_29615,N_28934);
or UO_3032 (O_3032,N_29496,N_29499);
and UO_3033 (O_3033,N_29452,N_29607);
xnor UO_3034 (O_3034,N_28896,N_29765);
nor UO_3035 (O_3035,N_29430,N_28594);
nor UO_3036 (O_3036,N_29726,N_29215);
nor UO_3037 (O_3037,N_29267,N_29483);
nand UO_3038 (O_3038,N_28608,N_29595);
xnor UO_3039 (O_3039,N_29588,N_29227);
and UO_3040 (O_3040,N_29194,N_28512);
xnor UO_3041 (O_3041,N_29454,N_28510);
and UO_3042 (O_3042,N_29807,N_28645);
nand UO_3043 (O_3043,N_29664,N_29246);
or UO_3044 (O_3044,N_29156,N_29759);
nor UO_3045 (O_3045,N_29185,N_29911);
or UO_3046 (O_3046,N_29162,N_28633);
or UO_3047 (O_3047,N_29808,N_28706);
and UO_3048 (O_3048,N_29723,N_29782);
nand UO_3049 (O_3049,N_29898,N_28851);
nand UO_3050 (O_3050,N_28760,N_29842);
and UO_3051 (O_3051,N_29500,N_28987);
nand UO_3052 (O_3052,N_28703,N_29821);
nand UO_3053 (O_3053,N_29736,N_29021);
nor UO_3054 (O_3054,N_28847,N_28729);
and UO_3055 (O_3055,N_28877,N_28926);
nand UO_3056 (O_3056,N_29940,N_28733);
xor UO_3057 (O_3057,N_28945,N_29251);
nand UO_3058 (O_3058,N_29127,N_29536);
xor UO_3059 (O_3059,N_29907,N_29650);
nor UO_3060 (O_3060,N_28938,N_29940);
and UO_3061 (O_3061,N_29979,N_28713);
xnor UO_3062 (O_3062,N_28562,N_29035);
xnor UO_3063 (O_3063,N_29895,N_28679);
or UO_3064 (O_3064,N_29678,N_29944);
xor UO_3065 (O_3065,N_28603,N_29540);
nor UO_3066 (O_3066,N_29890,N_28537);
nand UO_3067 (O_3067,N_29987,N_29037);
or UO_3068 (O_3068,N_29073,N_28934);
and UO_3069 (O_3069,N_28529,N_28612);
nor UO_3070 (O_3070,N_28759,N_29207);
nand UO_3071 (O_3071,N_28813,N_28500);
nor UO_3072 (O_3072,N_29495,N_28519);
nor UO_3073 (O_3073,N_29064,N_28635);
nand UO_3074 (O_3074,N_28787,N_28521);
or UO_3075 (O_3075,N_28943,N_29155);
nor UO_3076 (O_3076,N_29572,N_28901);
or UO_3077 (O_3077,N_29616,N_29546);
nor UO_3078 (O_3078,N_29719,N_29475);
xnor UO_3079 (O_3079,N_29031,N_29991);
nor UO_3080 (O_3080,N_29025,N_28815);
nand UO_3081 (O_3081,N_29416,N_29154);
nor UO_3082 (O_3082,N_29481,N_29947);
nand UO_3083 (O_3083,N_29526,N_29050);
nand UO_3084 (O_3084,N_28807,N_29343);
or UO_3085 (O_3085,N_28666,N_29797);
nor UO_3086 (O_3086,N_29311,N_29209);
nor UO_3087 (O_3087,N_29657,N_28598);
nand UO_3088 (O_3088,N_28632,N_29210);
or UO_3089 (O_3089,N_29899,N_29189);
nor UO_3090 (O_3090,N_29248,N_29858);
nor UO_3091 (O_3091,N_28877,N_29556);
nor UO_3092 (O_3092,N_29865,N_29273);
and UO_3093 (O_3093,N_29053,N_28859);
nand UO_3094 (O_3094,N_28968,N_29370);
or UO_3095 (O_3095,N_28847,N_29518);
nor UO_3096 (O_3096,N_29255,N_28684);
nand UO_3097 (O_3097,N_29984,N_29172);
and UO_3098 (O_3098,N_28828,N_29991);
or UO_3099 (O_3099,N_29241,N_28621);
nor UO_3100 (O_3100,N_28562,N_29920);
or UO_3101 (O_3101,N_29742,N_29979);
nor UO_3102 (O_3102,N_29255,N_28833);
or UO_3103 (O_3103,N_29356,N_29551);
and UO_3104 (O_3104,N_29481,N_28728);
or UO_3105 (O_3105,N_28647,N_29591);
nand UO_3106 (O_3106,N_29436,N_29503);
nand UO_3107 (O_3107,N_29587,N_28529);
nand UO_3108 (O_3108,N_28534,N_29753);
xnor UO_3109 (O_3109,N_28604,N_29267);
nand UO_3110 (O_3110,N_29633,N_29443);
nor UO_3111 (O_3111,N_29824,N_28798);
and UO_3112 (O_3112,N_28973,N_28719);
or UO_3113 (O_3113,N_29799,N_29920);
nor UO_3114 (O_3114,N_28887,N_29223);
xor UO_3115 (O_3115,N_29585,N_28779);
xor UO_3116 (O_3116,N_28695,N_29188);
nor UO_3117 (O_3117,N_29505,N_28554);
xnor UO_3118 (O_3118,N_29663,N_28850);
nor UO_3119 (O_3119,N_29385,N_29231);
or UO_3120 (O_3120,N_29580,N_29794);
xnor UO_3121 (O_3121,N_29388,N_28734);
or UO_3122 (O_3122,N_29305,N_28548);
nor UO_3123 (O_3123,N_29568,N_29718);
or UO_3124 (O_3124,N_28749,N_28967);
nor UO_3125 (O_3125,N_29094,N_29244);
or UO_3126 (O_3126,N_29352,N_28644);
nand UO_3127 (O_3127,N_28979,N_29500);
nor UO_3128 (O_3128,N_29075,N_29863);
and UO_3129 (O_3129,N_29143,N_29345);
xor UO_3130 (O_3130,N_29528,N_29904);
and UO_3131 (O_3131,N_29838,N_28859);
nor UO_3132 (O_3132,N_28593,N_29837);
or UO_3133 (O_3133,N_29689,N_28889);
or UO_3134 (O_3134,N_29497,N_28777);
or UO_3135 (O_3135,N_29939,N_29712);
xnor UO_3136 (O_3136,N_29425,N_29302);
xor UO_3137 (O_3137,N_29799,N_28901);
xor UO_3138 (O_3138,N_29635,N_29736);
nand UO_3139 (O_3139,N_29484,N_29022);
xor UO_3140 (O_3140,N_28745,N_29320);
and UO_3141 (O_3141,N_28645,N_29225);
nand UO_3142 (O_3142,N_29952,N_29587);
or UO_3143 (O_3143,N_28888,N_29739);
nand UO_3144 (O_3144,N_28856,N_29466);
xor UO_3145 (O_3145,N_28765,N_29040);
or UO_3146 (O_3146,N_29546,N_28776);
nor UO_3147 (O_3147,N_28639,N_28627);
nor UO_3148 (O_3148,N_28993,N_29415);
xnor UO_3149 (O_3149,N_29257,N_29497);
or UO_3150 (O_3150,N_29717,N_29714);
nor UO_3151 (O_3151,N_28695,N_29630);
nand UO_3152 (O_3152,N_29284,N_29764);
or UO_3153 (O_3153,N_29764,N_29651);
or UO_3154 (O_3154,N_28635,N_29958);
and UO_3155 (O_3155,N_29717,N_28939);
nand UO_3156 (O_3156,N_29840,N_29437);
nand UO_3157 (O_3157,N_29322,N_29832);
or UO_3158 (O_3158,N_28594,N_29185);
nand UO_3159 (O_3159,N_29632,N_28784);
or UO_3160 (O_3160,N_29955,N_29765);
nand UO_3161 (O_3161,N_29168,N_29736);
nor UO_3162 (O_3162,N_29048,N_28780);
nand UO_3163 (O_3163,N_29268,N_28882);
nor UO_3164 (O_3164,N_29320,N_28767);
xnor UO_3165 (O_3165,N_28692,N_29276);
xnor UO_3166 (O_3166,N_29993,N_29940);
and UO_3167 (O_3167,N_29508,N_28797);
and UO_3168 (O_3168,N_28555,N_29698);
and UO_3169 (O_3169,N_28928,N_28945);
nand UO_3170 (O_3170,N_28882,N_29676);
nor UO_3171 (O_3171,N_28701,N_29548);
and UO_3172 (O_3172,N_29923,N_28516);
or UO_3173 (O_3173,N_29542,N_28520);
xnor UO_3174 (O_3174,N_28651,N_28659);
and UO_3175 (O_3175,N_28837,N_29394);
nand UO_3176 (O_3176,N_29613,N_28720);
xnor UO_3177 (O_3177,N_29224,N_29727);
nor UO_3178 (O_3178,N_29508,N_29399);
xor UO_3179 (O_3179,N_29416,N_29112);
and UO_3180 (O_3180,N_29340,N_28800);
and UO_3181 (O_3181,N_28717,N_29674);
or UO_3182 (O_3182,N_29703,N_28540);
and UO_3183 (O_3183,N_29325,N_29092);
nor UO_3184 (O_3184,N_28603,N_29569);
or UO_3185 (O_3185,N_28744,N_29180);
nor UO_3186 (O_3186,N_28917,N_29565);
nand UO_3187 (O_3187,N_28575,N_29471);
nor UO_3188 (O_3188,N_28589,N_28585);
or UO_3189 (O_3189,N_28643,N_29444);
xor UO_3190 (O_3190,N_29374,N_29115);
nand UO_3191 (O_3191,N_28819,N_29787);
or UO_3192 (O_3192,N_28874,N_29634);
or UO_3193 (O_3193,N_28536,N_28647);
nand UO_3194 (O_3194,N_28873,N_29638);
or UO_3195 (O_3195,N_28788,N_29762);
nor UO_3196 (O_3196,N_28633,N_29243);
xor UO_3197 (O_3197,N_28998,N_29272);
nand UO_3198 (O_3198,N_29783,N_28918);
xor UO_3199 (O_3199,N_29614,N_29325);
nand UO_3200 (O_3200,N_29685,N_29786);
xnor UO_3201 (O_3201,N_29816,N_29564);
or UO_3202 (O_3202,N_29205,N_28727);
xnor UO_3203 (O_3203,N_29432,N_29338);
or UO_3204 (O_3204,N_29170,N_29664);
nor UO_3205 (O_3205,N_29342,N_28665);
nand UO_3206 (O_3206,N_29712,N_29668);
nor UO_3207 (O_3207,N_29594,N_29084);
nand UO_3208 (O_3208,N_29349,N_29917);
or UO_3209 (O_3209,N_29252,N_29094);
nand UO_3210 (O_3210,N_29056,N_28750);
nor UO_3211 (O_3211,N_29716,N_29763);
and UO_3212 (O_3212,N_28615,N_29265);
and UO_3213 (O_3213,N_29742,N_29876);
nor UO_3214 (O_3214,N_29010,N_29924);
and UO_3215 (O_3215,N_28992,N_29621);
and UO_3216 (O_3216,N_29809,N_28693);
and UO_3217 (O_3217,N_29319,N_29479);
and UO_3218 (O_3218,N_28871,N_28522);
nand UO_3219 (O_3219,N_28686,N_29287);
and UO_3220 (O_3220,N_28983,N_28596);
nor UO_3221 (O_3221,N_29951,N_28721);
or UO_3222 (O_3222,N_29347,N_29814);
and UO_3223 (O_3223,N_29169,N_29724);
nor UO_3224 (O_3224,N_29305,N_28967);
nand UO_3225 (O_3225,N_29435,N_29053);
or UO_3226 (O_3226,N_29727,N_29288);
xor UO_3227 (O_3227,N_29020,N_28523);
nor UO_3228 (O_3228,N_29094,N_29205);
or UO_3229 (O_3229,N_28799,N_28733);
and UO_3230 (O_3230,N_28793,N_29113);
or UO_3231 (O_3231,N_29291,N_29663);
nor UO_3232 (O_3232,N_29848,N_28879);
and UO_3233 (O_3233,N_28593,N_29499);
and UO_3234 (O_3234,N_29596,N_28975);
nor UO_3235 (O_3235,N_29967,N_29655);
nand UO_3236 (O_3236,N_28892,N_28907);
xnor UO_3237 (O_3237,N_29577,N_28679);
or UO_3238 (O_3238,N_28503,N_29060);
or UO_3239 (O_3239,N_28999,N_29039);
and UO_3240 (O_3240,N_29975,N_29226);
or UO_3241 (O_3241,N_29726,N_29463);
or UO_3242 (O_3242,N_29446,N_29907);
nand UO_3243 (O_3243,N_29491,N_29852);
xnor UO_3244 (O_3244,N_29721,N_29103);
or UO_3245 (O_3245,N_29698,N_29237);
xnor UO_3246 (O_3246,N_29880,N_29742);
nand UO_3247 (O_3247,N_29192,N_29725);
and UO_3248 (O_3248,N_29761,N_28772);
nand UO_3249 (O_3249,N_28781,N_28945);
nand UO_3250 (O_3250,N_29100,N_29668);
nor UO_3251 (O_3251,N_29795,N_28521);
xnor UO_3252 (O_3252,N_29340,N_29240);
nand UO_3253 (O_3253,N_28757,N_29473);
and UO_3254 (O_3254,N_28501,N_28634);
xnor UO_3255 (O_3255,N_29897,N_28808);
or UO_3256 (O_3256,N_29464,N_29453);
nor UO_3257 (O_3257,N_29067,N_29454);
xnor UO_3258 (O_3258,N_28912,N_28776);
nand UO_3259 (O_3259,N_29205,N_29634);
and UO_3260 (O_3260,N_29360,N_29257);
and UO_3261 (O_3261,N_29554,N_29313);
and UO_3262 (O_3262,N_29749,N_29067);
and UO_3263 (O_3263,N_28559,N_29383);
xnor UO_3264 (O_3264,N_29136,N_29209);
nand UO_3265 (O_3265,N_29485,N_29770);
or UO_3266 (O_3266,N_28886,N_29456);
xnor UO_3267 (O_3267,N_29317,N_29454);
nand UO_3268 (O_3268,N_29513,N_29277);
and UO_3269 (O_3269,N_29658,N_28926);
xor UO_3270 (O_3270,N_28735,N_29072);
and UO_3271 (O_3271,N_29463,N_29954);
nor UO_3272 (O_3272,N_29624,N_28722);
xor UO_3273 (O_3273,N_29180,N_29566);
xor UO_3274 (O_3274,N_29327,N_29924);
or UO_3275 (O_3275,N_29468,N_29930);
nor UO_3276 (O_3276,N_29684,N_28810);
or UO_3277 (O_3277,N_29442,N_29364);
nand UO_3278 (O_3278,N_29252,N_28781);
and UO_3279 (O_3279,N_29377,N_28580);
xnor UO_3280 (O_3280,N_28514,N_29665);
and UO_3281 (O_3281,N_29724,N_29964);
and UO_3282 (O_3282,N_29120,N_29532);
xnor UO_3283 (O_3283,N_28788,N_29418);
xnor UO_3284 (O_3284,N_29637,N_29358);
nor UO_3285 (O_3285,N_29100,N_29960);
xnor UO_3286 (O_3286,N_29744,N_28590);
xnor UO_3287 (O_3287,N_28583,N_29474);
or UO_3288 (O_3288,N_28997,N_29298);
and UO_3289 (O_3289,N_29855,N_29713);
nor UO_3290 (O_3290,N_29961,N_29657);
or UO_3291 (O_3291,N_28906,N_28510);
xor UO_3292 (O_3292,N_29974,N_28743);
and UO_3293 (O_3293,N_28862,N_29369);
and UO_3294 (O_3294,N_28808,N_28851);
and UO_3295 (O_3295,N_29316,N_29202);
and UO_3296 (O_3296,N_29913,N_28789);
xor UO_3297 (O_3297,N_29124,N_29453);
xnor UO_3298 (O_3298,N_29884,N_28703);
nor UO_3299 (O_3299,N_28805,N_28657);
nor UO_3300 (O_3300,N_29180,N_29446);
nor UO_3301 (O_3301,N_28552,N_28627);
xor UO_3302 (O_3302,N_29623,N_28579);
nand UO_3303 (O_3303,N_29881,N_29197);
and UO_3304 (O_3304,N_28952,N_28763);
xor UO_3305 (O_3305,N_29357,N_28782);
xor UO_3306 (O_3306,N_29793,N_28783);
and UO_3307 (O_3307,N_29471,N_29698);
and UO_3308 (O_3308,N_29215,N_29723);
xor UO_3309 (O_3309,N_29472,N_29677);
or UO_3310 (O_3310,N_29240,N_29487);
or UO_3311 (O_3311,N_29336,N_29043);
or UO_3312 (O_3312,N_29417,N_29727);
or UO_3313 (O_3313,N_29949,N_29570);
nor UO_3314 (O_3314,N_28929,N_28559);
nor UO_3315 (O_3315,N_28540,N_28885);
nand UO_3316 (O_3316,N_29863,N_28886);
and UO_3317 (O_3317,N_28777,N_29080);
xnor UO_3318 (O_3318,N_29404,N_29564);
xnor UO_3319 (O_3319,N_29576,N_29658);
nand UO_3320 (O_3320,N_29735,N_28944);
nor UO_3321 (O_3321,N_28847,N_29212);
or UO_3322 (O_3322,N_29408,N_28625);
and UO_3323 (O_3323,N_29568,N_28683);
nor UO_3324 (O_3324,N_29257,N_29158);
or UO_3325 (O_3325,N_28942,N_28784);
or UO_3326 (O_3326,N_29685,N_29723);
nand UO_3327 (O_3327,N_29906,N_28586);
xor UO_3328 (O_3328,N_29423,N_29695);
xnor UO_3329 (O_3329,N_28636,N_29394);
or UO_3330 (O_3330,N_28516,N_29335);
or UO_3331 (O_3331,N_28942,N_28529);
nand UO_3332 (O_3332,N_29080,N_28853);
xor UO_3333 (O_3333,N_29471,N_29621);
or UO_3334 (O_3334,N_29124,N_29877);
nand UO_3335 (O_3335,N_28935,N_28581);
or UO_3336 (O_3336,N_28923,N_28873);
nand UO_3337 (O_3337,N_29207,N_28569);
and UO_3338 (O_3338,N_28719,N_28900);
or UO_3339 (O_3339,N_29480,N_29574);
nand UO_3340 (O_3340,N_28798,N_29906);
and UO_3341 (O_3341,N_28523,N_29353);
or UO_3342 (O_3342,N_29359,N_29747);
or UO_3343 (O_3343,N_29574,N_29068);
or UO_3344 (O_3344,N_28727,N_29044);
nor UO_3345 (O_3345,N_29701,N_29725);
nor UO_3346 (O_3346,N_29234,N_29745);
nor UO_3347 (O_3347,N_29133,N_28915);
or UO_3348 (O_3348,N_28778,N_29142);
nand UO_3349 (O_3349,N_29795,N_29818);
xnor UO_3350 (O_3350,N_28518,N_29655);
xnor UO_3351 (O_3351,N_29915,N_29354);
nor UO_3352 (O_3352,N_28842,N_29301);
xnor UO_3353 (O_3353,N_29304,N_29666);
xor UO_3354 (O_3354,N_29514,N_29137);
and UO_3355 (O_3355,N_28759,N_29494);
xnor UO_3356 (O_3356,N_29507,N_28982);
or UO_3357 (O_3357,N_29099,N_28898);
nor UO_3358 (O_3358,N_29569,N_29566);
and UO_3359 (O_3359,N_29162,N_29336);
xnor UO_3360 (O_3360,N_29796,N_28932);
or UO_3361 (O_3361,N_29513,N_28967);
nand UO_3362 (O_3362,N_29456,N_29395);
nor UO_3363 (O_3363,N_29658,N_28946);
xnor UO_3364 (O_3364,N_29434,N_29253);
nor UO_3365 (O_3365,N_29198,N_28780);
nand UO_3366 (O_3366,N_28869,N_28702);
nand UO_3367 (O_3367,N_29468,N_29633);
or UO_3368 (O_3368,N_29112,N_29716);
nor UO_3369 (O_3369,N_29820,N_28741);
nand UO_3370 (O_3370,N_29478,N_28878);
xor UO_3371 (O_3371,N_29406,N_29962);
nor UO_3372 (O_3372,N_29195,N_29490);
nand UO_3373 (O_3373,N_29001,N_29628);
xor UO_3374 (O_3374,N_28849,N_29134);
xor UO_3375 (O_3375,N_28513,N_28584);
xnor UO_3376 (O_3376,N_29669,N_29737);
nor UO_3377 (O_3377,N_29440,N_28598);
xnor UO_3378 (O_3378,N_28520,N_29146);
nor UO_3379 (O_3379,N_29236,N_29743);
nand UO_3380 (O_3380,N_29679,N_29606);
or UO_3381 (O_3381,N_29167,N_29961);
nand UO_3382 (O_3382,N_28874,N_28752);
and UO_3383 (O_3383,N_28759,N_28845);
nand UO_3384 (O_3384,N_28600,N_28693);
or UO_3385 (O_3385,N_28782,N_28786);
nor UO_3386 (O_3386,N_28569,N_29074);
or UO_3387 (O_3387,N_29219,N_29016);
or UO_3388 (O_3388,N_29386,N_28609);
nor UO_3389 (O_3389,N_29509,N_29151);
nand UO_3390 (O_3390,N_28809,N_29914);
nor UO_3391 (O_3391,N_29318,N_29867);
nor UO_3392 (O_3392,N_29154,N_29830);
nor UO_3393 (O_3393,N_29619,N_28995);
nor UO_3394 (O_3394,N_29474,N_28525);
nor UO_3395 (O_3395,N_29499,N_29468);
nand UO_3396 (O_3396,N_29958,N_29381);
nand UO_3397 (O_3397,N_28521,N_28522);
xnor UO_3398 (O_3398,N_28886,N_29732);
xor UO_3399 (O_3399,N_29172,N_28778);
nor UO_3400 (O_3400,N_29660,N_29744);
and UO_3401 (O_3401,N_29005,N_28882);
xor UO_3402 (O_3402,N_28926,N_29238);
nor UO_3403 (O_3403,N_29237,N_29063);
xor UO_3404 (O_3404,N_28910,N_29666);
and UO_3405 (O_3405,N_29923,N_28961);
nor UO_3406 (O_3406,N_28955,N_28869);
nand UO_3407 (O_3407,N_28707,N_28934);
and UO_3408 (O_3408,N_29909,N_29605);
nand UO_3409 (O_3409,N_28888,N_29584);
nor UO_3410 (O_3410,N_29382,N_29884);
xnor UO_3411 (O_3411,N_28503,N_28943);
or UO_3412 (O_3412,N_28935,N_29715);
or UO_3413 (O_3413,N_29311,N_28561);
nor UO_3414 (O_3414,N_28678,N_29043);
nor UO_3415 (O_3415,N_29468,N_29962);
nand UO_3416 (O_3416,N_29719,N_29325);
and UO_3417 (O_3417,N_28805,N_29773);
or UO_3418 (O_3418,N_29978,N_28598);
or UO_3419 (O_3419,N_29105,N_29860);
nand UO_3420 (O_3420,N_29801,N_28751);
nand UO_3421 (O_3421,N_29336,N_29173);
and UO_3422 (O_3422,N_29487,N_29135);
xnor UO_3423 (O_3423,N_29528,N_29552);
and UO_3424 (O_3424,N_29727,N_28945);
and UO_3425 (O_3425,N_29810,N_29631);
nor UO_3426 (O_3426,N_28602,N_28977);
and UO_3427 (O_3427,N_28569,N_29811);
nor UO_3428 (O_3428,N_29945,N_29012);
or UO_3429 (O_3429,N_28506,N_29350);
or UO_3430 (O_3430,N_29302,N_28615);
xnor UO_3431 (O_3431,N_28731,N_28555);
nor UO_3432 (O_3432,N_28516,N_28701);
xnor UO_3433 (O_3433,N_28661,N_28897);
nand UO_3434 (O_3434,N_28592,N_28723);
nor UO_3435 (O_3435,N_29934,N_28753);
nor UO_3436 (O_3436,N_28553,N_29026);
and UO_3437 (O_3437,N_29072,N_29818);
nand UO_3438 (O_3438,N_29147,N_29502);
nor UO_3439 (O_3439,N_29835,N_29803);
or UO_3440 (O_3440,N_28508,N_29146);
nor UO_3441 (O_3441,N_28726,N_29698);
nor UO_3442 (O_3442,N_29336,N_28736);
nor UO_3443 (O_3443,N_29274,N_29234);
or UO_3444 (O_3444,N_28763,N_29279);
xor UO_3445 (O_3445,N_28676,N_29470);
nand UO_3446 (O_3446,N_29094,N_28521);
and UO_3447 (O_3447,N_28851,N_28996);
and UO_3448 (O_3448,N_28573,N_29637);
xor UO_3449 (O_3449,N_29771,N_29793);
and UO_3450 (O_3450,N_28696,N_28858);
or UO_3451 (O_3451,N_28906,N_29057);
nor UO_3452 (O_3452,N_28803,N_29365);
nand UO_3453 (O_3453,N_29509,N_29199);
nand UO_3454 (O_3454,N_29758,N_28589);
nand UO_3455 (O_3455,N_29961,N_28952);
xnor UO_3456 (O_3456,N_28851,N_28593);
and UO_3457 (O_3457,N_28945,N_29988);
and UO_3458 (O_3458,N_29371,N_29198);
nor UO_3459 (O_3459,N_29809,N_29779);
xor UO_3460 (O_3460,N_29807,N_29760);
and UO_3461 (O_3461,N_28568,N_29165);
xor UO_3462 (O_3462,N_28882,N_29824);
xor UO_3463 (O_3463,N_28593,N_28949);
and UO_3464 (O_3464,N_29972,N_29748);
xnor UO_3465 (O_3465,N_28626,N_29041);
and UO_3466 (O_3466,N_29518,N_29876);
or UO_3467 (O_3467,N_29273,N_29847);
nand UO_3468 (O_3468,N_29675,N_29013);
nand UO_3469 (O_3469,N_29238,N_29912);
nand UO_3470 (O_3470,N_29746,N_28549);
xor UO_3471 (O_3471,N_29965,N_29280);
nor UO_3472 (O_3472,N_29698,N_29545);
xnor UO_3473 (O_3473,N_29456,N_28780);
and UO_3474 (O_3474,N_28832,N_28614);
xnor UO_3475 (O_3475,N_28756,N_29140);
and UO_3476 (O_3476,N_29159,N_29414);
nor UO_3477 (O_3477,N_29245,N_28592);
nor UO_3478 (O_3478,N_28560,N_29625);
nor UO_3479 (O_3479,N_29623,N_29827);
nand UO_3480 (O_3480,N_29178,N_28842);
and UO_3481 (O_3481,N_28995,N_29762);
and UO_3482 (O_3482,N_29076,N_29378);
and UO_3483 (O_3483,N_28620,N_29676);
xor UO_3484 (O_3484,N_28796,N_28533);
or UO_3485 (O_3485,N_28837,N_29774);
xnor UO_3486 (O_3486,N_28598,N_29019);
and UO_3487 (O_3487,N_29582,N_28895);
and UO_3488 (O_3488,N_29839,N_28724);
nand UO_3489 (O_3489,N_29141,N_28633);
or UO_3490 (O_3490,N_28769,N_28854);
or UO_3491 (O_3491,N_29177,N_29487);
xor UO_3492 (O_3492,N_29071,N_28839);
and UO_3493 (O_3493,N_28597,N_29848);
xnor UO_3494 (O_3494,N_29831,N_28806);
or UO_3495 (O_3495,N_28634,N_29538);
or UO_3496 (O_3496,N_28894,N_28910);
nand UO_3497 (O_3497,N_29461,N_29203);
or UO_3498 (O_3498,N_28546,N_28745);
and UO_3499 (O_3499,N_28557,N_28661);
endmodule