module basic_500_3000_500_4_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xnor U0 (N_0,In_156,In_451);
nor U1 (N_1,In_323,In_258);
nand U2 (N_2,In_340,In_267);
xor U3 (N_3,In_63,In_118);
nand U4 (N_4,In_10,In_394);
and U5 (N_5,In_275,In_273);
nand U6 (N_6,In_165,In_288);
nor U7 (N_7,In_274,In_265);
nor U8 (N_8,In_281,In_349);
or U9 (N_9,In_49,In_373);
nand U10 (N_10,In_271,In_370);
and U11 (N_11,In_22,In_270);
and U12 (N_12,In_160,In_131);
and U13 (N_13,In_364,In_97);
nor U14 (N_14,In_80,In_282);
nor U15 (N_15,In_99,In_426);
nand U16 (N_16,In_64,In_93);
or U17 (N_17,In_135,In_257);
and U18 (N_18,In_54,In_313);
and U19 (N_19,In_14,In_461);
nand U20 (N_20,In_89,In_293);
and U21 (N_21,In_72,In_185);
and U22 (N_22,In_286,In_92);
nor U23 (N_23,In_154,In_27);
nand U24 (N_24,In_48,In_177);
and U25 (N_25,In_37,In_170);
nor U26 (N_26,In_200,In_439);
nor U27 (N_27,In_161,In_29);
nor U28 (N_28,In_330,In_263);
nand U29 (N_29,In_175,In_212);
and U30 (N_30,In_479,In_476);
and U31 (N_31,In_58,In_489);
nor U32 (N_32,In_109,In_147);
or U33 (N_33,In_346,In_39);
nand U34 (N_34,In_42,In_291);
nand U35 (N_35,In_26,In_298);
nor U36 (N_36,In_254,In_40);
or U37 (N_37,In_457,In_17);
nor U38 (N_38,In_81,In_223);
nor U39 (N_39,In_18,In_126);
nor U40 (N_40,In_325,In_35);
and U41 (N_41,In_381,In_466);
nand U42 (N_42,In_380,In_382);
nand U43 (N_43,In_192,In_322);
or U44 (N_44,In_85,In_202);
or U45 (N_45,In_378,In_153);
and U46 (N_46,In_480,In_82);
xor U47 (N_47,In_152,In_83);
nor U48 (N_48,In_24,In_218);
or U49 (N_49,In_279,In_132);
and U50 (N_50,In_383,In_314);
or U51 (N_51,In_395,In_401);
and U52 (N_52,In_419,In_62);
nor U53 (N_53,In_342,In_148);
and U54 (N_54,In_403,In_32);
nor U55 (N_55,In_45,In_169);
or U56 (N_56,In_84,In_449);
nand U57 (N_57,In_320,In_71);
nand U58 (N_58,In_341,In_348);
and U59 (N_59,In_41,In_137);
or U60 (N_60,In_377,In_438);
or U61 (N_61,In_125,In_174);
nand U62 (N_62,In_262,In_53);
or U63 (N_63,In_484,In_43);
or U64 (N_64,In_283,In_151);
nand U65 (N_65,In_74,In_201);
or U66 (N_66,In_213,In_198);
nor U67 (N_67,In_297,In_87);
nand U68 (N_68,In_136,In_442);
xor U69 (N_69,In_197,In_240);
nand U70 (N_70,In_337,In_88);
nand U71 (N_71,In_114,In_123);
nor U72 (N_72,In_164,In_408);
nor U73 (N_73,In_65,In_232);
or U74 (N_74,In_235,In_344);
or U75 (N_75,In_352,In_79);
xor U76 (N_76,In_446,In_171);
nor U77 (N_77,In_482,In_145);
nor U78 (N_78,In_440,In_6);
or U79 (N_79,In_431,In_219);
nand U80 (N_80,In_491,In_425);
nor U81 (N_81,In_243,In_113);
nand U82 (N_82,In_241,In_221);
nand U83 (N_83,In_374,In_407);
and U84 (N_84,In_253,In_475);
and U85 (N_85,In_23,In_104);
or U86 (N_86,In_339,In_115);
xnor U87 (N_87,In_3,In_420);
xor U88 (N_88,In_412,In_168);
nand U89 (N_89,In_266,In_448);
or U90 (N_90,In_255,In_110);
and U91 (N_91,In_358,In_55);
nand U92 (N_92,In_259,In_434);
xnor U93 (N_93,In_304,In_230);
nor U94 (N_94,In_7,In_276);
nor U95 (N_95,In_214,In_28);
nor U96 (N_96,In_492,In_172);
and U97 (N_97,In_0,In_157);
and U98 (N_98,In_410,In_95);
and U99 (N_99,In_67,In_498);
nor U100 (N_100,In_415,In_238);
nor U101 (N_101,In_237,In_264);
nor U102 (N_102,In_445,In_309);
nor U103 (N_103,In_75,In_469);
nor U104 (N_104,In_31,In_496);
or U105 (N_105,In_470,In_376);
or U106 (N_106,In_56,In_452);
and U107 (N_107,In_331,In_73);
nand U108 (N_108,In_361,In_68);
nor U109 (N_109,In_351,In_363);
and U110 (N_110,In_312,In_494);
xor U111 (N_111,In_473,In_430);
nor U112 (N_112,In_371,In_308);
and U113 (N_113,In_398,In_261);
nand U114 (N_114,In_455,In_302);
nand U115 (N_115,In_216,In_453);
or U116 (N_116,In_411,In_359);
or U117 (N_117,In_182,In_188);
or U118 (N_118,In_44,In_248);
or U119 (N_119,In_269,In_196);
nand U120 (N_120,In_396,In_464);
and U121 (N_121,In_233,In_250);
or U122 (N_122,In_36,In_2);
nand U123 (N_123,In_159,In_60);
nor U124 (N_124,In_400,In_19);
nor U125 (N_125,In_173,In_292);
nor U126 (N_126,In_90,In_217);
nor U127 (N_127,In_33,In_404);
nand U128 (N_128,In_328,In_450);
or U129 (N_129,In_354,In_481);
nor U130 (N_130,In_335,In_163);
and U131 (N_131,In_301,In_38);
and U132 (N_132,In_76,In_140);
and U133 (N_133,In_416,In_167);
and U134 (N_134,In_290,In_247);
nand U135 (N_135,In_379,In_134);
nor U136 (N_136,In_497,In_278);
nand U137 (N_137,In_189,In_181);
or U138 (N_138,In_319,In_318);
xor U139 (N_139,In_471,In_487);
and U140 (N_140,In_386,In_366);
nor U141 (N_141,In_252,In_34);
nand U142 (N_142,In_428,In_144);
or U143 (N_143,In_389,In_332);
and U144 (N_144,In_338,In_205);
or U145 (N_145,In_311,In_204);
and U146 (N_146,In_143,In_409);
nand U147 (N_147,In_384,In_94);
xor U148 (N_148,In_108,In_317);
or U149 (N_149,In_133,In_46);
nor U150 (N_150,In_299,In_443);
or U151 (N_151,In_287,In_119);
or U152 (N_152,In_350,In_413);
or U153 (N_153,In_245,In_227);
or U154 (N_154,In_324,In_176);
or U155 (N_155,In_329,In_316);
nor U156 (N_156,In_120,In_493);
or U157 (N_157,In_210,In_333);
or U158 (N_158,In_208,In_405);
and U159 (N_159,In_249,In_495);
nand U160 (N_160,In_393,In_52);
nor U161 (N_161,In_392,In_96);
or U162 (N_162,In_9,In_146);
nor U163 (N_163,In_1,In_477);
and U164 (N_164,In_424,In_195);
and U165 (N_165,In_468,In_69);
nor U166 (N_166,In_142,In_234);
nor U167 (N_167,In_305,In_483);
and U168 (N_168,In_414,In_465);
nor U169 (N_169,In_390,In_485);
and U170 (N_170,In_4,In_321);
nand U171 (N_171,In_421,In_490);
nand U172 (N_172,In_180,In_51);
and U173 (N_173,In_260,In_315);
nand U174 (N_174,In_190,In_59);
nor U175 (N_175,In_231,In_436);
nand U176 (N_176,In_66,In_220);
or U177 (N_177,In_15,In_166);
nand U178 (N_178,In_459,In_300);
and U179 (N_179,In_207,In_327);
nand U180 (N_180,In_375,In_447);
nand U181 (N_181,In_467,In_357);
xnor U182 (N_182,In_139,In_25);
nand U183 (N_183,In_116,In_70);
and U184 (N_184,In_347,In_345);
nor U185 (N_185,In_86,In_178);
nor U186 (N_186,In_388,In_368);
nor U187 (N_187,In_365,In_343);
and U188 (N_188,In_122,In_130);
and U189 (N_189,In_402,In_57);
or U190 (N_190,In_391,In_423);
or U191 (N_191,In_179,In_360);
nor U192 (N_192,In_106,In_307);
or U193 (N_193,In_399,In_117);
nand U194 (N_194,In_211,In_226);
and U195 (N_195,In_454,In_499);
nand U196 (N_196,In_289,In_129);
nor U197 (N_197,In_303,In_474);
and U198 (N_198,In_100,In_246);
nand U199 (N_199,In_256,In_418);
nand U200 (N_200,In_107,In_272);
xor U201 (N_201,In_78,In_268);
and U202 (N_202,In_77,In_150);
nor U203 (N_203,In_155,In_203);
or U204 (N_204,In_215,In_224);
or U205 (N_205,In_225,In_367);
nand U206 (N_206,In_30,In_437);
xnor U207 (N_207,In_310,In_295);
or U208 (N_208,In_228,In_242);
or U209 (N_209,In_429,In_284);
or U210 (N_210,In_353,In_91);
or U211 (N_211,In_191,In_372);
nor U212 (N_212,In_326,In_277);
xor U213 (N_213,In_20,In_138);
nor U214 (N_214,In_5,In_103);
or U215 (N_215,In_362,In_334);
xnor U216 (N_216,In_193,In_432);
or U217 (N_217,In_13,In_162);
or U218 (N_218,In_183,In_111);
nand U219 (N_219,In_458,In_422);
xor U220 (N_220,In_184,In_385);
nor U221 (N_221,In_488,In_462);
nand U222 (N_222,In_11,In_98);
and U223 (N_223,In_199,In_8);
nand U224 (N_224,In_444,In_236);
or U225 (N_225,In_194,In_355);
and U226 (N_226,In_406,In_187);
xor U227 (N_227,In_61,In_433);
nand U228 (N_228,In_460,In_463);
nand U229 (N_229,In_435,In_369);
nand U230 (N_230,In_47,In_105);
nand U231 (N_231,In_206,In_124);
and U232 (N_232,In_456,In_141);
xnor U233 (N_233,In_222,In_280);
and U234 (N_234,In_128,In_417);
and U235 (N_235,In_397,In_336);
nor U236 (N_236,In_21,In_441);
nand U237 (N_237,In_229,In_12);
or U238 (N_238,In_486,In_251);
nor U239 (N_239,In_209,In_427);
or U240 (N_240,In_244,In_387);
and U241 (N_241,In_16,In_478);
xor U242 (N_242,In_356,In_239);
or U243 (N_243,In_285,In_102);
nor U244 (N_244,In_127,In_121);
or U245 (N_245,In_294,In_101);
and U246 (N_246,In_112,In_149);
nor U247 (N_247,In_158,In_186);
nand U248 (N_248,In_472,In_306);
nand U249 (N_249,In_296,In_50);
nor U250 (N_250,In_208,In_387);
nor U251 (N_251,In_36,In_185);
nor U252 (N_252,In_5,In_259);
nor U253 (N_253,In_231,In_179);
and U254 (N_254,In_354,In_401);
nand U255 (N_255,In_121,In_242);
and U256 (N_256,In_205,In_26);
or U257 (N_257,In_134,In_36);
nor U258 (N_258,In_116,In_94);
nor U259 (N_259,In_172,In_399);
or U260 (N_260,In_415,In_139);
nor U261 (N_261,In_383,In_451);
nand U262 (N_262,In_391,In_473);
or U263 (N_263,In_415,In_79);
and U264 (N_264,In_277,In_268);
nor U265 (N_265,In_238,In_167);
and U266 (N_266,In_323,In_352);
xnor U267 (N_267,In_174,In_124);
or U268 (N_268,In_250,In_432);
nand U269 (N_269,In_52,In_288);
or U270 (N_270,In_307,In_158);
or U271 (N_271,In_468,In_381);
or U272 (N_272,In_189,In_397);
and U273 (N_273,In_47,In_491);
and U274 (N_274,In_369,In_302);
nor U275 (N_275,In_326,In_350);
nand U276 (N_276,In_465,In_454);
or U277 (N_277,In_398,In_164);
nand U278 (N_278,In_432,In_426);
and U279 (N_279,In_239,In_248);
nand U280 (N_280,In_68,In_322);
nand U281 (N_281,In_2,In_432);
nand U282 (N_282,In_463,In_223);
xnor U283 (N_283,In_18,In_405);
or U284 (N_284,In_472,In_13);
or U285 (N_285,In_229,In_175);
or U286 (N_286,In_442,In_231);
or U287 (N_287,In_499,In_253);
nand U288 (N_288,In_37,In_446);
nand U289 (N_289,In_30,In_495);
xor U290 (N_290,In_205,In_299);
xor U291 (N_291,In_258,In_279);
nor U292 (N_292,In_343,In_479);
nor U293 (N_293,In_290,In_426);
nor U294 (N_294,In_101,In_158);
nand U295 (N_295,In_62,In_25);
xnor U296 (N_296,In_488,In_402);
or U297 (N_297,In_7,In_161);
nand U298 (N_298,In_384,In_46);
nor U299 (N_299,In_111,In_205);
or U300 (N_300,In_147,In_359);
nand U301 (N_301,In_262,In_401);
and U302 (N_302,In_30,In_380);
or U303 (N_303,In_65,In_44);
nor U304 (N_304,In_199,In_253);
xnor U305 (N_305,In_495,In_466);
or U306 (N_306,In_365,In_191);
and U307 (N_307,In_434,In_356);
nor U308 (N_308,In_374,In_359);
and U309 (N_309,In_387,In_95);
nand U310 (N_310,In_388,In_304);
and U311 (N_311,In_341,In_319);
or U312 (N_312,In_67,In_74);
xnor U313 (N_313,In_175,In_272);
nand U314 (N_314,In_289,In_317);
xnor U315 (N_315,In_477,In_180);
and U316 (N_316,In_257,In_164);
nor U317 (N_317,In_99,In_494);
and U318 (N_318,In_418,In_100);
nor U319 (N_319,In_150,In_16);
or U320 (N_320,In_218,In_443);
nor U321 (N_321,In_202,In_369);
or U322 (N_322,In_436,In_413);
and U323 (N_323,In_326,In_43);
nor U324 (N_324,In_6,In_163);
nor U325 (N_325,In_356,In_326);
or U326 (N_326,In_485,In_144);
nand U327 (N_327,In_236,In_122);
xnor U328 (N_328,In_123,In_126);
or U329 (N_329,In_301,In_462);
or U330 (N_330,In_124,In_226);
nand U331 (N_331,In_497,In_345);
and U332 (N_332,In_337,In_110);
or U333 (N_333,In_408,In_68);
or U334 (N_334,In_24,In_395);
and U335 (N_335,In_239,In_353);
nor U336 (N_336,In_494,In_165);
and U337 (N_337,In_445,In_332);
nor U338 (N_338,In_337,In_363);
or U339 (N_339,In_19,In_218);
nand U340 (N_340,In_272,In_400);
xnor U341 (N_341,In_20,In_86);
or U342 (N_342,In_244,In_383);
and U343 (N_343,In_325,In_359);
nand U344 (N_344,In_478,In_37);
xor U345 (N_345,In_276,In_36);
and U346 (N_346,In_21,In_481);
xnor U347 (N_347,In_264,In_466);
or U348 (N_348,In_449,In_316);
nand U349 (N_349,In_144,In_380);
xnor U350 (N_350,In_292,In_65);
or U351 (N_351,In_112,In_69);
and U352 (N_352,In_146,In_100);
nand U353 (N_353,In_67,In_450);
and U354 (N_354,In_435,In_183);
and U355 (N_355,In_37,In_4);
nor U356 (N_356,In_5,In_115);
and U357 (N_357,In_189,In_315);
xor U358 (N_358,In_244,In_173);
nand U359 (N_359,In_46,In_334);
or U360 (N_360,In_310,In_156);
or U361 (N_361,In_104,In_93);
or U362 (N_362,In_52,In_446);
xnor U363 (N_363,In_383,In_256);
and U364 (N_364,In_404,In_104);
or U365 (N_365,In_367,In_147);
or U366 (N_366,In_431,In_112);
nor U367 (N_367,In_153,In_258);
nand U368 (N_368,In_321,In_225);
or U369 (N_369,In_466,In_238);
nand U370 (N_370,In_96,In_287);
and U371 (N_371,In_17,In_459);
xor U372 (N_372,In_119,In_464);
xor U373 (N_373,In_488,In_434);
nand U374 (N_374,In_403,In_90);
nand U375 (N_375,In_477,In_177);
or U376 (N_376,In_240,In_82);
nand U377 (N_377,In_327,In_36);
and U378 (N_378,In_443,In_332);
nor U379 (N_379,In_234,In_333);
or U380 (N_380,In_208,In_48);
and U381 (N_381,In_468,In_52);
or U382 (N_382,In_441,In_230);
and U383 (N_383,In_334,In_404);
or U384 (N_384,In_100,In_494);
and U385 (N_385,In_81,In_49);
nand U386 (N_386,In_271,In_341);
nor U387 (N_387,In_375,In_119);
xnor U388 (N_388,In_459,In_251);
and U389 (N_389,In_19,In_362);
or U390 (N_390,In_70,In_492);
and U391 (N_391,In_241,In_25);
and U392 (N_392,In_97,In_153);
or U393 (N_393,In_358,In_243);
or U394 (N_394,In_301,In_431);
or U395 (N_395,In_471,In_314);
nand U396 (N_396,In_208,In_299);
nor U397 (N_397,In_273,In_266);
nand U398 (N_398,In_342,In_334);
and U399 (N_399,In_350,In_26);
and U400 (N_400,In_291,In_423);
or U401 (N_401,In_165,In_255);
xnor U402 (N_402,In_235,In_264);
or U403 (N_403,In_395,In_337);
or U404 (N_404,In_472,In_397);
nor U405 (N_405,In_374,In_323);
and U406 (N_406,In_191,In_285);
or U407 (N_407,In_175,In_315);
nand U408 (N_408,In_220,In_150);
and U409 (N_409,In_449,In_94);
nor U410 (N_410,In_344,In_18);
or U411 (N_411,In_82,In_129);
xor U412 (N_412,In_345,In_324);
nand U413 (N_413,In_352,In_238);
nor U414 (N_414,In_380,In_64);
and U415 (N_415,In_314,In_466);
xnor U416 (N_416,In_340,In_315);
or U417 (N_417,In_75,In_322);
nor U418 (N_418,In_223,In_301);
nor U419 (N_419,In_11,In_373);
and U420 (N_420,In_291,In_20);
xor U421 (N_421,In_113,In_216);
nand U422 (N_422,In_91,In_181);
and U423 (N_423,In_484,In_347);
and U424 (N_424,In_192,In_70);
and U425 (N_425,In_453,In_119);
nand U426 (N_426,In_100,In_421);
nor U427 (N_427,In_40,In_15);
nand U428 (N_428,In_440,In_89);
nor U429 (N_429,In_305,In_162);
nand U430 (N_430,In_302,In_381);
nand U431 (N_431,In_141,In_478);
xor U432 (N_432,In_349,In_348);
nand U433 (N_433,In_191,In_32);
or U434 (N_434,In_334,In_183);
or U435 (N_435,In_160,In_334);
and U436 (N_436,In_284,In_468);
nand U437 (N_437,In_363,In_356);
or U438 (N_438,In_377,In_142);
nor U439 (N_439,In_182,In_309);
nor U440 (N_440,In_356,In_338);
xor U441 (N_441,In_155,In_340);
nor U442 (N_442,In_324,In_441);
nand U443 (N_443,In_69,In_291);
nand U444 (N_444,In_234,In_331);
and U445 (N_445,In_212,In_279);
or U446 (N_446,In_467,In_77);
nand U447 (N_447,In_278,In_153);
nand U448 (N_448,In_29,In_322);
xnor U449 (N_449,In_450,In_276);
and U450 (N_450,In_232,In_408);
xnor U451 (N_451,In_395,In_1);
xnor U452 (N_452,In_4,In_405);
nand U453 (N_453,In_289,In_37);
nand U454 (N_454,In_372,In_367);
nand U455 (N_455,In_44,In_353);
nand U456 (N_456,In_64,In_368);
or U457 (N_457,In_430,In_119);
xor U458 (N_458,In_143,In_242);
or U459 (N_459,In_242,In_277);
nor U460 (N_460,In_294,In_479);
or U461 (N_461,In_319,In_387);
nor U462 (N_462,In_389,In_370);
nand U463 (N_463,In_327,In_9);
nand U464 (N_464,In_76,In_396);
nor U465 (N_465,In_192,In_13);
and U466 (N_466,In_44,In_390);
xor U467 (N_467,In_132,In_437);
or U468 (N_468,In_401,In_31);
nand U469 (N_469,In_419,In_84);
and U470 (N_470,In_38,In_272);
nand U471 (N_471,In_96,In_440);
xor U472 (N_472,In_311,In_405);
or U473 (N_473,In_412,In_123);
nand U474 (N_474,In_436,In_437);
and U475 (N_475,In_80,In_135);
or U476 (N_476,In_396,In_33);
xnor U477 (N_477,In_200,In_211);
nand U478 (N_478,In_489,In_8);
nand U479 (N_479,In_277,In_265);
or U480 (N_480,In_166,In_237);
nor U481 (N_481,In_289,In_403);
or U482 (N_482,In_354,In_417);
nand U483 (N_483,In_423,In_499);
nand U484 (N_484,In_354,In_362);
or U485 (N_485,In_489,In_138);
or U486 (N_486,In_267,In_487);
nor U487 (N_487,In_166,In_161);
or U488 (N_488,In_403,In_71);
or U489 (N_489,In_308,In_259);
or U490 (N_490,In_33,In_174);
nand U491 (N_491,In_361,In_373);
or U492 (N_492,In_202,In_80);
nor U493 (N_493,In_145,In_345);
xnor U494 (N_494,In_157,In_203);
nor U495 (N_495,In_107,In_258);
or U496 (N_496,In_129,In_226);
nand U497 (N_497,In_129,In_370);
or U498 (N_498,In_197,In_496);
nand U499 (N_499,In_321,In_352);
and U500 (N_500,In_44,In_223);
nor U501 (N_501,In_171,In_431);
or U502 (N_502,In_221,In_187);
and U503 (N_503,In_344,In_495);
xnor U504 (N_504,In_294,In_6);
nand U505 (N_505,In_384,In_287);
or U506 (N_506,In_268,In_242);
nor U507 (N_507,In_222,In_425);
nor U508 (N_508,In_14,In_434);
and U509 (N_509,In_274,In_384);
nand U510 (N_510,In_107,In_488);
nor U511 (N_511,In_422,In_459);
and U512 (N_512,In_298,In_404);
or U513 (N_513,In_344,In_130);
nand U514 (N_514,In_228,In_75);
and U515 (N_515,In_274,In_499);
nand U516 (N_516,In_16,In_84);
nor U517 (N_517,In_496,In_357);
and U518 (N_518,In_225,In_258);
xor U519 (N_519,In_150,In_158);
nand U520 (N_520,In_44,In_192);
nand U521 (N_521,In_135,In_371);
and U522 (N_522,In_469,In_344);
nor U523 (N_523,In_323,In_417);
nor U524 (N_524,In_442,In_343);
nand U525 (N_525,In_170,In_449);
or U526 (N_526,In_298,In_470);
nand U527 (N_527,In_218,In_405);
or U528 (N_528,In_394,In_262);
or U529 (N_529,In_468,In_490);
or U530 (N_530,In_156,In_470);
or U531 (N_531,In_116,In_310);
xnor U532 (N_532,In_484,In_252);
nor U533 (N_533,In_423,In_1);
nor U534 (N_534,In_182,In_422);
nand U535 (N_535,In_74,In_153);
and U536 (N_536,In_78,In_67);
xor U537 (N_537,In_444,In_119);
and U538 (N_538,In_170,In_309);
nor U539 (N_539,In_134,In_57);
or U540 (N_540,In_347,In_166);
nor U541 (N_541,In_406,In_250);
nand U542 (N_542,In_403,In_297);
and U543 (N_543,In_309,In_101);
or U544 (N_544,In_398,In_83);
nor U545 (N_545,In_387,In_255);
and U546 (N_546,In_169,In_402);
nand U547 (N_547,In_44,In_23);
nor U548 (N_548,In_116,In_215);
and U549 (N_549,In_54,In_210);
and U550 (N_550,In_159,In_268);
or U551 (N_551,In_254,In_160);
and U552 (N_552,In_438,In_154);
nand U553 (N_553,In_409,In_122);
nor U554 (N_554,In_22,In_243);
nor U555 (N_555,In_194,In_5);
nand U556 (N_556,In_481,In_370);
nor U557 (N_557,In_423,In_6);
nor U558 (N_558,In_268,In_387);
nand U559 (N_559,In_123,In_150);
nand U560 (N_560,In_358,In_154);
nor U561 (N_561,In_332,In_375);
or U562 (N_562,In_70,In_357);
nor U563 (N_563,In_8,In_63);
nand U564 (N_564,In_463,In_493);
nor U565 (N_565,In_298,In_426);
nor U566 (N_566,In_408,In_330);
and U567 (N_567,In_317,In_259);
or U568 (N_568,In_423,In_465);
or U569 (N_569,In_167,In_162);
and U570 (N_570,In_50,In_44);
and U571 (N_571,In_50,In_11);
or U572 (N_572,In_217,In_332);
nor U573 (N_573,In_41,In_76);
nand U574 (N_574,In_273,In_331);
nand U575 (N_575,In_263,In_460);
or U576 (N_576,In_246,In_268);
nor U577 (N_577,In_207,In_274);
xnor U578 (N_578,In_256,In_122);
or U579 (N_579,In_207,In_258);
nand U580 (N_580,In_77,In_364);
nor U581 (N_581,In_419,In_231);
and U582 (N_582,In_252,In_154);
or U583 (N_583,In_335,In_381);
or U584 (N_584,In_32,In_272);
nor U585 (N_585,In_362,In_299);
nand U586 (N_586,In_79,In_392);
and U587 (N_587,In_81,In_281);
and U588 (N_588,In_172,In_481);
or U589 (N_589,In_341,In_209);
xor U590 (N_590,In_279,In_199);
xor U591 (N_591,In_327,In_144);
and U592 (N_592,In_239,In_390);
or U593 (N_593,In_419,In_224);
or U594 (N_594,In_311,In_193);
and U595 (N_595,In_250,In_170);
or U596 (N_596,In_354,In_224);
nor U597 (N_597,In_143,In_424);
or U598 (N_598,In_130,In_223);
xnor U599 (N_599,In_464,In_149);
or U600 (N_600,In_246,In_328);
nand U601 (N_601,In_293,In_108);
or U602 (N_602,In_268,In_428);
nor U603 (N_603,In_107,In_386);
nand U604 (N_604,In_219,In_192);
or U605 (N_605,In_93,In_151);
nor U606 (N_606,In_63,In_14);
or U607 (N_607,In_153,In_396);
and U608 (N_608,In_85,In_427);
and U609 (N_609,In_174,In_473);
and U610 (N_610,In_424,In_410);
and U611 (N_611,In_431,In_308);
xnor U612 (N_612,In_385,In_131);
and U613 (N_613,In_346,In_249);
nor U614 (N_614,In_483,In_65);
or U615 (N_615,In_179,In_312);
xnor U616 (N_616,In_426,In_178);
or U617 (N_617,In_354,In_243);
or U618 (N_618,In_486,In_344);
and U619 (N_619,In_390,In_25);
and U620 (N_620,In_31,In_203);
nand U621 (N_621,In_20,In_87);
and U622 (N_622,In_174,In_273);
or U623 (N_623,In_366,In_274);
nor U624 (N_624,In_165,In_227);
and U625 (N_625,In_494,In_362);
nor U626 (N_626,In_397,In_183);
or U627 (N_627,In_18,In_339);
and U628 (N_628,In_111,In_49);
and U629 (N_629,In_74,In_182);
nand U630 (N_630,In_287,In_386);
or U631 (N_631,In_111,In_70);
nand U632 (N_632,In_81,In_286);
nor U633 (N_633,In_259,In_499);
nand U634 (N_634,In_35,In_298);
nor U635 (N_635,In_388,In_81);
nor U636 (N_636,In_410,In_162);
nor U637 (N_637,In_46,In_263);
nor U638 (N_638,In_11,In_432);
or U639 (N_639,In_57,In_348);
nand U640 (N_640,In_332,In_382);
and U641 (N_641,In_223,In_244);
nor U642 (N_642,In_155,In_64);
xor U643 (N_643,In_56,In_81);
xnor U644 (N_644,In_148,In_291);
nor U645 (N_645,In_7,In_401);
and U646 (N_646,In_254,In_338);
nor U647 (N_647,In_318,In_263);
and U648 (N_648,In_215,In_489);
or U649 (N_649,In_170,In_498);
nor U650 (N_650,In_343,In_302);
nand U651 (N_651,In_109,In_245);
nor U652 (N_652,In_72,In_334);
xor U653 (N_653,In_123,In_368);
and U654 (N_654,In_457,In_379);
and U655 (N_655,In_8,In_59);
or U656 (N_656,In_68,In_188);
nand U657 (N_657,In_139,In_306);
nand U658 (N_658,In_71,In_143);
nand U659 (N_659,In_243,In_233);
nand U660 (N_660,In_260,In_41);
or U661 (N_661,In_131,In_90);
and U662 (N_662,In_215,In_406);
nor U663 (N_663,In_454,In_140);
nand U664 (N_664,In_90,In_16);
nor U665 (N_665,In_10,In_291);
xor U666 (N_666,In_266,In_87);
or U667 (N_667,In_485,In_105);
xnor U668 (N_668,In_311,In_342);
nand U669 (N_669,In_498,In_259);
and U670 (N_670,In_92,In_461);
nand U671 (N_671,In_19,In_121);
or U672 (N_672,In_186,In_449);
nor U673 (N_673,In_111,In_399);
nand U674 (N_674,In_37,In_108);
nor U675 (N_675,In_97,In_490);
nor U676 (N_676,In_461,In_35);
and U677 (N_677,In_454,In_390);
nand U678 (N_678,In_161,In_171);
nand U679 (N_679,In_387,In_3);
nor U680 (N_680,In_468,In_455);
and U681 (N_681,In_340,In_391);
or U682 (N_682,In_415,In_444);
nor U683 (N_683,In_149,In_252);
nand U684 (N_684,In_361,In_345);
xnor U685 (N_685,In_68,In_182);
xor U686 (N_686,In_458,In_376);
nand U687 (N_687,In_222,In_24);
nor U688 (N_688,In_253,In_72);
xor U689 (N_689,In_110,In_417);
nand U690 (N_690,In_425,In_59);
and U691 (N_691,In_418,In_467);
or U692 (N_692,In_477,In_259);
and U693 (N_693,In_485,In_13);
nor U694 (N_694,In_2,In_386);
xnor U695 (N_695,In_485,In_164);
nor U696 (N_696,In_478,In_164);
and U697 (N_697,In_118,In_164);
nor U698 (N_698,In_206,In_55);
and U699 (N_699,In_61,In_447);
or U700 (N_700,In_359,In_134);
and U701 (N_701,In_117,In_496);
nand U702 (N_702,In_440,In_93);
xnor U703 (N_703,In_388,In_359);
nand U704 (N_704,In_336,In_68);
and U705 (N_705,In_243,In_327);
nor U706 (N_706,In_391,In_23);
and U707 (N_707,In_437,In_123);
and U708 (N_708,In_436,In_466);
nand U709 (N_709,In_68,In_427);
and U710 (N_710,In_209,In_476);
xnor U711 (N_711,In_125,In_230);
nor U712 (N_712,In_138,In_66);
nor U713 (N_713,In_327,In_393);
nor U714 (N_714,In_218,In_407);
or U715 (N_715,In_460,In_146);
and U716 (N_716,In_183,In_478);
and U717 (N_717,In_11,In_310);
and U718 (N_718,In_413,In_188);
nor U719 (N_719,In_443,In_340);
and U720 (N_720,In_192,In_260);
and U721 (N_721,In_211,In_495);
or U722 (N_722,In_430,In_414);
nand U723 (N_723,In_271,In_177);
nor U724 (N_724,In_454,In_275);
or U725 (N_725,In_466,In_422);
nand U726 (N_726,In_272,In_446);
nand U727 (N_727,In_141,In_458);
nor U728 (N_728,In_239,In_346);
and U729 (N_729,In_114,In_344);
nand U730 (N_730,In_169,In_13);
xor U731 (N_731,In_64,In_451);
and U732 (N_732,In_26,In_73);
or U733 (N_733,In_449,In_415);
and U734 (N_734,In_486,In_142);
nand U735 (N_735,In_319,In_25);
or U736 (N_736,In_346,In_285);
nand U737 (N_737,In_172,In_383);
nor U738 (N_738,In_110,In_72);
nand U739 (N_739,In_338,In_343);
or U740 (N_740,In_397,In_201);
or U741 (N_741,In_290,In_461);
and U742 (N_742,In_389,In_138);
xor U743 (N_743,In_235,In_110);
and U744 (N_744,In_428,In_114);
nor U745 (N_745,In_331,In_248);
or U746 (N_746,In_194,In_127);
or U747 (N_747,In_39,In_118);
nand U748 (N_748,In_186,In_348);
or U749 (N_749,In_492,In_205);
or U750 (N_750,N_268,N_617);
or U751 (N_751,N_40,N_53);
and U752 (N_752,N_726,N_701);
nand U753 (N_753,N_76,N_517);
and U754 (N_754,N_524,N_662);
nand U755 (N_755,N_485,N_78);
or U756 (N_756,N_318,N_528);
nor U757 (N_757,N_738,N_716);
xnor U758 (N_758,N_699,N_3);
nand U759 (N_759,N_746,N_704);
nand U760 (N_760,N_461,N_741);
nor U761 (N_761,N_543,N_276);
nor U762 (N_762,N_2,N_630);
xor U763 (N_763,N_436,N_719);
and U764 (N_764,N_739,N_643);
nor U765 (N_765,N_179,N_170);
nand U766 (N_766,N_545,N_359);
nor U767 (N_767,N_23,N_456);
nor U768 (N_768,N_642,N_167);
nor U769 (N_769,N_408,N_293);
and U770 (N_770,N_392,N_618);
nor U771 (N_771,N_526,N_396);
nor U772 (N_772,N_475,N_64);
or U773 (N_773,N_164,N_422);
nor U774 (N_774,N_652,N_674);
xor U775 (N_775,N_549,N_284);
and U776 (N_776,N_532,N_636);
and U777 (N_777,N_369,N_554);
nor U778 (N_778,N_41,N_469);
and U779 (N_779,N_627,N_609);
and U780 (N_780,N_468,N_244);
nand U781 (N_781,N_356,N_625);
nand U782 (N_782,N_177,N_105);
xnor U783 (N_783,N_731,N_744);
or U784 (N_784,N_459,N_671);
xor U785 (N_785,N_591,N_593);
or U786 (N_786,N_334,N_620);
nand U787 (N_787,N_142,N_339);
and U788 (N_788,N_711,N_421);
nor U789 (N_789,N_663,N_646);
or U790 (N_790,N_202,N_95);
nor U791 (N_791,N_127,N_218);
or U792 (N_792,N_564,N_264);
nand U793 (N_793,N_375,N_668);
or U794 (N_794,N_444,N_92);
and U795 (N_795,N_709,N_196);
nand U796 (N_796,N_603,N_145);
nor U797 (N_797,N_180,N_495);
xnor U798 (N_798,N_217,N_614);
nand U799 (N_799,N_346,N_581);
and U800 (N_800,N_515,N_353);
or U801 (N_801,N_171,N_498);
or U802 (N_802,N_189,N_83);
or U803 (N_803,N_133,N_670);
nor U804 (N_804,N_60,N_633);
nor U805 (N_805,N_109,N_67);
and U806 (N_806,N_404,N_393);
nand U807 (N_807,N_479,N_123);
nor U808 (N_808,N_350,N_374);
xor U809 (N_809,N_44,N_156);
nor U810 (N_810,N_132,N_598);
nand U811 (N_811,N_52,N_11);
nor U812 (N_812,N_727,N_190);
and U813 (N_813,N_286,N_558);
nand U814 (N_814,N_223,N_693);
or U815 (N_815,N_557,N_735);
nor U816 (N_816,N_706,N_490);
nand U817 (N_817,N_653,N_397);
and U818 (N_818,N_313,N_601);
nor U819 (N_819,N_446,N_702);
nand U820 (N_820,N_120,N_358);
and U821 (N_821,N_106,N_722);
nand U822 (N_822,N_616,N_429);
nor U823 (N_823,N_417,N_426);
and U824 (N_824,N_107,N_473);
and U825 (N_825,N_519,N_172);
and U826 (N_826,N_206,N_118);
nor U827 (N_827,N_541,N_610);
and U828 (N_828,N_457,N_724);
and U829 (N_829,N_466,N_125);
nor U830 (N_830,N_730,N_624);
nand U831 (N_831,N_667,N_146);
nor U832 (N_832,N_553,N_450);
nor U833 (N_833,N_277,N_483);
nand U834 (N_834,N_523,N_471);
and U835 (N_835,N_732,N_599);
nand U836 (N_836,N_338,N_654);
and U837 (N_837,N_607,N_569);
nand U838 (N_838,N_292,N_579);
and U839 (N_839,N_74,N_715);
nor U840 (N_840,N_342,N_666);
and U841 (N_841,N_373,N_305);
or U842 (N_842,N_583,N_477);
nor U843 (N_843,N_198,N_147);
and U844 (N_844,N_410,N_93);
nand U845 (N_845,N_150,N_547);
xor U846 (N_846,N_207,N_291);
or U847 (N_847,N_447,N_182);
nand U848 (N_848,N_345,N_22);
xor U849 (N_849,N_298,N_499);
nor U850 (N_850,N_413,N_559);
or U851 (N_851,N_476,N_259);
xor U852 (N_852,N_655,N_637);
and U853 (N_853,N_534,N_449);
nor U854 (N_854,N_173,N_327);
and U855 (N_855,N_234,N_194);
or U856 (N_856,N_605,N_256);
nand U857 (N_857,N_341,N_491);
nand U858 (N_858,N_337,N_565);
nand U859 (N_859,N_721,N_432);
and U860 (N_860,N_503,N_104);
and U861 (N_861,N_357,N_333);
nand U862 (N_862,N_352,N_219);
nand U863 (N_863,N_33,N_175);
and U864 (N_864,N_14,N_378);
and U865 (N_865,N_29,N_214);
nor U866 (N_866,N_425,N_650);
nor U867 (N_867,N_84,N_336);
nand U868 (N_868,N_690,N_343);
and U869 (N_869,N_227,N_560);
nand U870 (N_870,N_148,N_312);
or U871 (N_871,N_297,N_65);
or U872 (N_872,N_283,N_696);
or U873 (N_873,N_710,N_188);
nor U874 (N_874,N_323,N_45);
nand U875 (N_875,N_428,N_486);
and U876 (N_876,N_191,N_243);
nor U877 (N_877,N_561,N_500);
and U878 (N_878,N_258,N_61);
nor U879 (N_879,N_497,N_159);
or U880 (N_880,N_280,N_440);
or U881 (N_881,N_31,N_448);
nor U882 (N_882,N_460,N_362);
nand U883 (N_883,N_20,N_508);
and U884 (N_884,N_600,N_433);
and U885 (N_885,N_394,N_376);
nor U886 (N_886,N_563,N_377);
nand U887 (N_887,N_664,N_400);
and U888 (N_888,N_493,N_262);
nor U889 (N_889,N_586,N_574);
nor U890 (N_890,N_472,N_686);
xnor U891 (N_891,N_529,N_749);
nand U892 (N_892,N_8,N_246);
nand U893 (N_893,N_71,N_665);
xor U894 (N_894,N_530,N_411);
and U895 (N_895,N_482,N_324);
nand U896 (N_896,N_689,N_678);
nand U897 (N_897,N_587,N_229);
nor U898 (N_898,N_58,N_301);
or U899 (N_899,N_521,N_615);
or U900 (N_900,N_208,N_86);
nand U901 (N_901,N_504,N_439);
nand U902 (N_902,N_679,N_306);
and U903 (N_903,N_251,N_101);
nor U904 (N_904,N_474,N_489);
nor U905 (N_905,N_568,N_114);
nand U906 (N_906,N_38,N_340);
or U907 (N_907,N_518,N_351);
nand U908 (N_908,N_103,N_10);
nor U909 (N_909,N_232,N_325);
and U910 (N_910,N_225,N_386);
or U911 (N_911,N_492,N_209);
or U912 (N_912,N_108,N_275);
or U913 (N_913,N_516,N_250);
nand U914 (N_914,N_228,N_718);
and U915 (N_915,N_512,N_619);
nand U916 (N_916,N_237,N_181);
nor U917 (N_917,N_431,N_302);
and U918 (N_918,N_94,N_349);
and U919 (N_919,N_274,N_418);
nand U920 (N_920,N_590,N_688);
nor U921 (N_921,N_612,N_72);
nand U922 (N_922,N_570,N_155);
or U923 (N_923,N_366,N_430);
nor U924 (N_924,N_698,N_119);
and U925 (N_925,N_454,N_49);
nand U926 (N_926,N_695,N_205);
or U927 (N_927,N_585,N_348);
nor U928 (N_928,N_645,N_131);
nand U929 (N_929,N_462,N_632);
and U930 (N_930,N_520,N_319);
xnor U931 (N_931,N_354,N_660);
nand U932 (N_932,N_314,N_389);
or U933 (N_933,N_21,N_405);
nor U934 (N_934,N_443,N_556);
nand U935 (N_935,N_287,N_494);
or U936 (N_936,N_531,N_562);
nand U937 (N_937,N_659,N_136);
or U938 (N_938,N_371,N_423);
or U939 (N_939,N_157,N_81);
nor U940 (N_940,N_282,N_143);
or U941 (N_941,N_121,N_658);
xor U942 (N_942,N_745,N_629);
nand U943 (N_943,N_737,N_365);
nand U944 (N_944,N_253,N_210);
or U945 (N_945,N_16,N_195);
nand U946 (N_946,N_192,N_395);
or U947 (N_947,N_183,N_437);
and U948 (N_948,N_154,N_149);
nand U949 (N_949,N_289,N_685);
or U950 (N_950,N_278,N_647);
or U951 (N_951,N_248,N_233);
or U952 (N_952,N_542,N_75);
nand U953 (N_953,N_46,N_743);
or U954 (N_954,N_728,N_481);
and U955 (N_955,N_380,N_139);
and U956 (N_956,N_162,N_204);
and U957 (N_957,N_55,N_129);
or U958 (N_958,N_240,N_267);
nand U959 (N_959,N_80,N_594);
nor U960 (N_960,N_317,N_384);
and U961 (N_961,N_546,N_263);
nor U962 (N_962,N_257,N_199);
and U963 (N_963,N_606,N_163);
nand U964 (N_964,N_17,N_288);
and U965 (N_965,N_115,N_220);
and U966 (N_966,N_368,N_300);
or U967 (N_967,N_187,N_303);
and U968 (N_968,N_128,N_506);
nand U969 (N_969,N_539,N_69);
nor U970 (N_970,N_725,N_370);
or U971 (N_971,N_551,N_420);
or U972 (N_972,N_91,N_124);
nand U973 (N_973,N_295,N_639);
or U974 (N_974,N_236,N_35);
xnor U975 (N_975,N_714,N_381);
nor U976 (N_976,N_403,N_501);
nand U977 (N_977,N_649,N_215);
and U978 (N_978,N_552,N_273);
nor U979 (N_979,N_672,N_505);
nand U980 (N_980,N_19,N_544);
nand U981 (N_981,N_153,N_322);
nor U982 (N_982,N_63,N_235);
xor U983 (N_983,N_224,N_510);
xor U984 (N_984,N_211,N_166);
or U985 (N_985,N_299,N_419);
nor U986 (N_986,N_496,N_379);
and U987 (N_987,N_613,N_56);
nand U988 (N_988,N_126,N_307);
nor U989 (N_989,N_705,N_51);
nor U990 (N_990,N_290,N_675);
nor U991 (N_991,N_608,N_144);
nand U992 (N_992,N_97,N_239);
xor U993 (N_993,N_241,N_548);
and U994 (N_994,N_623,N_245);
or U995 (N_995,N_242,N_85);
xor U996 (N_996,N_635,N_644);
nand U997 (N_997,N_39,N_116);
nor U998 (N_998,N_382,N_390);
and U999 (N_999,N_222,N_113);
or U1000 (N_1000,N_648,N_112);
nand U1001 (N_1001,N_28,N_742);
or U1002 (N_1002,N_596,N_626);
and U1003 (N_1003,N_509,N_576);
nand U1004 (N_1004,N_406,N_36);
nor U1005 (N_1005,N_470,N_455);
and U1006 (N_1006,N_255,N_463);
and U1007 (N_1007,N_582,N_513);
and U1008 (N_1008,N_178,N_174);
or U1009 (N_1009,N_584,N_73);
xor U1010 (N_1010,N_458,N_18);
and U1011 (N_1011,N_117,N_604);
nor U1012 (N_1012,N_82,N_185);
nand U1013 (N_1013,N_684,N_331);
or U1014 (N_1014,N_270,N_90);
or U1015 (N_1015,N_522,N_733);
or U1016 (N_1016,N_628,N_151);
and U1017 (N_1017,N_260,N_507);
nand U1018 (N_1018,N_427,N_575);
nor U1019 (N_1019,N_577,N_525);
and U1020 (N_1020,N_538,N_141);
or U1021 (N_1021,N_445,N_669);
nor U1022 (N_1022,N_661,N_310);
or U1023 (N_1023,N_621,N_514);
nor U1024 (N_1024,N_186,N_567);
nor U1025 (N_1025,N_453,N_111);
or U1026 (N_1026,N_388,N_98);
xnor U1027 (N_1027,N_311,N_79);
nor U1028 (N_1028,N_533,N_578);
nor U1029 (N_1029,N_168,N_32);
nor U1030 (N_1030,N_50,N_502);
xnor U1031 (N_1031,N_611,N_140);
xnor U1032 (N_1032,N_9,N_296);
xnor U1033 (N_1033,N_634,N_638);
nand U1034 (N_1034,N_309,N_326);
nor U1035 (N_1035,N_595,N_673);
nand U1036 (N_1036,N_321,N_62);
nor U1037 (N_1037,N_30,N_385);
nand U1038 (N_1038,N_713,N_285);
nand U1039 (N_1039,N_691,N_102);
and U1040 (N_1040,N_47,N_230);
xor U1041 (N_1041,N_27,N_720);
and U1042 (N_1042,N_320,N_201);
nor U1043 (N_1043,N_137,N_54);
xor U1044 (N_1044,N_57,N_527);
xor U1045 (N_1045,N_100,N_451);
and U1046 (N_1046,N_70,N_740);
and U1047 (N_1047,N_435,N_1);
xnor U1048 (N_1048,N_484,N_398);
and U1049 (N_1049,N_48,N_99);
or U1050 (N_1050,N_316,N_4);
or U1051 (N_1051,N_364,N_572);
xor U1052 (N_1052,N_238,N_434);
or U1053 (N_1053,N_87,N_399);
and U1054 (N_1054,N_536,N_573);
xor U1055 (N_1055,N_347,N_169);
and U1056 (N_1056,N_640,N_387);
nand U1057 (N_1057,N_37,N_330);
nor U1058 (N_1058,N_703,N_416);
nand U1059 (N_1059,N_414,N_452);
xor U1060 (N_1060,N_708,N_602);
nor U1061 (N_1061,N_135,N_252);
or U1062 (N_1062,N_261,N_656);
nor U1063 (N_1063,N_5,N_465);
nor U1064 (N_1064,N_747,N_161);
or U1065 (N_1065,N_26,N_367);
nor U1066 (N_1066,N_25,N_402);
and U1067 (N_1067,N_77,N_335);
or U1068 (N_1068,N_677,N_328);
and U1069 (N_1069,N_265,N_226);
nor U1070 (N_1070,N_681,N_729);
nor U1071 (N_1071,N_193,N_736);
xor U1072 (N_1072,N_221,N_355);
nand U1073 (N_1073,N_308,N_130);
nand U1074 (N_1074,N_247,N_134);
or U1075 (N_1075,N_372,N_160);
xor U1076 (N_1076,N_203,N_271);
nand U1077 (N_1077,N_580,N_279);
or U1078 (N_1078,N_329,N_0);
and U1079 (N_1079,N_680,N_24);
nand U1080 (N_1080,N_266,N_361);
or U1081 (N_1081,N_651,N_566);
nor U1082 (N_1082,N_478,N_409);
or U1083 (N_1083,N_734,N_687);
and U1084 (N_1084,N_294,N_487);
xor U1085 (N_1085,N_212,N_692);
nor U1086 (N_1086,N_571,N_415);
nand U1087 (N_1087,N_200,N_269);
and U1088 (N_1088,N_344,N_412);
or U1089 (N_1089,N_438,N_138);
xnor U1090 (N_1090,N_12,N_272);
or U1091 (N_1091,N_34,N_657);
or U1092 (N_1092,N_712,N_676);
nand U1093 (N_1093,N_537,N_363);
nand U1094 (N_1094,N_68,N_42);
or U1095 (N_1095,N_480,N_360);
and U1096 (N_1096,N_122,N_697);
or U1097 (N_1097,N_231,N_592);
or U1098 (N_1098,N_110,N_622);
and U1099 (N_1099,N_249,N_213);
or U1100 (N_1100,N_281,N_424);
xor U1101 (N_1101,N_184,N_641);
nand U1102 (N_1102,N_401,N_89);
and U1103 (N_1103,N_723,N_707);
or U1104 (N_1104,N_13,N_165);
nor U1105 (N_1105,N_682,N_748);
or U1106 (N_1106,N_597,N_152);
or U1107 (N_1107,N_588,N_7);
nand U1108 (N_1108,N_464,N_304);
or U1109 (N_1109,N_158,N_550);
nand U1110 (N_1110,N_683,N_511);
nor U1111 (N_1111,N_332,N_555);
and U1112 (N_1112,N_467,N_694);
or U1113 (N_1113,N_631,N_717);
and U1114 (N_1114,N_407,N_176);
xor U1115 (N_1115,N_315,N_383);
nand U1116 (N_1116,N_589,N_216);
nand U1117 (N_1117,N_700,N_59);
nor U1118 (N_1118,N_540,N_391);
and U1119 (N_1119,N_441,N_6);
nand U1120 (N_1120,N_254,N_96);
and U1121 (N_1121,N_442,N_43);
and U1122 (N_1122,N_197,N_488);
or U1123 (N_1123,N_88,N_66);
nor U1124 (N_1124,N_535,N_15);
nor U1125 (N_1125,N_562,N_81);
and U1126 (N_1126,N_303,N_536);
and U1127 (N_1127,N_258,N_440);
and U1128 (N_1128,N_559,N_577);
or U1129 (N_1129,N_480,N_484);
or U1130 (N_1130,N_706,N_605);
xor U1131 (N_1131,N_646,N_467);
xnor U1132 (N_1132,N_479,N_619);
or U1133 (N_1133,N_400,N_48);
or U1134 (N_1134,N_538,N_280);
nand U1135 (N_1135,N_45,N_354);
nor U1136 (N_1136,N_530,N_742);
nor U1137 (N_1137,N_409,N_477);
nor U1138 (N_1138,N_696,N_602);
or U1139 (N_1139,N_208,N_455);
and U1140 (N_1140,N_139,N_439);
nand U1141 (N_1141,N_434,N_419);
nor U1142 (N_1142,N_520,N_260);
nand U1143 (N_1143,N_543,N_615);
nand U1144 (N_1144,N_360,N_223);
nor U1145 (N_1145,N_212,N_445);
or U1146 (N_1146,N_149,N_551);
or U1147 (N_1147,N_693,N_225);
nand U1148 (N_1148,N_474,N_525);
or U1149 (N_1149,N_250,N_390);
and U1150 (N_1150,N_581,N_212);
nand U1151 (N_1151,N_199,N_64);
nand U1152 (N_1152,N_560,N_45);
and U1153 (N_1153,N_665,N_701);
nand U1154 (N_1154,N_256,N_5);
nand U1155 (N_1155,N_126,N_698);
nor U1156 (N_1156,N_529,N_696);
and U1157 (N_1157,N_173,N_428);
or U1158 (N_1158,N_580,N_471);
nand U1159 (N_1159,N_177,N_569);
and U1160 (N_1160,N_446,N_93);
and U1161 (N_1161,N_252,N_378);
and U1162 (N_1162,N_382,N_472);
nor U1163 (N_1163,N_206,N_560);
or U1164 (N_1164,N_568,N_511);
and U1165 (N_1165,N_301,N_604);
nor U1166 (N_1166,N_370,N_73);
nand U1167 (N_1167,N_201,N_326);
xnor U1168 (N_1168,N_411,N_684);
nand U1169 (N_1169,N_641,N_551);
nor U1170 (N_1170,N_631,N_304);
nor U1171 (N_1171,N_676,N_499);
or U1172 (N_1172,N_87,N_654);
nor U1173 (N_1173,N_411,N_298);
or U1174 (N_1174,N_697,N_655);
nand U1175 (N_1175,N_556,N_57);
or U1176 (N_1176,N_420,N_465);
nor U1177 (N_1177,N_351,N_181);
xor U1178 (N_1178,N_699,N_282);
and U1179 (N_1179,N_712,N_75);
nand U1180 (N_1180,N_164,N_689);
and U1181 (N_1181,N_20,N_559);
nor U1182 (N_1182,N_410,N_582);
and U1183 (N_1183,N_337,N_743);
nor U1184 (N_1184,N_190,N_297);
or U1185 (N_1185,N_326,N_71);
and U1186 (N_1186,N_649,N_402);
or U1187 (N_1187,N_681,N_208);
nor U1188 (N_1188,N_76,N_170);
or U1189 (N_1189,N_344,N_593);
and U1190 (N_1190,N_309,N_65);
nand U1191 (N_1191,N_561,N_212);
nor U1192 (N_1192,N_709,N_614);
and U1193 (N_1193,N_683,N_674);
and U1194 (N_1194,N_627,N_103);
nand U1195 (N_1195,N_629,N_572);
nand U1196 (N_1196,N_577,N_611);
nor U1197 (N_1197,N_129,N_704);
nand U1198 (N_1198,N_243,N_146);
and U1199 (N_1199,N_547,N_680);
nor U1200 (N_1200,N_226,N_325);
and U1201 (N_1201,N_695,N_88);
or U1202 (N_1202,N_350,N_52);
nor U1203 (N_1203,N_740,N_694);
and U1204 (N_1204,N_267,N_336);
and U1205 (N_1205,N_438,N_700);
xor U1206 (N_1206,N_265,N_395);
xnor U1207 (N_1207,N_83,N_712);
nand U1208 (N_1208,N_415,N_316);
and U1209 (N_1209,N_627,N_221);
and U1210 (N_1210,N_587,N_544);
nand U1211 (N_1211,N_25,N_639);
nand U1212 (N_1212,N_690,N_273);
nor U1213 (N_1213,N_63,N_359);
and U1214 (N_1214,N_147,N_588);
and U1215 (N_1215,N_516,N_744);
nor U1216 (N_1216,N_540,N_348);
or U1217 (N_1217,N_221,N_336);
and U1218 (N_1218,N_749,N_28);
nand U1219 (N_1219,N_525,N_67);
nor U1220 (N_1220,N_188,N_235);
or U1221 (N_1221,N_563,N_109);
or U1222 (N_1222,N_304,N_527);
xnor U1223 (N_1223,N_37,N_545);
or U1224 (N_1224,N_474,N_647);
nand U1225 (N_1225,N_576,N_634);
and U1226 (N_1226,N_311,N_733);
nand U1227 (N_1227,N_86,N_426);
and U1228 (N_1228,N_558,N_276);
nand U1229 (N_1229,N_46,N_264);
or U1230 (N_1230,N_115,N_490);
and U1231 (N_1231,N_563,N_289);
or U1232 (N_1232,N_710,N_101);
nor U1233 (N_1233,N_527,N_576);
nand U1234 (N_1234,N_21,N_399);
nor U1235 (N_1235,N_558,N_135);
or U1236 (N_1236,N_481,N_18);
nand U1237 (N_1237,N_96,N_552);
or U1238 (N_1238,N_743,N_301);
nand U1239 (N_1239,N_296,N_59);
or U1240 (N_1240,N_112,N_576);
nand U1241 (N_1241,N_708,N_154);
nor U1242 (N_1242,N_549,N_497);
nor U1243 (N_1243,N_437,N_257);
xor U1244 (N_1244,N_660,N_661);
and U1245 (N_1245,N_240,N_318);
nor U1246 (N_1246,N_458,N_593);
nor U1247 (N_1247,N_429,N_223);
xor U1248 (N_1248,N_260,N_453);
nor U1249 (N_1249,N_548,N_722);
and U1250 (N_1250,N_317,N_214);
or U1251 (N_1251,N_380,N_407);
xnor U1252 (N_1252,N_262,N_668);
nand U1253 (N_1253,N_353,N_489);
and U1254 (N_1254,N_86,N_508);
nand U1255 (N_1255,N_191,N_195);
nor U1256 (N_1256,N_538,N_30);
or U1257 (N_1257,N_487,N_632);
nor U1258 (N_1258,N_420,N_195);
or U1259 (N_1259,N_359,N_47);
or U1260 (N_1260,N_166,N_89);
nor U1261 (N_1261,N_59,N_361);
and U1262 (N_1262,N_323,N_73);
nor U1263 (N_1263,N_68,N_535);
and U1264 (N_1264,N_270,N_223);
nor U1265 (N_1265,N_468,N_663);
and U1266 (N_1266,N_460,N_721);
or U1267 (N_1267,N_707,N_675);
nand U1268 (N_1268,N_456,N_464);
and U1269 (N_1269,N_143,N_184);
or U1270 (N_1270,N_507,N_551);
and U1271 (N_1271,N_140,N_61);
xor U1272 (N_1272,N_404,N_585);
and U1273 (N_1273,N_183,N_632);
or U1274 (N_1274,N_219,N_42);
and U1275 (N_1275,N_354,N_36);
nor U1276 (N_1276,N_369,N_112);
or U1277 (N_1277,N_160,N_743);
nand U1278 (N_1278,N_46,N_196);
or U1279 (N_1279,N_556,N_681);
nor U1280 (N_1280,N_300,N_59);
nor U1281 (N_1281,N_652,N_382);
or U1282 (N_1282,N_15,N_49);
nor U1283 (N_1283,N_265,N_618);
nor U1284 (N_1284,N_273,N_632);
nor U1285 (N_1285,N_559,N_373);
or U1286 (N_1286,N_749,N_399);
and U1287 (N_1287,N_644,N_661);
or U1288 (N_1288,N_583,N_322);
nand U1289 (N_1289,N_92,N_381);
or U1290 (N_1290,N_714,N_557);
nand U1291 (N_1291,N_80,N_89);
nor U1292 (N_1292,N_307,N_707);
nand U1293 (N_1293,N_278,N_615);
and U1294 (N_1294,N_176,N_351);
xnor U1295 (N_1295,N_682,N_668);
and U1296 (N_1296,N_161,N_315);
and U1297 (N_1297,N_212,N_572);
and U1298 (N_1298,N_704,N_684);
or U1299 (N_1299,N_390,N_71);
or U1300 (N_1300,N_551,N_433);
or U1301 (N_1301,N_561,N_712);
and U1302 (N_1302,N_444,N_263);
or U1303 (N_1303,N_115,N_339);
nand U1304 (N_1304,N_203,N_607);
or U1305 (N_1305,N_209,N_620);
nor U1306 (N_1306,N_736,N_539);
nor U1307 (N_1307,N_106,N_480);
nor U1308 (N_1308,N_404,N_113);
nand U1309 (N_1309,N_91,N_116);
and U1310 (N_1310,N_265,N_172);
nor U1311 (N_1311,N_343,N_550);
nand U1312 (N_1312,N_245,N_622);
nor U1313 (N_1313,N_294,N_510);
or U1314 (N_1314,N_502,N_36);
nor U1315 (N_1315,N_238,N_262);
and U1316 (N_1316,N_274,N_62);
xnor U1317 (N_1317,N_342,N_487);
nand U1318 (N_1318,N_659,N_388);
and U1319 (N_1319,N_78,N_387);
nor U1320 (N_1320,N_706,N_506);
nand U1321 (N_1321,N_698,N_10);
nand U1322 (N_1322,N_141,N_117);
and U1323 (N_1323,N_624,N_475);
and U1324 (N_1324,N_261,N_678);
and U1325 (N_1325,N_730,N_533);
or U1326 (N_1326,N_690,N_382);
or U1327 (N_1327,N_148,N_675);
nand U1328 (N_1328,N_660,N_701);
nand U1329 (N_1329,N_600,N_30);
and U1330 (N_1330,N_620,N_90);
and U1331 (N_1331,N_59,N_460);
nand U1332 (N_1332,N_263,N_337);
nor U1333 (N_1333,N_202,N_237);
nor U1334 (N_1334,N_492,N_477);
nand U1335 (N_1335,N_180,N_96);
nor U1336 (N_1336,N_19,N_361);
xor U1337 (N_1337,N_577,N_550);
or U1338 (N_1338,N_644,N_104);
nor U1339 (N_1339,N_487,N_565);
or U1340 (N_1340,N_223,N_59);
nor U1341 (N_1341,N_335,N_426);
and U1342 (N_1342,N_95,N_277);
or U1343 (N_1343,N_24,N_9);
or U1344 (N_1344,N_73,N_581);
xnor U1345 (N_1345,N_545,N_220);
nor U1346 (N_1346,N_666,N_657);
and U1347 (N_1347,N_380,N_388);
or U1348 (N_1348,N_529,N_561);
and U1349 (N_1349,N_743,N_499);
or U1350 (N_1350,N_66,N_507);
nor U1351 (N_1351,N_624,N_482);
nor U1352 (N_1352,N_135,N_89);
and U1353 (N_1353,N_287,N_361);
and U1354 (N_1354,N_552,N_558);
nand U1355 (N_1355,N_665,N_604);
or U1356 (N_1356,N_434,N_204);
and U1357 (N_1357,N_234,N_0);
or U1358 (N_1358,N_665,N_296);
nand U1359 (N_1359,N_78,N_476);
xnor U1360 (N_1360,N_287,N_380);
nor U1361 (N_1361,N_573,N_222);
nor U1362 (N_1362,N_190,N_657);
and U1363 (N_1363,N_317,N_393);
and U1364 (N_1364,N_307,N_201);
nand U1365 (N_1365,N_283,N_446);
nand U1366 (N_1366,N_91,N_260);
and U1367 (N_1367,N_669,N_322);
nand U1368 (N_1368,N_690,N_141);
or U1369 (N_1369,N_85,N_668);
nor U1370 (N_1370,N_168,N_731);
nor U1371 (N_1371,N_744,N_143);
xnor U1372 (N_1372,N_340,N_246);
or U1373 (N_1373,N_513,N_715);
nand U1374 (N_1374,N_231,N_695);
nand U1375 (N_1375,N_388,N_695);
xor U1376 (N_1376,N_304,N_1);
or U1377 (N_1377,N_0,N_225);
nor U1378 (N_1378,N_130,N_701);
nor U1379 (N_1379,N_260,N_672);
and U1380 (N_1380,N_162,N_735);
nor U1381 (N_1381,N_656,N_414);
nor U1382 (N_1382,N_387,N_677);
or U1383 (N_1383,N_484,N_722);
and U1384 (N_1384,N_439,N_440);
nor U1385 (N_1385,N_659,N_439);
nor U1386 (N_1386,N_679,N_463);
or U1387 (N_1387,N_507,N_287);
nand U1388 (N_1388,N_488,N_670);
nand U1389 (N_1389,N_234,N_684);
xor U1390 (N_1390,N_438,N_117);
nor U1391 (N_1391,N_314,N_529);
nand U1392 (N_1392,N_183,N_323);
nor U1393 (N_1393,N_82,N_594);
nand U1394 (N_1394,N_722,N_307);
nand U1395 (N_1395,N_618,N_147);
nor U1396 (N_1396,N_221,N_347);
nor U1397 (N_1397,N_174,N_612);
or U1398 (N_1398,N_350,N_36);
or U1399 (N_1399,N_246,N_671);
or U1400 (N_1400,N_694,N_718);
and U1401 (N_1401,N_460,N_591);
xnor U1402 (N_1402,N_334,N_430);
or U1403 (N_1403,N_631,N_90);
xor U1404 (N_1404,N_473,N_604);
nand U1405 (N_1405,N_344,N_600);
nor U1406 (N_1406,N_747,N_107);
nand U1407 (N_1407,N_73,N_577);
and U1408 (N_1408,N_135,N_225);
and U1409 (N_1409,N_277,N_593);
nor U1410 (N_1410,N_368,N_124);
nand U1411 (N_1411,N_488,N_16);
and U1412 (N_1412,N_150,N_443);
nand U1413 (N_1413,N_434,N_361);
nand U1414 (N_1414,N_173,N_735);
and U1415 (N_1415,N_213,N_511);
or U1416 (N_1416,N_227,N_65);
nor U1417 (N_1417,N_557,N_479);
and U1418 (N_1418,N_67,N_584);
nand U1419 (N_1419,N_604,N_463);
nor U1420 (N_1420,N_521,N_507);
and U1421 (N_1421,N_737,N_413);
nor U1422 (N_1422,N_261,N_144);
or U1423 (N_1423,N_23,N_440);
and U1424 (N_1424,N_303,N_601);
or U1425 (N_1425,N_284,N_134);
nor U1426 (N_1426,N_259,N_594);
or U1427 (N_1427,N_384,N_520);
nor U1428 (N_1428,N_711,N_657);
or U1429 (N_1429,N_715,N_491);
and U1430 (N_1430,N_302,N_702);
or U1431 (N_1431,N_575,N_423);
nand U1432 (N_1432,N_165,N_331);
nor U1433 (N_1433,N_263,N_374);
or U1434 (N_1434,N_623,N_179);
nand U1435 (N_1435,N_478,N_632);
nor U1436 (N_1436,N_561,N_373);
nor U1437 (N_1437,N_684,N_527);
nand U1438 (N_1438,N_546,N_94);
xor U1439 (N_1439,N_558,N_685);
nand U1440 (N_1440,N_160,N_694);
or U1441 (N_1441,N_225,N_316);
nor U1442 (N_1442,N_79,N_265);
and U1443 (N_1443,N_549,N_472);
nor U1444 (N_1444,N_696,N_331);
and U1445 (N_1445,N_678,N_461);
nor U1446 (N_1446,N_535,N_650);
nand U1447 (N_1447,N_526,N_300);
nor U1448 (N_1448,N_299,N_130);
nor U1449 (N_1449,N_372,N_596);
nor U1450 (N_1450,N_526,N_458);
and U1451 (N_1451,N_9,N_633);
nand U1452 (N_1452,N_624,N_225);
or U1453 (N_1453,N_424,N_737);
and U1454 (N_1454,N_564,N_322);
or U1455 (N_1455,N_631,N_74);
nor U1456 (N_1456,N_344,N_301);
or U1457 (N_1457,N_470,N_601);
and U1458 (N_1458,N_273,N_542);
or U1459 (N_1459,N_75,N_394);
or U1460 (N_1460,N_128,N_677);
xnor U1461 (N_1461,N_483,N_223);
nand U1462 (N_1462,N_111,N_153);
nand U1463 (N_1463,N_575,N_183);
or U1464 (N_1464,N_34,N_91);
nand U1465 (N_1465,N_713,N_626);
or U1466 (N_1466,N_105,N_490);
nand U1467 (N_1467,N_309,N_202);
and U1468 (N_1468,N_330,N_34);
or U1469 (N_1469,N_93,N_212);
nand U1470 (N_1470,N_458,N_398);
and U1471 (N_1471,N_493,N_51);
and U1472 (N_1472,N_355,N_574);
and U1473 (N_1473,N_289,N_575);
or U1474 (N_1474,N_199,N_105);
or U1475 (N_1475,N_94,N_520);
nand U1476 (N_1476,N_343,N_326);
xnor U1477 (N_1477,N_244,N_157);
and U1478 (N_1478,N_75,N_440);
or U1479 (N_1479,N_144,N_286);
and U1480 (N_1480,N_188,N_450);
nand U1481 (N_1481,N_149,N_142);
or U1482 (N_1482,N_205,N_453);
and U1483 (N_1483,N_108,N_17);
nand U1484 (N_1484,N_361,N_9);
and U1485 (N_1485,N_668,N_449);
nor U1486 (N_1486,N_59,N_248);
or U1487 (N_1487,N_225,N_240);
and U1488 (N_1488,N_531,N_269);
nor U1489 (N_1489,N_725,N_734);
nand U1490 (N_1490,N_633,N_291);
xor U1491 (N_1491,N_579,N_62);
or U1492 (N_1492,N_508,N_4);
and U1493 (N_1493,N_380,N_652);
xnor U1494 (N_1494,N_152,N_160);
or U1495 (N_1495,N_55,N_242);
xor U1496 (N_1496,N_434,N_110);
or U1497 (N_1497,N_549,N_685);
nor U1498 (N_1498,N_552,N_608);
nor U1499 (N_1499,N_427,N_318);
nand U1500 (N_1500,N_995,N_1362);
or U1501 (N_1501,N_1369,N_883);
and U1502 (N_1502,N_896,N_1234);
or U1503 (N_1503,N_1038,N_844);
nand U1504 (N_1504,N_1037,N_1498);
nand U1505 (N_1505,N_937,N_1046);
xor U1506 (N_1506,N_822,N_1044);
or U1507 (N_1507,N_841,N_814);
and U1508 (N_1508,N_833,N_942);
nand U1509 (N_1509,N_1226,N_1488);
nor U1510 (N_1510,N_792,N_1131);
and U1511 (N_1511,N_1461,N_754);
nor U1512 (N_1512,N_1349,N_1394);
xor U1513 (N_1513,N_1413,N_1393);
nor U1514 (N_1514,N_1221,N_1055);
or U1515 (N_1515,N_864,N_1476);
nor U1516 (N_1516,N_852,N_1104);
or U1517 (N_1517,N_1162,N_1333);
or U1518 (N_1518,N_1191,N_1199);
and U1519 (N_1519,N_1134,N_1093);
and U1520 (N_1520,N_750,N_1177);
nand U1521 (N_1521,N_970,N_1088);
nand U1522 (N_1522,N_1174,N_897);
nor U1523 (N_1523,N_1278,N_818);
xnor U1524 (N_1524,N_1314,N_1499);
nand U1525 (N_1525,N_755,N_965);
and U1526 (N_1526,N_1357,N_1193);
or U1527 (N_1527,N_1281,N_945);
or U1528 (N_1528,N_1245,N_1015);
nand U1529 (N_1529,N_1183,N_858);
and U1530 (N_1530,N_1027,N_1477);
or U1531 (N_1531,N_1255,N_1095);
or U1532 (N_1532,N_1067,N_1051);
xor U1533 (N_1533,N_943,N_1277);
nand U1534 (N_1534,N_1425,N_1090);
or U1535 (N_1535,N_875,N_1448);
and U1536 (N_1536,N_1423,N_1118);
or U1537 (N_1537,N_1462,N_1220);
and U1538 (N_1538,N_1382,N_1227);
nor U1539 (N_1539,N_1170,N_1132);
nand U1540 (N_1540,N_950,N_913);
nor U1541 (N_1541,N_920,N_805);
nor U1542 (N_1542,N_1092,N_1456);
or U1543 (N_1543,N_879,N_892);
nor U1544 (N_1544,N_1381,N_1209);
nand U1545 (N_1545,N_932,N_803);
nor U1546 (N_1546,N_981,N_1474);
nand U1547 (N_1547,N_850,N_1304);
or U1548 (N_1548,N_802,N_772);
and U1549 (N_1549,N_1271,N_1124);
or U1550 (N_1550,N_1250,N_762);
xor U1551 (N_1551,N_900,N_1270);
or U1552 (N_1552,N_1068,N_1383);
nand U1553 (N_1553,N_1291,N_1453);
nor U1554 (N_1554,N_1181,N_1378);
or U1555 (N_1555,N_992,N_1190);
nand U1556 (N_1556,N_1103,N_1350);
and U1557 (N_1557,N_829,N_1328);
nor U1558 (N_1558,N_1036,N_1115);
and U1559 (N_1559,N_966,N_1003);
nand U1560 (N_1560,N_1323,N_1424);
nand U1561 (N_1561,N_813,N_1265);
or U1562 (N_1562,N_935,N_1263);
and U1563 (N_1563,N_1133,N_1089);
nor U1564 (N_1564,N_1111,N_977);
nor U1565 (N_1565,N_866,N_1283);
and U1566 (N_1566,N_972,N_1455);
nor U1567 (N_1567,N_1479,N_1346);
nor U1568 (N_1568,N_1211,N_1406);
nor U1569 (N_1569,N_1481,N_1097);
and U1570 (N_1570,N_946,N_1155);
or U1571 (N_1571,N_1302,N_1184);
nor U1572 (N_1572,N_1450,N_1404);
nor U1573 (N_1573,N_783,N_1315);
or U1574 (N_1574,N_1065,N_765);
nand U1575 (N_1575,N_1402,N_949);
nand U1576 (N_1576,N_1251,N_1126);
nor U1577 (N_1577,N_827,N_1398);
nor U1578 (N_1578,N_1136,N_914);
and U1579 (N_1579,N_839,N_1043);
and U1580 (N_1580,N_1129,N_1492);
or U1581 (N_1581,N_902,N_1142);
or U1582 (N_1582,N_1484,N_1151);
nor U1583 (N_1583,N_1218,N_1224);
or U1584 (N_1584,N_1222,N_905);
and U1585 (N_1585,N_1012,N_1143);
nor U1586 (N_1586,N_1007,N_1475);
nor U1587 (N_1587,N_807,N_1070);
nor U1588 (N_1588,N_1363,N_1483);
nor U1589 (N_1589,N_1201,N_856);
nand U1590 (N_1590,N_1309,N_774);
nand U1591 (N_1591,N_1085,N_921);
nand U1592 (N_1592,N_986,N_782);
nand U1593 (N_1593,N_1496,N_1337);
nand U1594 (N_1594,N_760,N_1082);
nand U1595 (N_1595,N_1495,N_1025);
nand U1596 (N_1596,N_1253,N_978);
and U1597 (N_1597,N_1313,N_793);
nand U1598 (N_1598,N_939,N_1004);
and U1599 (N_1599,N_854,N_1358);
nor U1600 (N_1600,N_1042,N_1083);
and U1601 (N_1601,N_847,N_874);
and U1602 (N_1602,N_1000,N_903);
and U1603 (N_1603,N_759,N_1237);
nor U1604 (N_1604,N_947,N_753);
and U1605 (N_1605,N_778,N_842);
nor U1606 (N_1606,N_893,N_1219);
and U1607 (N_1607,N_1144,N_1138);
nor U1608 (N_1608,N_930,N_1242);
or U1609 (N_1609,N_1268,N_846);
or U1610 (N_1610,N_961,N_979);
nor U1611 (N_1611,N_859,N_1331);
xor U1612 (N_1612,N_787,N_1367);
or U1613 (N_1613,N_1141,N_764);
nor U1614 (N_1614,N_1169,N_1340);
nor U1615 (N_1615,N_1139,N_1230);
xor U1616 (N_1616,N_1079,N_835);
or U1617 (N_1617,N_1254,N_1303);
or U1618 (N_1618,N_1342,N_1194);
xor U1619 (N_1619,N_938,N_1391);
nand U1620 (N_1620,N_904,N_1011);
nand U1621 (N_1621,N_1354,N_997);
nor U1622 (N_1622,N_1440,N_1119);
nor U1623 (N_1623,N_1166,N_1215);
and U1624 (N_1624,N_887,N_809);
nand U1625 (N_1625,N_928,N_1117);
nand U1626 (N_1626,N_1076,N_819);
nand U1627 (N_1627,N_1021,N_1260);
nand U1628 (N_1628,N_779,N_1062);
or U1629 (N_1629,N_1001,N_1100);
nand U1630 (N_1630,N_1348,N_1473);
or U1631 (N_1631,N_1186,N_1063);
or U1632 (N_1632,N_797,N_1470);
and U1633 (N_1633,N_990,N_1344);
nand U1634 (N_1634,N_1157,N_1310);
or U1635 (N_1635,N_828,N_1457);
or U1636 (N_1636,N_1325,N_1293);
and U1637 (N_1637,N_812,N_1438);
and U1638 (N_1638,N_964,N_926);
and U1639 (N_1639,N_911,N_1212);
and U1640 (N_1640,N_1324,N_1326);
nand U1641 (N_1641,N_777,N_843);
xnor U1642 (N_1642,N_1236,N_1057);
nand U1643 (N_1643,N_1454,N_873);
nor U1644 (N_1644,N_810,N_830);
nand U1645 (N_1645,N_857,N_967);
or U1646 (N_1646,N_1204,N_1202);
or U1647 (N_1647,N_1074,N_1319);
nand U1648 (N_1648,N_1116,N_1264);
nor U1649 (N_1649,N_1013,N_1494);
and U1650 (N_1650,N_1307,N_1207);
and U1651 (N_1651,N_862,N_1441);
and U1652 (N_1652,N_757,N_971);
and U1653 (N_1653,N_1109,N_840);
nor U1654 (N_1654,N_951,N_878);
nand U1655 (N_1655,N_1374,N_1073);
and U1656 (N_1656,N_1429,N_1182);
nand U1657 (N_1657,N_1485,N_871);
nor U1658 (N_1658,N_955,N_789);
or U1659 (N_1659,N_1463,N_1322);
nand U1660 (N_1660,N_1343,N_1298);
and U1661 (N_1661,N_953,N_1120);
or U1662 (N_1662,N_1016,N_1443);
nand U1663 (N_1663,N_1329,N_1290);
or U1664 (N_1664,N_1014,N_1414);
nand U1665 (N_1665,N_1266,N_1239);
or U1666 (N_1666,N_1377,N_1153);
or U1667 (N_1667,N_791,N_1370);
nor U1668 (N_1668,N_1468,N_1179);
or U1669 (N_1669,N_838,N_1206);
and U1670 (N_1670,N_1029,N_1299);
and U1671 (N_1671,N_1053,N_957);
nor U1672 (N_1672,N_1289,N_918);
or U1673 (N_1673,N_795,N_1469);
nor U1674 (N_1674,N_924,N_1318);
xor U1675 (N_1675,N_882,N_1482);
nor U1676 (N_1676,N_1122,N_1105);
and U1677 (N_1677,N_927,N_816);
and U1678 (N_1678,N_999,N_1336);
and U1679 (N_1679,N_1433,N_1335);
nor U1680 (N_1680,N_1189,N_1276);
nand U1681 (N_1681,N_1114,N_794);
xor U1682 (N_1682,N_1026,N_948);
and U1683 (N_1683,N_1019,N_1345);
nor U1684 (N_1684,N_788,N_1075);
nor U1685 (N_1685,N_1285,N_989);
nand U1686 (N_1686,N_1368,N_767);
and U1687 (N_1687,N_984,N_910);
and U1688 (N_1688,N_936,N_1228);
or U1689 (N_1689,N_888,N_1421);
and U1690 (N_1690,N_1172,N_1410);
nor U1691 (N_1691,N_959,N_1408);
xor U1692 (N_1692,N_1020,N_1041);
nor U1693 (N_1693,N_1415,N_1113);
or U1694 (N_1694,N_899,N_1417);
nand U1695 (N_1695,N_867,N_1320);
nor U1696 (N_1696,N_1176,N_1168);
and U1697 (N_1697,N_832,N_1486);
nor U1698 (N_1698,N_1446,N_923);
nand U1699 (N_1699,N_1034,N_1274);
xnor U1700 (N_1700,N_801,N_863);
and U1701 (N_1701,N_820,N_1431);
nor U1702 (N_1702,N_1102,N_1223);
or U1703 (N_1703,N_1360,N_1040);
and U1704 (N_1704,N_898,N_1497);
xor U1705 (N_1705,N_1301,N_808);
nand U1706 (N_1706,N_1148,N_941);
and U1707 (N_1707,N_1405,N_1389);
or U1708 (N_1708,N_1399,N_1030);
nor U1709 (N_1709,N_1444,N_1208);
nand U1710 (N_1710,N_1422,N_1039);
or U1711 (N_1711,N_1478,N_1247);
and U1712 (N_1712,N_1379,N_1359);
and U1713 (N_1713,N_916,N_996);
xor U1714 (N_1714,N_1447,N_1248);
or U1715 (N_1715,N_1490,N_868);
nor U1716 (N_1716,N_1292,N_1244);
nor U1717 (N_1717,N_1022,N_853);
nand U1718 (N_1718,N_1366,N_1355);
or U1719 (N_1719,N_1099,N_790);
or U1720 (N_1720,N_761,N_1137);
or U1721 (N_1721,N_962,N_889);
and U1722 (N_1722,N_885,N_1235);
nor U1723 (N_1723,N_1297,N_952);
and U1724 (N_1724,N_1371,N_1054);
nor U1725 (N_1725,N_991,N_1198);
nor U1726 (N_1726,N_1436,N_1430);
or U1727 (N_1727,N_1480,N_1146);
nand U1728 (N_1728,N_1069,N_786);
nor U1729 (N_1729,N_870,N_1262);
or U1730 (N_1730,N_1300,N_1364);
nand U1731 (N_1731,N_976,N_994);
xor U1732 (N_1732,N_1311,N_1471);
or U1733 (N_1733,N_985,N_1066);
nor U1734 (N_1734,N_933,N_1240);
nand U1735 (N_1735,N_1491,N_1380);
nor U1736 (N_1736,N_1225,N_929);
or U1737 (N_1737,N_825,N_1449);
nand U1738 (N_1738,N_1229,N_1295);
nor U1739 (N_1739,N_1238,N_1197);
and U1740 (N_1740,N_998,N_1002);
and U1741 (N_1741,N_1330,N_974);
and U1742 (N_1742,N_1390,N_1192);
and U1743 (N_1743,N_1164,N_799);
and U1744 (N_1744,N_1023,N_1098);
or U1745 (N_1745,N_969,N_1493);
or U1746 (N_1746,N_1005,N_1384);
nand U1747 (N_1747,N_1200,N_1256);
xnor U1748 (N_1748,N_1130,N_1280);
and U1749 (N_1749,N_1288,N_1165);
nand U1750 (N_1750,N_826,N_1006);
xor U1751 (N_1751,N_785,N_1187);
nand U1752 (N_1752,N_1284,N_1401);
or U1753 (N_1753,N_1231,N_1261);
and U1754 (N_1754,N_1108,N_1150);
and U1755 (N_1755,N_1059,N_1306);
nand U1756 (N_1756,N_1467,N_1465);
or U1757 (N_1757,N_960,N_891);
nor U1758 (N_1758,N_1356,N_1178);
or U1759 (N_1759,N_1395,N_983);
nor U1760 (N_1760,N_1434,N_954);
nand U1761 (N_1761,N_848,N_845);
and U1762 (N_1762,N_1052,N_925);
and U1763 (N_1763,N_1312,N_815);
or U1764 (N_1764,N_876,N_980);
or U1765 (N_1765,N_1418,N_849);
or U1766 (N_1766,N_1460,N_1035);
or U1767 (N_1767,N_1338,N_1411);
or U1768 (N_1768,N_1152,N_1110);
or U1769 (N_1769,N_1400,N_1028);
and U1770 (N_1770,N_1321,N_1196);
or U1771 (N_1771,N_758,N_1442);
nand U1772 (N_1772,N_781,N_1388);
nor U1773 (N_1773,N_1428,N_1259);
nor U1774 (N_1774,N_1216,N_917);
nand U1775 (N_1775,N_1050,N_804);
and U1776 (N_1776,N_973,N_1106);
nor U1777 (N_1777,N_1112,N_988);
xnor U1778 (N_1778,N_1128,N_1086);
or U1779 (N_1779,N_1249,N_1275);
nor U1780 (N_1780,N_1332,N_1272);
or U1781 (N_1781,N_1412,N_1175);
and U1782 (N_1782,N_1024,N_880);
and U1783 (N_1783,N_1018,N_1094);
nand U1784 (N_1784,N_1416,N_1246);
nand U1785 (N_1785,N_1396,N_1386);
nor U1786 (N_1786,N_823,N_1140);
nor U1787 (N_1787,N_1159,N_1397);
nand U1788 (N_1788,N_940,N_1171);
xor U1789 (N_1789,N_1173,N_1084);
and U1790 (N_1790,N_1048,N_1031);
and U1791 (N_1791,N_1273,N_1352);
nand U1792 (N_1792,N_837,N_1373);
xnor U1793 (N_1793,N_1279,N_907);
or U1794 (N_1794,N_836,N_1049);
nor U1795 (N_1795,N_975,N_1147);
nand U1796 (N_1796,N_1101,N_1213);
or U1797 (N_1797,N_1233,N_1437);
and U1798 (N_1798,N_958,N_1252);
xnor U1799 (N_1799,N_922,N_1161);
nor U1800 (N_1800,N_1008,N_1472);
or U1801 (N_1801,N_1464,N_1107);
and U1802 (N_1802,N_1217,N_1033);
or U1803 (N_1803,N_773,N_1045);
nand U1804 (N_1804,N_901,N_1214);
and U1805 (N_1805,N_1351,N_798);
nand U1806 (N_1806,N_780,N_915);
or U1807 (N_1807,N_1387,N_1096);
nor U1808 (N_1808,N_1432,N_1409);
nand U1809 (N_1809,N_811,N_963);
or U1810 (N_1810,N_824,N_1267);
or U1811 (N_1811,N_1009,N_751);
nand U1812 (N_1812,N_1010,N_834);
or U1813 (N_1813,N_1087,N_769);
nor U1814 (N_1814,N_1426,N_1294);
nor U1815 (N_1815,N_968,N_763);
or U1816 (N_1816,N_1353,N_776);
and U1817 (N_1817,N_1375,N_1257);
nand U1818 (N_1818,N_1160,N_756);
and U1819 (N_1819,N_1056,N_1071);
nand U1820 (N_1820,N_1339,N_1205);
nor U1821 (N_1821,N_1149,N_1407);
nor U1822 (N_1822,N_861,N_1458);
nor U1823 (N_1823,N_1282,N_1403);
nor U1824 (N_1824,N_1317,N_895);
and U1825 (N_1825,N_1195,N_1081);
and U1826 (N_1826,N_1185,N_855);
nand U1827 (N_1827,N_1145,N_1072);
nand U1828 (N_1828,N_1210,N_931);
and U1829 (N_1829,N_784,N_1180);
nand U1830 (N_1830,N_831,N_1420);
nor U1831 (N_1831,N_1188,N_1167);
or U1832 (N_1832,N_1017,N_806);
nand U1833 (N_1833,N_768,N_1080);
nand U1834 (N_1834,N_817,N_1316);
nor U1835 (N_1835,N_1376,N_1287);
nor U1836 (N_1836,N_1060,N_1156);
nand U1837 (N_1837,N_851,N_860);
and U1838 (N_1838,N_993,N_1451);
nor U1839 (N_1839,N_1452,N_1327);
and U1840 (N_1840,N_1121,N_1361);
nand U1841 (N_1841,N_1296,N_1385);
nor U1842 (N_1842,N_1078,N_1158);
and U1843 (N_1843,N_1154,N_1419);
nand U1844 (N_1844,N_909,N_770);
nor U1845 (N_1845,N_1308,N_1286);
nor U1846 (N_1846,N_1258,N_771);
or U1847 (N_1847,N_1163,N_1372);
or U1848 (N_1848,N_1232,N_796);
nand U1849 (N_1849,N_934,N_919);
or U1850 (N_1850,N_886,N_877);
or U1851 (N_1851,N_766,N_1047);
or U1852 (N_1852,N_1064,N_1466);
nand U1853 (N_1853,N_800,N_1341);
or U1854 (N_1854,N_908,N_1445);
nor U1855 (N_1855,N_956,N_1241);
nand U1856 (N_1856,N_872,N_1123);
nand U1857 (N_1857,N_1032,N_1334);
or U1858 (N_1858,N_1127,N_1489);
nand U1859 (N_1859,N_1487,N_1077);
or U1860 (N_1860,N_1459,N_1061);
or U1861 (N_1861,N_906,N_890);
nand U1862 (N_1862,N_1091,N_982);
and U1863 (N_1863,N_1243,N_894);
nor U1864 (N_1864,N_869,N_1439);
and U1865 (N_1865,N_1203,N_881);
xor U1866 (N_1866,N_1135,N_752);
or U1867 (N_1867,N_987,N_1427);
and U1868 (N_1868,N_884,N_865);
nor U1869 (N_1869,N_1269,N_821);
nor U1870 (N_1870,N_1392,N_1305);
nor U1871 (N_1871,N_1435,N_944);
and U1872 (N_1872,N_1125,N_1058);
nand U1873 (N_1873,N_1365,N_912);
nand U1874 (N_1874,N_1347,N_775);
and U1875 (N_1875,N_1397,N_809);
and U1876 (N_1876,N_1468,N_938);
xnor U1877 (N_1877,N_1357,N_981);
nand U1878 (N_1878,N_1359,N_1308);
nor U1879 (N_1879,N_1401,N_943);
and U1880 (N_1880,N_940,N_912);
and U1881 (N_1881,N_914,N_1294);
nor U1882 (N_1882,N_1406,N_1338);
and U1883 (N_1883,N_840,N_843);
and U1884 (N_1884,N_979,N_874);
nand U1885 (N_1885,N_908,N_1311);
or U1886 (N_1886,N_1325,N_1362);
or U1887 (N_1887,N_1162,N_892);
nand U1888 (N_1888,N_1065,N_1079);
xor U1889 (N_1889,N_809,N_795);
nand U1890 (N_1890,N_837,N_1310);
or U1891 (N_1891,N_914,N_1388);
nor U1892 (N_1892,N_968,N_1091);
and U1893 (N_1893,N_1133,N_1048);
or U1894 (N_1894,N_938,N_1301);
nand U1895 (N_1895,N_909,N_1308);
or U1896 (N_1896,N_1046,N_1272);
xnor U1897 (N_1897,N_1110,N_998);
nor U1898 (N_1898,N_1113,N_986);
and U1899 (N_1899,N_977,N_812);
and U1900 (N_1900,N_1218,N_1206);
and U1901 (N_1901,N_927,N_1103);
and U1902 (N_1902,N_773,N_1020);
and U1903 (N_1903,N_1178,N_1030);
or U1904 (N_1904,N_1339,N_1455);
nor U1905 (N_1905,N_1115,N_1341);
or U1906 (N_1906,N_866,N_1386);
nand U1907 (N_1907,N_1123,N_1298);
nor U1908 (N_1908,N_1387,N_878);
and U1909 (N_1909,N_1293,N_944);
nor U1910 (N_1910,N_1464,N_1050);
and U1911 (N_1911,N_1333,N_770);
or U1912 (N_1912,N_1025,N_1004);
or U1913 (N_1913,N_1288,N_1089);
nand U1914 (N_1914,N_993,N_1438);
nor U1915 (N_1915,N_1209,N_1058);
nand U1916 (N_1916,N_1051,N_1409);
or U1917 (N_1917,N_1011,N_1206);
nand U1918 (N_1918,N_1131,N_1227);
nand U1919 (N_1919,N_1171,N_1357);
nor U1920 (N_1920,N_824,N_855);
and U1921 (N_1921,N_767,N_1224);
and U1922 (N_1922,N_784,N_1277);
nor U1923 (N_1923,N_1264,N_795);
and U1924 (N_1924,N_842,N_1188);
and U1925 (N_1925,N_830,N_922);
or U1926 (N_1926,N_1242,N_765);
nand U1927 (N_1927,N_1476,N_1081);
and U1928 (N_1928,N_1276,N_808);
nand U1929 (N_1929,N_787,N_1249);
nand U1930 (N_1930,N_1375,N_1167);
nor U1931 (N_1931,N_1036,N_902);
nor U1932 (N_1932,N_1236,N_1197);
nor U1933 (N_1933,N_986,N_1114);
nor U1934 (N_1934,N_1040,N_1106);
xnor U1935 (N_1935,N_1462,N_1036);
nand U1936 (N_1936,N_756,N_1371);
nand U1937 (N_1937,N_869,N_1065);
nand U1938 (N_1938,N_824,N_1277);
nor U1939 (N_1939,N_907,N_1353);
nor U1940 (N_1940,N_1268,N_1235);
and U1941 (N_1941,N_960,N_1499);
and U1942 (N_1942,N_753,N_761);
nand U1943 (N_1943,N_859,N_822);
nor U1944 (N_1944,N_1348,N_1303);
and U1945 (N_1945,N_972,N_1360);
and U1946 (N_1946,N_1384,N_836);
nand U1947 (N_1947,N_863,N_1032);
and U1948 (N_1948,N_901,N_1177);
xnor U1949 (N_1949,N_927,N_1433);
nor U1950 (N_1950,N_1382,N_925);
nand U1951 (N_1951,N_1169,N_816);
nand U1952 (N_1952,N_1191,N_1412);
nand U1953 (N_1953,N_1317,N_1034);
nor U1954 (N_1954,N_932,N_1177);
and U1955 (N_1955,N_976,N_758);
nand U1956 (N_1956,N_965,N_1158);
nor U1957 (N_1957,N_805,N_839);
or U1958 (N_1958,N_1395,N_1394);
nor U1959 (N_1959,N_952,N_860);
nand U1960 (N_1960,N_1255,N_1272);
nand U1961 (N_1961,N_853,N_1333);
or U1962 (N_1962,N_1141,N_963);
nor U1963 (N_1963,N_1173,N_1148);
and U1964 (N_1964,N_936,N_1298);
or U1965 (N_1965,N_1328,N_1329);
nor U1966 (N_1966,N_1365,N_1485);
nand U1967 (N_1967,N_1177,N_1068);
and U1968 (N_1968,N_1160,N_966);
xnor U1969 (N_1969,N_801,N_1104);
nor U1970 (N_1970,N_943,N_1485);
and U1971 (N_1971,N_1413,N_1249);
and U1972 (N_1972,N_862,N_1165);
and U1973 (N_1973,N_846,N_1028);
and U1974 (N_1974,N_956,N_1150);
or U1975 (N_1975,N_1489,N_816);
nor U1976 (N_1976,N_1312,N_750);
and U1977 (N_1977,N_1221,N_1083);
nand U1978 (N_1978,N_1342,N_1390);
nand U1979 (N_1979,N_1230,N_1278);
or U1980 (N_1980,N_1371,N_1215);
and U1981 (N_1981,N_933,N_968);
nor U1982 (N_1982,N_1342,N_1325);
or U1983 (N_1983,N_809,N_1470);
nand U1984 (N_1984,N_1414,N_1338);
and U1985 (N_1985,N_1033,N_998);
nand U1986 (N_1986,N_1332,N_771);
nor U1987 (N_1987,N_1038,N_1448);
nor U1988 (N_1988,N_1430,N_1247);
nand U1989 (N_1989,N_1257,N_1488);
nor U1990 (N_1990,N_1259,N_1169);
nor U1991 (N_1991,N_1360,N_1184);
xnor U1992 (N_1992,N_1121,N_1349);
nor U1993 (N_1993,N_769,N_891);
nor U1994 (N_1994,N_847,N_1244);
xor U1995 (N_1995,N_1124,N_759);
and U1996 (N_1996,N_1390,N_1446);
nand U1997 (N_1997,N_1051,N_1027);
nor U1998 (N_1998,N_1141,N_1304);
nand U1999 (N_1999,N_949,N_977);
nor U2000 (N_2000,N_1054,N_1005);
nand U2001 (N_2001,N_1330,N_1315);
nand U2002 (N_2002,N_1027,N_1498);
nand U2003 (N_2003,N_1271,N_962);
nand U2004 (N_2004,N_1197,N_758);
or U2005 (N_2005,N_1027,N_1138);
nor U2006 (N_2006,N_830,N_844);
nor U2007 (N_2007,N_1393,N_1005);
nand U2008 (N_2008,N_842,N_969);
nor U2009 (N_2009,N_1314,N_986);
nand U2010 (N_2010,N_859,N_1086);
xnor U2011 (N_2011,N_1378,N_1001);
or U2012 (N_2012,N_1182,N_1261);
nor U2013 (N_2013,N_1012,N_772);
and U2014 (N_2014,N_1179,N_950);
and U2015 (N_2015,N_789,N_1159);
nand U2016 (N_2016,N_1382,N_1137);
nor U2017 (N_2017,N_777,N_1047);
nand U2018 (N_2018,N_1006,N_1428);
nor U2019 (N_2019,N_1388,N_1030);
nor U2020 (N_2020,N_1227,N_1100);
xor U2021 (N_2021,N_1259,N_915);
nand U2022 (N_2022,N_1487,N_1033);
and U2023 (N_2023,N_1289,N_1308);
nor U2024 (N_2024,N_1499,N_1172);
or U2025 (N_2025,N_1266,N_1463);
nand U2026 (N_2026,N_1012,N_1052);
nand U2027 (N_2027,N_1176,N_1140);
nand U2028 (N_2028,N_1118,N_1414);
and U2029 (N_2029,N_1387,N_1038);
or U2030 (N_2030,N_1042,N_892);
nor U2031 (N_2031,N_1383,N_1081);
nor U2032 (N_2032,N_1438,N_1433);
nand U2033 (N_2033,N_1477,N_991);
nor U2034 (N_2034,N_1247,N_1018);
or U2035 (N_2035,N_1282,N_1350);
xor U2036 (N_2036,N_943,N_836);
and U2037 (N_2037,N_1183,N_880);
or U2038 (N_2038,N_1134,N_876);
and U2039 (N_2039,N_1466,N_1220);
or U2040 (N_2040,N_925,N_1354);
or U2041 (N_2041,N_1368,N_1122);
xnor U2042 (N_2042,N_1422,N_1167);
nand U2043 (N_2043,N_1395,N_962);
or U2044 (N_2044,N_1399,N_1031);
nand U2045 (N_2045,N_1366,N_965);
nor U2046 (N_2046,N_795,N_899);
xnor U2047 (N_2047,N_1473,N_1057);
xor U2048 (N_2048,N_774,N_1476);
or U2049 (N_2049,N_1028,N_930);
and U2050 (N_2050,N_918,N_795);
nand U2051 (N_2051,N_1238,N_1236);
xor U2052 (N_2052,N_1034,N_1396);
and U2053 (N_2053,N_807,N_1378);
xor U2054 (N_2054,N_1379,N_1204);
nor U2055 (N_2055,N_1468,N_1378);
and U2056 (N_2056,N_1226,N_892);
or U2057 (N_2057,N_1411,N_784);
nor U2058 (N_2058,N_860,N_1353);
nor U2059 (N_2059,N_1429,N_1318);
nand U2060 (N_2060,N_1017,N_1310);
nand U2061 (N_2061,N_819,N_763);
and U2062 (N_2062,N_918,N_1043);
and U2063 (N_2063,N_901,N_763);
nand U2064 (N_2064,N_799,N_956);
xnor U2065 (N_2065,N_1061,N_997);
or U2066 (N_2066,N_1110,N_765);
and U2067 (N_2067,N_1063,N_950);
and U2068 (N_2068,N_1126,N_1177);
or U2069 (N_2069,N_1080,N_1254);
nand U2070 (N_2070,N_1437,N_1293);
and U2071 (N_2071,N_1015,N_892);
and U2072 (N_2072,N_1379,N_1355);
xor U2073 (N_2073,N_1062,N_1043);
or U2074 (N_2074,N_1182,N_1234);
or U2075 (N_2075,N_1490,N_1147);
nor U2076 (N_2076,N_1474,N_826);
nand U2077 (N_2077,N_888,N_768);
xnor U2078 (N_2078,N_1378,N_1267);
or U2079 (N_2079,N_1317,N_1069);
nand U2080 (N_2080,N_1004,N_759);
nor U2081 (N_2081,N_798,N_1056);
and U2082 (N_2082,N_999,N_1435);
or U2083 (N_2083,N_1106,N_1239);
or U2084 (N_2084,N_1300,N_900);
nor U2085 (N_2085,N_897,N_836);
and U2086 (N_2086,N_1099,N_1158);
or U2087 (N_2087,N_1210,N_1378);
and U2088 (N_2088,N_1465,N_1270);
nor U2089 (N_2089,N_920,N_921);
and U2090 (N_2090,N_846,N_1177);
xor U2091 (N_2091,N_1149,N_1405);
nor U2092 (N_2092,N_1498,N_1135);
or U2093 (N_2093,N_982,N_1345);
and U2094 (N_2094,N_1410,N_1158);
and U2095 (N_2095,N_978,N_1187);
and U2096 (N_2096,N_788,N_1428);
and U2097 (N_2097,N_1023,N_869);
and U2098 (N_2098,N_1114,N_1170);
nor U2099 (N_2099,N_1241,N_1082);
nor U2100 (N_2100,N_1221,N_1235);
nor U2101 (N_2101,N_1205,N_1132);
nand U2102 (N_2102,N_803,N_1279);
and U2103 (N_2103,N_1081,N_1013);
or U2104 (N_2104,N_788,N_982);
and U2105 (N_2105,N_1469,N_813);
nor U2106 (N_2106,N_812,N_1354);
or U2107 (N_2107,N_899,N_928);
or U2108 (N_2108,N_1249,N_1273);
nand U2109 (N_2109,N_1258,N_991);
or U2110 (N_2110,N_1451,N_773);
and U2111 (N_2111,N_1243,N_861);
nand U2112 (N_2112,N_807,N_1011);
and U2113 (N_2113,N_1346,N_1058);
nand U2114 (N_2114,N_773,N_905);
xor U2115 (N_2115,N_940,N_1397);
nor U2116 (N_2116,N_1045,N_1357);
nor U2117 (N_2117,N_1353,N_1303);
nand U2118 (N_2118,N_999,N_1349);
nand U2119 (N_2119,N_1180,N_1007);
nor U2120 (N_2120,N_1238,N_1015);
nor U2121 (N_2121,N_1124,N_883);
nor U2122 (N_2122,N_1176,N_1255);
nor U2123 (N_2123,N_783,N_1268);
nand U2124 (N_2124,N_836,N_1416);
nand U2125 (N_2125,N_926,N_1432);
and U2126 (N_2126,N_1023,N_1437);
nor U2127 (N_2127,N_1323,N_903);
or U2128 (N_2128,N_870,N_756);
nor U2129 (N_2129,N_1125,N_949);
xor U2130 (N_2130,N_1178,N_928);
and U2131 (N_2131,N_1423,N_842);
nor U2132 (N_2132,N_964,N_1470);
xor U2133 (N_2133,N_1458,N_894);
and U2134 (N_2134,N_1024,N_870);
and U2135 (N_2135,N_786,N_1148);
nor U2136 (N_2136,N_915,N_1222);
or U2137 (N_2137,N_1174,N_876);
or U2138 (N_2138,N_1288,N_977);
nor U2139 (N_2139,N_1217,N_753);
xor U2140 (N_2140,N_1270,N_1238);
nor U2141 (N_2141,N_1155,N_1194);
nor U2142 (N_2142,N_1292,N_1388);
and U2143 (N_2143,N_950,N_1351);
nand U2144 (N_2144,N_1113,N_1015);
xor U2145 (N_2145,N_805,N_924);
and U2146 (N_2146,N_837,N_828);
or U2147 (N_2147,N_1109,N_942);
nand U2148 (N_2148,N_1046,N_922);
nand U2149 (N_2149,N_790,N_1330);
nand U2150 (N_2150,N_1192,N_1331);
and U2151 (N_2151,N_931,N_772);
or U2152 (N_2152,N_919,N_936);
or U2153 (N_2153,N_1070,N_751);
nor U2154 (N_2154,N_1208,N_1234);
nor U2155 (N_2155,N_964,N_1060);
or U2156 (N_2156,N_1289,N_1451);
or U2157 (N_2157,N_1245,N_1155);
xnor U2158 (N_2158,N_1013,N_845);
and U2159 (N_2159,N_1389,N_861);
and U2160 (N_2160,N_1293,N_1121);
and U2161 (N_2161,N_1036,N_917);
and U2162 (N_2162,N_1093,N_1137);
nor U2163 (N_2163,N_898,N_764);
nand U2164 (N_2164,N_941,N_1159);
or U2165 (N_2165,N_1354,N_1476);
nand U2166 (N_2166,N_1452,N_1111);
or U2167 (N_2167,N_836,N_818);
and U2168 (N_2168,N_1363,N_1466);
nor U2169 (N_2169,N_768,N_1369);
nand U2170 (N_2170,N_828,N_1452);
nand U2171 (N_2171,N_1136,N_1323);
or U2172 (N_2172,N_1449,N_1350);
and U2173 (N_2173,N_1067,N_1397);
nand U2174 (N_2174,N_948,N_767);
nand U2175 (N_2175,N_901,N_754);
nand U2176 (N_2176,N_1301,N_1272);
and U2177 (N_2177,N_1437,N_753);
and U2178 (N_2178,N_918,N_1422);
nor U2179 (N_2179,N_1019,N_1319);
nor U2180 (N_2180,N_1184,N_1424);
nor U2181 (N_2181,N_761,N_1238);
or U2182 (N_2182,N_1156,N_1262);
nor U2183 (N_2183,N_844,N_1493);
nand U2184 (N_2184,N_1270,N_1257);
or U2185 (N_2185,N_1169,N_1358);
nand U2186 (N_2186,N_964,N_1293);
nand U2187 (N_2187,N_1234,N_952);
or U2188 (N_2188,N_1219,N_1202);
nor U2189 (N_2189,N_1476,N_989);
xnor U2190 (N_2190,N_797,N_1283);
nand U2191 (N_2191,N_875,N_1066);
nand U2192 (N_2192,N_810,N_1176);
nand U2193 (N_2193,N_924,N_1118);
or U2194 (N_2194,N_775,N_1076);
and U2195 (N_2195,N_803,N_943);
nor U2196 (N_2196,N_814,N_986);
or U2197 (N_2197,N_1255,N_1172);
nand U2198 (N_2198,N_1381,N_1383);
and U2199 (N_2199,N_780,N_1452);
xor U2200 (N_2200,N_1217,N_1400);
nor U2201 (N_2201,N_1085,N_1235);
nand U2202 (N_2202,N_1421,N_1267);
nor U2203 (N_2203,N_1414,N_781);
and U2204 (N_2204,N_1406,N_888);
nand U2205 (N_2205,N_1443,N_1232);
xor U2206 (N_2206,N_983,N_1159);
nor U2207 (N_2207,N_976,N_1227);
xnor U2208 (N_2208,N_1276,N_1120);
or U2209 (N_2209,N_1359,N_1468);
xnor U2210 (N_2210,N_997,N_991);
or U2211 (N_2211,N_1476,N_1179);
nor U2212 (N_2212,N_937,N_933);
or U2213 (N_2213,N_914,N_1210);
and U2214 (N_2214,N_820,N_1025);
or U2215 (N_2215,N_1153,N_1103);
and U2216 (N_2216,N_1002,N_778);
nor U2217 (N_2217,N_1381,N_1028);
nor U2218 (N_2218,N_873,N_1085);
and U2219 (N_2219,N_1074,N_1444);
nand U2220 (N_2220,N_924,N_1319);
nor U2221 (N_2221,N_1031,N_1182);
and U2222 (N_2222,N_889,N_1102);
or U2223 (N_2223,N_1218,N_874);
and U2224 (N_2224,N_1391,N_1162);
nor U2225 (N_2225,N_1384,N_928);
and U2226 (N_2226,N_1182,N_1357);
nand U2227 (N_2227,N_887,N_831);
nor U2228 (N_2228,N_1099,N_771);
nor U2229 (N_2229,N_1379,N_890);
or U2230 (N_2230,N_782,N_866);
nor U2231 (N_2231,N_1044,N_918);
or U2232 (N_2232,N_1289,N_1182);
and U2233 (N_2233,N_1243,N_1021);
and U2234 (N_2234,N_834,N_1499);
nand U2235 (N_2235,N_801,N_1403);
nand U2236 (N_2236,N_954,N_1360);
nor U2237 (N_2237,N_896,N_948);
nand U2238 (N_2238,N_1365,N_756);
nand U2239 (N_2239,N_1284,N_902);
nor U2240 (N_2240,N_923,N_803);
nand U2241 (N_2241,N_942,N_1345);
nor U2242 (N_2242,N_948,N_799);
and U2243 (N_2243,N_887,N_1039);
nor U2244 (N_2244,N_932,N_773);
or U2245 (N_2245,N_1214,N_971);
or U2246 (N_2246,N_1170,N_1217);
and U2247 (N_2247,N_1159,N_1237);
or U2248 (N_2248,N_1197,N_1252);
nand U2249 (N_2249,N_1163,N_1475);
nor U2250 (N_2250,N_1940,N_1976);
or U2251 (N_2251,N_1729,N_2028);
or U2252 (N_2252,N_2126,N_1581);
nand U2253 (N_2253,N_2240,N_2065);
xor U2254 (N_2254,N_1832,N_1840);
nor U2255 (N_2255,N_2022,N_1901);
nor U2256 (N_2256,N_1596,N_1509);
and U2257 (N_2257,N_2169,N_1859);
or U2258 (N_2258,N_2044,N_2093);
or U2259 (N_2259,N_2220,N_1970);
and U2260 (N_2260,N_1728,N_1689);
nand U2261 (N_2261,N_1672,N_1784);
xnor U2262 (N_2262,N_1587,N_1772);
and U2263 (N_2263,N_1933,N_1585);
and U2264 (N_2264,N_1968,N_1530);
xor U2265 (N_2265,N_2109,N_1516);
and U2266 (N_2266,N_2144,N_1872);
or U2267 (N_2267,N_1814,N_2108);
xnor U2268 (N_2268,N_1868,N_1550);
and U2269 (N_2269,N_2066,N_1654);
nor U2270 (N_2270,N_2225,N_1870);
nor U2271 (N_2271,N_1992,N_1644);
xnor U2272 (N_2272,N_1572,N_2201);
or U2273 (N_2273,N_2016,N_2143);
and U2274 (N_2274,N_1950,N_1759);
or U2275 (N_2275,N_1993,N_1515);
or U2276 (N_2276,N_1565,N_1836);
nand U2277 (N_2277,N_1892,N_1916);
xor U2278 (N_2278,N_1605,N_2026);
nand U2279 (N_2279,N_1563,N_2202);
or U2280 (N_2280,N_1567,N_1623);
nor U2281 (N_2281,N_1982,N_2161);
or U2282 (N_2282,N_1747,N_1591);
nand U2283 (N_2283,N_1527,N_1812);
xor U2284 (N_2284,N_1726,N_1925);
nand U2285 (N_2285,N_1560,N_2042);
or U2286 (N_2286,N_2122,N_2062);
or U2287 (N_2287,N_1830,N_1883);
nand U2288 (N_2288,N_1896,N_1756);
nand U2289 (N_2289,N_1642,N_1721);
nand U2290 (N_2290,N_1730,N_1743);
nor U2291 (N_2291,N_2103,N_2189);
nand U2292 (N_2292,N_1790,N_1540);
and U2293 (N_2293,N_2014,N_1939);
nor U2294 (N_2294,N_2068,N_1874);
and U2295 (N_2295,N_2205,N_1804);
nor U2296 (N_2296,N_1904,N_2153);
and U2297 (N_2297,N_1808,N_1504);
nor U2298 (N_2298,N_1974,N_2160);
or U2299 (N_2299,N_1511,N_1879);
nand U2300 (N_2300,N_2056,N_1652);
xor U2301 (N_2301,N_2011,N_1785);
nand U2302 (N_2302,N_2097,N_2137);
nand U2303 (N_2303,N_2000,N_1782);
and U2304 (N_2304,N_1696,N_2190);
nor U2305 (N_2305,N_1589,N_1526);
and U2306 (N_2306,N_1675,N_2147);
and U2307 (N_2307,N_1841,N_2218);
or U2308 (N_2308,N_2083,N_2239);
nand U2309 (N_2309,N_1690,N_1746);
and U2310 (N_2310,N_2032,N_2158);
nor U2311 (N_2311,N_1778,N_2178);
nor U2312 (N_2312,N_2074,N_1910);
nand U2313 (N_2313,N_1574,N_2193);
xnor U2314 (N_2314,N_2211,N_1914);
nand U2315 (N_2315,N_2245,N_1903);
and U2316 (N_2316,N_1599,N_1691);
or U2317 (N_2317,N_1665,N_2199);
and U2318 (N_2318,N_2145,N_2033);
or U2319 (N_2319,N_1650,N_1763);
nor U2320 (N_2320,N_2157,N_1631);
or U2321 (N_2321,N_1533,N_2174);
nand U2322 (N_2322,N_2210,N_1881);
and U2323 (N_2323,N_1717,N_1789);
and U2324 (N_2324,N_1984,N_1573);
and U2325 (N_2325,N_2249,N_1986);
xor U2326 (N_2326,N_2094,N_1657);
nand U2327 (N_2327,N_1532,N_1518);
nand U2328 (N_2328,N_1542,N_1851);
nor U2329 (N_2329,N_2204,N_1658);
or U2330 (N_2330,N_1956,N_1577);
nand U2331 (N_2331,N_2163,N_2060);
and U2332 (N_2332,N_1547,N_1924);
xnor U2333 (N_2333,N_2127,N_1655);
or U2334 (N_2334,N_2077,N_1604);
and U2335 (N_2335,N_1523,N_1628);
or U2336 (N_2336,N_2188,N_1568);
nor U2337 (N_2337,N_1662,N_2013);
nand U2338 (N_2338,N_1683,N_2207);
nor U2339 (N_2339,N_1781,N_1713);
and U2340 (N_2340,N_2168,N_1794);
and U2341 (N_2341,N_1783,N_1816);
or U2342 (N_2342,N_2246,N_1704);
and U2343 (N_2343,N_1770,N_1624);
nand U2344 (N_2344,N_2002,N_1674);
nor U2345 (N_2345,N_2140,N_1556);
nand U2346 (N_2346,N_1699,N_1817);
or U2347 (N_2347,N_1752,N_2006);
nor U2348 (N_2348,N_1811,N_2206);
or U2349 (N_2349,N_1776,N_2233);
xor U2350 (N_2350,N_1813,N_2047);
nand U2351 (N_2351,N_1935,N_2175);
nor U2352 (N_2352,N_2131,N_1918);
xnor U2353 (N_2353,N_2012,N_1797);
nor U2354 (N_2354,N_2120,N_2133);
xnor U2355 (N_2355,N_2228,N_1519);
and U2356 (N_2356,N_2155,N_1963);
or U2357 (N_2357,N_2197,N_1942);
and U2358 (N_2358,N_1653,N_1952);
nor U2359 (N_2359,N_2184,N_1663);
xnor U2360 (N_2360,N_1768,N_1825);
nand U2361 (N_2361,N_1948,N_1849);
nor U2362 (N_2362,N_2100,N_2194);
and U2363 (N_2363,N_1700,N_2209);
and U2364 (N_2364,N_1844,N_1975);
nor U2365 (N_2365,N_1994,N_2113);
and U2366 (N_2366,N_1678,N_2118);
nand U2367 (N_2367,N_1562,N_1549);
xor U2368 (N_2368,N_2067,N_1638);
xor U2369 (N_2369,N_1671,N_1514);
or U2370 (N_2370,N_1936,N_2090);
and U2371 (N_2371,N_1934,N_1848);
nor U2372 (N_2372,N_2111,N_1866);
or U2373 (N_2373,N_1983,N_2151);
and U2374 (N_2374,N_1688,N_1742);
or U2375 (N_2375,N_2009,N_1648);
nor U2376 (N_2376,N_1679,N_1737);
and U2377 (N_2377,N_1753,N_2167);
or U2378 (N_2378,N_1601,N_2064);
and U2379 (N_2379,N_1660,N_1805);
xnor U2380 (N_2380,N_1593,N_2052);
and U2381 (N_2381,N_1769,N_2173);
nor U2382 (N_2382,N_1643,N_1787);
nor U2383 (N_2383,N_1641,N_1684);
and U2384 (N_2384,N_2171,N_1981);
or U2385 (N_2385,N_1588,N_1877);
nand U2386 (N_2386,N_1831,N_2055);
nand U2387 (N_2387,N_1922,N_1850);
or U2388 (N_2388,N_1796,N_1720);
xnor U2389 (N_2389,N_1754,N_2136);
xnor U2390 (N_2390,N_1537,N_2244);
and U2391 (N_2391,N_1508,N_1579);
nor U2392 (N_2392,N_2248,N_2095);
and U2393 (N_2393,N_2148,N_1615);
and U2394 (N_2394,N_2196,N_1923);
xnor U2395 (N_2395,N_1538,N_1580);
or U2396 (N_2396,N_1535,N_1553);
nor U2397 (N_2397,N_2092,N_2079);
nand U2398 (N_2398,N_1863,N_1960);
nand U2399 (N_2399,N_1749,N_1893);
nand U2400 (N_2400,N_1930,N_1978);
nor U2401 (N_2401,N_2063,N_2085);
and U2402 (N_2402,N_1712,N_2236);
or U2403 (N_2403,N_1570,N_1685);
nand U2404 (N_2404,N_1997,N_2101);
or U2405 (N_2405,N_1627,N_1810);
nand U2406 (N_2406,N_1899,N_1894);
nor U2407 (N_2407,N_2213,N_1854);
nor U2408 (N_2408,N_1611,N_1987);
or U2409 (N_2409,N_1898,N_1736);
xnor U2410 (N_2410,N_2142,N_2183);
nor U2411 (N_2411,N_1632,N_1773);
and U2412 (N_2412,N_1502,N_1600);
and U2413 (N_2413,N_2010,N_1900);
and U2414 (N_2414,N_1711,N_2080);
xnor U2415 (N_2415,N_1965,N_1792);
nand U2416 (N_2416,N_2082,N_2152);
nand U2417 (N_2417,N_2180,N_2069);
and U2418 (N_2418,N_2200,N_1998);
nor U2419 (N_2419,N_1815,N_2115);
or U2420 (N_2420,N_2104,N_1732);
xor U2421 (N_2421,N_1517,N_1907);
and U2422 (N_2422,N_1501,N_2051);
nor U2423 (N_2423,N_1858,N_1528);
nor U2424 (N_2424,N_1833,N_1557);
nand U2425 (N_2425,N_1838,N_1764);
nand U2426 (N_2426,N_2223,N_1546);
or U2427 (N_2427,N_2027,N_2238);
or U2428 (N_2428,N_2048,N_2181);
xor U2429 (N_2429,N_1578,N_1758);
nor U2430 (N_2430,N_1937,N_1788);
nor U2431 (N_2431,N_1766,N_1677);
nor U2432 (N_2432,N_1719,N_1902);
and U2433 (N_2433,N_1731,N_1767);
or U2434 (N_2434,N_1503,N_1548);
and U2435 (N_2435,N_1541,N_1964);
and U2436 (N_2436,N_1739,N_2224);
nor U2437 (N_2437,N_1839,N_1705);
nor U2438 (N_2438,N_2035,N_2138);
xnor U2439 (N_2439,N_1897,N_1919);
nor U2440 (N_2440,N_2182,N_1908);
and U2441 (N_2441,N_1861,N_1694);
nand U2442 (N_2442,N_1536,N_1584);
or U2443 (N_2443,N_2231,N_2017);
and U2444 (N_2444,N_1626,N_1799);
nand U2445 (N_2445,N_1703,N_1669);
nand U2446 (N_2446,N_2030,N_1980);
nand U2447 (N_2447,N_1500,N_2081);
and U2448 (N_2448,N_2162,N_1826);
or U2449 (N_2449,N_1807,N_1822);
or U2450 (N_2450,N_1595,N_2075);
xor U2451 (N_2451,N_2215,N_1608);
and U2452 (N_2452,N_1798,N_2191);
or U2453 (N_2453,N_1820,N_1966);
nor U2454 (N_2454,N_1661,N_1864);
nand U2455 (N_2455,N_1727,N_2088);
and U2456 (N_2456,N_2154,N_1941);
nand U2457 (N_2457,N_2005,N_1692);
nor U2458 (N_2458,N_1534,N_2020);
nand U2459 (N_2459,N_1707,N_1915);
nor U2460 (N_2460,N_2237,N_1771);
nor U2461 (N_2461,N_2135,N_1630);
or U2462 (N_2462,N_1979,N_1803);
nor U2463 (N_2463,N_1929,N_1603);
xor U2464 (N_2464,N_1529,N_1640);
or U2465 (N_2465,N_1621,N_1738);
nand U2466 (N_2466,N_1955,N_1846);
nor U2467 (N_2467,N_2123,N_2185);
and U2468 (N_2468,N_1828,N_1716);
or U2469 (N_2469,N_1639,N_2221);
xor U2470 (N_2470,N_2124,N_1522);
nor U2471 (N_2471,N_1668,N_1651);
nand U2472 (N_2472,N_1757,N_2156);
nor U2473 (N_2473,N_1913,N_1607);
nor U2474 (N_2474,N_1635,N_2177);
nand U2475 (N_2475,N_1748,N_1741);
and U2476 (N_2476,N_1912,N_2216);
nor U2477 (N_2477,N_2139,N_1552);
nand U2478 (N_2478,N_2089,N_1701);
and U2479 (N_2479,N_2214,N_2203);
nor U2480 (N_2480,N_1762,N_1634);
nor U2481 (N_2481,N_2078,N_2102);
nor U2482 (N_2482,N_2070,N_2179);
nand U2483 (N_2483,N_1853,N_1876);
or U2484 (N_2484,N_2242,N_1760);
nand U2485 (N_2485,N_1506,N_2247);
nand U2486 (N_2486,N_1967,N_2038);
xnor U2487 (N_2487,N_2105,N_2061);
nor U2488 (N_2488,N_1800,N_2125);
nor U2489 (N_2489,N_1745,N_2050);
nor U2490 (N_2490,N_1695,N_1680);
nand U2491 (N_2491,N_1895,N_1735);
or U2492 (N_2492,N_1761,N_2187);
nor U2493 (N_2493,N_1878,N_1666);
nand U2494 (N_2494,N_1602,N_1687);
nand U2495 (N_2495,N_2008,N_1718);
nand U2496 (N_2496,N_1946,N_2018);
nor U2497 (N_2497,N_1673,N_2235);
and U2498 (N_2498,N_1555,N_1885);
xor U2499 (N_2499,N_1860,N_1613);
nand U2500 (N_2500,N_2087,N_1834);
nor U2501 (N_2501,N_1583,N_2037);
or U2502 (N_2502,N_1667,N_1962);
nor U2503 (N_2503,N_2071,N_2058);
nand U2504 (N_2504,N_1709,N_2043);
nor U2505 (N_2505,N_1809,N_1697);
nor U2506 (N_2506,N_2036,N_2001);
nor U2507 (N_2507,N_1586,N_1610);
xor U2508 (N_2508,N_1744,N_1681);
and U2509 (N_2509,N_1750,N_2129);
nand U2510 (N_2510,N_1888,N_1999);
xnor U2511 (N_2511,N_1510,N_1958);
nand U2512 (N_2512,N_2166,N_1592);
or U2513 (N_2513,N_1647,N_1646);
and U2514 (N_2514,N_1953,N_2031);
or U2515 (N_2515,N_1645,N_1633);
or U2516 (N_2516,N_1724,N_1911);
and U2517 (N_2517,N_1777,N_1943);
nor U2518 (N_2518,N_2024,N_1676);
xnor U2519 (N_2519,N_2116,N_2243);
or U2520 (N_2520,N_1710,N_1722);
and U2521 (N_2521,N_1835,N_2096);
xor U2522 (N_2522,N_1544,N_1917);
or U2523 (N_2523,N_1875,N_1909);
nand U2524 (N_2524,N_1606,N_1715);
or U2525 (N_2525,N_1755,N_1571);
nor U2526 (N_2526,N_1886,N_1521);
and U2527 (N_2527,N_1921,N_1871);
or U2528 (N_2528,N_1906,N_1884);
or U2529 (N_2529,N_1597,N_2112);
and U2530 (N_2530,N_1590,N_1801);
nor U2531 (N_2531,N_2107,N_1829);
or U2532 (N_2532,N_1734,N_2106);
xnor U2533 (N_2533,N_1845,N_2040);
and U2534 (N_2534,N_2119,N_1971);
nor U2535 (N_2535,N_1554,N_1622);
nor U2536 (N_2536,N_1616,N_1867);
and U2537 (N_2537,N_1905,N_2046);
nor U2538 (N_2538,N_1629,N_2114);
or U2539 (N_2539,N_2186,N_1618);
or U2540 (N_2540,N_1954,N_2054);
and U2541 (N_2541,N_1889,N_1786);
or U2542 (N_2542,N_1869,N_2176);
nand U2543 (N_2543,N_1543,N_1791);
xor U2544 (N_2544,N_2076,N_1664);
xnor U2545 (N_2545,N_2023,N_1512);
nor U2546 (N_2546,N_1949,N_2086);
and U2547 (N_2547,N_2084,N_1857);
nor U2548 (N_2548,N_1614,N_1823);
or U2549 (N_2549,N_1852,N_2049);
and U2550 (N_2550,N_2019,N_1847);
nand U2551 (N_2551,N_2004,N_1531);
or U2552 (N_2552,N_1751,N_1887);
nand U2553 (N_2553,N_2021,N_1670);
nand U2554 (N_2554,N_1972,N_1880);
or U2555 (N_2555,N_1843,N_2025);
xnor U2556 (N_2556,N_1926,N_2232);
nor U2557 (N_2557,N_1539,N_1821);
or U2558 (N_2558,N_2091,N_1649);
xor U2559 (N_2559,N_1873,N_1865);
nor U2560 (N_2560,N_1569,N_1636);
xor U2561 (N_2561,N_2029,N_1686);
nand U2562 (N_2562,N_1545,N_1637);
xor U2563 (N_2563,N_2241,N_1990);
nor U2564 (N_2564,N_1780,N_1582);
nor U2565 (N_2565,N_1513,N_1617);
and U2566 (N_2566,N_2146,N_1708);
nand U2567 (N_2567,N_2121,N_1698);
nand U2568 (N_2568,N_2212,N_1507);
nand U2569 (N_2569,N_2164,N_1988);
nor U2570 (N_2570,N_1505,N_2222);
nor U2571 (N_2571,N_1945,N_1920);
nand U2572 (N_2572,N_1733,N_1927);
nor U2573 (N_2573,N_1938,N_1779);
xor U2574 (N_2574,N_1706,N_2098);
nor U2575 (N_2575,N_2219,N_1564);
nand U2576 (N_2576,N_2226,N_1806);
and U2577 (N_2577,N_1625,N_1969);
or U2578 (N_2578,N_1693,N_1559);
nand U2579 (N_2579,N_1891,N_2217);
nor U2580 (N_2580,N_2130,N_1520);
nor U2581 (N_2581,N_2132,N_1656);
nand U2582 (N_2582,N_1932,N_1795);
and U2583 (N_2583,N_2141,N_2057);
or U2584 (N_2584,N_1802,N_2099);
or U2585 (N_2585,N_1827,N_1793);
nor U2586 (N_2586,N_2059,N_1837);
nand U2587 (N_2587,N_2159,N_2227);
and U2588 (N_2588,N_2117,N_1819);
nor U2589 (N_2589,N_2165,N_2007);
or U2590 (N_2590,N_1575,N_1775);
or U2591 (N_2591,N_2149,N_1774);
nor U2592 (N_2592,N_2003,N_1524);
nand U2593 (N_2593,N_2150,N_1944);
nand U2594 (N_2594,N_1566,N_1598);
nand U2595 (N_2595,N_1765,N_2072);
or U2596 (N_2596,N_1856,N_1612);
nand U2597 (N_2597,N_1824,N_1702);
or U2598 (N_2598,N_1957,N_1973);
nor U2599 (N_2599,N_2034,N_2134);
nand U2600 (N_2600,N_1842,N_1558);
and U2601 (N_2601,N_1928,N_2234);
nor U2602 (N_2602,N_2195,N_2041);
nand U2603 (N_2603,N_1961,N_1740);
nand U2604 (N_2604,N_2073,N_2208);
and U2605 (N_2605,N_1855,N_2230);
or U2606 (N_2606,N_1561,N_1609);
and U2607 (N_2607,N_2192,N_1620);
and U2608 (N_2608,N_2198,N_1989);
nand U2609 (N_2609,N_1723,N_1951);
xor U2610 (N_2610,N_1576,N_1682);
nor U2611 (N_2611,N_1882,N_2229);
or U2612 (N_2612,N_1991,N_1977);
nor U2613 (N_2613,N_1594,N_1862);
nor U2614 (N_2614,N_2039,N_1818);
xor U2615 (N_2615,N_1551,N_1959);
and U2616 (N_2616,N_2045,N_1995);
or U2617 (N_2617,N_1725,N_1996);
nand U2618 (N_2618,N_2015,N_1931);
nor U2619 (N_2619,N_1619,N_2172);
or U2620 (N_2620,N_2128,N_1985);
or U2621 (N_2621,N_2170,N_1947);
xnor U2622 (N_2622,N_2110,N_1659);
nor U2623 (N_2623,N_1890,N_2053);
and U2624 (N_2624,N_1714,N_1525);
nor U2625 (N_2625,N_1986,N_1916);
xor U2626 (N_2626,N_2001,N_2035);
nand U2627 (N_2627,N_2119,N_2105);
nor U2628 (N_2628,N_2224,N_2062);
or U2629 (N_2629,N_1736,N_1826);
and U2630 (N_2630,N_2220,N_1647);
or U2631 (N_2631,N_2098,N_2069);
or U2632 (N_2632,N_1722,N_2033);
nand U2633 (N_2633,N_2139,N_1921);
and U2634 (N_2634,N_1550,N_2159);
nand U2635 (N_2635,N_2002,N_1778);
and U2636 (N_2636,N_1552,N_1598);
and U2637 (N_2637,N_2011,N_1987);
and U2638 (N_2638,N_1612,N_2166);
nand U2639 (N_2639,N_2213,N_1827);
nor U2640 (N_2640,N_1526,N_1752);
xor U2641 (N_2641,N_1893,N_1712);
or U2642 (N_2642,N_2211,N_1832);
nand U2643 (N_2643,N_1731,N_2104);
and U2644 (N_2644,N_1647,N_2149);
and U2645 (N_2645,N_2246,N_2012);
or U2646 (N_2646,N_2202,N_2095);
or U2647 (N_2647,N_1732,N_2167);
and U2648 (N_2648,N_1862,N_1890);
or U2649 (N_2649,N_2115,N_1557);
nor U2650 (N_2650,N_1901,N_1744);
nand U2651 (N_2651,N_1600,N_1764);
nor U2652 (N_2652,N_1863,N_1516);
nor U2653 (N_2653,N_1654,N_1996);
or U2654 (N_2654,N_2027,N_1511);
xor U2655 (N_2655,N_2134,N_2190);
or U2656 (N_2656,N_2099,N_1996);
nor U2657 (N_2657,N_1947,N_1916);
nor U2658 (N_2658,N_1703,N_1570);
nand U2659 (N_2659,N_1983,N_2133);
or U2660 (N_2660,N_2238,N_1762);
or U2661 (N_2661,N_1611,N_2063);
or U2662 (N_2662,N_1559,N_2221);
nor U2663 (N_2663,N_1808,N_1839);
xor U2664 (N_2664,N_2154,N_1884);
and U2665 (N_2665,N_2021,N_2220);
or U2666 (N_2666,N_1965,N_2211);
and U2667 (N_2667,N_2034,N_1941);
nor U2668 (N_2668,N_1940,N_2166);
xor U2669 (N_2669,N_1539,N_2060);
nand U2670 (N_2670,N_1535,N_1752);
and U2671 (N_2671,N_1905,N_2089);
nor U2672 (N_2672,N_1747,N_2170);
or U2673 (N_2673,N_1995,N_1582);
nor U2674 (N_2674,N_1552,N_1926);
or U2675 (N_2675,N_2117,N_1991);
and U2676 (N_2676,N_1571,N_1795);
or U2677 (N_2677,N_1967,N_1860);
nor U2678 (N_2678,N_1690,N_1942);
nand U2679 (N_2679,N_1629,N_2050);
or U2680 (N_2680,N_2158,N_1969);
nand U2681 (N_2681,N_1728,N_1536);
and U2682 (N_2682,N_1872,N_1619);
nand U2683 (N_2683,N_1947,N_1951);
or U2684 (N_2684,N_2199,N_2166);
or U2685 (N_2685,N_2148,N_1895);
nor U2686 (N_2686,N_2193,N_1826);
nand U2687 (N_2687,N_2046,N_2217);
nand U2688 (N_2688,N_1984,N_2011);
or U2689 (N_2689,N_1848,N_1744);
xor U2690 (N_2690,N_1889,N_2237);
xor U2691 (N_2691,N_2195,N_1899);
nor U2692 (N_2692,N_2164,N_1831);
xor U2693 (N_2693,N_1941,N_2017);
or U2694 (N_2694,N_1616,N_1668);
nor U2695 (N_2695,N_1760,N_1771);
nand U2696 (N_2696,N_1947,N_1866);
nor U2697 (N_2697,N_2126,N_1764);
or U2698 (N_2698,N_1752,N_1620);
xor U2699 (N_2699,N_1634,N_1837);
or U2700 (N_2700,N_2086,N_1546);
nand U2701 (N_2701,N_2077,N_2101);
nor U2702 (N_2702,N_1545,N_2197);
nand U2703 (N_2703,N_2038,N_1748);
and U2704 (N_2704,N_1932,N_1756);
or U2705 (N_2705,N_1697,N_1851);
xor U2706 (N_2706,N_2194,N_2169);
nand U2707 (N_2707,N_1913,N_1835);
xnor U2708 (N_2708,N_2031,N_1934);
nand U2709 (N_2709,N_2029,N_1956);
nor U2710 (N_2710,N_2177,N_1821);
and U2711 (N_2711,N_2047,N_2173);
nand U2712 (N_2712,N_2200,N_1680);
or U2713 (N_2713,N_1741,N_1674);
nand U2714 (N_2714,N_1709,N_1500);
nor U2715 (N_2715,N_2150,N_1928);
nor U2716 (N_2716,N_1525,N_2093);
or U2717 (N_2717,N_2148,N_1996);
and U2718 (N_2718,N_1944,N_2091);
or U2719 (N_2719,N_1828,N_2113);
or U2720 (N_2720,N_1868,N_2191);
and U2721 (N_2721,N_2057,N_1903);
xor U2722 (N_2722,N_1994,N_1675);
or U2723 (N_2723,N_2013,N_1764);
nand U2724 (N_2724,N_2206,N_1552);
and U2725 (N_2725,N_2211,N_2145);
or U2726 (N_2726,N_1881,N_1997);
or U2727 (N_2727,N_2144,N_1512);
nor U2728 (N_2728,N_2014,N_1878);
nand U2729 (N_2729,N_2238,N_1536);
and U2730 (N_2730,N_1569,N_2045);
nor U2731 (N_2731,N_1788,N_1844);
or U2732 (N_2732,N_1607,N_1579);
nor U2733 (N_2733,N_1617,N_1571);
nand U2734 (N_2734,N_2076,N_1788);
nor U2735 (N_2735,N_1625,N_1566);
xor U2736 (N_2736,N_1660,N_1749);
nor U2737 (N_2737,N_1527,N_1802);
and U2738 (N_2738,N_2171,N_1953);
xnor U2739 (N_2739,N_1596,N_2115);
and U2740 (N_2740,N_2030,N_1595);
nand U2741 (N_2741,N_1520,N_1978);
and U2742 (N_2742,N_2198,N_1591);
nor U2743 (N_2743,N_1678,N_2164);
or U2744 (N_2744,N_1655,N_1989);
nand U2745 (N_2745,N_1993,N_1613);
or U2746 (N_2746,N_2052,N_1928);
or U2747 (N_2747,N_1516,N_1710);
nand U2748 (N_2748,N_1713,N_1529);
and U2749 (N_2749,N_2239,N_1521);
nand U2750 (N_2750,N_2095,N_1532);
nor U2751 (N_2751,N_1742,N_2139);
xnor U2752 (N_2752,N_1938,N_2107);
or U2753 (N_2753,N_1880,N_1613);
nor U2754 (N_2754,N_1556,N_1777);
nor U2755 (N_2755,N_1900,N_1545);
or U2756 (N_2756,N_1779,N_1791);
and U2757 (N_2757,N_1733,N_2038);
nor U2758 (N_2758,N_1781,N_2235);
or U2759 (N_2759,N_2017,N_1856);
and U2760 (N_2760,N_1655,N_1845);
nand U2761 (N_2761,N_1932,N_1821);
and U2762 (N_2762,N_1952,N_1979);
nor U2763 (N_2763,N_2020,N_1853);
nand U2764 (N_2764,N_1881,N_2191);
and U2765 (N_2765,N_2150,N_2032);
and U2766 (N_2766,N_1637,N_1729);
nor U2767 (N_2767,N_1887,N_2082);
and U2768 (N_2768,N_1892,N_2190);
nand U2769 (N_2769,N_1569,N_1724);
nor U2770 (N_2770,N_1737,N_2194);
or U2771 (N_2771,N_2095,N_1765);
or U2772 (N_2772,N_1843,N_1846);
nand U2773 (N_2773,N_2048,N_1761);
nor U2774 (N_2774,N_1791,N_1733);
nor U2775 (N_2775,N_1643,N_1741);
or U2776 (N_2776,N_1593,N_2197);
nor U2777 (N_2777,N_2188,N_2108);
and U2778 (N_2778,N_1620,N_1814);
xnor U2779 (N_2779,N_2162,N_1955);
and U2780 (N_2780,N_1613,N_1733);
or U2781 (N_2781,N_1859,N_1901);
and U2782 (N_2782,N_1792,N_1555);
xor U2783 (N_2783,N_1665,N_1961);
nor U2784 (N_2784,N_1562,N_2114);
or U2785 (N_2785,N_1779,N_1824);
nand U2786 (N_2786,N_1685,N_2209);
or U2787 (N_2787,N_1909,N_1623);
or U2788 (N_2788,N_1758,N_1741);
and U2789 (N_2789,N_1807,N_1561);
or U2790 (N_2790,N_2237,N_2070);
or U2791 (N_2791,N_1697,N_1649);
nor U2792 (N_2792,N_1620,N_2045);
or U2793 (N_2793,N_1832,N_2168);
nand U2794 (N_2794,N_2099,N_2240);
nor U2795 (N_2795,N_2004,N_2075);
nand U2796 (N_2796,N_1684,N_2225);
nand U2797 (N_2797,N_1605,N_1602);
and U2798 (N_2798,N_1553,N_1509);
nor U2799 (N_2799,N_2052,N_1634);
xor U2800 (N_2800,N_2204,N_2052);
or U2801 (N_2801,N_1605,N_1693);
nand U2802 (N_2802,N_2103,N_2044);
nor U2803 (N_2803,N_1744,N_1724);
nor U2804 (N_2804,N_1547,N_1692);
and U2805 (N_2805,N_1867,N_1713);
and U2806 (N_2806,N_1616,N_2121);
nand U2807 (N_2807,N_1735,N_1615);
or U2808 (N_2808,N_1694,N_1646);
nor U2809 (N_2809,N_2241,N_1627);
or U2810 (N_2810,N_1943,N_2120);
xnor U2811 (N_2811,N_1733,N_1648);
xor U2812 (N_2812,N_1838,N_1926);
nand U2813 (N_2813,N_1847,N_1630);
xor U2814 (N_2814,N_1757,N_1759);
nor U2815 (N_2815,N_2164,N_1951);
and U2816 (N_2816,N_1898,N_1502);
and U2817 (N_2817,N_2114,N_1616);
or U2818 (N_2818,N_1553,N_1773);
xnor U2819 (N_2819,N_1724,N_1955);
nor U2820 (N_2820,N_2155,N_1718);
and U2821 (N_2821,N_1763,N_2050);
or U2822 (N_2822,N_1527,N_1606);
nor U2823 (N_2823,N_1861,N_1909);
nand U2824 (N_2824,N_1685,N_1730);
xnor U2825 (N_2825,N_2072,N_1669);
or U2826 (N_2826,N_2222,N_1912);
and U2827 (N_2827,N_1588,N_1642);
or U2828 (N_2828,N_1825,N_2082);
nand U2829 (N_2829,N_1518,N_2000);
nor U2830 (N_2830,N_1621,N_1931);
or U2831 (N_2831,N_2176,N_1819);
nor U2832 (N_2832,N_1906,N_2178);
xnor U2833 (N_2833,N_1551,N_2153);
nor U2834 (N_2834,N_1923,N_1737);
xnor U2835 (N_2835,N_1894,N_1699);
or U2836 (N_2836,N_1784,N_1669);
or U2837 (N_2837,N_1692,N_1871);
nor U2838 (N_2838,N_1601,N_1812);
and U2839 (N_2839,N_2067,N_1511);
nand U2840 (N_2840,N_2091,N_1792);
nand U2841 (N_2841,N_2152,N_1758);
nor U2842 (N_2842,N_1875,N_2163);
nor U2843 (N_2843,N_1992,N_1952);
or U2844 (N_2844,N_1641,N_1994);
and U2845 (N_2845,N_1674,N_2226);
or U2846 (N_2846,N_1680,N_1959);
and U2847 (N_2847,N_2060,N_1944);
and U2848 (N_2848,N_1984,N_1718);
nor U2849 (N_2849,N_2118,N_1569);
or U2850 (N_2850,N_1986,N_1974);
xor U2851 (N_2851,N_1989,N_1512);
nand U2852 (N_2852,N_1877,N_1563);
nand U2853 (N_2853,N_1611,N_1766);
nand U2854 (N_2854,N_1535,N_2230);
and U2855 (N_2855,N_1618,N_1717);
nor U2856 (N_2856,N_1683,N_1662);
or U2857 (N_2857,N_1645,N_1913);
nand U2858 (N_2858,N_1742,N_1579);
and U2859 (N_2859,N_1878,N_1982);
and U2860 (N_2860,N_1531,N_1616);
or U2861 (N_2861,N_1513,N_2206);
and U2862 (N_2862,N_1729,N_2071);
and U2863 (N_2863,N_2094,N_2069);
nor U2864 (N_2864,N_1903,N_1695);
xnor U2865 (N_2865,N_1723,N_1631);
nand U2866 (N_2866,N_1777,N_1954);
xnor U2867 (N_2867,N_2144,N_1847);
or U2868 (N_2868,N_1982,N_1730);
xnor U2869 (N_2869,N_1608,N_1547);
nor U2870 (N_2870,N_2123,N_2137);
nor U2871 (N_2871,N_1937,N_1503);
nand U2872 (N_2872,N_1501,N_1874);
nand U2873 (N_2873,N_2005,N_1568);
nand U2874 (N_2874,N_1755,N_2159);
nand U2875 (N_2875,N_2163,N_2173);
and U2876 (N_2876,N_2137,N_2128);
or U2877 (N_2877,N_1894,N_1574);
and U2878 (N_2878,N_1653,N_2010);
and U2879 (N_2879,N_1553,N_1578);
and U2880 (N_2880,N_1535,N_1695);
or U2881 (N_2881,N_2173,N_1934);
nand U2882 (N_2882,N_2137,N_1708);
or U2883 (N_2883,N_1512,N_1896);
nor U2884 (N_2884,N_1909,N_1991);
nand U2885 (N_2885,N_2013,N_1775);
and U2886 (N_2886,N_1990,N_1625);
and U2887 (N_2887,N_1614,N_1603);
nand U2888 (N_2888,N_1963,N_1850);
xnor U2889 (N_2889,N_2184,N_2129);
and U2890 (N_2890,N_1932,N_1586);
nand U2891 (N_2891,N_2005,N_1596);
or U2892 (N_2892,N_1661,N_1741);
and U2893 (N_2893,N_2246,N_1609);
and U2894 (N_2894,N_1987,N_1509);
or U2895 (N_2895,N_1945,N_1541);
nand U2896 (N_2896,N_2134,N_1668);
or U2897 (N_2897,N_1720,N_2050);
or U2898 (N_2898,N_2076,N_1986);
nor U2899 (N_2899,N_1600,N_1627);
nor U2900 (N_2900,N_1656,N_1900);
xor U2901 (N_2901,N_1546,N_2082);
nand U2902 (N_2902,N_1909,N_1970);
nor U2903 (N_2903,N_1792,N_1740);
and U2904 (N_2904,N_2205,N_2081);
nor U2905 (N_2905,N_2041,N_1886);
and U2906 (N_2906,N_1802,N_2114);
xnor U2907 (N_2907,N_1987,N_1912);
or U2908 (N_2908,N_1572,N_2160);
xor U2909 (N_2909,N_1583,N_2140);
and U2910 (N_2910,N_2054,N_1562);
or U2911 (N_2911,N_1894,N_1981);
or U2912 (N_2912,N_2024,N_1592);
and U2913 (N_2913,N_2100,N_2246);
nor U2914 (N_2914,N_2081,N_2249);
nand U2915 (N_2915,N_2149,N_1734);
or U2916 (N_2916,N_2068,N_1814);
or U2917 (N_2917,N_2045,N_1972);
or U2918 (N_2918,N_1743,N_2214);
nand U2919 (N_2919,N_2158,N_2040);
nor U2920 (N_2920,N_2004,N_1707);
nand U2921 (N_2921,N_1815,N_1972);
nand U2922 (N_2922,N_2003,N_2075);
nor U2923 (N_2923,N_1727,N_2083);
nor U2924 (N_2924,N_1987,N_1648);
nor U2925 (N_2925,N_1689,N_1913);
or U2926 (N_2926,N_1913,N_1756);
xor U2927 (N_2927,N_2162,N_1559);
xor U2928 (N_2928,N_1918,N_1837);
and U2929 (N_2929,N_2212,N_2064);
or U2930 (N_2930,N_2091,N_2181);
and U2931 (N_2931,N_2059,N_2004);
nor U2932 (N_2932,N_1661,N_1558);
nand U2933 (N_2933,N_1656,N_2061);
and U2934 (N_2934,N_2075,N_2076);
nor U2935 (N_2935,N_1638,N_1622);
or U2936 (N_2936,N_1736,N_2245);
and U2937 (N_2937,N_1929,N_1752);
nand U2938 (N_2938,N_2235,N_1555);
or U2939 (N_2939,N_2044,N_2030);
nand U2940 (N_2940,N_2057,N_1967);
nor U2941 (N_2941,N_1955,N_1667);
nand U2942 (N_2942,N_2248,N_1722);
and U2943 (N_2943,N_1892,N_1554);
or U2944 (N_2944,N_1741,N_1720);
nor U2945 (N_2945,N_1969,N_2001);
nor U2946 (N_2946,N_1931,N_1542);
nor U2947 (N_2947,N_2130,N_1874);
nand U2948 (N_2948,N_1628,N_1619);
nor U2949 (N_2949,N_2056,N_1960);
and U2950 (N_2950,N_1573,N_1770);
or U2951 (N_2951,N_1538,N_1777);
and U2952 (N_2952,N_1512,N_1639);
or U2953 (N_2953,N_2101,N_1872);
nor U2954 (N_2954,N_2041,N_1980);
and U2955 (N_2955,N_1594,N_1652);
nor U2956 (N_2956,N_1955,N_1840);
or U2957 (N_2957,N_1620,N_1843);
nand U2958 (N_2958,N_2064,N_2189);
and U2959 (N_2959,N_1657,N_1871);
nor U2960 (N_2960,N_2001,N_1607);
or U2961 (N_2961,N_2102,N_2248);
nand U2962 (N_2962,N_1842,N_1930);
nand U2963 (N_2963,N_1823,N_1642);
and U2964 (N_2964,N_1562,N_1935);
and U2965 (N_2965,N_1533,N_1863);
nor U2966 (N_2966,N_1929,N_1841);
xor U2967 (N_2967,N_2183,N_2148);
nand U2968 (N_2968,N_1661,N_1629);
or U2969 (N_2969,N_1974,N_2093);
or U2970 (N_2970,N_2246,N_2177);
or U2971 (N_2971,N_1799,N_2114);
nand U2972 (N_2972,N_1756,N_2040);
and U2973 (N_2973,N_1675,N_1838);
nand U2974 (N_2974,N_1695,N_1561);
and U2975 (N_2975,N_2019,N_1786);
and U2976 (N_2976,N_1563,N_2062);
or U2977 (N_2977,N_1768,N_1530);
nor U2978 (N_2978,N_2222,N_1570);
nor U2979 (N_2979,N_1968,N_1773);
and U2980 (N_2980,N_1526,N_1677);
nor U2981 (N_2981,N_1976,N_1938);
or U2982 (N_2982,N_2212,N_2056);
and U2983 (N_2983,N_2086,N_1968);
nor U2984 (N_2984,N_1827,N_2043);
nor U2985 (N_2985,N_2233,N_1628);
nor U2986 (N_2986,N_1779,N_1792);
nor U2987 (N_2987,N_2017,N_1902);
xnor U2988 (N_2988,N_1631,N_2023);
nand U2989 (N_2989,N_2057,N_1653);
nand U2990 (N_2990,N_1846,N_1690);
nand U2991 (N_2991,N_2033,N_1659);
nand U2992 (N_2992,N_1983,N_1934);
and U2993 (N_2993,N_1726,N_1626);
and U2994 (N_2994,N_1732,N_2186);
nor U2995 (N_2995,N_1854,N_1913);
nand U2996 (N_2996,N_1667,N_2097);
xor U2997 (N_2997,N_1776,N_2037);
and U2998 (N_2998,N_1834,N_2119);
nor U2999 (N_2999,N_2186,N_2225);
nand UO_0 (O_0,N_2918,N_2990);
and UO_1 (O_1,N_2789,N_2259);
and UO_2 (O_2,N_2598,N_2654);
xnor UO_3 (O_3,N_2633,N_2402);
and UO_4 (O_4,N_2413,N_2296);
and UO_5 (O_5,N_2982,N_2279);
nor UO_6 (O_6,N_2362,N_2341);
nor UO_7 (O_7,N_2912,N_2860);
xnor UO_8 (O_8,N_2826,N_2611);
nand UO_9 (O_9,N_2671,N_2426);
xnor UO_10 (O_10,N_2624,N_2457);
nor UO_11 (O_11,N_2439,N_2669);
xnor UO_12 (O_12,N_2460,N_2967);
xor UO_13 (O_13,N_2861,N_2307);
nor UO_14 (O_14,N_2746,N_2272);
or UO_15 (O_15,N_2438,N_2262);
nand UO_16 (O_16,N_2305,N_2779);
xnor UO_17 (O_17,N_2753,N_2549);
nor UO_18 (O_18,N_2672,N_2981);
or UO_19 (O_19,N_2911,N_2588);
nor UO_20 (O_20,N_2530,N_2686);
and UO_21 (O_21,N_2877,N_2468);
nand UO_22 (O_22,N_2936,N_2899);
nand UO_23 (O_23,N_2821,N_2476);
and UO_24 (O_24,N_2784,N_2927);
xnor UO_25 (O_25,N_2776,N_2359);
nand UO_26 (O_26,N_2792,N_2443);
nor UO_27 (O_27,N_2309,N_2519);
nor UO_28 (O_28,N_2794,N_2721);
and UO_29 (O_29,N_2803,N_2915);
and UO_30 (O_30,N_2540,N_2858);
nor UO_31 (O_31,N_2634,N_2348);
nor UO_32 (O_32,N_2594,N_2928);
nor UO_33 (O_33,N_2571,N_2833);
and UO_34 (O_34,N_2284,N_2730);
nand UO_35 (O_35,N_2683,N_2499);
or UO_36 (O_36,N_2707,N_2815);
nor UO_37 (O_37,N_2433,N_2698);
nand UO_38 (O_38,N_2573,N_2289);
and UO_39 (O_39,N_2497,N_2414);
nand UO_40 (O_40,N_2910,N_2609);
nor UO_41 (O_41,N_2649,N_2926);
nor UO_42 (O_42,N_2589,N_2836);
nand UO_43 (O_43,N_2572,N_2435);
nor UO_44 (O_44,N_2665,N_2660);
nand UO_45 (O_45,N_2664,N_2253);
and UO_46 (O_46,N_2908,N_2366);
xor UO_47 (O_47,N_2642,N_2448);
or UO_48 (O_48,N_2632,N_2937);
xnor UO_49 (O_49,N_2989,N_2700);
nand UO_50 (O_50,N_2873,N_2749);
nand UO_51 (O_51,N_2480,N_2430);
nor UO_52 (O_52,N_2478,N_2380);
or UO_53 (O_53,N_2635,N_2825);
or UO_54 (O_54,N_2945,N_2995);
nor UO_55 (O_55,N_2879,N_2627);
and UO_56 (O_56,N_2935,N_2570);
and UO_57 (O_57,N_2616,N_2934);
and UO_58 (O_58,N_2379,N_2451);
nand UO_59 (O_59,N_2333,N_2893);
and UO_60 (O_60,N_2736,N_2703);
or UO_61 (O_61,N_2276,N_2404);
nor UO_62 (O_62,N_2486,N_2331);
nand UO_63 (O_63,N_2613,N_2473);
xor UO_64 (O_64,N_2264,N_2574);
nand UO_65 (O_65,N_2959,N_2623);
xnor UO_66 (O_66,N_2976,N_2285);
and UO_67 (O_67,N_2891,N_2865);
nand UO_68 (O_68,N_2752,N_2733);
nor UO_69 (O_69,N_2410,N_2527);
and UO_70 (O_70,N_2647,N_2428);
nand UO_71 (O_71,N_2687,N_2718);
nor UO_72 (O_72,N_2550,N_2850);
nor UO_73 (O_73,N_2561,N_2351);
nand UO_74 (O_74,N_2846,N_2342);
and UO_75 (O_75,N_2868,N_2339);
nand UO_76 (O_76,N_2273,N_2742);
or UO_77 (O_77,N_2896,N_2626);
xnor UO_78 (O_78,N_2691,N_2267);
and UO_79 (O_79,N_2444,N_2859);
or UO_80 (O_80,N_2492,N_2724);
nand UO_81 (O_81,N_2886,N_2958);
nor UO_82 (O_82,N_2955,N_2900);
nor UO_83 (O_83,N_2324,N_2754);
xor UO_84 (O_84,N_2261,N_2799);
and UO_85 (O_85,N_2881,N_2951);
and UO_86 (O_86,N_2696,N_2648);
or UO_87 (O_87,N_2596,N_2930);
or UO_88 (O_88,N_2628,N_2406);
or UO_89 (O_89,N_2418,N_2904);
or UO_90 (O_90,N_2994,N_2536);
and UO_91 (O_91,N_2838,N_2941);
or UO_92 (O_92,N_2909,N_2310);
nand UO_93 (O_93,N_2767,N_2897);
and UO_94 (O_94,N_2885,N_2498);
and UO_95 (O_95,N_2411,N_2867);
and UO_96 (O_96,N_2993,N_2681);
and UO_97 (O_97,N_2947,N_2306);
nor UO_98 (O_98,N_2374,N_2997);
nand UO_99 (O_99,N_2602,N_2405);
or UO_100 (O_100,N_2349,N_2521);
nand UO_101 (O_101,N_2764,N_2985);
nor UO_102 (O_102,N_2791,N_2999);
nand UO_103 (O_103,N_2270,N_2729);
nand UO_104 (O_104,N_2802,N_2801);
nand UO_105 (O_105,N_2851,N_2652);
or UO_106 (O_106,N_2932,N_2944);
nand UO_107 (O_107,N_2394,N_2517);
or UO_108 (O_108,N_2383,N_2745);
and UO_109 (O_109,N_2644,N_2670);
or UO_110 (O_110,N_2514,N_2946);
nand UO_111 (O_111,N_2352,N_2505);
or UO_112 (O_112,N_2808,N_2544);
nor UO_113 (O_113,N_2576,N_2922);
nor UO_114 (O_114,N_2365,N_2520);
nand UO_115 (O_115,N_2903,N_2988);
and UO_116 (O_116,N_2513,N_2979);
or UO_117 (O_117,N_2710,N_2583);
nand UO_118 (O_118,N_2254,N_2416);
or UO_119 (O_119,N_2436,N_2759);
nor UO_120 (O_120,N_2998,N_2612);
and UO_121 (O_121,N_2577,N_2363);
or UO_122 (O_122,N_2780,N_2692);
and UO_123 (O_123,N_2373,N_2870);
xnor UO_124 (O_124,N_2697,N_2822);
nor UO_125 (O_125,N_2695,N_2823);
or UO_126 (O_126,N_2914,N_2526);
nand UO_127 (O_127,N_2452,N_2318);
nand UO_128 (O_128,N_2839,N_2898);
nor UO_129 (O_129,N_2747,N_2834);
or UO_130 (O_130,N_2630,N_2370);
xor UO_131 (O_131,N_2377,N_2388);
nor UO_132 (O_132,N_2770,N_2312);
nor UO_133 (O_133,N_2292,N_2639);
nand UO_134 (O_134,N_2470,N_2939);
and UO_135 (O_135,N_2678,N_2554);
and UO_136 (O_136,N_2508,N_2471);
or UO_137 (O_137,N_2645,N_2694);
or UO_138 (O_138,N_2711,N_2481);
and UO_139 (O_139,N_2689,N_2328);
nor UO_140 (O_140,N_2828,N_2975);
or UO_141 (O_141,N_2919,N_2293);
and UO_142 (O_142,N_2895,N_2464);
nor UO_143 (O_143,N_2842,N_2288);
and UO_144 (O_144,N_2579,N_2463);
or UO_145 (O_145,N_2804,N_2263);
or UO_146 (O_146,N_2924,N_2638);
nand UO_147 (O_147,N_2523,N_2278);
or UO_148 (O_148,N_2403,N_2774);
nor UO_149 (O_149,N_2814,N_2316);
nand UO_150 (O_150,N_2586,N_2442);
or UO_151 (O_151,N_2763,N_2677);
nand UO_152 (O_152,N_2827,N_2256);
or UO_153 (O_153,N_2938,N_2668);
xnor UO_154 (O_154,N_2992,N_2358);
nand UO_155 (O_155,N_2948,N_2369);
nand UO_156 (O_156,N_2597,N_2676);
and UO_157 (O_157,N_2738,N_2706);
nand UO_158 (O_158,N_2943,N_2542);
and UO_159 (O_159,N_2485,N_2811);
nand UO_160 (O_160,N_2655,N_2384);
nor UO_161 (O_161,N_2489,N_2287);
and UO_162 (O_162,N_2608,N_2674);
and UO_163 (O_163,N_2964,N_2758);
or UO_164 (O_164,N_2841,N_2303);
xor UO_165 (O_165,N_2923,N_2875);
nor UO_166 (O_166,N_2666,N_2420);
or UO_167 (O_167,N_2500,N_2581);
nor UO_168 (O_168,N_2739,N_2277);
xnor UO_169 (O_169,N_2568,N_2472);
xor UO_170 (O_170,N_2831,N_2378);
or UO_171 (O_171,N_2806,N_2429);
or UO_172 (O_172,N_2512,N_2952);
or UO_173 (O_173,N_2344,N_2422);
nor UO_174 (O_174,N_2569,N_2887);
and UO_175 (O_175,N_2357,N_2297);
nand UO_176 (O_176,N_2506,N_2447);
xor UO_177 (O_177,N_2793,N_2356);
and UO_178 (O_178,N_2317,N_2563);
nand UO_179 (O_179,N_2539,N_2493);
or UO_180 (O_180,N_2960,N_2503);
or UO_181 (O_181,N_2962,N_2725);
and UO_182 (O_182,N_2343,N_2321);
nor UO_183 (O_183,N_2268,N_2528);
or UO_184 (O_184,N_2606,N_2490);
nand UO_185 (O_185,N_2713,N_2580);
nor UO_186 (O_186,N_2902,N_2425);
and UO_187 (O_187,N_2322,N_2364);
nor UO_188 (O_188,N_2501,N_2640);
or UO_189 (O_189,N_2869,N_2590);
and UO_190 (O_190,N_2332,N_2354);
nor UO_191 (O_191,N_2345,N_2385);
nand UO_192 (O_192,N_2876,N_2762);
xor UO_193 (O_193,N_2607,N_2323);
and UO_194 (O_194,N_2441,N_2734);
nand UO_195 (O_195,N_2302,N_2797);
or UO_196 (O_196,N_2788,N_2996);
xor UO_197 (O_197,N_2856,N_2889);
xor UO_198 (O_198,N_2313,N_2529);
nand UO_199 (O_199,N_2916,N_2751);
nor UO_200 (O_200,N_2266,N_2461);
nand UO_201 (O_201,N_2401,N_2469);
nand UO_202 (O_202,N_2818,N_2775);
nor UO_203 (O_203,N_2685,N_2809);
nand UO_204 (O_204,N_2798,N_2755);
nand UO_205 (O_205,N_2740,N_2761);
nor UO_206 (O_206,N_2984,N_2545);
nand UO_207 (O_207,N_2737,N_2773);
nand UO_208 (O_208,N_2882,N_2320);
or UO_209 (O_209,N_2969,N_2769);
xor UO_210 (O_210,N_2682,N_2983);
or UO_211 (O_211,N_2625,N_2294);
xnor UO_212 (O_212,N_2963,N_2731);
or UO_213 (O_213,N_2595,N_2974);
and UO_214 (O_214,N_2462,N_2314);
or UO_215 (O_215,N_2547,N_2601);
and UO_216 (O_216,N_2980,N_2515);
nor UO_217 (O_217,N_2949,N_2705);
nand UO_218 (O_218,N_2866,N_2853);
and UO_219 (O_219,N_2389,N_2884);
and UO_220 (O_220,N_2399,N_2744);
nand UO_221 (O_221,N_2525,N_2835);
xor UO_222 (O_222,N_2484,N_2355);
nor UO_223 (O_223,N_2662,N_2699);
nand UO_224 (O_224,N_2496,N_2494);
or UO_225 (O_225,N_2467,N_2587);
nand UO_226 (O_226,N_2298,N_2466);
nor UO_227 (O_227,N_2653,N_2453);
xnor UO_228 (O_228,N_2986,N_2620);
or UO_229 (O_229,N_2518,N_2714);
or UO_230 (O_230,N_2338,N_2712);
or UO_231 (O_231,N_2874,N_2781);
nand UO_232 (O_232,N_2325,N_2719);
or UO_233 (O_233,N_2757,N_2704);
or UO_234 (O_234,N_2778,N_2409);
and UO_235 (O_235,N_2311,N_2748);
nor UO_236 (O_236,N_2847,N_2970);
nand UO_237 (O_237,N_2631,N_2621);
nand UO_238 (O_238,N_2575,N_2387);
nand UO_239 (O_239,N_2925,N_2812);
or UO_240 (O_240,N_2371,N_2560);
nand UO_241 (O_241,N_2255,N_2680);
nor UO_242 (O_242,N_2541,N_2720);
or UO_243 (O_243,N_2667,N_2396);
nor UO_244 (O_244,N_2271,N_2455);
nand UO_245 (O_245,N_2728,N_2820);
and UO_246 (O_246,N_2330,N_2977);
and UO_247 (O_247,N_2954,N_2454);
or UO_248 (O_248,N_2618,N_2931);
and UO_249 (O_249,N_2701,N_2295);
or UO_250 (O_250,N_2603,N_2291);
nor UO_251 (O_251,N_2591,N_2578);
or UO_252 (O_252,N_2347,N_2872);
or UO_253 (O_253,N_2423,N_2906);
nand UO_254 (O_254,N_2646,N_2871);
xor UO_255 (O_255,N_2832,N_2350);
and UO_256 (O_256,N_2474,N_2551);
nand UO_257 (O_257,N_2709,N_2599);
nor UO_258 (O_258,N_2483,N_2957);
and UO_259 (O_259,N_2391,N_2750);
and UO_260 (O_260,N_2415,N_2290);
nand UO_261 (O_261,N_2741,N_2663);
or UO_262 (O_262,N_2593,N_2782);
or UO_263 (O_263,N_2562,N_2382);
nand UO_264 (O_264,N_2684,N_2538);
xor UO_265 (O_265,N_2552,N_2883);
nand UO_266 (O_266,N_2723,N_2548);
nor UO_267 (O_267,N_2787,N_2637);
or UO_268 (O_268,N_2269,N_2805);
or UO_269 (O_269,N_2619,N_2315);
and UO_270 (O_270,N_2319,N_2656);
xor UO_271 (O_271,N_2301,N_2449);
or UO_272 (O_272,N_2434,N_2732);
or UO_273 (O_273,N_2532,N_2968);
xnor UO_274 (O_274,N_2973,N_2796);
nor UO_275 (O_275,N_2392,N_2477);
or UO_276 (O_276,N_2274,N_2708);
nand UO_277 (O_277,N_2488,N_2286);
nand UO_278 (O_278,N_2534,N_2987);
nand UO_279 (O_279,N_2845,N_2622);
and UO_280 (O_280,N_2304,N_2813);
xnor UO_281 (O_281,N_2617,N_2991);
or UO_282 (O_282,N_2543,N_2659);
or UO_283 (O_283,N_2783,N_2440);
nand UO_284 (O_284,N_2495,N_2283);
and UO_285 (O_285,N_2308,N_2427);
or UO_286 (O_286,N_2265,N_2450);
nor UO_287 (O_287,N_2824,N_2398);
or UO_288 (O_288,N_2917,N_2956);
nor UO_289 (O_289,N_2393,N_2837);
and UO_290 (O_290,N_2819,N_2282);
and UO_291 (O_291,N_2675,N_2657);
nand UO_292 (O_292,N_2252,N_2516);
and UO_293 (O_293,N_2800,N_2465);
nor UO_294 (O_294,N_2795,N_2857);
and UO_295 (O_295,N_2864,N_2531);
and UO_296 (O_296,N_2913,N_2966);
and UO_297 (O_297,N_2862,N_2281);
nand UO_298 (O_298,N_2397,N_2848);
nand UO_299 (O_299,N_2375,N_2673);
or UO_300 (O_300,N_2641,N_2786);
nor UO_301 (O_301,N_2961,N_2614);
xnor UO_302 (O_302,N_2407,N_2722);
nor UO_303 (O_303,N_2901,N_2300);
and UO_304 (O_304,N_2565,N_2972);
and UO_305 (O_305,N_2905,N_2566);
and UO_306 (O_306,N_2768,N_2894);
nand UO_307 (O_307,N_2412,N_2336);
xor UO_308 (O_308,N_2971,N_2340);
nand UO_309 (O_309,N_2688,N_2502);
or UO_310 (O_310,N_2491,N_2479);
or UO_311 (O_311,N_2807,N_2650);
or UO_312 (O_312,N_2376,N_2702);
and UO_313 (O_313,N_2735,N_2921);
and UO_314 (O_314,N_2772,N_2756);
and UO_315 (O_315,N_2533,N_2810);
or UO_316 (O_316,N_2417,N_2585);
or UO_317 (O_317,N_2432,N_2816);
and UO_318 (O_318,N_2326,N_2257);
and UO_319 (O_319,N_2715,N_2854);
nand UO_320 (O_320,N_2830,N_2610);
or UO_321 (O_321,N_2978,N_2511);
or UO_322 (O_322,N_2717,N_2840);
xnor UO_323 (O_323,N_2537,N_2892);
or UO_324 (O_324,N_2933,N_2456);
or UO_325 (O_325,N_2555,N_2880);
or UO_326 (O_326,N_2368,N_2482);
nor UO_327 (O_327,N_2386,N_2337);
or UO_328 (O_328,N_2475,N_2716);
nand UO_329 (O_329,N_2727,N_2258);
xnor UO_330 (O_330,N_2346,N_2890);
nand UO_331 (O_331,N_2658,N_2334);
or UO_332 (O_332,N_2446,N_2636);
nor UO_333 (O_333,N_2509,N_2395);
xor UO_334 (O_334,N_2329,N_2280);
nor UO_335 (O_335,N_2251,N_2615);
nor UO_336 (O_336,N_2299,N_2522);
nand UO_337 (O_337,N_2760,N_2584);
nor UO_338 (O_338,N_2327,N_2556);
or UO_339 (O_339,N_2459,N_2524);
nor UO_340 (O_340,N_2390,N_2852);
nand UO_341 (O_341,N_2275,N_2940);
and UO_342 (O_342,N_2367,N_2829);
nor UO_343 (O_343,N_2679,N_2965);
or UO_344 (O_344,N_2950,N_2643);
nand UO_345 (O_345,N_2953,N_2766);
or UO_346 (O_346,N_2629,N_2693);
nand UO_347 (O_347,N_2250,N_2559);
or UO_348 (O_348,N_2564,N_2817);
nand UO_349 (O_349,N_2424,N_2765);
xnor UO_350 (O_350,N_2419,N_2360);
xor UO_351 (O_351,N_2843,N_2849);
or UO_352 (O_352,N_2431,N_2942);
or UO_353 (O_353,N_2557,N_2487);
nand UO_354 (O_354,N_2582,N_2510);
or UO_355 (O_355,N_2726,N_2863);
nand UO_356 (O_356,N_2771,N_2605);
or UO_357 (O_357,N_2888,N_2408);
xor UO_358 (O_358,N_2855,N_2604);
and UO_359 (O_359,N_2535,N_2553);
or UO_360 (O_360,N_2592,N_2600);
and UO_361 (O_361,N_2907,N_2507);
nand UO_362 (O_362,N_2445,N_2690);
or UO_363 (O_363,N_2777,N_2651);
nand UO_364 (O_364,N_2437,N_2661);
and UO_365 (O_365,N_2400,N_2546);
nor UO_366 (O_366,N_2567,N_2381);
and UO_367 (O_367,N_2421,N_2844);
and UO_368 (O_368,N_2743,N_2504);
or UO_369 (O_369,N_2372,N_2558);
or UO_370 (O_370,N_2785,N_2353);
nand UO_371 (O_371,N_2929,N_2458);
nand UO_372 (O_372,N_2878,N_2361);
and UO_373 (O_373,N_2790,N_2920);
nand UO_374 (O_374,N_2260,N_2335);
nand UO_375 (O_375,N_2820,N_2751);
nand UO_376 (O_376,N_2658,N_2438);
nor UO_377 (O_377,N_2936,N_2790);
nor UO_378 (O_378,N_2533,N_2775);
and UO_379 (O_379,N_2530,N_2814);
nand UO_380 (O_380,N_2824,N_2337);
and UO_381 (O_381,N_2517,N_2469);
nor UO_382 (O_382,N_2759,N_2351);
nand UO_383 (O_383,N_2514,N_2971);
nor UO_384 (O_384,N_2601,N_2731);
xnor UO_385 (O_385,N_2418,N_2622);
nor UO_386 (O_386,N_2447,N_2322);
and UO_387 (O_387,N_2262,N_2801);
or UO_388 (O_388,N_2543,N_2457);
nand UO_389 (O_389,N_2428,N_2650);
and UO_390 (O_390,N_2452,N_2909);
nand UO_391 (O_391,N_2664,N_2866);
or UO_392 (O_392,N_2682,N_2386);
and UO_393 (O_393,N_2555,N_2702);
or UO_394 (O_394,N_2609,N_2826);
nand UO_395 (O_395,N_2325,N_2391);
nor UO_396 (O_396,N_2954,N_2792);
nor UO_397 (O_397,N_2292,N_2329);
or UO_398 (O_398,N_2792,N_2541);
nand UO_399 (O_399,N_2549,N_2798);
nor UO_400 (O_400,N_2750,N_2442);
or UO_401 (O_401,N_2847,N_2302);
and UO_402 (O_402,N_2562,N_2832);
xor UO_403 (O_403,N_2624,N_2425);
nor UO_404 (O_404,N_2727,N_2559);
or UO_405 (O_405,N_2722,N_2342);
and UO_406 (O_406,N_2866,N_2800);
and UO_407 (O_407,N_2678,N_2908);
and UO_408 (O_408,N_2651,N_2343);
nand UO_409 (O_409,N_2696,N_2370);
and UO_410 (O_410,N_2672,N_2401);
or UO_411 (O_411,N_2973,N_2733);
or UO_412 (O_412,N_2361,N_2987);
or UO_413 (O_413,N_2621,N_2332);
and UO_414 (O_414,N_2736,N_2695);
or UO_415 (O_415,N_2790,N_2682);
nand UO_416 (O_416,N_2817,N_2472);
nand UO_417 (O_417,N_2851,N_2922);
nor UO_418 (O_418,N_2567,N_2862);
xor UO_419 (O_419,N_2436,N_2292);
nand UO_420 (O_420,N_2392,N_2628);
nor UO_421 (O_421,N_2397,N_2527);
and UO_422 (O_422,N_2594,N_2684);
xor UO_423 (O_423,N_2982,N_2710);
nor UO_424 (O_424,N_2333,N_2505);
nand UO_425 (O_425,N_2802,N_2672);
and UO_426 (O_426,N_2718,N_2361);
and UO_427 (O_427,N_2771,N_2665);
nor UO_428 (O_428,N_2626,N_2457);
nand UO_429 (O_429,N_2380,N_2313);
and UO_430 (O_430,N_2372,N_2506);
nor UO_431 (O_431,N_2471,N_2739);
xor UO_432 (O_432,N_2564,N_2313);
or UO_433 (O_433,N_2515,N_2594);
nand UO_434 (O_434,N_2333,N_2769);
and UO_435 (O_435,N_2937,N_2391);
nor UO_436 (O_436,N_2311,N_2511);
nor UO_437 (O_437,N_2528,N_2804);
xnor UO_438 (O_438,N_2536,N_2260);
and UO_439 (O_439,N_2263,N_2386);
and UO_440 (O_440,N_2381,N_2470);
or UO_441 (O_441,N_2862,N_2409);
nor UO_442 (O_442,N_2371,N_2782);
or UO_443 (O_443,N_2294,N_2869);
nand UO_444 (O_444,N_2423,N_2400);
and UO_445 (O_445,N_2458,N_2452);
nor UO_446 (O_446,N_2822,N_2967);
nand UO_447 (O_447,N_2608,N_2712);
xnor UO_448 (O_448,N_2295,N_2927);
and UO_449 (O_449,N_2439,N_2822);
xor UO_450 (O_450,N_2531,N_2458);
nor UO_451 (O_451,N_2937,N_2353);
xnor UO_452 (O_452,N_2743,N_2334);
nand UO_453 (O_453,N_2978,N_2593);
xnor UO_454 (O_454,N_2980,N_2372);
nand UO_455 (O_455,N_2520,N_2811);
and UO_456 (O_456,N_2844,N_2457);
or UO_457 (O_457,N_2588,N_2681);
or UO_458 (O_458,N_2509,N_2625);
nand UO_459 (O_459,N_2376,N_2288);
and UO_460 (O_460,N_2258,N_2778);
and UO_461 (O_461,N_2637,N_2731);
and UO_462 (O_462,N_2362,N_2865);
or UO_463 (O_463,N_2945,N_2709);
nor UO_464 (O_464,N_2346,N_2306);
and UO_465 (O_465,N_2921,N_2948);
xor UO_466 (O_466,N_2669,N_2755);
nor UO_467 (O_467,N_2836,N_2982);
nor UO_468 (O_468,N_2596,N_2253);
nor UO_469 (O_469,N_2735,N_2641);
nand UO_470 (O_470,N_2854,N_2837);
or UO_471 (O_471,N_2786,N_2624);
and UO_472 (O_472,N_2281,N_2352);
nor UO_473 (O_473,N_2433,N_2460);
nand UO_474 (O_474,N_2883,N_2418);
nor UO_475 (O_475,N_2294,N_2795);
and UO_476 (O_476,N_2362,N_2547);
nand UO_477 (O_477,N_2789,N_2925);
nand UO_478 (O_478,N_2791,N_2767);
and UO_479 (O_479,N_2256,N_2568);
or UO_480 (O_480,N_2814,N_2416);
nand UO_481 (O_481,N_2443,N_2711);
nand UO_482 (O_482,N_2399,N_2410);
and UO_483 (O_483,N_2629,N_2399);
nor UO_484 (O_484,N_2439,N_2909);
or UO_485 (O_485,N_2810,N_2672);
or UO_486 (O_486,N_2363,N_2827);
nor UO_487 (O_487,N_2846,N_2490);
and UO_488 (O_488,N_2693,N_2440);
and UO_489 (O_489,N_2259,N_2484);
xnor UO_490 (O_490,N_2513,N_2711);
and UO_491 (O_491,N_2367,N_2304);
or UO_492 (O_492,N_2713,N_2506);
nand UO_493 (O_493,N_2453,N_2310);
xnor UO_494 (O_494,N_2418,N_2470);
and UO_495 (O_495,N_2389,N_2686);
nand UO_496 (O_496,N_2798,N_2880);
and UO_497 (O_497,N_2733,N_2644);
or UO_498 (O_498,N_2654,N_2657);
nor UO_499 (O_499,N_2369,N_2600);
endmodule